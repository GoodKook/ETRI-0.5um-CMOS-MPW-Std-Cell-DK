magic
tech scmos
timestamp 1719894731
<< checkpaint >>
rect 7 781 80 855
rect 7 680 80 781
rect 7 659 80 680
rect 6 353 80 659
rect 8 -20 79 280
<< nwell >>
rect 0 700 60 761
rect 0 373 60 639
<< psubstratepdiff >>
rect 4 780 55 835
rect 4 0 55 260
<< nsubstratendiff >>
rect 4 703 55 758
rect 4 376 55 636
<< genericcontact >>
rect 8 821 10 823
rect 18 821 20 823
rect 32 821 34 823
rect 43 821 45 823
rect 8 810 10 812
rect 18 810 20 812
rect 32 810 34 812
rect 43 810 45 812
rect 8 799 10 801
rect 18 799 20 801
rect 32 799 34 801
rect 43 799 45 801
rect 8 789 10 791
rect 18 789 20 791
rect 32 789 34 791
rect 43 789 45 791
rect 8 741 10 743
rect 18 741 20 743
rect 32 741 34 743
rect 43 741 45 743
rect 8 731 10 733
rect 18 731 20 733
rect 32 731 34 733
rect 43 731 45 733
rect 8 720 10 722
rect 18 720 20 722
rect 32 720 34 722
rect 43 720 45 722
rect 8 709 10 711
rect 18 709 20 711
rect 32 709 34 711
rect 43 709 45 711
rect 8 627 10 629
rect 18 627 20 629
rect 32 627 34 629
rect 43 627 45 629
rect 8 617 10 619
rect 18 617 20 619
rect 32 617 34 619
rect 43 617 45 619
rect 8 606 10 608
rect 18 606 20 608
rect 32 606 34 608
rect 43 606 45 608
rect 8 595 10 597
rect 18 595 20 597
rect 32 595 34 597
rect 43 595 45 597
rect 8 585 10 587
rect 18 585 20 587
rect 32 585 34 587
rect 43 585 45 587
rect 8 574 10 576
rect 18 574 20 576
rect 32 574 34 576
rect 43 574 45 576
rect 8 563 10 565
rect 18 563 20 565
rect 32 563 34 565
rect 43 563 45 565
rect 8 553 10 555
rect 18 553 20 555
rect 32 553 34 555
rect 43 553 45 555
rect 8 542 10 544
rect 18 542 20 544
rect 32 542 34 544
rect 43 542 45 544
rect 8 531 10 533
rect 18 531 20 533
rect 32 531 34 533
rect 43 531 45 533
rect 8 521 10 523
rect 18 521 20 523
rect 32 521 34 523
rect 43 521 45 523
rect 8 510 10 512
rect 18 510 20 512
rect 32 510 34 512
rect 43 510 45 512
rect 8 499 10 501
rect 18 499 20 501
rect 32 499 34 501
rect 43 499 45 501
rect 8 489 10 491
rect 18 489 20 491
rect 32 489 34 491
rect 43 489 45 491
rect 8 478 10 480
rect 18 478 20 480
rect 32 478 34 480
rect 43 478 45 480
rect 8 467 10 469
rect 18 467 20 469
rect 32 467 34 469
rect 43 467 45 469
rect 8 457 10 459
rect 18 457 20 459
rect 32 457 34 459
rect 43 457 45 459
rect 8 446 10 448
rect 18 446 20 448
rect 32 446 34 448
rect 43 446 45 448
rect 8 435 10 437
rect 18 435 20 437
rect 32 435 34 437
rect 43 435 45 437
rect 8 425 10 427
rect 18 425 20 427
rect 32 425 34 427
rect 43 425 45 427
rect 8 414 10 416
rect 18 414 20 416
rect 32 414 34 416
rect 43 414 45 416
rect 8 403 10 405
rect 18 403 20 405
rect 32 403 34 405
rect 43 403 45 405
rect 8 393 10 395
rect 18 393 20 395
rect 32 393 34 395
rect 43 393 45 395
rect 8 382 10 384
rect 18 382 20 384
rect 32 382 34 384
rect 43 382 45 384
rect 9 248 11 250
rect 19 248 21 250
rect 33 248 35 250
rect 44 248 46 250
rect 9 237 11 239
rect 19 237 21 239
rect 33 237 35 239
rect 44 237 46 239
rect 9 226 11 228
rect 19 226 21 228
rect 33 226 35 228
rect 44 226 46 228
rect 9 216 11 218
rect 19 216 21 218
rect 33 216 35 218
rect 44 216 46 218
rect 9 205 11 207
rect 19 205 21 207
rect 33 205 35 207
rect 44 205 46 207
rect 9 194 11 196
rect 19 194 21 196
rect 33 194 35 196
rect 44 194 46 196
rect 9 184 11 186
rect 19 184 21 186
rect 33 184 35 186
rect 44 184 46 186
rect 9 173 11 175
rect 19 173 21 175
rect 33 173 35 175
rect 44 173 46 175
rect 9 162 11 164
rect 19 162 21 164
rect 33 162 35 164
rect 44 162 46 164
rect 9 152 11 154
rect 19 152 21 154
rect 33 152 35 154
rect 44 152 46 154
rect 9 141 11 143
rect 19 141 21 143
rect 33 141 35 143
rect 44 141 46 143
rect 9 130 11 132
rect 19 130 21 132
rect 33 130 35 132
rect 44 130 46 132
rect 9 120 11 122
rect 19 120 21 122
rect 33 120 35 122
rect 44 120 46 122
rect 9 109 11 111
rect 19 109 21 111
rect 33 109 35 111
rect 44 109 46 111
rect 9 98 11 100
rect 19 98 21 100
rect 33 98 35 100
rect 44 98 46 100
rect 9 88 11 90
rect 19 88 21 90
rect 33 88 35 90
rect 44 88 46 90
rect 9 77 11 79
rect 19 77 21 79
rect 33 77 35 79
rect 44 77 46 79
rect 9 66 11 68
rect 19 66 21 68
rect 33 66 35 68
rect 44 66 46 68
rect 9 56 11 58
rect 19 56 21 58
rect 33 56 35 58
rect 44 56 46 58
rect 9 45 11 47
rect 19 45 21 47
rect 33 45 35 47
rect 44 45 46 47
rect 9 34 11 36
rect 19 34 21 36
rect 33 34 35 36
rect 44 34 46 36
rect 9 24 11 26
rect 19 24 21 26
rect 33 24 35 26
rect 44 24 46 26
rect 9 13 11 15
rect 19 13 21 15
rect 33 13 35 15
rect 44 13 46 15
rect 9 2 11 4
rect 19 2 21 4
rect 33 2 35 4
rect 44 2 46 4
<< metal1 >>
rect 1 780 59 835
rect 1 703 59 758
rect 1 376 59 636
rect 1 0 59 260
<< metal2 >>
rect 1 780 59 835
rect 1 703 59 758
rect 1 376 59 636
rect 1 0 59 260
<< gv1 >>
rect 13 815 15 818
rect 23 815 26 818
rect 37 815 40 818
rect 48 815 51 818
rect 13 804 15 807
rect 23 804 26 807
rect 37 804 40 807
rect 48 804 51 807
rect 13 794 15 796
rect 23 794 26 796
rect 37 794 40 796
rect 48 794 51 796
rect 13 736 15 738
rect 23 736 26 738
rect 37 736 40 738
rect 48 736 51 738
rect 13 725 15 728
rect 23 725 26 728
rect 37 725 40 728
rect 48 725 51 728
rect 13 714 15 717
rect 23 714 26 717
rect 37 714 40 717
rect 48 714 51 717
rect 13 622 15 624
rect 23 622 26 624
rect 37 622 40 624
rect 48 622 51 624
rect 13 611 15 614
rect 23 611 26 614
rect 37 611 40 614
rect 48 611 51 614
rect 13 600 15 603
rect 23 600 26 603
rect 37 600 40 603
rect 48 600 51 603
rect 13 590 15 592
rect 23 590 26 592
rect 37 590 40 592
rect 48 590 51 592
rect 13 579 15 582
rect 23 579 26 582
rect 37 579 40 582
rect 48 579 51 582
rect 13 568 15 571
rect 23 568 26 571
rect 37 568 40 571
rect 48 568 51 571
rect 13 558 15 560
rect 23 558 26 560
rect 37 558 40 560
rect 48 558 51 560
rect 13 547 15 550
rect 23 547 26 550
rect 37 547 40 550
rect 48 547 51 550
rect 13 536 15 539
rect 23 536 26 539
rect 37 536 40 539
rect 48 536 51 539
rect 13 526 15 528
rect 23 526 26 528
rect 37 526 40 528
rect 48 526 51 528
rect 13 515 15 518
rect 23 515 26 518
rect 37 515 40 518
rect 48 515 51 518
rect 13 504 15 507
rect 23 504 26 507
rect 37 504 40 507
rect 48 504 51 507
rect 13 494 15 496
rect 23 494 26 496
rect 37 494 40 496
rect 48 494 51 496
rect 13 483 15 486
rect 23 483 26 486
rect 37 483 40 486
rect 48 483 51 486
rect 13 472 15 475
rect 23 472 26 475
rect 37 472 40 475
rect 48 472 51 475
rect 13 462 15 464
rect 23 462 26 464
rect 37 462 40 464
rect 48 462 51 464
rect 13 451 15 454
rect 23 451 26 454
rect 37 451 40 454
rect 48 451 51 454
rect 13 440 15 443
rect 23 440 26 443
rect 37 440 40 443
rect 48 440 51 443
rect 13 430 15 432
rect 23 430 26 432
rect 37 430 40 432
rect 48 430 51 432
rect 13 419 15 422
rect 23 419 26 422
rect 37 419 40 422
rect 48 419 51 422
rect 13 408 15 411
rect 23 408 26 411
rect 37 408 40 411
rect 48 408 51 411
rect 13 398 15 400
rect 23 398 26 400
rect 37 398 40 400
rect 48 398 51 400
rect 13 387 15 390
rect 23 387 26 390
rect 37 387 40 390
rect 48 387 51 390
rect 14 242 16 245
rect 24 242 27 245
rect 38 242 41 245
rect 49 242 52 245
rect 14 231 16 234
rect 24 231 27 234
rect 38 231 41 234
rect 49 231 52 234
rect 14 221 16 223
rect 24 221 27 223
rect 38 221 41 223
rect 49 221 52 223
rect 14 210 16 213
rect 24 210 27 213
rect 38 210 41 213
rect 49 210 52 213
rect 14 199 16 202
rect 24 199 27 202
rect 38 199 41 202
rect 49 199 52 202
rect 14 189 16 191
rect 24 189 27 191
rect 38 189 41 191
rect 49 189 52 191
rect 14 178 16 181
rect 24 178 27 181
rect 38 178 41 181
rect 49 178 52 181
rect 14 167 16 170
rect 24 167 27 170
rect 38 167 41 170
rect 49 167 52 170
rect 14 157 16 159
rect 24 157 27 159
rect 38 157 41 159
rect 49 157 52 159
rect 14 146 16 149
rect 24 146 27 149
rect 38 146 41 149
rect 49 146 52 149
rect 14 135 16 138
rect 24 135 27 138
rect 38 135 41 138
rect 49 135 52 138
rect 14 125 16 127
rect 24 125 27 127
rect 38 125 41 127
rect 49 125 52 127
rect 14 114 16 117
rect 24 114 27 117
rect 38 114 41 117
rect 49 114 52 117
rect 14 103 16 106
rect 24 103 27 106
rect 38 103 41 106
rect 49 103 52 106
rect 14 93 16 95
rect 24 93 27 95
rect 38 93 41 95
rect 49 93 52 95
rect 14 82 16 85
rect 24 82 27 85
rect 38 82 41 85
rect 49 82 52 85
rect 14 71 16 74
rect 24 71 27 74
rect 38 71 41 74
rect 49 71 52 74
rect 14 61 16 63
rect 24 61 27 63
rect 38 61 41 63
rect 49 61 52 63
rect 14 50 16 53
rect 24 50 27 53
rect 38 50 41 53
rect 49 50 52 53
rect 14 39 16 42
rect 24 39 27 42
rect 38 39 41 42
rect 49 39 52 42
rect 14 29 16 31
rect 24 29 27 31
rect 38 29 41 31
rect 49 29 52 31
rect 14 18 16 21
rect 24 18 27 21
rect 38 18 41 21
rect 49 18 52 21
rect 14 7 16 10
rect 24 7 27 10
rect 38 7 41 10
rect 49 7 52 10
<< metal3 >>
rect 1 780 59 835
rect 1 703 59 758
rect 1 376 59 636
rect 1 0 59 260
<< gv2 >>
rect 7 820 10 823
rect 18 820 21 823
rect 32 820 35 823
rect 43 820 45 823
rect 7 810 10 812
rect 18 810 21 812
rect 32 810 35 812
rect 43 810 45 812
rect 7 799 10 802
rect 18 799 21 802
rect 32 799 35 802
rect 43 799 45 802
rect 7 788 10 791
rect 18 788 21 791
rect 32 788 35 791
rect 43 788 45 791
rect 7 741 10 744
rect 18 741 21 744
rect 32 741 35 744
rect 43 741 45 744
rect 7 730 10 733
rect 18 730 21 733
rect 32 730 35 733
rect 43 730 45 733
rect 7 720 10 722
rect 18 720 21 722
rect 32 720 35 722
rect 43 720 45 722
rect 7 709 10 712
rect 18 709 21 712
rect 32 709 35 712
rect 43 709 45 712
rect 7 627 10 630
rect 18 627 21 630
rect 32 627 35 630
rect 43 627 45 630
rect 7 616 10 619
rect 18 616 21 619
rect 32 616 35 619
rect 43 616 45 619
rect 7 606 10 608
rect 18 606 21 608
rect 32 606 35 608
rect 43 606 45 608
rect 7 595 10 598
rect 18 595 21 598
rect 32 595 35 598
rect 43 595 45 598
rect 7 584 10 587
rect 18 584 21 587
rect 32 584 35 587
rect 43 584 45 587
rect 7 574 10 576
rect 18 574 21 576
rect 32 574 35 576
rect 43 574 45 576
rect 7 563 10 566
rect 18 563 21 566
rect 32 563 35 566
rect 43 563 45 566
rect 7 552 10 555
rect 18 552 21 555
rect 32 552 35 555
rect 43 552 45 555
rect 7 542 10 544
rect 18 542 21 544
rect 32 542 35 544
rect 43 542 45 544
rect 7 531 10 534
rect 18 531 21 534
rect 32 531 35 534
rect 43 531 45 534
rect 7 520 10 523
rect 18 520 21 523
rect 32 520 35 523
rect 43 520 45 523
rect 7 510 10 512
rect 18 510 21 512
rect 32 510 35 512
rect 43 510 45 512
rect 7 499 10 502
rect 18 499 21 502
rect 32 499 35 502
rect 43 499 45 502
rect 7 488 10 491
rect 18 488 21 491
rect 32 488 35 491
rect 43 488 45 491
rect 7 478 10 480
rect 18 478 21 480
rect 32 478 35 480
rect 43 478 45 480
rect 7 467 10 470
rect 18 467 21 470
rect 32 467 35 470
rect 43 467 45 470
rect 7 456 10 459
rect 18 456 21 459
rect 32 456 35 459
rect 43 456 45 459
rect 7 446 10 448
rect 18 446 21 448
rect 32 446 35 448
rect 43 446 45 448
rect 7 435 10 438
rect 18 435 21 438
rect 32 435 35 438
rect 43 435 45 438
rect 7 424 10 427
rect 18 424 21 427
rect 32 424 35 427
rect 43 424 45 427
rect 7 414 10 416
rect 18 414 21 416
rect 32 414 35 416
rect 43 414 45 416
rect 7 403 10 406
rect 18 403 21 406
rect 32 403 35 406
rect 43 403 45 406
rect 7 392 10 395
rect 18 392 21 395
rect 32 392 35 395
rect 43 392 45 395
rect 7 382 10 384
rect 18 382 21 384
rect 32 382 35 384
rect 43 382 45 384
rect 8 247 11 250
rect 19 247 22 250
rect 33 247 36 250
rect 44 247 46 250
rect 8 237 11 239
rect 19 237 22 239
rect 33 237 36 239
rect 44 237 46 239
rect 8 226 11 229
rect 19 226 22 229
rect 33 226 36 229
rect 44 226 46 229
rect 8 215 11 218
rect 19 215 22 218
rect 33 215 36 218
rect 44 215 46 218
rect 8 205 11 207
rect 19 205 22 207
rect 33 205 36 207
rect 44 205 46 207
rect 8 194 11 197
rect 19 194 22 197
rect 33 194 36 197
rect 44 194 46 197
rect 8 183 11 186
rect 19 183 22 186
rect 33 183 36 186
rect 44 183 46 186
rect 8 173 11 175
rect 19 173 22 175
rect 33 173 36 175
rect 44 173 46 175
rect 8 162 11 165
rect 19 162 22 165
rect 33 162 36 165
rect 44 162 46 165
rect 8 151 11 154
rect 19 151 22 154
rect 33 151 36 154
rect 44 151 46 154
rect 8 141 11 143
rect 19 141 22 143
rect 33 141 36 143
rect 44 141 46 143
rect 8 130 11 133
rect 19 130 22 133
rect 33 130 36 133
rect 44 130 46 133
rect 8 119 11 122
rect 19 119 22 122
rect 33 119 36 122
rect 44 119 46 122
rect 8 109 11 111
rect 19 109 22 111
rect 33 109 36 111
rect 44 109 46 111
rect 8 98 11 101
rect 19 98 22 101
rect 33 98 36 101
rect 44 98 46 101
rect 8 87 11 90
rect 19 87 22 90
rect 33 87 36 90
rect 44 87 46 90
rect 8 77 11 79
rect 19 77 22 79
rect 33 77 36 79
rect 44 77 46 79
rect 8 66 11 69
rect 19 66 22 69
rect 33 66 36 69
rect 44 66 46 69
rect 8 55 11 58
rect 19 55 22 58
rect 33 55 36 58
rect 44 55 46 58
rect 8 45 11 47
rect 19 45 22 47
rect 33 45 36 47
rect 44 45 46 47
rect 8 34 11 37
rect 19 34 22 37
rect 33 34 36 37
rect 44 34 46 37
rect 8 23 11 26
rect 19 23 22 26
rect 33 23 36 26
rect 44 23 46 26
rect 8 13 11 15
rect 19 13 22 15
rect 33 13 36 15
rect 44 13 46 15
rect 8 2 11 5
rect 19 2 22 5
rect 33 2 36 5
rect 44 2 46 5
<< end >>
