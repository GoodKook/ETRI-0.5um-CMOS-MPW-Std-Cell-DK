magic
tech scmos
magscale 1 2
timestamp 1727572430
<< nwell >>
rect -12 154 192 272
<< ntransistor >>
rect 40 14 44 34
rect 60 14 64 34
rect 80 14 84 34
<< ptransistor >>
rect 20 186 24 246
rect 40 186 44 246
rect 60 186 64 246
rect 80 186 84 246
rect 124 178 128 238
rect 144 178 148 238
<< ndiffusion >>
rect 38 14 40 34
rect 44 14 46 34
rect 58 14 60 34
rect 64 14 66 34
rect 78 14 80 34
rect 84 14 86 34
<< pdiffusion >>
rect 18 186 20 246
rect 24 186 26 246
rect 38 186 40 246
rect 44 186 46 246
rect 58 186 60 246
rect 64 234 80 246
rect 64 186 66 234
rect 78 186 80 234
rect 84 188 86 246
rect 84 186 98 188
rect 122 178 124 238
rect 128 234 144 238
rect 128 182 130 234
rect 142 182 144 234
rect 128 178 144 182
rect 148 178 150 238
<< ndcontact >>
rect 24 14 38 34
rect 46 14 58 34
rect 66 14 78 34
rect 86 14 98 34
<< pdcontact >>
rect 6 186 18 246
rect 26 186 38 246
rect 46 186 58 246
rect 66 186 78 234
rect 86 188 98 246
rect 110 178 122 238
rect 130 182 142 234
rect 150 178 162 238
<< psubstratepcontact >>
rect -6 -6 186 6
<< nsubstratencontact >>
rect -6 254 186 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 60 246 64 250
rect 80 246 84 250
rect 124 238 128 242
rect 144 238 148 242
rect 20 182 24 186
rect 40 182 44 186
rect 20 178 44 182
rect 40 128 44 178
rect 36 116 44 128
rect 40 34 44 116
rect 60 182 64 186
rect 80 182 84 186
rect 60 178 84 182
rect 60 34 64 178
rect 124 170 128 178
rect 144 170 148 178
rect 98 166 148 170
rect 98 128 104 166
rect 96 116 104 128
rect 98 56 104 116
rect 80 50 104 56
rect 80 34 84 50
rect 40 10 44 14
rect 60 10 64 14
rect 80 10 84 14
<< polycontact >>
rect 24 116 36 128
rect 64 110 76 122
rect 84 116 96 128
<< metal1 >>
rect -6 266 186 268
rect -6 252 186 254
rect 26 246 38 252
rect 58 240 86 246
rect 6 180 18 186
rect 46 180 58 186
rect 6 174 58 180
rect 110 240 162 246
rect 110 238 122 240
rect 66 182 78 186
rect 66 178 110 182
rect 150 238 162 240
rect 66 176 122 178
rect 130 166 138 182
rect 115 158 138 166
rect 115 46 123 158
rect 51 40 123 46
rect 51 34 58 40
rect 91 34 98 40
rect 24 8 38 14
rect 66 8 78 14
rect -6 6 186 8
rect -6 -8 186 -6
<< m2contact >>
rect 63 122 77 136
rect 23 102 37 116
rect 83 102 97 116
rect 123 102 137 116
<< metal2 >>
rect 63 136 77 156
rect 123 116 137 136
rect 23 82 37 102
rect 83 82 97 102
<< m2p >>
rect 63 142 77 156
rect 123 122 137 136
rect 23 82 37 96
rect 83 82 97 96
<< labels >>
rlabel metal2 23 82 37 96 0 A
port 0 nsew signal input
rlabel metal2 63 142 77 156 0 B
port 1 nsew signal input
rlabel metal2 83 82 97 96 0 C
port 2 nsew signal input
rlabel metal2 123 122 137 136 0 Y
port 3 nsew signal output
rlabel metal1 -6 252 186 268 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 -6 -8 186 8 0 gnd
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 180 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
