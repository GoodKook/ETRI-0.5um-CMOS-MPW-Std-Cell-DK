magic
tech scmos
magscale 1 3
timestamp 1554524574
<< checkpaint >>
rect -52 -52 1092 88
<< pseudo_rpoly2 >>
rect 8 8 1032 28
use poly2cont_CDNS_7230122529125  poly2cont_CDNS_7230122529125_0
timestamp 1554524574
transform 1 0 1014 0 1 8
box 0 0 18 20
use poly2cont_CDNS_7230122529125  poly2cont_CDNS_7230122529125_1
timestamp 1554524574
transform 1 0 8 0 1 8
box 0 0 18 20
<< end >>
