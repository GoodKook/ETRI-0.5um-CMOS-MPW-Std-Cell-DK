magic
tech scmos
magscale 1 6
timestamp 1726646557
<< checkpaint >>
rect 8700 8700 29300 29300
<< metal1 >>
rect 8840 27133 10240 27160
rect 8840 27115 8855 27133
rect 8873 27115 8891 27133
rect 8909 27115 8927 27133
rect 8945 27115 8963 27133
rect 8981 27115 8999 27133
rect 9017 27115 9035 27133
rect 9053 27115 9071 27133
rect 9089 27115 9107 27133
rect 9125 27115 10240 27133
rect 8840 27097 10240 27115
rect 8840 27079 8855 27097
rect 8873 27079 8891 27097
rect 8909 27079 8927 27097
rect 8945 27079 8963 27097
rect 8981 27079 8999 27097
rect 9017 27079 9035 27097
rect 9053 27079 9071 27097
rect 9089 27079 9107 27097
rect 9125 27079 10240 27097
rect 8840 27061 10240 27079
rect 8840 27043 8855 27061
rect 8873 27043 8891 27061
rect 8909 27043 8927 27061
rect 8945 27043 8963 27061
rect 8981 27043 8999 27061
rect 9017 27043 9035 27061
rect 9053 27043 9071 27061
rect 9089 27043 9107 27061
rect 9125 27043 10240 27061
rect 8840 27025 10240 27043
rect 8840 27007 8855 27025
rect 8873 27007 8891 27025
rect 8909 27007 8927 27025
rect 8945 27007 8963 27025
rect 8981 27007 8999 27025
rect 9017 27007 9035 27025
rect 9053 27007 9071 27025
rect 9089 27007 9107 27025
rect 9125 27007 10240 27025
rect 8840 26989 10240 27007
rect 8840 26971 8855 26989
rect 8873 26971 8891 26989
rect 8909 26971 8927 26989
rect 8945 26971 8963 26989
rect 8981 26971 8999 26989
rect 9017 26971 9035 26989
rect 9053 26971 9071 26989
rect 9089 26971 9107 26989
rect 9125 26971 10240 26989
rect 8840 26953 10240 26971
rect 8840 26935 8855 26953
rect 8873 26935 8891 26953
rect 8909 26935 8927 26953
rect 8945 26935 8963 26953
rect 8981 26935 8999 26953
rect 9017 26935 9035 26953
rect 9053 26935 9071 26953
rect 9089 26935 9107 26953
rect 9125 26935 10240 26953
rect 8840 26917 10240 26935
rect 8840 26899 8855 26917
rect 8873 26899 8891 26917
rect 8909 26899 8927 26917
rect 8945 26899 8963 26917
rect 8981 26899 8999 26917
rect 9017 26899 9035 26917
rect 9053 26899 9071 26917
rect 9089 26899 9107 26917
rect 9125 26899 10240 26917
rect 8840 26881 10240 26899
rect 8840 26863 8855 26881
rect 8873 26863 8891 26881
rect 8909 26863 8927 26881
rect 8945 26863 8963 26881
rect 8981 26863 8999 26881
rect 9017 26863 9035 26881
rect 9053 26863 9071 26881
rect 9089 26863 9107 26881
rect 9125 26863 10240 26881
rect 8840 26845 10240 26863
rect 8840 26827 8855 26845
rect 8873 26827 8891 26845
rect 8909 26827 8927 26845
rect 8945 26827 8963 26845
rect 8981 26827 8999 26845
rect 9017 26827 9035 26845
rect 9053 26827 9071 26845
rect 9089 26827 9107 26845
rect 9125 26827 10240 26845
rect 8840 26809 10240 26827
rect 8840 26791 8855 26809
rect 8873 26791 8891 26809
rect 8909 26791 8927 26809
rect 8945 26791 8963 26809
rect 8981 26791 8999 26809
rect 9017 26791 9035 26809
rect 9053 26791 9071 26809
rect 9089 26791 9107 26809
rect 9125 26791 10240 26809
rect 8840 26773 10240 26791
rect 8840 26755 8855 26773
rect 8873 26755 8891 26773
rect 8909 26755 8927 26773
rect 8945 26755 8963 26773
rect 8981 26755 8999 26773
rect 9017 26755 9035 26773
rect 9053 26755 9071 26773
rect 9089 26755 9107 26773
rect 9125 26755 10240 26773
rect 8840 26737 10240 26755
rect 8840 26719 8855 26737
rect 8873 26719 8891 26737
rect 8909 26719 8927 26737
rect 8945 26719 8963 26737
rect 8981 26719 8999 26737
rect 9017 26719 9035 26737
rect 9053 26719 9071 26737
rect 9089 26719 9107 26737
rect 9125 26719 10240 26737
rect 8840 26701 10240 26719
rect 8840 26683 8855 26701
rect 8873 26683 8891 26701
rect 8909 26683 8927 26701
rect 8945 26683 8963 26701
rect 8981 26683 8999 26701
rect 9017 26683 9035 26701
rect 9053 26683 9071 26701
rect 9089 26683 9107 26701
rect 9125 26683 10240 26701
rect 8840 26665 10240 26683
rect 8840 26647 8855 26665
rect 8873 26647 8891 26665
rect 8909 26647 8927 26665
rect 8945 26647 8963 26665
rect 8981 26647 8999 26665
rect 9017 26647 9035 26665
rect 9053 26647 9071 26665
rect 9089 26647 9107 26665
rect 9125 26647 10240 26665
rect 8840 26629 10240 26647
rect 8840 26611 8855 26629
rect 8873 26611 8891 26629
rect 8909 26611 8927 26629
rect 8945 26611 8963 26629
rect 8981 26611 8999 26629
rect 9017 26611 9035 26629
rect 9053 26611 9071 26629
rect 9089 26611 9107 26629
rect 9125 26611 10240 26629
rect 8840 26593 10240 26611
rect 8840 26575 8855 26593
rect 8873 26575 8891 26593
rect 8909 26575 8927 26593
rect 8945 26575 8963 26593
rect 8981 26575 8999 26593
rect 9017 26575 9035 26593
rect 9053 26575 9071 26593
rect 9089 26575 9107 26593
rect 9125 26575 10240 26593
rect 8840 26557 10240 26575
rect 8840 26539 8855 26557
rect 8873 26539 8891 26557
rect 8909 26539 8927 26557
rect 8945 26539 8963 26557
rect 8981 26539 8999 26557
rect 9017 26539 9035 26557
rect 9053 26539 9071 26557
rect 9089 26539 9107 26557
rect 9125 26539 10240 26557
rect 8840 26521 10240 26539
rect 8840 26503 8855 26521
rect 8873 26503 8891 26521
rect 8909 26503 8927 26521
rect 8945 26503 8963 26521
rect 8981 26503 8999 26521
rect 9017 26503 9035 26521
rect 9053 26503 9071 26521
rect 9089 26503 9107 26521
rect 9125 26503 10240 26521
rect 8840 26485 10240 26503
rect 8840 26467 8855 26485
rect 8873 26467 8891 26485
rect 8909 26467 8927 26485
rect 8945 26467 8963 26485
rect 8981 26467 8999 26485
rect 9017 26467 9035 26485
rect 9053 26467 9071 26485
rect 9089 26467 9107 26485
rect 9125 26467 10240 26485
rect 8840 26440 10240 26467
rect 27820 19927 29100 19940
rect 27820 19909 28767 19927
rect 28785 19909 28803 19927
rect 28821 19909 28839 19927
rect 28857 19909 28875 19927
rect 28893 19909 28911 19927
rect 28929 19909 28947 19927
rect 28965 19909 28983 19927
rect 29001 19909 29019 19927
rect 29037 19909 29055 19927
rect 29073 19909 29100 19927
rect 27820 19891 29100 19909
rect 27820 19873 28767 19891
rect 28785 19873 28803 19891
rect 28821 19873 28839 19891
rect 28857 19873 28875 19891
rect 28893 19873 28911 19891
rect 28929 19873 28947 19891
rect 28965 19873 28983 19891
rect 29001 19873 29019 19891
rect 29037 19873 29055 19891
rect 29073 19873 29100 19891
rect 27820 19855 29100 19873
rect 27820 19837 28767 19855
rect 28785 19837 28803 19855
rect 28821 19837 28839 19855
rect 28857 19837 28875 19855
rect 28893 19837 28911 19855
rect 28929 19837 28947 19855
rect 28965 19837 28983 19855
rect 29001 19837 29019 19855
rect 29037 19837 29055 19855
rect 29073 19837 29100 19855
rect 27820 19819 29100 19837
rect 27820 19801 28767 19819
rect 28785 19801 28803 19819
rect 28821 19801 28839 19819
rect 28857 19801 28875 19819
rect 28893 19801 28911 19819
rect 28929 19801 28947 19819
rect 28965 19801 28983 19819
rect 29001 19801 29019 19819
rect 29037 19801 29055 19819
rect 29073 19801 29100 19819
rect 27820 19783 29100 19801
rect 27820 19765 28767 19783
rect 28785 19765 28803 19783
rect 28821 19765 28839 19783
rect 28857 19765 28875 19783
rect 28893 19765 28911 19783
rect 28929 19765 28947 19783
rect 28965 19765 28983 19783
rect 29001 19765 29019 19783
rect 29037 19765 29055 19783
rect 29073 19765 29100 19783
rect 27820 19747 29100 19765
rect 27820 19729 28767 19747
rect 28785 19729 28803 19747
rect 28821 19729 28839 19747
rect 28857 19729 28875 19747
rect 28893 19729 28911 19747
rect 28929 19729 28947 19747
rect 28965 19729 28983 19747
rect 29001 19729 29019 19747
rect 29037 19729 29055 19747
rect 29073 19729 29100 19747
rect 27820 19711 29100 19729
rect 27820 19693 28767 19711
rect 28785 19693 28803 19711
rect 28821 19693 28839 19711
rect 28857 19693 28875 19711
rect 28893 19693 28911 19711
rect 28929 19693 28947 19711
rect 28965 19693 28983 19711
rect 29001 19693 29019 19711
rect 29037 19693 29055 19711
rect 29073 19693 29100 19711
rect 27820 19675 29100 19693
rect 27820 19657 28767 19675
rect 28785 19657 28803 19675
rect 28821 19657 28839 19675
rect 28857 19657 28875 19675
rect 28893 19657 28911 19675
rect 28929 19657 28947 19675
rect 28965 19657 28983 19675
rect 29001 19657 29019 19675
rect 29037 19657 29055 19675
rect 29073 19657 29100 19675
rect 27820 19639 29100 19657
rect 27820 19621 28767 19639
rect 28785 19621 28803 19639
rect 28821 19621 28839 19639
rect 28857 19621 28875 19639
rect 28893 19621 28911 19639
rect 28929 19621 28947 19639
rect 28965 19621 28983 19639
rect 29001 19621 29019 19639
rect 29037 19621 29055 19639
rect 29073 19621 29100 19639
rect 27820 19603 29100 19621
rect 27820 19585 28767 19603
rect 28785 19585 28803 19603
rect 28821 19585 28839 19603
rect 28857 19585 28875 19603
rect 28893 19585 28911 19603
rect 28929 19585 28947 19603
rect 28965 19585 28983 19603
rect 29001 19585 29019 19603
rect 29037 19585 29055 19603
rect 29073 19585 29100 19603
rect 27820 19567 29100 19585
rect 27820 19549 28767 19567
rect 28785 19549 28803 19567
rect 28821 19549 28839 19567
rect 28857 19549 28875 19567
rect 28893 19549 28911 19567
rect 28929 19549 28947 19567
rect 28965 19549 28983 19567
rect 29001 19549 29019 19567
rect 29037 19549 29055 19567
rect 29073 19549 29100 19567
rect 27820 19531 29100 19549
rect 27820 19513 28767 19531
rect 28785 19513 28803 19531
rect 28821 19513 28839 19531
rect 28857 19513 28875 19531
rect 28893 19513 28911 19531
rect 28929 19513 28947 19531
rect 28965 19513 28983 19531
rect 29001 19513 29019 19531
rect 29037 19513 29055 19531
rect 29073 19513 29100 19531
rect 27820 19495 29100 19513
rect 27820 19477 28767 19495
rect 28785 19477 28803 19495
rect 28821 19477 28839 19495
rect 28857 19477 28875 19495
rect 28893 19477 28911 19495
rect 28929 19477 28947 19495
rect 28965 19477 28983 19495
rect 29001 19477 29019 19495
rect 29037 19477 29055 19495
rect 29073 19477 29100 19495
rect 27820 19459 29100 19477
rect 27820 19441 28767 19459
rect 28785 19441 28803 19459
rect 28821 19441 28839 19459
rect 28857 19441 28875 19459
rect 28893 19441 28911 19459
rect 28929 19441 28947 19459
rect 28965 19441 28983 19459
rect 29001 19441 29019 19459
rect 29037 19441 29055 19459
rect 29073 19441 29100 19459
rect 27820 19423 29100 19441
rect 27820 19405 28767 19423
rect 28785 19405 28803 19423
rect 28821 19405 28839 19423
rect 28857 19405 28875 19423
rect 28893 19405 28911 19423
rect 28929 19405 28947 19423
rect 28965 19405 28983 19423
rect 29001 19405 29019 19423
rect 29037 19405 29055 19423
rect 29073 19405 29100 19423
rect 27820 19387 29100 19405
rect 27820 19369 28767 19387
rect 28785 19369 28803 19387
rect 28821 19369 28839 19387
rect 28857 19369 28875 19387
rect 28893 19369 28911 19387
rect 28929 19369 28947 19387
rect 28965 19369 28983 19387
rect 29001 19369 29019 19387
rect 29037 19369 29055 19387
rect 29073 19369 29100 19387
rect 27820 19351 29100 19369
rect 27820 19333 28767 19351
rect 28785 19333 28803 19351
rect 28821 19333 28839 19351
rect 28857 19333 28875 19351
rect 28893 19333 28911 19351
rect 28929 19333 28947 19351
rect 28965 19333 28983 19351
rect 29001 19333 29019 19351
rect 29037 19333 29055 19351
rect 29073 19333 29100 19351
rect 27820 19315 29100 19333
rect 27820 19297 28767 19315
rect 28785 19297 28803 19315
rect 28821 19297 28839 19315
rect 28857 19297 28875 19315
rect 28893 19297 28911 19315
rect 28929 19297 28947 19315
rect 28965 19297 28983 19315
rect 29001 19297 29019 19315
rect 29037 19297 29055 19315
rect 29073 19297 29100 19315
rect 27820 19279 29100 19297
rect 27820 19261 28767 19279
rect 28785 19261 28803 19279
rect 28821 19261 28839 19279
rect 28857 19261 28875 19279
rect 28893 19261 28911 19279
rect 28929 19261 28947 19279
rect 28965 19261 28983 19279
rect 29001 19261 29019 19279
rect 29037 19261 29055 19279
rect 29073 19261 29100 19279
rect 27820 19243 29100 19261
rect 27820 19225 28767 19243
rect 28785 19225 28803 19243
rect 28821 19225 28839 19243
rect 28857 19225 28875 19243
rect 28893 19225 28911 19243
rect 28929 19225 28947 19243
rect 28965 19225 28983 19243
rect 29001 19225 29019 19243
rect 29037 19225 29055 19243
rect 29073 19225 29100 19243
rect 27820 19207 29100 19225
rect 27820 19189 28767 19207
rect 28785 19189 28803 19207
rect 28821 19189 28839 19207
rect 28857 19189 28875 19207
rect 28893 19189 28911 19207
rect 28929 19189 28947 19207
rect 28965 19189 28983 19207
rect 29001 19189 29019 19207
rect 29037 19189 29055 19207
rect 29073 19189 29100 19207
rect 27820 19171 29100 19189
rect 27820 19153 28767 19171
rect 28785 19153 28803 19171
rect 28821 19153 28839 19171
rect 28857 19153 28875 19171
rect 28893 19153 28911 19171
rect 28929 19153 28947 19171
rect 28965 19153 28983 19171
rect 29001 19153 29019 19171
rect 29037 19153 29055 19171
rect 29073 19153 29100 19171
rect 27820 19135 29100 19153
rect 27820 19117 28767 19135
rect 28785 19117 28803 19135
rect 28821 19117 28839 19135
rect 28857 19117 28875 19135
rect 28893 19117 28911 19135
rect 28929 19117 28947 19135
rect 28965 19117 28983 19135
rect 29001 19117 29019 19135
rect 29037 19117 29055 19135
rect 29073 19117 29100 19135
rect 27820 19099 29100 19117
rect 27820 19081 28767 19099
rect 28785 19081 28803 19099
rect 28821 19081 28839 19099
rect 28857 19081 28875 19099
rect 28893 19081 28911 19099
rect 28929 19081 28947 19099
rect 28965 19081 28983 19099
rect 29001 19081 29019 19099
rect 29037 19081 29055 19099
rect 29073 19081 29100 19099
rect 27820 19063 29100 19081
rect 27820 19045 28767 19063
rect 28785 19045 28803 19063
rect 28821 19045 28839 19063
rect 28857 19045 28875 19063
rect 28893 19045 28911 19063
rect 28929 19045 28947 19063
rect 28965 19045 28983 19063
rect 29001 19045 29019 19063
rect 29037 19045 29055 19063
rect 29073 19045 29100 19063
rect 27820 19027 29100 19045
rect 27820 19009 28767 19027
rect 28785 19009 28803 19027
rect 28821 19009 28839 19027
rect 28857 19009 28875 19027
rect 28893 19009 28911 19027
rect 28929 19009 28947 19027
rect 28965 19009 28983 19027
rect 29001 19009 29019 19027
rect 29037 19009 29055 19027
rect 29073 19009 29100 19027
rect 27820 18991 29100 19009
rect 27820 18973 28767 18991
rect 28785 18973 28803 18991
rect 28821 18973 28839 18991
rect 28857 18973 28875 18991
rect 28893 18973 28911 18991
rect 28929 18973 28947 18991
rect 28965 18973 28983 18991
rect 29001 18973 29019 18991
rect 29037 18973 29055 18991
rect 29073 18973 29100 18991
rect 27820 18955 29100 18973
rect 27820 18937 28767 18955
rect 28785 18937 28803 18955
rect 28821 18937 28839 18955
rect 28857 18937 28875 18955
rect 28893 18937 28911 18955
rect 28929 18937 28947 18955
rect 28965 18937 28983 18955
rect 29001 18937 29019 18955
rect 29037 18937 29055 18955
rect 29073 18937 29100 18955
rect 27820 18919 29100 18937
rect 27820 18901 28767 18919
rect 28785 18901 28803 18919
rect 28821 18901 28839 18919
rect 28857 18901 28875 18919
rect 28893 18901 28911 18919
rect 28929 18901 28947 18919
rect 28965 18901 28983 18919
rect 29001 18901 29019 18919
rect 29037 18901 29055 18919
rect 29073 18901 29100 18919
rect 27820 18883 29100 18901
rect 27820 18865 28767 18883
rect 28785 18865 28803 18883
rect 28821 18865 28839 18883
rect 28857 18865 28875 18883
rect 28893 18865 28911 18883
rect 28929 18865 28947 18883
rect 28965 18865 28983 18883
rect 29001 18865 29019 18883
rect 29037 18865 29055 18883
rect 29073 18865 29100 18883
rect 27820 18847 29100 18865
rect 27820 18829 28767 18847
rect 28785 18829 28803 18847
rect 28821 18829 28839 18847
rect 28857 18829 28875 18847
rect 28893 18829 28911 18847
rect 28929 18829 28947 18847
rect 28965 18829 28983 18847
rect 29001 18829 29019 18847
rect 29037 18829 29055 18847
rect 29073 18829 29100 18847
rect 27820 18811 29100 18829
rect 27820 18793 28767 18811
rect 28785 18793 28803 18811
rect 28821 18793 28839 18811
rect 28857 18793 28875 18811
rect 28893 18793 28911 18811
rect 28929 18793 28947 18811
rect 28965 18793 28983 18811
rect 29001 18793 29019 18811
rect 29037 18793 29055 18811
rect 29073 18793 29100 18811
rect 27820 18775 29100 18793
rect 27820 18757 28767 18775
rect 28785 18757 28803 18775
rect 28821 18757 28839 18775
rect 28857 18757 28875 18775
rect 28893 18757 28911 18775
rect 28929 18757 28947 18775
rect 28965 18757 28983 18775
rect 29001 18757 29019 18775
rect 29037 18757 29055 18775
rect 29073 18757 29100 18775
rect 27820 18739 29100 18757
rect 27820 18721 28767 18739
rect 28785 18721 28803 18739
rect 28821 18721 28839 18739
rect 28857 18721 28875 18739
rect 28893 18721 28911 18739
rect 28929 18721 28947 18739
rect 28965 18721 28983 18739
rect 29001 18721 29019 18739
rect 29037 18721 29055 18739
rect 29073 18721 29100 18739
rect 27820 18703 29100 18721
rect 27820 18685 28767 18703
rect 28785 18685 28803 18703
rect 28821 18685 28839 18703
rect 28857 18685 28875 18703
rect 28893 18685 28911 18703
rect 28929 18685 28947 18703
rect 28965 18685 28983 18703
rect 29001 18685 29019 18703
rect 29037 18685 29055 18703
rect 29073 18685 29100 18703
rect 27820 18667 29100 18685
rect 27820 18649 28767 18667
rect 28785 18649 28803 18667
rect 28821 18649 28839 18667
rect 28857 18649 28875 18667
rect 28893 18649 28911 18667
rect 28929 18649 28947 18667
rect 28965 18649 28983 18667
rect 29001 18649 29019 18667
rect 29037 18649 29055 18667
rect 29073 18649 29100 18667
rect 27820 18631 29100 18649
rect 27820 18613 28767 18631
rect 28785 18613 28803 18631
rect 28821 18613 28839 18631
rect 28857 18613 28875 18631
rect 28893 18613 28911 18631
rect 28929 18613 28947 18631
rect 28965 18613 28983 18631
rect 29001 18613 29019 18631
rect 29037 18613 29055 18631
rect 29073 18613 29100 18631
rect 27820 18595 29100 18613
rect 27820 18577 28767 18595
rect 28785 18577 28803 18595
rect 28821 18577 28839 18595
rect 28857 18577 28875 18595
rect 28893 18577 28911 18595
rect 28929 18577 28947 18595
rect 28965 18577 28983 18595
rect 29001 18577 29019 18595
rect 29037 18577 29055 18595
rect 29073 18577 29100 18595
rect 27820 18559 29100 18577
rect 27820 18541 28767 18559
rect 28785 18541 28803 18559
rect 28821 18541 28839 18559
rect 28857 18541 28875 18559
rect 28893 18541 28911 18559
rect 28929 18541 28947 18559
rect 28965 18541 28983 18559
rect 29001 18541 29019 18559
rect 29037 18541 29055 18559
rect 29073 18541 29100 18559
rect 27820 18523 29100 18541
rect 27820 18505 28767 18523
rect 28785 18505 28803 18523
rect 28821 18505 28839 18523
rect 28857 18505 28875 18523
rect 28893 18505 28911 18523
rect 28929 18505 28947 18523
rect 28965 18505 28983 18523
rect 29001 18505 29019 18523
rect 29037 18505 29055 18523
rect 29073 18505 29100 18523
rect 27820 18487 29100 18505
rect 27820 18469 28767 18487
rect 28785 18469 28803 18487
rect 28821 18469 28839 18487
rect 28857 18469 28875 18487
rect 28893 18469 28911 18487
rect 28929 18469 28947 18487
rect 28965 18469 28983 18487
rect 29001 18469 29019 18487
rect 29037 18469 29055 18487
rect 29073 18469 29100 18487
rect 27820 18451 29100 18469
rect 27820 18433 28767 18451
rect 28785 18433 28803 18451
rect 28821 18433 28839 18451
rect 28857 18433 28875 18451
rect 28893 18433 28911 18451
rect 28929 18433 28947 18451
rect 28965 18433 28983 18451
rect 29001 18433 29019 18451
rect 29037 18433 29055 18451
rect 29073 18433 29100 18451
rect 27820 18415 29100 18433
rect 27820 18397 28767 18415
rect 28785 18397 28803 18415
rect 28821 18397 28839 18415
rect 28857 18397 28875 18415
rect 28893 18397 28911 18415
rect 28929 18397 28947 18415
rect 28965 18397 28983 18415
rect 29001 18397 29019 18415
rect 29037 18397 29055 18415
rect 29073 18397 29100 18415
rect 27820 18379 29100 18397
rect 27820 18361 28767 18379
rect 28785 18361 28803 18379
rect 28821 18361 28839 18379
rect 28857 18361 28875 18379
rect 28893 18361 28911 18379
rect 28929 18361 28947 18379
rect 28965 18361 28983 18379
rect 29001 18361 29019 18379
rect 29037 18361 29055 18379
rect 29073 18361 29100 18379
rect 27820 18343 29100 18361
rect 27820 18325 28767 18343
rect 28785 18325 28803 18343
rect 28821 18325 28839 18343
rect 28857 18325 28875 18343
rect 28893 18325 28911 18343
rect 28929 18325 28947 18343
rect 28965 18325 28983 18343
rect 29001 18325 29019 18343
rect 29037 18325 29055 18343
rect 29073 18325 29100 18343
rect 27820 18307 29100 18325
rect 27820 18289 28767 18307
rect 28785 18289 28803 18307
rect 28821 18289 28839 18307
rect 28857 18289 28875 18307
rect 28893 18289 28911 18307
rect 28929 18289 28947 18307
rect 28965 18289 28983 18307
rect 29001 18289 29019 18307
rect 29037 18289 29055 18307
rect 29073 18289 29100 18307
rect 27820 18271 29100 18289
rect 27820 18253 28767 18271
rect 28785 18253 28803 18271
rect 28821 18253 28839 18271
rect 28857 18253 28875 18271
rect 28893 18253 28911 18271
rect 28929 18253 28947 18271
rect 28965 18253 28983 18271
rect 29001 18253 29019 18271
rect 29037 18253 29055 18271
rect 29073 18253 29100 18271
rect 27820 18235 29100 18253
rect 27820 18217 28767 18235
rect 28785 18217 28803 18235
rect 28821 18217 28839 18235
rect 28857 18217 28875 18235
rect 28893 18217 28911 18235
rect 28929 18217 28947 18235
rect 28965 18217 28983 18235
rect 29001 18217 29019 18235
rect 29037 18217 29055 18235
rect 29073 18217 29100 18235
rect 27820 18199 29100 18217
rect 27820 18181 28767 18199
rect 28785 18181 28803 18199
rect 28821 18181 28839 18199
rect 28857 18181 28875 18199
rect 28893 18181 28911 18199
rect 28929 18181 28947 18199
rect 28965 18181 28983 18199
rect 29001 18181 29019 18199
rect 29037 18181 29055 18199
rect 29073 18181 29100 18199
rect 27820 18163 29100 18181
rect 27820 18145 28767 18163
rect 28785 18145 28803 18163
rect 28821 18145 28839 18163
rect 28857 18145 28875 18163
rect 28893 18145 28911 18163
rect 28929 18145 28947 18163
rect 28965 18145 28983 18163
rect 29001 18145 29019 18163
rect 29037 18145 29055 18163
rect 29073 18145 29100 18163
rect 27820 18127 29100 18145
rect 27820 18109 28767 18127
rect 28785 18109 28803 18127
rect 28821 18109 28839 18127
rect 28857 18109 28875 18127
rect 28893 18109 28911 18127
rect 28929 18109 28947 18127
rect 28965 18109 28983 18127
rect 29001 18109 29019 18127
rect 29037 18109 29055 18127
rect 29073 18109 29100 18127
rect 27820 18091 29100 18109
rect 27820 18073 28767 18091
rect 28785 18073 28803 18091
rect 28821 18073 28839 18091
rect 28857 18073 28875 18091
rect 28893 18073 28911 18091
rect 28929 18073 28947 18091
rect 28965 18073 28983 18091
rect 29001 18073 29019 18091
rect 29037 18073 29055 18091
rect 29073 18073 29100 18091
rect 27820 18060 29100 18073
rect 8840 11565 10240 11580
rect 8840 11547 8855 11565
rect 8873 11547 8891 11565
rect 8909 11547 8927 11565
rect 8945 11547 8963 11565
rect 8981 11547 8999 11565
rect 9017 11547 9035 11565
rect 9053 11547 9071 11565
rect 9089 11547 9107 11565
rect 9125 11547 10240 11565
rect 8840 11529 10240 11547
rect 8840 11511 8855 11529
rect 8873 11511 8891 11529
rect 8909 11511 8927 11529
rect 8945 11511 8963 11529
rect 8981 11511 8999 11529
rect 9017 11511 9035 11529
rect 9053 11511 9071 11529
rect 9089 11511 9107 11529
rect 9125 11511 10240 11529
rect 8840 11493 10240 11511
rect 8840 11475 8855 11493
rect 8873 11475 8891 11493
rect 8909 11475 8927 11493
rect 8945 11475 8963 11493
rect 8981 11475 8999 11493
rect 9017 11475 9035 11493
rect 9053 11475 9071 11493
rect 9089 11475 9107 11493
rect 9125 11475 10240 11493
rect 8840 11457 10240 11475
rect 8840 11439 8855 11457
rect 8873 11439 8891 11457
rect 8909 11439 8927 11457
rect 8945 11439 8963 11457
rect 8981 11439 8999 11457
rect 9017 11439 9035 11457
rect 9053 11439 9071 11457
rect 9089 11439 9107 11457
rect 9125 11439 10240 11457
rect 8840 11421 10240 11439
rect 8840 11403 8855 11421
rect 8873 11403 8891 11421
rect 8909 11403 8927 11421
rect 8945 11403 8963 11421
rect 8981 11403 8999 11421
rect 9017 11403 9035 11421
rect 9053 11403 9071 11421
rect 9089 11403 9107 11421
rect 9125 11403 10240 11421
rect 8840 11385 10240 11403
rect 8840 11367 8855 11385
rect 8873 11367 8891 11385
rect 8909 11367 8927 11385
rect 8945 11367 8963 11385
rect 8981 11367 8999 11385
rect 9017 11367 9035 11385
rect 9053 11367 9071 11385
rect 9089 11367 9107 11385
rect 9125 11367 10240 11385
rect 8840 11349 10240 11367
rect 8840 11331 8855 11349
rect 8873 11331 8891 11349
rect 8909 11331 8927 11349
rect 8945 11331 8963 11349
rect 8981 11331 8999 11349
rect 9017 11331 9035 11349
rect 9053 11331 9071 11349
rect 9089 11331 9107 11349
rect 9125 11331 10240 11349
rect 8840 11313 10240 11331
rect 8840 11295 8855 11313
rect 8873 11295 8891 11313
rect 8909 11295 8927 11313
rect 8945 11295 8963 11313
rect 8981 11295 8999 11313
rect 9017 11295 9035 11313
rect 9053 11295 9071 11313
rect 9089 11295 9107 11313
rect 9125 11295 10240 11313
rect 8840 11277 10240 11295
rect 8840 11259 8855 11277
rect 8873 11259 8891 11277
rect 8909 11259 8927 11277
rect 8945 11259 8963 11277
rect 8981 11259 8999 11277
rect 9017 11259 9035 11277
rect 9053 11259 9071 11277
rect 9089 11259 9107 11277
rect 9125 11259 10240 11277
rect 8840 11241 10240 11259
rect 8840 11223 8855 11241
rect 8873 11223 8891 11241
rect 8909 11223 8927 11241
rect 8945 11223 8963 11241
rect 8981 11223 8999 11241
rect 9017 11223 9035 11241
rect 9053 11223 9071 11241
rect 9089 11223 9107 11241
rect 9125 11223 10240 11241
rect 8840 11205 10240 11223
rect 8840 11187 8855 11205
rect 8873 11187 8891 11205
rect 8909 11187 8927 11205
rect 8945 11187 8963 11205
rect 8981 11187 8999 11205
rect 9017 11187 9035 11205
rect 9053 11187 9071 11205
rect 9089 11187 9107 11205
rect 9125 11187 10240 11205
rect 8840 11169 10240 11187
rect 8840 11151 8855 11169
rect 8873 11151 8891 11169
rect 8909 11151 8927 11169
rect 8945 11151 8963 11169
rect 8981 11151 8999 11169
rect 9017 11151 9035 11169
rect 9053 11151 9071 11169
rect 9089 11151 9107 11169
rect 9125 11151 10240 11169
rect 8840 11133 10240 11151
rect 8840 11115 8855 11133
rect 8873 11115 8891 11133
rect 8909 11115 8927 11133
rect 8945 11115 8963 11133
rect 8981 11115 8999 11133
rect 9017 11115 9035 11133
rect 9053 11115 9071 11133
rect 9089 11115 9107 11133
rect 9125 11115 10240 11133
rect 8840 11097 10240 11115
rect 8840 11079 8855 11097
rect 8873 11079 8891 11097
rect 8909 11079 8927 11097
rect 8945 11079 8963 11097
rect 8981 11079 8999 11097
rect 9017 11079 9035 11097
rect 9053 11079 9071 11097
rect 9089 11079 9107 11097
rect 9125 11079 10240 11097
rect 8840 11061 10240 11079
rect 8840 11043 8855 11061
rect 8873 11043 8891 11061
rect 8909 11043 8927 11061
rect 8945 11043 8963 11061
rect 8981 11043 8999 11061
rect 9017 11043 9035 11061
rect 9053 11043 9071 11061
rect 9089 11043 9107 11061
rect 9125 11043 10240 11061
rect 8840 11025 10240 11043
rect 8840 11007 8855 11025
rect 8873 11007 8891 11025
rect 8909 11007 8927 11025
rect 8945 11007 8963 11025
rect 8981 11007 8999 11025
rect 9017 11007 9035 11025
rect 9053 11007 9071 11025
rect 9089 11007 9107 11025
rect 9125 11007 10240 11025
rect 8840 10989 10240 11007
rect 8840 10971 8855 10989
rect 8873 10971 8891 10989
rect 8909 10971 8927 10989
rect 8945 10971 8963 10989
rect 8981 10971 8999 10989
rect 9017 10971 9035 10989
rect 9053 10971 9071 10989
rect 9089 10971 9107 10989
rect 9125 10971 10240 10989
rect 8840 10953 10240 10971
rect 8840 10935 8855 10953
rect 8873 10935 8891 10953
rect 8909 10935 8927 10953
rect 8945 10935 8963 10953
rect 8981 10935 8999 10953
rect 9017 10935 9035 10953
rect 9053 10935 9071 10953
rect 9089 10935 9107 10953
rect 9125 10935 10240 10953
rect 8840 10917 10240 10935
rect 8840 10899 8855 10917
rect 8873 10899 8891 10917
rect 8909 10899 8927 10917
rect 8945 10899 8963 10917
rect 8981 10899 8999 10917
rect 9017 10899 9035 10917
rect 9053 10899 9071 10917
rect 9089 10899 9107 10917
rect 9125 10899 10240 10917
rect 8840 10881 10240 10899
rect 8840 10863 8855 10881
rect 8873 10863 8891 10881
rect 8909 10863 8927 10881
rect 8945 10863 8963 10881
rect 8981 10863 8999 10881
rect 9017 10863 9035 10881
rect 9053 10863 9071 10881
rect 9089 10863 9107 10881
rect 9125 10863 10240 10881
rect 8840 10845 10240 10863
rect 8840 10827 8855 10845
rect 8873 10827 8891 10845
rect 8909 10827 8927 10845
rect 8945 10827 8963 10845
rect 8981 10827 8999 10845
rect 9017 10827 9035 10845
rect 9053 10827 9071 10845
rect 9089 10827 9107 10845
rect 9125 10827 10240 10845
rect 8840 10809 10240 10827
rect 8840 10791 8855 10809
rect 8873 10791 8891 10809
rect 8909 10791 8927 10809
rect 8945 10791 8963 10809
rect 8981 10791 8999 10809
rect 9017 10791 9035 10809
rect 9053 10791 9071 10809
rect 9089 10791 9107 10809
rect 9125 10791 10240 10809
rect 8840 10773 10240 10791
rect 8840 10755 8855 10773
rect 8873 10755 8891 10773
rect 8909 10755 8927 10773
rect 8945 10755 8963 10773
rect 8981 10755 8999 10773
rect 9017 10755 9035 10773
rect 9053 10755 9071 10773
rect 9089 10755 9107 10773
rect 9125 10755 10240 10773
rect 8840 10740 10240 10755
<< m2contact >>
rect 8855 27115 8873 27133
rect 8891 27115 8909 27133
rect 8927 27115 8945 27133
rect 8963 27115 8981 27133
rect 8999 27115 9017 27133
rect 9035 27115 9053 27133
rect 9071 27115 9089 27133
rect 9107 27115 9125 27133
rect 8855 27079 8873 27097
rect 8891 27079 8909 27097
rect 8927 27079 8945 27097
rect 8963 27079 8981 27097
rect 8999 27079 9017 27097
rect 9035 27079 9053 27097
rect 9071 27079 9089 27097
rect 9107 27079 9125 27097
rect 8855 27043 8873 27061
rect 8891 27043 8909 27061
rect 8927 27043 8945 27061
rect 8963 27043 8981 27061
rect 8999 27043 9017 27061
rect 9035 27043 9053 27061
rect 9071 27043 9089 27061
rect 9107 27043 9125 27061
rect 8855 27007 8873 27025
rect 8891 27007 8909 27025
rect 8927 27007 8945 27025
rect 8963 27007 8981 27025
rect 8999 27007 9017 27025
rect 9035 27007 9053 27025
rect 9071 27007 9089 27025
rect 9107 27007 9125 27025
rect 8855 26971 8873 26989
rect 8891 26971 8909 26989
rect 8927 26971 8945 26989
rect 8963 26971 8981 26989
rect 8999 26971 9017 26989
rect 9035 26971 9053 26989
rect 9071 26971 9089 26989
rect 9107 26971 9125 26989
rect 8855 26935 8873 26953
rect 8891 26935 8909 26953
rect 8927 26935 8945 26953
rect 8963 26935 8981 26953
rect 8999 26935 9017 26953
rect 9035 26935 9053 26953
rect 9071 26935 9089 26953
rect 9107 26935 9125 26953
rect 8855 26899 8873 26917
rect 8891 26899 8909 26917
rect 8927 26899 8945 26917
rect 8963 26899 8981 26917
rect 8999 26899 9017 26917
rect 9035 26899 9053 26917
rect 9071 26899 9089 26917
rect 9107 26899 9125 26917
rect 8855 26863 8873 26881
rect 8891 26863 8909 26881
rect 8927 26863 8945 26881
rect 8963 26863 8981 26881
rect 8999 26863 9017 26881
rect 9035 26863 9053 26881
rect 9071 26863 9089 26881
rect 9107 26863 9125 26881
rect 8855 26827 8873 26845
rect 8891 26827 8909 26845
rect 8927 26827 8945 26845
rect 8963 26827 8981 26845
rect 8999 26827 9017 26845
rect 9035 26827 9053 26845
rect 9071 26827 9089 26845
rect 9107 26827 9125 26845
rect 8855 26791 8873 26809
rect 8891 26791 8909 26809
rect 8927 26791 8945 26809
rect 8963 26791 8981 26809
rect 8999 26791 9017 26809
rect 9035 26791 9053 26809
rect 9071 26791 9089 26809
rect 9107 26791 9125 26809
rect 8855 26755 8873 26773
rect 8891 26755 8909 26773
rect 8927 26755 8945 26773
rect 8963 26755 8981 26773
rect 8999 26755 9017 26773
rect 9035 26755 9053 26773
rect 9071 26755 9089 26773
rect 9107 26755 9125 26773
rect 8855 26719 8873 26737
rect 8891 26719 8909 26737
rect 8927 26719 8945 26737
rect 8963 26719 8981 26737
rect 8999 26719 9017 26737
rect 9035 26719 9053 26737
rect 9071 26719 9089 26737
rect 9107 26719 9125 26737
rect 8855 26683 8873 26701
rect 8891 26683 8909 26701
rect 8927 26683 8945 26701
rect 8963 26683 8981 26701
rect 8999 26683 9017 26701
rect 9035 26683 9053 26701
rect 9071 26683 9089 26701
rect 9107 26683 9125 26701
rect 8855 26647 8873 26665
rect 8891 26647 8909 26665
rect 8927 26647 8945 26665
rect 8963 26647 8981 26665
rect 8999 26647 9017 26665
rect 9035 26647 9053 26665
rect 9071 26647 9089 26665
rect 9107 26647 9125 26665
rect 8855 26611 8873 26629
rect 8891 26611 8909 26629
rect 8927 26611 8945 26629
rect 8963 26611 8981 26629
rect 8999 26611 9017 26629
rect 9035 26611 9053 26629
rect 9071 26611 9089 26629
rect 9107 26611 9125 26629
rect 8855 26575 8873 26593
rect 8891 26575 8909 26593
rect 8927 26575 8945 26593
rect 8963 26575 8981 26593
rect 8999 26575 9017 26593
rect 9035 26575 9053 26593
rect 9071 26575 9089 26593
rect 9107 26575 9125 26593
rect 8855 26539 8873 26557
rect 8891 26539 8909 26557
rect 8927 26539 8945 26557
rect 8963 26539 8981 26557
rect 8999 26539 9017 26557
rect 9035 26539 9053 26557
rect 9071 26539 9089 26557
rect 9107 26539 9125 26557
rect 8855 26503 8873 26521
rect 8891 26503 8909 26521
rect 8927 26503 8945 26521
rect 8963 26503 8981 26521
rect 8999 26503 9017 26521
rect 9035 26503 9053 26521
rect 9071 26503 9089 26521
rect 9107 26503 9125 26521
rect 8855 26467 8873 26485
rect 8891 26467 8909 26485
rect 8927 26467 8945 26485
rect 8963 26467 8981 26485
rect 8999 26467 9017 26485
rect 9035 26467 9053 26485
rect 9071 26467 9089 26485
rect 9107 26467 9125 26485
rect 28767 19909 28785 19927
rect 28803 19909 28821 19927
rect 28839 19909 28857 19927
rect 28875 19909 28893 19927
rect 28911 19909 28929 19927
rect 28947 19909 28965 19927
rect 28983 19909 29001 19927
rect 29019 19909 29037 19927
rect 29055 19909 29073 19927
rect 28767 19873 28785 19891
rect 28803 19873 28821 19891
rect 28839 19873 28857 19891
rect 28875 19873 28893 19891
rect 28911 19873 28929 19891
rect 28947 19873 28965 19891
rect 28983 19873 29001 19891
rect 29019 19873 29037 19891
rect 29055 19873 29073 19891
rect 28767 19837 28785 19855
rect 28803 19837 28821 19855
rect 28839 19837 28857 19855
rect 28875 19837 28893 19855
rect 28911 19837 28929 19855
rect 28947 19837 28965 19855
rect 28983 19837 29001 19855
rect 29019 19837 29037 19855
rect 29055 19837 29073 19855
rect 28767 19801 28785 19819
rect 28803 19801 28821 19819
rect 28839 19801 28857 19819
rect 28875 19801 28893 19819
rect 28911 19801 28929 19819
rect 28947 19801 28965 19819
rect 28983 19801 29001 19819
rect 29019 19801 29037 19819
rect 29055 19801 29073 19819
rect 28767 19765 28785 19783
rect 28803 19765 28821 19783
rect 28839 19765 28857 19783
rect 28875 19765 28893 19783
rect 28911 19765 28929 19783
rect 28947 19765 28965 19783
rect 28983 19765 29001 19783
rect 29019 19765 29037 19783
rect 29055 19765 29073 19783
rect 28767 19729 28785 19747
rect 28803 19729 28821 19747
rect 28839 19729 28857 19747
rect 28875 19729 28893 19747
rect 28911 19729 28929 19747
rect 28947 19729 28965 19747
rect 28983 19729 29001 19747
rect 29019 19729 29037 19747
rect 29055 19729 29073 19747
rect 28767 19693 28785 19711
rect 28803 19693 28821 19711
rect 28839 19693 28857 19711
rect 28875 19693 28893 19711
rect 28911 19693 28929 19711
rect 28947 19693 28965 19711
rect 28983 19693 29001 19711
rect 29019 19693 29037 19711
rect 29055 19693 29073 19711
rect 28767 19657 28785 19675
rect 28803 19657 28821 19675
rect 28839 19657 28857 19675
rect 28875 19657 28893 19675
rect 28911 19657 28929 19675
rect 28947 19657 28965 19675
rect 28983 19657 29001 19675
rect 29019 19657 29037 19675
rect 29055 19657 29073 19675
rect 28767 19621 28785 19639
rect 28803 19621 28821 19639
rect 28839 19621 28857 19639
rect 28875 19621 28893 19639
rect 28911 19621 28929 19639
rect 28947 19621 28965 19639
rect 28983 19621 29001 19639
rect 29019 19621 29037 19639
rect 29055 19621 29073 19639
rect 28767 19585 28785 19603
rect 28803 19585 28821 19603
rect 28839 19585 28857 19603
rect 28875 19585 28893 19603
rect 28911 19585 28929 19603
rect 28947 19585 28965 19603
rect 28983 19585 29001 19603
rect 29019 19585 29037 19603
rect 29055 19585 29073 19603
rect 28767 19549 28785 19567
rect 28803 19549 28821 19567
rect 28839 19549 28857 19567
rect 28875 19549 28893 19567
rect 28911 19549 28929 19567
rect 28947 19549 28965 19567
rect 28983 19549 29001 19567
rect 29019 19549 29037 19567
rect 29055 19549 29073 19567
rect 28767 19513 28785 19531
rect 28803 19513 28821 19531
rect 28839 19513 28857 19531
rect 28875 19513 28893 19531
rect 28911 19513 28929 19531
rect 28947 19513 28965 19531
rect 28983 19513 29001 19531
rect 29019 19513 29037 19531
rect 29055 19513 29073 19531
rect 28767 19477 28785 19495
rect 28803 19477 28821 19495
rect 28839 19477 28857 19495
rect 28875 19477 28893 19495
rect 28911 19477 28929 19495
rect 28947 19477 28965 19495
rect 28983 19477 29001 19495
rect 29019 19477 29037 19495
rect 29055 19477 29073 19495
rect 28767 19441 28785 19459
rect 28803 19441 28821 19459
rect 28839 19441 28857 19459
rect 28875 19441 28893 19459
rect 28911 19441 28929 19459
rect 28947 19441 28965 19459
rect 28983 19441 29001 19459
rect 29019 19441 29037 19459
rect 29055 19441 29073 19459
rect 28767 19405 28785 19423
rect 28803 19405 28821 19423
rect 28839 19405 28857 19423
rect 28875 19405 28893 19423
rect 28911 19405 28929 19423
rect 28947 19405 28965 19423
rect 28983 19405 29001 19423
rect 29019 19405 29037 19423
rect 29055 19405 29073 19423
rect 28767 19369 28785 19387
rect 28803 19369 28821 19387
rect 28839 19369 28857 19387
rect 28875 19369 28893 19387
rect 28911 19369 28929 19387
rect 28947 19369 28965 19387
rect 28983 19369 29001 19387
rect 29019 19369 29037 19387
rect 29055 19369 29073 19387
rect 28767 19333 28785 19351
rect 28803 19333 28821 19351
rect 28839 19333 28857 19351
rect 28875 19333 28893 19351
rect 28911 19333 28929 19351
rect 28947 19333 28965 19351
rect 28983 19333 29001 19351
rect 29019 19333 29037 19351
rect 29055 19333 29073 19351
rect 28767 19297 28785 19315
rect 28803 19297 28821 19315
rect 28839 19297 28857 19315
rect 28875 19297 28893 19315
rect 28911 19297 28929 19315
rect 28947 19297 28965 19315
rect 28983 19297 29001 19315
rect 29019 19297 29037 19315
rect 29055 19297 29073 19315
rect 28767 19261 28785 19279
rect 28803 19261 28821 19279
rect 28839 19261 28857 19279
rect 28875 19261 28893 19279
rect 28911 19261 28929 19279
rect 28947 19261 28965 19279
rect 28983 19261 29001 19279
rect 29019 19261 29037 19279
rect 29055 19261 29073 19279
rect 28767 19225 28785 19243
rect 28803 19225 28821 19243
rect 28839 19225 28857 19243
rect 28875 19225 28893 19243
rect 28911 19225 28929 19243
rect 28947 19225 28965 19243
rect 28983 19225 29001 19243
rect 29019 19225 29037 19243
rect 29055 19225 29073 19243
rect 28767 19189 28785 19207
rect 28803 19189 28821 19207
rect 28839 19189 28857 19207
rect 28875 19189 28893 19207
rect 28911 19189 28929 19207
rect 28947 19189 28965 19207
rect 28983 19189 29001 19207
rect 29019 19189 29037 19207
rect 29055 19189 29073 19207
rect 28767 19153 28785 19171
rect 28803 19153 28821 19171
rect 28839 19153 28857 19171
rect 28875 19153 28893 19171
rect 28911 19153 28929 19171
rect 28947 19153 28965 19171
rect 28983 19153 29001 19171
rect 29019 19153 29037 19171
rect 29055 19153 29073 19171
rect 28767 19117 28785 19135
rect 28803 19117 28821 19135
rect 28839 19117 28857 19135
rect 28875 19117 28893 19135
rect 28911 19117 28929 19135
rect 28947 19117 28965 19135
rect 28983 19117 29001 19135
rect 29019 19117 29037 19135
rect 29055 19117 29073 19135
rect 28767 19081 28785 19099
rect 28803 19081 28821 19099
rect 28839 19081 28857 19099
rect 28875 19081 28893 19099
rect 28911 19081 28929 19099
rect 28947 19081 28965 19099
rect 28983 19081 29001 19099
rect 29019 19081 29037 19099
rect 29055 19081 29073 19099
rect 28767 19045 28785 19063
rect 28803 19045 28821 19063
rect 28839 19045 28857 19063
rect 28875 19045 28893 19063
rect 28911 19045 28929 19063
rect 28947 19045 28965 19063
rect 28983 19045 29001 19063
rect 29019 19045 29037 19063
rect 29055 19045 29073 19063
rect 28767 19009 28785 19027
rect 28803 19009 28821 19027
rect 28839 19009 28857 19027
rect 28875 19009 28893 19027
rect 28911 19009 28929 19027
rect 28947 19009 28965 19027
rect 28983 19009 29001 19027
rect 29019 19009 29037 19027
rect 29055 19009 29073 19027
rect 28767 18973 28785 18991
rect 28803 18973 28821 18991
rect 28839 18973 28857 18991
rect 28875 18973 28893 18991
rect 28911 18973 28929 18991
rect 28947 18973 28965 18991
rect 28983 18973 29001 18991
rect 29019 18973 29037 18991
rect 29055 18973 29073 18991
rect 28767 18937 28785 18955
rect 28803 18937 28821 18955
rect 28839 18937 28857 18955
rect 28875 18937 28893 18955
rect 28911 18937 28929 18955
rect 28947 18937 28965 18955
rect 28983 18937 29001 18955
rect 29019 18937 29037 18955
rect 29055 18937 29073 18955
rect 28767 18901 28785 18919
rect 28803 18901 28821 18919
rect 28839 18901 28857 18919
rect 28875 18901 28893 18919
rect 28911 18901 28929 18919
rect 28947 18901 28965 18919
rect 28983 18901 29001 18919
rect 29019 18901 29037 18919
rect 29055 18901 29073 18919
rect 28767 18865 28785 18883
rect 28803 18865 28821 18883
rect 28839 18865 28857 18883
rect 28875 18865 28893 18883
rect 28911 18865 28929 18883
rect 28947 18865 28965 18883
rect 28983 18865 29001 18883
rect 29019 18865 29037 18883
rect 29055 18865 29073 18883
rect 28767 18829 28785 18847
rect 28803 18829 28821 18847
rect 28839 18829 28857 18847
rect 28875 18829 28893 18847
rect 28911 18829 28929 18847
rect 28947 18829 28965 18847
rect 28983 18829 29001 18847
rect 29019 18829 29037 18847
rect 29055 18829 29073 18847
rect 28767 18793 28785 18811
rect 28803 18793 28821 18811
rect 28839 18793 28857 18811
rect 28875 18793 28893 18811
rect 28911 18793 28929 18811
rect 28947 18793 28965 18811
rect 28983 18793 29001 18811
rect 29019 18793 29037 18811
rect 29055 18793 29073 18811
rect 28767 18757 28785 18775
rect 28803 18757 28821 18775
rect 28839 18757 28857 18775
rect 28875 18757 28893 18775
rect 28911 18757 28929 18775
rect 28947 18757 28965 18775
rect 28983 18757 29001 18775
rect 29019 18757 29037 18775
rect 29055 18757 29073 18775
rect 28767 18721 28785 18739
rect 28803 18721 28821 18739
rect 28839 18721 28857 18739
rect 28875 18721 28893 18739
rect 28911 18721 28929 18739
rect 28947 18721 28965 18739
rect 28983 18721 29001 18739
rect 29019 18721 29037 18739
rect 29055 18721 29073 18739
rect 28767 18685 28785 18703
rect 28803 18685 28821 18703
rect 28839 18685 28857 18703
rect 28875 18685 28893 18703
rect 28911 18685 28929 18703
rect 28947 18685 28965 18703
rect 28983 18685 29001 18703
rect 29019 18685 29037 18703
rect 29055 18685 29073 18703
rect 28767 18649 28785 18667
rect 28803 18649 28821 18667
rect 28839 18649 28857 18667
rect 28875 18649 28893 18667
rect 28911 18649 28929 18667
rect 28947 18649 28965 18667
rect 28983 18649 29001 18667
rect 29019 18649 29037 18667
rect 29055 18649 29073 18667
rect 28767 18613 28785 18631
rect 28803 18613 28821 18631
rect 28839 18613 28857 18631
rect 28875 18613 28893 18631
rect 28911 18613 28929 18631
rect 28947 18613 28965 18631
rect 28983 18613 29001 18631
rect 29019 18613 29037 18631
rect 29055 18613 29073 18631
rect 28767 18577 28785 18595
rect 28803 18577 28821 18595
rect 28839 18577 28857 18595
rect 28875 18577 28893 18595
rect 28911 18577 28929 18595
rect 28947 18577 28965 18595
rect 28983 18577 29001 18595
rect 29019 18577 29037 18595
rect 29055 18577 29073 18595
rect 28767 18541 28785 18559
rect 28803 18541 28821 18559
rect 28839 18541 28857 18559
rect 28875 18541 28893 18559
rect 28911 18541 28929 18559
rect 28947 18541 28965 18559
rect 28983 18541 29001 18559
rect 29019 18541 29037 18559
rect 29055 18541 29073 18559
rect 28767 18505 28785 18523
rect 28803 18505 28821 18523
rect 28839 18505 28857 18523
rect 28875 18505 28893 18523
rect 28911 18505 28929 18523
rect 28947 18505 28965 18523
rect 28983 18505 29001 18523
rect 29019 18505 29037 18523
rect 29055 18505 29073 18523
rect 28767 18469 28785 18487
rect 28803 18469 28821 18487
rect 28839 18469 28857 18487
rect 28875 18469 28893 18487
rect 28911 18469 28929 18487
rect 28947 18469 28965 18487
rect 28983 18469 29001 18487
rect 29019 18469 29037 18487
rect 29055 18469 29073 18487
rect 28767 18433 28785 18451
rect 28803 18433 28821 18451
rect 28839 18433 28857 18451
rect 28875 18433 28893 18451
rect 28911 18433 28929 18451
rect 28947 18433 28965 18451
rect 28983 18433 29001 18451
rect 29019 18433 29037 18451
rect 29055 18433 29073 18451
rect 28767 18397 28785 18415
rect 28803 18397 28821 18415
rect 28839 18397 28857 18415
rect 28875 18397 28893 18415
rect 28911 18397 28929 18415
rect 28947 18397 28965 18415
rect 28983 18397 29001 18415
rect 29019 18397 29037 18415
rect 29055 18397 29073 18415
rect 28767 18361 28785 18379
rect 28803 18361 28821 18379
rect 28839 18361 28857 18379
rect 28875 18361 28893 18379
rect 28911 18361 28929 18379
rect 28947 18361 28965 18379
rect 28983 18361 29001 18379
rect 29019 18361 29037 18379
rect 29055 18361 29073 18379
rect 28767 18325 28785 18343
rect 28803 18325 28821 18343
rect 28839 18325 28857 18343
rect 28875 18325 28893 18343
rect 28911 18325 28929 18343
rect 28947 18325 28965 18343
rect 28983 18325 29001 18343
rect 29019 18325 29037 18343
rect 29055 18325 29073 18343
rect 28767 18289 28785 18307
rect 28803 18289 28821 18307
rect 28839 18289 28857 18307
rect 28875 18289 28893 18307
rect 28911 18289 28929 18307
rect 28947 18289 28965 18307
rect 28983 18289 29001 18307
rect 29019 18289 29037 18307
rect 29055 18289 29073 18307
rect 28767 18253 28785 18271
rect 28803 18253 28821 18271
rect 28839 18253 28857 18271
rect 28875 18253 28893 18271
rect 28911 18253 28929 18271
rect 28947 18253 28965 18271
rect 28983 18253 29001 18271
rect 29019 18253 29037 18271
rect 29055 18253 29073 18271
rect 28767 18217 28785 18235
rect 28803 18217 28821 18235
rect 28839 18217 28857 18235
rect 28875 18217 28893 18235
rect 28911 18217 28929 18235
rect 28947 18217 28965 18235
rect 28983 18217 29001 18235
rect 29019 18217 29037 18235
rect 29055 18217 29073 18235
rect 28767 18181 28785 18199
rect 28803 18181 28821 18199
rect 28839 18181 28857 18199
rect 28875 18181 28893 18199
rect 28911 18181 28929 18199
rect 28947 18181 28965 18199
rect 28983 18181 29001 18199
rect 29019 18181 29037 18199
rect 29055 18181 29073 18199
rect 28767 18145 28785 18163
rect 28803 18145 28821 18163
rect 28839 18145 28857 18163
rect 28875 18145 28893 18163
rect 28911 18145 28929 18163
rect 28947 18145 28965 18163
rect 28983 18145 29001 18163
rect 29019 18145 29037 18163
rect 29055 18145 29073 18163
rect 28767 18109 28785 18127
rect 28803 18109 28821 18127
rect 28839 18109 28857 18127
rect 28875 18109 28893 18127
rect 28911 18109 28929 18127
rect 28947 18109 28965 18127
rect 28983 18109 29001 18127
rect 29019 18109 29037 18127
rect 29055 18109 29073 18127
rect 28767 18073 28785 18091
rect 28803 18073 28821 18091
rect 28839 18073 28857 18091
rect 28875 18073 28893 18091
rect 28911 18073 28929 18091
rect 28947 18073 28965 18091
rect 28983 18073 29001 18091
rect 29019 18073 29037 18091
rect 29055 18073 29073 18091
rect 8855 11547 8873 11565
rect 8891 11547 8909 11565
rect 8927 11547 8945 11565
rect 8963 11547 8981 11565
rect 8999 11547 9017 11565
rect 9035 11547 9053 11565
rect 9071 11547 9089 11565
rect 9107 11547 9125 11565
rect 8855 11511 8873 11529
rect 8891 11511 8909 11529
rect 8927 11511 8945 11529
rect 8963 11511 8981 11529
rect 8999 11511 9017 11529
rect 9035 11511 9053 11529
rect 9071 11511 9089 11529
rect 9107 11511 9125 11529
rect 8855 11475 8873 11493
rect 8891 11475 8909 11493
rect 8927 11475 8945 11493
rect 8963 11475 8981 11493
rect 8999 11475 9017 11493
rect 9035 11475 9053 11493
rect 9071 11475 9089 11493
rect 9107 11475 9125 11493
rect 8855 11439 8873 11457
rect 8891 11439 8909 11457
rect 8927 11439 8945 11457
rect 8963 11439 8981 11457
rect 8999 11439 9017 11457
rect 9035 11439 9053 11457
rect 9071 11439 9089 11457
rect 9107 11439 9125 11457
rect 8855 11403 8873 11421
rect 8891 11403 8909 11421
rect 8927 11403 8945 11421
rect 8963 11403 8981 11421
rect 8999 11403 9017 11421
rect 9035 11403 9053 11421
rect 9071 11403 9089 11421
rect 9107 11403 9125 11421
rect 8855 11367 8873 11385
rect 8891 11367 8909 11385
rect 8927 11367 8945 11385
rect 8963 11367 8981 11385
rect 8999 11367 9017 11385
rect 9035 11367 9053 11385
rect 9071 11367 9089 11385
rect 9107 11367 9125 11385
rect 8855 11331 8873 11349
rect 8891 11331 8909 11349
rect 8927 11331 8945 11349
rect 8963 11331 8981 11349
rect 8999 11331 9017 11349
rect 9035 11331 9053 11349
rect 9071 11331 9089 11349
rect 9107 11331 9125 11349
rect 8855 11295 8873 11313
rect 8891 11295 8909 11313
rect 8927 11295 8945 11313
rect 8963 11295 8981 11313
rect 8999 11295 9017 11313
rect 9035 11295 9053 11313
rect 9071 11295 9089 11313
rect 9107 11295 9125 11313
rect 8855 11259 8873 11277
rect 8891 11259 8909 11277
rect 8927 11259 8945 11277
rect 8963 11259 8981 11277
rect 8999 11259 9017 11277
rect 9035 11259 9053 11277
rect 9071 11259 9089 11277
rect 9107 11259 9125 11277
rect 8855 11223 8873 11241
rect 8891 11223 8909 11241
rect 8927 11223 8945 11241
rect 8963 11223 8981 11241
rect 8999 11223 9017 11241
rect 9035 11223 9053 11241
rect 9071 11223 9089 11241
rect 9107 11223 9125 11241
rect 8855 11187 8873 11205
rect 8891 11187 8909 11205
rect 8927 11187 8945 11205
rect 8963 11187 8981 11205
rect 8999 11187 9017 11205
rect 9035 11187 9053 11205
rect 9071 11187 9089 11205
rect 9107 11187 9125 11205
rect 8855 11151 8873 11169
rect 8891 11151 8909 11169
rect 8927 11151 8945 11169
rect 8963 11151 8981 11169
rect 8999 11151 9017 11169
rect 9035 11151 9053 11169
rect 9071 11151 9089 11169
rect 9107 11151 9125 11169
rect 8855 11115 8873 11133
rect 8891 11115 8909 11133
rect 8927 11115 8945 11133
rect 8963 11115 8981 11133
rect 8999 11115 9017 11133
rect 9035 11115 9053 11133
rect 9071 11115 9089 11133
rect 9107 11115 9125 11133
rect 8855 11079 8873 11097
rect 8891 11079 8909 11097
rect 8927 11079 8945 11097
rect 8963 11079 8981 11097
rect 8999 11079 9017 11097
rect 9035 11079 9053 11097
rect 9071 11079 9089 11097
rect 9107 11079 9125 11097
rect 8855 11043 8873 11061
rect 8891 11043 8909 11061
rect 8927 11043 8945 11061
rect 8963 11043 8981 11061
rect 8999 11043 9017 11061
rect 9035 11043 9053 11061
rect 9071 11043 9089 11061
rect 9107 11043 9125 11061
rect 8855 11007 8873 11025
rect 8891 11007 8909 11025
rect 8927 11007 8945 11025
rect 8963 11007 8981 11025
rect 8999 11007 9017 11025
rect 9035 11007 9053 11025
rect 9071 11007 9089 11025
rect 9107 11007 9125 11025
rect 8855 10971 8873 10989
rect 8891 10971 8909 10989
rect 8927 10971 8945 10989
rect 8963 10971 8981 10989
rect 8999 10971 9017 10989
rect 9035 10971 9053 10989
rect 9071 10971 9089 10989
rect 9107 10971 9125 10989
rect 8855 10935 8873 10953
rect 8891 10935 8909 10953
rect 8927 10935 8945 10953
rect 8963 10935 8981 10953
rect 8999 10935 9017 10953
rect 9035 10935 9053 10953
rect 9071 10935 9089 10953
rect 9107 10935 9125 10953
rect 8855 10899 8873 10917
rect 8891 10899 8909 10917
rect 8927 10899 8945 10917
rect 8963 10899 8981 10917
rect 8999 10899 9017 10917
rect 9035 10899 9053 10917
rect 9071 10899 9089 10917
rect 9107 10899 9125 10917
rect 8855 10863 8873 10881
rect 8891 10863 8909 10881
rect 8927 10863 8945 10881
rect 8963 10863 8981 10881
rect 8999 10863 9017 10881
rect 9035 10863 9053 10881
rect 9071 10863 9089 10881
rect 9107 10863 9125 10881
rect 8855 10827 8873 10845
rect 8891 10827 8909 10845
rect 8927 10827 8945 10845
rect 8963 10827 8981 10845
rect 8999 10827 9017 10845
rect 9035 10827 9053 10845
rect 9071 10827 9089 10845
rect 9107 10827 9125 10845
rect 8855 10791 8873 10809
rect 8891 10791 8909 10809
rect 8927 10791 8945 10809
rect 8963 10791 8981 10809
rect 8999 10791 9017 10809
rect 9035 10791 9053 10809
rect 9071 10791 9089 10809
rect 9107 10791 9125 10809
rect 8855 10755 8873 10773
rect 8891 10755 8909 10773
rect 8927 10755 8945 10773
rect 8963 10755 8981 10773
rect 8999 10755 9017 10773
rect 9035 10755 9053 10773
rect 9071 10755 9089 10773
rect 9107 10755 9125 10773
<< metal2 >>
rect 11960 28160 12040 29180
rect 11960 28147 12200 28160
rect 11960 28129 11981 28147
rect 11999 28129 12017 28147
rect 12035 28129 12053 28147
rect 12071 28129 12089 28147
rect 12107 28129 12125 28147
rect 12143 28129 12161 28147
rect 12179 28129 12200 28147
rect 11960 28111 12200 28129
rect 11960 28093 11981 28111
rect 11999 28093 12017 28111
rect 12035 28093 12053 28111
rect 12071 28093 12089 28111
rect 12107 28093 12125 28111
rect 12143 28093 12161 28111
rect 12179 28093 12200 28111
rect 11960 28080 12200 28093
rect 14660 27960 14740 29180
rect 17360 28380 17440 29180
rect 20060 28600 20140 29180
rect 20060 28520 20700 28600
rect 17360 28367 17560 28380
rect 17360 28349 17379 28367
rect 17397 28349 17415 28367
rect 17433 28349 17451 28367
rect 17469 28349 17487 28367
rect 17505 28349 17523 28367
rect 17541 28349 17560 28367
rect 17360 28331 17560 28349
rect 17360 28313 17379 28331
rect 17397 28313 17415 28331
rect 17433 28313 17451 28331
rect 17469 28313 17487 28331
rect 17505 28313 17523 28331
rect 17541 28313 17560 28331
rect 17360 28300 17560 28313
rect 19880 28367 20080 28380
rect 19880 28349 19899 28367
rect 19917 28349 19935 28367
rect 19953 28349 19971 28367
rect 19989 28349 20007 28367
rect 20025 28349 20043 28367
rect 20061 28349 20080 28367
rect 19880 28331 20080 28349
rect 19880 28313 19899 28331
rect 19917 28313 19935 28331
rect 19953 28313 19971 28331
rect 19989 28313 20007 28331
rect 20025 28313 20043 28331
rect 20061 28313 20080 28331
rect 19880 28300 20080 28313
rect 15960 28147 19620 28160
rect 15960 28129 15983 28147
rect 16001 28129 16019 28147
rect 16037 28129 16055 28147
rect 16073 28129 16091 28147
rect 16109 28129 16127 28147
rect 16145 28129 16163 28147
rect 16181 28129 16199 28147
rect 16217 28129 19620 28147
rect 15960 28111 19620 28129
rect 15960 28093 15983 28111
rect 16001 28093 16019 28111
rect 16037 28093 16055 28111
rect 16073 28093 16091 28111
rect 16109 28093 16127 28111
rect 16145 28093 16163 28111
rect 16181 28093 16199 28111
rect 16217 28093 19620 28111
rect 15960 28080 19620 28093
rect 14660 27937 14960 27960
rect 14660 27919 14675 27937
rect 14693 27919 14711 27937
rect 14729 27919 14747 27937
rect 14765 27919 14783 27937
rect 14801 27919 14819 27937
rect 14837 27919 14855 27937
rect 14873 27919 14891 27937
rect 14909 27919 14927 27937
rect 14945 27919 14960 27937
rect 14660 27901 14960 27919
rect 14660 27883 14675 27901
rect 14693 27883 14711 27901
rect 14729 27883 14747 27901
rect 14765 27883 14783 27901
rect 14801 27883 14819 27901
rect 14837 27883 14855 27901
rect 14873 27883 14891 27901
rect 14909 27883 14927 27901
rect 14945 27883 14960 27901
rect 14660 27860 14960 27883
rect 17280 27937 19120 27960
rect 17280 27919 17303 27937
rect 17321 27919 17339 27937
rect 17357 27919 17375 27937
rect 17393 27919 17411 27937
rect 17429 27919 17447 27937
rect 17465 27919 17483 27937
rect 17501 27919 17519 27937
rect 17537 27919 19120 27937
rect 17280 27901 19120 27919
rect 17280 27883 17303 27901
rect 17321 27883 17339 27901
rect 17357 27883 17375 27901
rect 17393 27883 17411 27901
rect 17429 27883 17447 27901
rect 17465 27883 17483 27901
rect 17501 27883 17519 27901
rect 17537 27883 19120 27901
rect 17280 27860 19120 27883
rect 19040 27280 19120 27860
rect 19540 27280 19620 28080
rect 20000 27280 20080 28300
rect 20620 27280 20700 28520
rect 21980 28587 22300 28600
rect 21980 28569 22005 28587
rect 22023 28569 22041 28587
rect 22059 28569 22077 28587
rect 22095 28569 22113 28587
rect 22131 28569 22149 28587
rect 22167 28569 22185 28587
rect 22203 28569 22221 28587
rect 22239 28569 22257 28587
rect 22275 28569 22300 28587
rect 21980 28551 22300 28569
rect 21980 28533 22005 28551
rect 22023 28533 22041 28551
rect 22059 28533 22077 28551
rect 22095 28533 22113 28551
rect 22131 28533 22149 28551
rect 22167 28533 22185 28551
rect 22203 28533 22221 28551
rect 22239 28533 22257 28551
rect 22275 28533 22300 28551
rect 21980 28520 22300 28533
rect 21980 27280 22060 28520
rect 22760 28320 22840 29180
rect 22120 28240 22840 28320
rect 22120 27280 22200 28240
rect 25460 28100 25540 29180
rect 28160 28600 28240 29180
rect 27980 28587 28240 28600
rect 27980 28569 27993 28587
rect 28011 28569 28029 28587
rect 28047 28569 28065 28587
rect 28083 28569 28101 28587
rect 28119 28569 28137 28587
rect 28155 28569 28173 28587
rect 28191 28569 28209 28587
rect 28227 28569 28240 28587
rect 27980 28551 28240 28569
rect 27980 28533 27993 28551
rect 28011 28533 28029 28551
rect 28047 28533 28065 28551
rect 28083 28533 28101 28551
rect 28119 28533 28137 28551
rect 28155 28533 28173 28551
rect 28191 28533 28209 28551
rect 28227 28533 28240 28551
rect 27980 28520 28240 28533
rect 22900 28087 23180 28100
rect 22900 28069 22923 28087
rect 22941 28069 22959 28087
rect 22977 28069 22995 28087
rect 23013 28069 23031 28087
rect 23049 28069 23067 28087
rect 23085 28069 23103 28087
rect 23121 28069 23139 28087
rect 23157 28069 23180 28087
rect 22900 28051 23180 28069
rect 22900 28033 22923 28051
rect 22941 28033 22959 28051
rect 22977 28033 22995 28051
rect 23013 28033 23031 28051
rect 23049 28033 23067 28051
rect 23085 28033 23103 28051
rect 23121 28033 23139 28051
rect 23157 28033 23180 28051
rect 22900 28020 23180 28033
rect 25260 28087 25540 28100
rect 25260 28069 25283 28087
rect 25301 28069 25319 28087
rect 25337 28069 25355 28087
rect 25373 28069 25391 28087
rect 25409 28069 25427 28087
rect 25445 28069 25463 28087
rect 25481 28069 25499 28087
rect 25517 28069 25540 28087
rect 25260 28051 25540 28069
rect 25260 28033 25283 28051
rect 25301 28033 25319 28051
rect 25337 28033 25355 28051
rect 25373 28033 25391 28051
rect 25409 28033 25427 28051
rect 25445 28033 25463 28051
rect 25481 28033 25499 28051
rect 25517 28033 25540 28051
rect 25260 28020 25540 28033
rect 22900 27280 22980 28020
rect 8840 27133 9140 27160
rect 8840 27115 8855 27133
rect 8873 27115 8891 27133
rect 8909 27115 8927 27133
rect 8945 27115 8963 27133
rect 8981 27115 8999 27133
rect 9017 27115 9035 27133
rect 9053 27115 9071 27133
rect 9089 27115 9107 27133
rect 9125 27115 9140 27133
rect 8840 27097 9140 27115
rect 8840 27079 8855 27097
rect 8873 27079 8891 27097
rect 8909 27079 8927 27097
rect 8945 27079 8963 27097
rect 8981 27079 8999 27097
rect 9017 27079 9035 27097
rect 9053 27079 9071 27097
rect 9089 27079 9107 27097
rect 9125 27079 9140 27097
rect 8840 27061 9140 27079
rect 8840 27043 8855 27061
rect 8873 27043 8891 27061
rect 8909 27043 8927 27061
rect 8945 27043 8963 27061
rect 8981 27043 8999 27061
rect 9017 27043 9035 27061
rect 9053 27043 9071 27061
rect 9089 27043 9107 27061
rect 9125 27043 9140 27061
rect 8840 27025 9140 27043
rect 8840 27007 8855 27025
rect 8873 27007 8891 27025
rect 8909 27007 8927 27025
rect 8945 27007 8963 27025
rect 8981 27007 8999 27025
rect 9017 27007 9035 27025
rect 9053 27007 9071 27025
rect 9089 27007 9107 27025
rect 9125 27007 9140 27025
rect 8840 26989 9140 27007
rect 8840 26971 8855 26989
rect 8873 26971 8891 26989
rect 8909 26971 8927 26989
rect 8945 26971 8963 26989
rect 8981 26971 8999 26989
rect 9017 26971 9035 26989
rect 9053 26971 9071 26989
rect 9089 26971 9107 26989
rect 9125 26971 9140 26989
rect 8840 26953 9140 26971
rect 8840 26935 8855 26953
rect 8873 26935 8891 26953
rect 8909 26935 8927 26953
rect 8945 26935 8963 26953
rect 8981 26935 8999 26953
rect 9017 26935 9035 26953
rect 9053 26935 9071 26953
rect 9089 26935 9107 26953
rect 9125 26935 9140 26953
rect 8840 26917 9140 26935
rect 8840 26899 8855 26917
rect 8873 26899 8891 26917
rect 8909 26899 8927 26917
rect 8945 26899 8963 26917
rect 8981 26899 8999 26917
rect 9017 26899 9035 26917
rect 9053 26899 9071 26917
rect 9089 26899 9107 26917
rect 9125 26899 9140 26917
rect 8840 26881 9140 26899
rect 8840 26863 8855 26881
rect 8873 26863 8891 26881
rect 8909 26863 8927 26881
rect 8945 26863 8963 26881
rect 8981 26863 8999 26881
rect 9017 26863 9035 26881
rect 9053 26863 9071 26881
rect 9089 26863 9107 26881
rect 9125 26863 9140 26881
rect 8840 26845 9140 26863
rect 8840 26827 8855 26845
rect 8873 26827 8891 26845
rect 8909 26827 8927 26845
rect 8945 26827 8963 26845
rect 8981 26827 8999 26845
rect 9017 26827 9035 26845
rect 9053 26827 9071 26845
rect 9089 26827 9107 26845
rect 9125 26827 9140 26845
rect 8840 26809 9140 26827
rect 8840 26791 8855 26809
rect 8873 26791 8891 26809
rect 8909 26791 8927 26809
rect 8945 26791 8963 26809
rect 8981 26791 8999 26809
rect 9017 26791 9035 26809
rect 9053 26791 9071 26809
rect 9089 26791 9107 26809
rect 9125 26791 9140 26809
rect 8840 26773 9140 26791
rect 8840 26755 8855 26773
rect 8873 26755 8891 26773
rect 8909 26755 8927 26773
rect 8945 26755 8963 26773
rect 8981 26755 8999 26773
rect 9017 26755 9035 26773
rect 9053 26755 9071 26773
rect 9089 26755 9107 26773
rect 9125 26755 9140 26773
rect 8840 26737 9140 26755
rect 8840 26719 8855 26737
rect 8873 26719 8891 26737
rect 8909 26719 8927 26737
rect 8945 26719 8963 26737
rect 8981 26719 8999 26737
rect 9017 26719 9035 26737
rect 9053 26719 9071 26737
rect 9089 26719 9107 26737
rect 9125 26719 9140 26737
rect 8840 26701 9140 26719
rect 8840 26683 8855 26701
rect 8873 26683 8891 26701
rect 8909 26683 8927 26701
rect 8945 26683 8963 26701
rect 8981 26683 8999 26701
rect 9017 26683 9035 26701
rect 9053 26683 9071 26701
rect 9089 26683 9107 26701
rect 9125 26683 9140 26701
rect 8840 26665 9140 26683
rect 8840 26647 8855 26665
rect 8873 26647 8891 26665
rect 8909 26647 8927 26665
rect 8945 26647 8963 26665
rect 8981 26647 8999 26665
rect 9017 26647 9035 26665
rect 9053 26647 9071 26665
rect 9089 26647 9107 26665
rect 9125 26647 9140 26665
rect 8840 26629 9140 26647
rect 8840 26611 8855 26629
rect 8873 26611 8891 26629
rect 8909 26611 8927 26629
rect 8945 26611 8963 26629
rect 8981 26611 8999 26629
rect 9017 26611 9035 26629
rect 9053 26611 9071 26629
rect 9089 26611 9107 26629
rect 9125 26611 9140 26629
rect 8840 26593 9140 26611
rect 8840 26575 8855 26593
rect 8873 26575 8891 26593
rect 8909 26575 8927 26593
rect 8945 26575 8963 26593
rect 8981 26575 8999 26593
rect 9017 26575 9035 26593
rect 9053 26575 9071 26593
rect 9089 26575 9107 26593
rect 9125 26575 9140 26593
rect 8840 26557 9140 26575
rect 8840 26539 8855 26557
rect 8873 26539 8891 26557
rect 8909 26539 8927 26557
rect 8945 26539 8963 26557
rect 8981 26539 8999 26557
rect 9017 26539 9035 26557
rect 9053 26539 9071 26557
rect 9089 26539 9107 26557
rect 9125 26539 9140 26557
rect 8840 26521 9140 26539
rect 8840 26503 8855 26521
rect 8873 26503 8891 26521
rect 8909 26503 8927 26521
rect 8945 26503 8963 26521
rect 8981 26503 8999 26521
rect 9017 26503 9035 26521
rect 9053 26503 9071 26521
rect 9089 26503 9107 26521
rect 9125 26503 9140 26521
rect 8840 26485 9140 26503
rect 8840 26467 8855 26485
rect 8873 26467 8891 26485
rect 8909 26467 8927 26485
rect 8945 26467 8963 26485
rect 8981 26467 8999 26485
rect 9017 26467 9035 26485
rect 9053 26467 9071 26485
rect 9089 26467 9107 26485
rect 9125 26467 9140 26485
rect 8840 26440 9140 26467
rect 28260 26057 29180 26080
rect 28260 26039 28273 26057
rect 28291 26039 28309 26057
rect 28327 26039 29180 26057
rect 28260 26021 29180 26039
rect 28260 26003 28273 26021
rect 28291 26003 28309 26021
rect 28327 26003 29180 26021
rect 28260 26000 29180 26003
rect 28260 25985 28340 26000
rect 28260 25967 28273 25985
rect 28291 25967 28309 25985
rect 28327 25967 28340 25985
rect 28260 25949 28340 25967
rect 28260 25931 28273 25949
rect 28291 25931 28309 25949
rect 28327 25931 28340 25949
rect 28260 25913 28340 25931
rect 28260 25895 28273 25913
rect 28291 25895 28309 25913
rect 28327 25895 28340 25913
rect 28260 25877 28340 25895
rect 28260 25859 28273 25877
rect 28291 25859 28309 25877
rect 28327 25859 28340 25877
rect 28260 25841 28340 25859
rect 28260 25823 28273 25841
rect 28291 25823 28309 25841
rect 28327 25823 28340 25841
rect 28260 25800 28340 25823
rect 28540 23367 29180 23380
rect 28540 23349 28553 23367
rect 28571 23349 28589 23367
rect 28607 23349 29180 23367
rect 8820 23319 9940 23340
rect 8820 23301 9873 23319
rect 9891 23301 9909 23319
rect 9927 23301 9940 23319
rect 8820 23283 9940 23301
rect 8820 23265 9873 23283
rect 9891 23265 9909 23283
rect 9927 23265 9940 23283
rect 8820 23260 9940 23265
rect 9860 23247 9940 23260
rect 9860 23229 9873 23247
rect 9891 23229 9909 23247
rect 9927 23229 9940 23247
rect 9860 23211 9940 23229
rect 9860 23193 9873 23211
rect 9891 23193 9909 23211
rect 9927 23193 9940 23211
rect 9860 23175 9940 23193
rect 9860 23157 9873 23175
rect 9891 23157 9909 23175
rect 9927 23157 9940 23175
rect 9860 23139 9940 23157
rect 9860 23121 9873 23139
rect 9891 23121 9909 23139
rect 9927 23121 9940 23139
rect 9860 23100 9940 23121
rect 28540 23331 29180 23349
rect 28540 23313 28553 23331
rect 28571 23313 28589 23331
rect 28607 23313 29180 23331
rect 28540 23300 29180 23313
rect 28540 23295 28620 23300
rect 28540 23277 28553 23295
rect 28571 23277 28589 23295
rect 28607 23277 28620 23295
rect 28540 23259 28620 23277
rect 28540 23241 28553 23259
rect 28571 23241 28589 23259
rect 28607 23241 28620 23259
rect 28540 23223 28620 23241
rect 28540 23205 28553 23223
rect 28571 23205 28589 23223
rect 28607 23205 28620 23223
rect 28540 23187 28620 23205
rect 28540 23169 28553 23187
rect 28571 23169 28589 23187
rect 28607 23169 28620 23187
rect 28540 23151 28620 23169
rect 28540 23133 28553 23151
rect 28571 23133 28589 23151
rect 28607 23133 28620 23151
rect 28540 23120 28620 23133
rect 28540 20885 28640 20900
rect 28540 20867 28563 20885
rect 28581 20867 28599 20885
rect 28617 20867 28640 20885
rect 28540 20849 28640 20867
rect 28540 20831 28563 20849
rect 28581 20831 28599 20849
rect 28617 20831 28640 20849
rect 28540 20813 28640 20831
rect 28540 20795 28563 20813
rect 28581 20795 28599 20813
rect 28617 20795 28640 20813
rect 9880 20751 9960 20780
rect 9880 20733 9893 20751
rect 9911 20733 9929 20751
rect 9947 20733 9960 20751
rect 9880 20715 9960 20733
rect 9880 20697 9893 20715
rect 9911 20697 9929 20715
rect 9947 20697 9960 20715
rect 9880 20679 9960 20697
rect 9880 20661 9893 20679
rect 9911 20661 9929 20679
rect 9947 20661 9960 20679
rect 9880 20643 9960 20661
rect 9880 20640 9893 20643
rect 8820 20625 9893 20640
rect 9911 20625 9929 20643
rect 9947 20625 9960 20643
rect 8820 20607 9960 20625
rect 8820 20589 9893 20607
rect 9911 20589 9929 20607
rect 9947 20589 9960 20607
rect 28540 20777 28640 20795
rect 28540 20759 28563 20777
rect 28581 20759 28599 20777
rect 28617 20759 28640 20777
rect 28540 20741 28640 20759
rect 28540 20723 28563 20741
rect 28581 20723 28599 20741
rect 28617 20723 28640 20741
rect 28540 20705 28640 20723
rect 28540 20687 28563 20705
rect 28581 20687 28599 20705
rect 28617 20687 28640 20705
rect 28540 20680 28640 20687
rect 28540 20669 29180 20680
rect 28540 20651 28563 20669
rect 28581 20651 28599 20669
rect 28617 20651 29180 20669
rect 28540 20633 29180 20651
rect 28540 20615 28563 20633
rect 28581 20615 28599 20633
rect 28617 20615 29180 20633
rect 28540 20600 29180 20615
rect 8820 20560 9960 20589
rect 28740 19927 29180 19940
rect 28740 19909 28767 19927
rect 28785 19909 28803 19927
rect 28821 19909 28839 19927
rect 28857 19909 28875 19927
rect 28893 19909 28911 19927
rect 28929 19909 28947 19927
rect 28965 19909 28983 19927
rect 29001 19909 29019 19927
rect 29037 19909 29055 19927
rect 29073 19909 29180 19927
rect 28740 19891 29180 19909
rect 28740 19873 28767 19891
rect 28785 19873 28803 19891
rect 28821 19873 28839 19891
rect 28857 19873 28875 19891
rect 28893 19873 28911 19891
rect 28929 19873 28947 19891
rect 28965 19873 28983 19891
rect 29001 19873 29019 19891
rect 29037 19873 29055 19891
rect 29073 19873 29180 19891
rect 28740 19855 29180 19873
rect 28740 19837 28767 19855
rect 28785 19837 28803 19855
rect 28821 19837 28839 19855
rect 28857 19837 28875 19855
rect 28893 19837 28911 19855
rect 28929 19837 28947 19855
rect 28965 19837 28983 19855
rect 29001 19837 29019 19855
rect 29037 19837 29055 19855
rect 29073 19837 29180 19855
rect 28740 19819 29180 19837
rect 28740 19801 28767 19819
rect 28785 19801 28803 19819
rect 28821 19801 28839 19819
rect 28857 19801 28875 19819
rect 28893 19801 28911 19819
rect 28929 19801 28947 19819
rect 28965 19801 28983 19819
rect 29001 19801 29019 19819
rect 29037 19801 29055 19819
rect 29073 19801 29180 19819
rect 28740 19783 29180 19801
rect 28740 19765 28767 19783
rect 28785 19765 28803 19783
rect 28821 19765 28839 19783
rect 28857 19765 28875 19783
rect 28893 19765 28911 19783
rect 28929 19765 28947 19783
rect 28965 19765 28983 19783
rect 29001 19765 29019 19783
rect 29037 19765 29055 19783
rect 29073 19765 29180 19783
rect 28740 19747 29180 19765
rect 28740 19729 28767 19747
rect 28785 19729 28803 19747
rect 28821 19729 28839 19747
rect 28857 19729 28875 19747
rect 28893 19729 28911 19747
rect 28929 19729 28947 19747
rect 28965 19729 28983 19747
rect 29001 19729 29019 19747
rect 29037 19729 29055 19747
rect 29073 19729 29180 19747
rect 28740 19711 29180 19729
rect 28740 19693 28767 19711
rect 28785 19693 28803 19711
rect 28821 19693 28839 19711
rect 28857 19693 28875 19711
rect 28893 19693 28911 19711
rect 28929 19693 28947 19711
rect 28965 19693 28983 19711
rect 29001 19693 29019 19711
rect 29037 19693 29055 19711
rect 29073 19693 29180 19711
rect 28740 19675 29180 19693
rect 28740 19657 28767 19675
rect 28785 19657 28803 19675
rect 28821 19657 28839 19675
rect 28857 19657 28875 19675
rect 28893 19657 28911 19675
rect 28929 19657 28947 19675
rect 28965 19657 28983 19675
rect 29001 19657 29019 19675
rect 29037 19657 29055 19675
rect 29073 19657 29180 19675
rect 28740 19639 29180 19657
rect 28740 19621 28767 19639
rect 28785 19621 28803 19639
rect 28821 19621 28839 19639
rect 28857 19621 28875 19639
rect 28893 19621 28911 19639
rect 28929 19621 28947 19639
rect 28965 19621 28983 19639
rect 29001 19621 29019 19639
rect 29037 19621 29055 19639
rect 29073 19621 29180 19639
rect 28740 19603 29180 19621
rect 28740 19585 28767 19603
rect 28785 19585 28803 19603
rect 28821 19585 28839 19603
rect 28857 19585 28875 19603
rect 28893 19585 28911 19603
rect 28929 19585 28947 19603
rect 28965 19585 28983 19603
rect 29001 19585 29019 19603
rect 29037 19585 29055 19603
rect 29073 19585 29180 19603
rect 28740 19567 29180 19585
rect 28740 19549 28767 19567
rect 28785 19549 28803 19567
rect 28821 19549 28839 19567
rect 28857 19549 28875 19567
rect 28893 19549 28911 19567
rect 28929 19549 28947 19567
rect 28965 19549 28983 19567
rect 29001 19549 29019 19567
rect 29037 19549 29055 19567
rect 29073 19549 29180 19567
rect 28740 19531 29180 19549
rect 28740 19513 28767 19531
rect 28785 19513 28803 19531
rect 28821 19513 28839 19531
rect 28857 19513 28875 19531
rect 28893 19513 28911 19531
rect 28929 19513 28947 19531
rect 28965 19513 28983 19531
rect 29001 19513 29019 19531
rect 29037 19513 29055 19531
rect 29073 19513 29180 19531
rect 28740 19495 29180 19513
rect 28740 19477 28767 19495
rect 28785 19477 28803 19495
rect 28821 19477 28839 19495
rect 28857 19477 28875 19495
rect 28893 19477 28911 19495
rect 28929 19477 28947 19495
rect 28965 19477 28983 19495
rect 29001 19477 29019 19495
rect 29037 19477 29055 19495
rect 29073 19477 29180 19495
rect 28740 19459 29180 19477
rect 28740 19441 28767 19459
rect 28785 19441 28803 19459
rect 28821 19441 28839 19459
rect 28857 19441 28875 19459
rect 28893 19441 28911 19459
rect 28929 19441 28947 19459
rect 28965 19441 28983 19459
rect 29001 19441 29019 19459
rect 29037 19441 29055 19459
rect 29073 19441 29180 19459
rect 28740 19423 29180 19441
rect 28740 19405 28767 19423
rect 28785 19405 28803 19423
rect 28821 19405 28839 19423
rect 28857 19405 28875 19423
rect 28893 19405 28911 19423
rect 28929 19405 28947 19423
rect 28965 19405 28983 19423
rect 29001 19405 29019 19423
rect 29037 19405 29055 19423
rect 29073 19405 29180 19423
rect 28740 19387 29180 19405
rect 28740 19369 28767 19387
rect 28785 19369 28803 19387
rect 28821 19369 28839 19387
rect 28857 19369 28875 19387
rect 28893 19369 28911 19387
rect 28929 19369 28947 19387
rect 28965 19369 28983 19387
rect 29001 19369 29019 19387
rect 29037 19369 29055 19387
rect 29073 19369 29180 19387
rect 28740 19351 29180 19369
rect 28740 19333 28767 19351
rect 28785 19333 28803 19351
rect 28821 19333 28839 19351
rect 28857 19333 28875 19351
rect 28893 19333 28911 19351
rect 28929 19333 28947 19351
rect 28965 19333 28983 19351
rect 29001 19333 29019 19351
rect 29037 19333 29055 19351
rect 29073 19333 29180 19351
rect 28740 19315 29180 19333
rect 28740 19297 28767 19315
rect 28785 19297 28803 19315
rect 28821 19297 28839 19315
rect 28857 19297 28875 19315
rect 28893 19297 28911 19315
rect 28929 19297 28947 19315
rect 28965 19297 28983 19315
rect 29001 19297 29019 19315
rect 29037 19297 29055 19315
rect 29073 19297 29180 19315
rect 28740 19279 29180 19297
rect 28740 19261 28767 19279
rect 28785 19261 28803 19279
rect 28821 19261 28839 19279
rect 28857 19261 28875 19279
rect 28893 19261 28911 19279
rect 28929 19261 28947 19279
rect 28965 19261 28983 19279
rect 29001 19261 29019 19279
rect 29037 19261 29055 19279
rect 29073 19261 29180 19279
rect 28740 19243 29180 19261
rect 28740 19225 28767 19243
rect 28785 19225 28803 19243
rect 28821 19225 28839 19243
rect 28857 19225 28875 19243
rect 28893 19225 28911 19243
rect 28929 19225 28947 19243
rect 28965 19225 28983 19243
rect 29001 19225 29019 19243
rect 29037 19225 29055 19243
rect 29073 19225 29180 19243
rect 28740 19207 29180 19225
rect 28740 19189 28767 19207
rect 28785 19189 28803 19207
rect 28821 19189 28839 19207
rect 28857 19189 28875 19207
rect 28893 19189 28911 19207
rect 28929 19189 28947 19207
rect 28965 19189 28983 19207
rect 29001 19189 29019 19207
rect 29037 19189 29055 19207
rect 29073 19189 29180 19207
rect 28740 19171 29180 19189
rect 28740 19153 28767 19171
rect 28785 19153 28803 19171
rect 28821 19153 28839 19171
rect 28857 19153 28875 19171
rect 28893 19153 28911 19171
rect 28929 19153 28947 19171
rect 28965 19153 28983 19171
rect 29001 19153 29019 19171
rect 29037 19153 29055 19171
rect 29073 19153 29180 19171
rect 28740 19135 29180 19153
rect 28740 19117 28767 19135
rect 28785 19117 28803 19135
rect 28821 19117 28839 19135
rect 28857 19117 28875 19135
rect 28893 19117 28911 19135
rect 28929 19117 28947 19135
rect 28965 19117 28983 19135
rect 29001 19117 29019 19135
rect 29037 19117 29055 19135
rect 29073 19117 29180 19135
rect 28740 19099 29180 19117
rect 28740 19081 28767 19099
rect 28785 19081 28803 19099
rect 28821 19081 28839 19099
rect 28857 19081 28875 19099
rect 28893 19081 28911 19099
rect 28929 19081 28947 19099
rect 28965 19081 28983 19099
rect 29001 19081 29019 19099
rect 29037 19081 29055 19099
rect 29073 19081 29180 19099
rect 28740 19063 29180 19081
rect 28740 19045 28767 19063
rect 28785 19045 28803 19063
rect 28821 19045 28839 19063
rect 28857 19045 28875 19063
rect 28893 19045 28911 19063
rect 28929 19045 28947 19063
rect 28965 19045 28983 19063
rect 29001 19045 29019 19063
rect 29037 19045 29055 19063
rect 29073 19045 29180 19063
rect 28740 19027 29180 19045
rect 28740 19009 28767 19027
rect 28785 19009 28803 19027
rect 28821 19009 28839 19027
rect 28857 19009 28875 19027
rect 28893 19009 28911 19027
rect 28929 19009 28947 19027
rect 28965 19009 28983 19027
rect 29001 19009 29019 19027
rect 29037 19009 29055 19027
rect 29073 19009 29180 19027
rect 28740 18991 29180 19009
rect 28740 18973 28767 18991
rect 28785 18973 28803 18991
rect 28821 18973 28839 18991
rect 28857 18973 28875 18991
rect 28893 18973 28911 18991
rect 28929 18973 28947 18991
rect 28965 18973 28983 18991
rect 29001 18973 29019 18991
rect 29037 18973 29055 18991
rect 29073 18973 29180 18991
rect 28740 18955 29180 18973
rect 28740 18937 28767 18955
rect 28785 18937 28803 18955
rect 28821 18937 28839 18955
rect 28857 18937 28875 18955
rect 28893 18937 28911 18955
rect 28929 18937 28947 18955
rect 28965 18937 28983 18955
rect 29001 18937 29019 18955
rect 29037 18937 29055 18955
rect 29073 18937 29180 18955
rect 28740 18919 29180 18937
rect 28740 18901 28767 18919
rect 28785 18901 28803 18919
rect 28821 18901 28839 18919
rect 28857 18901 28875 18919
rect 28893 18901 28911 18919
rect 28929 18901 28947 18919
rect 28965 18901 28983 18919
rect 29001 18901 29019 18919
rect 29037 18901 29055 18919
rect 29073 18901 29180 18919
rect 28740 18883 29180 18901
rect 28740 18865 28767 18883
rect 28785 18865 28803 18883
rect 28821 18865 28839 18883
rect 28857 18865 28875 18883
rect 28893 18865 28911 18883
rect 28929 18865 28947 18883
rect 28965 18865 28983 18883
rect 29001 18865 29019 18883
rect 29037 18865 29055 18883
rect 29073 18865 29180 18883
rect 28740 18847 29180 18865
rect 28740 18829 28767 18847
rect 28785 18829 28803 18847
rect 28821 18829 28839 18847
rect 28857 18829 28875 18847
rect 28893 18829 28911 18847
rect 28929 18829 28947 18847
rect 28965 18829 28983 18847
rect 29001 18829 29019 18847
rect 29037 18829 29055 18847
rect 29073 18829 29180 18847
rect 28740 18811 29180 18829
rect 28740 18793 28767 18811
rect 28785 18793 28803 18811
rect 28821 18793 28839 18811
rect 28857 18793 28875 18811
rect 28893 18793 28911 18811
rect 28929 18793 28947 18811
rect 28965 18793 28983 18811
rect 29001 18793 29019 18811
rect 29037 18793 29055 18811
rect 29073 18793 29180 18811
rect 28740 18775 29180 18793
rect 28740 18757 28767 18775
rect 28785 18757 28803 18775
rect 28821 18757 28839 18775
rect 28857 18757 28875 18775
rect 28893 18757 28911 18775
rect 28929 18757 28947 18775
rect 28965 18757 28983 18775
rect 29001 18757 29019 18775
rect 29037 18757 29055 18775
rect 29073 18757 29180 18775
rect 28740 18739 29180 18757
rect 28740 18721 28767 18739
rect 28785 18721 28803 18739
rect 28821 18721 28839 18739
rect 28857 18721 28875 18739
rect 28893 18721 28911 18739
rect 28929 18721 28947 18739
rect 28965 18721 28983 18739
rect 29001 18721 29019 18739
rect 29037 18721 29055 18739
rect 29073 18721 29180 18739
rect 28740 18703 29180 18721
rect 28740 18685 28767 18703
rect 28785 18685 28803 18703
rect 28821 18685 28839 18703
rect 28857 18685 28875 18703
rect 28893 18685 28911 18703
rect 28929 18685 28947 18703
rect 28965 18685 28983 18703
rect 29001 18685 29019 18703
rect 29037 18685 29055 18703
rect 29073 18685 29180 18703
rect 28740 18667 29180 18685
rect 28740 18649 28767 18667
rect 28785 18649 28803 18667
rect 28821 18649 28839 18667
rect 28857 18649 28875 18667
rect 28893 18649 28911 18667
rect 28929 18649 28947 18667
rect 28965 18649 28983 18667
rect 29001 18649 29019 18667
rect 29037 18649 29055 18667
rect 29073 18649 29180 18667
rect 28740 18631 29180 18649
rect 28740 18613 28767 18631
rect 28785 18613 28803 18631
rect 28821 18613 28839 18631
rect 28857 18613 28875 18631
rect 28893 18613 28911 18631
rect 28929 18613 28947 18631
rect 28965 18613 28983 18631
rect 29001 18613 29019 18631
rect 29037 18613 29055 18631
rect 29073 18613 29180 18631
rect 28740 18595 29180 18613
rect 28740 18577 28767 18595
rect 28785 18577 28803 18595
rect 28821 18577 28839 18595
rect 28857 18577 28875 18595
rect 28893 18577 28911 18595
rect 28929 18577 28947 18595
rect 28965 18577 28983 18595
rect 29001 18577 29019 18595
rect 29037 18577 29055 18595
rect 29073 18577 29180 18595
rect 28740 18559 29180 18577
rect 28740 18541 28767 18559
rect 28785 18541 28803 18559
rect 28821 18541 28839 18559
rect 28857 18541 28875 18559
rect 28893 18541 28911 18559
rect 28929 18541 28947 18559
rect 28965 18541 28983 18559
rect 29001 18541 29019 18559
rect 29037 18541 29055 18559
rect 29073 18541 29180 18559
rect 28740 18523 29180 18541
rect 28740 18505 28767 18523
rect 28785 18505 28803 18523
rect 28821 18505 28839 18523
rect 28857 18505 28875 18523
rect 28893 18505 28911 18523
rect 28929 18505 28947 18523
rect 28965 18505 28983 18523
rect 29001 18505 29019 18523
rect 29037 18505 29055 18523
rect 29073 18505 29180 18523
rect 28740 18487 29180 18505
rect 28740 18469 28767 18487
rect 28785 18469 28803 18487
rect 28821 18469 28839 18487
rect 28857 18469 28875 18487
rect 28893 18469 28911 18487
rect 28929 18469 28947 18487
rect 28965 18469 28983 18487
rect 29001 18469 29019 18487
rect 29037 18469 29055 18487
rect 29073 18469 29180 18487
rect 28740 18451 29180 18469
rect 28740 18433 28767 18451
rect 28785 18433 28803 18451
rect 28821 18433 28839 18451
rect 28857 18433 28875 18451
rect 28893 18433 28911 18451
rect 28929 18433 28947 18451
rect 28965 18433 28983 18451
rect 29001 18433 29019 18451
rect 29037 18433 29055 18451
rect 29073 18433 29180 18451
rect 28740 18415 29180 18433
rect 28740 18397 28767 18415
rect 28785 18397 28803 18415
rect 28821 18397 28839 18415
rect 28857 18397 28875 18415
rect 28893 18397 28911 18415
rect 28929 18397 28947 18415
rect 28965 18397 28983 18415
rect 29001 18397 29019 18415
rect 29037 18397 29055 18415
rect 29073 18397 29180 18415
rect 28740 18379 29180 18397
rect 28740 18361 28767 18379
rect 28785 18361 28803 18379
rect 28821 18361 28839 18379
rect 28857 18361 28875 18379
rect 28893 18361 28911 18379
rect 28929 18361 28947 18379
rect 28965 18361 28983 18379
rect 29001 18361 29019 18379
rect 29037 18361 29055 18379
rect 29073 18361 29180 18379
rect 28740 18343 29180 18361
rect 28740 18325 28767 18343
rect 28785 18325 28803 18343
rect 28821 18325 28839 18343
rect 28857 18325 28875 18343
rect 28893 18325 28911 18343
rect 28929 18325 28947 18343
rect 28965 18325 28983 18343
rect 29001 18325 29019 18343
rect 29037 18325 29055 18343
rect 29073 18325 29180 18343
rect 28740 18307 29180 18325
rect 28740 18289 28767 18307
rect 28785 18289 28803 18307
rect 28821 18289 28839 18307
rect 28857 18289 28875 18307
rect 28893 18289 28911 18307
rect 28929 18289 28947 18307
rect 28965 18289 28983 18307
rect 29001 18289 29019 18307
rect 29037 18289 29055 18307
rect 29073 18289 29180 18307
rect 28740 18271 29180 18289
rect 28740 18253 28767 18271
rect 28785 18253 28803 18271
rect 28821 18253 28839 18271
rect 28857 18253 28875 18271
rect 28893 18253 28911 18271
rect 28929 18253 28947 18271
rect 28965 18253 28983 18271
rect 29001 18253 29019 18271
rect 29037 18253 29055 18271
rect 29073 18253 29180 18271
rect 28740 18235 29180 18253
rect 28740 18217 28767 18235
rect 28785 18217 28803 18235
rect 28821 18217 28839 18235
rect 28857 18217 28875 18235
rect 28893 18217 28911 18235
rect 28929 18217 28947 18235
rect 28965 18217 28983 18235
rect 29001 18217 29019 18235
rect 29037 18217 29055 18235
rect 29073 18217 29180 18235
rect 28740 18199 29180 18217
rect 28740 18181 28767 18199
rect 28785 18181 28803 18199
rect 28821 18181 28839 18199
rect 28857 18181 28875 18199
rect 28893 18181 28911 18199
rect 28929 18181 28947 18199
rect 28965 18181 28983 18199
rect 29001 18181 29019 18199
rect 29037 18181 29055 18199
rect 29073 18181 29180 18199
rect 28740 18163 29180 18181
rect 28740 18145 28767 18163
rect 28785 18145 28803 18163
rect 28821 18145 28839 18163
rect 28857 18145 28875 18163
rect 28893 18145 28911 18163
rect 28929 18145 28947 18163
rect 28965 18145 28983 18163
rect 29001 18145 29019 18163
rect 29037 18145 29055 18163
rect 29073 18145 29180 18163
rect 28740 18127 29180 18145
rect 28740 18109 28767 18127
rect 28785 18109 28803 18127
rect 28821 18109 28839 18127
rect 28857 18109 28875 18127
rect 28893 18109 28911 18127
rect 28929 18109 28947 18127
rect 28965 18109 28983 18127
rect 29001 18109 29019 18127
rect 29037 18109 29055 18127
rect 29073 18109 29180 18127
rect 28740 18091 29180 18109
rect 9400 18051 9480 18080
rect 28740 18073 28767 18091
rect 28785 18073 28803 18091
rect 28821 18073 28839 18091
rect 28857 18073 28875 18091
rect 28893 18073 28911 18091
rect 28929 18073 28947 18091
rect 28965 18073 28983 18091
rect 29001 18073 29019 18091
rect 29037 18073 29055 18091
rect 29073 18073 29180 18091
rect 28740 18060 29180 18073
rect 9400 18033 9413 18051
rect 9431 18033 9449 18051
rect 9467 18033 9480 18051
rect 9400 18015 9480 18033
rect 9400 17997 9413 18015
rect 9431 17997 9449 18015
rect 9467 17997 9480 18015
rect 9400 17979 9480 17997
rect 9400 17961 9413 17979
rect 9431 17961 9449 17979
rect 9467 17961 9480 17979
rect 9400 17943 9480 17961
rect 9400 17940 9413 17943
rect 8820 17925 9413 17940
rect 9431 17925 9449 17943
rect 9467 17925 9480 17943
rect 8820 17907 9480 17925
rect 8820 17889 9413 17907
rect 9431 17889 9449 17907
rect 9467 17889 9480 17907
rect 8820 17860 9480 17889
rect 9620 17651 9700 17680
rect 9620 17633 9633 17651
rect 9651 17633 9669 17651
rect 9687 17633 9700 17651
rect 9620 17615 9700 17633
rect 9620 17597 9633 17615
rect 9651 17597 9669 17615
rect 9687 17597 9700 17615
rect 9620 17579 9700 17597
rect 9620 17561 9633 17579
rect 9651 17561 9669 17579
rect 9687 17561 9700 17579
rect 9620 17543 9700 17561
rect 9620 17525 9633 17543
rect 9651 17525 9669 17543
rect 9687 17525 9700 17543
rect 9620 17507 9700 17525
rect 9620 17489 9633 17507
rect 9651 17489 9669 17507
rect 9687 17489 9700 17507
rect 9620 15240 9700 17489
rect 8820 15160 9700 15240
rect 28380 15447 28460 15460
rect 28380 15429 28393 15447
rect 28411 15429 28429 15447
rect 28447 15429 28460 15447
rect 28380 15411 28460 15429
rect 28380 15393 28393 15411
rect 28411 15393 28429 15411
rect 28447 15393 28460 15411
rect 28380 15375 28460 15393
rect 28380 15357 28393 15375
rect 28411 15357 28429 15375
rect 28447 15357 28460 15375
rect 28380 15339 28460 15357
rect 28380 15321 28393 15339
rect 28411 15321 28429 15339
rect 28447 15321 28460 15339
rect 28380 15303 28460 15321
rect 28380 15285 28393 15303
rect 28411 15285 28429 15303
rect 28447 15285 28460 15303
rect 28380 15280 28460 15285
rect 28380 15267 29180 15280
rect 28380 15249 28393 15267
rect 28411 15249 28429 15267
rect 28447 15249 29180 15267
rect 28380 15231 29180 15249
rect 28380 15213 28393 15231
rect 28411 15213 28429 15231
rect 28447 15213 29180 15231
rect 28380 15200 29180 15213
rect 9880 14437 9960 14460
rect 9880 14419 9893 14437
rect 9911 14419 9929 14437
rect 9947 14419 9960 14437
rect 9880 14401 9960 14419
rect 9880 14383 9893 14401
rect 9911 14383 9929 14401
rect 9947 14383 9960 14401
rect 9880 14365 9960 14383
rect 9880 14347 9893 14365
rect 9911 14347 9929 14365
rect 9947 14347 9960 14365
rect 9880 14329 9960 14347
rect 9880 14311 9893 14329
rect 9911 14311 9929 14329
rect 9947 14311 9960 14329
rect 9880 14293 9960 14311
rect 9880 14275 9893 14293
rect 9911 14275 9929 14293
rect 9947 14275 9960 14293
rect 9880 14257 9960 14275
rect 9880 14239 9893 14257
rect 9911 14239 9929 14257
rect 9947 14239 9960 14257
rect 9880 14221 9960 14239
rect 9880 14203 9893 14221
rect 9911 14203 9929 14221
rect 9947 14203 9960 14221
rect 9880 12540 9960 14203
rect 8820 12460 9960 12540
rect 28160 12747 28240 12760
rect 28160 12729 28173 12747
rect 28191 12729 28209 12747
rect 28227 12729 28240 12747
rect 28160 12711 28240 12729
rect 28160 12693 28173 12711
rect 28191 12693 28209 12711
rect 28227 12693 28240 12711
rect 28160 12675 28240 12693
rect 28160 12657 28173 12675
rect 28191 12657 28209 12675
rect 28227 12657 28240 12675
rect 28160 12639 28240 12657
rect 28160 12621 28173 12639
rect 28191 12621 28209 12639
rect 28227 12621 28240 12639
rect 28160 12603 28240 12621
rect 28160 12585 28173 12603
rect 28191 12585 28209 12603
rect 28227 12585 28240 12603
rect 28160 12580 28240 12585
rect 28160 12567 29180 12580
rect 28160 12549 28173 12567
rect 28191 12549 28209 12567
rect 28227 12549 29180 12567
rect 28160 12531 29180 12549
rect 28160 12513 28173 12531
rect 28191 12513 28209 12531
rect 28227 12513 29180 12531
rect 28160 12500 29180 12513
rect 8820 11565 9140 11580
rect 8820 11547 8855 11565
rect 8873 11547 8891 11565
rect 8909 11547 8927 11565
rect 8945 11547 8963 11565
rect 8981 11547 8999 11565
rect 9017 11547 9035 11565
rect 9053 11547 9071 11565
rect 9089 11547 9107 11565
rect 9125 11547 9140 11565
rect 8820 11529 9140 11547
rect 8820 11511 8855 11529
rect 8873 11511 8891 11529
rect 8909 11511 8927 11529
rect 8945 11511 8963 11529
rect 8981 11511 8999 11529
rect 9017 11511 9035 11529
rect 9053 11511 9071 11529
rect 9089 11511 9107 11529
rect 9125 11511 9140 11529
rect 8820 11493 9140 11511
rect 8820 11475 8855 11493
rect 8873 11475 8891 11493
rect 8909 11475 8927 11493
rect 8945 11475 8963 11493
rect 8981 11475 8999 11493
rect 9017 11475 9035 11493
rect 9053 11475 9071 11493
rect 9089 11475 9107 11493
rect 9125 11475 9140 11493
rect 8820 11457 9140 11475
rect 8820 11439 8855 11457
rect 8873 11439 8891 11457
rect 8909 11439 8927 11457
rect 8945 11439 8963 11457
rect 8981 11439 8999 11457
rect 9017 11439 9035 11457
rect 9053 11439 9071 11457
rect 9089 11439 9107 11457
rect 9125 11439 9140 11457
rect 8820 11421 9140 11439
rect 8820 11403 8855 11421
rect 8873 11403 8891 11421
rect 8909 11403 8927 11421
rect 8945 11403 8963 11421
rect 8981 11403 8999 11421
rect 9017 11403 9035 11421
rect 9053 11403 9071 11421
rect 9089 11403 9107 11421
rect 9125 11403 9140 11421
rect 8820 11385 9140 11403
rect 8820 11367 8855 11385
rect 8873 11367 8891 11385
rect 8909 11367 8927 11385
rect 8945 11367 8963 11385
rect 8981 11367 8999 11385
rect 9017 11367 9035 11385
rect 9053 11367 9071 11385
rect 9089 11367 9107 11385
rect 9125 11367 9140 11385
rect 8820 11349 9140 11367
rect 8820 11331 8855 11349
rect 8873 11331 8891 11349
rect 8909 11331 8927 11349
rect 8945 11331 8963 11349
rect 8981 11331 8999 11349
rect 9017 11331 9035 11349
rect 9053 11331 9071 11349
rect 9089 11331 9107 11349
rect 9125 11331 9140 11349
rect 8820 11313 9140 11331
rect 8820 11295 8855 11313
rect 8873 11295 8891 11313
rect 8909 11295 8927 11313
rect 8945 11295 8963 11313
rect 8981 11295 8999 11313
rect 9017 11295 9035 11313
rect 9053 11295 9071 11313
rect 9089 11295 9107 11313
rect 9125 11295 9140 11313
rect 8820 11277 9140 11295
rect 8820 11259 8855 11277
rect 8873 11259 8891 11277
rect 8909 11259 8927 11277
rect 8945 11259 8963 11277
rect 8981 11259 8999 11277
rect 9017 11259 9035 11277
rect 9053 11259 9071 11277
rect 9089 11259 9107 11277
rect 9125 11259 9140 11277
rect 8820 11241 9140 11259
rect 8820 11223 8855 11241
rect 8873 11223 8891 11241
rect 8909 11223 8927 11241
rect 8945 11223 8963 11241
rect 8981 11223 8999 11241
rect 9017 11223 9035 11241
rect 9053 11223 9071 11241
rect 9089 11223 9107 11241
rect 9125 11223 9140 11241
rect 8820 11205 9140 11223
rect 8820 11187 8855 11205
rect 8873 11187 8891 11205
rect 8909 11187 8927 11205
rect 8945 11187 8963 11205
rect 8981 11187 8999 11205
rect 9017 11187 9035 11205
rect 9053 11187 9071 11205
rect 9089 11187 9107 11205
rect 9125 11187 9140 11205
rect 8820 11169 9140 11187
rect 8820 11151 8855 11169
rect 8873 11151 8891 11169
rect 8909 11151 8927 11169
rect 8945 11151 8963 11169
rect 8981 11151 8999 11169
rect 9017 11151 9035 11169
rect 9053 11151 9071 11169
rect 9089 11151 9107 11169
rect 9125 11151 9140 11169
rect 8820 11133 9140 11151
rect 8820 11115 8855 11133
rect 8873 11115 8891 11133
rect 8909 11115 8927 11133
rect 8945 11115 8963 11133
rect 8981 11115 8999 11133
rect 9017 11115 9035 11133
rect 9053 11115 9071 11133
rect 9089 11115 9107 11133
rect 9125 11115 9140 11133
rect 8820 11097 9140 11115
rect 8820 11079 8855 11097
rect 8873 11079 8891 11097
rect 8909 11079 8927 11097
rect 8945 11079 8963 11097
rect 8981 11079 8999 11097
rect 9017 11079 9035 11097
rect 9053 11079 9071 11097
rect 9089 11079 9107 11097
rect 9125 11079 9140 11097
rect 8820 11061 9140 11079
rect 8820 11043 8855 11061
rect 8873 11043 8891 11061
rect 8909 11043 8927 11061
rect 8945 11043 8963 11061
rect 8981 11043 8999 11061
rect 9017 11043 9035 11061
rect 9053 11043 9071 11061
rect 9089 11043 9107 11061
rect 9125 11043 9140 11061
rect 8820 11025 9140 11043
rect 8820 11007 8855 11025
rect 8873 11007 8891 11025
rect 8909 11007 8927 11025
rect 8945 11007 8963 11025
rect 8981 11007 8999 11025
rect 9017 11007 9035 11025
rect 9053 11007 9071 11025
rect 9089 11007 9107 11025
rect 9125 11007 9140 11025
rect 8820 10989 9140 11007
rect 8820 10971 8855 10989
rect 8873 10971 8891 10989
rect 8909 10971 8927 10989
rect 8945 10971 8963 10989
rect 8981 10971 8999 10989
rect 9017 10971 9035 10989
rect 9053 10971 9071 10989
rect 9089 10971 9107 10989
rect 9125 10971 9140 10989
rect 8820 10953 9140 10971
rect 8820 10935 8855 10953
rect 8873 10935 8891 10953
rect 8909 10935 8927 10953
rect 8945 10935 8963 10953
rect 8981 10935 8999 10953
rect 9017 10935 9035 10953
rect 9053 10935 9071 10953
rect 9089 10935 9107 10953
rect 9125 10935 9140 10953
rect 8820 10917 9140 10935
rect 8820 10899 8855 10917
rect 8873 10899 8891 10917
rect 8909 10899 8927 10917
rect 8945 10899 8963 10917
rect 8981 10899 8999 10917
rect 9017 10899 9035 10917
rect 9053 10899 9071 10917
rect 9089 10899 9107 10917
rect 9125 10899 9140 10917
rect 8820 10881 9140 10899
rect 8820 10863 8855 10881
rect 8873 10863 8891 10881
rect 8909 10863 8927 10881
rect 8945 10863 8963 10881
rect 8981 10863 8999 10881
rect 9017 10863 9035 10881
rect 9053 10863 9071 10881
rect 9089 10863 9107 10881
rect 9125 10863 9140 10881
rect 8820 10845 9140 10863
rect 8820 10827 8855 10845
rect 8873 10827 8891 10845
rect 8909 10827 8927 10845
rect 8945 10827 8963 10845
rect 8981 10827 8999 10845
rect 9017 10827 9035 10845
rect 9053 10827 9071 10845
rect 9089 10827 9107 10845
rect 9125 10827 9140 10845
rect 8820 10809 9140 10827
rect 8820 10791 8855 10809
rect 8873 10791 8891 10809
rect 8909 10791 8927 10809
rect 8945 10791 8963 10809
rect 8981 10791 8999 10809
rect 9017 10791 9035 10809
rect 9053 10791 9071 10809
rect 9089 10791 9107 10809
rect 9125 10791 9140 10809
rect 8820 10773 9140 10791
rect 8820 10755 8855 10773
rect 8873 10755 8891 10773
rect 8909 10755 8927 10773
rect 8945 10755 8963 10773
rect 8981 10755 8999 10773
rect 9017 10755 9035 10773
rect 9053 10755 9071 10773
rect 9089 10755 9107 10773
rect 9125 10755 9140 10773
rect 8820 10740 9140 10755
rect 17560 10360 17620 10680
rect 11960 10347 12180 10360
rect 11960 10329 11989 10347
rect 12007 10329 12025 10347
rect 12043 10329 12061 10347
rect 12079 10329 12097 10347
rect 12115 10329 12133 10347
rect 12151 10329 12180 10347
rect 11960 10311 12180 10329
rect 11960 10293 11989 10311
rect 12007 10293 12025 10311
rect 12043 10293 12061 10311
rect 12079 10293 12097 10311
rect 12115 10293 12133 10311
rect 12151 10293 12180 10311
rect 11960 10280 12180 10293
rect 15040 10347 17620 10360
rect 15040 10329 15069 10347
rect 15087 10329 15105 10347
rect 15123 10329 15141 10347
rect 15159 10329 15177 10347
rect 15195 10329 15213 10347
rect 15231 10329 17620 10347
rect 15040 10311 17620 10329
rect 15040 10293 15069 10311
rect 15087 10293 15105 10311
rect 15123 10293 15141 10311
rect 15159 10293 15177 10311
rect 15195 10293 15213 10311
rect 15231 10293 17620 10311
rect 15040 10280 17620 10293
rect 11960 8820 12040 10280
rect 17860 10140 17920 10680
rect 14660 10127 14880 10140
rect 14660 10109 14689 10127
rect 14707 10109 14725 10127
rect 14743 10109 14761 10127
rect 14779 10109 14797 10127
rect 14815 10109 14833 10127
rect 14851 10109 14880 10127
rect 14660 10091 14880 10109
rect 14660 10073 14689 10091
rect 14707 10073 14725 10091
rect 14743 10073 14761 10091
rect 14779 10073 14797 10091
rect 14815 10073 14833 10091
rect 14851 10073 14880 10091
rect 14660 10060 14880 10073
rect 17700 10127 17920 10140
rect 17700 10109 17729 10127
rect 17747 10109 17765 10127
rect 17783 10109 17801 10127
rect 17819 10109 17837 10127
rect 17855 10109 17873 10127
rect 17891 10109 17920 10127
rect 17700 10091 17920 10109
rect 20260 10100 20320 10680
rect 17700 10073 17729 10091
rect 17747 10073 17765 10091
rect 17783 10073 17801 10091
rect 17819 10073 17837 10091
rect 17855 10073 17873 10091
rect 17891 10073 17920 10091
rect 17700 10060 17920 10073
rect 14660 8820 14740 10060
rect 20060 10020 20320 10100
rect 17360 9827 17540 9840
rect 17360 9809 17387 9827
rect 17405 9809 17423 9827
rect 17441 9809 17459 9827
rect 17477 9809 17495 9827
rect 17513 9809 17540 9827
rect 17360 9791 17540 9809
rect 17360 9773 17387 9791
rect 17405 9773 17423 9791
rect 17441 9773 17459 9791
rect 17477 9773 17495 9791
rect 17513 9773 17540 9791
rect 17360 9760 17540 9773
rect 17360 8820 17440 9760
rect 20060 8820 20140 10020
rect 20380 9840 20440 10680
rect 20260 9827 20440 9840
rect 20260 9809 20287 9827
rect 20305 9809 20323 9827
rect 20341 9809 20359 9827
rect 20377 9809 20395 9827
rect 20413 9809 20440 9827
rect 20260 9791 20440 9809
rect 20260 9773 20287 9791
rect 20305 9773 20323 9791
rect 20341 9773 20359 9791
rect 20377 9773 20395 9791
rect 20413 9773 20440 9791
rect 20260 9760 20440 9773
rect 22720 9640 22780 10680
rect 22840 9880 22900 10680
rect 22840 9867 23040 9880
rect 22840 9849 22859 9867
rect 22877 9849 22895 9867
rect 22913 9849 22931 9867
rect 22949 9849 22967 9867
rect 22985 9849 23003 9867
rect 23021 9849 23040 9867
rect 22840 9831 23040 9849
rect 22840 9813 22859 9831
rect 22877 9813 22895 9831
rect 22913 9813 22931 9831
rect 22949 9813 22967 9831
rect 22985 9813 23003 9831
rect 23021 9813 23040 9831
rect 22840 9800 23040 9813
rect 20600 9560 22780 9640
rect 23140 9640 23200 10680
rect 23140 9627 23340 9640
rect 23140 9609 23159 9627
rect 23177 9609 23195 9627
rect 23213 9609 23231 9627
rect 23249 9609 23267 9627
rect 23285 9609 23303 9627
rect 23321 9609 23340 9627
rect 23140 9591 23340 9609
rect 23140 9573 23159 9591
rect 23177 9573 23195 9591
rect 23213 9573 23231 9591
rect 23249 9573 23267 9591
rect 23285 9573 23303 9591
rect 23321 9573 23340 9591
rect 23140 9560 23340 9573
rect 20600 8820 20680 9560
rect 23380 9220 23440 10680
rect 26420 9867 29180 9880
rect 26420 9849 26433 9867
rect 26451 9849 26469 9867
rect 26487 9849 26505 9867
rect 26523 9849 26541 9867
rect 26559 9849 26577 9867
rect 26595 9849 26613 9867
rect 26631 9849 26649 9867
rect 26667 9849 29180 9867
rect 26420 9831 29180 9849
rect 26420 9813 26433 9831
rect 26451 9813 26469 9831
rect 26487 9813 26505 9831
rect 26523 9813 26541 9831
rect 26559 9813 26577 9831
rect 26595 9813 26613 9831
rect 26631 9813 26649 9831
rect 26667 9813 29180 9831
rect 26420 9800 29180 9813
rect 25820 9627 26080 9640
rect 25820 9609 25833 9627
rect 25851 9609 25869 9627
rect 25887 9609 25905 9627
rect 25923 9609 25941 9627
rect 25959 9609 25977 9627
rect 25995 9609 26013 9627
rect 26031 9609 26049 9627
rect 26067 9609 26080 9627
rect 25820 9591 26080 9609
rect 25820 9573 25833 9591
rect 25851 9573 25869 9591
rect 25887 9573 25905 9591
rect 25923 9573 25941 9591
rect 25959 9573 25977 9591
rect 25995 9573 26013 9591
rect 26031 9573 26049 9591
rect 26067 9573 26080 9591
rect 25820 9560 26080 9573
rect 23300 9140 23440 9220
rect 23300 8820 23380 9140
rect 26000 8820 26080 9560
<< m3contact >>
rect 11981 28129 11999 28147
rect 12017 28129 12035 28147
rect 12053 28129 12071 28147
rect 12089 28129 12107 28147
rect 12125 28129 12143 28147
rect 12161 28129 12179 28147
rect 11981 28093 11999 28111
rect 12017 28093 12035 28111
rect 12053 28093 12071 28111
rect 12089 28093 12107 28111
rect 12125 28093 12143 28111
rect 12161 28093 12179 28111
rect 17379 28349 17397 28367
rect 17415 28349 17433 28367
rect 17451 28349 17469 28367
rect 17487 28349 17505 28367
rect 17523 28349 17541 28367
rect 17379 28313 17397 28331
rect 17415 28313 17433 28331
rect 17451 28313 17469 28331
rect 17487 28313 17505 28331
rect 17523 28313 17541 28331
rect 19899 28349 19917 28367
rect 19935 28349 19953 28367
rect 19971 28349 19989 28367
rect 20007 28349 20025 28367
rect 20043 28349 20061 28367
rect 19899 28313 19917 28331
rect 19935 28313 19953 28331
rect 19971 28313 19989 28331
rect 20007 28313 20025 28331
rect 20043 28313 20061 28331
rect 15983 28129 16001 28147
rect 16019 28129 16037 28147
rect 16055 28129 16073 28147
rect 16091 28129 16109 28147
rect 16127 28129 16145 28147
rect 16163 28129 16181 28147
rect 16199 28129 16217 28147
rect 15983 28093 16001 28111
rect 16019 28093 16037 28111
rect 16055 28093 16073 28111
rect 16091 28093 16109 28111
rect 16127 28093 16145 28111
rect 16163 28093 16181 28111
rect 16199 28093 16217 28111
rect 14675 27919 14693 27937
rect 14711 27919 14729 27937
rect 14747 27919 14765 27937
rect 14783 27919 14801 27937
rect 14819 27919 14837 27937
rect 14855 27919 14873 27937
rect 14891 27919 14909 27937
rect 14927 27919 14945 27937
rect 14675 27883 14693 27901
rect 14711 27883 14729 27901
rect 14747 27883 14765 27901
rect 14783 27883 14801 27901
rect 14819 27883 14837 27901
rect 14855 27883 14873 27901
rect 14891 27883 14909 27901
rect 14927 27883 14945 27901
rect 17303 27919 17321 27937
rect 17339 27919 17357 27937
rect 17375 27919 17393 27937
rect 17411 27919 17429 27937
rect 17447 27919 17465 27937
rect 17483 27919 17501 27937
rect 17519 27919 17537 27937
rect 17303 27883 17321 27901
rect 17339 27883 17357 27901
rect 17375 27883 17393 27901
rect 17411 27883 17429 27901
rect 17447 27883 17465 27901
rect 17483 27883 17501 27901
rect 17519 27883 17537 27901
rect 22005 28569 22023 28587
rect 22041 28569 22059 28587
rect 22077 28569 22095 28587
rect 22113 28569 22131 28587
rect 22149 28569 22167 28587
rect 22185 28569 22203 28587
rect 22221 28569 22239 28587
rect 22257 28569 22275 28587
rect 22005 28533 22023 28551
rect 22041 28533 22059 28551
rect 22077 28533 22095 28551
rect 22113 28533 22131 28551
rect 22149 28533 22167 28551
rect 22185 28533 22203 28551
rect 22221 28533 22239 28551
rect 22257 28533 22275 28551
rect 27993 28569 28011 28587
rect 28029 28569 28047 28587
rect 28065 28569 28083 28587
rect 28101 28569 28119 28587
rect 28137 28569 28155 28587
rect 28173 28569 28191 28587
rect 28209 28569 28227 28587
rect 27993 28533 28011 28551
rect 28029 28533 28047 28551
rect 28065 28533 28083 28551
rect 28101 28533 28119 28551
rect 28137 28533 28155 28551
rect 28173 28533 28191 28551
rect 28209 28533 28227 28551
rect 22923 28069 22941 28087
rect 22959 28069 22977 28087
rect 22995 28069 23013 28087
rect 23031 28069 23049 28087
rect 23067 28069 23085 28087
rect 23103 28069 23121 28087
rect 23139 28069 23157 28087
rect 22923 28033 22941 28051
rect 22959 28033 22977 28051
rect 22995 28033 23013 28051
rect 23031 28033 23049 28051
rect 23067 28033 23085 28051
rect 23103 28033 23121 28051
rect 23139 28033 23157 28051
rect 25283 28069 25301 28087
rect 25319 28069 25337 28087
rect 25355 28069 25373 28087
rect 25391 28069 25409 28087
rect 25427 28069 25445 28087
rect 25463 28069 25481 28087
rect 25499 28069 25517 28087
rect 25283 28033 25301 28051
rect 25319 28033 25337 28051
rect 25355 28033 25373 28051
rect 25391 28033 25409 28051
rect 25427 28033 25445 28051
rect 25463 28033 25481 28051
rect 25499 28033 25517 28051
rect 28273 26039 28291 26057
rect 28309 26039 28327 26057
rect 28273 26003 28291 26021
rect 28309 26003 28327 26021
rect 28273 25967 28291 25985
rect 28309 25967 28327 25985
rect 28273 25931 28291 25949
rect 28309 25931 28327 25949
rect 28273 25895 28291 25913
rect 28309 25895 28327 25913
rect 28273 25859 28291 25877
rect 28309 25859 28327 25877
rect 28273 25823 28291 25841
rect 28309 25823 28327 25841
rect 28553 23349 28571 23367
rect 28589 23349 28607 23367
rect 9873 23301 9891 23319
rect 9909 23301 9927 23319
rect 9873 23265 9891 23283
rect 9909 23265 9927 23283
rect 9873 23229 9891 23247
rect 9909 23229 9927 23247
rect 9873 23193 9891 23211
rect 9909 23193 9927 23211
rect 9873 23157 9891 23175
rect 9909 23157 9927 23175
rect 9873 23121 9891 23139
rect 9909 23121 9927 23139
rect 28553 23313 28571 23331
rect 28589 23313 28607 23331
rect 28553 23277 28571 23295
rect 28589 23277 28607 23295
rect 28553 23241 28571 23259
rect 28589 23241 28607 23259
rect 28553 23205 28571 23223
rect 28589 23205 28607 23223
rect 28553 23169 28571 23187
rect 28589 23169 28607 23187
rect 28553 23133 28571 23151
rect 28589 23133 28607 23151
rect 28563 20867 28581 20885
rect 28599 20867 28617 20885
rect 28563 20831 28581 20849
rect 28599 20831 28617 20849
rect 28563 20795 28581 20813
rect 28599 20795 28617 20813
rect 9893 20733 9911 20751
rect 9929 20733 9947 20751
rect 9893 20697 9911 20715
rect 9929 20697 9947 20715
rect 9893 20661 9911 20679
rect 9929 20661 9947 20679
rect 9893 20625 9911 20643
rect 9929 20625 9947 20643
rect 9893 20589 9911 20607
rect 9929 20589 9947 20607
rect 28563 20759 28581 20777
rect 28599 20759 28617 20777
rect 28563 20723 28581 20741
rect 28599 20723 28617 20741
rect 28563 20687 28581 20705
rect 28599 20687 28617 20705
rect 28563 20651 28581 20669
rect 28599 20651 28617 20669
rect 28563 20615 28581 20633
rect 28599 20615 28617 20633
rect 9413 18033 9431 18051
rect 9449 18033 9467 18051
rect 9413 17997 9431 18015
rect 9449 17997 9467 18015
rect 9413 17961 9431 17979
rect 9449 17961 9467 17979
rect 9413 17925 9431 17943
rect 9449 17925 9467 17943
rect 9413 17889 9431 17907
rect 9449 17889 9467 17907
rect 9633 17633 9651 17651
rect 9669 17633 9687 17651
rect 9633 17597 9651 17615
rect 9669 17597 9687 17615
rect 9633 17561 9651 17579
rect 9669 17561 9687 17579
rect 9633 17525 9651 17543
rect 9669 17525 9687 17543
rect 9633 17489 9651 17507
rect 9669 17489 9687 17507
rect 28393 15429 28411 15447
rect 28429 15429 28447 15447
rect 28393 15393 28411 15411
rect 28429 15393 28447 15411
rect 28393 15357 28411 15375
rect 28429 15357 28447 15375
rect 28393 15321 28411 15339
rect 28429 15321 28447 15339
rect 28393 15285 28411 15303
rect 28429 15285 28447 15303
rect 28393 15249 28411 15267
rect 28429 15249 28447 15267
rect 28393 15213 28411 15231
rect 28429 15213 28447 15231
rect 9893 14419 9911 14437
rect 9929 14419 9947 14437
rect 9893 14383 9911 14401
rect 9929 14383 9947 14401
rect 9893 14347 9911 14365
rect 9929 14347 9947 14365
rect 9893 14311 9911 14329
rect 9929 14311 9947 14329
rect 9893 14275 9911 14293
rect 9929 14275 9947 14293
rect 9893 14239 9911 14257
rect 9929 14239 9947 14257
rect 9893 14203 9911 14221
rect 9929 14203 9947 14221
rect 28173 12729 28191 12747
rect 28209 12729 28227 12747
rect 28173 12693 28191 12711
rect 28209 12693 28227 12711
rect 28173 12657 28191 12675
rect 28209 12657 28227 12675
rect 28173 12621 28191 12639
rect 28209 12621 28227 12639
rect 28173 12585 28191 12603
rect 28209 12585 28227 12603
rect 28173 12549 28191 12567
rect 28209 12549 28227 12567
rect 28173 12513 28191 12531
rect 28209 12513 28227 12531
rect 11989 10329 12007 10347
rect 12025 10329 12043 10347
rect 12061 10329 12079 10347
rect 12097 10329 12115 10347
rect 12133 10329 12151 10347
rect 11989 10293 12007 10311
rect 12025 10293 12043 10311
rect 12061 10293 12079 10311
rect 12097 10293 12115 10311
rect 12133 10293 12151 10311
rect 15069 10329 15087 10347
rect 15105 10329 15123 10347
rect 15141 10329 15159 10347
rect 15177 10329 15195 10347
rect 15213 10329 15231 10347
rect 15069 10293 15087 10311
rect 15105 10293 15123 10311
rect 15141 10293 15159 10311
rect 15177 10293 15195 10311
rect 15213 10293 15231 10311
rect 14689 10109 14707 10127
rect 14725 10109 14743 10127
rect 14761 10109 14779 10127
rect 14797 10109 14815 10127
rect 14833 10109 14851 10127
rect 14689 10073 14707 10091
rect 14725 10073 14743 10091
rect 14761 10073 14779 10091
rect 14797 10073 14815 10091
rect 14833 10073 14851 10091
rect 17729 10109 17747 10127
rect 17765 10109 17783 10127
rect 17801 10109 17819 10127
rect 17837 10109 17855 10127
rect 17873 10109 17891 10127
rect 17729 10073 17747 10091
rect 17765 10073 17783 10091
rect 17801 10073 17819 10091
rect 17837 10073 17855 10091
rect 17873 10073 17891 10091
rect 17387 9809 17405 9827
rect 17423 9809 17441 9827
rect 17459 9809 17477 9827
rect 17495 9809 17513 9827
rect 17387 9773 17405 9791
rect 17423 9773 17441 9791
rect 17459 9773 17477 9791
rect 17495 9773 17513 9791
rect 20287 9809 20305 9827
rect 20323 9809 20341 9827
rect 20359 9809 20377 9827
rect 20395 9809 20413 9827
rect 20287 9773 20305 9791
rect 20323 9773 20341 9791
rect 20359 9773 20377 9791
rect 20395 9773 20413 9791
rect 22859 9849 22877 9867
rect 22895 9849 22913 9867
rect 22931 9849 22949 9867
rect 22967 9849 22985 9867
rect 23003 9849 23021 9867
rect 22859 9813 22877 9831
rect 22895 9813 22913 9831
rect 22931 9813 22949 9831
rect 22967 9813 22985 9831
rect 23003 9813 23021 9831
rect 23159 9609 23177 9627
rect 23195 9609 23213 9627
rect 23231 9609 23249 9627
rect 23267 9609 23285 9627
rect 23303 9609 23321 9627
rect 23159 9573 23177 9591
rect 23195 9573 23213 9591
rect 23231 9573 23249 9591
rect 23267 9573 23285 9591
rect 23303 9573 23321 9591
rect 26433 9849 26451 9867
rect 26469 9849 26487 9867
rect 26505 9849 26523 9867
rect 26541 9849 26559 9867
rect 26577 9849 26595 9867
rect 26613 9849 26631 9867
rect 26649 9849 26667 9867
rect 26433 9813 26451 9831
rect 26469 9813 26487 9831
rect 26505 9813 26523 9831
rect 26541 9813 26559 9831
rect 26577 9813 26595 9831
rect 26613 9813 26631 9831
rect 26649 9813 26667 9831
rect 25833 9609 25851 9627
rect 25869 9609 25887 9627
rect 25905 9609 25923 9627
rect 25941 9609 25959 9627
rect 25977 9609 25995 9627
rect 26013 9609 26031 9627
rect 26049 9609 26067 9627
rect 25833 9573 25851 9591
rect 25869 9573 25887 9591
rect 25905 9573 25923 9591
rect 25941 9573 25959 9591
rect 25977 9573 25995 9591
rect 26013 9573 26031 9591
rect 26049 9573 26067 9591
<< metal3 >>
rect 21980 28587 28240 28600
rect 21980 28569 22005 28587
rect 22023 28569 22041 28587
rect 22059 28569 22077 28587
rect 22095 28569 22113 28587
rect 22131 28569 22149 28587
rect 22167 28569 22185 28587
rect 22203 28569 22221 28587
rect 22239 28569 22257 28587
rect 22275 28569 27993 28587
rect 28011 28569 28029 28587
rect 28047 28569 28065 28587
rect 28083 28569 28101 28587
rect 28119 28569 28137 28587
rect 28155 28569 28173 28587
rect 28191 28569 28209 28587
rect 28227 28569 28240 28587
rect 21980 28551 28240 28569
rect 21980 28533 22005 28551
rect 22023 28533 22041 28551
rect 22059 28533 22077 28551
rect 22095 28533 22113 28551
rect 22131 28533 22149 28551
rect 22167 28533 22185 28551
rect 22203 28533 22221 28551
rect 22239 28533 22257 28551
rect 22275 28533 27993 28551
rect 28011 28533 28029 28551
rect 28047 28533 28065 28551
rect 28083 28533 28101 28551
rect 28119 28533 28137 28551
rect 28155 28533 28173 28551
rect 28191 28533 28209 28551
rect 28227 28533 28240 28551
rect 21980 28520 28240 28533
rect 17360 28367 20080 28380
rect 17360 28349 17379 28367
rect 17397 28349 17415 28367
rect 17433 28349 17451 28367
rect 17469 28349 17487 28367
rect 17505 28349 17523 28367
rect 17541 28349 19899 28367
rect 19917 28349 19935 28367
rect 19953 28349 19971 28367
rect 19989 28349 20007 28367
rect 20025 28349 20043 28367
rect 20061 28349 20080 28367
rect 17360 28331 20080 28349
rect 17360 28313 17379 28331
rect 17397 28313 17415 28331
rect 17433 28313 17451 28331
rect 17469 28313 17487 28331
rect 17505 28313 17523 28331
rect 17541 28313 19899 28331
rect 19917 28313 19935 28331
rect 19953 28313 19971 28331
rect 19989 28313 20007 28331
rect 20025 28313 20043 28331
rect 20061 28313 20080 28331
rect 17360 28300 20080 28313
rect 11960 28147 16240 28160
rect 11960 28129 11981 28147
rect 11999 28129 12017 28147
rect 12035 28129 12053 28147
rect 12071 28129 12089 28147
rect 12107 28129 12125 28147
rect 12143 28129 12161 28147
rect 12179 28129 15983 28147
rect 16001 28129 16019 28147
rect 16037 28129 16055 28147
rect 16073 28129 16091 28147
rect 16109 28129 16127 28147
rect 16145 28129 16163 28147
rect 16181 28129 16199 28147
rect 16217 28129 16240 28147
rect 11960 28111 16240 28129
rect 11960 28093 11981 28111
rect 11999 28093 12017 28111
rect 12035 28093 12053 28111
rect 12071 28093 12089 28111
rect 12107 28093 12125 28111
rect 12143 28093 12161 28111
rect 12179 28093 15983 28111
rect 16001 28093 16019 28111
rect 16037 28093 16055 28111
rect 16073 28093 16091 28111
rect 16109 28093 16127 28111
rect 16145 28093 16163 28111
rect 16181 28093 16199 28111
rect 16217 28093 16240 28111
rect 11960 28080 16240 28093
rect 22900 28087 25540 28100
rect 22900 28069 22923 28087
rect 22941 28069 22959 28087
rect 22977 28069 22995 28087
rect 23013 28069 23031 28087
rect 23049 28069 23067 28087
rect 23085 28069 23103 28087
rect 23121 28069 23139 28087
rect 23157 28069 25283 28087
rect 25301 28069 25319 28087
rect 25337 28069 25355 28087
rect 25373 28069 25391 28087
rect 25409 28069 25427 28087
rect 25445 28069 25463 28087
rect 25481 28069 25499 28087
rect 25517 28069 25540 28087
rect 22900 28051 25540 28069
rect 22900 28033 22923 28051
rect 22941 28033 22959 28051
rect 22977 28033 22995 28051
rect 23013 28033 23031 28051
rect 23049 28033 23067 28051
rect 23085 28033 23103 28051
rect 23121 28033 23139 28051
rect 23157 28033 25283 28051
rect 25301 28033 25319 28051
rect 25337 28033 25355 28051
rect 25373 28033 25391 28051
rect 25409 28033 25427 28051
rect 25445 28033 25463 28051
rect 25481 28033 25499 28051
rect 25517 28033 25540 28051
rect 22900 28020 25540 28033
rect 14660 27937 17560 27960
rect 14660 27919 14675 27937
rect 14693 27919 14711 27937
rect 14729 27919 14747 27937
rect 14765 27919 14783 27937
rect 14801 27919 14819 27937
rect 14837 27919 14855 27937
rect 14873 27919 14891 27937
rect 14909 27919 14927 27937
rect 14945 27919 17303 27937
rect 17321 27919 17339 27937
rect 17357 27919 17375 27937
rect 17393 27919 17411 27937
rect 17429 27919 17447 27937
rect 17465 27919 17483 27937
rect 17501 27919 17519 27937
rect 17537 27919 17560 27937
rect 14660 27901 17560 27919
rect 14660 27883 14675 27901
rect 14693 27883 14711 27901
rect 14729 27883 14747 27901
rect 14765 27883 14783 27901
rect 14801 27883 14819 27901
rect 14837 27883 14855 27901
rect 14873 27883 14891 27901
rect 14909 27883 14927 27901
rect 14945 27883 17303 27901
rect 17321 27883 17339 27901
rect 17357 27883 17375 27901
rect 17393 27883 17411 27901
rect 17429 27883 17447 27901
rect 17465 27883 17483 27901
rect 17501 27883 17519 27901
rect 17537 27883 17560 27901
rect 14660 27860 17560 27883
rect 28260 26057 28340 26080
rect 28260 26039 28273 26057
rect 28291 26039 28309 26057
rect 28327 26039 28340 26057
rect 28260 26021 28340 26039
rect 28260 26003 28273 26021
rect 28291 26003 28309 26021
rect 28327 26003 28340 26021
rect 28260 25985 28340 26003
rect 28260 25967 28273 25985
rect 28291 25967 28309 25985
rect 28327 25967 28340 25985
rect 28260 25949 28340 25967
rect 28260 25931 28273 25949
rect 28291 25931 28309 25949
rect 28327 25931 28340 25949
rect 28260 25913 28340 25931
rect 28260 25895 28273 25913
rect 28291 25895 28309 25913
rect 28327 25895 28340 25913
rect 28260 25877 28340 25895
rect 28260 25859 28273 25877
rect 28291 25859 28309 25877
rect 28327 25859 28340 25877
rect 28260 25841 28340 25859
rect 28260 25823 28273 25841
rect 28291 25823 28309 25841
rect 28327 25823 28340 25841
rect 9860 23319 9940 23340
rect 9860 23301 9873 23319
rect 9891 23301 9909 23319
rect 9927 23301 9940 23319
rect 9860 23283 9940 23301
rect 9860 23265 9873 23283
rect 9891 23265 9909 23283
rect 9927 23265 9940 23283
rect 9860 23247 9940 23265
rect 9860 23229 9873 23247
rect 9891 23229 9909 23247
rect 9927 23229 9940 23247
rect 9860 23211 9940 23229
rect 9860 23193 9873 23211
rect 9891 23193 9909 23211
rect 9927 23193 9940 23211
rect 9860 23175 9940 23193
rect 9860 23157 9873 23175
rect 9891 23157 9909 23175
rect 9927 23157 9940 23175
rect 9860 23139 9940 23157
rect 9860 23121 9873 23139
rect 9891 23121 9909 23139
rect 9927 23121 9940 23139
rect 9860 21440 9940 23121
rect 28260 23020 28340 25823
rect 27780 22940 28340 23020
rect 28540 23367 28620 23380
rect 28540 23349 28553 23367
rect 28571 23349 28589 23367
rect 28607 23349 28620 23367
rect 28540 23331 28620 23349
rect 28540 23313 28553 23331
rect 28571 23313 28589 23331
rect 28607 23313 28620 23331
rect 28540 23295 28620 23313
rect 28540 23277 28553 23295
rect 28571 23277 28589 23295
rect 28607 23277 28620 23295
rect 28540 23259 28620 23277
rect 28540 23241 28553 23259
rect 28571 23241 28589 23259
rect 28607 23241 28620 23259
rect 28540 23223 28620 23241
rect 28540 23205 28553 23223
rect 28571 23205 28589 23223
rect 28607 23205 28620 23223
rect 28540 23187 28620 23205
rect 28540 23169 28553 23187
rect 28571 23169 28589 23187
rect 28607 23169 28620 23187
rect 28540 23151 28620 23169
rect 28540 23133 28553 23151
rect 28571 23133 28589 23151
rect 28607 23133 28620 23151
rect 28540 22880 28620 23133
rect 27780 22800 28620 22880
rect 27780 22040 28640 22120
rect 9860 21380 10340 21440
rect 9880 21260 10340 21320
rect 9880 20751 9960 21260
rect 9880 20733 9893 20751
rect 9911 20733 9929 20751
rect 9947 20733 9960 20751
rect 9880 20715 9960 20733
rect 9880 20697 9893 20715
rect 9911 20697 9929 20715
rect 9947 20697 9960 20715
rect 9880 20679 9960 20697
rect 9880 20661 9893 20679
rect 9911 20661 9929 20679
rect 9947 20661 9960 20679
rect 9880 20643 9960 20661
rect 9880 20625 9893 20643
rect 9911 20625 9929 20643
rect 9947 20625 9960 20643
rect 9880 20607 9960 20625
rect 9880 20589 9893 20607
rect 9911 20589 9929 20607
rect 9947 20589 9960 20607
rect 28540 20885 28640 22040
rect 28540 20867 28563 20885
rect 28581 20867 28599 20885
rect 28617 20867 28640 20885
rect 28540 20849 28640 20867
rect 28540 20831 28563 20849
rect 28581 20831 28599 20849
rect 28617 20831 28640 20849
rect 28540 20813 28640 20831
rect 28540 20795 28563 20813
rect 28581 20795 28599 20813
rect 28617 20795 28640 20813
rect 28540 20777 28640 20795
rect 28540 20759 28563 20777
rect 28581 20759 28599 20777
rect 28617 20759 28640 20777
rect 28540 20741 28640 20759
rect 28540 20723 28563 20741
rect 28581 20723 28599 20741
rect 28617 20723 28640 20741
rect 28540 20705 28640 20723
rect 28540 20687 28563 20705
rect 28581 20687 28599 20705
rect 28617 20687 28640 20705
rect 28540 20669 28640 20687
rect 28540 20651 28563 20669
rect 28581 20651 28599 20669
rect 28617 20651 28640 20669
rect 28540 20633 28640 20651
rect 28540 20615 28563 20633
rect 28581 20615 28599 20633
rect 28617 20615 28640 20633
rect 28540 20600 28640 20615
rect 9880 20560 9960 20589
rect 9400 19820 10340 19880
rect 9400 18051 9480 19820
rect 9400 18033 9413 18051
rect 9431 18033 9449 18051
rect 9467 18033 9480 18051
rect 9400 18015 9480 18033
rect 9400 17997 9413 18015
rect 9431 17997 9449 18015
rect 9467 17997 9480 18015
rect 9400 17979 9480 17997
rect 9400 17961 9413 17979
rect 9431 17961 9449 17979
rect 9467 17961 9480 17979
rect 9400 17943 9480 17961
rect 9400 17925 9413 17943
rect 9431 17925 9449 17943
rect 9467 17925 9480 17943
rect 9400 17907 9480 17925
rect 9400 17889 9413 17907
rect 9431 17889 9449 17907
rect 9467 17889 9480 17907
rect 9400 17860 9480 17889
rect 9620 19700 10340 19760
rect 27760 19700 28460 19780
rect 9620 17651 9700 19700
rect 27760 18920 28240 19000
rect 9620 17633 9633 17651
rect 9651 17633 9669 17651
rect 9687 17633 9700 17651
rect 9620 17615 9700 17633
rect 9620 17597 9633 17615
rect 9651 17597 9669 17615
rect 9687 17597 9700 17615
rect 9620 17579 9700 17597
rect 9620 17561 9633 17579
rect 9651 17561 9669 17579
rect 9687 17561 9700 17579
rect 9620 17543 9700 17561
rect 9620 17525 9633 17543
rect 9651 17525 9669 17543
rect 9687 17525 9700 17543
rect 9620 17507 9700 17525
rect 9620 17489 9633 17507
rect 9651 17489 9669 17507
rect 9687 17489 9700 17507
rect 9620 17460 9700 17489
rect 9880 16580 10340 16640
rect 9880 14437 9960 16580
rect 9880 14419 9893 14437
rect 9911 14419 9929 14437
rect 9947 14419 9960 14437
rect 9880 14401 9960 14419
rect 9880 14383 9893 14401
rect 9911 14383 9929 14401
rect 9947 14383 9960 14401
rect 9880 14365 9960 14383
rect 9880 14347 9893 14365
rect 9911 14347 9929 14365
rect 9947 14347 9960 14365
rect 9880 14329 9960 14347
rect 9880 14311 9893 14329
rect 9911 14311 9929 14329
rect 9947 14311 9960 14329
rect 9880 14293 9960 14311
rect 9880 14275 9893 14293
rect 9911 14275 9929 14293
rect 9947 14275 9960 14293
rect 9880 14257 9960 14275
rect 9880 14239 9893 14257
rect 9911 14239 9929 14257
rect 9947 14239 9960 14257
rect 9880 14221 9960 14239
rect 9880 14203 9893 14221
rect 9911 14203 9929 14221
rect 9947 14203 9960 14221
rect 9880 14180 9960 14203
rect 28160 12747 28240 18920
rect 28380 15447 28460 19700
rect 28380 15429 28393 15447
rect 28411 15429 28429 15447
rect 28447 15429 28460 15447
rect 28380 15411 28460 15429
rect 28380 15393 28393 15411
rect 28411 15393 28429 15411
rect 28447 15393 28460 15411
rect 28380 15375 28460 15393
rect 28380 15357 28393 15375
rect 28411 15357 28429 15375
rect 28447 15357 28460 15375
rect 28380 15339 28460 15357
rect 28380 15321 28393 15339
rect 28411 15321 28429 15339
rect 28447 15321 28460 15339
rect 28380 15303 28460 15321
rect 28380 15285 28393 15303
rect 28411 15285 28429 15303
rect 28447 15285 28460 15303
rect 28380 15267 28460 15285
rect 28380 15249 28393 15267
rect 28411 15249 28429 15267
rect 28447 15249 28460 15267
rect 28380 15231 28460 15249
rect 28380 15213 28393 15231
rect 28411 15213 28429 15231
rect 28447 15213 28460 15231
rect 28380 15200 28460 15213
rect 28160 12729 28173 12747
rect 28191 12729 28209 12747
rect 28227 12729 28240 12747
rect 28160 12711 28240 12729
rect 28160 12693 28173 12711
rect 28191 12693 28209 12711
rect 28227 12693 28240 12711
rect 28160 12675 28240 12693
rect 28160 12657 28173 12675
rect 28191 12657 28209 12675
rect 28227 12657 28240 12675
rect 28160 12639 28240 12657
rect 28160 12621 28173 12639
rect 28191 12621 28209 12639
rect 28227 12621 28240 12639
rect 28160 12603 28240 12621
rect 28160 12585 28173 12603
rect 28191 12585 28209 12603
rect 28227 12585 28240 12603
rect 28160 12567 28240 12585
rect 28160 12549 28173 12567
rect 28191 12549 28209 12567
rect 28227 12549 28240 12567
rect 28160 12531 28240 12549
rect 28160 12513 28173 12531
rect 28191 12513 28209 12531
rect 28227 12513 28240 12531
rect 28160 12500 28240 12513
rect 11960 10347 15260 10360
rect 11960 10329 11989 10347
rect 12007 10329 12025 10347
rect 12043 10329 12061 10347
rect 12079 10329 12097 10347
rect 12115 10329 12133 10347
rect 12151 10329 15069 10347
rect 15087 10329 15105 10347
rect 15123 10329 15141 10347
rect 15159 10329 15177 10347
rect 15195 10329 15213 10347
rect 15231 10329 15260 10347
rect 11960 10311 15260 10329
rect 11960 10293 11989 10311
rect 12007 10293 12025 10311
rect 12043 10293 12061 10311
rect 12079 10293 12097 10311
rect 12115 10293 12133 10311
rect 12151 10293 15069 10311
rect 15087 10293 15105 10311
rect 15123 10293 15141 10311
rect 15159 10293 15177 10311
rect 15195 10293 15213 10311
rect 15231 10293 15260 10311
rect 11960 10280 15260 10293
rect 14660 10127 17920 10140
rect 14660 10109 14689 10127
rect 14707 10109 14725 10127
rect 14743 10109 14761 10127
rect 14779 10109 14797 10127
rect 14815 10109 14833 10127
rect 14851 10109 17729 10127
rect 17747 10109 17765 10127
rect 17783 10109 17801 10127
rect 17819 10109 17837 10127
rect 17855 10109 17873 10127
rect 17891 10109 17920 10127
rect 14660 10091 17920 10109
rect 14660 10073 14689 10091
rect 14707 10073 14725 10091
rect 14743 10073 14761 10091
rect 14779 10073 14797 10091
rect 14815 10073 14833 10091
rect 14851 10073 17729 10091
rect 17747 10073 17765 10091
rect 17783 10073 17801 10091
rect 17819 10073 17837 10091
rect 17855 10073 17873 10091
rect 17891 10073 17920 10091
rect 14660 10060 17920 10073
rect 22840 9867 26680 9880
rect 22840 9849 22859 9867
rect 22877 9849 22895 9867
rect 22913 9849 22931 9867
rect 22949 9849 22967 9867
rect 22985 9849 23003 9867
rect 23021 9849 26433 9867
rect 26451 9849 26469 9867
rect 26487 9849 26505 9867
rect 26523 9849 26541 9867
rect 26559 9849 26577 9867
rect 26595 9849 26613 9867
rect 26631 9849 26649 9867
rect 26667 9849 26680 9867
rect 17360 9827 20440 9840
rect 17360 9809 17387 9827
rect 17405 9809 17423 9827
rect 17441 9809 17459 9827
rect 17477 9809 17495 9827
rect 17513 9809 20287 9827
rect 20305 9809 20323 9827
rect 20341 9809 20359 9827
rect 20377 9809 20395 9827
rect 20413 9809 20440 9827
rect 17360 9791 20440 9809
rect 22840 9831 26680 9849
rect 22840 9813 22859 9831
rect 22877 9813 22895 9831
rect 22913 9813 22931 9831
rect 22949 9813 22967 9831
rect 22985 9813 23003 9831
rect 23021 9813 26433 9831
rect 26451 9813 26469 9831
rect 26487 9813 26505 9831
rect 26523 9813 26541 9831
rect 26559 9813 26577 9831
rect 26595 9813 26613 9831
rect 26631 9813 26649 9831
rect 26667 9813 26680 9831
rect 22840 9800 26680 9813
rect 17360 9773 17387 9791
rect 17405 9773 17423 9791
rect 17441 9773 17459 9791
rect 17477 9773 17495 9791
rect 17513 9773 20287 9791
rect 20305 9773 20323 9791
rect 20341 9773 20359 9791
rect 20377 9773 20395 9791
rect 20413 9773 20440 9791
rect 17360 9760 20440 9773
rect 23140 9627 26080 9640
rect 23140 9609 23159 9627
rect 23177 9609 23195 9627
rect 23213 9609 23231 9627
rect 23249 9609 23267 9627
rect 23285 9609 23303 9627
rect 23321 9609 25833 9627
rect 25851 9609 25869 9627
rect 25887 9609 25905 9627
rect 25923 9609 25941 9627
rect 25959 9609 25977 9627
rect 25995 9609 26013 9627
rect 26031 9609 26049 9627
rect 26067 9609 26080 9627
rect 23140 9591 26080 9609
rect 23140 9573 23159 9591
rect 23177 9573 23195 9591
rect 23213 9573 23231 9591
rect 23249 9573 23267 9591
rect 23285 9573 23303 9591
rect 23321 9573 25833 9591
rect 25851 9573 25869 9591
rect 25887 9573 25905 9591
rect 25923 9573 25941 9591
rect 25959 9573 25977 9591
rect 25995 9573 26013 9591
rect 26031 9573 26049 9591
rect 26067 9573 26080 9591
rect 23140 9560 26080 9573
<< end >>
