magic
tech scmos
timestamp 1537935238
<< checkpaint >>
rect -21 -21 21 21
<< genericcontact >>
rect -1 -1 1 1
<< end >>
