magic
tech scmos
magscale 1 2
timestamp 1728304421
<< nwell >>
rect -12 134 212 252
<< ntransistor >>
rect 21 14 25 54
rect 41 14 45 54
rect 61 14 65 54
rect 81 14 85 54
rect 101 14 105 54
rect 121 14 125 54
rect 141 14 145 54
rect 161 14 165 54
<< ptransistor >>
rect 21 146 25 226
rect 41 146 45 226
rect 61 146 65 226
rect 81 146 85 226
rect 101 146 105 226
rect 121 146 125 226
rect 141 146 145 226
rect 161 146 165 226
<< ndiffusion >>
rect 19 14 21 54
rect 25 14 27 54
rect 39 14 41 54
rect 45 14 47 54
rect 59 14 61 54
rect 65 14 67 54
rect 79 14 81 54
rect 85 14 87 54
rect 99 14 101 54
rect 105 14 107 54
rect 119 14 121 54
rect 125 14 127 54
rect 139 14 141 54
rect 145 14 147 54
rect 159 14 161 54
rect 165 14 167 54
<< pdiffusion >>
rect 19 146 21 226
rect 25 146 27 226
rect 39 146 41 226
rect 45 146 47 226
rect 59 146 61 226
rect 65 146 67 226
rect 79 146 81 226
rect 85 146 87 226
rect 99 146 101 226
rect 105 146 107 226
rect 119 146 121 226
rect 125 146 127 226
rect 139 146 141 226
rect 145 146 147 226
rect 159 146 161 226
rect 165 146 167 226
<< ndcontact >>
rect 7 14 19 54
rect 27 14 39 54
rect 47 14 59 54
rect 67 14 79 54
rect 87 14 99 54
rect 107 14 119 54
rect 127 14 139 54
rect 147 14 159 54
rect 167 14 179 54
<< pdcontact >>
rect 7 146 19 226
rect 27 146 39 226
rect 47 146 59 226
rect 67 146 79 226
rect 87 146 99 226
rect 107 146 119 226
rect 127 146 139 226
rect 147 146 159 226
rect 167 146 179 226
<< psubstratepcontact >>
rect -6 -6 206 6
<< nsubstratencontact >>
rect -6 234 206 246
<< polysilicon >>
rect 21 226 25 230
rect 41 226 45 230
rect 61 226 65 230
rect 81 226 85 230
rect 101 226 105 230
rect 121 226 125 230
rect 141 226 145 230
rect 161 226 165 230
rect 21 89 25 146
rect 41 89 45 146
rect 21 77 24 89
rect 36 77 45 89
rect 61 86 65 146
rect 81 86 85 146
rect 101 86 105 146
rect 121 86 125 146
rect 141 86 145 146
rect 161 86 165 146
rect 21 54 25 77
rect 41 54 45 77
rect 72 74 85 86
rect 112 74 125 86
rect 152 74 165 86
rect 61 54 65 74
rect 81 54 85 74
rect 101 54 105 74
rect 121 54 125 74
rect 141 54 145 74
rect 161 54 165 74
rect 21 10 25 14
rect 41 10 45 14
rect 61 10 65 14
rect 81 10 85 14
rect 101 10 105 14
rect 121 10 125 14
rect 141 10 145 14
rect 161 10 165 14
<< polycontact >>
rect 24 77 36 89
rect 60 74 72 86
rect 100 74 112 86
rect 140 74 152 86
<< metal1 >>
rect -6 246 206 248
rect -6 232 206 234
rect 7 226 19 232
rect 47 226 59 232
rect 87 226 99 232
rect 127 226 139 232
rect 167 226 179 232
rect 27 140 39 146
rect 67 140 79 146
rect 107 140 119 146
rect 147 140 159 146
rect 27 132 53 140
rect 67 132 92 140
rect 107 132 132 140
rect 147 132 165 140
rect 45 86 53 132
rect 84 86 92 132
rect 124 86 132 132
rect 158 103 165 132
rect 158 89 163 103
rect 45 74 60 86
rect 84 74 100 86
rect 124 74 140 86
rect 45 68 53 74
rect 84 68 92 74
rect 124 68 132 74
rect 158 68 165 89
rect 26 60 53 68
rect 67 60 92 68
rect 106 60 132 68
rect 146 61 165 68
rect 146 60 164 61
rect 26 54 38 60
rect 67 54 79 60
rect 106 54 118 60
rect 146 54 158 60
rect 7 8 19 14
rect 47 8 59 14
rect 87 8 99 14
rect 127 8 139 14
rect 167 8 179 14
rect -6 6 206 8
rect -6 -8 206 -6
<< m2contact >>
rect 23 89 37 103
rect 163 89 177 103
<< metal2 >>
rect 23 103 37 117
rect 163 103 177 117
<< m1p >>
rect -6 232 206 248
rect -6 -8 206 8
<< m2p >>
rect 23 103 37 117
rect 163 103 177 117
<< labels >>
rlabel metal1 -6 -8 206 8 0 gnd
port 3 nsew ground bidirectional abutment
rlabel metal1 -6 232 206 248 0 vdd
port 2 nsew power bidirectional abutment
rlabel metal2 23 103 37 117 0 A
port 0 nsew signal input
rlabel metal2 163 103 177 117 0 Y
port 1 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 200 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
