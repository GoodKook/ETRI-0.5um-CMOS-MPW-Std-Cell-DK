VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fir_pe
  CLASS BLOCK ;
  FOREIGN fir_pe ;
  ORIGIN 6.000 6.000 ;
  SIZE 924.000 BY 912.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 1.500 897.300 920.550 899.700 ;
        RECT 22.800 887.400 24.600 897.300 ;
        RECT 36.000 890.400 37.800 897.300 ;
        RECT 43.800 893.400 45.600 897.300 ;
        RECT 70.800 887.400 72.600 897.300 ;
        RECT 94.800 887.400 96.600 897.300 ;
        RECT 115.800 892.200 117.600 897.300 ;
        RECT 139.800 892.200 141.600 897.300 ;
        RECT 155.400 893.400 157.200 897.300 ;
        RECT 173.400 893.400 175.200 897.300 ;
        RECT 192.000 890.400 193.800 897.300 ;
        RECT 199.800 893.400 201.600 897.300 ;
        RECT 223.500 890.400 225.300 897.300 ;
        RECT 239.400 892.200 241.200 897.300 ;
        RECT 260.700 890.400 262.500 897.300 ;
        RECT 286.500 890.400 288.300 897.300 ;
        RECT 305.700 890.400 307.500 897.300 ;
        RECT 331.500 890.400 333.300 897.300 ;
        RECT 348.900 890.400 350.700 897.300 ;
        RECT 376.500 890.400 378.300 897.300 ;
        RECT 389.700 890.400 391.500 897.300 ;
        RECT 412.800 893.400 414.600 897.300 ;
        RECT 418.800 893.400 420.600 897.300 ;
        RECT 431.700 890.400 433.500 897.300 ;
        RECT 455.700 890.400 457.500 897.300 ;
        RECT 480.300 890.400 482.100 897.300 ;
        RECT 500.400 893.400 502.200 897.300 ;
        RECT 508.200 890.400 510.000 897.300 ;
        RECT 532.800 887.400 534.600 897.300 ;
        RECT 545.700 890.400 547.500 897.300 ;
        RECT 577.800 887.400 579.600 897.300 ;
        RECT 598.500 890.400 600.300 897.300 ;
        RECT 614.700 890.400 616.500 897.300 ;
        RECT 637.500 890.400 639.300 897.300 ;
        RECT 646.500 890.400 648.300 897.300 ;
        RECT 664.500 890.400 666.300 897.300 ;
        RECT 685.800 893.400 687.600 897.300 ;
        RECT 701.700 890.400 703.500 897.300 ;
        RECT 726.300 890.400 728.100 897.300 ;
        RECT 743.700 890.400 745.500 897.300 ;
        RECT 752.700 890.400 754.500 897.300 ;
        RECT 774.900 890.400 776.700 897.300 ;
        RECT 799.500 890.400 801.300 897.300 ;
        RECT 808.500 890.400 810.300 897.300 ;
        RECT 821.700 890.400 823.500 897.300 ;
        RECT 845.400 892.200 847.200 897.300 ;
        RECT 866.400 893.400 868.200 897.300 ;
        RECT 884.400 896.400 885.600 897.300 ;
        RECT 884.400 893.400 886.200 896.400 ;
        RECT 890.400 893.400 892.200 897.300 ;
        RECT 22.800 821.700 24.600 831.600 ;
        RECT 36.000 821.700 37.800 828.600 ;
        RECT 43.800 821.700 45.600 825.600 ;
        RECT 70.800 821.700 72.600 831.600 ;
        RECT 84.000 821.700 85.800 828.600 ;
        RECT 91.800 821.700 93.600 825.600 ;
        RECT 110.400 821.700 112.200 825.600 ;
        RECT 118.200 821.700 120.000 828.600 ;
        RECT 136.800 821.700 138.600 825.600 ;
        RECT 152.400 821.700 154.200 826.800 ;
        RECT 181.800 821.700 183.600 826.800 ;
        RECT 197.400 821.700 199.200 825.600 ;
        RECT 203.400 821.700 205.200 825.600 ;
        RECT 218.400 821.700 220.200 825.600 ;
        RECT 224.400 821.700 226.200 825.600 ;
        RECT 239.700 821.700 241.500 828.600 ;
        RECT 260.700 821.700 262.500 828.600 ;
        RECT 269.700 821.700 271.500 828.600 ;
        RECT 294.300 821.700 296.100 828.600 ;
        RECT 316.500 821.700 318.300 828.600 ;
        RECT 325.500 821.700 327.300 828.600 ;
        RECT 343.500 821.700 345.300 828.600 ;
        RECT 362.400 821.700 364.200 825.600 ;
        RECT 370.200 821.700 372.000 828.600 ;
        RECT 394.800 821.700 396.600 831.600 ;
        RECT 407.700 821.700 409.500 828.600 ;
        RECT 436.800 821.700 438.600 826.800 ;
        RECT 452.700 821.700 454.500 828.600 ;
        RECT 461.700 821.700 463.500 828.600 ;
        RECT 479.400 821.700 481.200 825.600 ;
        RECT 497.700 821.700 499.500 828.600 ;
        RECT 521.400 821.700 523.200 825.600 ;
        RECT 529.200 821.700 531.000 828.600 ;
        RECT 547.800 821.700 549.600 825.600 ;
        RECT 560.700 821.700 562.500 828.600 ;
        RECT 584.400 821.700 586.200 826.800 ;
        RECT 608.400 821.700 610.200 826.800 ;
        RECT 636.300 821.700 638.100 828.600 ;
        RECT 658.800 821.700 660.600 828.600 ;
        RECT 679.800 821.700 681.600 826.800 ;
        RECT 703.500 821.700 705.300 828.600 ;
        RECT 716.700 821.700 718.500 828.600 ;
        RECT 725.700 821.700 727.500 828.600 ;
        RECT 743.400 821.700 745.200 831.600 ;
        RECT 771.900 821.700 773.700 828.600 ;
        RECT 799.500 821.700 801.300 828.600 ;
        RECT 813.000 821.700 814.800 828.600 ;
        RECT 820.800 821.700 822.600 825.600 ;
        RECT 836.400 821.700 838.200 825.600 ;
        RECT 842.400 821.700 844.200 825.600 ;
        RECT 865.500 821.700 867.300 828.600 ;
        RECT 878.700 821.700 880.500 828.600 ;
        RECT 899.700 821.700 901.500 828.600 ;
        RECT 911.550 821.700 920.550 897.300 ;
        RECT 1.500 819.300 920.550 821.700 ;
        RECT 14.400 815.400 16.200 819.300 ;
        RECT 22.200 812.400 24.000 819.300 ;
        RECT 43.800 814.200 45.600 819.300 ;
        RECT 67.800 814.200 69.600 819.300 ;
        RECT 94.800 809.400 96.600 819.300 ;
        RECT 110.400 815.400 112.200 819.300 ;
        RECT 118.200 812.400 120.000 819.300 ;
        RECT 136.800 815.400 138.600 819.300 ;
        RECT 157.500 812.400 159.300 819.300 ;
        RECT 178.800 814.200 180.600 819.300 ;
        RECT 202.500 812.400 204.300 819.300 ;
        RECT 222.300 812.400 224.100 819.300 ;
        RECT 244.500 812.400 246.300 819.300 ;
        RECT 271.800 809.400 273.600 819.300 ;
        RECT 292.800 814.200 294.600 819.300 ;
        RECT 316.800 814.200 318.600 819.300 ;
        RECT 335.400 815.400 337.200 819.300 ;
        RECT 343.200 812.400 345.000 819.300 ;
        RECT 367.800 809.400 369.600 819.300 ;
        RECT 385.800 815.400 387.600 819.300 ;
        RECT 399.000 812.400 400.800 819.300 ;
        RECT 406.800 815.400 408.600 819.300 ;
        RECT 430.800 814.200 432.600 819.300 ;
        RECT 454.800 814.200 456.600 819.300 ;
        RECT 481.800 809.400 483.600 819.300 ;
        RECT 499.500 812.400 501.300 819.300 ;
        RECT 508.500 812.400 510.300 819.300 ;
        RECT 529.800 814.200 531.600 819.300 ;
        RECT 550.500 812.400 552.300 819.300 ;
        RECT 559.500 812.400 561.300 819.300 ;
        RECT 576.900 812.400 578.700 819.300 ;
        RECT 604.500 812.400 606.300 819.300 ;
        RECT 628.800 809.400 630.600 819.300 ;
        RECT 644.400 815.400 646.200 819.300 ;
        RECT 652.200 812.400 654.000 819.300 ;
        RECT 670.800 815.400 672.600 819.300 ;
        RECT 687.900 812.400 689.700 819.300 ;
        RECT 718.800 809.400 720.600 819.300 ;
        RECT 731.700 812.400 733.500 819.300 ;
        RECT 755.400 815.400 757.200 819.300 ;
        RECT 763.200 812.400 765.000 819.300 ;
        RECT 784.500 812.400 786.300 819.300 ;
        RECT 802.800 815.400 804.600 819.300 ;
        RECT 818.400 814.200 820.200 819.300 ;
        RECT 842.400 814.200 844.200 819.300 ;
        RECT 865.800 815.400 867.600 819.300 ;
        RECT 871.800 815.400 873.600 819.300 ;
        RECT 885.000 812.400 886.800 819.300 ;
        RECT 892.800 815.400 894.600 819.300 ;
        RECT 16.800 743.700 18.600 747.600 ;
        RECT 29.400 743.700 31.200 753.600 ;
        RECT 61.800 743.700 63.600 748.800 ;
        RECT 88.800 743.700 90.600 753.600 ;
        RECT 112.800 743.700 114.600 753.600 ;
        RECT 126.000 743.700 127.800 750.600 ;
        RECT 133.800 743.700 135.600 747.600 ;
        RECT 160.800 743.700 162.600 753.600 ;
        RECT 176.400 743.700 178.200 747.600 ;
        RECT 184.200 743.700 186.000 750.600 ;
        RECT 197.700 743.700 199.500 750.600 ;
        RECT 226.800 743.700 228.600 748.800 ;
        RECT 247.800 743.700 249.600 750.600 ;
        RECT 271.800 743.700 273.600 753.600 ;
        RECT 285.000 743.700 286.800 750.600 ;
        RECT 292.800 743.700 294.600 747.600 ;
        RECT 308.400 743.700 310.200 753.600 ;
        RECT 340.800 743.700 342.600 748.800 ;
        RECT 359.400 743.700 361.200 747.600 ;
        RECT 367.200 743.700 369.000 750.600 ;
        RECT 391.800 743.700 393.600 753.600 ;
        RECT 415.800 743.700 417.600 753.600 ;
        RECT 428.400 743.700 430.200 753.600 ;
        RECT 455.400 743.700 457.200 748.800 ;
        RECT 477.000 743.700 478.800 750.600 ;
        RECT 484.800 743.700 486.600 747.600 ;
        RECT 508.800 743.700 510.600 748.800 ;
        RECT 529.800 743.700 531.600 750.600 ;
        RECT 553.800 743.700 555.600 753.600 ;
        RECT 567.000 743.700 568.800 750.600 ;
        RECT 574.800 743.700 576.600 747.600 ;
        RECT 598.800 743.700 600.600 748.800 ;
        RECT 622.500 743.700 624.300 750.600 ;
        RECT 643.800 743.700 645.600 748.800 ;
        RECT 659.400 743.700 661.200 747.600 ;
        RECT 665.400 743.700 667.200 747.600 ;
        RECT 683.400 743.700 685.200 749.100 ;
        RECT 712.800 743.700 714.600 747.600 ;
        RECT 726.000 743.700 727.800 750.600 ;
        RECT 733.800 743.700 735.600 747.600 ;
        RECT 754.800 743.700 756.600 750.600 ;
        RECT 767.700 743.700 769.500 750.600 ;
        RECT 791.400 743.700 793.200 748.800 ;
        RECT 820.500 743.700 822.300 750.600 ;
        RECT 836.700 743.700 838.500 750.600 ;
        RECT 857.400 743.700 859.200 748.800 ;
        RECT 881.700 743.700 883.500 750.600 ;
        RECT 899.400 743.700 901.200 747.600 ;
        RECT 905.400 743.700 907.200 747.600 ;
        RECT 911.550 743.700 920.550 819.300 ;
        RECT 1.500 741.300 920.550 743.700 ;
        RECT 16.800 737.400 18.600 741.300 ;
        RECT 32.400 736.200 34.200 741.300 ;
        RECT 54.000 734.400 55.800 741.300 ;
        RECT 61.800 737.400 63.600 741.300 ;
        RECT 82.800 737.400 84.600 741.300 ;
        RECT 103.800 736.200 105.600 741.300 ;
        RECT 122.400 736.200 124.200 741.300 ;
        RECT 146.400 736.200 148.200 741.300 ;
        RECT 168.000 734.400 169.800 741.300 ;
        RECT 175.800 737.400 177.600 741.300 ;
        RECT 191.400 737.400 193.200 741.300 ;
        RECT 197.400 737.400 199.200 741.300 ;
        RECT 212.400 737.400 214.200 741.300 ;
        RECT 230.700 734.400 232.500 741.300 ;
        RECT 259.800 736.200 261.600 741.300 ;
        RECT 275.700 734.400 277.500 741.300 ;
        RECT 304.800 736.200 306.600 741.300 ;
        RECT 320.700 734.400 322.500 741.300 ;
        RECT 341.700 734.400 343.500 741.300 ;
        RECT 366.900 734.400 368.700 741.300 ;
        RECT 386.400 731.400 388.200 741.300 ;
        RECT 411.000 734.400 412.800 741.300 ;
        RECT 418.800 737.400 420.600 741.300 ;
        RECT 434.400 737.400 436.200 741.300 ;
        RECT 452.400 734.400 454.200 741.300 ;
        RECT 473.400 736.200 475.200 741.300 ;
        RECT 494.700 734.400 496.500 741.300 ;
        RECT 518.400 736.200 520.200 741.300 ;
        RECT 546.300 734.400 548.100 741.300 ;
        RECT 570.300 734.400 572.100 741.300 ;
        RECT 595.800 736.200 597.600 741.300 ;
        RECT 614.400 736.200 616.200 741.300 ;
        RECT 643.500 734.400 645.300 741.300 ;
        RECT 664.800 736.200 666.600 741.300 ;
        RECT 688.500 734.400 690.300 741.300 ;
        RECT 704.400 736.200 706.200 741.300 ;
        RECT 725.400 737.400 727.200 741.300 ;
        RECT 731.400 737.400 733.200 741.300 ;
        RECT 749.400 736.200 751.200 741.300 ;
        RECT 770.700 734.400 772.500 741.300 ;
        RECT 791.700 734.400 793.500 741.300 ;
        RECT 817.800 734.400 819.600 741.300 ;
        RECT 830.400 737.400 832.200 741.300 ;
        RECT 851.700 734.400 853.500 741.300 ;
        RECT 869.700 734.400 871.500 741.300 ;
        RECT 890.400 731.400 892.200 741.300 ;
        RECT 16.800 665.700 18.600 669.600 ;
        RECT 40.800 665.700 42.600 675.600 ;
        RECT 64.800 665.700 66.600 675.600 ;
        RECT 82.800 665.700 84.600 669.600 ;
        RECT 106.800 665.700 108.600 675.600 ;
        RECT 122.400 665.700 124.200 670.800 ;
        RECT 143.700 665.700 145.500 672.600 ;
        RECT 152.700 665.700 154.500 672.600 ;
        RECT 178.500 665.700 180.300 672.600 ;
        RECT 199.800 665.700 201.600 670.800 ;
        RECT 218.400 665.700 220.200 670.800 ;
        RECT 239.700 665.700 241.500 672.600 ;
        RECT 265.800 665.700 267.600 669.600 ;
        RECT 278.400 665.700 280.200 675.600 ;
        RECT 302.400 665.700 304.200 675.600 ;
        RECT 329.400 665.700 331.200 670.800 ;
        RECT 350.700 665.700 352.500 672.600 ;
        RECT 371.700 665.700 373.500 672.600 ;
        RECT 395.400 665.700 397.200 670.800 ;
        RECT 421.800 665.700 423.600 669.600 ;
        RECT 434.700 665.700 436.500 672.600 ;
        RECT 455.400 665.700 457.200 675.600 ;
        RECT 484.800 665.700 486.600 672.600 ;
        RECT 502.800 665.700 504.600 672.600 ;
        RECT 520.800 665.700 522.600 672.600 ;
        RECT 544.800 665.700 546.600 675.600 ;
        RECT 557.400 665.700 559.200 675.600 ;
        RECT 582.000 665.700 583.800 672.600 ;
        RECT 589.800 665.700 591.600 669.600 ;
        RECT 605.400 665.700 607.200 672.600 ;
        RECT 623.700 665.700 625.500 672.600 ;
        RECT 647.400 665.700 649.200 670.800 ;
        RECT 668.700 665.700 670.500 672.600 ;
        RECT 691.800 665.700 693.600 669.600 ;
        RECT 697.800 665.700 699.600 669.600 ;
        RECT 713.400 665.700 715.200 670.800 ;
        RECT 742.500 665.700 744.300 672.600 ;
        RECT 763.800 665.700 765.600 670.800 ;
        RECT 779.400 665.700 781.200 675.600 ;
        RECT 803.700 665.700 805.500 672.600 ;
        RECT 825.000 665.700 826.800 672.600 ;
        RECT 832.800 665.700 834.600 669.600 ;
        RECT 856.800 665.700 858.600 670.800 ;
        RECT 875.400 665.700 877.200 670.800 ;
        RECT 896.400 665.700 898.200 669.600 ;
        RECT 911.550 665.700 920.550 741.300 ;
        RECT 1.500 663.300 920.550 665.700 ;
        RECT 22.800 653.400 24.600 663.300 ;
        RECT 36.000 656.400 37.800 663.300 ;
        RECT 43.800 659.400 45.600 663.300 ;
        RECT 64.800 659.400 66.600 663.300 ;
        RECT 79.800 659.400 81.600 663.300 ;
        RECT 85.800 659.400 87.600 663.300 ;
        RECT 101.400 659.400 103.200 663.300 ;
        RECT 109.200 656.400 111.000 663.300 ;
        RECT 122.400 653.400 124.200 663.300 ;
        RECT 141.150 659.400 142.950 663.300 ;
        RECT 150.450 659.400 152.250 663.300 ;
        RECT 157.350 659.400 159.150 663.300 ;
        RECT 166.350 659.400 168.150 663.300 ;
        RECT 182.400 659.400 184.200 663.300 ;
        RECT 188.400 659.400 190.200 663.300 ;
        RECT 203.700 656.400 205.500 663.300 ;
        RECT 229.800 659.400 231.600 663.300 ;
        RECT 250.800 658.200 252.600 663.300 ;
        RECT 270.900 656.400 272.700 663.300 ;
        RECT 298.500 656.400 300.300 663.300 ;
        RECT 319.800 658.200 321.600 663.300 ;
        RECT 338.400 658.200 340.200 663.300 ;
        RECT 367.800 658.200 369.600 663.300 ;
        RECT 378.150 659.400 379.950 663.300 ;
        RECT 387.450 659.400 389.250 663.300 ;
        RECT 394.350 659.400 396.150 663.300 ;
        RECT 403.350 659.400 405.150 663.300 ;
        RECT 419.400 653.400 421.200 663.300 ;
        RECT 450.300 656.400 452.100 663.300 ;
        RECT 467.700 656.400 469.500 663.300 ;
        RECT 493.800 659.400 495.600 663.300 ;
        RECT 514.800 658.200 516.600 663.300 ;
        RECT 525.150 659.400 526.950 663.300 ;
        RECT 534.450 659.400 536.250 663.300 ;
        RECT 541.350 659.400 543.150 663.300 ;
        RECT 550.350 659.400 552.150 663.300 ;
        RECT 570.900 656.400 572.700 663.300 ;
        RECT 598.800 658.200 600.600 663.300 ;
        RECT 625.800 653.400 627.600 663.300 ;
        RECT 638.400 659.400 640.200 663.300 ;
        RECT 659.400 658.200 661.200 663.300 ;
        RECT 684.900 656.400 686.700 663.300 ;
        RECT 704.400 659.400 706.200 663.300 ;
        RECT 710.400 659.400 712.200 663.300 ;
        RECT 728.400 658.200 730.200 663.300 ;
        RECT 752.400 658.200 754.200 663.300 ;
        RECT 781.800 658.200 783.600 663.300 ;
        RECT 797.700 656.400 799.500 663.300 ;
        RECT 826.500 656.400 828.300 663.300 ;
        RECT 839.400 662.400 840.600 663.300 ;
        RECT 839.400 659.400 841.200 662.400 ;
        RECT 845.400 659.400 847.200 663.300 ;
        RECT 874.800 653.400 876.600 663.300 ;
        RECT 887.400 653.400 889.200 663.300 ;
        RECT 19.500 587.700 21.300 594.600 ;
        RECT 43.800 587.700 45.600 597.600 ;
        RECT 64.500 587.700 66.300 594.600 ;
        RECT 85.800 587.700 87.600 592.800 ;
        RECT 95.850 587.700 97.650 591.600 ;
        RECT 104.850 587.700 106.650 591.600 ;
        RECT 111.750 587.700 113.550 591.600 ;
        RECT 121.050 587.700 122.850 591.600 ;
        RECT 145.800 587.700 147.600 592.800 ;
        RECT 156.150 587.700 157.950 591.600 ;
        RECT 165.450 587.700 167.250 591.600 ;
        RECT 172.350 587.700 174.150 591.600 ;
        RECT 181.350 587.700 183.150 591.600 ;
        RECT 205.800 587.700 207.600 592.800 ;
        RECT 221.700 587.700 223.500 594.600 ;
        RECT 242.700 587.700 244.500 594.600 ;
        RECT 263.700 587.700 265.500 594.600 ;
        RECT 288.900 587.700 290.700 594.600 ;
        RECT 319.800 587.700 321.600 597.600 ;
        RECT 340.800 587.700 342.600 592.800 ;
        RECT 359.400 587.700 361.200 592.800 ;
        RECT 391.800 587.700 393.600 597.600 ;
        RECT 407.400 587.700 409.200 591.600 ;
        RECT 415.200 587.700 417.000 594.600 ;
        RECT 423.150 587.700 424.950 591.600 ;
        RECT 432.450 587.700 434.250 591.600 ;
        RECT 439.350 587.700 441.150 591.600 ;
        RECT 448.350 587.700 450.150 591.600 ;
        RECT 465.000 587.700 466.800 594.600 ;
        RECT 472.800 587.700 474.600 591.600 ;
        RECT 496.800 587.700 498.600 592.800 ;
        RECT 507.150 587.700 508.950 591.600 ;
        RECT 516.450 587.700 518.250 591.600 ;
        RECT 523.350 587.700 525.150 591.600 ;
        RECT 532.350 587.700 534.150 591.600 ;
        RECT 551.400 587.700 553.200 591.600 ;
        RECT 559.200 587.700 561.000 594.600 ;
        RECT 583.800 587.700 585.600 597.600 ;
        RECT 604.800 587.700 606.600 592.800 ;
        RECT 628.500 587.700 630.300 594.600 ;
        RECT 652.800 587.700 654.600 597.600 ;
        RECT 665.700 587.700 667.500 594.600 ;
        RECT 694.800 587.700 696.600 592.800 ;
        RECT 713.400 587.700 715.200 592.800 ;
        RECT 734.700 587.700 736.500 594.600 ;
        RECT 755.700 587.700 757.500 594.600 ;
        RECT 779.400 587.700 781.200 592.800 ;
        RECT 803.400 587.700 805.200 592.800 ;
        RECT 827.400 587.700 829.200 592.800 ;
        RECT 848.700 587.700 850.500 594.600 ;
        RECT 872.400 587.700 874.200 591.600 ;
        RECT 880.200 587.700 882.000 594.600 ;
        RECT 893.400 587.700 895.200 597.600 ;
        RECT 911.550 587.700 920.550 663.300 ;
        RECT 1.500 585.300 920.550 587.700 ;
        RECT 19.500 578.400 21.300 585.300 ;
        RECT 32.400 575.400 34.200 585.300 ;
        RECT 64.500 578.400 66.300 585.300 ;
        RECT 85.500 578.400 87.300 585.300 ;
        RECT 101.400 581.400 103.200 585.300 ;
        RECT 109.200 578.400 111.000 585.300 ;
        RECT 133.800 575.400 135.600 585.300 ;
        RECT 146.700 578.400 148.500 585.300 ;
        RECT 172.800 581.400 174.600 585.300 ;
        RECT 185.400 581.400 187.200 585.300 ;
        RECT 214.800 575.400 216.600 585.300 ;
        RECT 238.800 575.400 240.600 585.300 ;
        RECT 251.700 578.400 253.500 585.300 ;
        RECT 275.400 581.400 277.200 585.300 ;
        RECT 283.200 578.400 285.000 585.300 ;
        RECT 307.800 575.400 309.600 585.300 ;
        RECT 325.800 581.400 327.600 585.300 ;
        RECT 341.400 581.400 343.200 585.300 ;
        RECT 349.200 578.400 351.000 585.300 ;
        RECT 373.800 575.400 375.600 585.300 ;
        RECT 394.500 578.400 396.300 585.300 ;
        RECT 407.700 578.400 409.500 585.300 ;
        RECT 436.800 580.200 438.600 585.300 ;
        RECT 460.500 578.400 462.300 585.300 ;
        RECT 481.800 580.200 483.600 585.300 ;
        RECT 500.400 580.200 502.200 585.300 ;
        RECT 524.400 581.400 526.200 585.300 ;
        RECT 532.200 578.400 534.000 585.300 ;
        RECT 556.800 575.400 558.600 585.300 ;
        RECT 574.800 581.400 576.600 585.300 ;
        RECT 588.000 578.400 589.800 585.300 ;
        RECT 595.800 581.400 597.600 585.300 ;
        RECT 618.300 578.400 620.100 585.300 ;
        RECT 635.700 578.400 637.500 585.300 ;
        RECT 664.800 580.200 666.600 585.300 ;
        RECT 691.800 575.400 693.600 585.300 ;
        RECT 707.400 581.400 709.200 585.300 ;
        RECT 715.200 578.400 717.000 585.300 ;
        RECT 728.400 575.400 730.200 585.300 ;
        RECT 752.400 581.400 754.200 585.300 ;
        RECT 758.400 581.400 760.200 585.300 ;
        RECT 773.400 581.400 775.200 585.300 ;
        RECT 802.800 575.400 804.600 585.300 ;
        RECT 815.400 575.400 817.200 585.300 ;
        RECT 844.800 581.400 846.600 585.300 ;
        RECT 865.800 580.200 867.600 585.300 ;
        RECT 881.400 581.400 883.200 585.300 ;
        RECT 902.700 578.400 904.500 585.300 ;
        RECT 16.800 509.700 18.600 513.600 ;
        RECT 30.000 509.700 31.800 516.600 ;
        RECT 37.800 509.700 39.600 513.600 ;
        RECT 58.800 509.700 60.600 513.600 ;
        RECT 71.400 509.700 73.200 519.600 ;
        RECT 98.400 509.700 100.200 514.800 ;
        RECT 122.700 509.700 124.500 516.600 ;
        RECT 135.150 509.700 136.950 513.600 ;
        RECT 144.450 509.700 146.250 513.600 ;
        RECT 151.350 509.700 153.150 513.600 ;
        RECT 160.350 509.700 162.150 513.600 ;
        RECT 179.400 509.700 181.200 514.800 ;
        RECT 208.500 509.700 210.300 516.600 ;
        RECT 229.800 509.700 231.600 514.800 ;
        RECT 253.800 509.700 255.600 514.800 ;
        RECT 272.400 509.700 274.200 513.600 ;
        RECT 280.200 509.700 282.000 516.600 ;
        RECT 304.800 509.700 306.600 519.600 ;
        RECT 317.400 509.700 319.200 519.600 ;
        RECT 344.400 509.700 346.200 514.800 ;
        RECT 365.700 509.700 367.500 516.600 ;
        RECT 374.700 509.700 376.500 516.600 ;
        RECT 397.500 509.700 399.300 516.600 ;
        RECT 424.800 509.700 426.600 519.600 ;
        RECT 448.800 509.700 450.600 519.600 ;
        RECT 472.800 509.700 474.600 519.600 ;
        RECT 496.800 509.700 498.600 519.600 ;
        RECT 510.000 509.700 511.800 516.600 ;
        RECT 517.800 509.700 519.600 513.600 ;
        RECT 541.800 509.700 543.600 514.800 ;
        RECT 560.400 509.700 562.200 513.600 ;
        RECT 568.200 509.700 570.000 516.600 ;
        RECT 581.400 509.700 583.200 519.600 ;
        RECT 605.400 509.700 607.200 513.600 ;
        RECT 626.400 509.700 628.200 513.600 ;
        RECT 634.200 509.700 636.000 516.600 ;
        RECT 658.800 509.700 660.600 519.600 ;
        RECT 682.800 509.700 684.600 519.600 ;
        RECT 698.400 509.700 700.200 514.800 ;
        RECT 719.700 509.700 721.500 516.600 ;
        RECT 745.500 509.700 747.300 516.600 ;
        RECT 754.500 509.700 756.300 516.600 ;
        RECT 778.800 509.700 780.600 519.600 ;
        RECT 796.800 509.700 798.600 513.600 ;
        RECT 809.400 509.700 811.200 519.600 ;
        RECT 838.800 509.700 840.600 513.600 ;
        RECT 862.800 509.700 864.600 519.600 ;
        RECT 876.000 509.700 877.800 516.600 ;
        RECT 883.800 509.700 885.600 513.600 ;
        RECT 899.400 509.700 901.200 513.600 ;
        RECT 911.550 509.700 920.550 585.300 ;
        RECT 1.500 507.300 920.550 509.700 ;
        RECT 14.400 503.400 16.200 507.300 ;
        RECT 22.200 500.400 24.000 507.300 ;
        RECT 35.400 497.400 37.200 507.300 ;
        RECT 59.400 503.400 61.200 507.300 ;
        RECT 85.500 500.400 87.300 507.300 ;
        RECT 103.500 500.400 105.300 507.300 ;
        RECT 112.500 500.400 114.300 507.300 ;
        RECT 122.700 500.400 124.500 507.300 ;
        RECT 143.400 506.400 144.600 507.300 ;
        RECT 143.400 503.400 145.200 506.400 ;
        RECT 149.400 503.400 151.200 507.300 ;
        RECT 169.800 500.400 171.600 507.300 ;
        RECT 175.800 500.400 177.600 507.300 ;
        RECT 181.800 500.400 183.600 507.300 ;
        RECT 187.800 500.400 189.600 507.300 ;
        RECT 193.800 500.400 195.600 507.300 ;
        RECT 211.800 503.400 213.600 507.300 ;
        RECT 219.150 503.400 220.950 507.300 ;
        RECT 228.450 503.400 230.250 507.300 ;
        RECT 235.350 503.400 237.150 507.300 ;
        RECT 244.350 503.400 246.150 507.300 ;
        RECT 260.400 503.400 262.200 507.300 ;
        RECT 283.800 503.400 285.600 507.300 ;
        RECT 290.850 503.400 292.650 507.300 ;
        RECT 299.850 503.400 301.650 507.300 ;
        RECT 306.750 503.400 308.550 507.300 ;
        RECT 316.050 503.400 317.850 507.300 ;
        RECT 339.300 500.400 341.100 507.300 ;
        RECT 356.400 497.400 358.200 507.300 ;
        RECT 382.800 503.400 384.600 507.300 ;
        RECT 388.800 503.400 390.600 507.300 ;
        RECT 404.400 503.400 406.200 507.300 ;
        RECT 412.200 500.400 414.000 507.300 ;
        RECT 425.400 497.400 427.200 507.300 ;
        RECT 454.800 503.400 456.600 507.300 ;
        RECT 467.400 497.400 469.200 507.300 ;
        RECT 502.800 497.400 504.600 507.300 ;
        RECT 526.800 497.400 528.600 507.300 ;
        RECT 539.400 503.400 541.200 507.300 ;
        RECT 560.400 502.200 562.200 507.300 ;
        RECT 586.800 503.400 588.600 507.300 ;
        RECT 599.400 497.400 601.200 507.300 ;
        RECT 631.500 500.400 633.300 507.300 ;
        RECT 646.800 503.400 648.600 507.300 ;
        RECT 652.800 503.400 654.600 507.300 ;
        RECT 673.500 500.400 675.300 507.300 ;
        RECT 689.400 502.200 691.200 507.300 ;
        RECT 721.800 497.400 723.600 507.300 ;
        RECT 734.400 503.400 736.200 507.300 ;
        RECT 740.400 503.400 742.200 507.300 ;
        RECT 758.400 503.400 760.200 507.300 ;
        RECT 766.200 500.400 768.000 507.300 ;
        RECT 787.500 500.400 789.300 507.300 ;
        RECT 804.900 500.400 806.700 507.300 ;
        RECT 835.800 497.400 837.600 507.300 ;
        RECT 856.500 500.400 858.300 507.300 ;
        RECT 880.800 497.400 882.600 507.300 ;
        RECT 893.700 500.400 895.500 507.300 ;
        RECT 22.800 431.700 24.600 437.100 ;
        RECT 38.700 431.700 40.500 438.600 ;
        RECT 67.500 431.700 69.300 438.600 ;
        RECT 88.500 431.700 90.300 438.600 ;
        RECT 109.800 431.700 111.600 436.800 ;
        RECT 127.800 431.700 129.600 435.600 ;
        RECT 133.800 431.700 135.600 435.600 ;
        RECT 146.400 431.700 148.200 435.600 ;
        RECT 167.400 431.700 169.200 436.800 ;
        RECT 199.800 431.700 201.600 441.600 ;
        RECT 220.800 431.700 222.600 436.800 ;
        RECT 241.500 431.700 243.300 438.600 ;
        RECT 260.400 431.700 262.200 437.100 ;
        RECT 284.400 431.700 286.200 435.600 ;
        RECT 290.400 431.700 292.200 435.600 ;
        RECT 313.500 431.700 315.300 438.600 ;
        RECT 329.400 431.700 331.200 436.800 ;
        RECT 358.800 431.700 360.600 436.800 ;
        RECT 374.400 431.700 376.200 435.600 ;
        RECT 395.400 431.700 397.200 436.800 ;
        RECT 416.400 431.700 418.200 435.600 ;
        RECT 424.200 431.700 426.000 438.600 ;
        RECT 437.400 431.700 439.200 441.600 ;
        RECT 469.500 431.700 471.300 438.600 ;
        RECT 482.700 431.700 484.500 438.600 ;
        RECT 503.700 431.700 505.500 438.600 ;
        RECT 525.000 431.700 526.800 438.600 ;
        RECT 532.800 431.700 534.600 435.600 ;
        RECT 556.500 431.700 558.300 438.600 ;
        RECT 572.400 431.700 574.200 436.800 ;
        RECT 596.400 431.700 598.200 436.800 ;
        RECT 617.400 431.700 619.200 435.600 ;
        RECT 638.400 431.700 640.200 435.600 ;
        RECT 646.200 431.700 648.000 438.600 ;
        RECT 659.400 431.700 661.200 441.600 ;
        RECT 688.500 431.700 690.300 438.600 ;
        RECT 704.400 431.700 706.200 435.600 ;
        RECT 733.800 431.700 735.600 441.600 ;
        RECT 746.700 431.700 748.500 438.600 ;
        RECT 775.800 431.700 777.600 436.800 ;
        RECT 791.400 431.700 793.200 435.600 ;
        RECT 820.800 431.700 822.600 441.600 ;
        RECT 833.400 431.700 835.200 435.600 ;
        RECT 851.700 431.700 853.500 438.600 ;
        RECT 872.400 432.600 874.200 435.600 ;
        RECT 872.400 431.700 873.600 432.600 ;
        RECT 878.400 431.700 880.200 435.600 ;
        RECT 896.700 431.700 898.500 438.600 ;
        RECT 911.550 431.700 920.550 507.300 ;
        RECT 1.500 429.300 920.550 431.700 ;
        RECT 6.150 425.400 7.950 429.300 ;
        RECT 15.450 425.400 17.250 429.300 ;
        RECT 22.350 425.400 24.150 429.300 ;
        RECT 31.350 425.400 33.150 429.300 ;
        RECT 58.800 423.900 60.600 429.300 ;
        RECT 69.150 425.400 70.950 429.300 ;
        RECT 78.450 425.400 80.250 429.300 ;
        RECT 85.350 425.400 87.150 429.300 ;
        RECT 94.350 425.400 96.150 429.300 ;
        RECT 115.800 425.400 117.600 429.300 ;
        RECT 130.800 425.400 132.600 429.300 ;
        RECT 136.800 425.400 138.600 429.300 ;
        RECT 143.850 425.400 145.650 429.300 ;
        RECT 152.850 425.400 154.650 429.300 ;
        RECT 159.750 425.400 161.550 429.300 ;
        RECT 169.050 425.400 170.850 429.300 ;
        RECT 179.850 425.400 181.650 429.300 ;
        RECT 188.850 425.400 190.650 429.300 ;
        RECT 195.750 425.400 197.550 429.300 ;
        RECT 205.050 425.400 206.850 429.300 ;
        RECT 216.150 425.400 217.950 429.300 ;
        RECT 225.450 425.400 227.250 429.300 ;
        RECT 232.350 425.400 234.150 429.300 ;
        RECT 241.350 425.400 243.150 429.300 ;
        RECT 257.400 425.400 259.200 429.300 ;
        RECT 275.400 425.400 277.200 429.300 ;
        RECT 281.400 425.400 283.200 429.300 ;
        RECT 298.800 425.400 300.600 429.300 ;
        RECT 304.800 425.400 306.600 429.300 ;
        RECT 317.400 425.400 319.200 429.300 ;
        RECT 338.700 422.400 340.500 429.300 ;
        RECT 364.500 422.400 366.300 429.300 ;
        RECT 377.700 422.400 379.500 429.300 ;
        RECT 400.800 425.400 402.600 429.300 ;
        RECT 406.800 425.400 408.600 429.300 ;
        RECT 422.400 424.200 424.200 429.300 ;
        RECT 446.700 422.400 448.500 429.300 ;
        RECT 469.500 422.400 471.300 429.300 ;
        RECT 488.400 424.200 490.200 429.300 ;
        RECT 520.800 419.400 522.600 429.300 ;
        RECT 544.800 419.400 546.600 429.300 ;
        RECT 565.500 422.400 567.300 429.300 ;
        RECT 589.800 419.400 591.600 429.300 ;
        RECT 604.800 425.400 606.600 429.300 ;
        RECT 622.800 425.400 624.600 429.300 ;
        RECT 638.400 424.200 640.200 429.300 ;
        RECT 659.400 425.400 661.200 429.300 ;
        RECT 682.800 425.400 684.600 429.300 ;
        RECT 697.800 425.400 699.600 429.300 ;
        RECT 703.800 425.400 705.600 429.300 ;
        RECT 719.400 424.200 721.200 429.300 ;
        RECT 745.800 425.400 747.600 429.300 ;
        RECT 760.800 425.400 762.600 429.300 ;
        RECT 766.800 425.400 768.600 429.300 ;
        RECT 781.800 425.400 783.600 429.300 ;
        RECT 787.800 425.400 789.600 429.300 ;
        RECT 803.400 424.200 805.200 429.300 ;
        RECT 824.400 425.400 826.200 429.300 ;
        RECT 830.400 425.400 832.200 429.300 ;
        RECT 845.400 425.400 847.200 429.300 ;
        RECT 851.400 425.400 853.200 429.300 ;
        RECT 873.300 422.400 875.100 429.300 ;
        RECT 890.400 425.400 892.200 429.300 ;
        RECT 896.400 425.400 898.200 429.300 ;
        RECT 5.850 353.700 7.650 357.600 ;
        RECT 14.850 353.700 16.650 357.600 ;
        RECT 21.750 353.700 23.550 357.600 ;
        RECT 31.050 353.700 32.850 357.600 ;
        RECT 42.150 353.700 43.950 357.600 ;
        RECT 51.450 353.700 53.250 357.600 ;
        RECT 58.350 353.700 60.150 357.600 ;
        RECT 67.350 353.700 69.150 357.600 ;
        RECT 88.800 353.700 90.600 357.600 ;
        RECT 104.400 353.700 106.200 357.600 ;
        RECT 112.200 353.700 114.000 360.600 ;
        RECT 127.800 353.700 129.600 357.600 ;
        RECT 133.800 353.700 135.600 357.600 ;
        RECT 146.400 354.600 148.200 357.600 ;
        RECT 146.400 353.700 147.600 354.600 ;
        RECT 152.400 353.700 154.200 357.600 ;
        RECT 170.700 353.700 172.500 360.600 ;
        RECT 191.700 353.700 193.500 360.600 ;
        RECT 220.800 353.700 222.600 358.800 ;
        RECT 236.400 353.700 238.200 357.600 ;
        RECT 242.400 353.700 244.200 357.600 ;
        RECT 259.800 353.700 261.600 357.600 ;
        RECT 265.800 353.700 267.600 357.600 ;
        RECT 286.500 353.700 288.300 360.600 ;
        RECT 302.400 353.700 304.200 358.800 ;
        RECT 323.700 353.700 325.500 360.600 ;
        RECT 352.500 353.700 354.300 360.600 ;
        RECT 367.800 353.700 369.600 357.600 ;
        RECT 373.800 353.700 375.600 357.600 ;
        RECT 389.400 353.700 391.200 357.600 ;
        RECT 397.200 353.700 399.000 360.600 ;
        RECT 404.850 353.700 406.650 357.600 ;
        RECT 413.850 353.700 415.650 357.600 ;
        RECT 420.750 353.700 422.550 357.600 ;
        RECT 430.050 353.700 431.850 357.600 ;
        RECT 449.400 353.700 451.200 358.800 ;
        RECT 471.000 353.700 472.800 360.600 ;
        RECT 478.800 353.700 480.600 357.600 ;
        RECT 489.150 353.700 490.950 357.600 ;
        RECT 498.450 353.700 500.250 357.600 ;
        RECT 505.350 353.700 507.150 357.600 ;
        RECT 514.350 353.700 516.150 357.600 ;
        RECT 530.400 353.700 532.200 357.600 ;
        RECT 536.400 353.700 538.200 357.600 ;
        RECT 559.500 353.700 561.300 360.600 ;
        RECT 580.800 353.700 582.600 358.800 ;
        RECT 596.400 353.700 598.200 357.600 ;
        RECT 608.850 353.700 610.650 357.600 ;
        RECT 617.850 353.700 619.650 357.600 ;
        RECT 624.750 353.700 626.550 357.600 ;
        RECT 634.050 353.700 635.850 357.600 ;
        RECT 653.400 353.700 655.200 359.100 ;
        RECT 677.400 353.700 679.200 357.600 ;
        RECT 683.400 353.700 685.200 357.600 ;
        RECT 699.000 353.700 700.800 360.600 ;
        RECT 706.800 353.700 708.600 357.600 ;
        RECT 723.000 353.700 724.800 360.600 ;
        RECT 730.800 353.700 732.600 357.600 ;
        RECT 741.150 353.700 742.950 357.600 ;
        RECT 750.450 353.700 752.250 357.600 ;
        RECT 757.350 353.700 759.150 357.600 ;
        RECT 766.350 353.700 768.150 357.600 ;
        RECT 782.700 353.700 784.500 360.600 ;
        RECT 791.700 353.700 793.500 360.600 ;
        RECT 809.700 353.700 811.500 360.600 ;
        RECT 835.800 353.700 837.600 357.600 ;
        RECT 841.800 354.600 843.600 357.600 ;
        RECT 842.400 353.700 843.600 354.600 ;
        RECT 857.400 353.700 859.200 358.800 ;
        RECT 873.150 353.700 874.950 357.600 ;
        RECT 882.450 353.700 884.250 357.600 ;
        RECT 889.350 353.700 891.150 357.600 ;
        RECT 898.350 353.700 900.150 357.600 ;
        RECT 911.550 353.700 920.550 429.300 ;
        RECT 1.500 351.300 920.550 353.700 ;
        RECT 11.400 347.400 13.200 351.300 ;
        RECT 34.800 347.400 36.600 351.300 ;
        RECT 52.800 347.400 54.600 351.300 ;
        RECT 67.800 347.400 69.600 351.300 ;
        RECT 73.800 347.400 75.600 351.300 ;
        RECT 88.800 347.400 90.600 351.300 ;
        RECT 94.800 347.400 96.600 351.300 ;
        RECT 112.800 347.400 114.600 351.300 ;
        RECT 119.850 347.400 121.650 351.300 ;
        RECT 128.850 347.400 130.650 351.300 ;
        RECT 135.750 347.400 137.550 351.300 ;
        RECT 145.050 347.400 146.850 351.300 ;
        RECT 169.800 346.200 171.600 351.300 ;
        RECT 180.150 347.400 181.950 351.300 ;
        RECT 189.450 347.400 191.250 351.300 ;
        RECT 196.350 347.400 198.150 351.300 ;
        RECT 205.350 347.400 207.150 351.300 ;
        RECT 221.400 347.400 223.200 351.300 ;
        RECT 242.400 346.200 244.200 351.300 ;
        RECT 266.700 344.400 268.500 351.300 ;
        RECT 284.700 344.400 286.500 351.300 ;
        RECT 310.500 344.400 312.300 351.300 ;
        RECT 331.500 344.400 333.300 351.300 ;
        RECT 349.800 347.400 351.600 351.300 ;
        RECT 355.800 347.400 357.600 351.300 ;
        RECT 362.850 347.400 364.650 351.300 ;
        RECT 371.850 347.400 373.650 351.300 ;
        RECT 378.750 347.400 380.550 351.300 ;
        RECT 388.050 347.400 389.850 351.300 ;
        RECT 406.800 347.400 408.600 351.300 ;
        RECT 412.800 347.400 414.600 351.300 ;
        RECT 428.400 347.400 430.200 351.300 ;
        RECT 436.200 344.400 438.000 351.300 ;
        RECT 444.150 347.400 445.950 351.300 ;
        RECT 453.450 347.400 455.250 351.300 ;
        RECT 460.350 347.400 462.150 351.300 ;
        RECT 469.350 347.400 471.150 351.300 ;
        RECT 486.000 344.400 487.800 351.300 ;
        RECT 493.800 347.400 495.600 351.300 ;
        RECT 511.800 347.400 513.600 351.300 ;
        RECT 517.800 347.400 519.600 351.300 ;
        RECT 524.850 347.400 526.650 351.300 ;
        RECT 533.850 347.400 535.650 351.300 ;
        RECT 540.750 347.400 542.550 351.300 ;
        RECT 550.050 347.400 551.850 351.300 ;
        RECT 561.150 347.400 562.950 351.300 ;
        RECT 570.450 347.400 572.250 351.300 ;
        RECT 577.350 347.400 579.150 351.300 ;
        RECT 586.350 347.400 588.150 351.300 ;
        RECT 602.400 347.400 604.200 351.300 ;
        RECT 608.400 347.400 610.200 351.300 ;
        RECT 623.400 347.400 625.200 351.300 ;
        RECT 641.400 347.400 643.200 351.300 ;
        RECT 647.400 347.400 649.200 351.300 ;
        RECT 663.000 344.400 664.800 351.300 ;
        RECT 670.800 347.400 672.600 351.300 ;
        RECT 686.700 344.400 688.500 351.300 ;
        RECT 695.700 344.400 697.500 351.300 ;
        RECT 713.400 350.400 714.600 351.300 ;
        RECT 713.400 347.400 715.200 350.400 ;
        RECT 719.400 347.400 721.200 351.300 ;
        RECT 732.150 347.400 733.950 351.300 ;
        RECT 741.450 347.400 743.250 351.300 ;
        RECT 748.350 347.400 750.150 351.300 ;
        RECT 757.350 347.400 759.150 351.300 ;
        RECT 773.400 347.400 775.200 351.300 ;
        RECT 793.800 347.400 795.600 351.300 ;
        RECT 799.800 347.400 801.600 351.300 ;
        RECT 812.400 347.400 814.200 351.300 ;
        RECT 838.500 344.400 840.300 351.300 ;
        RECT 851.400 347.400 853.200 351.300 ;
        RECT 880.800 345.900 882.600 351.300 ;
        RECT 901.800 347.400 903.600 351.300 ;
        RECT 13.800 275.700 15.600 279.600 ;
        RECT 19.800 275.700 21.600 279.600 ;
        RECT 43.800 275.700 45.600 285.600 ;
        RECT 64.800 275.700 66.600 280.800 ;
        RECT 85.800 275.700 87.600 279.600 ;
        RECT 101.400 275.700 103.200 280.800 ;
        RECT 122.700 275.700 124.500 282.600 ;
        RECT 143.400 275.700 145.200 279.600 ;
        RECT 155.850 275.700 157.650 279.600 ;
        RECT 164.850 275.700 166.650 279.600 ;
        RECT 171.750 275.700 173.550 279.600 ;
        RECT 181.050 275.700 182.850 279.600 ;
        RECT 200.400 275.700 202.200 280.800 ;
        RECT 221.700 275.700 223.500 282.600 ;
        RECT 244.800 275.700 246.600 279.600 ;
        RECT 250.800 275.700 252.600 279.600 ;
        RECT 257.850 275.700 259.650 279.600 ;
        RECT 266.850 275.700 268.650 279.600 ;
        RECT 273.750 275.700 275.550 279.600 ;
        RECT 283.050 275.700 284.850 279.600 ;
        RECT 302.400 275.700 304.200 279.600 ;
        RECT 310.200 275.700 312.000 282.600 ;
        RECT 325.800 275.700 327.600 282.600 ;
        RECT 331.800 275.700 333.600 282.600 ;
        RECT 337.800 275.700 339.600 282.600 ;
        RECT 343.800 275.700 345.600 282.600 ;
        RECT 349.800 275.700 351.600 282.600 ;
        RECT 363.000 275.700 364.800 282.600 ;
        RECT 370.800 275.700 372.600 279.600 ;
        RECT 381.150 275.700 382.950 279.600 ;
        RECT 390.450 275.700 392.250 279.600 ;
        RECT 397.350 275.700 399.150 279.600 ;
        RECT 406.350 275.700 408.150 279.600 ;
        RECT 416.850 275.700 418.650 279.600 ;
        RECT 425.850 275.700 427.650 279.600 ;
        RECT 432.750 275.700 434.550 279.600 ;
        RECT 442.050 275.700 443.850 279.600 ;
        RECT 463.800 275.700 465.600 279.600 ;
        RECT 470.850 275.700 472.650 279.600 ;
        RECT 479.850 275.700 481.650 279.600 ;
        RECT 486.750 275.700 488.550 279.600 ;
        RECT 496.050 275.700 497.850 279.600 ;
        RECT 512.700 275.700 514.500 282.600 ;
        RECT 527.850 275.700 529.650 279.600 ;
        RECT 536.850 275.700 538.650 279.600 ;
        RECT 543.750 275.700 545.550 279.600 ;
        RECT 553.050 275.700 554.850 279.600 ;
        RECT 571.800 275.700 573.600 282.600 ;
        RECT 577.800 275.700 579.600 282.600 ;
        RECT 583.800 275.700 585.600 282.600 ;
        RECT 589.800 275.700 591.600 282.600 ;
        RECT 595.800 275.700 597.600 282.600 ;
        RECT 611.400 275.700 613.200 280.800 ;
        RECT 627.150 275.700 628.950 279.600 ;
        RECT 636.450 275.700 638.250 279.600 ;
        RECT 643.350 275.700 645.150 279.600 ;
        RECT 652.350 275.700 654.150 279.600 ;
        RECT 668.700 275.700 670.500 282.600 ;
        RECT 683.850 275.700 685.650 279.600 ;
        RECT 692.850 275.700 694.650 279.600 ;
        RECT 699.750 275.700 701.550 279.600 ;
        RECT 709.050 275.700 710.850 279.600 ;
        RECT 725.700 275.700 727.500 282.600 ;
        RECT 741.150 275.700 742.950 279.600 ;
        RECT 750.450 275.700 752.250 279.600 ;
        RECT 757.350 275.700 759.150 279.600 ;
        RECT 766.350 275.700 768.150 279.600 ;
        RECT 790.800 275.700 792.600 280.800 ;
        RECT 808.800 275.700 810.600 279.600 ;
        RECT 814.800 275.700 816.600 279.600 ;
        RECT 822.150 275.700 823.950 279.600 ;
        RECT 831.450 275.700 833.250 279.600 ;
        RECT 838.350 275.700 840.150 279.600 ;
        RECT 847.350 275.700 849.150 279.600 ;
        RECT 863.400 275.700 865.200 282.600 ;
        RECT 869.400 275.700 871.200 282.600 ;
        RECT 875.400 275.700 877.200 282.600 ;
        RECT 881.400 275.700 883.200 282.600 ;
        RECT 887.400 275.700 889.200 282.600 ;
        RECT 911.550 275.700 920.550 351.300 ;
        RECT 1.500 273.300 920.550 275.700 ;
        RECT 13.800 269.400 15.600 273.300 ;
        RECT 19.800 269.400 21.600 273.300 ;
        RECT 37.800 269.400 39.600 273.300 ;
        RECT 44.850 269.400 46.650 273.300 ;
        RECT 53.850 269.400 55.650 273.300 ;
        RECT 60.750 269.400 62.550 273.300 ;
        RECT 70.050 269.400 71.850 273.300 ;
        RECT 89.400 268.200 91.200 273.300 ;
        RECT 112.800 269.400 114.600 273.300 ;
        RECT 118.800 269.400 120.600 273.300 ;
        RECT 136.800 269.400 138.600 273.300 ;
        RECT 143.850 269.400 145.650 273.300 ;
        RECT 152.850 269.400 154.650 273.300 ;
        RECT 159.750 269.400 161.550 273.300 ;
        RECT 169.050 269.400 170.850 273.300 ;
        RECT 188.400 268.200 190.200 273.300 ;
        RECT 209.400 269.400 211.200 273.300 ;
        RECT 235.500 266.400 237.300 273.300 ;
        RECT 248.700 266.400 250.500 273.300 ;
        RECT 277.800 268.200 279.600 273.300 ;
        RECT 287.850 269.400 289.650 273.300 ;
        RECT 296.850 269.400 298.650 273.300 ;
        RECT 303.750 269.400 305.550 273.300 ;
        RECT 313.050 269.400 314.850 273.300 ;
        RECT 337.800 268.200 339.600 273.300 ;
        RECT 356.400 268.200 358.200 273.300 ;
        RECT 385.800 268.200 387.600 273.300 ;
        RECT 401.400 269.400 403.200 273.300 ;
        RECT 424.800 266.400 426.600 273.300 ;
        RECT 439.800 269.400 441.600 273.300 ;
        RECT 445.800 269.400 447.600 273.300 ;
        RECT 460.800 269.400 462.600 273.300 ;
        RECT 466.800 269.400 468.600 273.300 ;
        RECT 479.400 269.400 481.200 273.300 ;
        RECT 500.400 268.200 502.200 273.300 ;
        RECT 524.700 266.400 526.500 273.300 ;
        RECT 537.150 269.400 538.950 273.300 ;
        RECT 546.450 269.400 548.250 273.300 ;
        RECT 553.350 269.400 555.150 273.300 ;
        RECT 562.350 269.400 564.150 273.300 ;
        RECT 581.400 268.200 583.200 273.300 ;
        RECT 602.700 266.400 604.500 273.300 ;
        RECT 623.400 269.400 625.200 273.300 ;
        RECT 629.400 269.400 631.200 273.300 ;
        RECT 644.400 266.400 646.200 273.300 ;
        RECT 650.400 266.400 652.200 273.300 ;
        RECT 656.400 266.400 658.200 273.300 ;
        RECT 662.400 266.400 664.200 273.300 ;
        RECT 668.400 266.400 670.200 273.300 ;
        RECT 683.400 269.400 685.200 273.300 ;
        RECT 704.400 268.200 706.200 273.300 ;
        RECT 733.500 266.400 735.300 273.300 ;
        RECT 754.500 266.400 756.300 273.300 ;
        RECT 775.500 266.400 777.300 273.300 ;
        RECT 791.400 268.200 793.200 273.300 ;
        RECT 820.800 268.200 822.600 273.300 ;
        RECT 841.800 269.400 843.600 273.300 ;
        RECT 854.400 269.400 856.200 273.300 ;
        RECT 860.400 269.400 862.200 273.300 ;
        RECT 875.400 269.400 877.200 273.300 ;
        RECT 881.400 269.400 883.200 273.300 ;
        RECT 899.700 266.400 901.500 273.300 ;
        RECT 19.500 197.700 21.300 204.600 ;
        RECT 40.800 197.700 42.600 202.800 ;
        RECT 58.800 197.700 60.600 201.600 ;
        RECT 64.800 197.700 66.600 201.600 ;
        RECT 79.800 197.700 81.600 201.600 ;
        RECT 85.800 197.700 87.600 201.600 ;
        RECT 92.850 197.700 94.650 201.600 ;
        RECT 101.850 197.700 103.650 201.600 ;
        RECT 108.750 197.700 110.550 201.600 ;
        RECT 118.050 197.700 119.850 201.600 ;
        RECT 137.400 197.700 139.200 202.800 ;
        RECT 158.700 197.700 160.500 204.600 ;
        RECT 173.850 197.700 175.650 201.600 ;
        RECT 182.850 197.700 184.650 201.600 ;
        RECT 189.750 197.700 191.550 201.600 ;
        RECT 199.050 197.700 200.850 201.600 ;
        RECT 223.800 197.700 225.600 202.800 ;
        RECT 247.800 197.700 249.600 202.800 ;
        RECT 266.400 197.700 268.200 202.800 ;
        RECT 289.800 197.700 291.600 201.600 ;
        RECT 295.800 197.700 297.600 201.600 ;
        RECT 316.800 197.700 318.600 202.800 ;
        RECT 337.800 197.700 339.600 201.600 ;
        RECT 347.700 197.700 349.500 204.600 ;
        RECT 362.850 197.700 364.650 201.600 ;
        RECT 371.850 197.700 373.650 201.600 ;
        RECT 378.750 197.700 380.550 201.600 ;
        RECT 388.050 197.700 389.850 201.600 ;
        RECT 407.400 197.700 409.200 201.600 ;
        RECT 415.200 197.700 417.000 204.600 ;
        RECT 428.400 197.700 430.200 201.600 ;
        RECT 434.400 197.700 436.200 201.600 ;
        RECT 450.000 197.700 451.800 204.600 ;
        RECT 457.800 197.700 459.600 201.600 ;
        RECT 468.150 197.700 469.950 201.600 ;
        RECT 477.450 197.700 479.250 201.600 ;
        RECT 484.350 197.700 486.150 201.600 ;
        RECT 493.350 197.700 495.150 201.600 ;
        RECT 509.400 197.700 511.200 201.600 ;
        RECT 515.400 197.700 517.200 201.600 ;
        RECT 538.500 197.700 540.300 204.600 ;
        RECT 559.800 197.700 561.600 202.800 ;
        RECT 570.150 197.700 571.950 201.600 ;
        RECT 579.450 197.700 581.250 201.600 ;
        RECT 586.350 197.700 588.150 201.600 ;
        RECT 595.350 197.700 597.150 201.600 ;
        RECT 611.400 197.700 613.200 201.600 ;
        RECT 632.400 197.700 634.200 202.800 ;
        RECT 661.800 197.700 663.600 202.800 ;
        RECT 677.400 197.700 679.200 201.600 ;
        RECT 683.400 197.700 685.200 201.600 ;
        RECT 698.400 197.700 700.200 201.600 ;
        RECT 704.400 197.700 706.200 201.600 ;
        RECT 722.400 197.700 724.200 202.800 ;
        RECT 751.500 197.700 753.300 204.600 ;
        RECT 764.700 197.700 766.500 204.600 ;
        RECT 779.850 197.700 781.650 201.600 ;
        RECT 788.850 197.700 790.650 201.600 ;
        RECT 795.750 197.700 797.550 201.600 ;
        RECT 805.050 197.700 806.850 201.600 ;
        RECT 815.850 197.700 817.650 201.600 ;
        RECT 824.850 197.700 826.650 201.600 ;
        RECT 831.750 197.700 833.550 201.600 ;
        RECT 841.050 197.700 842.850 201.600 ;
        RECT 852.150 197.700 853.950 201.600 ;
        RECT 861.450 197.700 863.250 201.600 ;
        RECT 868.350 197.700 870.150 201.600 ;
        RECT 877.350 197.700 879.150 201.600 ;
        RECT 896.400 197.700 898.200 201.600 ;
        RECT 904.200 197.700 906.000 204.600 ;
        RECT 911.550 197.700 920.550 273.300 ;
        RECT 1.500 195.300 920.550 197.700 ;
        RECT 13.800 191.400 15.600 195.300 ;
        RECT 19.800 191.400 21.600 195.300 ;
        RECT 35.400 190.200 37.200 195.300 ;
        RECT 56.400 191.400 58.200 195.300 ;
        RECT 74.700 188.400 76.500 195.300 ;
        RECT 95.400 191.400 97.200 195.300 ;
        RECT 101.400 191.400 103.200 195.300 ;
        RECT 116.400 191.400 118.200 195.300 ;
        RECT 134.400 191.400 136.200 195.300 ;
        RECT 146.850 191.400 148.650 195.300 ;
        RECT 155.850 191.400 157.650 195.300 ;
        RECT 162.750 191.400 164.550 195.300 ;
        RECT 172.050 191.400 173.850 195.300 ;
        RECT 191.400 190.200 193.200 195.300 ;
        RECT 214.800 188.400 216.600 195.300 ;
        RECT 220.800 188.400 222.600 195.300 ;
        RECT 226.800 188.400 228.600 195.300 ;
        RECT 232.800 188.400 234.600 195.300 ;
        RECT 238.800 188.400 240.600 195.300 ;
        RECT 259.500 188.400 261.300 195.300 ;
        RECT 277.500 188.400 279.300 195.300 ;
        RECT 287.850 191.400 289.650 195.300 ;
        RECT 296.850 191.400 298.650 195.300 ;
        RECT 303.750 191.400 305.550 195.300 ;
        RECT 313.050 191.400 314.850 195.300 ;
        RECT 332.400 190.200 334.200 195.300 ;
        RECT 353.700 188.400 355.500 195.300 ;
        RECT 376.800 188.400 378.600 195.300 ;
        RECT 382.800 188.400 384.600 195.300 ;
        RECT 388.800 188.400 390.600 195.300 ;
        RECT 394.800 188.400 396.600 195.300 ;
        RECT 400.800 188.400 402.600 195.300 ;
        RECT 413.700 188.400 415.500 195.300 ;
        RECT 434.400 191.400 436.200 195.300 ;
        RECT 452.400 188.400 454.200 195.300 ;
        RECT 458.400 188.400 460.200 195.300 ;
        RECT 464.400 188.400 466.200 195.300 ;
        RECT 470.400 188.400 472.200 195.300 ;
        RECT 476.400 188.400 478.200 195.300 ;
        RECT 499.500 188.400 501.300 195.300 ;
        RECT 512.700 188.400 514.500 195.300 ;
        RECT 527.850 191.400 529.650 195.300 ;
        RECT 536.850 191.400 538.650 195.300 ;
        RECT 543.750 191.400 545.550 195.300 ;
        RECT 553.050 191.400 554.850 195.300 ;
        RECT 574.800 191.400 576.600 195.300 ;
        RECT 590.400 191.400 592.200 195.300 ;
        RECT 598.200 188.400 600.000 195.300 ;
        RECT 613.800 191.400 615.600 195.300 ;
        RECT 619.800 191.400 621.600 195.300 ;
        RECT 639.300 188.400 641.100 195.300 ;
        RECT 657.000 188.400 658.800 195.300 ;
        RECT 664.800 191.400 666.600 195.300 ;
        RECT 680.400 191.400 682.200 195.300 ;
        RECT 686.400 191.400 688.200 195.300 ;
        RECT 703.800 191.400 705.600 195.300 ;
        RECT 709.800 191.400 711.600 195.300 ;
        RECT 726.900 188.400 728.700 195.300 ;
        RECT 751.800 191.400 753.600 195.300 ;
        RECT 772.800 190.200 774.600 195.300 ;
        RECT 788.400 191.400 790.200 195.300 ;
        RECT 794.400 191.400 796.200 195.300 ;
        RECT 820.800 185.400 822.600 195.300 ;
        RECT 833.400 191.400 835.200 195.300 ;
        RECT 851.400 191.400 853.200 195.300 ;
        RECT 871.800 191.400 873.600 195.300 ;
        RECT 877.800 191.400 879.600 195.300 ;
        RECT 895.800 191.400 897.600 195.300 ;
        RECT 14.400 119.700 16.200 123.600 ;
        RECT 22.200 119.700 24.000 126.600 ;
        RECT 35.700 119.700 37.500 126.600 ;
        RECT 56.400 119.700 58.200 129.600 ;
        RECT 81.000 119.700 82.800 126.600 ;
        RECT 88.800 119.700 90.600 123.600 ;
        RECT 108.900 119.700 110.700 126.600 ;
        RECT 128.400 119.700 130.200 123.600 ;
        RECT 134.400 119.700 136.200 123.600 ;
        RECT 151.800 119.700 153.600 123.600 ;
        RECT 157.800 119.700 159.600 123.600 ;
        RECT 170.400 119.700 172.200 123.600 ;
        RECT 191.400 119.700 193.200 124.800 ;
        RECT 215.400 119.700 217.200 124.800 ;
        RECT 231.150 119.700 232.950 123.600 ;
        RECT 240.450 119.700 242.250 123.600 ;
        RECT 247.350 119.700 249.150 123.600 ;
        RECT 256.350 119.700 258.150 123.600 ;
        RECT 267.150 119.700 268.950 123.600 ;
        RECT 276.450 119.700 278.250 123.600 ;
        RECT 283.350 119.700 285.150 123.600 ;
        RECT 292.350 119.700 294.150 123.600 ;
        RECT 303.150 119.700 304.950 123.600 ;
        RECT 312.450 119.700 314.250 123.600 ;
        RECT 319.350 119.700 321.150 123.600 ;
        RECT 328.350 119.700 330.150 123.600 ;
        RECT 352.800 119.700 354.600 124.800 ;
        RECT 368.400 119.700 370.200 123.600 ;
        RECT 391.800 119.700 393.600 123.600 ;
        RECT 406.800 119.700 408.600 123.600 ;
        RECT 412.800 119.700 414.600 123.600 ;
        RECT 425.400 119.700 427.200 123.600 ;
        RECT 431.400 119.700 433.200 123.600 ;
        RECT 447.000 119.700 448.800 126.600 ;
        RECT 454.800 119.700 456.600 123.600 ;
        RECT 478.800 119.700 480.600 124.800 ;
        RECT 494.400 119.700 496.200 123.600 ;
        RECT 500.400 119.700 502.200 123.600 ;
        RECT 515.700 119.700 517.500 126.600 ;
        RECT 544.500 119.700 546.300 126.600 ;
        RECT 565.800 119.700 567.600 124.800 ;
        RECT 589.500 119.700 591.300 126.600 ;
        RECT 607.800 119.700 609.600 123.600 ;
        RECT 623.400 119.700 625.200 124.800 ;
        RECT 652.500 119.700 654.300 126.600 ;
        RECT 659.850 119.700 661.650 123.600 ;
        RECT 668.850 119.700 670.650 123.600 ;
        RECT 675.750 119.700 677.550 123.600 ;
        RECT 685.050 119.700 686.850 123.600 ;
        RECT 706.500 119.700 708.300 126.600 ;
        RECT 725.400 119.700 727.200 124.800 ;
        RECT 754.500 119.700 756.300 126.600 ;
        RECT 775.800 119.700 777.600 124.800 ;
        RECT 799.800 119.700 801.600 124.800 ;
        RECT 818.400 119.700 820.200 124.800 ;
        RECT 847.800 119.700 849.600 124.800 ;
        RECT 863.400 119.700 865.200 123.600 ;
        RECT 884.400 119.700 886.200 124.800 ;
        RECT 911.550 119.700 920.550 195.300 ;
        RECT 1.500 117.300 920.550 119.700 ;
        RECT 15.900 110.400 17.700 117.300 ;
        RECT 36.000 110.400 37.800 117.300 ;
        RECT 43.800 113.400 45.600 117.300 ;
        RECT 61.800 113.400 63.600 117.300 ;
        RECT 67.800 113.400 69.600 117.300 ;
        RECT 88.800 112.200 90.600 117.300 ;
        RECT 109.800 113.400 111.600 117.300 ;
        RECT 130.800 112.200 132.600 117.300 ;
        RECT 146.400 113.400 148.200 117.300 ;
        RECT 152.400 113.400 154.200 117.300 ;
        RECT 161.850 113.400 163.650 117.300 ;
        RECT 170.850 113.400 172.650 117.300 ;
        RECT 177.750 113.400 179.550 117.300 ;
        RECT 187.050 113.400 188.850 117.300 ;
        RECT 203.400 113.400 205.200 117.300 ;
        RECT 209.400 113.400 211.200 117.300 ;
        RECT 232.500 110.400 234.300 117.300 ;
        RECT 248.400 112.200 250.200 117.300 ;
        RECT 269.700 110.400 271.500 117.300 ;
        RECT 295.500 110.400 297.300 117.300 ;
        RECT 304.500 110.400 306.300 117.300 ;
        RECT 322.500 110.400 324.300 117.300 ;
        RECT 340.800 110.400 342.600 117.300 ;
        RECT 346.800 110.400 348.600 117.300 ;
        RECT 352.800 110.400 354.600 117.300 ;
        RECT 370.800 113.400 372.600 117.300 ;
        RECT 391.800 112.200 393.600 117.300 ;
        RECT 409.800 113.400 411.600 117.300 ;
        RECT 415.800 113.400 417.600 117.300 ;
        RECT 428.400 113.400 430.200 117.300 ;
        RECT 450.900 110.400 452.700 117.300 ;
        RECT 473.400 112.200 475.200 117.300 ;
        RECT 502.500 110.400 504.300 117.300 ;
        RECT 510.150 113.400 511.950 117.300 ;
        RECT 519.450 113.400 521.250 117.300 ;
        RECT 526.350 113.400 528.150 117.300 ;
        RECT 535.350 113.400 537.150 117.300 ;
        RECT 554.400 112.200 556.200 117.300 ;
        RECT 570.150 113.400 571.950 117.300 ;
        RECT 579.450 113.400 581.250 117.300 ;
        RECT 586.350 113.400 588.150 117.300 ;
        RECT 595.350 113.400 597.150 117.300 ;
        RECT 611.400 113.400 613.200 117.300 ;
        RECT 617.400 113.400 619.200 117.300 ;
        RECT 632.400 107.400 634.200 117.300 ;
        RECT 659.400 112.200 661.200 117.300 ;
        RECT 682.800 113.400 684.600 117.300 ;
        RECT 688.800 113.400 690.600 117.300 ;
        RECT 701.400 116.400 702.600 117.300 ;
        RECT 701.400 113.400 703.200 116.400 ;
        RECT 707.400 113.400 709.200 117.300 ;
        RECT 733.800 112.200 735.600 117.300 ;
        RECT 752.700 110.400 754.500 117.300 ;
        RECT 764.850 113.400 766.650 117.300 ;
        RECT 773.850 113.400 775.650 117.300 ;
        RECT 780.750 113.400 782.550 117.300 ;
        RECT 790.050 113.400 791.850 117.300 ;
        RECT 806.700 110.400 808.500 117.300 ;
        RECT 830.400 113.400 832.200 117.300 ;
        RECT 838.200 110.400 840.000 117.300 ;
        RECT 853.800 113.400 855.600 117.300 ;
        RECT 859.800 113.400 861.600 117.300 ;
        RECT 880.800 112.200 882.600 117.300 ;
        RECT 896.400 113.400 898.200 117.300 ;
        RECT 902.400 113.400 904.200 117.300 ;
        RECT 13.800 41.700 15.600 45.600 ;
        RECT 19.800 41.700 21.600 45.600 ;
        RECT 35.400 41.700 37.200 46.800 ;
        RECT 60.900 41.700 62.700 48.600 ;
        RECT 85.800 41.700 87.600 45.600 ;
        RECT 105.300 41.700 107.100 48.600 ;
        RECT 127.800 41.700 129.600 45.600 ;
        RECT 148.500 41.700 150.300 48.600 ;
        RECT 161.400 42.600 163.200 45.600 ;
        RECT 161.400 41.700 162.600 42.600 ;
        RECT 167.400 41.700 169.200 45.600 ;
        RECT 185.700 41.700 187.500 48.600 ;
        RECT 209.400 41.700 211.200 46.800 ;
        RECT 225.150 41.700 226.950 45.600 ;
        RECT 234.450 41.700 236.250 45.600 ;
        RECT 241.350 41.700 243.150 45.600 ;
        RECT 250.350 41.700 252.150 45.600 ;
        RECT 266.700 41.700 268.500 48.600 ;
        RECT 282.150 41.700 283.950 45.600 ;
        RECT 291.450 41.700 293.250 45.600 ;
        RECT 298.350 41.700 300.150 45.600 ;
        RECT 307.350 41.700 309.150 45.600 ;
        RECT 323.700 41.700 325.500 48.600 ;
        RECT 332.700 41.700 334.500 48.600 ;
        RECT 353.700 41.700 355.500 48.600 ;
        RECT 374.700 41.700 376.500 48.600 ;
        RECT 393.000 41.700 394.800 48.600 ;
        RECT 400.800 41.700 402.600 45.600 ;
        RECT 416.400 42.600 418.200 45.600 ;
        RECT 416.400 41.700 417.600 42.600 ;
        RECT 422.400 41.700 424.200 45.600 ;
        RECT 435.150 41.700 436.950 45.600 ;
        RECT 444.450 41.700 446.250 45.600 ;
        RECT 451.350 41.700 453.150 45.600 ;
        RECT 460.350 41.700 462.150 45.600 ;
        RECT 476.400 41.700 478.200 45.600 ;
        RECT 482.400 41.700 484.200 45.600 ;
        RECT 502.800 41.700 504.600 45.600 ;
        RECT 520.800 41.700 522.600 45.600 ;
        RECT 535.800 41.700 537.600 45.600 ;
        RECT 541.800 41.700 543.600 45.600 ;
        RECT 554.400 41.700 556.200 45.600 ;
        RECT 567.150 41.700 568.950 45.600 ;
        RECT 576.450 41.700 578.250 45.600 ;
        RECT 583.350 41.700 585.150 45.600 ;
        RECT 592.350 41.700 594.150 45.600 ;
        RECT 616.800 41.700 618.600 46.800 ;
        RECT 632.400 41.700 634.200 45.600 ;
        RECT 638.400 41.700 640.200 45.600 ;
        RECT 661.800 41.700 663.600 46.800 ;
        RECT 672.150 41.700 673.950 45.600 ;
        RECT 681.450 41.700 683.250 45.600 ;
        RECT 688.350 41.700 690.150 45.600 ;
        RECT 697.350 41.700 699.150 45.600 ;
        RECT 713.400 41.700 715.200 45.600 ;
        RECT 731.400 41.700 733.200 45.600 ;
        RECT 737.400 41.700 739.200 45.600 ;
        RECT 755.700 41.700 757.500 48.600 ;
        RECT 781.800 41.700 783.600 46.800 ;
        RECT 805.500 41.700 807.300 48.600 ;
        RECT 812.850 41.700 814.650 45.600 ;
        RECT 821.850 41.700 823.650 45.600 ;
        RECT 828.750 41.700 830.550 45.600 ;
        RECT 838.050 41.700 839.850 45.600 ;
        RECT 857.400 41.700 859.200 46.800 ;
        RECT 881.400 41.700 883.200 45.600 ;
        RECT 889.200 41.700 891.000 48.600 ;
        RECT 899.400 41.700 901.200 45.600 ;
        RECT 911.550 41.700 920.550 117.300 ;
        RECT 1.500 39.300 920.550 41.700 ;
        RECT 16.800 35.400 18.600 39.300 ;
        RECT 32.400 34.200 34.200 39.300 ;
        RECT 47.850 35.400 49.650 39.300 ;
        RECT 56.850 35.400 58.650 39.300 ;
        RECT 63.750 35.400 65.550 39.300 ;
        RECT 73.050 35.400 74.850 39.300 ;
        RECT 97.800 34.200 99.600 39.300 ;
        RECT 117.900 32.400 119.700 39.300 ;
        RECT 140.400 34.200 142.200 39.300 ;
        RECT 156.150 35.400 157.950 39.300 ;
        RECT 165.450 35.400 167.250 39.300 ;
        RECT 172.350 35.400 174.150 39.300 ;
        RECT 181.350 35.400 183.150 39.300 ;
        RECT 197.700 32.400 199.500 39.300 ;
        RECT 221.400 34.200 223.200 39.300 ;
        RECT 237.150 35.400 238.950 39.300 ;
        RECT 246.450 35.400 248.250 39.300 ;
        RECT 253.350 35.400 255.150 39.300 ;
        RECT 262.350 35.400 264.150 39.300 ;
        RECT 278.700 32.400 280.500 39.300 ;
        RECT 299.700 32.400 301.500 39.300 ;
        RECT 308.700 32.400 310.500 39.300 ;
        RECT 331.500 32.400 333.300 39.300 ;
        RECT 340.500 32.400 342.300 39.300 ;
        RECT 361.500 32.400 363.300 39.300 ;
        RECT 382.800 34.200 384.600 39.300 ;
        RECT 392.850 35.400 394.650 39.300 ;
        RECT 401.850 35.400 403.650 39.300 ;
        RECT 408.750 35.400 410.550 39.300 ;
        RECT 418.050 35.400 419.850 39.300 ;
        RECT 434.400 35.400 436.200 39.300 ;
        RECT 457.500 32.400 459.300 39.300 ;
        RECT 466.500 32.400 468.300 39.300 ;
        RECT 474.150 35.400 475.950 39.300 ;
        RECT 483.450 35.400 485.250 39.300 ;
        RECT 490.350 35.400 492.150 39.300 ;
        RECT 499.350 35.400 501.150 39.300 ;
        RECT 515.400 35.400 517.200 39.300 ;
        RECT 541.500 32.400 543.300 39.300 ;
        RECT 562.800 34.200 564.600 39.300 ;
        RECT 586.800 34.200 588.600 39.300 ;
        RECT 602.400 35.400 604.200 39.300 ;
        RECT 628.800 34.200 630.600 39.300 ;
        RECT 647.700 32.400 649.500 39.300 ;
        RECT 668.700 32.400 670.500 39.300 ;
        RECT 689.700 32.400 691.500 39.300 ;
        RECT 710.700 32.400 712.500 39.300 ;
        RECT 736.500 32.400 738.300 39.300 ;
        RECT 757.800 34.200 759.600 39.300 ;
        RECT 773.700 32.400 775.500 39.300 ;
        RECT 788.850 35.400 790.650 39.300 ;
        RECT 797.850 35.400 799.650 39.300 ;
        RECT 804.750 35.400 806.550 39.300 ;
        RECT 814.050 35.400 815.850 39.300 ;
        RECT 824.850 35.400 826.650 39.300 ;
        RECT 833.850 35.400 835.650 39.300 ;
        RECT 840.750 35.400 842.550 39.300 ;
        RECT 850.050 35.400 851.850 39.300 ;
        RECT 866.400 35.400 868.200 39.300 ;
        RECT 884.700 32.400 886.500 39.300 ;
        RECT 893.700 32.400 895.500 39.300 ;
        RECT 911.550 0.300 920.550 39.300 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -8.550 860.700 0.450 899.700 ;
        RECT 16.800 860.700 18.600 867.000 ;
        RECT 22.800 860.700 24.600 867.600 ;
        RECT 38.400 860.700 40.200 871.800 ;
        RECT 64.800 860.700 66.600 867.000 ;
        RECT 70.800 860.700 72.600 867.600 ;
        RECT 88.800 860.700 90.600 867.000 ;
        RECT 94.800 860.700 96.600 867.600 ;
        RECT 110.400 860.700 112.200 867.600 ;
        RECT 118.500 860.700 120.300 873.600 ;
        RECT 134.400 860.700 136.200 867.600 ;
        RECT 142.500 860.700 144.300 873.600 ;
        RECT 155.400 860.700 157.200 867.600 ;
        RECT 173.400 860.700 175.200 867.600 ;
        RECT 194.400 860.700 196.200 871.800 ;
        RECT 217.800 860.700 219.600 867.600 ;
        RECT 223.800 860.700 225.600 867.600 ;
        RECT 236.700 860.700 238.500 873.600 ;
        RECT 244.800 860.700 246.600 867.600 ;
        RECT 260.400 860.700 262.200 867.600 ;
        RECT 266.400 860.700 268.200 867.600 ;
        RECT 286.500 860.700 288.300 873.600 ;
        RECT 305.700 860.700 307.500 873.600 ;
        RECT 325.800 860.700 327.600 867.600 ;
        RECT 331.800 860.700 333.600 867.600 ;
        RECT 344.400 860.700 346.200 867.600 ;
        RECT 350.700 860.700 352.500 873.600 ;
        RECT 370.800 860.700 372.600 867.600 ;
        RECT 376.800 860.700 378.600 867.600 ;
        RECT 389.400 860.700 391.200 867.600 ;
        RECT 395.400 860.700 397.200 867.600 ;
        RECT 418.800 860.700 420.600 873.600 ;
        RECT 431.400 860.700 433.200 867.600 ;
        RECT 437.400 860.700 439.200 867.600 ;
        RECT 455.700 860.700 457.500 873.600 ;
        RECT 478.500 860.700 480.300 873.600 ;
        RECT 484.800 860.700 486.600 867.600 ;
        RECT 505.800 860.700 507.600 871.800 ;
        RECT 526.800 860.700 528.600 867.000 ;
        RECT 532.800 860.700 534.600 867.600 ;
        RECT 545.400 860.700 547.200 867.600 ;
        RECT 551.400 860.700 553.200 867.600 ;
        RECT 571.800 860.700 573.600 867.000 ;
        RECT 577.800 860.700 579.600 867.600 ;
        RECT 592.800 860.700 594.600 867.600 ;
        RECT 598.800 860.700 600.600 867.600 ;
        RECT 614.700 860.700 616.500 873.600 ;
        RECT 643.800 860.700 645.600 871.500 ;
        RECT 664.500 860.700 666.300 873.600 ;
        RECT 685.800 860.700 687.600 867.600 ;
        RECT 701.700 860.700 703.500 873.600 ;
        RECT 724.500 860.700 726.300 873.600 ;
        RECT 730.800 860.700 732.600 867.600 ;
        RECT 746.400 860.700 748.200 871.500 ;
        RECT 770.400 860.700 772.200 867.600 ;
        RECT 776.700 860.700 778.500 873.600 ;
        RECT 805.800 860.700 807.600 871.500 ;
        RECT 821.400 860.700 823.200 867.600 ;
        RECT 827.400 860.700 829.200 867.600 ;
        RECT 842.700 860.700 844.500 873.600 ;
        RECT 850.800 860.700 852.600 867.600 ;
        RECT 866.400 860.700 868.200 867.600 ;
        RECT 888.900 860.700 890.700 873.600 ;
        RECT -8.550 858.300 910.500 860.700 ;
        RECT -8.550 782.700 0.450 858.300 ;
        RECT 16.800 852.000 18.600 858.300 ;
        RECT 22.800 851.400 24.600 858.300 ;
        RECT 38.400 847.200 40.200 858.300 ;
        RECT 64.800 852.000 66.600 858.300 ;
        RECT 70.800 851.400 72.600 858.300 ;
        RECT 86.400 847.200 88.200 858.300 ;
        RECT 115.800 847.200 117.600 858.300 ;
        RECT 136.800 851.400 138.600 858.300 ;
        RECT 149.700 845.400 151.500 858.300 ;
        RECT 157.800 851.400 159.600 858.300 ;
        RECT 176.400 851.400 178.200 858.300 ;
        RECT 184.500 845.400 186.300 858.300 ;
        RECT 197.400 845.400 199.200 858.300 ;
        RECT 218.400 845.400 220.200 858.300 ;
        RECT 239.400 851.400 241.200 858.300 ;
        RECT 245.400 851.400 247.200 858.300 ;
        RECT 263.400 847.500 265.200 858.300 ;
        RECT 292.500 845.400 294.300 858.300 ;
        RECT 298.800 851.400 300.600 858.300 ;
        RECT 322.800 847.500 324.600 858.300 ;
        RECT 343.500 845.400 345.300 858.300 ;
        RECT 367.800 847.200 369.600 858.300 ;
        RECT 388.800 852.000 390.600 858.300 ;
        RECT 394.800 851.400 396.600 858.300 ;
        RECT 407.400 851.400 409.200 858.300 ;
        RECT 413.400 851.400 415.200 858.300 ;
        RECT 431.400 851.400 433.200 858.300 ;
        RECT 439.500 845.400 441.300 858.300 ;
        RECT 455.400 847.500 457.200 858.300 ;
        RECT 479.400 851.400 481.200 858.300 ;
        RECT 497.400 851.400 499.200 858.300 ;
        RECT 503.400 851.400 505.200 858.300 ;
        RECT 526.800 847.200 528.600 858.300 ;
        RECT 547.800 851.400 549.600 858.300 ;
        RECT 560.400 851.400 562.200 858.300 ;
        RECT 566.400 851.400 568.200 858.300 ;
        RECT 581.700 845.400 583.500 858.300 ;
        RECT 589.800 851.400 591.600 858.300 ;
        RECT 605.700 845.400 607.500 858.300 ;
        RECT 613.800 851.400 615.600 858.300 ;
        RECT 634.500 845.400 636.300 858.300 ;
        RECT 640.800 851.400 642.600 858.300 ;
        RECT 658.800 845.400 660.600 858.300 ;
        RECT 674.400 851.400 676.200 858.300 ;
        RECT 682.500 845.400 684.300 858.300 ;
        RECT 697.800 851.400 699.600 858.300 ;
        RECT 703.800 851.400 705.600 858.300 ;
        RECT 719.400 847.500 721.200 858.300 ;
        RECT 743.400 851.400 745.200 858.300 ;
        RECT 749.400 852.000 751.200 858.300 ;
        RECT 767.400 851.400 769.200 858.300 ;
        RECT 773.700 845.400 775.500 858.300 ;
        RECT 793.800 851.400 795.600 858.300 ;
        RECT 799.800 851.400 801.600 858.300 ;
        RECT 815.400 847.200 817.200 858.300 ;
        RECT 836.400 845.400 838.200 858.300 ;
        RECT 859.800 851.400 861.600 858.300 ;
        RECT 865.800 851.400 867.600 858.300 ;
        RECT 878.400 851.400 880.200 858.300 ;
        RECT 884.400 851.400 886.200 858.300 ;
        RECT 899.400 851.400 901.200 858.300 ;
        RECT 905.400 851.400 907.200 858.300 ;
        RECT 19.800 782.700 21.600 793.800 ;
        RECT 38.400 782.700 40.200 789.600 ;
        RECT 46.500 782.700 48.300 795.600 ;
        RECT 62.400 782.700 64.200 789.600 ;
        RECT 70.500 782.700 72.300 795.600 ;
        RECT 88.800 782.700 90.600 789.000 ;
        RECT 94.800 782.700 96.600 789.600 ;
        RECT 115.800 782.700 117.600 793.800 ;
        RECT 136.800 782.700 138.600 789.600 ;
        RECT 151.800 782.700 153.600 789.600 ;
        RECT 157.800 782.700 159.600 789.600 ;
        RECT 173.400 782.700 175.200 789.600 ;
        RECT 181.500 782.700 183.300 795.600 ;
        RECT 196.800 782.700 198.600 789.600 ;
        RECT 202.800 782.700 204.600 789.600 ;
        RECT 220.500 782.700 222.300 795.600 ;
        RECT 226.800 782.700 228.600 789.600 ;
        RECT 244.500 782.700 246.300 795.600 ;
        RECT 265.800 782.700 267.600 789.000 ;
        RECT 271.800 782.700 273.600 789.600 ;
        RECT 287.400 782.700 289.200 789.600 ;
        RECT 295.500 782.700 297.300 795.600 ;
        RECT 311.400 782.700 313.200 789.600 ;
        RECT 319.500 782.700 321.300 795.600 ;
        RECT 340.800 782.700 342.600 793.800 ;
        RECT 361.800 782.700 363.600 789.000 ;
        RECT 367.800 782.700 369.600 789.600 ;
        RECT 385.800 782.700 387.600 789.600 ;
        RECT 401.400 782.700 403.200 793.800 ;
        RECT 425.400 782.700 427.200 789.600 ;
        RECT 433.500 782.700 435.300 795.600 ;
        RECT 449.400 782.700 451.200 789.600 ;
        RECT 457.500 782.700 459.300 795.600 ;
        RECT 475.800 782.700 477.600 789.000 ;
        RECT 481.800 782.700 483.600 789.600 ;
        RECT 505.800 782.700 507.600 793.500 ;
        RECT 524.400 782.700 526.200 789.600 ;
        RECT 532.500 782.700 534.300 795.600 ;
        RECT 556.800 782.700 558.600 793.500 ;
        RECT 572.400 782.700 574.200 789.600 ;
        RECT 578.700 782.700 580.500 795.600 ;
        RECT 598.800 782.700 600.600 789.600 ;
        RECT 604.800 782.700 606.600 789.600 ;
        RECT 622.800 782.700 624.600 789.000 ;
        RECT 628.800 782.700 630.600 789.600 ;
        RECT 649.800 782.700 651.600 793.800 ;
        RECT 670.800 782.700 672.600 789.600 ;
        RECT 683.400 782.700 685.200 789.600 ;
        RECT 689.700 782.700 691.500 795.600 ;
        RECT 712.800 782.700 714.600 789.000 ;
        RECT 718.800 782.700 720.600 789.600 ;
        RECT 731.400 782.700 733.200 789.600 ;
        RECT 737.400 782.700 739.200 789.600 ;
        RECT 760.800 782.700 762.600 793.800 ;
        RECT 778.800 782.700 780.600 789.600 ;
        RECT 784.800 782.700 786.600 789.600 ;
        RECT 802.800 782.700 804.600 789.600 ;
        RECT 815.700 782.700 817.500 795.600 ;
        RECT 823.800 782.700 825.600 789.600 ;
        RECT 839.700 782.700 841.500 795.600 ;
        RECT 847.800 782.700 849.600 789.600 ;
        RECT 871.800 782.700 873.600 795.600 ;
        RECT 887.400 782.700 889.200 793.800 ;
        RECT -8.550 780.300 910.500 782.700 ;
        RECT -8.550 704.700 0.450 780.300 ;
        RECT 16.800 773.400 18.600 780.300 ;
        RECT 29.400 773.400 31.200 780.300 ;
        RECT 35.400 774.000 37.200 780.300 ;
        RECT 56.400 773.400 58.200 780.300 ;
        RECT 64.500 767.400 66.300 780.300 ;
        RECT 82.800 774.000 84.600 780.300 ;
        RECT 88.800 773.400 90.600 780.300 ;
        RECT 106.800 774.000 108.600 780.300 ;
        RECT 112.800 773.400 114.600 780.300 ;
        RECT 128.400 769.200 130.200 780.300 ;
        RECT 154.800 774.000 156.600 780.300 ;
        RECT 160.800 773.400 162.600 780.300 ;
        RECT 181.800 769.200 183.600 780.300 ;
        RECT 197.400 773.400 199.200 780.300 ;
        RECT 203.400 773.400 205.200 780.300 ;
        RECT 221.400 773.400 223.200 780.300 ;
        RECT 229.500 767.400 231.300 780.300 ;
        RECT 247.800 767.400 249.600 780.300 ;
        RECT 265.800 774.000 267.600 780.300 ;
        RECT 271.800 773.400 273.600 780.300 ;
        RECT 287.400 769.200 289.200 780.300 ;
        RECT 308.400 773.400 310.200 780.300 ;
        RECT 314.400 774.000 316.200 780.300 ;
        RECT 335.400 773.400 337.200 780.300 ;
        RECT 343.500 767.400 345.300 780.300 ;
        RECT 364.800 769.200 366.600 780.300 ;
        RECT 385.800 774.000 387.600 780.300 ;
        RECT 391.800 773.400 393.600 780.300 ;
        RECT 409.800 774.000 411.600 780.300 ;
        RECT 415.800 773.400 417.600 780.300 ;
        RECT 428.400 773.400 430.200 780.300 ;
        RECT 434.400 774.000 436.200 780.300 ;
        RECT 452.700 767.400 454.500 780.300 ;
        RECT 460.800 773.400 462.600 780.300 ;
        RECT 479.400 769.200 481.200 780.300 ;
        RECT 503.400 773.400 505.200 780.300 ;
        RECT 511.500 767.400 513.300 780.300 ;
        RECT 529.800 767.400 531.600 780.300 ;
        RECT 547.800 774.000 549.600 780.300 ;
        RECT 553.800 773.400 555.600 780.300 ;
        RECT 569.400 769.200 571.200 780.300 ;
        RECT 593.400 773.400 595.200 780.300 ;
        RECT 601.500 767.400 603.300 780.300 ;
        RECT 616.800 773.400 618.600 780.300 ;
        RECT 622.800 773.400 624.600 780.300 ;
        RECT 638.400 773.400 640.200 780.300 ;
        RECT 646.500 767.400 648.300 780.300 ;
        RECT 659.400 767.400 661.200 780.300 ;
        RECT 680.400 767.400 682.200 780.300 ;
        RECT 690.900 767.400 692.700 780.300 ;
        RECT 712.800 773.400 714.600 780.300 ;
        RECT 728.400 769.200 730.200 780.300 ;
        RECT 754.800 767.400 756.600 780.300 ;
        RECT 767.400 773.400 769.200 780.300 ;
        RECT 773.400 773.400 775.200 780.300 ;
        RECT 788.700 767.400 790.500 780.300 ;
        RECT 796.800 773.400 798.600 780.300 ;
        RECT 814.800 773.400 816.600 780.300 ;
        RECT 820.800 773.400 822.600 780.300 ;
        RECT 836.700 767.400 838.500 780.300 ;
        RECT 854.700 767.400 856.500 780.300 ;
        RECT 862.800 773.400 864.600 780.300 ;
        RECT 881.700 767.400 883.500 780.300 ;
        RECT 899.400 767.400 901.200 780.300 ;
        RECT 16.800 704.700 18.600 711.600 ;
        RECT 29.700 704.700 31.500 717.600 ;
        RECT 37.800 704.700 39.600 711.600 ;
        RECT 56.400 704.700 58.200 715.800 ;
        RECT 82.800 704.700 84.600 711.600 ;
        RECT 98.400 704.700 100.200 711.600 ;
        RECT 106.500 704.700 108.300 717.600 ;
        RECT 119.700 704.700 121.500 717.600 ;
        RECT 127.800 704.700 129.600 711.600 ;
        RECT 143.700 704.700 145.500 717.600 ;
        RECT 151.800 704.700 153.600 711.600 ;
        RECT 170.400 704.700 172.200 715.800 ;
        RECT 191.400 704.700 193.200 717.600 ;
        RECT 212.400 704.700 214.200 711.600 ;
        RECT 230.400 704.700 232.200 711.600 ;
        RECT 236.400 704.700 238.200 711.600 ;
        RECT 254.400 704.700 256.200 711.600 ;
        RECT 262.500 704.700 264.300 717.600 ;
        RECT 275.400 704.700 277.200 711.600 ;
        RECT 281.400 704.700 283.200 711.600 ;
        RECT 299.400 704.700 301.200 711.600 ;
        RECT 307.500 704.700 309.300 717.600 ;
        RECT 320.400 704.700 322.200 711.600 ;
        RECT 326.400 704.700 328.200 711.600 ;
        RECT 341.400 704.700 343.200 711.600 ;
        RECT 347.400 704.700 349.200 711.600 ;
        RECT 362.400 704.700 364.200 711.600 ;
        RECT 368.700 704.700 370.500 717.600 ;
        RECT 386.400 704.700 388.200 711.600 ;
        RECT 392.400 704.700 394.200 711.000 ;
        RECT 413.400 704.700 415.200 715.800 ;
        RECT 434.400 704.700 436.200 711.600 ;
        RECT 452.400 704.700 454.200 717.600 ;
        RECT 470.700 704.700 472.500 717.600 ;
        RECT 478.800 704.700 480.600 711.600 ;
        RECT 494.400 704.700 496.200 711.600 ;
        RECT 500.400 704.700 502.200 711.600 ;
        RECT 515.700 704.700 517.500 717.600 ;
        RECT 523.800 704.700 525.600 711.600 ;
        RECT 544.500 704.700 546.300 717.600 ;
        RECT 550.800 704.700 552.600 711.600 ;
        RECT 568.500 704.700 570.300 717.600 ;
        RECT 574.800 704.700 576.600 711.600 ;
        RECT 590.400 704.700 592.200 711.600 ;
        RECT 598.500 704.700 600.300 717.600 ;
        RECT 611.700 704.700 613.500 717.600 ;
        RECT 619.800 704.700 621.600 711.600 ;
        RECT 637.800 704.700 639.600 711.600 ;
        RECT 643.800 704.700 645.600 711.600 ;
        RECT 659.400 704.700 661.200 711.600 ;
        RECT 667.500 704.700 669.300 717.600 ;
        RECT 682.800 704.700 684.600 711.600 ;
        RECT 688.800 704.700 690.600 711.600 ;
        RECT 701.700 704.700 703.500 717.600 ;
        RECT 709.800 704.700 711.600 711.600 ;
        RECT 725.400 704.700 727.200 717.600 ;
        RECT 746.700 704.700 748.500 717.600 ;
        RECT 754.800 704.700 756.600 711.600 ;
        RECT 770.400 704.700 772.200 711.600 ;
        RECT 776.400 704.700 778.200 711.600 ;
        RECT 791.400 704.700 793.200 711.600 ;
        RECT 797.400 704.700 799.200 711.600 ;
        RECT 817.800 704.700 819.600 717.600 ;
        RECT 830.400 704.700 832.200 711.600 ;
        RECT 851.700 704.700 853.500 717.600 ;
        RECT 869.400 704.700 871.200 711.600 ;
        RECT 875.400 704.700 877.200 711.600 ;
        RECT 890.400 704.700 892.200 711.600 ;
        RECT 896.400 704.700 898.200 711.000 ;
        RECT -8.550 702.300 910.500 704.700 ;
        RECT -8.550 626.700 0.450 702.300 ;
        RECT 16.800 695.400 18.600 702.300 ;
        RECT 34.800 696.000 36.600 702.300 ;
        RECT 40.800 695.400 42.600 702.300 ;
        RECT 58.800 696.000 60.600 702.300 ;
        RECT 64.800 695.400 66.600 702.300 ;
        RECT 82.800 695.400 84.600 702.300 ;
        RECT 100.800 696.000 102.600 702.300 ;
        RECT 106.800 695.400 108.600 702.300 ;
        RECT 119.700 689.400 121.500 702.300 ;
        RECT 127.800 695.400 129.600 702.300 ;
        RECT 146.400 691.500 148.200 702.300 ;
        RECT 172.800 695.400 174.600 702.300 ;
        RECT 178.800 695.400 180.600 702.300 ;
        RECT 194.400 695.400 196.200 702.300 ;
        RECT 202.500 689.400 204.300 702.300 ;
        RECT 215.700 689.400 217.500 702.300 ;
        RECT 223.800 695.400 225.600 702.300 ;
        RECT 239.400 695.400 241.200 702.300 ;
        RECT 245.400 695.400 247.200 702.300 ;
        RECT 265.800 695.400 267.600 702.300 ;
        RECT 278.400 695.400 280.200 702.300 ;
        RECT 284.400 696.000 286.200 702.300 ;
        RECT 302.400 695.400 304.200 702.300 ;
        RECT 308.400 696.000 310.200 702.300 ;
        RECT 326.700 689.400 328.500 702.300 ;
        RECT 334.800 695.400 336.600 702.300 ;
        RECT 350.400 695.400 352.200 702.300 ;
        RECT 356.400 695.400 358.200 702.300 ;
        RECT 371.400 695.400 373.200 702.300 ;
        RECT 377.400 695.400 379.200 702.300 ;
        RECT 392.700 689.400 394.500 702.300 ;
        RECT 400.800 695.400 402.600 702.300 ;
        RECT 421.800 695.400 423.600 702.300 ;
        RECT 434.400 695.400 436.200 702.300 ;
        RECT 440.400 695.400 442.200 702.300 ;
        RECT 455.400 695.400 457.200 702.300 ;
        RECT 461.400 696.000 463.200 702.300 ;
        RECT 484.800 689.400 486.600 702.300 ;
        RECT 502.800 689.400 504.600 702.300 ;
        RECT 520.800 689.400 522.600 702.300 ;
        RECT 538.800 696.000 540.600 702.300 ;
        RECT 544.800 695.400 546.600 702.300 ;
        RECT 557.400 695.400 559.200 702.300 ;
        RECT 563.400 696.000 565.200 702.300 ;
        RECT 584.400 691.200 586.200 702.300 ;
        RECT 605.400 689.400 607.200 702.300 ;
        RECT 623.400 695.400 625.200 702.300 ;
        RECT 629.400 695.400 631.200 702.300 ;
        RECT 644.700 689.400 646.500 702.300 ;
        RECT 652.800 695.400 654.600 702.300 ;
        RECT 668.400 695.400 670.200 702.300 ;
        RECT 674.400 695.400 676.200 702.300 ;
        RECT 697.800 689.400 699.600 702.300 ;
        RECT 710.700 689.400 712.500 702.300 ;
        RECT 718.800 695.400 720.600 702.300 ;
        RECT 736.800 695.400 738.600 702.300 ;
        RECT 742.800 695.400 744.600 702.300 ;
        RECT 758.400 695.400 760.200 702.300 ;
        RECT 766.500 689.400 768.300 702.300 ;
        RECT 779.400 695.400 781.200 702.300 ;
        RECT 785.400 696.000 787.200 702.300 ;
        RECT 803.400 695.400 805.200 702.300 ;
        RECT 809.400 695.400 811.200 702.300 ;
        RECT 827.400 691.200 829.200 702.300 ;
        RECT 851.400 695.400 853.200 702.300 ;
        RECT 859.500 689.400 861.300 702.300 ;
        RECT 872.700 689.400 874.500 702.300 ;
        RECT 880.800 695.400 882.600 702.300 ;
        RECT 896.400 695.400 898.200 702.300 ;
        RECT 16.800 626.700 18.600 633.000 ;
        RECT 22.800 626.700 24.600 633.600 ;
        RECT 38.400 626.700 40.200 637.800 ;
        RECT 64.800 626.700 66.600 633.600 ;
        RECT 85.800 626.700 87.600 639.600 ;
        RECT 106.800 626.700 108.600 637.800 ;
        RECT 122.400 626.700 124.200 633.600 ;
        RECT 128.400 626.700 130.200 633.000 ;
        RECT 141.150 626.700 142.950 633.600 ;
        RECT 151.350 626.700 153.150 633.600 ;
        RECT 157.950 626.700 159.750 633.600 ;
        RECT 166.650 626.700 168.450 630.600 ;
        RECT 182.400 626.700 184.200 639.600 ;
        RECT 203.400 626.700 205.200 633.600 ;
        RECT 209.400 626.700 211.200 633.600 ;
        RECT 229.800 626.700 231.600 633.600 ;
        RECT 245.400 626.700 247.200 633.600 ;
        RECT 253.500 626.700 255.300 639.600 ;
        RECT 266.400 626.700 268.200 633.600 ;
        RECT 272.700 626.700 274.500 639.600 ;
        RECT 292.800 626.700 294.600 633.600 ;
        RECT 298.800 626.700 300.600 633.600 ;
        RECT 314.400 626.700 316.200 633.600 ;
        RECT 322.500 626.700 324.300 639.600 ;
        RECT 335.700 626.700 337.500 639.600 ;
        RECT 343.800 626.700 345.600 633.600 ;
        RECT 362.400 626.700 364.200 633.600 ;
        RECT 370.500 626.700 372.300 639.600 ;
        RECT 378.150 626.700 379.950 633.600 ;
        RECT 388.350 626.700 390.150 633.600 ;
        RECT 394.950 626.700 396.750 633.600 ;
        RECT 403.650 626.700 405.450 630.600 ;
        RECT 419.400 626.700 421.200 633.600 ;
        RECT 425.400 626.700 427.200 633.000 ;
        RECT 448.500 626.700 450.300 639.600 ;
        RECT 454.800 626.700 456.600 633.600 ;
        RECT 467.400 626.700 469.200 633.600 ;
        RECT 473.400 626.700 475.200 633.600 ;
        RECT 493.800 626.700 495.600 633.600 ;
        RECT 509.400 626.700 511.200 633.600 ;
        RECT 517.500 626.700 519.300 639.600 ;
        RECT 525.150 626.700 526.950 633.600 ;
        RECT 535.350 626.700 537.150 633.600 ;
        RECT 541.950 626.700 543.750 633.600 ;
        RECT 550.650 626.700 552.450 630.600 ;
        RECT 566.400 626.700 568.200 633.600 ;
        RECT 572.700 626.700 574.500 639.600 ;
        RECT 593.400 626.700 595.200 633.600 ;
        RECT 601.500 626.700 603.300 639.600 ;
        RECT 619.800 626.700 621.600 633.000 ;
        RECT 625.800 626.700 627.600 633.600 ;
        RECT 638.400 626.700 640.200 633.600 ;
        RECT 656.700 626.700 658.500 639.600 ;
        RECT 664.800 626.700 666.600 633.600 ;
        RECT 680.400 626.700 682.200 633.600 ;
        RECT 686.700 626.700 688.500 639.600 ;
        RECT 704.400 626.700 706.200 639.600 ;
        RECT 725.700 626.700 727.500 639.600 ;
        RECT 733.800 626.700 735.600 633.600 ;
        RECT 749.700 626.700 751.500 639.600 ;
        RECT 757.800 626.700 759.600 633.600 ;
        RECT 776.400 626.700 778.200 633.600 ;
        RECT 784.500 626.700 786.300 639.600 ;
        RECT 797.400 626.700 799.200 633.600 ;
        RECT 803.400 626.700 805.200 633.600 ;
        RECT 820.800 626.700 822.600 633.600 ;
        RECT 826.800 626.700 828.600 633.600 ;
        RECT 843.900 626.700 845.700 639.600 ;
        RECT 868.800 626.700 870.600 633.000 ;
        RECT 874.800 626.700 876.600 633.600 ;
        RECT 887.400 626.700 889.200 633.600 ;
        RECT 893.400 626.700 895.200 633.000 ;
        RECT -8.550 624.300 910.500 626.700 ;
        RECT -8.550 548.700 0.450 624.300 ;
        RECT 13.800 617.400 15.600 624.300 ;
        RECT 19.800 617.400 21.600 624.300 ;
        RECT 37.800 618.000 39.600 624.300 ;
        RECT 43.800 617.400 45.600 624.300 ;
        RECT 58.800 617.400 60.600 624.300 ;
        RECT 64.800 617.400 66.600 624.300 ;
        RECT 80.400 617.400 82.200 624.300 ;
        RECT 88.500 611.400 90.300 624.300 ;
        RECT 95.550 620.400 97.350 624.300 ;
        RECT 104.250 617.400 106.050 624.300 ;
        RECT 110.850 617.400 112.650 624.300 ;
        RECT 121.050 617.400 122.850 624.300 ;
        RECT 140.400 617.400 142.200 624.300 ;
        RECT 148.500 611.400 150.300 624.300 ;
        RECT 156.150 617.400 157.950 624.300 ;
        RECT 166.350 617.400 168.150 624.300 ;
        RECT 172.950 617.400 174.750 624.300 ;
        RECT 181.650 620.400 183.450 624.300 ;
        RECT 200.400 617.400 202.200 624.300 ;
        RECT 208.500 611.400 210.300 624.300 ;
        RECT 221.400 617.400 223.200 624.300 ;
        RECT 227.400 617.400 229.200 624.300 ;
        RECT 242.400 617.400 244.200 624.300 ;
        RECT 248.400 617.400 250.200 624.300 ;
        RECT 263.400 617.400 265.200 624.300 ;
        RECT 269.400 617.400 271.200 624.300 ;
        RECT 284.400 617.400 286.200 624.300 ;
        RECT 290.700 611.400 292.500 624.300 ;
        RECT 313.800 618.000 315.600 624.300 ;
        RECT 319.800 617.400 321.600 624.300 ;
        RECT 335.400 617.400 337.200 624.300 ;
        RECT 343.500 611.400 345.300 624.300 ;
        RECT 356.700 611.400 358.500 624.300 ;
        RECT 364.800 617.400 366.600 624.300 ;
        RECT 385.800 618.000 387.600 624.300 ;
        RECT 391.800 617.400 393.600 624.300 ;
        RECT 412.800 613.200 414.600 624.300 ;
        RECT 423.150 617.400 424.950 624.300 ;
        RECT 433.350 617.400 435.150 624.300 ;
        RECT 439.950 617.400 441.750 624.300 ;
        RECT 448.650 620.400 450.450 624.300 ;
        RECT 467.400 613.200 469.200 624.300 ;
        RECT 491.400 617.400 493.200 624.300 ;
        RECT 499.500 611.400 501.300 624.300 ;
        RECT 507.150 617.400 508.950 624.300 ;
        RECT 517.350 617.400 519.150 624.300 ;
        RECT 523.950 617.400 525.750 624.300 ;
        RECT 532.650 620.400 534.450 624.300 ;
        RECT 556.800 613.200 558.600 624.300 ;
        RECT 577.800 618.000 579.600 624.300 ;
        RECT 583.800 617.400 585.600 624.300 ;
        RECT 599.400 617.400 601.200 624.300 ;
        RECT 607.500 611.400 609.300 624.300 ;
        RECT 622.800 617.400 624.600 624.300 ;
        RECT 628.800 617.400 630.600 624.300 ;
        RECT 646.800 618.000 648.600 624.300 ;
        RECT 652.800 617.400 654.600 624.300 ;
        RECT 665.400 617.400 667.200 624.300 ;
        RECT 671.400 617.400 673.200 624.300 ;
        RECT 689.400 617.400 691.200 624.300 ;
        RECT 697.500 611.400 699.300 624.300 ;
        RECT 710.700 611.400 712.500 624.300 ;
        RECT 718.800 617.400 720.600 624.300 ;
        RECT 734.400 617.400 736.200 624.300 ;
        RECT 740.400 617.400 742.200 624.300 ;
        RECT 755.400 617.400 757.200 624.300 ;
        RECT 761.400 617.400 763.200 624.300 ;
        RECT 776.700 611.400 778.500 624.300 ;
        RECT 784.800 617.400 786.600 624.300 ;
        RECT 800.700 611.400 802.500 624.300 ;
        RECT 808.800 617.400 810.600 624.300 ;
        RECT 824.700 611.400 826.500 624.300 ;
        RECT 832.800 617.400 834.600 624.300 ;
        RECT 848.400 617.400 850.200 624.300 ;
        RECT 854.400 617.400 856.200 624.300 ;
        RECT 877.800 613.200 879.600 624.300 ;
        RECT 893.400 617.400 895.200 624.300 ;
        RECT 899.400 618.000 901.200 624.300 ;
        RECT 13.800 548.700 15.600 555.600 ;
        RECT 19.800 548.700 21.600 555.600 ;
        RECT 32.400 548.700 34.200 555.600 ;
        RECT 38.400 548.700 40.200 555.000 ;
        RECT 58.800 548.700 60.600 555.600 ;
        RECT 64.800 548.700 66.600 555.600 ;
        RECT 79.800 548.700 81.600 555.600 ;
        RECT 85.800 548.700 87.600 555.600 ;
        RECT 106.800 548.700 108.600 559.800 ;
        RECT 127.800 548.700 129.600 555.000 ;
        RECT 133.800 548.700 135.600 555.600 ;
        RECT 146.400 548.700 148.200 555.600 ;
        RECT 152.400 548.700 154.200 555.600 ;
        RECT 172.800 548.700 174.600 555.600 ;
        RECT 185.400 548.700 187.200 555.600 ;
        RECT 208.800 548.700 210.600 555.000 ;
        RECT 214.800 548.700 216.600 555.600 ;
        RECT 232.800 548.700 234.600 555.000 ;
        RECT 238.800 548.700 240.600 555.600 ;
        RECT 251.400 548.700 253.200 555.600 ;
        RECT 257.400 548.700 259.200 555.600 ;
        RECT 280.800 548.700 282.600 559.800 ;
        RECT 301.800 548.700 303.600 555.000 ;
        RECT 307.800 548.700 309.600 555.600 ;
        RECT 325.800 548.700 327.600 555.600 ;
        RECT 346.800 548.700 348.600 559.800 ;
        RECT 367.800 548.700 369.600 555.000 ;
        RECT 373.800 548.700 375.600 555.600 ;
        RECT 388.800 548.700 390.600 555.600 ;
        RECT 394.800 548.700 396.600 555.600 ;
        RECT 407.400 548.700 409.200 555.600 ;
        RECT 413.400 548.700 415.200 555.600 ;
        RECT 431.400 548.700 433.200 555.600 ;
        RECT 439.500 548.700 441.300 561.600 ;
        RECT 454.800 548.700 456.600 555.600 ;
        RECT 460.800 548.700 462.600 555.600 ;
        RECT 476.400 548.700 478.200 555.600 ;
        RECT 484.500 548.700 486.300 561.600 ;
        RECT 497.700 548.700 499.500 561.600 ;
        RECT 505.800 548.700 507.600 555.600 ;
        RECT 529.800 548.700 531.600 559.800 ;
        RECT 550.800 548.700 552.600 555.000 ;
        RECT 556.800 548.700 558.600 555.600 ;
        RECT 574.800 548.700 576.600 555.600 ;
        RECT 590.400 548.700 592.200 559.800 ;
        RECT 616.500 548.700 618.300 561.600 ;
        RECT 622.800 548.700 624.600 555.600 ;
        RECT 635.400 548.700 637.200 555.600 ;
        RECT 641.400 548.700 643.200 555.600 ;
        RECT 659.400 548.700 661.200 555.600 ;
        RECT 667.500 548.700 669.300 561.600 ;
        RECT 685.800 548.700 687.600 555.000 ;
        RECT 691.800 548.700 693.600 555.600 ;
        RECT 712.800 548.700 714.600 559.800 ;
        RECT 728.400 548.700 730.200 555.600 ;
        RECT 734.400 548.700 736.200 555.000 ;
        RECT 752.400 548.700 754.200 561.600 ;
        RECT 773.400 548.700 775.200 555.600 ;
        RECT 796.800 548.700 798.600 555.000 ;
        RECT 802.800 548.700 804.600 555.600 ;
        RECT 815.400 548.700 817.200 555.600 ;
        RECT 821.400 548.700 823.200 555.000 ;
        RECT 844.800 548.700 846.600 555.600 ;
        RECT 860.400 548.700 862.200 555.600 ;
        RECT 868.500 548.700 870.300 561.600 ;
        RECT 881.400 548.700 883.200 555.600 ;
        RECT 902.700 548.700 904.500 561.600 ;
        RECT -8.550 546.300 910.500 548.700 ;
        RECT -8.550 470.700 0.450 546.300 ;
        RECT 16.800 539.400 18.600 546.300 ;
        RECT 32.400 535.200 34.200 546.300 ;
        RECT 58.800 539.400 60.600 546.300 ;
        RECT 71.400 539.400 73.200 546.300 ;
        RECT 77.400 540.000 79.200 546.300 ;
        RECT 95.700 533.400 97.500 546.300 ;
        RECT 103.800 539.400 105.600 546.300 ;
        RECT 122.700 533.400 124.500 546.300 ;
        RECT 135.150 539.400 136.950 546.300 ;
        RECT 145.350 539.400 147.150 546.300 ;
        RECT 151.950 539.400 153.750 546.300 ;
        RECT 160.650 542.400 162.450 546.300 ;
        RECT 176.700 533.400 178.500 546.300 ;
        RECT 184.800 539.400 186.600 546.300 ;
        RECT 202.800 539.400 204.600 546.300 ;
        RECT 208.800 539.400 210.600 546.300 ;
        RECT 224.400 539.400 226.200 546.300 ;
        RECT 232.500 533.400 234.300 546.300 ;
        RECT 248.400 539.400 250.200 546.300 ;
        RECT 256.500 533.400 258.300 546.300 ;
        RECT 277.800 535.200 279.600 546.300 ;
        RECT 298.800 540.000 300.600 546.300 ;
        RECT 304.800 539.400 306.600 546.300 ;
        RECT 317.400 539.400 319.200 546.300 ;
        RECT 323.400 540.000 325.200 546.300 ;
        RECT 341.700 533.400 343.500 546.300 ;
        RECT 349.800 539.400 351.600 546.300 ;
        RECT 368.400 535.500 370.200 546.300 ;
        RECT 397.500 533.400 399.300 546.300 ;
        RECT 418.800 540.000 420.600 546.300 ;
        RECT 424.800 539.400 426.600 546.300 ;
        RECT 442.800 540.000 444.600 546.300 ;
        RECT 448.800 539.400 450.600 546.300 ;
        RECT 466.800 540.000 468.600 546.300 ;
        RECT 472.800 539.400 474.600 546.300 ;
        RECT 490.800 540.000 492.600 546.300 ;
        RECT 496.800 539.400 498.600 546.300 ;
        RECT 512.400 535.200 514.200 546.300 ;
        RECT 536.400 539.400 538.200 546.300 ;
        RECT 544.500 533.400 546.300 546.300 ;
        RECT 565.800 535.200 567.600 546.300 ;
        RECT 581.400 539.400 583.200 546.300 ;
        RECT 587.400 540.000 589.200 546.300 ;
        RECT 605.400 539.400 607.200 546.300 ;
        RECT 631.800 535.200 633.600 546.300 ;
        RECT 652.800 540.000 654.600 546.300 ;
        RECT 658.800 539.400 660.600 546.300 ;
        RECT 676.800 540.000 678.600 546.300 ;
        RECT 682.800 539.400 684.600 546.300 ;
        RECT 695.700 533.400 697.500 546.300 ;
        RECT 703.800 539.400 705.600 546.300 ;
        RECT 719.400 539.400 721.200 546.300 ;
        RECT 725.400 539.400 727.200 546.300 ;
        RECT 751.800 535.500 753.600 546.300 ;
        RECT 772.800 540.000 774.600 546.300 ;
        RECT 778.800 539.400 780.600 546.300 ;
        RECT 796.800 539.400 798.600 546.300 ;
        RECT 809.400 539.400 811.200 546.300 ;
        RECT 815.400 540.000 817.200 546.300 ;
        RECT 838.800 539.400 840.600 546.300 ;
        RECT 856.800 540.000 858.600 546.300 ;
        RECT 862.800 539.400 864.600 546.300 ;
        RECT 878.400 535.200 880.200 546.300 ;
        RECT 899.400 539.400 901.200 546.300 ;
        RECT 19.800 470.700 21.600 481.800 ;
        RECT 35.400 470.700 37.200 477.600 ;
        RECT 41.400 470.700 43.200 477.000 ;
        RECT 59.400 470.700 61.200 477.600 ;
        RECT 79.800 470.700 81.600 477.600 ;
        RECT 85.800 470.700 87.600 477.600 ;
        RECT 109.800 470.700 111.600 481.500 ;
        RECT 122.400 470.700 124.200 477.600 ;
        RECT 128.400 470.700 130.200 477.600 ;
        RECT 147.900 470.700 149.700 483.600 ;
        RECT 169.800 470.700 171.600 483.600 ;
        RECT 175.800 470.700 177.600 483.600 ;
        RECT 181.800 470.700 183.600 483.600 ;
        RECT 187.800 470.700 189.600 483.600 ;
        RECT 193.800 470.700 195.600 483.600 ;
        RECT 211.800 470.700 213.600 477.600 ;
        RECT 219.150 470.700 220.950 477.600 ;
        RECT 229.350 470.700 231.150 477.600 ;
        RECT 235.950 470.700 237.750 477.600 ;
        RECT 244.650 470.700 246.450 474.600 ;
        RECT 260.400 470.700 262.200 477.600 ;
        RECT 283.800 470.700 285.600 477.600 ;
        RECT 290.550 470.700 292.350 474.600 ;
        RECT 299.250 470.700 301.050 477.600 ;
        RECT 305.850 470.700 307.650 477.600 ;
        RECT 316.050 470.700 317.850 477.600 ;
        RECT 337.500 470.700 339.300 483.600 ;
        RECT 343.800 470.700 345.600 477.600 ;
        RECT 356.400 470.700 358.200 477.600 ;
        RECT 362.400 470.700 364.200 477.000 ;
        RECT 388.800 470.700 390.600 483.600 ;
        RECT 409.800 470.700 411.600 481.800 ;
        RECT 425.400 470.700 427.200 477.600 ;
        RECT 431.400 470.700 433.200 477.000 ;
        RECT 454.800 470.700 456.600 477.600 ;
        RECT 467.400 470.700 469.200 477.600 ;
        RECT 473.400 470.700 475.200 477.000 ;
        RECT 496.800 470.700 498.600 477.000 ;
        RECT 502.800 470.700 504.600 477.600 ;
        RECT 520.800 470.700 522.600 477.000 ;
        RECT 526.800 470.700 528.600 477.600 ;
        RECT 539.400 470.700 541.200 477.600 ;
        RECT 557.700 470.700 559.500 483.600 ;
        RECT 565.800 470.700 567.600 477.600 ;
        RECT 586.800 470.700 588.600 477.600 ;
        RECT 599.400 470.700 601.200 477.600 ;
        RECT 605.400 470.700 607.200 477.000 ;
        RECT 625.800 470.700 627.600 477.600 ;
        RECT 631.800 470.700 633.600 477.600 ;
        RECT 652.800 470.700 654.600 483.600 ;
        RECT 667.800 470.700 669.600 477.600 ;
        RECT 673.800 470.700 675.600 477.600 ;
        RECT 686.700 470.700 688.500 483.600 ;
        RECT 694.800 470.700 696.600 477.600 ;
        RECT 715.800 470.700 717.600 477.000 ;
        RECT 721.800 470.700 723.600 477.600 ;
        RECT 734.400 470.700 736.200 483.600 ;
        RECT 763.800 470.700 765.600 481.800 ;
        RECT 781.800 470.700 783.600 477.600 ;
        RECT 787.800 470.700 789.600 477.600 ;
        RECT 800.400 470.700 802.200 477.600 ;
        RECT 806.700 470.700 808.500 483.600 ;
        RECT 829.800 470.700 831.600 477.000 ;
        RECT 835.800 470.700 837.600 477.600 ;
        RECT 850.800 470.700 852.600 477.600 ;
        RECT 856.800 470.700 858.600 477.600 ;
        RECT 874.800 470.700 876.600 477.000 ;
        RECT 880.800 470.700 882.600 477.600 ;
        RECT 893.400 470.700 895.200 477.600 ;
        RECT 899.400 470.700 901.200 477.600 ;
        RECT -8.550 468.300 910.500 470.700 ;
        RECT -8.550 392.700 0.450 468.300 ;
        RECT 15.300 455.400 17.100 468.300 ;
        RECT 25.800 455.400 27.600 468.300 ;
        RECT 38.400 461.400 40.200 468.300 ;
        RECT 44.400 461.400 46.200 468.300 ;
        RECT 61.800 461.400 63.600 468.300 ;
        RECT 67.800 461.400 69.600 468.300 ;
        RECT 82.800 461.400 84.600 468.300 ;
        RECT 88.800 461.400 90.600 468.300 ;
        RECT 104.400 461.400 106.200 468.300 ;
        RECT 112.500 455.400 114.300 468.300 ;
        RECT 133.800 455.400 135.600 468.300 ;
        RECT 146.400 461.400 148.200 468.300 ;
        RECT 164.700 455.400 166.500 468.300 ;
        RECT 172.800 461.400 174.600 468.300 ;
        RECT 193.800 462.000 195.600 468.300 ;
        RECT 199.800 461.400 201.600 468.300 ;
        RECT 215.400 461.400 217.200 468.300 ;
        RECT 223.500 455.400 225.300 468.300 ;
        RECT 241.500 455.400 243.300 468.300 ;
        RECT 257.400 455.400 259.200 468.300 ;
        RECT 267.900 455.400 269.700 468.300 ;
        RECT 284.400 455.400 286.200 468.300 ;
        RECT 307.800 461.400 309.600 468.300 ;
        RECT 313.800 461.400 315.600 468.300 ;
        RECT 326.700 455.400 328.500 468.300 ;
        RECT 334.800 461.400 336.600 468.300 ;
        RECT 353.400 461.400 355.200 468.300 ;
        RECT 361.500 455.400 363.300 468.300 ;
        RECT 374.400 461.400 376.200 468.300 ;
        RECT 392.700 455.400 394.500 468.300 ;
        RECT 400.800 461.400 402.600 468.300 ;
        RECT 421.800 457.200 423.600 468.300 ;
        RECT 437.400 461.400 439.200 468.300 ;
        RECT 443.400 462.000 445.200 468.300 ;
        RECT 463.800 461.400 465.600 468.300 ;
        RECT 469.800 461.400 471.600 468.300 ;
        RECT 482.400 461.400 484.200 468.300 ;
        RECT 488.400 461.400 490.200 468.300 ;
        RECT 503.400 461.400 505.200 468.300 ;
        RECT 509.400 461.400 511.200 468.300 ;
        RECT 527.400 457.200 529.200 468.300 ;
        RECT 550.800 461.400 552.600 468.300 ;
        RECT 556.800 461.400 558.600 468.300 ;
        RECT 569.700 455.400 571.500 468.300 ;
        RECT 577.800 461.400 579.600 468.300 ;
        RECT 593.700 455.400 595.500 468.300 ;
        RECT 601.800 461.400 603.600 468.300 ;
        RECT 617.400 461.400 619.200 468.300 ;
        RECT 643.800 457.200 645.600 468.300 ;
        RECT 659.400 461.400 661.200 468.300 ;
        RECT 665.400 462.000 667.200 468.300 ;
        RECT 688.500 455.400 690.300 468.300 ;
        RECT 704.400 461.400 706.200 468.300 ;
        RECT 727.800 462.000 729.600 468.300 ;
        RECT 733.800 461.400 735.600 468.300 ;
        RECT 746.400 461.400 748.200 468.300 ;
        RECT 752.400 461.400 754.200 468.300 ;
        RECT 770.400 461.400 772.200 468.300 ;
        RECT 778.500 455.400 780.300 468.300 ;
        RECT 791.400 461.400 793.200 468.300 ;
        RECT 814.800 462.000 816.600 468.300 ;
        RECT 820.800 461.400 822.600 468.300 ;
        RECT 833.400 461.400 835.200 468.300 ;
        RECT 851.400 461.400 853.200 468.300 ;
        RECT 857.400 461.400 859.200 468.300 ;
        RECT 876.900 455.400 878.700 468.300 ;
        RECT 896.400 461.400 898.200 468.300 ;
        RECT 902.400 461.400 904.200 468.300 ;
        RECT 6.150 392.700 7.950 399.600 ;
        RECT 16.350 392.700 18.150 399.600 ;
        RECT 22.950 392.700 24.750 399.600 ;
        RECT 31.650 392.700 33.450 396.600 ;
        RECT 51.300 392.700 53.100 405.600 ;
        RECT 61.800 392.700 63.600 405.600 ;
        RECT 69.150 392.700 70.950 399.600 ;
        RECT 79.350 392.700 81.150 399.600 ;
        RECT 85.950 392.700 87.750 399.600 ;
        RECT 94.650 392.700 96.450 396.600 ;
        RECT 115.800 392.700 117.600 399.600 ;
        RECT 136.800 392.700 138.600 405.600 ;
        RECT 143.550 392.700 145.350 396.600 ;
        RECT 152.250 392.700 154.050 399.600 ;
        RECT 158.850 392.700 160.650 399.600 ;
        RECT 169.050 392.700 170.850 399.600 ;
        RECT 179.550 392.700 181.350 396.600 ;
        RECT 188.250 392.700 190.050 399.600 ;
        RECT 194.850 392.700 196.650 399.600 ;
        RECT 205.050 392.700 206.850 399.600 ;
        RECT 216.150 392.700 217.950 399.600 ;
        RECT 226.350 392.700 228.150 399.600 ;
        RECT 232.950 392.700 234.750 399.600 ;
        RECT 241.650 392.700 243.450 396.600 ;
        RECT 257.400 392.700 259.200 399.600 ;
        RECT 275.400 392.700 277.200 405.600 ;
        RECT 304.800 392.700 306.600 405.600 ;
        RECT 317.400 392.700 319.200 399.600 ;
        RECT 338.700 392.700 340.500 405.600 ;
        RECT 358.800 392.700 360.600 399.600 ;
        RECT 364.800 392.700 366.600 399.600 ;
        RECT 377.400 392.700 379.200 399.600 ;
        RECT 383.400 392.700 385.200 399.600 ;
        RECT 406.800 392.700 408.600 405.600 ;
        RECT 419.700 392.700 421.500 405.600 ;
        RECT 427.800 392.700 429.600 399.600 ;
        RECT 446.700 392.700 448.500 405.600 ;
        RECT 469.500 392.700 471.300 405.600 ;
        RECT 485.700 392.700 487.500 405.600 ;
        RECT 493.800 392.700 495.600 399.600 ;
        RECT 514.800 392.700 516.600 399.000 ;
        RECT 520.800 392.700 522.600 399.600 ;
        RECT 538.800 392.700 540.600 399.000 ;
        RECT 544.800 392.700 546.600 399.600 ;
        RECT 559.800 392.700 561.600 399.600 ;
        RECT 565.800 392.700 567.600 399.600 ;
        RECT 583.800 392.700 585.600 399.000 ;
        RECT 589.800 392.700 591.600 399.600 ;
        RECT 604.800 392.700 606.600 399.600 ;
        RECT 622.800 392.700 624.600 399.600 ;
        RECT 635.700 392.700 637.500 405.600 ;
        RECT 643.800 392.700 645.600 399.600 ;
        RECT 659.400 392.700 661.200 399.600 ;
        RECT 682.800 392.700 684.600 399.600 ;
        RECT 703.800 392.700 705.600 405.600 ;
        RECT 716.700 392.700 718.500 405.600 ;
        RECT 724.800 392.700 726.600 399.600 ;
        RECT 745.800 392.700 747.600 399.600 ;
        RECT 766.800 392.700 768.600 405.600 ;
        RECT 787.800 392.700 789.600 405.600 ;
        RECT 800.700 392.700 802.500 405.600 ;
        RECT 808.800 392.700 810.600 399.600 ;
        RECT 824.400 392.700 826.200 405.600 ;
        RECT 845.400 392.700 847.200 405.600 ;
        RECT 871.500 392.700 873.300 405.600 ;
        RECT 877.800 392.700 879.600 399.600 ;
        RECT 890.400 392.700 892.200 405.600 ;
        RECT -8.550 390.300 910.500 392.700 ;
        RECT -8.550 314.700 0.450 390.300 ;
        RECT 5.550 386.400 7.350 390.300 ;
        RECT 14.250 383.400 16.050 390.300 ;
        RECT 20.850 383.400 22.650 390.300 ;
        RECT 31.050 383.400 32.850 390.300 ;
        RECT 42.150 383.400 43.950 390.300 ;
        RECT 52.350 383.400 54.150 390.300 ;
        RECT 58.950 383.400 60.750 390.300 ;
        RECT 67.650 386.400 69.450 390.300 ;
        RECT 88.800 383.400 90.600 390.300 ;
        RECT 109.800 379.200 111.600 390.300 ;
        RECT 133.800 377.400 135.600 390.300 ;
        RECT 150.900 377.400 152.700 390.300 ;
        RECT 170.400 383.400 172.200 390.300 ;
        RECT 176.400 383.400 178.200 390.300 ;
        RECT 191.400 383.400 193.200 390.300 ;
        RECT 197.400 383.400 199.200 390.300 ;
        RECT 215.400 383.400 217.200 390.300 ;
        RECT 223.500 377.400 225.300 390.300 ;
        RECT 236.400 377.400 238.200 390.300 ;
        RECT 265.800 377.400 267.600 390.300 ;
        RECT 280.800 383.400 282.600 390.300 ;
        RECT 286.800 383.400 288.600 390.300 ;
        RECT 299.700 377.400 301.500 390.300 ;
        RECT 307.800 383.400 309.600 390.300 ;
        RECT 323.400 383.400 325.200 390.300 ;
        RECT 329.400 383.400 331.200 390.300 ;
        RECT 346.800 383.400 348.600 390.300 ;
        RECT 352.800 383.400 354.600 390.300 ;
        RECT 373.800 377.400 375.600 390.300 ;
        RECT 394.800 379.200 396.600 390.300 ;
        RECT 404.550 386.400 406.350 390.300 ;
        RECT 413.250 383.400 415.050 390.300 ;
        RECT 419.850 383.400 421.650 390.300 ;
        RECT 430.050 383.400 431.850 390.300 ;
        RECT 446.700 377.400 448.500 390.300 ;
        RECT 454.800 383.400 456.600 390.300 ;
        RECT 473.400 379.200 475.200 390.300 ;
        RECT 489.150 383.400 490.950 390.300 ;
        RECT 499.350 383.400 501.150 390.300 ;
        RECT 505.950 383.400 507.750 390.300 ;
        RECT 514.650 386.400 516.450 390.300 ;
        RECT 530.400 377.400 532.200 390.300 ;
        RECT 553.800 383.400 555.600 390.300 ;
        RECT 559.800 383.400 561.600 390.300 ;
        RECT 575.400 383.400 577.200 390.300 ;
        RECT 583.500 377.400 585.300 390.300 ;
        RECT 596.400 383.400 598.200 390.300 ;
        RECT 608.550 386.400 610.350 390.300 ;
        RECT 617.250 383.400 619.050 390.300 ;
        RECT 623.850 383.400 625.650 390.300 ;
        RECT 634.050 383.400 635.850 390.300 ;
        RECT 650.400 377.400 652.200 390.300 ;
        RECT 660.900 377.400 662.700 390.300 ;
        RECT 677.400 377.400 679.200 390.300 ;
        RECT 701.400 379.200 703.200 390.300 ;
        RECT 725.400 379.200 727.200 390.300 ;
        RECT 741.150 383.400 742.950 390.300 ;
        RECT 751.350 383.400 753.150 390.300 ;
        RECT 757.950 383.400 759.750 390.300 ;
        RECT 766.650 386.400 768.450 390.300 ;
        RECT 785.400 379.500 787.200 390.300 ;
        RECT 809.400 383.400 811.200 390.300 ;
        RECT 815.400 383.400 817.200 390.300 ;
        RECT 837.300 377.400 839.100 390.300 ;
        RECT 854.700 377.400 856.500 390.300 ;
        RECT 862.800 383.400 864.600 390.300 ;
        RECT 873.150 383.400 874.950 390.300 ;
        RECT 883.350 383.400 885.150 390.300 ;
        RECT 889.950 383.400 891.750 390.300 ;
        RECT 898.650 386.400 900.450 390.300 ;
        RECT 11.400 314.700 13.200 321.600 ;
        RECT 34.800 314.700 36.600 321.600 ;
        RECT 52.800 314.700 54.600 321.600 ;
        RECT 73.800 314.700 75.600 327.600 ;
        RECT 94.800 314.700 96.600 327.600 ;
        RECT 112.800 314.700 114.600 321.600 ;
        RECT 119.550 314.700 121.350 318.600 ;
        RECT 128.250 314.700 130.050 321.600 ;
        RECT 134.850 314.700 136.650 321.600 ;
        RECT 145.050 314.700 146.850 321.600 ;
        RECT 164.400 314.700 166.200 321.600 ;
        RECT 172.500 314.700 174.300 327.600 ;
        RECT 180.150 314.700 181.950 321.600 ;
        RECT 190.350 314.700 192.150 321.600 ;
        RECT 196.950 314.700 198.750 321.600 ;
        RECT 205.650 314.700 207.450 318.600 ;
        RECT 221.400 314.700 223.200 321.600 ;
        RECT 239.700 314.700 241.500 327.600 ;
        RECT 247.800 314.700 249.600 321.600 ;
        RECT 266.700 314.700 268.500 327.600 ;
        RECT 284.400 314.700 286.200 321.600 ;
        RECT 290.400 314.700 292.200 321.600 ;
        RECT 310.500 314.700 312.300 327.600 ;
        RECT 331.500 314.700 333.300 327.600 ;
        RECT 355.800 314.700 357.600 327.600 ;
        RECT 362.550 314.700 364.350 318.600 ;
        RECT 371.250 314.700 373.050 321.600 ;
        RECT 377.850 314.700 379.650 321.600 ;
        RECT 388.050 314.700 389.850 321.600 ;
        RECT 412.800 314.700 414.600 327.600 ;
        RECT 433.800 314.700 435.600 325.800 ;
        RECT 444.150 314.700 445.950 321.600 ;
        RECT 454.350 314.700 456.150 321.600 ;
        RECT 460.950 314.700 462.750 321.600 ;
        RECT 469.650 314.700 471.450 318.600 ;
        RECT 488.400 314.700 490.200 325.800 ;
        RECT 517.800 314.700 519.600 327.600 ;
        RECT 524.550 314.700 526.350 318.600 ;
        RECT 533.250 314.700 535.050 321.600 ;
        RECT 539.850 314.700 541.650 321.600 ;
        RECT 550.050 314.700 551.850 321.600 ;
        RECT 561.150 314.700 562.950 321.600 ;
        RECT 571.350 314.700 573.150 321.600 ;
        RECT 577.950 314.700 579.750 321.600 ;
        RECT 586.650 314.700 588.450 318.600 ;
        RECT 602.400 314.700 604.200 327.600 ;
        RECT 623.400 314.700 625.200 321.600 ;
        RECT 641.400 314.700 643.200 327.600 ;
        RECT 665.400 314.700 667.200 325.800 ;
        RECT 689.400 314.700 691.200 325.500 ;
        RECT 717.900 314.700 719.700 327.600 ;
        RECT 732.150 314.700 733.950 321.600 ;
        RECT 742.350 314.700 744.150 321.600 ;
        RECT 748.950 314.700 750.750 321.600 ;
        RECT 757.650 314.700 759.450 318.600 ;
        RECT 773.400 314.700 775.200 321.600 ;
        RECT 799.800 314.700 801.600 327.600 ;
        RECT 812.400 314.700 814.200 321.600 ;
        RECT 832.800 314.700 834.600 321.600 ;
        RECT 838.800 314.700 840.600 321.600 ;
        RECT 851.400 314.700 853.200 321.600 ;
        RECT 873.300 314.700 875.100 327.600 ;
        RECT 883.800 314.700 885.600 327.600 ;
        RECT 901.800 314.700 903.600 321.600 ;
        RECT -8.550 312.300 910.500 314.700 ;
        RECT -8.550 236.700 0.450 312.300 ;
        RECT 19.800 299.400 21.600 312.300 ;
        RECT 37.800 306.000 39.600 312.300 ;
        RECT 43.800 305.400 45.600 312.300 ;
        RECT 59.400 305.400 61.200 312.300 ;
        RECT 67.500 299.400 69.300 312.300 ;
        RECT 85.800 305.400 87.600 312.300 ;
        RECT 98.700 299.400 100.500 312.300 ;
        RECT 106.800 305.400 108.600 312.300 ;
        RECT 122.400 305.400 124.200 312.300 ;
        RECT 128.400 305.400 130.200 312.300 ;
        RECT 143.400 305.400 145.200 312.300 ;
        RECT 155.550 308.400 157.350 312.300 ;
        RECT 164.250 305.400 166.050 312.300 ;
        RECT 170.850 305.400 172.650 312.300 ;
        RECT 181.050 305.400 182.850 312.300 ;
        RECT 197.700 299.400 199.500 312.300 ;
        RECT 205.800 305.400 207.600 312.300 ;
        RECT 221.400 305.400 223.200 312.300 ;
        RECT 227.400 305.400 229.200 312.300 ;
        RECT 250.800 299.400 252.600 312.300 ;
        RECT 257.550 308.400 259.350 312.300 ;
        RECT 266.250 305.400 268.050 312.300 ;
        RECT 272.850 305.400 274.650 312.300 ;
        RECT 283.050 305.400 284.850 312.300 ;
        RECT 307.800 301.200 309.600 312.300 ;
        RECT 325.800 299.400 327.600 312.300 ;
        RECT 331.800 299.400 333.600 312.300 ;
        RECT 337.800 299.400 339.600 312.300 ;
        RECT 343.800 299.400 345.600 312.300 ;
        RECT 349.800 299.400 351.600 312.300 ;
        RECT 365.400 301.200 367.200 312.300 ;
        RECT 381.150 305.400 382.950 312.300 ;
        RECT 391.350 305.400 393.150 312.300 ;
        RECT 397.950 305.400 399.750 312.300 ;
        RECT 406.650 308.400 408.450 312.300 ;
        RECT 416.550 308.400 418.350 312.300 ;
        RECT 425.250 305.400 427.050 312.300 ;
        RECT 431.850 305.400 433.650 312.300 ;
        RECT 442.050 305.400 443.850 312.300 ;
        RECT 463.800 305.400 465.600 312.300 ;
        RECT 470.550 308.400 472.350 312.300 ;
        RECT 479.250 305.400 481.050 312.300 ;
        RECT 485.850 305.400 487.650 312.300 ;
        RECT 496.050 305.400 497.850 312.300 ;
        RECT 512.400 305.400 514.200 312.300 ;
        RECT 518.400 305.400 520.200 312.300 ;
        RECT 527.550 308.400 529.350 312.300 ;
        RECT 536.250 305.400 538.050 312.300 ;
        RECT 542.850 305.400 544.650 312.300 ;
        RECT 553.050 305.400 554.850 312.300 ;
        RECT 571.800 299.400 573.600 312.300 ;
        RECT 577.800 299.400 579.600 312.300 ;
        RECT 583.800 299.400 585.600 312.300 ;
        RECT 589.800 299.400 591.600 312.300 ;
        RECT 595.800 299.400 597.600 312.300 ;
        RECT 608.700 299.400 610.500 312.300 ;
        RECT 616.800 305.400 618.600 312.300 ;
        RECT 627.150 305.400 628.950 312.300 ;
        RECT 637.350 305.400 639.150 312.300 ;
        RECT 643.950 305.400 645.750 312.300 ;
        RECT 652.650 308.400 654.450 312.300 ;
        RECT 668.400 305.400 670.200 312.300 ;
        RECT 674.400 305.400 676.200 312.300 ;
        RECT 683.550 308.400 685.350 312.300 ;
        RECT 692.250 305.400 694.050 312.300 ;
        RECT 698.850 305.400 700.650 312.300 ;
        RECT 709.050 305.400 710.850 312.300 ;
        RECT 725.400 305.400 727.200 312.300 ;
        RECT 731.400 305.400 733.200 312.300 ;
        RECT 741.150 305.400 742.950 312.300 ;
        RECT 751.350 305.400 753.150 312.300 ;
        RECT 757.950 305.400 759.750 312.300 ;
        RECT 766.650 308.400 768.450 312.300 ;
        RECT 785.400 305.400 787.200 312.300 ;
        RECT 793.500 299.400 795.300 312.300 ;
        RECT 814.800 299.400 816.600 312.300 ;
        RECT 822.150 305.400 823.950 312.300 ;
        RECT 832.350 305.400 834.150 312.300 ;
        RECT 838.950 305.400 840.750 312.300 ;
        RECT 847.650 308.400 849.450 312.300 ;
        RECT 863.400 299.400 865.200 312.300 ;
        RECT 869.400 299.400 871.200 312.300 ;
        RECT 875.400 299.400 877.200 312.300 ;
        RECT 881.400 299.400 883.200 312.300 ;
        RECT 887.400 299.400 889.200 312.300 ;
        RECT 19.800 236.700 21.600 249.600 ;
        RECT 37.800 236.700 39.600 243.600 ;
        RECT 44.550 236.700 46.350 240.600 ;
        RECT 53.250 236.700 55.050 243.600 ;
        RECT 59.850 236.700 61.650 243.600 ;
        RECT 70.050 236.700 71.850 243.600 ;
        RECT 86.700 236.700 88.500 249.600 ;
        RECT 94.800 236.700 96.600 243.600 ;
        RECT 118.800 236.700 120.600 249.600 ;
        RECT 136.800 236.700 138.600 243.600 ;
        RECT 143.550 236.700 145.350 240.600 ;
        RECT 152.250 236.700 154.050 243.600 ;
        RECT 158.850 236.700 160.650 243.600 ;
        RECT 169.050 236.700 170.850 243.600 ;
        RECT 185.700 236.700 187.500 249.600 ;
        RECT 193.800 236.700 195.600 243.600 ;
        RECT 209.400 236.700 211.200 243.600 ;
        RECT 229.800 236.700 231.600 243.600 ;
        RECT 235.800 236.700 237.600 243.600 ;
        RECT 248.400 236.700 250.200 243.600 ;
        RECT 254.400 236.700 256.200 243.600 ;
        RECT 272.400 236.700 274.200 243.600 ;
        RECT 280.500 236.700 282.300 249.600 ;
        RECT 287.550 236.700 289.350 240.600 ;
        RECT 296.250 236.700 298.050 243.600 ;
        RECT 302.850 236.700 304.650 243.600 ;
        RECT 313.050 236.700 314.850 243.600 ;
        RECT 332.400 236.700 334.200 243.600 ;
        RECT 340.500 236.700 342.300 249.600 ;
        RECT 353.700 236.700 355.500 249.600 ;
        RECT 361.800 236.700 363.600 243.600 ;
        RECT 380.400 236.700 382.200 243.600 ;
        RECT 388.500 236.700 390.300 249.600 ;
        RECT 401.400 236.700 403.200 243.600 ;
        RECT 424.800 236.700 426.600 249.600 ;
        RECT 445.800 236.700 447.600 249.600 ;
        RECT 466.800 236.700 468.600 249.600 ;
        RECT 479.400 236.700 481.200 243.600 ;
        RECT 497.700 236.700 499.500 249.600 ;
        RECT 505.800 236.700 507.600 243.600 ;
        RECT 524.700 236.700 526.500 249.600 ;
        RECT 537.150 236.700 538.950 243.600 ;
        RECT 547.350 236.700 549.150 243.600 ;
        RECT 553.950 236.700 555.750 243.600 ;
        RECT 562.650 236.700 564.450 240.600 ;
        RECT 578.700 236.700 580.500 249.600 ;
        RECT 586.800 236.700 588.600 243.600 ;
        RECT 602.400 236.700 604.200 243.600 ;
        RECT 608.400 236.700 610.200 243.600 ;
        RECT 623.400 236.700 625.200 249.600 ;
        RECT 644.400 236.700 646.200 249.600 ;
        RECT 650.400 236.700 652.200 249.600 ;
        RECT 656.400 236.700 658.200 249.600 ;
        RECT 662.400 236.700 664.200 249.600 ;
        RECT 668.400 236.700 670.200 249.600 ;
        RECT 683.400 236.700 685.200 243.600 ;
        RECT 701.700 236.700 703.500 249.600 ;
        RECT 709.800 236.700 711.600 243.600 ;
        RECT 727.800 236.700 729.600 243.600 ;
        RECT 733.800 236.700 735.600 243.600 ;
        RECT 748.800 236.700 750.600 243.600 ;
        RECT 754.800 236.700 756.600 243.600 ;
        RECT 769.800 236.700 771.600 243.600 ;
        RECT 775.800 236.700 777.600 243.600 ;
        RECT 788.700 236.700 790.500 249.600 ;
        RECT 796.800 236.700 798.600 243.600 ;
        RECT 815.400 236.700 817.200 243.600 ;
        RECT 823.500 236.700 825.300 249.600 ;
        RECT 841.800 236.700 843.600 243.600 ;
        RECT 854.400 236.700 856.200 249.600 ;
        RECT 875.400 236.700 877.200 249.600 ;
        RECT 899.700 236.700 901.500 249.600 ;
        RECT -8.550 234.300 910.500 236.700 ;
        RECT -8.550 158.700 0.450 234.300 ;
        RECT 13.800 227.400 15.600 234.300 ;
        RECT 19.800 227.400 21.600 234.300 ;
        RECT 35.400 227.400 37.200 234.300 ;
        RECT 43.500 221.400 45.300 234.300 ;
        RECT 64.800 221.400 66.600 234.300 ;
        RECT 85.800 221.400 87.600 234.300 ;
        RECT 92.550 230.400 94.350 234.300 ;
        RECT 101.250 227.400 103.050 234.300 ;
        RECT 107.850 227.400 109.650 234.300 ;
        RECT 118.050 227.400 119.850 234.300 ;
        RECT 134.700 221.400 136.500 234.300 ;
        RECT 142.800 227.400 144.600 234.300 ;
        RECT 158.400 227.400 160.200 234.300 ;
        RECT 164.400 227.400 166.200 234.300 ;
        RECT 173.550 230.400 175.350 234.300 ;
        RECT 182.250 227.400 184.050 234.300 ;
        RECT 188.850 227.400 190.650 234.300 ;
        RECT 199.050 227.400 200.850 234.300 ;
        RECT 218.400 227.400 220.200 234.300 ;
        RECT 226.500 221.400 228.300 234.300 ;
        RECT 242.400 227.400 244.200 234.300 ;
        RECT 250.500 221.400 252.300 234.300 ;
        RECT 263.700 221.400 265.500 234.300 ;
        RECT 271.800 227.400 273.600 234.300 ;
        RECT 295.800 221.400 297.600 234.300 ;
        RECT 311.400 227.400 313.200 234.300 ;
        RECT 319.500 221.400 321.300 234.300 ;
        RECT 337.800 227.400 339.600 234.300 ;
        RECT 347.400 227.400 349.200 234.300 ;
        RECT 353.400 227.400 355.200 234.300 ;
        RECT 362.550 230.400 364.350 234.300 ;
        RECT 371.250 227.400 373.050 234.300 ;
        RECT 377.850 227.400 379.650 234.300 ;
        RECT 388.050 227.400 389.850 234.300 ;
        RECT 412.800 223.200 414.600 234.300 ;
        RECT 428.400 221.400 430.200 234.300 ;
        RECT 452.400 223.200 454.200 234.300 ;
        RECT 468.150 227.400 469.950 234.300 ;
        RECT 478.350 227.400 480.150 234.300 ;
        RECT 484.950 227.400 486.750 234.300 ;
        RECT 493.650 230.400 495.450 234.300 ;
        RECT 509.400 221.400 511.200 234.300 ;
        RECT 532.800 227.400 534.600 234.300 ;
        RECT 538.800 227.400 540.600 234.300 ;
        RECT 554.400 227.400 556.200 234.300 ;
        RECT 562.500 221.400 564.300 234.300 ;
        RECT 570.150 227.400 571.950 234.300 ;
        RECT 580.350 227.400 582.150 234.300 ;
        RECT 586.950 227.400 588.750 234.300 ;
        RECT 595.650 230.400 597.450 234.300 ;
        RECT 611.400 227.400 613.200 234.300 ;
        RECT 629.700 221.400 631.500 234.300 ;
        RECT 637.800 227.400 639.600 234.300 ;
        RECT 656.400 227.400 658.200 234.300 ;
        RECT 664.500 221.400 666.300 234.300 ;
        RECT 677.400 221.400 679.200 234.300 ;
        RECT 698.400 221.400 700.200 234.300 ;
        RECT 719.700 221.400 721.500 234.300 ;
        RECT 727.800 227.400 729.600 234.300 ;
        RECT 745.800 227.400 747.600 234.300 ;
        RECT 751.800 227.400 753.600 234.300 ;
        RECT 764.400 227.400 766.200 234.300 ;
        RECT 770.400 227.400 772.200 234.300 ;
        RECT 779.550 230.400 781.350 234.300 ;
        RECT 788.250 227.400 790.050 234.300 ;
        RECT 794.850 227.400 796.650 234.300 ;
        RECT 805.050 227.400 806.850 234.300 ;
        RECT 815.550 230.400 817.350 234.300 ;
        RECT 824.250 227.400 826.050 234.300 ;
        RECT 830.850 227.400 832.650 234.300 ;
        RECT 841.050 227.400 842.850 234.300 ;
        RECT 852.150 227.400 853.950 234.300 ;
        RECT 862.350 227.400 864.150 234.300 ;
        RECT 868.950 227.400 870.750 234.300 ;
        RECT 877.650 230.400 879.450 234.300 ;
        RECT 901.800 223.200 903.600 234.300 ;
        RECT 19.800 158.700 21.600 171.600 ;
        RECT 32.700 158.700 34.500 171.600 ;
        RECT 40.800 158.700 42.600 165.600 ;
        RECT 56.400 158.700 58.200 165.600 ;
        RECT 74.400 158.700 76.200 165.600 ;
        RECT 80.400 158.700 82.200 165.600 ;
        RECT 95.400 158.700 97.200 171.600 ;
        RECT 116.400 158.700 118.200 165.600 ;
        RECT 134.400 158.700 136.200 165.600 ;
        RECT 146.550 158.700 148.350 162.600 ;
        RECT 155.250 158.700 157.050 165.600 ;
        RECT 161.850 158.700 163.650 165.600 ;
        RECT 172.050 158.700 173.850 165.600 ;
        RECT 188.700 158.700 190.500 171.600 ;
        RECT 196.800 158.700 198.600 165.600 ;
        RECT 214.800 158.700 216.600 171.600 ;
        RECT 220.800 158.700 222.600 171.600 ;
        RECT 226.800 158.700 228.600 171.600 ;
        RECT 232.800 158.700 234.600 171.600 ;
        RECT 238.800 158.700 240.600 171.600 ;
        RECT 253.800 158.700 255.600 165.600 ;
        RECT 259.800 158.700 261.600 165.600 ;
        RECT 277.500 158.700 279.300 171.600 ;
        RECT 287.550 158.700 289.350 162.600 ;
        RECT 296.250 158.700 298.050 165.600 ;
        RECT 302.850 158.700 304.650 165.600 ;
        RECT 313.050 158.700 314.850 165.600 ;
        RECT 329.700 158.700 331.500 171.600 ;
        RECT 337.800 158.700 339.600 165.600 ;
        RECT 353.400 158.700 355.200 165.600 ;
        RECT 359.400 158.700 361.200 165.600 ;
        RECT 376.800 158.700 378.600 171.600 ;
        RECT 382.800 158.700 384.600 171.600 ;
        RECT 388.800 158.700 390.600 171.600 ;
        RECT 394.800 158.700 396.600 171.600 ;
        RECT 400.800 158.700 402.600 171.600 ;
        RECT 413.400 158.700 415.200 165.600 ;
        RECT 419.400 158.700 421.200 165.600 ;
        RECT 434.400 158.700 436.200 165.600 ;
        RECT 452.400 158.700 454.200 171.600 ;
        RECT 458.400 158.700 460.200 171.600 ;
        RECT 464.400 158.700 466.200 171.600 ;
        RECT 470.400 158.700 472.200 171.600 ;
        RECT 476.400 158.700 478.200 171.600 ;
        RECT 493.800 158.700 495.600 165.600 ;
        RECT 499.800 158.700 501.600 165.600 ;
        RECT 512.400 158.700 514.200 165.600 ;
        RECT 518.400 158.700 520.200 165.600 ;
        RECT 527.550 158.700 529.350 162.600 ;
        RECT 536.250 158.700 538.050 165.600 ;
        RECT 542.850 158.700 544.650 165.600 ;
        RECT 553.050 158.700 554.850 165.600 ;
        RECT 574.800 158.700 576.600 165.600 ;
        RECT 595.800 158.700 597.600 169.800 ;
        RECT 619.800 158.700 621.600 171.600 ;
        RECT 637.500 158.700 639.300 171.600 ;
        RECT 643.800 158.700 645.600 165.600 ;
        RECT 659.400 158.700 661.200 169.800 ;
        RECT 680.400 158.700 682.200 171.600 ;
        RECT 709.800 158.700 711.600 171.600 ;
        RECT 722.400 158.700 724.200 165.600 ;
        RECT 728.700 158.700 730.500 171.600 ;
        RECT 751.800 158.700 753.600 165.600 ;
        RECT 767.400 158.700 769.200 165.600 ;
        RECT 775.500 158.700 777.300 171.600 ;
        RECT 788.400 158.700 790.200 171.600 ;
        RECT 814.800 158.700 816.600 165.000 ;
        RECT 820.800 158.700 822.600 165.600 ;
        RECT 833.400 158.700 835.200 165.600 ;
        RECT 851.400 158.700 853.200 165.600 ;
        RECT 877.800 158.700 879.600 171.600 ;
        RECT 895.800 158.700 897.600 165.600 ;
        RECT -8.550 156.300 910.500 158.700 ;
        RECT -8.550 80.700 0.450 156.300 ;
        RECT 19.800 145.200 21.600 156.300 ;
        RECT 35.400 149.400 37.200 156.300 ;
        RECT 41.400 149.400 43.200 156.300 ;
        RECT 56.400 149.400 58.200 156.300 ;
        RECT 62.400 150.000 64.200 156.300 ;
        RECT 83.400 145.200 85.200 156.300 ;
        RECT 104.400 149.400 106.200 156.300 ;
        RECT 110.700 143.400 112.500 156.300 ;
        RECT 128.400 143.400 130.200 156.300 ;
        RECT 157.800 143.400 159.600 156.300 ;
        RECT 170.400 149.400 172.200 156.300 ;
        RECT 188.700 143.400 190.500 156.300 ;
        RECT 196.800 149.400 198.600 156.300 ;
        RECT 212.700 143.400 214.500 156.300 ;
        RECT 220.800 149.400 222.600 156.300 ;
        RECT 231.150 149.400 232.950 156.300 ;
        RECT 241.350 149.400 243.150 156.300 ;
        RECT 247.950 149.400 249.750 156.300 ;
        RECT 256.650 152.400 258.450 156.300 ;
        RECT 267.150 149.400 268.950 156.300 ;
        RECT 277.350 149.400 279.150 156.300 ;
        RECT 283.950 149.400 285.750 156.300 ;
        RECT 292.650 152.400 294.450 156.300 ;
        RECT 303.150 149.400 304.950 156.300 ;
        RECT 313.350 149.400 315.150 156.300 ;
        RECT 319.950 149.400 321.750 156.300 ;
        RECT 328.650 152.400 330.450 156.300 ;
        RECT 347.400 149.400 349.200 156.300 ;
        RECT 355.500 143.400 357.300 156.300 ;
        RECT 368.400 149.400 370.200 156.300 ;
        RECT 391.800 149.400 393.600 156.300 ;
        RECT 412.800 143.400 414.600 156.300 ;
        RECT 425.400 143.400 427.200 156.300 ;
        RECT 449.400 145.200 451.200 156.300 ;
        RECT 473.400 149.400 475.200 156.300 ;
        RECT 481.500 143.400 483.300 156.300 ;
        RECT 494.400 143.400 496.200 156.300 ;
        RECT 515.400 149.400 517.200 156.300 ;
        RECT 521.400 149.400 523.200 156.300 ;
        RECT 538.800 149.400 540.600 156.300 ;
        RECT 544.800 149.400 546.600 156.300 ;
        RECT 560.400 149.400 562.200 156.300 ;
        RECT 568.500 143.400 570.300 156.300 ;
        RECT 583.800 149.400 585.600 156.300 ;
        RECT 589.800 149.400 591.600 156.300 ;
        RECT 607.800 149.400 609.600 156.300 ;
        RECT 620.700 143.400 622.500 156.300 ;
        RECT 628.800 149.400 630.600 156.300 ;
        RECT 646.800 149.400 648.600 156.300 ;
        RECT 652.800 149.400 654.600 156.300 ;
        RECT 659.550 152.400 661.350 156.300 ;
        RECT 668.250 149.400 670.050 156.300 ;
        RECT 674.850 149.400 676.650 156.300 ;
        RECT 685.050 149.400 686.850 156.300 ;
        RECT 706.500 143.400 708.300 156.300 ;
        RECT 722.700 143.400 724.500 156.300 ;
        RECT 730.800 149.400 732.600 156.300 ;
        RECT 748.800 149.400 750.600 156.300 ;
        RECT 754.800 149.400 756.600 156.300 ;
        RECT 770.400 149.400 772.200 156.300 ;
        RECT 778.500 143.400 780.300 156.300 ;
        RECT 794.400 149.400 796.200 156.300 ;
        RECT 802.500 143.400 804.300 156.300 ;
        RECT 815.700 143.400 817.500 156.300 ;
        RECT 823.800 149.400 825.600 156.300 ;
        RECT 842.400 149.400 844.200 156.300 ;
        RECT 850.500 143.400 852.300 156.300 ;
        RECT 863.400 149.400 865.200 156.300 ;
        RECT 881.700 143.400 883.500 156.300 ;
        RECT 889.800 149.400 891.600 156.300 ;
        RECT 11.400 80.700 13.200 87.600 ;
        RECT 17.700 80.700 19.500 93.600 ;
        RECT 38.400 80.700 40.200 91.800 ;
        RECT 67.800 80.700 69.600 93.600 ;
        RECT 83.400 80.700 85.200 87.600 ;
        RECT 91.500 80.700 93.300 93.600 ;
        RECT 109.800 80.700 111.600 87.600 ;
        RECT 125.400 80.700 127.200 87.600 ;
        RECT 133.500 80.700 135.300 93.600 ;
        RECT 146.400 80.700 148.200 93.600 ;
        RECT 161.550 80.700 163.350 84.600 ;
        RECT 170.250 80.700 172.050 87.600 ;
        RECT 176.850 80.700 178.650 87.600 ;
        RECT 187.050 80.700 188.850 87.600 ;
        RECT 203.400 80.700 205.200 93.600 ;
        RECT 226.800 80.700 228.600 87.600 ;
        RECT 232.800 80.700 234.600 87.600 ;
        RECT 245.700 80.700 247.500 93.600 ;
        RECT 253.800 80.700 255.600 87.600 ;
        RECT 269.400 80.700 271.200 87.600 ;
        RECT 275.400 80.700 277.200 87.600 ;
        RECT 301.800 80.700 303.600 91.500 ;
        RECT 322.500 80.700 324.300 93.600 ;
        RECT 340.800 80.700 342.600 93.600 ;
        RECT 346.800 80.700 348.600 93.600 ;
        RECT 352.800 80.700 354.600 93.600 ;
        RECT 370.800 80.700 372.600 87.600 ;
        RECT 386.400 80.700 388.200 87.600 ;
        RECT 394.500 80.700 396.300 93.600 ;
        RECT 415.800 80.700 417.600 93.600 ;
        RECT 428.400 80.700 430.200 87.600 ;
        RECT 446.400 80.700 448.200 87.600 ;
        RECT 452.700 80.700 454.500 93.600 ;
        RECT 470.700 80.700 472.500 93.600 ;
        RECT 478.800 80.700 480.600 87.600 ;
        RECT 496.800 80.700 498.600 87.600 ;
        RECT 502.800 80.700 504.600 87.600 ;
        RECT 510.150 80.700 511.950 87.600 ;
        RECT 520.350 80.700 522.150 87.600 ;
        RECT 526.950 80.700 528.750 87.600 ;
        RECT 535.650 80.700 537.450 84.600 ;
        RECT 551.700 80.700 553.500 93.600 ;
        RECT 559.800 80.700 561.600 87.600 ;
        RECT 570.150 80.700 571.950 87.600 ;
        RECT 580.350 80.700 582.150 87.600 ;
        RECT 586.950 80.700 588.750 87.600 ;
        RECT 595.650 80.700 597.450 84.600 ;
        RECT 611.400 80.700 613.200 93.600 ;
        RECT 632.400 80.700 634.200 87.600 ;
        RECT 638.400 80.700 640.200 87.000 ;
        RECT 656.700 80.700 658.500 93.600 ;
        RECT 664.800 80.700 666.600 87.600 ;
        RECT 688.800 80.700 690.600 93.600 ;
        RECT 705.900 80.700 707.700 93.600 ;
        RECT 728.400 80.700 730.200 87.600 ;
        RECT 736.500 80.700 738.300 93.600 ;
        RECT 752.700 80.700 754.500 93.600 ;
        RECT 764.550 80.700 766.350 84.600 ;
        RECT 773.250 80.700 775.050 87.600 ;
        RECT 779.850 80.700 781.650 87.600 ;
        RECT 790.050 80.700 791.850 87.600 ;
        RECT 806.400 80.700 808.200 87.600 ;
        RECT 812.400 80.700 814.200 87.600 ;
        RECT 835.800 80.700 837.600 91.800 ;
        RECT 859.800 80.700 861.600 93.600 ;
        RECT 875.400 80.700 877.200 87.600 ;
        RECT 883.500 80.700 885.300 93.600 ;
        RECT 896.400 80.700 898.200 93.600 ;
        RECT -8.550 78.300 910.500 80.700 ;
        RECT -8.550 2.700 0.450 78.300 ;
        RECT 19.800 65.400 21.600 78.300 ;
        RECT 32.700 65.400 34.500 78.300 ;
        RECT 40.800 71.400 42.600 78.300 ;
        RECT 56.400 71.400 58.200 78.300 ;
        RECT 62.700 65.400 64.500 78.300 ;
        RECT 85.800 71.400 87.600 78.300 ;
        RECT 103.500 65.400 105.300 78.300 ;
        RECT 109.800 71.400 111.600 78.300 ;
        RECT 127.800 71.400 129.600 78.300 ;
        RECT 142.800 71.400 144.600 78.300 ;
        RECT 148.800 71.400 150.600 78.300 ;
        RECT 165.900 65.400 167.700 78.300 ;
        RECT 185.400 71.400 187.200 78.300 ;
        RECT 191.400 71.400 193.200 78.300 ;
        RECT 206.700 65.400 208.500 78.300 ;
        RECT 214.800 71.400 216.600 78.300 ;
        RECT 225.150 71.400 226.950 78.300 ;
        RECT 235.350 71.400 237.150 78.300 ;
        RECT 241.950 71.400 243.750 78.300 ;
        RECT 250.650 74.400 252.450 78.300 ;
        RECT 266.400 71.400 268.200 78.300 ;
        RECT 272.400 71.400 274.200 78.300 ;
        RECT 282.150 71.400 283.950 78.300 ;
        RECT 292.350 71.400 294.150 78.300 ;
        RECT 298.950 71.400 300.750 78.300 ;
        RECT 307.650 74.400 309.450 78.300 ;
        RECT 326.400 67.500 328.200 78.300 ;
        RECT 353.700 65.400 355.500 78.300 ;
        RECT 374.700 65.400 376.500 78.300 ;
        RECT 395.400 67.200 397.200 78.300 ;
        RECT 420.900 65.400 422.700 78.300 ;
        RECT 435.150 71.400 436.950 78.300 ;
        RECT 445.350 71.400 447.150 78.300 ;
        RECT 451.950 71.400 453.750 78.300 ;
        RECT 460.650 74.400 462.450 78.300 ;
        RECT 476.400 65.400 478.200 78.300 ;
        RECT 502.800 71.400 504.600 78.300 ;
        RECT 520.800 71.400 522.600 78.300 ;
        RECT 541.800 65.400 543.600 78.300 ;
        RECT 554.400 71.400 556.200 78.300 ;
        RECT 567.150 71.400 568.950 78.300 ;
        RECT 577.350 71.400 579.150 78.300 ;
        RECT 583.950 71.400 585.750 78.300 ;
        RECT 592.650 74.400 594.450 78.300 ;
        RECT 611.400 71.400 613.200 78.300 ;
        RECT 619.500 65.400 621.300 78.300 ;
        RECT 632.400 65.400 634.200 78.300 ;
        RECT 656.400 71.400 658.200 78.300 ;
        RECT 664.500 65.400 666.300 78.300 ;
        RECT 672.150 71.400 673.950 78.300 ;
        RECT 682.350 71.400 684.150 78.300 ;
        RECT 688.950 71.400 690.750 78.300 ;
        RECT 697.650 74.400 699.450 78.300 ;
        RECT 713.400 71.400 715.200 78.300 ;
        RECT 731.400 65.400 733.200 78.300 ;
        RECT 755.700 65.400 757.500 78.300 ;
        RECT 776.400 71.400 778.200 78.300 ;
        RECT 784.500 65.400 786.300 78.300 ;
        RECT 799.800 71.400 801.600 78.300 ;
        RECT 805.800 71.400 807.600 78.300 ;
        RECT 812.550 74.400 814.350 78.300 ;
        RECT 821.250 71.400 823.050 78.300 ;
        RECT 827.850 71.400 829.650 78.300 ;
        RECT 838.050 71.400 839.850 78.300 ;
        RECT 854.700 65.400 856.500 78.300 ;
        RECT 862.800 71.400 864.600 78.300 ;
        RECT 886.800 67.200 888.600 78.300 ;
        RECT 899.400 71.400 901.200 78.300 ;
        RECT 16.800 2.700 18.600 9.600 ;
        RECT 29.700 2.700 31.500 15.600 ;
        RECT 37.800 2.700 39.600 9.600 ;
        RECT 47.550 2.700 49.350 6.600 ;
        RECT 56.250 2.700 58.050 9.600 ;
        RECT 62.850 2.700 64.650 9.600 ;
        RECT 73.050 2.700 74.850 9.600 ;
        RECT 92.400 2.700 94.200 9.600 ;
        RECT 100.500 2.700 102.300 15.600 ;
        RECT 113.400 2.700 115.200 9.600 ;
        RECT 119.700 2.700 121.500 15.600 ;
        RECT 137.700 2.700 139.500 15.600 ;
        RECT 145.800 2.700 147.600 9.600 ;
        RECT 156.150 2.700 157.950 9.600 ;
        RECT 166.350 2.700 168.150 9.600 ;
        RECT 172.950 2.700 174.750 9.600 ;
        RECT 181.650 2.700 183.450 6.600 ;
        RECT 197.400 2.700 199.200 9.600 ;
        RECT 203.400 2.700 205.200 9.600 ;
        RECT 218.700 2.700 220.500 15.600 ;
        RECT 226.800 2.700 228.600 9.600 ;
        RECT 237.150 2.700 238.950 9.600 ;
        RECT 247.350 2.700 249.150 9.600 ;
        RECT 253.950 2.700 255.750 9.600 ;
        RECT 262.650 2.700 264.450 6.600 ;
        RECT 278.400 2.700 280.200 9.600 ;
        RECT 284.400 2.700 286.200 9.600 ;
        RECT 302.400 2.700 304.200 13.500 ;
        RECT 337.800 2.700 339.600 13.500 ;
        RECT 355.800 2.700 357.600 9.600 ;
        RECT 361.800 2.700 363.600 9.600 ;
        RECT 377.400 2.700 379.200 9.600 ;
        RECT 385.500 2.700 387.300 15.600 ;
        RECT 392.550 2.700 394.350 6.600 ;
        RECT 401.250 2.700 403.050 9.600 ;
        RECT 407.850 2.700 409.650 9.600 ;
        RECT 418.050 2.700 419.850 9.600 ;
        RECT 434.400 2.700 436.200 9.600 ;
        RECT 463.800 2.700 465.600 13.500 ;
        RECT 474.150 2.700 475.950 9.600 ;
        RECT 484.350 2.700 486.150 9.600 ;
        RECT 490.950 2.700 492.750 9.600 ;
        RECT 499.650 2.700 501.450 6.600 ;
        RECT 515.400 2.700 517.200 9.600 ;
        RECT 535.800 2.700 537.600 9.600 ;
        RECT 541.800 2.700 543.600 9.600 ;
        RECT 557.400 2.700 559.200 9.600 ;
        RECT 565.500 2.700 567.300 15.600 ;
        RECT 581.400 2.700 583.200 9.600 ;
        RECT 589.500 2.700 591.300 15.600 ;
        RECT 602.400 2.700 604.200 9.600 ;
        RECT 623.400 2.700 625.200 9.600 ;
        RECT 631.500 2.700 633.300 15.600 ;
        RECT 647.700 2.700 649.500 15.600 ;
        RECT 668.700 2.700 670.500 15.600 ;
        RECT 689.700 2.700 691.500 15.600 ;
        RECT 710.700 2.700 712.500 15.600 ;
        RECT 730.800 2.700 732.600 9.600 ;
        RECT 736.800 2.700 738.600 9.600 ;
        RECT 752.400 2.700 754.200 9.600 ;
        RECT 760.500 2.700 762.300 15.600 ;
        RECT 773.400 2.700 775.200 9.600 ;
        RECT 779.400 2.700 781.200 9.600 ;
        RECT 788.550 2.700 790.350 6.600 ;
        RECT 797.250 2.700 799.050 9.600 ;
        RECT 803.850 2.700 805.650 9.600 ;
        RECT 814.050 2.700 815.850 9.600 ;
        RECT 824.550 2.700 826.350 6.600 ;
        RECT 833.250 2.700 835.050 9.600 ;
        RECT 839.850 2.700 841.650 9.600 ;
        RECT 850.050 2.700 851.850 9.600 ;
        RECT 866.400 2.700 868.200 9.600 ;
        RECT 887.400 2.700 889.200 13.500 ;
        RECT -8.550 0.300 910.500 2.700 ;
    END
  END vdd
  PIN Cin[5]
    PORT
      LAYER metal1 ;
        RECT 814.950 892.950 817.050 895.050 ;
        RECT 815.550 865.050 816.450 892.950 ;
        RECT 814.950 862.950 817.050 865.050 ;
        RECT 784.950 850.950 787.050 853.050 ;
        RECT 785.550 826.050 786.450 850.950 ;
        RECT 784.950 823.950 787.050 826.050 ;
        RECT 490.950 712.950 493.050 715.050 ;
        RECT 491.550 709.050 492.450 712.950 ;
        RECT 490.950 706.950 493.050 709.050 ;
        RECT 382.950 697.950 385.050 700.050 ;
        RECT 383.550 673.050 384.450 697.950 ;
        RECT 382.950 670.950 385.050 673.050 ;
      LAYER metal2 ;
        RECT 814.950 894.450 817.050 895.050 ;
        RECT 820.950 894.450 823.050 895.050 ;
        RECT 814.950 893.400 823.050 894.450 ;
        RECT 814.950 892.950 817.050 893.400 ;
        RECT 820.950 892.950 823.050 893.400 ;
        RECT 791.100 864.450 793.200 865.050 ;
        RECT 814.950 864.450 817.050 865.050 ;
        RECT 791.100 863.400 817.050 864.450 ;
        RECT 791.100 862.950 793.200 863.400 ;
        RECT 814.950 862.950 817.050 863.400 ;
        RECT 784.950 852.450 787.050 853.050 ;
        RECT 790.950 852.450 793.050 853.050 ;
        RECT 784.950 851.400 793.050 852.450 ;
        RECT 784.950 850.950 787.050 851.400 ;
        RECT 790.950 850.950 793.050 851.400 ;
        RECT 742.950 822.450 745.050 823.050 ;
        RECT 784.950 822.450 787.050 826.050 ;
        RECT 742.950 822.000 787.050 822.450 ;
        RECT 742.950 821.400 786.450 822.000 ;
        RECT 742.950 820.950 745.050 821.400 ;
        RECT 742.950 765.450 745.050 766.050 ;
        RECT 754.950 765.450 757.050 766.050 ;
        RECT 742.950 764.400 757.050 765.450 ;
        RECT 742.950 763.950 745.050 764.400 ;
        RECT 754.950 763.950 757.050 764.400 ;
        RECT 718.950 747.450 721.050 748.050 ;
        RECT 754.950 747.450 757.050 748.050 ;
        RECT 760.950 747.450 763.050 748.050 ;
        RECT 718.950 746.400 763.050 747.450 ;
        RECT 718.950 745.950 721.050 746.400 ;
        RECT 754.950 745.950 757.050 746.400 ;
        RECT 760.950 745.950 763.050 746.400 ;
        RECT 676.950 741.450 679.050 742.050 ;
        RECT 718.800 741.450 720.900 742.200 ;
        RECT 676.950 740.400 720.900 741.450 ;
        RECT 676.950 739.950 679.050 740.400 ;
        RECT 718.800 740.100 720.900 740.400 ;
        RECT 490.950 714.450 493.050 715.050 ;
        RECT 470.400 713.400 493.050 714.450 ;
        RECT 454.950 711.450 457.050 712.050 ;
        RECT 470.400 711.450 471.450 713.400 ;
        RECT 490.950 712.950 493.050 713.400 ;
        RECT 454.950 710.400 471.450 711.450 ;
        RECT 454.950 709.950 457.050 710.400 ;
        RECT 490.950 708.450 493.050 709.050 ;
        RECT 490.950 707.400 519.450 708.450 ;
        RECT 490.950 706.950 493.050 707.400 ;
        RECT 518.400 705.450 519.450 707.400 ;
        RECT 628.950 705.450 631.050 706.050 ;
        RECT 676.950 705.450 679.050 706.050 ;
        RECT 518.400 704.400 540.450 705.450 ;
        RECT 539.400 702.450 540.450 704.400 ;
        RECT 584.400 704.400 679.050 705.450 ;
        RECT 584.400 702.450 585.450 704.400 ;
        RECT 628.950 703.950 631.050 704.400 ;
        RECT 676.950 703.950 679.050 704.400 ;
        RECT 539.400 701.400 585.450 702.450 ;
        RECT 382.950 699.450 385.050 700.050 ;
        RECT 439.950 699.450 442.050 700.050 ;
        RECT 454.950 699.450 457.050 700.050 ;
        RECT 382.950 698.400 457.050 699.450 ;
        RECT 382.950 697.950 385.050 698.400 ;
        RECT 439.950 697.950 442.050 698.400 ;
        RECT 454.950 697.950 457.050 698.400 ;
        RECT 760.950 696.450 763.050 697.050 ;
        RECT 808.950 696.450 811.050 697.050 ;
        RECT 760.950 695.400 811.050 696.450 ;
        RECT 760.950 694.950 763.050 695.400 ;
        RECT 808.950 694.950 811.050 695.400 ;
        RECT 376.950 685.950 379.050 688.050 ;
        RECT 439.950 685.950 442.050 691.050 ;
        RECT 628.950 685.950 631.050 688.050 ;
        RECT 808.950 685.950 811.050 688.050 ;
        RECT 376.950 672.450 379.050 673.050 ;
        RECT 382.950 672.450 385.050 673.050 ;
        RECT 376.950 671.400 385.050 672.450 ;
        RECT 376.950 670.950 379.050 671.400 ;
        RECT 382.950 670.950 385.050 671.400 ;
      LAYER metal3 ;
        RECT 821.400 895.050 822.600 906.600 ;
        RECT 820.950 892.950 823.050 895.050 ;
        RECT 791.100 862.950 793.200 865.050 ;
        RECT 791.400 853.050 792.600 862.950 ;
        RECT 790.950 850.950 793.050 853.050 ;
        RECT 742.950 820.950 745.050 823.050 ;
        RECT 743.400 766.050 744.600 820.950 ;
        RECT 742.950 763.950 745.050 766.050 ;
        RECT 754.950 763.950 757.050 766.050 ;
        RECT 755.400 748.050 756.600 763.950 ;
        RECT 718.950 745.950 721.050 748.050 ;
        RECT 754.950 745.950 757.050 748.050 ;
        RECT 760.950 745.950 763.050 748.050 ;
        RECT 719.400 742.200 720.600 745.950 ;
        RECT 676.950 739.950 679.050 742.050 ;
        RECT 718.800 740.100 720.900 742.200 ;
        RECT 454.950 709.950 457.050 712.050 ;
        RECT 455.400 700.050 456.600 709.950 ;
        RECT 677.400 706.050 678.600 739.950 ;
        RECT 628.950 703.950 631.050 706.050 ;
        RECT 676.950 703.950 679.050 706.050 ;
        RECT 439.950 697.950 442.050 700.050 ;
        RECT 454.950 697.950 457.050 700.050 ;
        RECT 440.400 691.050 441.600 697.950 ;
        RECT 439.950 688.950 442.050 691.050 ;
        RECT 629.400 688.050 630.600 703.950 ;
        RECT 761.400 697.050 762.600 745.950 ;
        RECT 760.950 694.950 763.050 697.050 ;
        RECT 808.950 694.950 811.050 697.050 ;
        RECT 809.400 688.050 810.600 694.950 ;
        RECT 376.950 685.950 379.050 688.050 ;
        RECT 628.950 685.950 631.050 688.050 ;
        RECT 808.950 685.950 811.050 688.050 ;
        RECT 377.400 673.050 378.600 685.950 ;
        RECT 376.950 670.950 379.050 673.050 ;
    END
  END Cin[5]
  PIN Cin[4]
    PORT
      LAYER metal1 ;
        RECT 736.950 889.950 739.050 892.050 ;
        RECT 737.550 868.050 738.450 889.950 ;
        RECT 787.950 883.950 790.050 886.050 ;
        RECT 736.950 865.950 739.050 868.050 ;
        RECT 788.550 865.050 789.450 883.950 ;
        RECT 787.800 862.950 789.900 865.050 ;
        RECT 733.950 829.950 736.050 832.050 ;
        RECT 734.550 826.050 735.450 829.950 ;
        RECT 733.800 823.950 735.900 826.050 ;
        RECT 379.950 733.950 382.050 736.050 ;
        RECT 380.550 715.050 381.450 733.950 ;
        RECT 784.950 724.950 787.050 727.050 ;
        RECT 785.550 715.050 786.450 724.950 ;
        RECT 379.950 712.950 382.050 715.050 ;
        RECT 785.100 712.950 787.200 715.050 ;
        RECT 796.950 697.950 799.050 700.050 ;
        RECT 598.950 691.950 601.050 694.050 ;
        RECT 599.550 670.050 600.450 691.950 ;
        RECT 797.550 670.050 798.450 697.950 ;
        RECT 599.100 667.950 601.200 670.050 ;
        RECT 796.950 667.950 799.050 670.050 ;
        RECT 260.100 658.950 262.200 661.050 ;
        RECT 260.550 631.050 261.450 658.950 ;
        RECT 769.950 652.950 772.050 655.050 ;
        RECT 770.550 631.050 771.450 652.950 ;
        RECT 259.950 628.950 262.050 631.050 ;
        RECT 769.950 628.950 772.050 631.050 ;
      LAYER metal2 ;
        RECT 742.950 897.450 745.050 898.050 ;
        RECT 781.950 897.450 784.050 898.050 ;
        RECT 742.950 896.400 784.050 897.450 ;
        RECT 742.950 895.950 745.050 896.400 ;
        RECT 781.950 895.950 784.050 896.400 ;
        RECT 736.950 891.450 739.050 892.050 ;
        RECT 742.950 891.450 745.050 892.050 ;
        RECT 736.950 890.400 745.050 891.450 ;
        RECT 736.950 889.950 739.050 890.400 ;
        RECT 742.950 889.950 745.050 890.400 ;
        RECT 745.950 886.950 748.050 889.050 ;
        RECT 781.950 885.450 784.050 886.050 ;
        RECT 787.950 885.450 790.050 886.050 ;
        RECT 781.950 884.400 790.050 885.450 ;
        RECT 781.950 883.950 784.050 884.400 ;
        RECT 787.950 883.950 790.050 884.400 ;
        RECT 815.100 873.000 817.200 874.050 ;
        RECT 814.950 871.950 817.200 873.000 ;
        RECT 814.950 871.050 817.050 871.950 ;
        RECT 811.950 870.000 817.050 871.050 ;
        RECT 811.950 869.400 816.600 870.000 ;
        RECT 811.950 868.950 816.000 869.400 ;
        RECT 713.100 867.450 715.200 868.050 ;
        RECT 736.950 867.450 739.050 868.050 ;
        RECT 713.100 866.400 739.050 867.450 ;
        RECT 713.100 865.950 715.200 866.400 ;
        RECT 736.950 865.950 739.050 866.400 ;
        RECT 787.800 864.000 789.900 865.050 ;
        RECT 787.800 862.950 790.050 864.000 ;
        RECT 787.950 861.450 790.050 862.950 ;
        RECT 811.950 861.450 814.050 862.050 ;
        RECT 787.950 861.000 814.050 861.450 ;
        RECT 788.400 860.400 814.050 861.000 ;
        RECT 811.950 859.950 814.050 860.400 ;
        RECT 745.950 832.950 748.050 835.050 ;
        RECT 733.950 831.450 736.050 832.050 ;
        RECT 742.950 831.450 745.050 832.050 ;
        RECT 733.950 830.400 745.050 831.450 ;
        RECT 733.950 829.950 736.050 830.400 ;
        RECT 742.950 829.950 745.050 830.400 ;
        RECT 712.950 825.450 715.050 826.050 ;
        RECT 724.950 825.450 727.050 826.050 ;
        RECT 733.800 825.450 735.900 826.050 ;
        RECT 712.950 824.400 735.900 825.450 ;
        RECT 712.950 823.950 715.050 824.400 ;
        RECT 724.950 823.950 727.050 824.400 ;
        RECT 733.800 823.950 735.900 824.400 ;
        RECT 724.950 780.450 727.050 781.050 ;
        RECT 769.950 780.450 772.050 781.050 ;
        RECT 724.950 779.400 772.050 780.450 ;
        RECT 724.950 778.950 727.050 779.400 ;
        RECT 769.950 778.950 772.050 779.400 ;
        RECT 769.950 747.450 772.050 748.050 ;
        RECT 778.950 747.450 781.050 748.050 ;
        RECT 769.950 746.400 781.050 747.450 ;
        RECT 769.950 745.950 772.050 746.400 ;
        RECT 778.950 745.950 781.050 746.400 ;
        RECT 442.950 744.450 445.050 745.050 ;
        RECT 514.950 744.450 517.050 745.050 ;
        RECT 562.950 744.450 565.050 745.050 ;
        RECT 568.950 744.450 571.050 745.050 ;
        RECT 442.950 743.400 571.050 744.450 ;
        RECT 442.950 742.950 445.050 743.400 ;
        RECT 514.950 742.950 517.050 743.400 ;
        RECT 562.950 742.950 565.050 743.400 ;
        RECT 568.950 742.950 571.050 743.400 ;
        RECT 379.950 735.450 382.050 736.050 ;
        RECT 442.950 735.450 445.050 736.050 ;
        RECT 379.950 734.400 445.050 735.450 ;
        RECT 379.950 733.950 382.050 734.400 ;
        RECT 442.950 733.950 445.050 734.400 ;
        RECT 568.950 727.950 571.050 730.050 ;
        RECT 778.950 726.450 781.050 727.050 ;
        RECT 784.950 726.450 787.050 727.050 ;
        RECT 778.950 725.400 787.050 726.450 ;
        RECT 778.950 724.950 781.050 725.400 ;
        RECT 784.950 724.950 787.050 725.400 ;
        RECT 325.950 718.950 328.050 721.050 ;
        RECT 775.950 718.950 778.050 721.050 ;
        RECT 275.100 714.450 277.200 715.050 ;
        RECT 325.950 714.450 328.050 715.050 ;
        RECT 346.950 714.450 349.050 715.050 ;
        RECT 379.950 714.450 382.050 715.050 ;
        RECT 275.100 713.400 382.050 714.450 ;
        RECT 275.100 712.950 277.200 713.400 ;
        RECT 325.950 712.950 328.050 713.400 ;
        RECT 346.950 712.950 349.050 713.400 ;
        RECT 379.950 712.950 382.050 713.400 ;
        RECT 785.100 714.450 787.200 715.050 ;
        RECT 805.950 714.450 808.050 715.050 ;
        RECT 785.100 713.400 808.050 714.450 ;
        RECT 785.100 712.950 787.200 713.400 ;
        RECT 805.950 712.950 808.050 713.400 ;
        RECT 502.950 705.450 505.050 706.050 ;
        RECT 514.950 705.450 517.050 706.050 ;
        RECT 502.950 704.400 517.050 705.450 ;
        RECT 502.950 703.950 505.050 704.400 ;
        RECT 514.950 703.950 517.050 704.400 ;
        RECT 347.100 699.450 349.200 700.050 ;
        RECT 361.950 699.450 364.050 699.900 ;
        RECT 347.100 698.400 364.050 699.450 ;
        RECT 347.100 697.950 349.200 698.400 ;
        RECT 361.950 697.800 364.050 698.400 ;
        RECT 796.950 699.450 799.050 700.050 ;
        RECT 805.950 699.450 808.050 700.050 ;
        RECT 796.950 698.400 808.050 699.450 ;
        RECT 796.950 697.950 799.050 698.400 ;
        RECT 805.950 697.950 808.050 698.400 ;
        RECT 562.950 693.450 565.050 694.050 ;
        RECT 598.950 693.450 601.050 694.050 ;
        RECT 562.950 692.400 601.050 693.450 ;
        RECT 562.950 691.950 565.050 692.400 ;
        RECT 598.950 691.950 601.050 692.400 ;
        RECT 355.950 687.450 358.050 688.050 ;
        RECT 360.000 687.450 364.050 688.050 ;
        RECT 355.950 686.400 364.050 687.450 ;
        RECT 355.950 685.950 358.050 686.400 ;
        RECT 360.000 685.950 364.050 686.400 ;
        RECT 502.950 685.950 505.050 688.050 ;
        RECT 599.100 669.000 601.200 670.050 ;
        RECT 598.950 667.950 601.200 669.000 ;
        RECT 776.100 669.450 778.200 670.050 ;
        RECT 796.950 669.450 799.050 670.050 ;
        RECT 808.950 669.450 811.050 670.050 ;
        RECT 776.100 668.400 811.050 669.450 ;
        RECT 776.100 667.950 778.200 668.400 ;
        RECT 796.950 667.950 799.050 668.400 ;
        RECT 808.950 667.950 811.050 668.400 ;
        RECT 571.950 666.450 574.050 667.050 ;
        RECT 598.950 666.450 601.050 667.950 ;
        RECT 571.950 666.000 601.050 666.450 ;
        RECT 571.950 665.400 600.450 666.000 ;
        RECT 571.950 664.950 574.050 665.400 ;
        RECT 260.100 660.450 262.200 661.050 ;
        RECT 274.950 660.450 277.050 661.050 ;
        RECT 260.100 659.400 277.050 660.450 ;
        RECT 260.100 658.950 262.200 659.400 ;
        RECT 274.950 658.950 277.050 659.400 ;
        RECT 769.950 654.900 774.000 655.050 ;
        RECT 769.950 652.950 775.050 654.900 ;
        RECT 772.950 652.800 775.050 652.950 ;
        RECT 571.950 649.950 574.050 652.050 ;
        RECT 820.950 640.950 823.050 643.050 ;
        RECT 808.950 639.450 811.050 640.200 ;
        RECT 808.950 638.400 816.450 639.450 ;
        RECT 808.950 638.100 811.050 638.400 ;
        RECT 815.400 636.450 816.450 638.400 ;
        RECT 820.950 636.450 823.050 637.050 ;
        RECT 815.400 635.400 823.050 636.450 ;
        RECT 820.950 634.950 823.050 635.400 ;
        RECT 571.950 633.450 574.050 634.050 ;
        RECT 685.950 633.450 688.050 634.050 ;
        RECT 571.950 632.400 688.050 633.450 ;
        RECT 571.950 631.950 574.050 632.400 ;
        RECT 685.950 631.950 688.050 632.400 ;
        RECT 259.950 630.450 262.050 631.050 ;
        RECT 289.950 630.450 292.050 631.050 ;
        RECT 259.950 629.400 292.050 630.450 ;
        RECT 259.950 628.950 262.050 629.400 ;
        RECT 289.950 628.950 292.050 629.400 ;
        RECT 760.950 630.450 763.050 631.050 ;
        RECT 769.950 630.450 772.050 631.050 ;
        RECT 760.950 629.400 772.050 630.450 ;
        RECT 760.950 628.950 763.050 629.400 ;
        RECT 769.950 628.950 772.050 629.400 ;
        RECT 685.950 615.450 688.050 616.050 ;
        RECT 760.950 615.450 763.050 616.050 ;
        RECT 685.950 614.400 763.050 615.450 ;
        RECT 685.950 613.950 688.050 614.400 ;
        RECT 760.950 613.950 763.050 614.400 ;
        RECT 760.950 607.950 763.050 610.050 ;
        RECT 289.950 598.950 292.050 601.050 ;
      LAYER metal3 ;
        RECT 812.400 905.400 816.600 906.600 ;
        RECT 742.950 895.950 745.050 898.050 ;
        RECT 781.950 895.950 784.050 898.050 ;
        RECT 743.400 892.050 744.600 895.950 ;
        RECT 742.950 889.050 745.050 892.050 ;
        RECT 742.950 888.000 748.050 889.050 ;
        RECT 743.400 887.400 748.050 888.000 ;
        RECT 744.000 886.950 748.050 887.400 ;
        RECT 782.400 886.050 783.600 895.950 ;
        RECT 812.400 894.600 813.600 905.400 ;
        RECT 812.400 893.400 816.600 894.600 ;
        RECT 781.950 883.950 784.050 886.050 ;
        RECT 815.400 874.050 816.600 893.400 ;
        RECT 815.100 871.950 817.200 874.050 ;
        RECT 811.950 868.950 814.050 871.050 ;
        RECT 713.100 865.950 715.200 868.050 ;
        RECT 713.400 826.050 714.600 865.950 ;
        RECT 812.400 862.050 813.600 868.950 ;
        RECT 811.950 859.950 814.050 862.050 ;
        RECT 744.000 834.600 748.050 835.050 ;
        RECT 743.400 834.000 748.050 834.600 ;
        RECT 742.950 832.950 748.050 834.000 ;
        RECT 742.950 829.950 745.050 832.950 ;
        RECT 712.950 823.950 715.050 826.050 ;
        RECT 724.950 823.950 727.050 826.050 ;
        RECT 725.400 781.050 726.600 823.950 ;
        RECT 724.950 778.950 727.050 781.050 ;
        RECT 769.950 778.950 772.050 781.050 ;
        RECT 770.400 748.050 771.600 778.950 ;
        RECT 769.950 745.950 772.050 748.050 ;
        RECT 778.950 745.950 781.050 748.050 ;
        RECT 442.950 742.950 445.050 745.050 ;
        RECT 514.950 742.950 517.050 745.050 ;
        RECT 562.950 742.950 565.050 745.050 ;
        RECT 568.950 742.950 571.050 745.050 ;
        RECT 443.400 736.050 444.600 742.950 ;
        RECT 442.950 733.950 445.050 736.050 ;
        RECT 325.950 718.950 328.050 721.050 ;
        RECT 326.400 715.050 327.600 718.950 ;
        RECT 275.100 712.950 277.200 715.050 ;
        RECT 325.950 712.950 328.050 715.050 ;
        RECT 346.950 712.950 349.050 715.050 ;
        RECT 275.400 661.050 276.600 712.950 ;
        RECT 347.400 700.050 348.600 712.950 ;
        RECT 515.400 706.050 516.600 742.950 ;
        RECT 502.950 703.950 505.050 706.050 ;
        RECT 514.950 703.950 517.050 706.050 ;
        RECT 347.100 697.950 349.200 700.050 ;
        RECT 361.950 697.800 364.050 699.900 ;
        RECT 362.400 688.050 363.600 697.800 ;
        RECT 503.400 688.050 504.600 703.950 ;
        RECT 563.400 694.050 564.600 742.950 ;
        RECT 569.400 730.050 570.600 742.950 ;
        RECT 568.950 727.950 571.050 730.050 ;
        RECT 779.400 727.050 780.600 745.950 ;
        RECT 778.950 724.950 781.050 727.050 ;
        RECT 779.400 721.050 780.600 724.950 ;
        RECT 775.950 719.400 780.600 721.050 ;
        RECT 775.950 718.950 780.000 719.400 ;
        RECT 805.950 712.950 808.050 715.050 ;
        RECT 806.400 700.050 807.600 712.950 ;
        RECT 805.950 697.950 808.050 700.050 ;
        RECT 562.950 691.950 565.050 694.050 ;
        RECT 361.950 685.950 364.050 688.050 ;
        RECT 502.950 685.950 505.050 688.050 ;
        RECT 776.100 667.950 778.200 670.050 ;
        RECT 808.950 667.950 811.050 670.050 ;
        RECT 571.950 664.950 574.050 667.050 ;
        RECT 274.950 658.950 277.050 661.050 ;
        RECT 572.400 652.050 573.600 664.950 ;
        RECT 776.400 655.050 777.600 667.950 ;
        RECT 774.000 654.900 777.600 655.050 ;
        RECT 772.950 653.400 777.600 654.900 ;
        RECT 772.950 652.950 777.000 653.400 ;
        RECT 772.950 652.800 775.050 652.950 ;
        RECT 571.950 649.950 574.050 652.050 ;
        RECT 572.400 634.050 573.600 649.950 ;
        RECT 809.400 640.200 810.600 667.950 ;
        RECT 820.950 640.950 823.050 643.050 ;
        RECT 808.950 638.100 811.050 640.200 ;
        RECT 821.400 637.050 822.600 640.950 ;
        RECT 820.950 634.950 823.050 637.050 ;
        RECT 571.950 631.950 574.050 634.050 ;
        RECT 685.950 631.950 688.050 634.050 ;
        RECT 289.950 628.950 292.050 631.050 ;
        RECT 290.400 601.050 291.600 628.950 ;
        RECT 686.400 616.050 687.600 631.950 ;
        RECT 760.950 628.950 763.050 631.050 ;
        RECT 761.400 616.050 762.600 628.950 ;
        RECT 685.950 613.950 688.050 616.050 ;
        RECT 760.950 613.950 763.050 616.050 ;
        RECT 761.400 610.050 762.600 613.950 ;
        RECT 760.950 607.950 763.050 610.050 ;
        RECT 289.950 598.950 292.050 601.050 ;
    END
  END Cin[4]
  PIN Cin[3]
    PORT
      LAYER metal1 ;
        RECT 605.100 733.950 607.200 736.050 ;
        RECT 605.550 712.050 606.450 733.950 ;
        RECT 604.950 709.950 607.050 712.050 ;
        RECT 286.950 658.950 289.050 661.050 ;
        RECT 325.950 660.450 330.000 661.050 ;
        RECT 325.950 660.000 330.450 660.450 ;
        RECT 325.950 658.950 331.050 660.000 ;
        RECT 287.550 652.050 288.450 658.950 ;
        RECT 328.950 658.050 331.050 658.950 ;
        RECT 328.950 657.000 331.200 658.050 ;
        RECT 329.100 655.950 331.200 657.000 ;
        RECT 286.950 649.950 289.050 652.050 ;
        RECT 409.950 649.950 412.050 652.050 ;
        RECT 410.550 631.050 411.450 649.950 ;
        RECT 409.800 628.950 411.900 631.050 ;
      LAYER metal2 ;
        RECT 793.950 897.450 796.050 898.050 ;
        RECT 802.950 897.450 805.050 898.050 ;
        RECT 793.950 896.400 805.050 897.450 ;
        RECT 793.950 895.950 796.050 896.400 ;
        RECT 802.950 895.950 805.050 896.400 ;
        RECT 751.950 886.950 754.050 889.050 ;
        RECT 793.950 870.450 796.050 871.200 ;
        RECT 788.400 869.400 796.050 870.450 ;
        RECT 745.950 867.450 748.050 868.050 ;
        RECT 772.950 867.450 775.050 868.050 ;
        RECT 788.400 867.450 789.450 869.400 ;
        RECT 793.950 869.100 796.050 869.400 ;
        RECT 745.950 866.400 789.450 867.450 ;
        RECT 745.950 865.950 748.050 866.400 ;
        RECT 772.950 865.950 775.050 866.400 ;
        RECT 739.950 852.450 742.050 853.050 ;
        RECT 745.800 852.450 747.900 853.050 ;
        RECT 739.950 851.400 747.900 852.450 ;
        RECT 739.950 850.950 742.050 851.400 ;
        RECT 745.800 850.950 747.900 851.400 ;
        RECT 772.950 832.950 775.050 835.050 ;
        RECT 739.950 774.450 742.050 775.200 ;
        RECT 781.950 774.450 784.050 775.050 ;
        RECT 739.950 773.400 784.050 774.450 ;
        RECT 739.950 773.100 742.050 773.400 ;
        RECT 781.950 772.950 784.050 773.400 ;
        RECT 583.950 771.450 586.050 772.050 ;
        RECT 607.950 771.450 610.050 772.050 ;
        RECT 583.950 770.400 610.050 771.450 ;
        RECT 583.950 769.950 586.050 770.400 ;
        RECT 607.950 769.950 610.050 770.400 ;
        RECT 583.800 750.450 585.900 751.050 ;
        RECT 575.400 749.400 585.900 750.450 ;
        RECT 418.950 747.450 421.050 748.050 ;
        RECT 433.950 747.450 436.050 748.050 ;
        RECT 418.950 746.400 436.050 747.450 ;
        RECT 418.950 745.950 421.050 746.400 ;
        RECT 433.950 745.950 436.050 746.400 ;
        RECT 506.100 747.450 508.200 748.050 ;
        RECT 547.950 747.450 550.050 748.050 ;
        RECT 575.400 747.450 576.450 749.400 ;
        RECT 583.800 748.950 585.900 749.400 ;
        RECT 506.100 746.400 576.450 747.450 ;
        RECT 506.100 745.950 508.200 746.400 ;
        RECT 547.950 745.950 550.050 746.400 ;
        RECT 434.100 741.450 436.200 742.050 ;
        RECT 505.950 741.450 508.050 742.050 ;
        RECT 434.100 740.400 508.050 741.450 ;
        RECT 434.100 739.950 436.200 740.400 ;
        RECT 505.950 739.950 508.050 740.400 ;
        RECT 605.100 733.950 610.050 736.050 ;
        RECT 544.950 727.950 550.050 730.050 ;
        RECT 280.950 718.950 283.050 721.050 ;
        RECT 604.950 711.450 607.050 712.050 ;
        RECT 610.950 711.450 613.050 712.050 ;
        RECT 604.950 710.400 613.050 711.450 ;
        RECT 604.950 709.950 607.050 710.400 ;
        RECT 610.950 709.950 613.050 710.400 ;
        RECT 673.950 708.450 676.050 709.050 ;
        RECT 706.950 708.450 709.050 709.050 ;
        RECT 673.950 707.400 709.050 708.450 ;
        RECT 673.950 706.950 676.050 707.400 ;
        RECT 706.950 706.950 709.050 707.400 ;
        RECT 280.950 705.450 283.050 706.050 ;
        RECT 784.950 705.450 787.050 706.050 ;
        RECT 790.950 705.450 793.050 706.050 ;
        RECT 269.400 704.400 283.050 705.450 ;
        RECT 244.950 702.450 247.050 703.050 ;
        RECT 269.400 702.450 270.450 704.400 ;
        RECT 280.950 703.950 283.050 704.400 ;
        RECT 770.400 704.400 793.050 705.450 ;
        RECT 244.950 701.400 270.450 702.450 ;
        RECT 706.950 702.450 709.050 703.050 ;
        RECT 736.950 702.450 739.050 702.900 ;
        RECT 770.400 702.450 771.450 704.400 ;
        RECT 784.950 703.950 787.050 704.400 ;
        RECT 790.950 703.950 793.050 704.400 ;
        RECT 706.950 701.400 771.450 702.450 ;
        RECT 244.950 700.950 247.050 701.400 ;
        RECT 706.950 700.950 709.050 701.400 ;
        RECT 736.950 700.800 739.050 701.400 ;
        RECT 604.950 693.450 607.050 694.050 ;
        RECT 610.800 693.450 612.900 694.050 ;
        RECT 604.950 692.400 612.900 693.450 ;
        RECT 604.950 691.950 607.050 692.400 ;
        RECT 610.800 691.950 612.900 692.400 ;
        RECT 244.950 685.950 247.050 688.050 ;
        RECT 604.950 687.450 607.050 688.050 ;
        RECT 616.950 687.450 619.050 688.050 ;
        RECT 604.950 686.400 619.050 687.450 ;
        RECT 604.950 685.950 607.050 686.400 ;
        RECT 616.950 685.950 619.050 686.400 ;
        RECT 673.950 685.950 676.050 688.050 ;
        RECT 736.950 685.950 739.050 688.050 ;
        RECT 793.950 678.450 796.050 679.050 ;
        RECT 799.950 678.450 802.050 679.050 ;
        RECT 793.950 677.400 802.050 678.450 ;
        RECT 793.950 676.950 796.050 677.400 ;
        RECT 799.950 676.950 802.050 677.400 ;
        RECT 247.950 666.450 250.050 667.050 ;
        RECT 286.950 666.450 289.050 667.050 ;
        RECT 673.950 666.450 676.050 667.050 ;
        RECT 247.950 665.400 289.050 666.450 ;
        RECT 247.950 664.950 250.050 665.400 ;
        RECT 286.950 664.950 289.050 665.400 ;
        RECT 665.400 665.400 676.050 666.450 ;
        RECT 616.950 663.450 619.050 664.050 ;
        RECT 665.400 663.450 666.450 665.400 ;
        RECT 673.950 664.950 676.050 665.400 ;
        RECT 616.950 662.400 666.450 663.450 ;
        RECT 616.950 661.950 619.050 662.400 ;
        RECT 286.950 660.450 289.050 661.050 ;
        RECT 325.950 660.450 328.050 661.050 ;
        RECT 286.950 659.400 328.050 660.450 ;
        RECT 286.950 658.950 289.050 659.400 ;
        RECT 325.950 658.950 328.050 659.400 ;
        RECT 673.950 660.450 676.050 661.050 ;
        RECT 685.950 660.450 688.050 660.900 ;
        RECT 673.950 659.400 688.050 660.450 ;
        RECT 673.950 658.950 676.050 659.400 ;
        RECT 685.950 658.800 688.050 659.400 ;
        RECT 329.100 657.450 331.200 658.050 ;
        RECT 352.950 657.450 355.050 658.050 ;
        RECT 329.100 656.400 355.050 657.450 ;
        RECT 329.100 655.950 331.200 656.400 ;
        RECT 352.950 655.950 355.050 656.400 ;
        RECT 271.950 649.950 274.050 652.050 ;
        RECT 277.950 651.450 280.050 652.050 ;
        RECT 286.950 651.450 289.050 652.050 ;
        RECT 277.950 650.400 289.050 651.450 ;
        RECT 277.950 649.950 280.050 650.400 ;
        RECT 286.950 649.950 289.050 650.400 ;
        RECT 409.950 651.450 412.050 652.050 ;
        RECT 415.950 651.450 418.050 652.050 ;
        RECT 409.950 650.400 418.050 651.450 ;
        RECT 409.950 649.950 412.050 650.400 ;
        RECT 415.950 649.950 418.050 650.400 ;
        RECT 685.950 649.950 688.050 652.050 ;
        RECT 802.950 640.950 805.050 643.050 ;
        RECT 400.950 630.450 403.050 631.050 ;
        RECT 409.800 630.450 411.900 631.050 ;
        RECT 400.950 629.400 411.900 630.450 ;
        RECT 400.950 628.950 403.050 629.400 ;
        RECT 409.800 628.950 411.900 629.400 ;
        RECT 352.950 627.450 355.050 628.050 ;
        RECT 352.950 627.000 366.450 627.450 ;
        RECT 352.950 626.400 367.050 627.000 ;
        RECT 352.950 625.950 355.050 626.400 ;
        RECT 364.950 625.050 367.050 626.400 ;
        RECT 364.950 624.000 367.200 625.050 ;
        RECT 365.100 622.950 367.200 624.000 ;
        RECT 364.950 618.450 367.050 619.050 ;
        RECT 400.950 618.450 403.050 619.050 ;
        RECT 364.950 617.400 403.050 618.450 ;
        RECT 364.950 616.950 367.050 617.400 ;
        RECT 400.950 616.950 403.050 617.400 ;
      LAYER metal3 ;
        RECT 803.400 905.400 807.600 906.600 ;
        RECT 803.400 898.050 804.600 905.400 ;
        RECT 793.950 895.950 796.050 898.050 ;
        RECT 802.950 895.950 805.050 898.050 ;
        RECT 751.950 885.600 754.050 889.050 ;
        RECT 746.400 885.000 754.050 885.600 ;
        RECT 746.400 884.400 753.600 885.000 ;
        RECT 746.400 868.050 747.600 884.400 ;
        RECT 794.400 871.200 795.600 895.950 ;
        RECT 793.950 869.100 796.050 871.200 ;
        RECT 745.950 865.950 748.050 868.050 ;
        RECT 772.950 865.950 775.050 868.050 ;
        RECT 746.400 853.050 747.600 865.950 ;
        RECT 773.400 855.600 774.600 865.950 ;
        RECT 770.400 854.400 774.600 855.600 ;
        RECT 739.950 850.950 742.050 853.050 ;
        RECT 745.800 850.950 747.900 853.050 ;
        RECT 740.400 775.200 741.600 850.950 ;
        RECT 770.400 835.050 771.600 854.400 ;
        RECT 770.400 833.400 775.050 835.050 ;
        RECT 771.000 832.950 775.050 833.400 ;
        RECT 739.950 773.100 742.050 775.200 ;
        RECT 781.950 772.950 784.050 775.050 ;
        RECT 583.950 769.950 586.050 772.050 ;
        RECT 607.950 769.950 610.050 772.050 ;
        RECT 584.400 751.050 585.600 769.950 ;
        RECT 583.800 748.950 585.900 751.050 ;
        RECT 418.950 745.950 421.050 748.050 ;
        RECT 433.950 745.950 436.050 748.050 ;
        RECT 506.100 745.950 508.200 748.050 ;
        RECT 547.950 745.950 550.050 748.050 ;
        RECT 419.400 723.600 420.600 745.950 ;
        RECT 434.400 742.050 435.600 745.950 ;
        RECT 506.400 742.050 507.600 745.950 ;
        RECT 434.100 739.950 436.200 742.050 ;
        RECT 505.950 739.950 508.050 742.050 ;
        RECT 548.400 730.050 549.600 745.950 ;
        RECT 608.400 736.050 609.600 769.950 ;
        RECT 607.950 733.950 610.050 736.050 ;
        RECT 547.950 727.950 550.050 730.050 ;
        RECT 413.400 722.400 420.600 723.600 ;
        RECT 280.950 718.950 283.050 721.050 ;
        RECT 281.400 706.050 282.600 718.950 ;
        RECT 413.400 708.600 414.600 722.400 ;
        RECT 782.400 720.600 783.600 772.950 ;
        RECT 782.400 719.400 786.600 720.600 ;
        RECT 610.950 709.950 613.050 712.050 ;
        RECT 413.400 707.400 417.600 708.600 ;
        RECT 280.950 703.950 283.050 706.050 ;
        RECT 244.950 700.950 247.050 703.050 ;
        RECT 245.400 688.050 246.600 700.950 ;
        RECT 244.950 687.600 249.000 688.050 ;
        RECT 244.950 685.950 249.600 687.600 ;
        RECT 248.400 667.050 249.600 685.950 ;
        RECT 247.950 664.950 250.050 667.050 ;
        RECT 286.950 664.950 289.050 667.050 ;
        RECT 287.400 661.050 288.600 664.950 ;
        RECT 286.950 658.950 289.050 661.050 ;
        RECT 352.950 655.950 355.050 658.050 ;
        RECT 271.950 651.600 274.050 652.050 ;
        RECT 277.950 651.600 280.050 652.050 ;
        RECT 271.950 650.400 280.050 651.600 ;
        RECT 271.950 649.950 274.050 650.400 ;
        RECT 277.950 649.950 280.050 650.400 ;
        RECT 353.400 628.050 354.600 655.950 ;
        RECT 416.400 652.050 417.600 707.400 ;
        RECT 611.400 694.050 612.600 709.950 ;
        RECT 673.950 706.950 676.050 709.050 ;
        RECT 706.950 706.950 709.050 709.050 ;
        RECT 674.400 696.600 675.600 706.950 ;
        RECT 707.400 703.050 708.600 706.950 ;
        RECT 785.400 706.050 786.600 719.400 ;
        RECT 784.950 703.950 787.050 706.050 ;
        RECT 790.950 703.950 793.050 706.050 ;
        RECT 706.950 700.950 709.050 703.050 ;
        RECT 736.950 700.800 739.050 702.900 ;
        RECT 671.400 695.400 675.600 696.600 ;
        RECT 604.950 691.950 607.050 694.050 ;
        RECT 610.800 691.950 612.900 694.050 ;
        RECT 605.400 688.050 606.600 691.950 ;
        RECT 671.400 690.600 672.600 695.400 ;
        RECT 671.400 689.400 675.600 690.600 ;
        RECT 674.400 688.050 675.600 689.400 ;
        RECT 737.400 688.050 738.600 700.800 ;
        RECT 604.950 685.950 607.050 688.050 ;
        RECT 616.950 685.950 619.050 688.050 ;
        RECT 673.950 685.950 676.050 688.050 ;
        RECT 736.950 685.950 739.050 688.050 ;
        RECT 617.400 664.050 618.600 685.950 ;
        RECT 674.400 667.050 675.600 685.950 ;
        RECT 791.400 681.600 792.600 703.950 ;
        RECT 791.400 681.000 795.600 681.600 ;
        RECT 791.400 680.400 796.050 681.000 ;
        RECT 793.950 676.950 796.050 680.400 ;
        RECT 799.950 676.950 802.050 679.050 ;
        RECT 673.950 664.950 676.050 667.050 ;
        RECT 616.950 661.950 619.050 664.050 ;
        RECT 674.400 661.050 675.600 664.950 ;
        RECT 673.950 658.950 676.050 661.050 ;
        RECT 685.950 658.800 688.050 660.900 ;
        RECT 686.400 652.050 687.600 658.800 ;
        RECT 415.950 649.950 418.050 652.050 ;
        RECT 685.950 649.950 688.050 652.050 ;
        RECT 800.400 643.050 801.600 676.950 ;
        RECT 800.400 641.400 805.050 643.050 ;
        RECT 801.000 640.950 805.050 641.400 ;
        RECT 400.950 628.950 403.050 631.050 ;
        RECT 352.950 625.950 355.050 628.050 ;
        RECT 365.100 622.950 367.200 625.050 ;
        RECT 365.400 619.050 366.600 622.950 ;
        RECT 401.400 619.050 402.600 628.950 ;
        RECT 364.950 616.950 367.050 619.050 ;
        RECT 400.950 616.950 403.050 619.050 ;
    END
  END Cin[3]
  PIN Cin[2]
    PORT
      LAYER metal1 ;
        RECT 791.100 892.950 793.200 895.050 ;
        RECT 791.550 868.050 792.450 892.950 ;
        RECT 790.950 865.950 793.050 868.050 ;
        RECT 553.800 855.000 555.900 856.050 ;
        RECT 553.800 853.950 556.050 855.000 ;
        RECT 553.950 853.050 556.050 853.950 ;
        RECT 553.950 852.000 559.050 853.050 ;
        RECT 554.550 851.550 559.050 852.000 ;
        RECT 555.000 850.950 559.050 851.550 ;
      LAYER metal2 ;
        RECT 217.950 900.450 220.050 901.050 ;
        RECT 217.950 899.400 528.450 900.450 ;
        RECT 217.950 898.950 220.050 899.400 ;
        RECT 527.400 897.450 528.450 899.400 ;
        RECT 556.950 897.450 559.050 898.050 ;
        RECT 527.400 896.400 559.050 897.450 ;
        RECT 556.950 895.950 559.050 896.400 ;
        RECT 791.100 894.450 793.200 895.050 ;
        RECT 799.950 894.450 802.050 895.050 ;
        RECT 805.950 894.450 808.050 895.050 ;
        RECT 791.100 893.400 808.050 894.450 ;
        RECT 791.100 892.950 793.200 893.400 ;
        RECT 799.950 892.950 802.050 893.400 ;
        RECT 805.950 892.950 808.050 893.400 ;
        RECT 805.950 886.950 808.050 889.050 ;
        RECT 217.950 874.950 220.050 877.050 ;
        RECT 550.950 876.450 553.050 877.050 ;
        RECT 555.000 876.450 559.050 877.050 ;
        RECT 550.950 875.400 559.050 876.450 ;
        RECT 550.950 871.950 553.050 875.400 ;
        RECT 555.000 874.950 559.050 875.400 ;
        RECT 790.950 867.900 795.000 868.050 ;
        RECT 790.950 865.950 796.050 867.900 ;
        RECT 793.950 865.800 796.050 865.950 ;
        RECT 217.950 861.450 220.050 862.050 ;
        RECT 256.950 861.450 259.050 862.050 ;
        RECT 217.950 860.400 259.050 861.450 ;
        RECT 217.950 859.950 220.050 860.400 ;
        RECT 256.950 859.950 259.050 860.400 ;
        RECT 550.950 856.050 553.050 856.200 ;
        RECT 499.950 855.450 502.050 856.050 ;
        RECT 550.950 855.450 555.900 856.050 ;
        RECT 499.950 854.400 555.900 855.450 ;
        RECT 499.950 853.950 502.050 854.400 ;
        RECT 550.950 854.100 555.900 854.400 ;
        RECT 552.000 853.950 555.900 854.100 ;
        RECT 556.950 850.950 562.050 853.050 ;
        RECT 697.950 849.450 700.050 850.050 ;
        RECT 793.950 849.450 796.050 850.050 ;
        RECT 697.950 848.400 796.050 849.450 ;
        RECT 697.950 847.950 700.050 848.400 ;
        RECT 793.950 847.950 796.050 848.400 ;
        RECT 502.950 841.950 505.050 844.050 ;
        RECT 697.950 841.950 700.050 844.050 ;
        RECT 793.950 841.950 796.050 844.050 ;
        RECT 562.950 822.450 565.050 823.050 ;
        RECT 697.950 822.450 700.050 823.050 ;
        RECT 562.950 821.400 700.050 822.450 ;
        RECT 562.950 820.950 565.050 821.400 ;
        RECT 697.950 820.950 700.050 821.400 ;
        RECT 205.950 771.450 208.050 772.050 ;
        RECT 235.950 771.450 238.050 772.050 ;
        RECT 256.950 771.450 259.050 772.050 ;
        RECT 205.950 770.400 259.050 771.450 ;
        RECT 205.950 769.950 208.050 770.400 ;
        RECT 235.950 769.950 238.050 770.400 ;
        RECT 256.950 769.950 259.050 770.400 ;
        RECT 202.950 763.950 205.050 766.050 ;
        RECT 235.950 718.950 238.050 721.050 ;
      LAYER metal3 ;
        RECT 217.950 898.950 220.050 901.050 ;
        RECT 218.400 877.050 219.600 898.950 ;
        RECT 556.950 895.950 559.050 898.050 ;
        RECT 557.400 877.050 558.600 895.950 ;
        RECT 800.400 895.050 801.600 906.600 ;
        RECT 799.950 892.950 802.050 895.050 ;
        RECT 805.950 892.950 808.050 895.050 ;
        RECT 806.400 889.050 807.600 892.950 ;
        RECT 805.950 886.950 808.050 889.050 ;
        RECT 217.950 874.950 220.050 877.050 ;
        RECT 556.950 874.950 559.050 877.050 ;
        RECT 218.400 862.050 219.600 874.950 ;
        RECT 550.950 871.950 553.050 874.050 ;
        RECT 217.950 859.950 220.050 862.050 ;
        RECT 256.950 859.950 259.050 862.050 ;
        RECT 257.400 772.050 258.600 859.950 ;
        RECT 551.400 856.200 552.600 871.950 ;
        RECT 793.950 865.800 796.050 867.900 ;
        RECT 499.950 853.950 502.050 856.050 ;
        RECT 550.950 854.100 553.050 856.200 ;
        RECT 500.400 844.050 501.600 853.950 ;
        RECT 559.950 850.950 562.050 853.050 ;
        RECT 500.400 842.400 505.050 844.050 ;
        RECT 501.000 841.950 505.050 842.400 ;
        RECT 560.400 825.600 561.600 850.950 ;
        RECT 794.400 850.050 795.600 865.800 ;
        RECT 697.950 847.950 700.050 850.050 ;
        RECT 793.950 847.950 796.050 850.050 ;
        RECT 698.400 844.050 699.600 847.950 ;
        RECT 794.400 844.050 795.600 847.950 ;
        RECT 697.950 841.950 700.050 844.050 ;
        RECT 793.950 841.950 796.050 844.050 ;
        RECT 560.400 825.000 564.600 825.600 ;
        RECT 560.400 824.400 565.050 825.000 ;
        RECT 562.950 820.950 565.050 824.400 ;
        RECT 698.400 823.050 699.600 841.950 ;
        RECT 697.950 820.950 700.050 823.050 ;
        RECT 205.950 769.950 208.050 772.050 ;
        RECT 235.950 769.950 238.050 772.050 ;
        RECT 256.950 769.950 259.050 772.050 ;
        RECT 206.400 766.050 207.600 769.950 ;
        RECT 202.950 764.400 207.600 766.050 ;
        RECT 202.950 763.950 207.000 764.400 ;
        RECT 236.400 721.050 237.600 769.950 ;
        RECT 235.950 718.950 238.050 721.050 ;
    END
  END Cin[2]
  PIN Cin[1]
    PORT
      LAYER metal2 ;
        RECT 289.950 894.450 292.050 895.050 ;
        RECT 301.950 894.450 304.050 895.050 ;
        RECT 613.950 894.450 616.050 895.050 ;
        RECT 289.950 893.400 648.450 894.450 ;
        RECT 289.950 892.950 292.050 893.400 ;
        RECT 301.950 892.950 304.050 893.400 ;
        RECT 613.950 892.950 616.050 893.400 ;
        RECT 647.400 891.450 648.450 893.400 ;
        RECT 697.950 891.450 700.050 892.050 ;
        RECT 647.400 890.400 700.050 891.450 ;
        RECT 668.400 886.050 669.450 890.400 ;
        RECT 697.950 889.950 700.050 890.400 ;
        RECT 289.950 883.950 292.050 886.050 ;
        RECT 301.950 883.950 304.050 886.050 ;
        RECT 667.950 883.950 670.050 886.050 ;
        RECT 697.950 883.950 700.050 886.050 ;
      LAYER metal3 ;
        RECT 614.400 895.050 615.600 906.600 ;
        RECT 289.950 892.950 292.050 895.050 ;
        RECT 301.950 892.950 304.050 895.050 ;
        RECT 613.950 892.950 616.050 895.050 ;
        RECT 290.400 886.050 291.600 892.950 ;
        RECT 302.400 886.050 303.600 892.950 ;
        RECT 697.950 889.950 700.050 892.050 ;
        RECT 698.400 886.050 699.600 889.950 ;
        RECT 289.950 883.950 292.050 886.050 ;
        RECT 301.950 883.950 304.050 886.050 ;
        RECT 697.950 883.950 700.050 886.050 ;
    END
  END Cin[1]
  PIN Cin[0]
    PORT
      LAYER metal2 ;
        RECT 451.950 883.950 454.050 886.050 ;
        RECT 607.950 883.950 613.050 886.050 ;
        RECT 250.950 870.450 253.050 871.050 ;
        RECT 346.950 870.450 349.050 871.050 ;
        RECT 451.950 870.450 454.050 871.050 ;
        RECT 610.950 870.450 613.050 871.200 ;
        RECT 250.950 869.400 613.050 870.450 ;
        RECT 250.950 868.950 253.050 869.400 ;
        RECT 346.950 868.950 349.050 869.400 ;
        RECT 451.950 868.950 454.050 869.400 ;
        RECT 610.950 869.100 613.050 869.400 ;
        RECT 346.950 832.950 349.050 835.050 ;
        RECT 247.950 805.950 250.050 808.050 ;
      LAYER metal3 ;
        RECT 608.400 886.050 609.600 906.600 ;
        RECT 451.950 883.950 454.050 886.050 ;
        RECT 607.950 883.950 610.050 886.050 ;
        RECT 610.950 883.950 613.050 886.050 ;
        RECT 452.400 871.050 453.600 883.950 ;
        RECT 611.400 871.200 612.600 883.950 ;
        RECT 250.950 868.950 253.050 871.050 ;
        RECT 346.950 868.950 349.050 871.050 ;
        RECT 451.950 868.950 454.050 871.050 ;
        RECT 610.950 869.100 613.050 871.200 ;
        RECT 251.400 810.600 252.600 868.950 ;
        RECT 347.400 835.050 348.600 868.950 ;
        RECT 346.950 832.950 349.050 835.050 ;
        RECT 248.400 810.000 252.600 810.600 ;
        RECT 247.950 809.400 252.600 810.000 ;
        RECT 247.950 805.950 250.050 809.400 ;
    END
  END Cin[0]
  PIN Rdy
    PORT
      LAYER metal2 ;
        RECT -3.600 405.450 -2.550 411.450 ;
        RECT 13.950 406.950 16.050 412.050 ;
        RECT 4.950 405.450 7.050 406.050 ;
        RECT -3.600 404.400 7.050 405.450 ;
        RECT 4.950 403.950 7.050 404.400 ;
      LAYER metal3 ;
        RECT 4.950 405.600 7.050 406.050 ;
        RECT 13.950 405.600 16.050 409.050 ;
        RECT 4.950 405.000 16.050 405.600 ;
        RECT 4.950 404.400 15.600 405.000 ;
        RECT 4.950 403.950 7.050 404.400 ;
    END
  END Rdy
  PIN Vld
    PORT
      LAYER metal2 ;
        RECT 901.950 255.450 904.050 256.050 ;
        RECT 901.950 254.400 918.450 255.450 ;
        RECT 901.950 253.950 904.050 254.400 ;
    END
  END Vld
  PIN Xin[3]
    PORT
      LAYER metal2 ;
        RECT 32.100 630.450 34.200 631.050 ;
        RECT 241.950 630.450 244.050 631.050 ;
        RECT 32.100 629.400 244.050 630.450 ;
        RECT 32.100 628.950 34.200 629.400 ;
        RECT 241.950 628.950 244.050 629.400 ;
        RECT 31.950 615.450 34.050 616.050 ;
        RECT 241.950 615.450 244.050 616.050 ;
        RECT -3.600 614.400 34.050 615.450 ;
        RECT -3.600 611.400 -2.550 614.400 ;
        RECT 31.950 613.950 34.050 614.400 ;
        RECT 227.400 614.400 244.050 615.450 ;
        RECT 227.400 610.050 228.450 614.400 ;
        RECT 241.950 613.950 244.050 614.400 ;
        RECT 226.950 607.950 229.050 610.050 ;
        RECT 241.950 607.950 244.050 610.050 ;
      LAYER metal3 ;
        RECT 32.100 628.950 34.200 631.050 ;
        RECT 241.950 628.950 244.050 631.050 ;
        RECT 32.400 616.050 33.600 628.950 ;
        RECT 242.400 616.050 243.600 628.950 ;
        RECT 31.950 613.950 34.050 616.050 ;
        RECT 241.950 613.950 244.050 616.050 ;
        RECT 242.400 610.050 243.600 613.950 ;
        RECT 241.950 607.950 244.050 610.050 ;
    END
  END Xin[3]
  PIN Xin[2]
    PORT
      LAYER metal2 ;
        RECT 1.950 618.450 4.050 619.050 ;
        RECT 49.950 618.450 52.050 619.050 ;
        RECT 1.950 617.400 52.050 618.450 ;
        RECT 1.950 616.950 4.050 617.400 ;
        RECT 49.950 616.950 52.050 617.400 ;
        RECT 49.950 609.450 52.050 610.050 ;
        RECT 58.950 609.450 61.050 610.050 ;
        RECT 49.950 608.400 61.050 609.450 ;
        RECT 49.950 607.950 52.050 608.400 ;
        RECT 58.950 607.950 61.050 608.400 ;
        RECT 262.950 607.950 265.050 610.050 ;
        RECT 1.950 606.450 4.050 607.050 ;
        RECT -3.600 605.400 4.050 606.450 ;
        RECT 1.950 604.950 4.050 605.400 ;
        RECT 61.950 588.450 64.050 589.050 ;
        RECT 262.950 588.450 265.050 589.050 ;
        RECT 61.950 587.400 265.050 588.450 ;
        RECT 61.950 586.950 64.050 587.400 ;
        RECT 262.950 586.950 265.050 587.400 ;
      LAYER metal3 ;
        RECT 1.950 616.950 4.050 619.050 ;
        RECT 49.950 616.950 52.050 619.050 ;
        RECT 2.400 607.050 3.600 616.950 ;
        RECT 50.400 610.050 51.600 616.950 ;
        RECT 49.950 607.950 52.050 610.050 ;
        RECT 1.950 604.950 4.050 607.050 ;
        RECT 58.950 606.600 61.050 610.050 ;
        RECT 262.950 607.950 265.050 610.050 ;
        RECT 58.950 606.000 63.600 606.600 ;
        RECT 59.400 605.400 63.600 606.000 ;
        RECT 62.400 589.050 63.600 605.400 ;
        RECT 263.400 589.050 264.600 607.950 ;
        RECT 61.950 586.950 64.050 589.050 ;
        RECT 262.950 586.950 265.050 589.050 ;
    END
  END Xin[2]
  PIN Xin[1]
    PORT
      LAYER metal1 ;
        RECT 163.950 562.950 166.050 565.050 ;
        RECT 164.550 553.050 165.450 562.950 ;
        RECT 163.950 550.950 166.050 553.050 ;
      LAYER metal2 ;
        RECT 1.950 567.450 4.050 568.050 ;
        RECT -3.600 566.400 4.050 567.450 ;
        RECT 1.950 565.950 4.050 566.400 ;
        RECT 151.950 564.450 154.050 565.050 ;
        RECT 163.950 564.450 166.050 565.050 ;
        RECT 151.950 563.400 166.050 564.450 ;
        RECT 151.950 559.950 154.050 563.400 ;
        RECT 163.950 562.950 166.050 563.400 ;
        RECT 250.950 562.950 253.050 565.050 ;
        RECT 163.950 552.450 166.050 553.050 ;
        RECT 250.950 552.450 253.050 553.050 ;
        RECT 163.950 551.400 253.050 552.450 ;
        RECT 163.950 550.950 166.050 551.400 ;
        RECT 250.950 550.950 253.050 551.400 ;
        RECT 1.950 549.450 4.050 550.050 ;
        RECT 1.950 548.400 81.450 549.450 ;
        RECT 1.950 547.950 4.050 548.400 ;
        RECT 80.400 546.450 81.450 548.400 ;
        RECT 151.950 546.450 154.050 547.050 ;
        RECT 80.400 545.400 154.050 546.450 ;
        RECT 151.950 544.950 154.050 545.400 ;
      LAYER metal3 ;
        RECT 1.950 565.950 4.050 568.050 ;
        RECT 2.400 550.050 3.600 565.950 ;
        RECT 250.950 562.950 253.050 565.050 ;
        RECT 151.950 559.950 154.050 562.050 ;
        RECT 1.950 547.950 4.050 550.050 ;
        RECT 152.400 547.050 153.600 559.950 ;
        RECT 251.400 553.050 252.600 562.950 ;
        RECT 250.950 550.950 253.050 553.050 ;
        RECT 151.950 544.950 154.050 547.050 ;
    END
  END Xin[1]
  PIN Xin[0]
    PORT
      LAYER metal1 ;
        RECT 190.950 541.950 193.050 544.050 ;
        RECT 191.550 532.050 192.450 541.950 ;
        RECT 190.950 529.950 193.050 532.050 ;
      LAYER metal2 ;
        RECT 406.950 562.950 409.050 565.050 ;
        RECT 406.950 546.450 409.050 547.050 ;
        RECT 341.400 545.400 409.050 546.450 ;
        RECT 1.950 543.450 4.050 544.050 ;
        RECT 190.950 543.450 193.050 544.050 ;
        RECT 341.400 543.450 342.450 545.400 ;
        RECT 406.950 544.950 409.050 545.400 ;
        RECT 1.950 542.400 342.450 543.450 ;
        RECT 1.950 541.950 4.050 542.400 ;
        RECT 190.950 541.950 193.050 542.400 ;
        RECT 1.950 531.450 4.050 532.050 ;
        RECT -3.600 530.400 4.050 531.450 ;
        RECT 1.950 529.950 4.050 530.400 ;
        RECT 190.950 531.450 193.050 532.050 ;
        RECT 202.950 531.450 205.050 532.050 ;
        RECT 190.950 530.400 205.050 531.450 ;
        RECT 190.950 529.950 193.050 530.400 ;
        RECT 202.950 529.950 205.050 530.400 ;
      LAYER metal3 ;
        RECT 406.950 562.950 409.050 565.050 ;
        RECT 407.400 547.050 408.600 562.950 ;
        RECT 406.950 544.950 409.050 547.050 ;
        RECT 1.950 541.950 4.050 544.050 ;
        RECT 2.400 532.050 3.600 541.950 ;
        RECT 1.950 529.950 4.050 532.050 ;
    END
  END Xin[0]
  PIN Xout[3]
    PORT
      LAYER metal2 ;
        RECT 895.950 777.450 898.050 778.050 ;
        RECT 895.950 776.400 912.450 777.450 ;
        RECT 895.950 775.950 898.050 776.400 ;
        RECT 911.400 774.450 912.450 776.400 ;
        RECT 911.400 773.400 918.450 774.450 ;
        RECT 917.400 767.400 918.450 773.400 ;
        RECT 883.950 762.450 886.050 763.050 ;
        RECT 895.950 762.450 898.050 763.200 ;
        RECT 883.950 761.400 898.050 762.450 ;
        RECT 883.950 760.950 886.050 761.400 ;
        RECT 895.950 761.100 898.050 761.400 ;
      LAYER metal3 ;
        RECT 895.950 775.950 898.050 778.050 ;
        RECT 896.400 763.200 897.600 775.950 ;
        RECT 895.950 761.100 898.050 763.200 ;
    END
  END Xout[3]
  PIN Xout[2]
    PORT
      LAYER metal1 ;
        RECT 850.950 772.950 853.050 775.050 ;
        RECT 907.950 772.950 910.050 775.050 ;
        RECT 851.550 763.050 852.450 772.950 ;
        RECT 908.550 766.050 909.450 772.950 ;
        RECT 907.950 763.950 910.050 766.050 ;
        RECT 850.950 760.950 853.050 763.050 ;
      LAYER metal2 ;
        RECT 850.950 774.450 853.050 775.050 ;
        RECT 907.950 774.450 910.050 775.050 ;
        RECT 850.950 773.400 910.050 774.450 ;
        RECT 850.950 772.950 853.050 773.400 ;
        RECT 907.950 772.950 910.050 773.400 ;
        RECT 907.950 765.450 910.050 766.050 ;
        RECT 907.950 764.400 915.450 765.450 ;
        RECT 907.950 763.950 910.050 764.400 ;
        RECT 838.950 762.450 841.050 763.050 ;
        RECT 850.950 762.450 853.050 763.050 ;
        RECT 838.950 761.400 853.050 762.450 ;
        RECT 914.400 762.450 915.450 764.400 ;
        RECT 914.400 761.400 918.450 762.450 ;
        RECT 838.950 760.950 841.050 761.400 ;
        RECT 850.950 760.950 853.050 761.400 ;
    END
  END Xout[2]
  PIN Xout[1]
    PORT
      LAYER metal1 ;
        RECT 904.950 715.950 907.050 718.050 ;
        RECT 905.550 709.050 906.450 715.950 ;
        RECT 904.800 706.950 906.900 709.050 ;
      LAYER metal2 ;
        RECT 853.950 723.450 856.050 724.050 ;
        RECT 862.950 723.450 865.050 724.050 ;
        RECT 853.950 722.400 865.050 723.450 ;
        RECT 853.950 721.950 856.050 722.400 ;
        RECT 862.950 721.950 865.050 722.400 ;
        RECT 908.100 723.450 910.200 724.050 ;
        RECT 908.100 722.400 918.450 723.450 ;
        RECT 908.100 721.950 910.200 722.400 ;
        RECT 904.950 715.950 910.050 718.050 ;
        RECT 862.950 708.450 865.050 709.050 ;
        RECT 904.800 708.450 906.900 709.050 ;
        RECT 862.950 707.400 906.900 708.450 ;
        RECT 862.950 706.950 865.050 707.400 ;
        RECT 904.800 706.950 906.900 707.400 ;
      LAYER metal3 ;
        RECT 862.950 721.950 865.050 724.050 ;
        RECT 908.100 721.950 910.200 724.050 ;
        RECT 863.400 709.050 864.600 721.950 ;
        RECT 908.400 718.050 909.600 721.950 ;
        RECT 907.950 715.950 910.050 718.050 ;
        RECT 862.950 706.950 865.050 709.050 ;
    END
  END Xout[1]
  PIN Xout[0]
    PORT
      LAYER metal2 ;
        RECT 904.950 567.450 907.050 568.050 ;
        RECT 904.950 566.400 918.450 567.450 ;
        RECT 904.950 565.950 907.050 566.400 ;
    END
  END Xout[0]
  PIN Yin[3]
    PORT
      LAYER metal2 ;
        RECT 520.950 52.950 526.050 55.050 ;
        RECT 517.950 3.450 520.050 4.050 ;
        RECT 523.950 3.450 526.050 4.050 ;
        RECT 517.950 2.400 526.050 3.450 ;
        RECT 517.950 1.950 520.050 2.400 ;
        RECT 523.950 1.950 526.050 2.400 ;
      LAYER metal3 ;
        RECT 523.950 52.950 526.050 55.050 ;
        RECT 524.400 4.050 525.600 52.950 ;
        RECT 517.950 1.950 520.050 4.050 ;
        RECT 523.950 1.950 526.050 4.050 ;
        RECT 518.400 -3.600 519.600 1.950 ;
    END
  END Yin[3]
  PIN Yin[2]
    PORT
      LAYER metal2 ;
        RECT 502.950 52.950 508.050 55.050 ;
        RECT 499.950 6.450 502.050 7.050 ;
        RECT 505.950 6.450 508.050 7.050 ;
        RECT 499.950 5.400 508.050 6.450 ;
        RECT 499.950 4.950 502.050 5.400 ;
        RECT 505.950 4.950 508.050 5.400 ;
      LAYER metal3 ;
        RECT 505.950 52.950 508.050 55.050 ;
        RECT 506.400 7.050 507.600 52.950 ;
        RECT 499.950 4.950 502.050 7.050 ;
        RECT 505.950 4.950 508.050 7.050 ;
        RECT 500.400 -3.600 501.600 4.950 ;
    END
  END Yin[2]
  PIN Yin[1]
    PORT
      LAYER metal2 ;
        RECT 433.950 25.950 439.050 28.050 ;
      LAYER metal3 ;
        RECT 436.950 25.950 439.050 28.050 ;
        RECT 437.400 -3.600 438.600 25.950 ;
    END
  END Yin[1]
  PIN Yin[0]
    PORT
      LAYER metal1 ;
        RECT 379.950 112.950 382.050 115.050 ;
        RECT 380.550 88.050 381.450 112.950 ;
        RECT 379.800 85.950 381.900 88.050 ;
      LAYER metal2 ;
        RECT 400.950 259.950 403.050 262.050 ;
        RECT 388.950 207.450 391.050 208.050 ;
        RECT 400.950 207.450 403.050 208.050 ;
        RECT 388.950 206.400 403.050 207.450 ;
        RECT 388.950 205.950 391.050 206.400 ;
        RECT 400.950 205.950 403.050 206.400 ;
        RECT 379.950 114.450 382.050 115.050 ;
        RECT 385.950 114.450 388.050 115.050 ;
        RECT 379.950 113.400 388.050 114.450 ;
        RECT 379.950 112.950 382.050 113.400 ;
        RECT 385.950 112.950 388.050 113.400 ;
        RECT 379.800 87.000 381.900 88.050 ;
        RECT 379.800 85.950 382.050 87.000 ;
        RECT 379.950 85.050 382.050 85.950 ;
        RECT 379.800 84.000 382.050 85.050 ;
        RECT 379.800 82.950 381.900 84.000 ;
        RECT 379.950 42.450 382.050 43.050 ;
        RECT 406.950 42.450 409.050 43.050 ;
        RECT 379.950 41.400 409.050 42.450 ;
        RECT 379.950 40.950 382.050 41.400 ;
        RECT 406.950 40.950 409.050 41.400 ;
      LAYER metal3 ;
        RECT 400.950 259.950 403.050 262.050 ;
        RECT 401.400 208.050 402.600 259.950 ;
        RECT 388.950 205.950 391.050 208.050 ;
        RECT 400.950 205.950 403.050 208.050 ;
        RECT 389.400 195.600 390.600 205.950 ;
        RECT 386.400 194.400 390.600 195.600 ;
        RECT 386.400 115.050 387.600 194.400 ;
        RECT 385.950 112.950 388.050 115.050 ;
        RECT 379.800 82.950 381.900 85.050 ;
        RECT 380.400 43.050 381.600 82.950 ;
        RECT 379.950 40.950 382.050 43.050 ;
        RECT 406.950 40.950 409.050 43.050 ;
        RECT 407.400 -2.400 408.600 40.950 ;
        RECT 404.400 -3.600 408.600 -2.400 ;
    END
  END Yin[0]
  PIN Yout[3]
    PORT
      LAYER metal2 ;
        RECT 649.950 19.950 652.050 22.050 ;
        RECT 650.400 15.450 651.450 19.950 ;
        RECT 715.950 15.450 718.050 16.050 ;
        RECT 650.400 14.400 718.050 15.450 ;
        RECT 715.950 13.950 718.050 14.400 ;
      LAYER metal3 ;
        RECT 715.950 13.950 718.050 16.050 ;
        RECT 716.400 -3.600 717.600 13.950 ;
    END
  END Yout[3]
  PIN Yout[2]
    PORT
      LAYER metal2 ;
        RECT 709.950 19.950 715.050 22.050 ;
      LAYER metal3 ;
        RECT 709.950 19.950 712.050 22.050 ;
        RECT 710.400 -3.600 711.600 19.950 ;
    END
  END Yout[2]
  PIN Yout[1]
    PORT
      LAYER metal2 ;
        RECT 688.950 19.950 694.050 22.050 ;
      LAYER metal3 ;
        RECT 688.950 19.950 691.050 22.050 ;
        RECT 689.400 -3.600 690.600 19.950 ;
    END
  END Yout[1]
  PIN Yout[0]
    PORT
      LAYER metal2 ;
        RECT 667.950 19.950 673.050 22.050 ;
      LAYER metal3 ;
        RECT 667.950 19.950 670.050 22.050 ;
        RECT 668.400 -3.600 669.600 19.950 ;
    END
  END Yout[0]
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 166.950 772.950 169.050 775.050 ;
        RECT 167.550 754.050 168.450 772.950 ;
        RECT 166.950 751.950 169.050 754.050 ;
      LAYER metal2 ;
        RECT 163.950 900.450 166.050 901.050 ;
        RECT 196.950 900.450 199.050 901.050 ;
        RECT 163.950 899.400 199.050 900.450 ;
        RECT 163.950 898.950 166.050 899.400 ;
        RECT 196.950 898.950 199.050 899.400 ;
        RECT 163.950 772.950 169.050 775.050 ;
        RECT 160.950 753.450 163.050 754.050 ;
        RECT 166.950 753.450 169.050 754.050 ;
        RECT 160.950 752.400 169.050 753.450 ;
        RECT 160.950 751.950 163.050 752.400 ;
        RECT 166.950 751.950 169.050 752.400 ;
        RECT 160.950 663.450 163.050 664.050 ;
        RECT 178.950 663.450 181.050 664.050 ;
        RECT 160.950 662.400 181.050 663.450 ;
        RECT 160.950 661.950 163.050 662.400 ;
        RECT 178.950 661.950 181.050 662.400 ;
        RECT 178.950 555.450 181.050 556.050 ;
        RECT 190.950 555.450 193.050 556.050 ;
        RECT 178.950 554.400 193.050 555.450 ;
        RECT 178.950 553.950 181.050 554.400 ;
        RECT 190.950 553.950 193.050 554.400 ;
        RECT 190.950 487.950 193.050 490.050 ;
        RECT 190.950 471.450 193.050 472.050 ;
        RECT 247.950 471.450 250.050 472.050 ;
        RECT 190.950 470.400 250.050 471.450 ;
        RECT 190.950 469.950 193.050 470.400 ;
        RECT 247.950 469.950 250.050 470.400 ;
        RECT 250.950 429.450 253.050 430.050 ;
        RECT 274.950 429.450 277.050 430.050 ;
        RECT 250.950 428.400 277.050 429.450 ;
        RECT 250.950 427.950 253.050 428.400 ;
        RECT 274.950 427.950 277.050 428.400 ;
        RECT 274.950 390.450 277.050 391.050 ;
        RECT 340.950 390.450 343.050 391.050 ;
        RECT 274.950 389.400 343.050 390.450 ;
        RECT 274.950 388.950 277.050 389.400 ;
        RECT 340.950 388.950 343.050 389.400 ;
        RECT 340.950 348.450 343.050 349.050 ;
        RECT 346.950 348.450 349.050 349.050 ;
        RECT 340.950 347.400 349.050 348.450 ;
        RECT 340.950 346.950 343.050 347.400 ;
        RECT 346.950 346.950 349.050 347.400 ;
        RECT 646.950 312.450 649.050 313.050 ;
        RECT 862.950 312.450 865.050 313.050 ;
        RECT 646.950 311.400 865.050 312.450 ;
        RECT 646.950 310.950 649.050 311.400 ;
        RECT 862.950 310.950 865.050 311.400 ;
        RECT 346.950 292.950 349.050 295.050 ;
        RECT 592.950 292.950 595.050 295.050 ;
        RECT 865.950 292.950 868.050 295.050 ;
        RECT 574.950 285.450 577.050 286.050 ;
        RECT 592.950 285.450 595.050 286.050 ;
        RECT 574.950 284.400 595.050 285.450 ;
        RECT 574.950 283.950 577.050 284.400 ;
        RECT 592.950 283.950 595.050 284.400 ;
        RECT 646.950 253.950 649.050 256.050 ;
        RECT 340.950 249.450 343.050 250.050 ;
        RECT 346.950 249.450 349.050 250.050 ;
        RECT 340.950 248.400 349.050 249.450 ;
        RECT 340.950 247.950 343.050 248.400 ;
        RECT 346.950 247.950 349.050 248.400 ;
        RECT 574.950 243.450 577.050 244.050 ;
        RECT 646.950 243.450 649.050 244.050 ;
        RECT 574.950 242.400 649.050 243.450 ;
        RECT 574.950 241.950 577.050 242.400 ;
        RECT 646.950 241.950 649.050 242.400 ;
        RECT 487.950 237.450 490.050 238.050 ;
        RECT 574.950 237.450 577.050 238.050 ;
        RECT 487.950 236.400 577.050 237.450 ;
        RECT 487.950 235.950 490.050 236.400 ;
        RECT 574.950 235.950 577.050 236.400 ;
        RECT 244.950 198.450 247.050 199.050 ;
        RECT 340.950 198.450 343.050 199.050 ;
        RECT 397.950 198.450 400.050 199.050 ;
        RECT 244.950 197.400 400.050 198.450 ;
        RECT 244.950 196.950 247.050 197.400 ;
        RECT 340.950 196.950 343.050 197.400 ;
        RECT 397.950 196.950 400.050 197.400 ;
        RECT 235.950 177.450 238.050 178.050 ;
        RECT 244.950 177.450 247.050 178.050 ;
        RECT 235.950 176.400 247.050 177.450 ;
        RECT 235.950 175.950 238.050 176.400 ;
        RECT 244.950 175.950 247.050 176.400 ;
        RECT 397.950 175.950 400.050 178.050 ;
        RECT 454.950 175.950 457.050 178.050 ;
        RECT 397.950 168.450 400.050 169.050 ;
        RECT 454.950 168.450 457.050 169.050 ;
        RECT 487.950 168.450 490.050 169.050 ;
        RECT 397.950 167.400 490.050 168.450 ;
        RECT 397.950 166.950 400.050 167.400 ;
        RECT 454.950 166.950 457.050 167.400 ;
        RECT 487.950 166.950 490.050 167.400 ;
      LAYER metal3 ;
        RECT 197.400 901.050 198.600 906.600 ;
        RECT 163.950 898.950 166.050 901.050 ;
        RECT 196.950 898.950 199.050 901.050 ;
        RECT 164.400 775.050 165.600 898.950 ;
        RECT 163.950 772.950 166.050 775.050 ;
        RECT 160.950 751.950 163.050 754.050 ;
        RECT 161.400 664.050 162.600 751.950 ;
        RECT 160.950 661.950 163.050 664.050 ;
        RECT 178.950 661.950 181.050 664.050 ;
        RECT 179.400 556.050 180.600 661.950 ;
        RECT 178.950 553.950 181.050 556.050 ;
        RECT 190.950 553.950 193.050 556.050 ;
        RECT 191.400 490.050 192.600 553.950 ;
        RECT 190.950 487.950 193.050 490.050 ;
        RECT 191.400 472.050 192.600 487.950 ;
        RECT 190.950 469.950 193.050 472.050 ;
        RECT 247.950 468.600 250.050 472.050 ;
        RECT 247.950 468.000 252.600 468.600 ;
        RECT 248.400 467.400 252.600 468.000 ;
        RECT 251.400 430.050 252.600 467.400 ;
        RECT 250.950 427.950 253.050 430.050 ;
        RECT 274.950 427.950 277.050 430.050 ;
        RECT 275.400 391.050 276.600 427.950 ;
        RECT 274.950 388.950 277.050 391.050 ;
        RECT 340.950 388.950 343.050 391.050 ;
        RECT 341.400 349.050 342.600 388.950 ;
        RECT 340.950 346.950 343.050 349.050 ;
        RECT 346.950 346.950 349.050 349.050 ;
        RECT 347.400 295.050 348.600 346.950 ;
        RECT 646.950 310.950 649.050 313.050 ;
        RECT 862.950 310.950 865.050 313.050 ;
        RECT 346.950 292.950 349.050 295.050 ;
        RECT 592.950 292.950 595.050 295.050 ;
        RECT 347.400 250.050 348.600 292.950 ;
        RECT 593.400 286.050 594.600 292.950 ;
        RECT 574.950 283.950 577.050 286.050 ;
        RECT 592.950 283.950 595.050 286.050 ;
        RECT 340.950 247.950 343.050 250.050 ;
        RECT 346.950 247.950 349.050 250.050 ;
        RECT 341.400 199.050 342.600 247.950 ;
        RECT 575.400 244.050 576.600 283.950 ;
        RECT 647.400 256.050 648.600 310.950 ;
        RECT 863.400 295.050 864.600 310.950 ;
        RECT 863.400 293.400 868.050 295.050 ;
        RECT 864.000 292.950 868.050 293.400 ;
        RECT 646.950 253.950 649.050 256.050 ;
        RECT 647.400 244.050 648.600 253.950 ;
        RECT 574.950 241.950 577.050 244.050 ;
        RECT 646.950 241.950 649.050 244.050 ;
        RECT 575.400 238.050 576.600 241.950 ;
        RECT 487.950 235.950 490.050 238.050 ;
        RECT 574.950 235.950 577.050 238.050 ;
        RECT 244.950 196.950 247.050 199.050 ;
        RECT 340.950 196.950 343.050 199.050 ;
        RECT 397.950 196.950 400.050 199.050 ;
        RECT 245.400 178.050 246.600 196.950 ;
        RECT 398.400 178.050 399.600 196.950 ;
        RECT 244.950 175.950 247.050 178.050 ;
        RECT 397.950 175.950 400.050 178.050 ;
        RECT 454.950 175.950 457.050 178.050 ;
        RECT 398.400 169.050 399.600 175.950 ;
        RECT 455.400 169.050 456.600 175.950 ;
        RECT 488.400 169.050 489.600 235.950 ;
        RECT 397.950 166.950 400.050 169.050 ;
        RECT 454.950 166.950 457.050 169.050 ;
        RECT 487.950 166.950 490.050 169.050 ;
    END
  END clk
  OBS
      LAYER metal1 ;
        RECT 16.200 888.000 18.000 896.400 ;
        RECT 40.500 891.600 42.300 896.400 ;
        RECT 40.500 890.400 45.600 891.600 ;
        RECT 14.700 886.800 18.000 888.000 ;
        RECT 14.700 883.050 15.600 886.800 ;
        RECT 44.400 883.050 45.600 890.400 ;
        RECT 64.200 888.000 66.000 896.400 ;
        RECT 76.950 892.950 79.050 895.050 ;
        RECT 62.700 886.800 66.000 888.000 ;
        RECT 46.800 885.450 51.000 886.050 ;
        RECT 46.800 883.950 51.450 885.450 ;
        RECT 13.950 880.950 16.050 883.050 ;
        RECT 14.700 868.800 15.600 880.950 ;
        RECT 17.100 880.050 18.900 881.850 ;
        RECT 19.950 880.950 22.050 883.050 ;
        RECT 16.950 877.950 19.050 880.050 ;
        RECT 20.100 879.150 21.900 880.950 ;
        RECT 23.100 880.050 24.900 881.850 ;
        RECT 35.100 880.050 36.900 881.850 ;
        RECT 37.950 880.950 40.050 883.050 ;
        RECT 22.950 877.950 25.050 880.050 ;
        RECT 34.950 877.950 37.050 880.050 ;
        RECT 38.100 879.150 39.900 880.950 ;
        RECT 41.100 880.050 42.900 881.850 ;
        RECT 43.950 880.950 46.050 883.050 ;
        RECT 40.950 877.950 43.050 880.050 ;
        RECT 44.400 873.600 45.600 880.950 ;
        RECT 35.400 872.700 43.200 873.600 ;
        RECT 14.700 867.900 21.300 868.800 ;
        RECT 14.700 867.600 15.600 867.900 ;
        RECT 13.800 861.600 15.600 867.600 ;
        RECT 19.800 867.600 21.300 867.900 ;
        RECT 19.800 861.600 21.600 867.600 ;
        RECT 35.400 861.600 37.200 872.700 ;
        RECT 41.400 861.600 43.200 872.700 ;
        RECT 44.400 861.600 46.200 873.600 ;
        RECT 50.550 865.050 51.450 883.950 ;
        RECT 62.700 883.050 63.600 886.800 ;
        RECT 61.950 880.950 64.050 883.050 ;
        RECT 62.700 868.800 63.600 880.950 ;
        RECT 65.100 880.050 66.900 881.850 ;
        RECT 67.950 880.950 70.050 883.050 ;
        RECT 64.950 877.950 67.050 880.050 ;
        RECT 68.100 879.150 69.900 880.950 ;
        RECT 71.100 880.050 72.900 881.850 ;
        RECT 70.950 877.950 73.050 880.050 ;
        RECT 77.550 871.050 78.450 892.950 ;
        RECT 88.200 888.000 90.000 896.400 ;
        RECT 109.800 890.400 111.600 896.400 ;
        RECT 86.700 886.800 90.000 888.000 ;
        RECT 110.400 888.300 111.600 890.400 ;
        RECT 112.800 891.300 114.600 896.400 ;
        RECT 118.800 891.300 120.600 896.400 ;
        RECT 112.800 889.950 120.600 891.300 ;
        RECT 133.800 890.400 135.600 896.400 ;
        RECT 134.400 888.300 135.600 890.400 ;
        RECT 136.800 891.300 138.600 896.400 ;
        RECT 142.800 891.300 144.600 896.400 ;
        RECT 136.800 889.950 144.600 891.300 ;
        RECT 158.400 893.400 160.200 896.400 ;
        RECT 176.400 893.400 178.200 896.400 ;
        RECT 110.400 887.250 114.150 888.300 ;
        RECT 134.400 887.250 138.150 888.300 ;
        RECT 81.000 885.450 85.050 886.050 ;
        RECT 80.550 883.950 85.050 885.450 ;
        RECT 76.950 868.950 79.050 871.050 ;
        RECT 62.700 867.900 69.300 868.800 ;
        RECT 62.700 867.600 63.600 867.900 ;
        RECT 49.950 862.950 52.050 865.050 ;
        RECT 61.800 861.600 63.600 867.600 ;
        RECT 67.800 867.600 69.300 867.900 ;
        RECT 67.800 861.600 69.600 867.600 ;
        RECT 80.550 865.050 81.450 883.950 ;
        RECT 86.700 883.050 87.600 886.800 ;
        RECT 103.950 883.950 106.050 886.050 ;
        RECT 85.950 880.950 88.050 883.050 ;
        RECT 86.700 868.800 87.600 880.950 ;
        RECT 89.100 880.050 90.900 881.850 ;
        RECT 91.950 880.950 94.050 883.050 ;
        RECT 88.950 877.950 91.050 880.050 ;
        RECT 92.100 879.150 93.900 880.950 ;
        RECT 95.100 880.050 96.900 881.850 ;
        RECT 100.950 880.950 103.050 883.050 ;
        RECT 94.950 877.950 97.050 880.050 ;
        RECT 101.550 871.050 102.450 880.950 ;
        RECT 100.950 868.950 103.050 871.050 ;
        RECT 86.700 867.900 93.300 868.800 ;
        RECT 86.700 867.600 87.600 867.900 ;
        RECT 79.800 862.950 81.900 865.050 ;
        RECT 85.800 861.600 87.600 867.600 ;
        RECT 91.800 867.600 93.300 867.900 ;
        RECT 91.800 861.600 93.600 867.600 ;
        RECT 104.550 865.050 105.450 883.950 ;
        RECT 112.950 883.050 114.150 887.250 ;
        RECT 136.950 883.050 138.150 887.250 ;
        RECT 110.100 880.050 111.900 881.850 ;
        RECT 112.950 880.950 115.050 883.050 ;
        RECT 109.950 877.950 112.050 880.050 ;
        RECT 113.850 867.600 115.050 880.950 ;
        RECT 116.100 880.050 117.900 881.850 ;
        RECT 118.950 880.950 121.050 883.050 ;
        RECT 127.950 880.950 130.050 883.050 ;
        RECT 115.950 877.950 118.050 880.050 ;
        RECT 119.100 879.150 120.900 880.950 ;
        RECT 128.550 871.050 129.450 880.950 ;
        RECT 134.100 880.050 135.900 881.850 ;
        RECT 136.950 880.950 139.050 883.050 ;
        RECT 133.950 877.950 136.050 880.050 ;
        RECT 127.950 868.950 130.050 871.050 ;
        RECT 137.850 867.600 139.050 880.950 ;
        RECT 140.100 880.050 141.900 881.850 ;
        RECT 142.950 880.950 145.050 883.050 ;
        RECT 154.950 880.950 157.050 883.050 ;
        RECT 139.950 877.950 142.050 880.050 ;
        RECT 143.100 879.150 144.900 880.950 ;
        RECT 155.100 879.150 156.900 880.950 ;
        RECT 158.400 880.050 159.600 893.400 ;
        RECT 172.950 880.950 175.050 883.050 ;
        RECT 157.950 874.950 160.050 880.050 ;
        RECT 173.100 879.150 174.900 880.950 ;
        RECT 176.400 880.050 177.600 893.400 ;
        RECT 196.500 891.600 198.300 896.400 ;
        RECT 196.500 890.400 201.600 891.600 ;
        RECT 200.400 883.050 201.600 890.400 ;
        RECT 218.400 889.200 220.200 896.400 ;
        RECT 236.400 891.300 238.200 896.400 ;
        RECT 242.400 891.300 244.200 896.400 ;
        RECT 236.400 889.950 244.200 891.300 ;
        RECT 245.400 890.400 247.200 896.400 ;
        RECT 218.400 888.300 222.600 889.200 ;
        RECT 245.400 888.300 246.600 890.400 ;
        RECT 265.800 889.200 267.600 896.400 ;
        RECT 221.400 883.050 222.600 888.300 ;
        RECT 242.850 887.250 246.600 888.300 ;
        RECT 263.400 888.300 267.600 889.200 ;
        RECT 283.500 890.400 285.300 896.400 ;
        RECT 289.800 893.400 291.600 896.400 ;
        RECT 242.850 883.050 244.050 887.250 ;
        RECT 263.400 883.050 264.600 888.300 ;
        RECT 283.500 883.050 284.700 890.400 ;
        RECT 290.400 889.500 291.600 893.400 ;
        RECT 285.600 888.600 291.600 889.500 ;
        RECT 302.400 893.400 304.200 896.400 ;
        RECT 302.400 889.500 303.600 893.400 ;
        RECT 308.700 890.400 310.500 896.400 ;
        RECT 302.400 888.600 308.400 889.500 ;
        RECT 285.600 887.700 287.850 888.600 ;
        RECT 191.100 880.050 192.900 881.850 ;
        RECT 193.950 880.950 196.050 883.050 ;
        RECT 175.950 874.950 178.050 880.050 ;
        RECT 190.950 877.950 193.050 880.050 ;
        RECT 194.100 879.150 195.900 880.950 ;
        RECT 197.100 880.050 198.900 881.850 ;
        RECT 199.950 880.950 202.050 883.050 ;
        RECT 196.950 877.950 199.050 880.050 ;
        RECT 158.400 867.600 159.600 874.950 ;
        RECT 176.400 867.600 177.600 874.950 ;
        RECT 200.400 873.600 201.600 880.950 ;
        RECT 218.100 880.050 219.900 881.850 ;
        RECT 220.950 880.950 223.050 883.050 ;
        RECT 217.950 877.950 220.050 880.050 ;
        RECT 191.400 872.700 199.200 873.600 ;
        RECT 103.950 862.950 106.050 865.050 ;
        RECT 113.400 861.600 115.200 867.600 ;
        RECT 137.400 861.600 139.200 867.600 ;
        RECT 158.400 861.600 160.200 867.600 ;
        RECT 176.400 861.600 178.200 867.600 ;
        RECT 191.400 861.600 193.200 872.700 ;
        RECT 197.400 861.600 199.200 872.700 ;
        RECT 200.400 861.600 202.200 873.600 ;
        RECT 221.400 867.600 222.600 880.950 ;
        RECT 224.100 880.050 225.900 881.850 ;
        RECT 235.950 880.950 238.050 883.050 ;
        RECT 223.950 877.950 226.050 880.050 ;
        RECT 236.100 879.150 237.900 880.950 ;
        RECT 239.100 880.050 240.900 881.850 ;
        RECT 241.950 880.950 244.050 883.050 ;
        RECT 238.950 877.950 241.050 880.050 ;
        RECT 241.950 867.600 243.150 880.950 ;
        RECT 245.100 880.050 246.900 881.850 ;
        RECT 260.100 880.050 261.900 881.850 ;
        RECT 262.950 880.950 265.050 883.050 ;
        RECT 244.950 877.950 247.050 880.050 ;
        RECT 259.950 877.950 262.050 880.050 ;
        RECT 263.400 867.600 264.600 880.950 ;
        RECT 266.100 880.050 267.900 881.850 ;
        RECT 283.500 880.950 286.050 883.050 ;
        RECT 265.950 877.950 268.050 880.050 ;
        RECT 283.500 873.600 284.700 880.950 ;
        RECT 286.950 876.300 287.850 887.700 ;
        RECT 306.150 887.700 308.400 888.600 ;
        RECT 289.950 880.950 292.050 883.050 ;
        RECT 301.950 880.950 304.050 883.050 ;
        RECT 290.100 879.150 291.900 880.950 ;
        RECT 302.100 879.150 303.900 880.950 ;
        RECT 285.600 875.400 287.850 876.300 ;
        RECT 306.150 876.300 307.050 887.700 ;
        RECT 309.300 883.050 310.500 890.400 ;
        RECT 326.400 889.200 328.200 896.400 ;
        RECT 326.400 888.300 330.600 889.200 ;
        RECT 329.400 883.050 330.600 888.300 ;
        RECT 344.400 888.600 346.200 896.400 ;
        RECT 351.900 892.200 353.700 896.400 ;
        RECT 351.900 890.400 354.600 892.200 ;
        RECT 350.100 888.600 351.900 889.500 ;
        RECT 344.400 887.700 351.900 888.600 ;
        RECT 344.100 883.050 345.900 884.850 ;
        RECT 307.950 880.950 310.500 883.050 ;
        RECT 306.150 875.400 308.400 876.300 ;
        RECT 285.600 874.500 291.600 875.400 ;
        RECT 220.800 861.600 222.600 867.600 ;
        RECT 241.800 861.600 243.600 867.600 ;
        RECT 263.400 861.600 265.200 867.600 ;
        RECT 283.500 861.600 285.300 873.600 ;
        RECT 290.400 867.600 291.600 874.500 ;
        RECT 289.800 861.600 291.600 867.600 ;
        RECT 302.400 874.500 308.400 875.400 ;
        RECT 302.400 867.600 303.600 874.500 ;
        RECT 309.300 873.600 310.500 880.950 ;
        RECT 326.100 880.050 327.900 881.850 ;
        RECT 328.950 880.950 331.050 883.050 ;
        RECT 325.950 877.950 328.050 880.050 ;
        RECT 302.400 861.600 304.200 867.600 ;
        RECT 308.700 861.600 310.500 873.600 ;
        RECT 329.400 867.600 330.600 880.950 ;
        RECT 332.100 880.050 333.900 881.850 ;
        RECT 343.950 880.950 346.050 883.050 ;
        RECT 331.950 877.950 334.050 880.050 ;
        RECT 328.800 861.600 330.600 867.600 ;
        RECT 347.400 867.600 348.300 887.700 ;
        RECT 353.700 883.050 354.600 890.400 ;
        RECT 371.400 889.200 373.200 896.400 ;
        RECT 394.800 889.200 396.600 896.400 ;
        RECT 415.800 893.400 417.600 896.400 ;
        RECT 371.400 888.300 375.600 889.200 ;
        RECT 374.400 883.050 375.600 888.300 ;
        RECT 392.400 888.300 396.600 889.200 ;
        RECT 382.950 883.950 385.050 886.050 ;
        RECT 349.950 880.950 352.050 883.050 ;
        RECT 352.950 880.950 355.050 883.050 ;
        RECT 350.100 879.150 351.900 880.950 ;
        RECT 353.700 873.600 354.600 880.950 ;
        RECT 371.100 880.050 372.900 881.850 ;
        RECT 373.950 880.950 376.050 883.050 ;
        RECT 370.950 877.950 373.050 880.050 ;
        RECT 347.400 861.600 349.200 867.600 ;
        RECT 353.700 861.600 355.500 873.600 ;
        RECT 374.400 867.600 375.600 880.950 ;
        RECT 377.100 880.050 378.900 881.850 ;
        RECT 376.950 877.950 379.050 880.050 ;
        RECT 383.550 877.050 384.450 883.950 ;
        RECT 392.400 883.050 393.600 888.300 ;
        RECT 400.950 886.950 403.050 889.050 ;
        RECT 389.100 880.050 390.900 881.850 ;
        RECT 391.950 880.950 394.050 883.050 ;
        RECT 388.950 877.950 391.050 880.050 ;
        RECT 382.950 874.950 385.050 877.050 ;
        RECT 373.800 861.600 375.600 867.600 ;
        RECT 392.400 867.600 393.600 880.950 ;
        RECT 395.100 880.050 396.900 881.850 ;
        RECT 394.950 877.950 397.050 880.050 ;
        RECT 392.400 861.600 394.200 867.600 ;
        RECT 401.550 865.050 402.450 886.950 ;
        RECT 406.950 883.950 409.050 886.050 ;
        RECT 412.950 883.950 415.050 886.050 ;
        RECT 407.550 865.050 408.450 883.950 ;
        RECT 413.100 882.150 414.900 883.950 ;
        RECT 416.400 883.050 417.300 893.400 ;
        RECT 436.800 889.200 438.600 896.400 ;
        RECT 434.400 888.300 438.600 889.200 ;
        RECT 452.400 893.400 454.200 896.400 ;
        RECT 452.400 889.500 453.600 893.400 ;
        RECT 458.700 890.400 460.500 896.400 ;
        RECT 477.300 892.200 479.100 896.400 ;
        RECT 452.400 888.600 458.400 889.500 ;
        RECT 418.950 883.950 421.050 886.050 ;
        RECT 415.950 880.950 418.050 883.050 ;
        RECT 419.100 882.150 420.900 883.950 ;
        RECT 434.400 883.050 435.600 888.300 ;
        RECT 456.150 887.700 458.400 888.600 ;
        RECT 416.400 873.600 417.300 880.950 ;
        RECT 431.100 880.050 432.900 881.850 ;
        RECT 433.950 880.950 436.050 883.050 ;
        RECT 430.950 877.950 433.050 880.050 ;
        RECT 413.700 872.400 417.300 873.600 ;
        RECT 400.950 862.950 403.050 865.050 ;
        RECT 406.950 862.950 409.050 865.050 ;
        RECT 413.700 861.600 415.500 872.400 ;
        RECT 434.400 867.600 435.600 880.950 ;
        RECT 437.100 880.050 438.900 881.850 ;
        RECT 451.950 880.950 454.050 883.050 ;
        RECT 436.950 877.950 439.050 880.050 ;
        RECT 452.100 879.150 453.900 880.950 ;
        RECT 456.150 876.300 457.050 887.700 ;
        RECT 459.300 883.050 460.500 890.400 ;
        RECT 476.400 890.400 479.100 892.200 ;
        RECT 476.400 883.050 477.300 890.400 ;
        RECT 479.100 888.600 480.900 889.500 ;
        RECT 484.800 888.600 486.600 896.400 ;
        RECT 503.700 891.600 505.500 896.400 ;
        RECT 479.100 887.700 486.600 888.600 ;
        RECT 500.400 890.400 505.500 891.600 ;
        RECT 457.950 880.950 460.500 883.050 ;
        RECT 475.950 880.950 478.050 883.050 ;
        RECT 478.950 880.950 481.050 883.050 ;
        RECT 456.150 875.400 458.400 876.300 ;
        RECT 452.400 874.500 458.400 875.400 ;
        RECT 452.400 867.600 453.600 874.500 ;
        RECT 459.300 873.600 460.500 880.950 ;
        RECT 476.400 873.600 477.300 880.950 ;
        RECT 479.100 879.150 480.900 880.950 ;
        RECT 434.400 861.600 436.200 867.600 ;
        RECT 452.400 861.600 454.200 867.600 ;
        RECT 458.700 861.600 460.500 873.600 ;
        RECT 475.500 861.600 477.300 873.600 ;
        RECT 482.700 867.600 483.600 887.700 ;
        RECT 485.100 883.050 486.900 884.850 ;
        RECT 500.400 883.050 501.600 890.400 ;
        RECT 514.950 889.950 517.050 892.050 ;
        RECT 484.950 880.950 487.050 883.050 ;
        RECT 499.950 880.950 502.050 883.050 ;
        RECT 500.400 873.600 501.600 880.950 ;
        RECT 503.100 880.050 504.900 881.850 ;
        RECT 505.950 880.950 508.050 883.050 ;
        RECT 502.950 877.950 505.050 880.050 ;
        RECT 506.100 879.150 507.900 880.950 ;
        RECT 509.100 880.050 510.900 881.850 ;
        RECT 508.950 877.950 511.050 880.050 ;
        RECT 515.550 877.050 516.450 889.950 ;
        RECT 526.200 888.000 528.000 896.400 ;
        RECT 538.950 889.950 541.050 892.050 ;
        RECT 524.700 886.800 528.000 888.000 ;
        RECT 524.700 883.050 525.600 886.800 ;
        RECT 523.950 880.950 526.050 883.050 ;
        RECT 514.950 874.950 517.050 877.050 ;
        RECT 481.800 861.600 483.600 867.600 ;
        RECT 499.800 861.600 501.600 873.600 ;
        RECT 502.800 872.700 510.600 873.600 ;
        RECT 502.800 861.600 504.600 872.700 ;
        RECT 508.800 861.600 510.600 872.700 ;
        RECT 524.700 868.800 525.600 880.950 ;
        RECT 527.100 880.050 528.900 881.850 ;
        RECT 529.950 880.950 532.050 883.050 ;
        RECT 526.950 877.950 529.050 880.050 ;
        RECT 530.100 879.150 531.900 880.950 ;
        RECT 533.100 880.050 534.900 881.850 ;
        RECT 532.950 877.950 535.050 880.050 ;
        RECT 539.550 877.050 540.450 889.950 ;
        RECT 550.800 889.200 552.600 896.400 ;
        RECT 548.400 888.300 552.600 889.200 ;
        RECT 548.400 883.050 549.600 888.300 ;
        RECT 571.200 888.000 573.000 896.400 ;
        RECT 593.400 889.200 595.200 896.400 ;
        RECT 611.400 893.400 613.200 896.400 ;
        RECT 611.400 889.500 612.600 893.400 ;
        RECT 617.700 890.400 619.500 896.400 ;
        RECT 593.400 888.300 597.600 889.200 ;
        RECT 611.400 888.600 617.400 889.500 ;
        RECT 569.700 886.800 573.000 888.000 ;
        RECT 569.700 883.050 570.600 886.800 ;
        RECT 596.400 883.050 597.600 888.300 ;
        RECT 615.150 887.700 617.400 888.600 ;
        RECT 545.100 880.050 546.900 881.850 ;
        RECT 547.950 880.950 550.050 883.050 ;
        RECT 544.950 877.950 547.050 880.050 ;
        RECT 538.950 874.950 541.050 877.050 ;
        RECT 524.700 867.900 531.300 868.800 ;
        RECT 524.700 867.600 525.600 867.900 ;
        RECT 523.800 861.600 525.600 867.600 ;
        RECT 529.800 867.600 531.300 867.900 ;
        RECT 529.800 861.600 531.600 867.600 ;
        RECT 539.550 865.050 540.450 874.950 ;
        RECT 535.800 863.550 540.450 865.050 ;
        RECT 548.400 867.600 549.600 880.950 ;
        RECT 551.100 880.050 552.900 881.850 ;
        RECT 568.950 880.950 571.050 883.050 ;
        RECT 550.950 877.950 553.050 880.050 ;
        RECT 569.700 868.800 570.600 880.950 ;
        RECT 572.100 880.050 573.900 881.850 ;
        RECT 574.950 880.950 577.050 883.050 ;
        RECT 571.950 877.950 574.050 880.050 ;
        RECT 575.100 879.150 576.900 880.950 ;
        RECT 578.100 880.050 579.900 881.850 ;
        RECT 593.100 880.050 594.900 881.850 ;
        RECT 595.950 880.950 598.050 883.050 ;
        RECT 577.950 877.950 580.050 880.050 ;
        RECT 592.950 877.950 595.050 880.050 ;
        RECT 580.950 874.950 583.050 877.050 ;
        RECT 569.700 867.900 576.300 868.800 ;
        RECT 569.700 867.600 570.600 867.900 ;
        RECT 535.800 862.950 540.000 863.550 ;
        RECT 548.400 861.600 550.200 867.600 ;
        RECT 568.800 861.600 570.600 867.600 ;
        RECT 574.800 867.600 576.300 867.900 ;
        RECT 574.800 861.600 576.600 867.600 ;
        RECT 581.550 865.050 582.450 874.950 ;
        RECT 596.400 867.600 597.600 880.950 ;
        RECT 599.100 880.050 600.900 881.850 ;
        RECT 610.950 880.950 613.050 883.050 ;
        RECT 598.950 877.950 601.050 880.050 ;
        RECT 611.100 879.150 612.900 880.950 ;
        RECT 615.150 876.300 616.050 887.700 ;
        RECT 618.300 883.050 619.500 890.400 ;
        RECT 642.000 890.400 643.800 896.400 ;
        RECT 661.500 890.400 663.300 896.400 ;
        RECT 667.800 893.400 669.600 896.400 ;
        RECT 682.800 893.400 684.600 896.400 ;
        RECT 635.100 883.050 636.900 884.850 ;
        RECT 637.950 883.950 640.050 886.050 ;
        RECT 616.950 880.950 619.500 883.050 ;
        RECT 634.950 880.950 637.050 883.050 ;
        RECT 638.100 882.150 639.900 883.950 ;
        RECT 642.000 883.050 643.050 890.400 ;
        RECT 643.950 883.950 646.050 886.050 ;
        RECT 640.950 880.950 643.050 883.050 ;
        RECT 644.100 882.150 645.900 883.950 ;
        RECT 647.100 883.050 648.900 884.850 ;
        RECT 661.500 883.050 662.700 890.400 ;
        RECT 668.400 889.500 669.600 893.400 ;
        RECT 663.600 888.600 669.600 889.500 ;
        RECT 663.600 887.700 665.850 888.600 ;
        RECT 646.950 880.950 649.050 883.050 ;
        RECT 661.500 880.950 664.050 883.050 ;
        RECT 615.150 875.400 617.400 876.300 ;
        RECT 580.950 862.950 583.050 865.050 ;
        RECT 595.800 861.600 597.600 867.600 ;
        RECT 611.400 874.500 617.400 875.400 ;
        RECT 611.400 867.600 612.600 874.500 ;
        RECT 618.300 873.600 619.500 880.950 ;
        RECT 642.000 875.400 642.900 880.950 ;
        RECT 637.800 874.500 642.900 875.400 ;
        RECT 611.400 861.600 613.200 867.600 ;
        RECT 617.700 861.600 619.500 873.600 ;
        RECT 634.800 862.500 636.600 873.600 ;
        RECT 637.800 863.400 639.600 874.500 ;
        RECT 661.500 873.600 662.700 880.950 ;
        RECT 664.950 876.300 665.850 887.700 ;
        RECT 667.950 880.950 670.050 883.050 ;
        RECT 668.100 879.150 669.900 880.950 ;
        RECT 683.400 880.050 684.600 893.400 ;
        RECT 698.400 893.400 700.200 896.400 ;
        RECT 698.400 889.500 699.600 893.400 ;
        RECT 704.700 890.400 706.500 896.400 ;
        RECT 723.300 892.200 725.100 896.400 ;
        RECT 698.400 888.600 704.400 889.500 ;
        RECT 702.150 887.700 704.400 888.600 ;
        RECT 685.950 880.950 688.050 883.050 ;
        RECT 697.950 880.950 700.050 883.050 ;
        RECT 663.600 875.400 665.850 876.300 ;
        RECT 663.600 874.500 669.600 875.400 ;
        RECT 682.950 874.950 685.050 880.050 ;
        RECT 686.100 879.150 687.900 880.950 ;
        RECT 698.100 879.150 699.900 880.950 ;
        RECT 702.150 876.300 703.050 887.700 ;
        RECT 705.300 883.050 706.500 890.400 ;
        RECT 709.950 889.950 712.050 892.050 ;
        RECT 722.400 890.400 725.100 892.200 ;
        RECT 703.950 880.950 706.500 883.050 ;
        RECT 702.150 875.400 704.400 876.300 ;
        RECT 640.800 872.400 648.600 873.300 ;
        RECT 640.800 862.500 642.600 872.400 ;
        RECT 634.800 861.600 642.600 862.500 ;
        RECT 646.800 861.600 648.600 872.400 ;
        RECT 661.500 861.600 663.300 873.600 ;
        RECT 668.400 867.600 669.600 874.500 ;
        RECT 683.400 867.600 684.600 874.950 ;
        RECT 667.800 861.600 669.600 867.600 ;
        RECT 682.800 861.600 684.600 867.600 ;
        RECT 698.400 874.500 704.400 875.400 ;
        RECT 698.400 867.600 699.600 874.500 ;
        RECT 705.300 873.600 706.500 880.950 ;
        RECT 698.400 861.600 700.200 867.600 ;
        RECT 704.700 861.600 706.500 873.600 ;
        RECT 710.550 868.050 711.450 889.950 ;
        RECT 722.400 883.050 723.300 890.400 ;
        RECT 725.100 888.600 726.900 889.500 ;
        RECT 730.800 888.600 732.600 896.400 ;
        RECT 748.200 890.400 750.000 896.400 ;
        RECT 766.950 892.950 769.050 895.050 ;
        RECT 725.100 887.700 732.600 888.600 ;
        RECT 721.950 880.950 724.050 883.050 ;
        RECT 724.950 880.950 727.050 883.050 ;
        RECT 722.400 873.600 723.300 880.950 ;
        RECT 725.100 879.150 726.900 880.950 ;
        RECT 709.800 865.950 711.900 868.050 ;
        RECT 721.500 861.600 723.300 873.600 ;
        RECT 728.700 867.600 729.600 887.700 ;
        RECT 731.100 883.050 732.900 884.850 ;
        RECT 743.100 883.050 744.900 884.850 ;
        RECT 745.950 883.950 748.050 886.050 ;
        RECT 730.950 880.950 733.050 883.050 ;
        RECT 742.950 880.950 745.050 883.050 ;
        RECT 746.100 882.150 747.900 883.950 ;
        RECT 748.950 883.050 750.000 890.400 ;
        RECT 767.550 889.050 768.450 892.950 ;
        RECT 766.950 886.950 769.050 889.050 ;
        RECT 770.400 888.600 772.200 896.400 ;
        RECT 777.900 892.200 779.700 896.400 ;
        RECT 777.900 890.400 780.600 892.200 ;
        RECT 776.100 888.600 777.900 889.500 ;
        RECT 770.400 887.700 777.900 888.600 ;
        RECT 751.950 883.950 754.050 886.050 ;
        RECT 748.950 880.950 751.050 883.050 ;
        RECT 752.100 882.150 753.900 883.950 ;
        RECT 755.100 883.050 756.900 884.850 ;
        RECT 770.100 883.050 771.900 884.850 ;
        RECT 754.950 880.950 757.050 883.050 ;
        RECT 769.950 880.950 772.050 883.050 ;
        RECT 749.100 875.400 750.000 880.950 ;
        RECT 749.100 874.500 754.200 875.400 ;
        RECT 727.800 861.600 729.600 867.600 ;
        RECT 743.400 872.400 751.200 873.300 ;
        RECT 743.400 861.600 745.200 872.400 ;
        RECT 749.400 862.500 751.200 872.400 ;
        RECT 752.400 863.400 754.200 874.500 ;
        RECT 755.400 862.500 757.200 873.600 ;
        RECT 749.400 861.600 757.200 862.500 ;
        RECT 773.400 867.600 774.300 887.700 ;
        RECT 779.700 883.050 780.600 890.400 ;
        RECT 804.000 890.400 805.800 896.400 ;
        RECT 797.100 883.050 798.900 884.850 ;
        RECT 799.950 883.950 802.050 886.050 ;
        RECT 775.950 880.950 778.050 883.050 ;
        RECT 778.950 880.950 781.050 883.050 ;
        RECT 796.950 880.950 799.050 883.050 ;
        RECT 800.100 882.150 801.900 883.950 ;
        RECT 804.000 883.050 805.050 890.400 ;
        RECT 826.800 889.200 828.600 896.400 ;
        RECT 842.400 891.300 844.200 896.400 ;
        RECT 848.400 891.300 850.200 896.400 ;
        RECT 842.400 889.950 850.200 891.300 ;
        RECT 851.400 890.400 853.200 896.400 ;
        RECT 869.400 893.400 871.200 896.400 ;
        RECT 887.400 893.400 889.200 896.400 ;
        RECT 824.400 888.300 828.600 889.200 ;
        RECT 851.400 888.300 852.600 890.400 ;
        RECT 805.950 883.950 808.050 886.050 ;
        RECT 802.950 880.950 805.050 883.050 ;
        RECT 806.100 882.150 807.900 883.950 ;
        RECT 809.100 883.050 810.900 884.850 ;
        RECT 824.400 883.050 825.600 888.300 ;
        RECT 848.850 887.250 852.600 888.300 ;
        RECT 848.850 883.050 850.050 887.250 ;
        RECT 808.950 880.950 811.050 883.050 ;
        RECT 776.100 879.150 777.900 880.950 ;
        RECT 779.700 873.600 780.600 880.950 ;
        RECT 804.000 875.400 804.900 880.950 ;
        RECT 821.100 880.050 822.900 881.850 ;
        RECT 823.950 880.950 826.050 883.050 ;
        RECT 820.950 877.950 823.050 880.050 ;
        RECT 799.800 874.500 804.900 875.400 ;
        RECT 773.400 861.600 775.200 867.600 ;
        RECT 779.700 861.600 781.500 873.600 ;
        RECT 796.800 862.500 798.600 873.600 ;
        RECT 799.800 863.400 801.600 874.500 ;
        RECT 802.800 872.400 810.600 873.300 ;
        RECT 802.800 862.500 804.600 872.400 ;
        RECT 796.800 861.600 804.600 862.500 ;
        RECT 808.800 861.600 810.600 872.400 ;
        RECT 811.800 871.950 813.900 874.050 ;
        RECT 812.550 868.050 813.450 871.950 ;
        RECT 811.950 865.950 814.050 868.050 ;
        RECT 824.400 867.600 825.600 880.950 ;
        RECT 827.100 880.050 828.900 881.850 ;
        RECT 841.950 880.950 844.050 883.050 ;
        RECT 826.950 877.950 829.050 880.050 ;
        RECT 842.100 879.150 843.900 880.950 ;
        RECT 845.100 880.050 846.900 881.850 ;
        RECT 847.950 880.950 850.050 883.050 ;
        RECT 844.950 877.950 847.050 880.050 ;
        RECT 847.950 867.600 849.150 880.950 ;
        RECT 851.100 880.050 852.900 881.850 ;
        RECT 865.950 880.950 868.050 883.050 ;
        RECT 850.950 877.950 853.050 880.050 ;
        RECT 866.100 879.150 867.900 880.950 ;
        RECT 869.400 880.050 870.600 893.400 ;
        RECT 888.300 889.200 889.200 893.400 ;
        RECT 893.400 890.400 895.200 896.400 ;
        RECT 888.300 888.300 891.600 889.200 ;
        RECT 889.800 887.400 891.600 888.300 ;
        RECT 884.100 880.050 885.900 881.850 ;
        RECT 886.950 880.950 889.050 883.050 ;
        RECT 868.950 874.950 871.050 880.050 ;
        RECT 883.950 877.950 886.050 880.050 ;
        RECT 887.100 879.150 888.900 880.950 ;
        RECT 890.700 876.900 891.600 887.400 ;
        RECT 894.000 883.050 895.050 890.400 ;
        RECT 889.800 876.300 891.600 876.900 ;
        RECT 884.400 875.100 891.600 876.300 ;
        RECT 892.950 880.950 895.050 883.050 ;
        RECT 869.400 867.600 870.600 874.950 ;
        RECT 884.400 873.600 885.600 875.100 ;
        RECT 892.950 873.600 894.300 880.950 ;
        RECT 824.400 861.600 826.200 867.600 ;
        RECT 847.800 861.600 849.600 867.600 ;
        RECT 869.400 861.600 871.200 867.600 ;
        RECT 884.400 861.600 886.200 873.600 ;
        RECT 891.900 872.100 894.300 873.600 ;
        RECT 891.900 861.600 893.700 872.100 ;
        RECT 13.800 851.400 15.600 857.400 ;
        RECT 14.700 851.100 15.600 851.400 ;
        RECT 19.800 851.400 21.600 857.400 ;
        RECT 19.800 851.100 21.300 851.400 ;
        RECT 14.700 850.200 21.300 851.100 ;
        RECT 14.700 838.050 15.600 850.200 ;
        RECT 35.400 846.300 37.200 857.400 ;
        RECT 41.400 846.300 43.200 857.400 ;
        RECT 35.400 845.400 43.200 846.300 ;
        RECT 44.400 845.400 46.200 857.400 ;
        RECT 61.800 851.400 63.600 857.400 ;
        RECT 62.700 851.100 63.600 851.400 ;
        RECT 67.800 851.400 69.600 857.400 ;
        RECT 67.800 851.100 69.300 851.400 ;
        RECT 62.700 850.200 69.300 851.100 ;
        RECT 16.950 838.950 19.050 841.050 ;
        RECT 13.950 835.950 16.050 838.050 ;
        RECT 17.100 837.150 18.900 838.950 ;
        RECT 20.100 838.050 21.900 839.850 ;
        RECT 22.950 838.950 25.050 841.050 ;
        RECT 34.950 838.950 37.050 841.050 ;
        RECT 19.950 835.950 22.050 838.050 ;
        RECT 23.100 837.150 24.900 838.950 ;
        RECT 35.100 837.150 36.900 838.950 ;
        RECT 38.100 838.050 39.900 839.850 ;
        RECT 40.950 838.950 43.050 841.050 ;
        RECT 37.950 835.950 40.050 838.050 ;
        RECT 41.100 837.150 42.900 838.950 ;
        RECT 44.400 838.050 45.600 845.400 ;
        RECT 62.700 838.050 63.600 850.200 ;
        RECT 83.400 846.300 85.200 857.400 ;
        RECT 89.400 846.300 91.200 857.400 ;
        RECT 83.400 845.400 91.200 846.300 ;
        RECT 92.400 845.400 94.200 857.400 ;
        RECT 109.800 845.400 111.600 857.400 ;
        RECT 112.800 846.300 114.600 857.400 ;
        RECT 118.800 846.300 120.600 857.400 ;
        RECT 133.800 851.400 135.600 857.400 ;
        RECT 154.800 851.400 156.600 857.400 ;
        RECT 179.400 851.400 181.200 857.400 ;
        RECT 112.800 845.400 120.600 846.300 ;
        RECT 64.950 838.950 67.050 841.050 ;
        RECT 43.950 835.950 46.050 838.050 ;
        RECT 61.950 835.950 64.050 838.050 ;
        RECT 65.100 837.150 66.900 838.950 ;
        RECT 68.100 838.050 69.900 839.850 ;
        RECT 70.950 838.950 73.050 841.050 ;
        RECT 82.950 838.950 85.050 841.050 ;
        RECT 67.950 835.950 70.050 838.050 ;
        RECT 71.100 837.150 72.900 838.950 ;
        RECT 83.100 837.150 84.900 838.950 ;
        RECT 86.100 838.050 87.900 839.850 ;
        RECT 88.950 838.950 91.050 841.050 ;
        RECT 85.950 835.950 88.050 838.050 ;
        RECT 89.100 837.150 90.900 838.950 ;
        RECT 92.400 838.050 93.600 845.400 ;
        RECT 97.950 841.950 100.050 844.050 ;
        RECT 91.950 835.950 94.050 838.050 ;
        RECT 14.700 832.200 15.600 835.950 ;
        RECT 14.700 831.000 18.000 832.200 ;
        RECT 16.200 822.600 18.000 831.000 ;
        RECT 44.400 828.600 45.600 835.950 ;
        RECT 62.700 832.200 63.600 835.950 ;
        RECT 62.700 831.000 66.000 832.200 ;
        RECT 40.500 827.400 45.600 828.600 ;
        RECT 40.500 822.600 42.300 827.400 ;
        RECT 64.200 822.600 66.000 831.000 ;
        RECT 92.400 828.600 93.600 835.950 ;
        RECT 88.500 827.400 93.600 828.600 ;
        RECT 88.500 822.600 90.300 827.400 ;
        RECT 98.550 826.050 99.450 841.950 ;
        RECT 110.400 838.050 111.600 845.400 ;
        RECT 134.400 844.050 135.600 851.400 ;
        RECT 124.950 841.950 127.050 844.050 ;
        RECT 112.950 838.950 115.050 841.050 ;
        RECT 109.950 835.950 112.050 838.050 ;
        RECT 113.100 837.150 114.900 838.950 ;
        RECT 116.100 838.050 117.900 839.850 ;
        RECT 118.950 838.950 121.050 841.050 ;
        RECT 115.950 835.950 118.050 838.050 ;
        RECT 119.100 837.150 120.900 838.950 ;
        RECT 110.400 828.600 111.600 835.950 ;
        RECT 125.550 829.050 126.450 841.950 ;
        RECT 133.950 838.950 136.050 844.050 ;
        RECT 110.400 827.400 115.500 828.600 ;
        RECT 97.950 823.950 100.050 826.050 ;
        RECT 113.700 822.600 115.500 827.400 ;
        RECT 124.950 826.950 127.050 829.050 ;
        RECT 134.400 825.600 135.600 838.950 ;
        RECT 137.100 838.050 138.900 839.850 ;
        RECT 149.100 838.050 150.900 839.850 ;
        RECT 151.950 838.950 154.050 841.050 ;
        RECT 136.950 835.950 139.050 838.050 ;
        RECT 148.950 835.950 151.050 838.050 ;
        RECT 152.100 837.150 153.900 838.950 ;
        RECT 154.950 838.050 156.150 851.400 ;
        RECT 157.950 838.950 160.050 841.050 ;
        RECT 175.950 838.950 178.050 841.050 ;
        RECT 154.950 835.950 157.050 838.050 ;
        RECT 158.100 837.150 159.900 838.950 ;
        RECT 176.100 837.150 177.900 838.950 ;
        RECT 179.850 838.050 181.050 851.400 ;
        RECT 202.500 846.600 204.300 857.400 ;
        RECT 205.950 850.950 208.050 853.050 ;
        RECT 200.700 845.400 204.300 846.600 ;
        RECT 181.950 838.950 184.050 841.050 ;
        RECT 155.850 831.750 157.050 835.950 ;
        RECT 178.950 835.950 181.050 838.050 ;
        RECT 182.100 837.150 183.900 838.950 ;
        RECT 185.100 838.050 186.900 839.850 ;
        RECT 200.700 838.050 201.600 845.400 ;
        RECT 206.550 841.050 207.450 850.950 ;
        RECT 223.500 846.600 225.300 857.400 ;
        RECT 221.700 845.400 225.300 846.600 ;
        RECT 242.400 851.400 244.200 857.400 ;
        RECT 250.950 853.950 253.050 856.050 ;
        RECT 205.950 838.950 208.050 841.050 ;
        RECT 221.700 838.050 222.600 845.400 ;
        RECT 238.950 838.950 241.050 841.050 ;
        RECT 184.950 835.950 187.050 838.050 ;
        RECT 178.950 831.750 180.150 835.950 ;
        RECT 197.100 835.050 198.900 836.850 ;
        RECT 199.950 835.950 202.050 838.050 ;
        RECT 196.950 832.950 199.050 835.050 ;
        RECT 155.850 830.700 159.600 831.750 ;
        RECT 133.800 822.600 135.600 825.600 ;
        RECT 149.400 827.700 157.200 829.050 ;
        RECT 149.400 822.600 151.200 827.700 ;
        RECT 155.400 822.600 157.200 827.700 ;
        RECT 158.400 828.600 159.600 830.700 ;
        RECT 176.400 830.700 180.150 831.750 ;
        RECT 176.400 828.600 177.600 830.700 ;
        RECT 158.400 822.600 160.200 828.600 ;
        RECT 175.800 822.600 177.600 828.600 ;
        RECT 178.800 827.700 186.600 829.050 ;
        RECT 178.800 822.600 180.600 827.700 ;
        RECT 184.800 822.600 186.600 827.700 ;
        RECT 200.700 825.600 201.600 835.950 ;
        RECT 203.100 835.050 204.900 836.850 ;
        RECT 218.100 835.050 219.900 836.850 ;
        RECT 220.950 835.950 223.050 838.050 ;
        RECT 239.100 837.150 240.900 838.950 ;
        RECT 242.400 838.050 243.600 851.400 ;
        RECT 251.550 847.050 252.450 853.950 ;
        RECT 250.950 844.950 253.050 847.050 ;
        RECT 260.400 846.600 262.200 857.400 ;
        RECT 266.400 856.500 274.200 857.400 ;
        RECT 266.400 846.600 268.200 856.500 ;
        RECT 260.400 845.700 268.200 846.600 ;
        RECT 269.400 844.500 271.200 855.600 ;
        RECT 272.400 845.400 274.200 856.500 ;
        RECT 289.500 845.400 291.300 857.400 ;
        RECT 295.800 851.400 297.600 857.400 ;
        RECT 266.100 843.600 271.200 844.500 ;
        RECT 244.950 838.950 247.050 841.050 ;
        RECT 202.950 832.950 205.050 835.050 ;
        RECT 217.950 832.950 220.050 835.050 ;
        RECT 221.700 825.600 222.600 835.950 ;
        RECT 224.100 835.050 225.900 836.850 ;
        RECT 241.950 835.950 244.050 838.050 ;
        RECT 245.100 837.150 246.900 838.950 ;
        RECT 266.100 838.050 267.000 843.600 ;
        RECT 290.400 838.050 291.300 845.400 ;
        RECT 293.100 838.050 294.900 839.850 ;
        RECT 259.950 835.950 262.050 838.050 ;
        RECT 223.950 832.950 226.050 835.050 ;
        RECT 242.400 830.700 243.600 835.950 ;
        RECT 260.100 834.150 261.900 835.950 ;
        RECT 263.100 835.050 264.900 836.850 ;
        RECT 265.950 835.950 268.050 838.050 ;
        RECT 262.950 832.950 265.050 835.050 ;
        RECT 242.400 829.800 246.600 830.700 ;
        RECT 200.400 822.600 202.200 825.600 ;
        RECT 221.400 822.600 223.200 825.600 ;
        RECT 244.800 822.600 246.600 829.800 ;
        RECT 265.950 828.600 267.000 835.950 ;
        RECT 269.100 835.050 270.900 836.850 ;
        RECT 271.950 835.950 274.050 838.050 ;
        RECT 289.950 835.950 292.050 838.050 ;
        RECT 292.950 835.950 295.050 838.050 ;
        RECT 268.950 832.950 271.050 835.050 ;
        RECT 272.100 834.150 273.900 835.950 ;
        RECT 265.200 822.600 267.000 828.600 ;
        RECT 290.400 828.600 291.300 835.950 ;
        RECT 296.700 831.300 297.600 851.400 ;
        RECT 313.800 856.500 321.600 857.400 ;
        RECT 313.800 845.400 315.600 856.500 ;
        RECT 316.800 844.500 318.600 855.600 ;
        RECT 319.800 846.600 321.600 856.500 ;
        RECT 325.800 846.600 327.600 857.400 ;
        RECT 319.800 845.700 327.600 846.600 ;
        RECT 340.500 845.400 342.300 857.400 ;
        RECT 346.800 851.400 348.600 857.400 ;
        RECT 316.800 843.600 321.900 844.500 ;
        RECT 321.000 838.050 321.900 843.600 ;
        RECT 340.500 838.050 341.700 845.400 ;
        RECT 347.400 844.500 348.600 851.400 ;
        RECT 361.800 845.400 363.600 857.400 ;
        RECT 364.800 846.300 366.600 857.400 ;
        RECT 370.800 846.300 372.600 857.400 ;
        RECT 385.800 851.400 387.600 857.400 ;
        RECT 364.800 845.400 372.600 846.300 ;
        RECT 386.700 851.100 387.600 851.400 ;
        RECT 391.800 851.400 393.600 857.400 ;
        RECT 397.950 853.950 400.050 856.050 ;
        RECT 391.800 851.100 393.300 851.400 ;
        RECT 386.700 850.200 393.300 851.100 ;
        RECT 342.600 843.600 348.600 844.500 ;
        RECT 342.600 842.700 344.850 843.600 ;
        RECT 298.950 835.950 301.050 838.050 ;
        RECT 313.950 835.950 316.050 838.050 ;
        RECT 299.100 834.150 300.900 835.950 ;
        RECT 314.100 834.150 315.900 835.950 ;
        RECT 317.100 835.050 318.900 836.850 ;
        RECT 319.950 835.950 322.050 838.050 ;
        RECT 316.950 832.950 319.050 835.050 ;
        RECT 293.100 830.400 300.600 831.300 ;
        RECT 293.100 829.500 294.900 830.400 ;
        RECT 290.400 826.800 293.100 828.600 ;
        RECT 291.300 822.600 293.100 826.800 ;
        RECT 298.800 822.600 300.600 830.400 ;
        RECT 321.000 828.600 322.050 835.950 ;
        RECT 323.100 835.050 324.900 836.850 ;
        RECT 325.950 835.950 328.050 838.050 ;
        RECT 340.500 835.950 343.050 838.050 ;
        RECT 322.950 832.950 325.050 835.050 ;
        RECT 326.100 834.150 327.900 835.950 ;
        RECT 340.500 828.600 341.700 835.950 ;
        RECT 343.950 831.300 344.850 842.700 ;
        RECT 347.100 838.050 348.900 839.850 ;
        RECT 362.400 838.050 363.600 845.400 ;
        RECT 364.950 838.950 367.050 841.050 ;
        RECT 346.950 835.950 349.050 838.050 ;
        RECT 361.950 835.950 364.050 838.050 ;
        RECT 365.100 837.150 366.900 838.950 ;
        RECT 368.100 838.050 369.900 839.850 ;
        RECT 370.950 838.950 373.050 841.050 ;
        RECT 367.950 835.950 370.050 838.050 ;
        RECT 371.100 837.150 372.900 838.950 ;
        RECT 386.700 838.050 387.600 850.200 ;
        RECT 398.550 850.050 399.450 853.950 ;
        RECT 410.400 851.400 412.200 857.400 ;
        RECT 434.400 851.400 436.200 857.400 ;
        RECT 442.950 853.950 445.050 856.050 ;
        RECT 397.950 847.950 400.050 850.050 ;
        RECT 398.550 844.050 399.450 847.950 ;
        RECT 397.950 841.950 400.050 844.050 ;
        RECT 388.950 838.950 391.050 841.050 ;
        RECT 385.950 835.950 388.050 838.050 ;
        RECT 389.100 837.150 390.900 838.950 ;
        RECT 392.100 838.050 393.900 839.850 ;
        RECT 394.950 838.950 397.050 841.050 ;
        RECT 406.950 838.950 409.050 841.050 ;
        RECT 391.950 835.950 394.050 838.050 ;
        RECT 395.100 837.150 396.900 838.950 ;
        RECT 407.100 837.150 408.900 838.950 ;
        RECT 410.400 838.050 411.600 851.400 ;
        RECT 412.950 838.950 415.050 841.050 ;
        RECT 430.950 838.950 433.050 841.050 ;
        RECT 409.950 835.950 412.050 838.050 ;
        RECT 413.100 837.150 414.900 838.950 ;
        RECT 431.100 837.150 432.900 838.950 ;
        RECT 434.850 838.050 436.050 851.400 ;
        RECT 443.550 844.050 444.450 853.950 ;
        RECT 452.400 846.600 454.200 857.400 ;
        RECT 458.400 856.500 466.200 857.400 ;
        RECT 458.400 846.600 460.200 856.500 ;
        RECT 452.400 845.700 460.200 846.600 ;
        RECT 461.400 844.500 463.200 855.600 ;
        RECT 464.400 845.400 466.200 856.500 ;
        RECT 482.400 851.400 484.200 857.400 ;
        RECT 487.950 853.950 490.050 856.050 ;
        RECT 469.950 847.950 472.050 850.050 ;
        RECT 442.950 841.950 445.050 844.050 ;
        RECT 458.100 843.600 463.200 844.500 ;
        RECT 436.950 838.950 439.050 841.050 ;
        RECT 433.950 835.950 436.050 838.050 ;
        RECT 437.100 837.150 438.900 838.950 ;
        RECT 440.100 838.050 441.900 839.850 ;
        RECT 458.100 838.050 459.000 843.600 ;
        RECT 439.950 835.950 442.050 838.050 ;
        RECT 451.950 835.950 454.050 838.050 ;
        RECT 342.600 830.400 344.850 831.300 ;
        RECT 342.600 829.500 348.600 830.400 ;
        RECT 321.000 822.600 322.800 828.600 ;
        RECT 340.500 822.600 342.300 828.600 ;
        RECT 347.400 825.600 348.600 829.500 ;
        RECT 362.400 828.600 363.600 835.950 ;
        RECT 386.700 832.200 387.600 835.950 ;
        RECT 386.700 831.000 390.000 832.200 ;
        RECT 362.400 827.400 367.500 828.600 ;
        RECT 346.800 822.600 348.600 825.600 ;
        RECT 365.700 822.600 367.500 827.400 ;
        RECT 388.200 822.600 390.000 831.000 ;
        RECT 410.400 830.700 411.600 835.950 ;
        RECT 424.950 832.950 427.050 835.050 ;
        RECT 410.400 829.800 414.600 830.700 ;
        RECT 412.800 822.600 414.600 829.800 ;
        RECT 425.550 826.050 426.450 832.950 ;
        RECT 433.950 831.750 435.150 835.950 ;
        RECT 452.100 834.150 453.900 835.950 ;
        RECT 455.100 835.050 456.900 836.850 ;
        RECT 457.950 835.950 460.050 838.050 ;
        RECT 454.950 832.950 457.050 835.050 ;
        RECT 431.400 830.700 435.150 831.750 ;
        RECT 431.400 828.600 432.600 830.700 ;
        RECT 424.950 823.950 427.050 826.050 ;
        RECT 430.800 822.600 432.600 828.600 ;
        RECT 433.800 827.700 441.600 829.050 ;
        RECT 457.950 828.600 459.000 835.950 ;
        RECT 461.100 835.050 462.900 836.850 ;
        RECT 463.950 835.950 466.050 838.050 ;
        RECT 460.950 832.950 463.050 835.050 ;
        RECT 464.100 834.150 465.900 835.950 ;
        RECT 470.550 829.050 471.450 847.950 ;
        RECT 482.400 844.050 483.600 851.400 ;
        RECT 479.100 838.050 480.900 839.850 ;
        RECT 481.950 838.950 484.050 844.050 ;
        RECT 478.950 835.950 481.050 838.050 ;
        RECT 433.800 822.600 435.600 827.700 ;
        RECT 439.800 822.600 441.600 827.700 ;
        RECT 457.200 822.600 459.000 828.600 ;
        RECT 469.950 826.950 472.050 829.050 ;
        RECT 482.400 825.600 483.600 838.950 ;
        RECT 488.550 826.050 489.450 853.950 ;
        RECT 500.400 851.400 502.200 857.400 ;
        RECT 496.950 838.950 499.050 841.050 ;
        RECT 497.100 837.150 498.900 838.950 ;
        RECT 500.400 838.050 501.600 851.400 ;
        RECT 520.800 845.400 522.600 857.400 ;
        RECT 523.800 846.300 525.600 857.400 ;
        RECT 529.800 846.300 531.600 857.400 ;
        RECT 544.800 851.400 546.600 857.400 ;
        RECT 523.800 845.400 531.600 846.300 ;
        RECT 502.950 838.950 505.050 841.050 ;
        RECT 499.950 835.950 502.050 838.050 ;
        RECT 503.100 837.150 504.900 838.950 ;
        RECT 521.400 838.050 522.600 845.400 ;
        RECT 545.400 844.050 546.600 851.400 ;
        RECT 563.400 851.400 565.200 857.400 ;
        RECT 586.800 851.400 588.600 857.400 ;
        RECT 610.800 851.400 612.600 857.400 ;
        RECT 535.950 841.950 538.050 844.050 ;
        RECT 523.950 838.950 526.050 841.050 ;
        RECT 520.950 835.950 523.050 838.050 ;
        RECT 524.100 837.150 525.900 838.950 ;
        RECT 527.100 838.050 528.900 839.850 ;
        RECT 529.950 838.950 532.050 841.050 ;
        RECT 526.950 835.950 529.050 838.050 ;
        RECT 530.100 837.150 531.900 838.950 ;
        RECT 500.400 830.700 501.600 835.950 ;
        RECT 500.400 829.800 504.600 830.700 ;
        RECT 482.400 822.600 484.200 825.600 ;
        RECT 487.950 823.950 490.050 826.050 ;
        RECT 502.800 822.600 504.600 829.800 ;
        RECT 521.400 828.600 522.600 835.950 ;
        RECT 536.550 829.050 537.450 841.950 ;
        RECT 544.950 838.950 547.050 844.050 ;
        RECT 521.400 827.400 526.500 828.600 ;
        RECT 524.700 822.600 526.500 827.400 ;
        RECT 532.800 827.550 537.450 829.050 ;
        RECT 532.800 826.950 537.000 827.550 ;
        RECT 545.400 825.600 546.600 838.950 ;
        RECT 548.100 838.050 549.900 839.850 ;
        RECT 559.950 838.950 562.050 841.050 ;
        RECT 547.950 835.950 550.050 838.050 ;
        RECT 560.100 837.150 561.900 838.950 ;
        RECT 563.400 838.050 564.600 851.400 ;
        RECT 565.950 838.950 568.050 841.050 ;
        RECT 562.950 835.950 565.050 838.050 ;
        RECT 566.100 837.150 567.900 838.950 ;
        RECT 581.100 838.050 582.900 839.850 ;
        RECT 583.950 838.950 586.050 841.050 ;
        RECT 580.950 835.950 583.050 838.050 ;
        RECT 584.100 837.150 585.900 838.950 ;
        RECT 586.950 838.050 588.150 851.400 ;
        RECT 589.950 838.950 592.050 841.050 ;
        RECT 586.950 835.950 589.050 838.050 ;
        RECT 590.100 837.150 591.900 838.950 ;
        RECT 605.100 838.050 606.900 839.850 ;
        RECT 607.950 838.950 610.050 841.050 ;
        RECT 604.950 835.950 607.050 838.050 ;
        RECT 608.100 837.150 609.900 838.950 ;
        RECT 610.950 838.050 612.150 851.400 ;
        RECT 631.500 845.400 633.300 857.400 ;
        RECT 637.800 851.400 639.600 857.400 ;
        RECT 649.950 853.950 652.050 856.050 ;
        RECT 613.950 838.950 616.050 841.050 ;
        RECT 610.950 835.950 613.050 838.050 ;
        RECT 614.100 837.150 615.900 838.950 ;
        RECT 632.400 838.050 633.300 845.400 ;
        RECT 635.100 838.050 636.900 839.850 ;
        RECT 631.950 835.950 634.050 838.050 ;
        RECT 634.950 835.950 637.050 838.050 ;
        RECT 563.400 830.700 564.600 835.950 ;
        RECT 587.850 831.750 589.050 835.950 ;
        RECT 611.850 831.750 613.050 835.950 ;
        RECT 587.850 830.700 591.600 831.750 ;
        RECT 611.850 830.700 615.600 831.750 ;
        RECT 563.400 829.800 567.600 830.700 ;
        RECT 544.800 822.600 546.600 825.600 ;
        RECT 565.800 822.600 567.600 829.800 ;
        RECT 581.400 827.700 589.200 829.050 ;
        RECT 581.400 822.600 583.200 827.700 ;
        RECT 587.400 822.600 589.200 827.700 ;
        RECT 590.400 828.600 591.600 830.700 ;
        RECT 590.400 822.600 592.200 828.600 ;
        RECT 605.400 827.700 613.200 829.050 ;
        RECT 605.400 822.600 607.200 827.700 ;
        RECT 611.400 822.600 613.200 827.700 ;
        RECT 614.400 828.600 615.600 830.700 ;
        RECT 632.400 828.600 633.300 835.950 ;
        RECT 638.700 831.300 639.600 851.400 ;
        RECT 640.950 835.950 643.050 838.050 ;
        RECT 641.100 834.150 642.900 835.950 ;
        RECT 650.550 832.050 651.450 853.950 ;
        RECT 655.800 845.400 657.600 857.400 ;
        RECT 677.400 851.400 679.200 857.400 ;
        RECT 700.800 851.400 702.600 857.400 ;
        RECT 709.950 853.950 712.050 856.050 ;
        RECT 656.400 838.050 657.600 845.400 ;
        RECT 658.950 838.950 661.050 841.050 ;
        RECT 673.950 838.950 676.050 841.050 ;
        RECT 655.950 835.950 658.050 838.050 ;
        RECT 659.100 837.150 660.900 838.950 ;
        RECT 674.100 837.150 675.900 838.950 ;
        RECT 677.850 838.050 679.050 851.400 ;
        RECT 679.950 838.950 682.050 841.050 ;
        RECT 676.950 835.950 679.050 838.050 ;
        RECT 680.100 837.150 681.900 838.950 ;
        RECT 683.100 838.050 684.900 839.850 ;
        RECT 697.950 838.950 700.050 841.050 ;
        RECT 682.950 835.950 685.050 838.050 ;
        RECT 698.100 837.150 699.900 838.950 ;
        RECT 701.400 838.050 702.600 851.400 ;
        RECT 703.950 838.950 706.050 841.050 ;
        RECT 700.950 835.950 703.050 838.050 ;
        RECT 704.100 837.150 705.900 838.950 ;
        RECT 635.100 830.400 642.600 831.300 ;
        RECT 635.100 829.500 636.900 830.400 ;
        RECT 614.400 822.600 616.200 828.600 ;
        RECT 632.400 826.800 635.100 828.600 ;
        RECT 633.300 822.600 635.100 826.800 ;
        RECT 640.800 822.600 642.600 830.400 ;
        RECT 649.950 829.950 652.050 832.050 ;
        RECT 656.400 828.600 657.600 835.950 ;
        RECT 676.950 831.750 678.150 835.950 ;
        RECT 674.400 830.700 678.150 831.750 ;
        RECT 701.400 830.700 702.600 835.950 ;
        RECT 710.550 832.050 711.450 853.950 ;
        RECT 716.400 846.600 718.200 857.400 ;
        RECT 722.400 856.500 730.200 857.400 ;
        RECT 722.400 846.600 724.200 856.500 ;
        RECT 716.400 845.700 724.200 846.600 ;
        RECT 725.400 844.500 727.200 855.600 ;
        RECT 728.400 845.400 730.200 856.500 ;
        RECT 746.400 851.400 748.200 857.400 ;
        RECT 746.700 851.100 748.200 851.400 ;
        RECT 752.400 851.400 754.200 857.400 ;
        RECT 757.950 853.950 760.050 856.050 ;
        RECT 752.400 851.100 753.300 851.400 ;
        RECT 746.700 850.200 753.300 851.100 ;
        RECT 736.950 844.950 739.050 847.050 ;
        RECT 722.100 843.600 727.200 844.500 ;
        RECT 722.100 838.050 723.000 843.600 ;
        RECT 715.950 835.950 718.050 838.050 ;
        RECT 716.100 834.150 717.900 835.950 ;
        RECT 719.100 835.050 720.900 836.850 ;
        RECT 721.950 835.950 724.050 838.050 ;
        RECT 718.950 832.950 721.050 835.050 ;
        RECT 674.400 828.600 675.600 830.700 ;
        RECT 698.400 829.800 702.600 830.700 ;
        RECT 709.950 829.950 712.050 832.050 ;
        RECT 655.800 822.600 657.600 828.600 ;
        RECT 673.800 822.600 675.600 828.600 ;
        RECT 676.800 827.700 684.600 829.050 ;
        RECT 676.800 822.600 678.600 827.700 ;
        RECT 682.800 822.600 684.600 827.700 ;
        RECT 698.400 822.600 700.200 829.800 ;
        RECT 721.950 828.600 723.000 835.950 ;
        RECT 725.100 835.050 726.900 836.850 ;
        RECT 727.950 835.950 730.050 838.050 ;
        RECT 724.950 832.950 727.050 835.050 ;
        RECT 728.100 834.150 729.900 835.950 ;
        RECT 737.550 829.050 738.450 844.950 ;
        RECT 742.950 838.950 745.050 841.050 ;
        RECT 743.100 837.150 744.900 838.950 ;
        RECT 746.100 838.050 747.900 839.850 ;
        RECT 748.950 838.950 751.050 841.050 ;
        RECT 745.950 835.950 748.050 838.050 ;
        RECT 749.100 837.150 750.900 838.950 ;
        RECT 752.400 838.050 753.300 850.200 ;
        RECT 751.950 835.950 754.050 838.050 ;
        RECT 752.400 832.200 753.300 835.950 ;
        RECT 758.550 835.050 759.450 853.950 ;
        RECT 770.400 851.400 772.200 857.400 ;
        RECT 766.950 835.950 769.050 838.050 ;
        RECT 757.950 832.950 760.050 835.050 ;
        RECT 767.100 834.150 768.900 835.950 ;
        RECT 750.000 831.000 753.300 832.200 ;
        RECT 770.400 831.300 771.300 851.400 ;
        RECT 776.700 845.400 778.500 857.400 ;
        RECT 796.800 851.400 798.600 857.400 ;
        RECT 773.100 838.050 774.900 839.850 ;
        RECT 776.700 838.050 777.600 845.400 ;
        RECT 793.950 838.950 796.050 841.050 ;
        RECT 772.950 835.950 775.050 838.050 ;
        RECT 775.950 835.950 778.050 838.050 ;
        RECT 794.100 837.150 795.900 838.950 ;
        RECT 797.400 838.050 798.600 851.400 ;
        RECT 805.950 847.950 808.050 850.050 ;
        RECT 799.950 838.950 802.050 841.050 ;
        RECT 796.950 835.950 799.050 838.050 ;
        RECT 800.100 837.150 801.900 838.950 ;
        RECT 721.200 822.600 723.000 828.600 ;
        RECT 736.950 826.950 739.050 829.050 ;
        RECT 750.000 822.600 751.800 831.000 ;
        RECT 767.400 830.400 774.900 831.300 ;
        RECT 767.400 822.600 769.200 830.400 ;
        RECT 773.100 829.500 774.900 830.400 ;
        RECT 776.700 828.600 777.600 835.950 ;
        RECT 797.400 830.700 798.600 835.950 ;
        RECT 774.900 826.800 777.600 828.600 ;
        RECT 794.400 829.800 798.600 830.700 ;
        RECT 774.900 822.600 776.700 826.800 ;
        RECT 794.400 822.600 796.200 829.800 ;
        RECT 806.550 826.050 807.450 847.950 ;
        RECT 812.400 846.300 814.200 857.400 ;
        RECT 818.400 846.300 820.200 857.400 ;
        RECT 812.400 845.400 820.200 846.300 ;
        RECT 821.400 845.400 823.200 857.400 ;
        RECT 841.500 846.600 843.300 857.400 ;
        RECT 850.950 853.950 853.050 856.050 ;
        RECT 839.700 845.400 843.300 846.600 ;
        RECT 811.950 838.950 814.050 841.050 ;
        RECT 812.100 837.150 813.900 838.950 ;
        RECT 815.100 838.050 816.900 839.850 ;
        RECT 817.950 838.950 820.050 841.050 ;
        RECT 814.950 835.950 817.050 838.050 ;
        RECT 818.100 837.150 819.900 838.950 ;
        RECT 821.400 838.050 822.600 845.400 ;
        RECT 839.700 838.050 840.600 845.400 ;
        RECT 820.950 835.950 823.050 838.050 ;
        RECT 821.400 828.600 822.600 835.950 ;
        RECT 836.100 835.050 837.900 836.850 ;
        RECT 838.950 835.950 841.050 838.050 ;
        RECT 835.950 832.950 838.050 835.050 ;
        RECT 817.500 827.400 822.600 828.600 ;
        RECT 805.950 823.950 808.050 826.050 ;
        RECT 817.500 822.600 819.300 827.400 ;
        RECT 839.700 825.600 840.600 835.950 ;
        RECT 842.100 835.050 843.900 836.850 ;
        RECT 841.950 832.950 844.050 835.050 ;
        RECT 851.550 826.050 852.450 853.950 ;
        RECT 862.800 851.400 864.600 857.400 ;
        RECT 859.950 838.950 862.050 841.050 ;
        RECT 860.100 837.150 861.900 838.950 ;
        RECT 863.400 838.050 864.600 851.400 ;
        RECT 881.400 851.400 883.200 857.400 ;
        RECT 902.400 851.400 904.200 857.400 ;
        RECT 871.950 841.950 874.050 844.050 ;
        RECT 865.950 838.950 868.050 841.050 ;
        RECT 862.950 835.950 865.050 838.050 ;
        RECT 866.100 837.150 867.900 838.950 ;
        RECT 872.550 838.050 873.450 841.950 ;
        RECT 877.950 838.950 880.050 841.050 ;
        RECT 871.950 835.950 874.050 838.050 ;
        RECT 878.100 837.150 879.900 838.950 ;
        RECT 881.400 838.050 882.600 851.400 ;
        RECT 883.950 838.950 886.050 841.050 ;
        RECT 898.950 838.950 901.050 841.050 ;
        RECT 880.950 835.950 883.050 838.050 ;
        RECT 884.100 837.150 885.900 838.950 ;
        RECT 899.100 837.150 900.900 838.950 ;
        RECT 902.400 838.050 903.600 851.400 ;
        RECT 904.950 838.950 907.050 841.050 ;
        RECT 901.950 835.950 904.050 838.050 ;
        RECT 905.100 837.150 906.900 838.950 ;
        RECT 863.400 830.700 864.600 835.950 ;
        RECT 839.400 822.600 841.200 825.600 ;
        RECT 847.950 824.550 852.450 826.050 ;
        RECT 860.400 829.800 864.600 830.700 ;
        RECT 881.400 830.700 882.600 835.950 ;
        RECT 902.400 830.700 903.600 835.950 ;
        RECT 881.400 829.800 885.600 830.700 ;
        RECT 902.400 829.800 906.600 830.700 ;
        RECT 907.950 829.950 910.050 832.050 ;
        RECT 847.950 823.950 852.000 824.550 ;
        RECT 860.400 822.600 862.200 829.800 ;
        RECT 883.800 822.600 885.600 829.800 ;
        RECT 904.800 822.600 906.600 829.800 ;
        RECT 908.550 826.050 909.450 829.950 ;
        RECT 907.950 823.950 910.050 826.050 ;
        RECT 17.700 813.600 19.500 818.400 ;
        RECT 28.950 814.950 31.050 817.050 ;
        RECT 14.400 812.400 19.500 813.600 ;
        RECT 14.400 805.050 15.600 812.400 ;
        RECT 13.950 802.950 16.050 805.050 ;
        RECT 14.400 795.600 15.600 802.950 ;
        RECT 17.100 802.050 18.900 803.850 ;
        RECT 19.950 802.950 22.050 805.050 ;
        RECT 16.950 799.950 19.050 802.050 ;
        RECT 20.100 801.150 21.900 802.950 ;
        RECT 23.100 802.050 24.900 803.850 ;
        RECT 22.950 799.950 25.050 802.050 ;
        RECT 13.800 783.600 15.600 795.600 ;
        RECT 16.800 794.700 24.600 795.600 ;
        RECT 16.800 783.600 18.600 794.700 ;
        RECT 22.800 783.600 24.600 794.700 ;
        RECT 29.550 790.050 30.450 814.950 ;
        RECT 37.800 812.400 39.600 818.400 ;
        RECT 38.400 810.300 39.600 812.400 ;
        RECT 40.800 813.300 42.600 818.400 ;
        RECT 46.800 813.300 48.600 818.400 ;
        RECT 40.800 811.950 48.600 813.300 ;
        RECT 61.800 812.400 63.600 818.400 ;
        RECT 62.400 810.300 63.600 812.400 ;
        RECT 64.800 813.300 66.600 818.400 ;
        RECT 70.800 813.300 72.600 818.400 ;
        RECT 64.800 811.950 72.600 813.300 ;
        RECT 38.400 809.250 42.150 810.300 ;
        RECT 62.400 809.250 66.150 810.300 ;
        RECT 88.200 810.000 90.000 818.400 ;
        RECT 100.950 811.950 103.050 814.050 ;
        RECT 113.700 813.600 115.500 818.400 ;
        RECT 124.950 814.950 127.050 817.050 ;
        RECT 133.800 815.400 135.600 818.400 ;
        RECT 110.400 812.400 115.500 813.600 ;
        RECT 40.950 805.050 42.150 809.250 ;
        RECT 64.950 805.050 66.150 809.250 ;
        RECT 86.700 808.800 90.000 810.000 ;
        RECT 86.700 805.050 87.600 808.800 ;
        RECT 38.100 802.050 39.900 803.850 ;
        RECT 40.950 802.950 43.050 805.050 ;
        RECT 37.950 799.950 40.050 802.050 ;
        RECT 28.950 787.950 31.050 790.050 ;
        RECT 41.850 789.600 43.050 802.950 ;
        RECT 44.100 802.050 45.900 803.850 ;
        RECT 46.950 802.950 49.050 805.050 ;
        RECT 43.950 799.950 46.050 802.050 ;
        RECT 47.100 801.150 48.900 802.950 ;
        RECT 62.100 802.050 63.900 803.850 ;
        RECT 64.950 802.950 67.050 805.050 ;
        RECT 61.950 799.950 64.050 802.050 ;
        RECT 65.850 789.600 67.050 802.950 ;
        RECT 68.100 802.050 69.900 803.850 ;
        RECT 70.950 802.950 73.050 805.050 ;
        RECT 85.950 802.950 88.050 805.050 ;
        RECT 67.950 799.950 70.050 802.050 ;
        RECT 71.100 801.150 72.900 802.950 ;
        RECT 86.700 790.800 87.600 802.950 ;
        RECT 89.100 802.050 90.900 803.850 ;
        RECT 91.950 802.950 94.050 805.050 ;
        RECT 88.950 799.950 91.050 802.050 ;
        RECT 92.100 801.150 93.900 802.950 ;
        RECT 95.100 802.050 96.900 803.850 ;
        RECT 94.950 799.950 97.050 802.050 ;
        RECT 86.700 789.900 93.300 790.800 ;
        RECT 86.700 789.600 87.600 789.900 ;
        RECT 41.400 783.600 43.200 789.600 ;
        RECT 65.400 783.600 67.200 789.600 ;
        RECT 85.800 783.600 87.600 789.600 ;
        RECT 91.800 789.600 93.300 789.900 ;
        RECT 91.800 783.600 93.600 789.600 ;
        RECT 101.550 787.050 102.450 811.950 ;
        RECT 110.400 805.050 111.600 812.400 ;
        RECT 109.950 802.950 112.050 805.050 ;
        RECT 110.400 795.600 111.600 802.950 ;
        RECT 113.100 802.050 114.900 803.850 ;
        RECT 115.950 802.950 118.050 805.050 ;
        RECT 112.950 799.950 115.050 802.050 ;
        RECT 116.100 801.150 117.900 802.950 ;
        RECT 119.100 802.050 120.900 803.850 ;
        RECT 118.950 799.950 121.050 802.050 ;
        RECT 125.550 799.050 126.450 814.950 ;
        RECT 134.400 802.050 135.600 815.400 ;
        RECT 152.400 811.200 154.200 818.400 ;
        RECT 163.950 814.950 166.050 817.050 ;
        RECT 152.400 810.300 156.600 811.200 ;
        RECT 155.400 805.050 156.600 810.300 ;
        RECT 136.950 802.950 139.050 805.050 ;
        RECT 124.950 796.950 127.050 799.050 ;
        RECT 133.950 796.950 136.050 802.050 ;
        RECT 137.100 801.150 138.900 802.950 ;
        RECT 152.100 802.050 153.900 803.850 ;
        RECT 154.950 802.950 157.050 805.050 ;
        RECT 151.950 799.950 154.050 802.050 ;
        RECT 100.950 784.950 103.050 787.050 ;
        RECT 109.800 783.600 111.600 795.600 ;
        RECT 112.800 794.700 120.600 795.600 ;
        RECT 112.800 783.600 114.600 794.700 ;
        RECT 118.800 783.600 120.600 794.700 ;
        RECT 134.400 789.600 135.600 796.950 ;
        RECT 155.400 789.600 156.600 802.950 ;
        RECT 158.100 802.050 159.900 803.850 ;
        RECT 157.950 799.950 160.050 802.050 ;
        RECT 164.550 799.050 165.450 814.950 ;
        RECT 172.800 812.400 174.600 818.400 ;
        RECT 173.400 810.300 174.600 812.400 ;
        RECT 175.800 813.300 177.600 818.400 ;
        RECT 181.800 813.300 183.600 818.400 ;
        RECT 175.800 811.950 183.600 813.300 ;
        RECT 197.400 811.200 199.200 818.400 ;
        RECT 219.300 814.200 221.100 818.400 ;
        RECT 218.400 812.400 221.100 814.200 ;
        RECT 197.400 810.300 201.600 811.200 ;
        RECT 173.400 809.250 177.150 810.300 ;
        RECT 166.950 805.950 169.050 808.050 ;
        RECT 163.950 796.950 166.050 799.050 ;
        RECT 164.550 793.050 165.450 796.950 ;
        RECT 163.950 790.950 166.050 793.050 ;
        RECT 133.800 783.600 135.600 789.600 ;
        RECT 154.800 783.600 156.600 789.600 ;
        RECT 167.550 787.050 168.450 805.950 ;
        RECT 175.950 805.050 177.150 809.250 ;
        RECT 200.400 805.050 201.600 810.300 ;
        RECT 211.950 808.950 214.050 811.050 ;
        RECT 173.100 802.050 174.900 803.850 ;
        RECT 175.950 802.950 178.050 805.050 ;
        RECT 172.950 799.950 175.050 802.050 ;
        RECT 176.850 789.600 178.050 802.950 ;
        RECT 179.100 802.050 180.900 803.850 ;
        RECT 181.950 802.950 184.050 805.050 ;
        RECT 178.950 799.950 181.050 802.050 ;
        RECT 182.100 801.150 183.900 802.950 ;
        RECT 197.100 802.050 198.900 803.850 ;
        RECT 199.950 802.950 202.050 805.050 ;
        RECT 196.950 799.950 199.050 802.050 ;
        RECT 200.400 789.600 201.600 802.950 ;
        RECT 203.100 802.050 204.900 803.850 ;
        RECT 202.950 799.950 205.050 802.050 ;
        RECT 212.550 790.050 213.450 808.950 ;
        RECT 218.400 805.050 219.300 812.400 ;
        RECT 221.100 810.600 222.900 811.500 ;
        RECT 226.800 810.600 228.600 818.400 ;
        RECT 221.100 809.700 228.600 810.600 ;
        RECT 241.500 812.400 243.300 818.400 ;
        RECT 247.800 815.400 249.600 818.400 ;
        RECT 217.950 802.950 220.050 805.050 ;
        RECT 220.950 802.950 223.050 805.050 ;
        RECT 218.400 795.600 219.300 802.950 ;
        RECT 221.100 801.150 222.900 802.950 ;
        RECT 166.950 784.950 169.050 787.050 ;
        RECT 176.400 783.600 178.200 789.600 ;
        RECT 199.800 783.600 201.600 789.600 ;
        RECT 212.100 787.950 214.200 790.050 ;
        RECT 217.500 783.600 219.300 795.600 ;
        RECT 224.700 789.600 225.600 809.700 ;
        RECT 227.100 805.050 228.900 806.850 ;
        RECT 241.500 805.050 242.700 812.400 ;
        RECT 248.400 811.500 249.600 815.400 ;
        RECT 256.950 814.950 259.050 817.050 ;
        RECT 243.600 810.600 249.600 811.500 ;
        RECT 243.600 809.700 245.850 810.600 ;
        RECT 226.950 802.950 229.050 805.050 ;
        RECT 241.500 802.950 244.050 805.050 ;
        RECT 223.800 783.600 225.600 789.600 ;
        RECT 241.500 795.600 242.700 802.950 ;
        RECT 244.950 798.300 245.850 809.700 ;
        RECT 247.950 802.950 250.050 805.050 ;
        RECT 248.100 801.150 249.900 802.950 ;
        RECT 243.600 797.400 245.850 798.300 ;
        RECT 243.600 796.500 249.600 797.400 ;
        RECT 241.500 783.600 243.300 795.600 ;
        RECT 248.400 789.600 249.600 796.500 ;
        RECT 257.550 793.050 258.450 814.950 ;
        RECT 265.200 810.000 267.000 818.400 ;
        RECT 286.800 812.400 288.600 818.400 ;
        RECT 263.700 808.800 267.000 810.000 ;
        RECT 287.400 810.300 288.600 812.400 ;
        RECT 289.800 813.300 291.600 818.400 ;
        RECT 295.800 813.300 297.600 818.400 ;
        RECT 289.800 811.950 297.600 813.300 ;
        RECT 310.800 812.400 312.600 818.400 ;
        RECT 311.400 810.300 312.600 812.400 ;
        RECT 313.800 813.300 315.600 818.400 ;
        RECT 319.800 813.300 321.600 818.400 ;
        RECT 338.700 813.600 340.500 818.400 ;
        RECT 313.800 811.950 321.600 813.300 ;
        RECT 335.400 812.400 340.500 813.600 ;
        RECT 287.400 809.250 291.150 810.300 ;
        RECT 311.400 809.250 315.150 810.300 ;
        RECT 263.700 805.050 264.600 808.800 ;
        RECT 277.950 805.950 280.050 808.050 ;
        RECT 262.950 802.950 265.050 805.050 ;
        RECT 256.950 790.950 259.050 793.050 ;
        RECT 263.700 790.800 264.600 802.950 ;
        RECT 266.100 802.050 267.900 803.850 ;
        RECT 268.950 802.950 271.050 805.050 ;
        RECT 265.950 799.950 268.050 802.050 ;
        RECT 269.100 801.150 270.900 802.950 ;
        RECT 272.100 802.050 273.900 803.850 ;
        RECT 271.950 799.950 274.050 802.050 ;
        RECT 263.700 789.900 270.300 790.800 ;
        RECT 263.700 789.600 264.600 789.900 ;
        RECT 247.800 783.600 249.600 789.600 ;
        RECT 262.800 783.600 264.600 789.600 ;
        RECT 268.800 789.600 270.300 789.900 ;
        RECT 268.800 783.600 270.600 789.600 ;
        RECT 278.550 787.050 279.450 805.950 ;
        RECT 289.950 805.050 291.150 809.250 ;
        RECT 313.950 805.050 315.150 809.250 ;
        RECT 335.400 805.050 336.600 812.400 ;
        RECT 361.200 810.000 363.000 818.400 ;
        RECT 382.800 815.400 384.600 818.400 ;
        RECT 359.700 808.800 363.000 810.000 ;
        RECT 359.700 805.050 360.600 808.800 ;
        RECT 287.100 802.050 288.900 803.850 ;
        RECT 289.950 802.950 292.050 805.050 ;
        RECT 286.950 799.950 289.050 802.050 ;
        RECT 290.850 789.600 292.050 802.950 ;
        RECT 293.100 802.050 294.900 803.850 ;
        RECT 295.950 802.950 298.050 805.050 ;
        RECT 292.950 799.950 295.050 802.050 ;
        RECT 296.100 801.150 297.900 802.950 ;
        RECT 311.100 802.050 312.900 803.850 ;
        RECT 313.950 802.950 316.050 805.050 ;
        RECT 310.950 799.950 313.050 802.050 ;
        RECT 314.850 789.600 316.050 802.950 ;
        RECT 317.100 802.050 318.900 803.850 ;
        RECT 319.950 802.950 322.050 805.050 ;
        RECT 334.950 802.950 337.050 805.050 ;
        RECT 316.950 799.950 319.050 802.050 ;
        RECT 320.100 801.150 321.900 802.950 ;
        RECT 335.400 795.600 336.600 802.950 ;
        RECT 338.100 802.050 339.900 803.850 ;
        RECT 340.950 802.950 343.050 805.050 ;
        RECT 337.950 799.950 340.050 802.050 ;
        RECT 341.100 801.150 342.900 802.950 ;
        RECT 344.100 802.050 345.900 803.850 ;
        RECT 358.950 802.950 361.050 805.050 ;
        RECT 343.950 799.950 346.050 802.050 ;
        RECT 274.800 785.550 279.450 787.050 ;
        RECT 274.800 784.950 279.000 785.550 ;
        RECT 290.400 783.600 292.200 789.600 ;
        RECT 314.400 783.600 316.200 789.600 ;
        RECT 334.800 783.600 336.600 795.600 ;
        RECT 337.800 794.700 345.600 795.600 ;
        RECT 337.800 783.600 339.600 794.700 ;
        RECT 343.800 783.600 345.600 794.700 ;
        RECT 346.950 790.950 349.050 793.050 ;
        RECT 347.550 787.050 348.450 790.950 ;
        RECT 359.700 790.800 360.600 802.950 ;
        RECT 362.100 802.050 363.900 803.850 ;
        RECT 364.950 802.950 367.050 805.050 ;
        RECT 361.950 799.950 364.050 802.050 ;
        RECT 365.100 801.150 366.900 802.950 ;
        RECT 368.100 802.050 369.900 803.850 ;
        RECT 383.400 802.050 384.600 815.400 ;
        RECT 403.500 813.600 405.300 818.400 ;
        RECT 418.950 814.950 421.050 817.050 ;
        RECT 403.500 812.400 408.600 813.600 ;
        RECT 407.400 805.050 408.600 812.400 ;
        RECT 412.950 805.950 415.050 808.050 ;
        RECT 385.950 802.950 388.050 805.050 ;
        RECT 367.950 799.950 370.050 802.050 ;
        RECT 382.950 796.950 385.050 802.050 ;
        RECT 386.100 801.150 387.900 802.950 ;
        RECT 398.100 802.050 399.900 803.850 ;
        RECT 400.950 802.950 403.050 805.050 ;
        RECT 397.950 799.950 400.050 802.050 ;
        RECT 401.100 801.150 402.900 802.950 ;
        RECT 404.100 802.050 405.900 803.850 ;
        RECT 406.950 802.950 409.050 805.050 ;
        RECT 403.950 799.950 406.050 802.050 ;
        RECT 359.700 789.900 366.300 790.800 ;
        RECT 359.700 789.600 360.600 789.900 ;
        RECT 346.950 784.950 349.050 787.050 ;
        RECT 358.800 783.600 360.600 789.600 ;
        RECT 364.800 789.600 366.300 789.900 ;
        RECT 383.400 789.600 384.600 796.950 ;
        RECT 407.400 795.600 408.600 802.950 ;
        RECT 364.800 783.600 366.600 789.600 ;
        RECT 382.800 783.600 384.600 789.600 ;
        RECT 398.400 794.700 406.200 795.600 ;
        RECT 398.400 783.600 400.200 794.700 ;
        RECT 404.400 783.600 406.200 794.700 ;
        RECT 407.400 783.600 409.200 795.600 ;
        RECT 413.550 790.050 414.450 805.950 ;
        RECT 415.950 793.950 418.050 796.050 ;
        RECT 412.800 787.950 414.900 790.050 ;
        RECT 416.550 787.050 417.450 793.950 ;
        RECT 419.550 790.050 420.450 814.950 ;
        RECT 424.800 812.400 426.600 818.400 ;
        RECT 425.400 810.300 426.600 812.400 ;
        RECT 427.800 813.300 429.600 818.400 ;
        RECT 433.800 813.300 435.600 818.400 ;
        RECT 427.800 811.950 435.600 813.300 ;
        RECT 439.950 811.950 442.050 814.050 ;
        RECT 448.800 812.400 450.600 818.400 ;
        RECT 425.400 809.250 429.150 810.300 ;
        RECT 427.950 805.050 429.150 809.250 ;
        RECT 425.100 802.050 426.900 803.850 ;
        RECT 427.950 802.950 430.050 805.050 ;
        RECT 424.950 799.950 427.050 802.050 ;
        RECT 418.950 787.950 421.050 790.050 ;
        RECT 428.850 789.600 430.050 802.950 ;
        RECT 431.100 802.050 432.900 803.850 ;
        RECT 433.950 802.950 436.050 805.050 ;
        RECT 430.950 799.950 433.050 802.050 ;
        RECT 434.100 801.150 435.900 802.950 ;
        RECT 436.950 796.950 439.050 799.050 ;
        RECT 437.550 790.050 438.450 796.950 ;
        RECT 415.950 784.950 418.050 787.050 ;
        RECT 428.400 783.600 430.200 789.600 ;
        RECT 436.800 787.950 438.900 790.050 ;
        RECT 440.550 787.050 441.450 811.950 ;
        RECT 449.400 810.300 450.600 812.400 ;
        RECT 451.800 813.300 453.600 818.400 ;
        RECT 457.800 813.300 459.600 818.400 ;
        RECT 467.100 814.950 469.200 817.050 ;
        RECT 451.800 811.950 459.600 813.300 ;
        RECT 449.400 809.250 453.150 810.300 ;
        RECT 451.950 805.050 453.150 809.250 ;
        RECT 449.100 802.050 450.900 803.850 ;
        RECT 451.950 802.950 454.050 805.050 ;
        RECT 448.950 799.950 451.050 802.050 ;
        RECT 452.850 789.600 454.050 802.950 ;
        RECT 455.100 802.050 456.900 803.850 ;
        RECT 457.950 802.950 460.050 805.050 ;
        RECT 454.950 799.950 457.050 802.050 ;
        RECT 458.100 801.150 459.900 802.950 ;
        RECT 467.550 799.050 468.450 814.950 ;
        RECT 475.200 810.000 477.000 818.400 ;
        RECT 473.700 808.800 477.000 810.000 ;
        RECT 504.000 812.400 505.800 818.400 ;
        RECT 523.800 812.400 525.600 818.400 ;
        RECT 473.700 805.050 474.600 808.800 ;
        RECT 497.100 805.050 498.900 806.850 ;
        RECT 499.950 805.950 502.050 808.050 ;
        RECT 472.950 802.950 475.050 805.050 ;
        RECT 466.950 796.950 469.050 799.050 ;
        RECT 473.700 790.800 474.600 802.950 ;
        RECT 476.100 802.050 477.900 803.850 ;
        RECT 478.950 802.950 481.050 805.050 ;
        RECT 475.950 799.950 478.050 802.050 ;
        RECT 479.100 801.150 480.900 802.950 ;
        RECT 482.100 802.050 483.900 803.850 ;
        RECT 496.950 802.950 499.050 805.050 ;
        RECT 500.100 804.150 501.900 805.950 ;
        RECT 504.000 805.050 505.050 812.400 ;
        RECT 514.950 808.950 517.050 811.050 ;
        RECT 524.400 810.300 525.600 812.400 ;
        RECT 526.800 813.300 528.600 818.400 ;
        RECT 532.800 813.300 534.600 818.400 ;
        RECT 526.800 811.950 534.600 813.300 ;
        RECT 541.950 811.950 544.050 814.050 ;
        RECT 555.000 812.400 556.800 818.400 ;
        RECT 524.400 809.250 528.150 810.300 ;
        RECT 505.950 805.950 508.050 808.050 ;
        RECT 502.950 802.950 505.050 805.050 ;
        RECT 506.100 804.150 507.900 805.950 ;
        RECT 509.100 805.050 510.900 806.850 ;
        RECT 508.950 802.950 511.050 805.050 ;
        RECT 481.950 799.950 484.050 802.050 ;
        RECT 504.000 797.400 504.900 802.950 ;
        RECT 499.800 796.500 504.900 797.400 ;
        RECT 473.700 789.900 480.300 790.800 ;
        RECT 473.700 789.600 474.600 789.900 ;
        RECT 439.950 784.950 442.050 787.050 ;
        RECT 452.400 783.600 454.200 789.600 ;
        RECT 472.800 783.600 474.600 789.600 ;
        RECT 478.800 789.600 480.300 789.900 ;
        RECT 478.800 783.600 480.600 789.600 ;
        RECT 496.800 784.500 498.600 795.600 ;
        RECT 499.800 785.400 501.600 796.500 ;
        RECT 502.800 794.400 510.600 795.300 ;
        RECT 502.800 784.500 504.600 794.400 ;
        RECT 496.800 783.600 504.600 784.500 ;
        RECT 508.800 783.600 510.600 794.400 ;
        RECT 515.550 793.050 516.450 808.950 ;
        RECT 526.950 805.050 528.150 809.250 ;
        RECT 524.100 802.050 525.900 803.850 ;
        RECT 526.950 802.950 529.050 805.050 ;
        RECT 523.950 799.950 526.050 802.050 ;
        RECT 517.950 793.950 520.050 796.050 ;
        RECT 514.950 790.950 517.050 793.050 ;
        RECT 518.550 790.050 519.450 793.950 ;
        RECT 517.950 787.950 520.050 790.050 ;
        RECT 527.850 789.600 529.050 802.950 ;
        RECT 530.100 802.050 531.900 803.850 ;
        RECT 532.950 802.950 535.050 805.050 ;
        RECT 529.950 799.950 532.050 802.050 ;
        RECT 533.100 801.150 534.900 802.950 ;
        RECT 527.400 783.600 529.200 789.600 ;
        RECT 542.550 787.050 543.450 811.950 ;
        RECT 548.100 805.050 549.900 806.850 ;
        RECT 550.950 805.950 553.050 808.050 ;
        RECT 547.950 802.950 550.050 805.050 ;
        RECT 551.100 804.150 552.900 805.950 ;
        RECT 555.000 805.050 556.050 812.400 ;
        RECT 572.400 810.600 574.200 818.400 ;
        RECT 579.900 814.200 581.700 818.400 ;
        RECT 579.900 812.400 582.600 814.200 ;
        RECT 578.100 810.600 579.900 811.500 ;
        RECT 572.400 809.700 579.900 810.600 ;
        RECT 556.950 805.950 559.050 808.050 ;
        RECT 553.950 802.950 556.050 805.050 ;
        RECT 557.100 804.150 558.900 805.950 ;
        RECT 560.100 805.050 561.900 806.850 ;
        RECT 572.100 805.050 573.900 806.850 ;
        RECT 559.950 802.950 562.050 805.050 ;
        RECT 571.950 802.950 574.050 805.050 ;
        RECT 555.000 797.400 555.900 802.950 ;
        RECT 550.800 796.500 555.900 797.400 ;
        RECT 541.950 784.950 544.050 787.050 ;
        RECT 547.800 784.500 549.600 795.600 ;
        RECT 550.800 785.400 552.600 796.500 ;
        RECT 553.800 794.400 561.600 795.300 ;
        RECT 553.800 784.500 555.600 794.400 ;
        RECT 547.800 783.600 555.600 784.500 ;
        RECT 559.800 783.600 561.600 794.400 ;
        RECT 575.400 789.600 576.300 809.700 ;
        RECT 581.700 805.050 582.600 812.400 ;
        RECT 599.400 811.200 601.200 818.400 ;
        RECT 610.950 814.950 613.050 817.050 ;
        RECT 599.400 810.300 603.600 811.200 ;
        RECT 602.400 805.050 603.600 810.300 ;
        RECT 611.550 808.050 612.450 814.950 ;
        RECT 614.100 811.950 616.200 814.050 ;
        RECT 610.950 805.950 613.050 808.050 ;
        RECT 577.950 802.950 580.050 805.050 ;
        RECT 580.950 802.950 583.050 805.050 ;
        RECT 578.100 801.150 579.900 802.950 ;
        RECT 581.700 795.600 582.600 802.950 ;
        RECT 599.100 802.050 600.900 803.850 ;
        RECT 601.950 802.950 604.050 805.050 ;
        RECT 598.950 799.950 601.050 802.050 ;
        RECT 575.400 783.600 577.200 789.600 ;
        RECT 581.700 783.600 583.500 795.600 ;
        RECT 602.400 789.600 603.600 802.950 ;
        RECT 605.100 802.050 606.900 803.850 ;
        RECT 604.950 799.950 607.050 802.050 ;
        RECT 614.550 790.050 615.450 811.950 ;
        RECT 622.200 810.000 624.000 818.400 ;
        RECT 647.700 813.600 649.500 818.400 ;
        RECT 667.800 815.400 669.600 818.400 ;
        RECT 644.400 812.400 649.500 813.600 ;
        RECT 620.700 808.800 624.000 810.000 ;
        RECT 634.950 808.950 637.050 811.050 ;
        RECT 620.700 805.050 621.600 808.800 ;
        RECT 619.950 802.950 622.050 805.050 ;
        RECT 620.700 790.800 621.600 802.950 ;
        RECT 623.100 802.050 624.900 803.850 ;
        RECT 625.950 802.950 628.050 805.050 ;
        RECT 622.950 799.950 625.050 802.050 ;
        RECT 626.100 801.150 627.900 802.950 ;
        RECT 629.100 802.050 630.900 803.850 ;
        RECT 628.950 799.950 631.050 802.050 ;
        RECT 601.800 783.600 603.600 789.600 ;
        RECT 613.950 787.950 616.050 790.050 ;
        RECT 620.700 789.900 627.300 790.800 ;
        RECT 635.550 790.050 636.450 808.950 ;
        RECT 644.400 805.050 645.600 812.400 ;
        RECT 658.950 811.950 661.050 814.050 ;
        RECT 643.950 802.950 646.050 805.050 ;
        RECT 637.950 799.950 640.050 802.050 ;
        RECT 638.550 796.050 639.450 799.950 ;
        RECT 637.950 793.950 640.050 796.050 ;
        RECT 644.400 795.600 645.600 802.950 ;
        RECT 647.100 802.050 648.900 803.850 ;
        RECT 649.950 802.950 652.050 805.050 ;
        RECT 646.950 799.950 649.050 802.050 ;
        RECT 650.100 801.150 651.900 802.950 ;
        RECT 653.100 802.050 654.900 803.850 ;
        RECT 652.950 799.950 655.050 802.050 ;
        RECT 659.550 799.050 660.450 811.950 ;
        RECT 668.400 802.050 669.600 815.400 ;
        RECT 683.400 810.600 685.200 818.400 ;
        RECT 690.900 814.200 692.700 818.400 ;
        RECT 703.950 814.950 706.050 817.050 ;
        RECT 690.900 812.400 693.600 814.200 ;
        RECT 689.100 810.600 690.900 811.500 ;
        RECT 683.400 809.700 690.900 810.600 ;
        RECT 683.100 805.050 684.900 806.850 ;
        RECT 670.950 802.950 673.050 805.050 ;
        RECT 682.950 802.950 685.050 805.050 ;
        RECT 658.950 796.950 661.050 799.050 ;
        RECT 667.950 796.950 670.050 802.050 ;
        RECT 671.100 801.150 672.900 802.950 ;
        RECT 620.700 789.600 621.600 789.900 ;
        RECT 619.800 783.600 621.600 789.600 ;
        RECT 625.800 789.600 627.300 789.900 ;
        RECT 625.800 783.600 627.600 789.600 ;
        RECT 634.950 787.950 637.050 790.050 ;
        RECT 643.800 783.600 645.600 795.600 ;
        RECT 646.800 794.700 654.600 795.600 ;
        RECT 646.800 783.600 648.600 794.700 ;
        RECT 652.800 783.600 654.600 794.700 ;
        RECT 668.400 789.600 669.600 796.950 ;
        RECT 667.800 783.600 669.600 789.600 ;
        RECT 686.400 789.600 687.300 809.700 ;
        RECT 692.700 805.050 693.600 812.400 ;
        RECT 700.950 808.950 703.050 811.050 ;
        RECT 688.950 802.950 691.050 805.050 ;
        RECT 691.950 802.950 694.050 805.050 ;
        RECT 689.100 801.150 690.900 802.950 ;
        RECT 692.700 795.600 693.600 802.950 ;
        RECT 686.400 783.600 688.200 789.600 ;
        RECT 692.700 783.600 694.500 795.600 ;
        RECT 701.550 790.050 702.450 808.950 ;
        RECT 700.950 787.950 703.050 790.050 ;
        RECT 704.550 787.050 705.450 814.950 ;
        RECT 712.200 810.000 714.000 818.400 ;
        RECT 724.950 811.950 727.050 814.050 ;
        RECT 710.700 808.800 714.000 810.000 ;
        RECT 710.700 805.050 711.600 808.800 ;
        RECT 709.950 802.950 712.050 805.050 ;
        RECT 710.700 790.800 711.600 802.950 ;
        RECT 713.100 802.050 714.900 803.850 ;
        RECT 715.950 802.950 718.050 805.050 ;
        RECT 712.950 799.950 715.050 802.050 ;
        RECT 716.100 801.150 717.900 802.950 ;
        RECT 719.100 802.050 720.900 803.850 ;
        RECT 718.950 799.950 721.050 802.050 ;
        RECT 710.700 789.900 717.300 790.800 ;
        RECT 710.700 789.600 711.600 789.900 ;
        RECT 703.950 784.950 706.050 787.050 ;
        RECT 709.800 783.600 711.600 789.600 ;
        RECT 715.800 789.600 717.300 789.900 ;
        RECT 715.800 783.600 717.600 789.600 ;
        RECT 725.550 787.050 726.450 811.950 ;
        RECT 736.800 811.200 738.600 818.400 ;
        RECT 742.950 814.950 745.050 817.050 ;
        RECT 734.400 810.300 738.600 811.200 ;
        RECT 734.400 805.050 735.600 810.300 ;
        RECT 731.100 802.050 732.900 803.850 ;
        RECT 733.950 802.950 736.050 805.050 ;
        RECT 730.950 799.950 733.050 802.050 ;
        RECT 734.400 789.600 735.600 802.950 ;
        RECT 737.100 802.050 738.900 803.850 ;
        RECT 736.950 799.950 739.050 802.050 ;
        RECT 743.550 793.050 744.450 814.950 ;
        RECT 758.700 813.600 760.500 818.400 ;
        RECT 755.400 812.400 760.500 813.600 ;
        RECT 755.400 805.050 756.600 812.400 ;
        RECT 779.400 811.200 781.200 818.400 ;
        RECT 799.800 815.400 801.600 818.400 ;
        RECT 779.400 810.300 783.600 811.200 ;
        RECT 782.400 805.050 783.600 810.300 ;
        RECT 754.950 802.950 757.050 805.050 ;
        RECT 755.400 795.600 756.600 802.950 ;
        RECT 758.100 802.050 759.900 803.850 ;
        RECT 760.950 802.950 763.050 805.050 ;
        RECT 757.950 799.950 760.050 802.050 ;
        RECT 761.100 801.150 762.900 802.950 ;
        RECT 764.100 802.050 765.900 803.850 ;
        RECT 779.100 802.050 780.900 803.850 ;
        RECT 781.950 802.950 784.050 805.050 ;
        RECT 763.950 799.950 766.050 802.050 ;
        RECT 778.950 799.950 781.050 802.050 ;
        RECT 742.950 790.950 745.050 793.050 ;
        RECT 724.950 784.950 727.050 787.050 ;
        RECT 734.400 783.600 736.200 789.600 ;
        RECT 754.800 783.600 756.600 795.600 ;
        RECT 757.800 794.700 765.600 795.600 ;
        RECT 757.800 783.600 759.600 794.700 ;
        RECT 763.800 783.600 765.600 794.700 ;
        RECT 782.400 789.600 783.600 802.950 ;
        RECT 785.100 802.050 786.900 803.850 ;
        RECT 800.400 802.050 801.600 815.400 ;
        RECT 815.400 813.300 817.200 818.400 ;
        RECT 821.400 813.300 823.200 818.400 ;
        RECT 815.400 811.950 823.200 813.300 ;
        RECT 824.400 812.400 826.200 818.400 ;
        RECT 839.400 813.300 841.200 818.400 ;
        RECT 845.400 813.300 847.200 818.400 ;
        RECT 824.400 810.300 825.600 812.400 ;
        RECT 839.400 811.950 847.200 813.300 ;
        RECT 848.400 812.400 850.200 818.400 ;
        RECT 860.100 814.950 862.200 817.050 ;
        RECT 868.800 815.400 870.600 818.400 ;
        RECT 848.400 810.300 849.600 812.400 ;
        RECT 821.850 809.250 825.600 810.300 ;
        RECT 845.850 809.250 849.600 810.300 ;
        RECT 821.850 805.050 823.050 809.250 ;
        RECT 845.850 805.050 847.050 809.250 ;
        RECT 802.950 802.950 805.050 805.050 ;
        RECT 814.950 802.950 817.050 805.050 ;
        RECT 784.950 799.950 787.050 802.050 ;
        RECT 793.800 796.950 795.900 799.050 ;
        RECT 799.950 796.950 802.050 802.050 ;
        RECT 803.100 801.150 804.900 802.950 ;
        RECT 815.100 801.150 816.900 802.950 ;
        RECT 818.100 802.050 819.900 803.850 ;
        RECT 820.950 802.950 823.050 805.050 ;
        RECT 817.950 799.950 820.050 802.050 ;
        RECT 781.800 783.600 783.600 789.600 ;
        RECT 794.550 787.050 795.450 796.950 ;
        RECT 800.400 789.600 801.600 796.950 ;
        RECT 820.950 789.600 822.150 802.950 ;
        RECT 824.100 802.050 825.900 803.850 ;
        RECT 838.950 802.950 841.050 805.050 ;
        RECT 823.950 799.950 826.050 802.050 ;
        RECT 839.100 801.150 840.900 802.950 ;
        RECT 842.100 802.050 843.900 803.850 ;
        RECT 844.950 802.950 847.050 805.050 ;
        RECT 841.950 799.950 844.050 802.050 ;
        RECT 844.950 789.600 846.150 802.950 ;
        RECT 848.100 802.050 849.900 803.850 ;
        RECT 847.950 799.950 850.050 802.050 ;
        RECT 790.950 785.550 795.450 787.050 ;
        RECT 790.950 784.950 795.000 785.550 ;
        RECT 799.800 783.600 801.600 789.600 ;
        RECT 820.800 783.600 822.600 789.600 ;
        RECT 844.800 783.600 846.600 789.600 ;
        RECT 860.550 787.050 861.450 814.950 ;
        RECT 865.950 805.950 868.050 808.050 ;
        RECT 866.100 804.150 867.900 805.950 ;
        RECT 869.400 805.050 870.300 815.400 ;
        RECT 889.500 813.600 891.300 818.400 ;
        RECT 901.950 814.950 904.050 817.050 ;
        RECT 889.500 812.400 894.600 813.600 ;
        RECT 871.950 805.950 874.050 808.050 ;
        RECT 868.950 802.950 871.050 805.050 ;
        RECT 872.100 804.150 873.900 805.950 ;
        RECT 893.400 805.050 894.600 812.400 ;
        RECT 898.950 805.950 901.050 808.050 ;
        RECT 869.400 795.600 870.300 802.950 ;
        RECT 884.100 802.050 885.900 803.850 ;
        RECT 886.950 802.950 889.050 805.050 ;
        RECT 883.950 799.950 886.050 802.050 ;
        RECT 887.100 801.150 888.900 802.950 ;
        RECT 890.100 802.050 891.900 803.850 ;
        RECT 892.950 802.950 895.050 805.050 ;
        RECT 889.950 799.950 892.050 802.050 ;
        RECT 893.400 795.600 894.600 802.950 ;
        RECT 866.700 794.400 870.300 795.600 ;
        RECT 884.400 794.700 892.200 795.600 ;
        RECT 859.950 784.950 862.050 787.050 ;
        RECT 866.700 783.600 868.500 794.400 ;
        RECT 884.400 783.600 886.200 794.700 ;
        RECT 890.400 783.600 892.200 794.700 ;
        RECT 893.400 783.600 895.200 795.600 ;
        RECT 899.550 787.050 900.450 805.950 ;
        RECT 902.550 793.050 903.450 814.950 ;
        RECT 901.950 790.950 904.050 793.050 ;
        RECT 898.950 784.950 901.050 787.050 ;
        RECT 13.800 773.400 15.600 779.400 ;
        RECT 32.400 773.400 34.200 779.400 ;
        RECT 14.400 766.050 15.600 773.400 ;
        RECT 32.700 773.100 34.200 773.400 ;
        RECT 38.400 773.400 40.200 779.400 ;
        RECT 59.400 773.400 61.200 779.400 ;
        RECT 79.800 773.400 81.600 779.400 ;
        RECT 38.400 773.100 39.300 773.400 ;
        RECT 32.700 772.200 39.300 773.100 ;
        RECT 13.950 760.950 16.050 766.050 ;
        RECT 14.400 747.600 15.600 760.950 ;
        RECT 17.100 760.050 18.900 761.850 ;
        RECT 28.950 760.950 31.050 763.050 ;
        RECT 16.950 757.950 19.050 760.050 ;
        RECT 29.100 759.150 30.900 760.950 ;
        RECT 32.100 760.050 33.900 761.850 ;
        RECT 34.950 760.950 37.050 763.050 ;
        RECT 31.950 757.950 34.050 760.050 ;
        RECT 35.100 759.150 36.900 760.950 ;
        RECT 38.400 760.050 39.300 772.200 ;
        RECT 55.950 760.950 58.050 763.050 ;
        RECT 37.950 757.950 40.050 760.050 ;
        RECT 56.100 759.150 57.900 760.950 ;
        RECT 59.850 760.050 61.050 773.400 ;
        RECT 80.700 773.100 81.600 773.400 ;
        RECT 85.800 773.400 87.600 779.400 ;
        RECT 103.800 773.400 105.600 779.400 ;
        RECT 85.800 773.100 87.300 773.400 ;
        RECT 80.700 772.200 87.300 773.100 ;
        RECT 104.700 773.100 105.600 773.400 ;
        RECT 109.800 773.400 111.600 779.400 ;
        RECT 109.800 773.100 111.300 773.400 ;
        RECT 104.700 772.200 111.300 773.100 ;
        RECT 61.950 760.950 64.050 763.050 ;
        RECT 58.950 757.950 61.050 760.050 ;
        RECT 62.100 759.150 63.900 760.950 ;
        RECT 65.100 760.050 66.900 761.850 ;
        RECT 80.700 760.050 81.600 772.200 ;
        RECT 97.950 769.950 100.050 772.050 ;
        RECT 82.950 760.950 85.050 763.050 ;
        RECT 64.950 757.950 67.050 760.050 ;
        RECT 79.950 757.950 82.050 760.050 ;
        RECT 83.100 759.150 84.900 760.950 ;
        RECT 86.100 760.050 87.900 761.850 ;
        RECT 88.950 760.950 91.050 763.050 ;
        RECT 85.950 757.950 88.050 760.050 ;
        RECT 89.100 759.150 90.900 760.950 ;
        RECT 38.400 754.200 39.300 757.950 ;
        RECT 13.800 744.600 15.600 747.600 ;
        RECT 36.000 753.000 39.300 754.200 ;
        RECT 58.950 753.750 60.150 757.950 ;
        RECT 36.000 744.600 37.800 753.000 ;
        RECT 56.400 752.700 60.150 753.750 ;
        RECT 80.700 754.200 81.600 757.950 ;
        RECT 80.700 753.000 84.000 754.200 ;
        RECT 56.400 750.600 57.600 752.700 ;
        RECT 55.800 744.600 57.600 750.600 ;
        RECT 58.800 749.700 66.600 751.050 ;
        RECT 58.800 744.600 60.600 749.700 ;
        RECT 64.800 744.600 66.600 749.700 ;
        RECT 82.200 744.600 84.000 753.000 ;
        RECT 98.550 748.050 99.450 769.950 ;
        RECT 104.700 760.050 105.600 772.200 ;
        RECT 125.400 768.300 127.200 779.400 ;
        RECT 131.400 768.300 133.200 779.400 ;
        RECT 125.400 767.400 133.200 768.300 ;
        RECT 134.400 767.400 136.200 779.400 ;
        RECT 151.800 773.400 153.600 779.400 ;
        RECT 152.700 773.100 153.600 773.400 ;
        RECT 157.800 773.400 159.600 779.400 ;
        RECT 157.800 773.100 159.300 773.400 ;
        RECT 152.700 772.200 159.300 773.100 ;
        RECT 106.950 760.950 109.050 763.050 ;
        RECT 103.950 757.950 106.050 760.050 ;
        RECT 107.100 759.150 108.900 760.950 ;
        RECT 110.100 760.050 111.900 761.850 ;
        RECT 112.950 760.950 115.050 763.050 ;
        RECT 124.950 760.950 127.050 763.050 ;
        RECT 109.950 757.950 112.050 760.050 ;
        RECT 113.100 759.150 114.900 760.950 ;
        RECT 118.950 757.950 121.050 760.050 ;
        RECT 125.100 759.150 126.900 760.950 ;
        RECT 128.100 760.050 129.900 761.850 ;
        RECT 130.950 760.950 133.050 763.050 ;
        RECT 127.950 757.950 130.050 760.050 ;
        RECT 131.100 759.150 132.900 760.950 ;
        RECT 134.400 760.050 135.600 767.400 ;
        RECT 152.700 760.050 153.600 772.200 ;
        RECT 175.800 767.400 177.600 779.400 ;
        RECT 178.800 768.300 180.600 779.400 ;
        RECT 184.800 768.300 186.600 779.400 ;
        RECT 200.400 773.400 202.200 779.400 ;
        RECT 210.000 774.450 214.050 775.050 ;
        RECT 188.100 769.950 190.200 772.050 ;
        RECT 178.800 767.400 186.600 768.300 ;
        RECT 154.950 760.950 157.050 763.050 ;
        RECT 133.950 757.950 136.050 760.050 ;
        RECT 145.950 757.950 148.050 760.050 ;
        RECT 151.950 757.950 154.050 760.050 ;
        RECT 155.100 759.150 156.900 760.950 ;
        RECT 158.100 760.050 159.900 761.850 ;
        RECT 160.950 760.950 163.050 763.050 ;
        RECT 157.950 757.950 160.050 760.050 ;
        RECT 161.100 759.150 162.900 760.950 ;
        RECT 176.400 760.050 177.600 767.400 ;
        RECT 188.550 766.050 189.450 769.950 ;
        RECT 187.950 763.950 190.050 766.050 ;
        RECT 178.950 760.950 181.050 763.050 ;
        RECT 169.950 757.950 172.050 760.050 ;
        RECT 175.950 757.950 178.050 760.050 ;
        RECT 179.100 759.150 180.900 760.950 ;
        RECT 182.100 760.050 183.900 761.850 ;
        RECT 184.950 760.950 187.050 763.050 ;
        RECT 196.950 760.950 199.050 763.050 ;
        RECT 181.950 757.950 184.050 760.050 ;
        RECT 185.100 759.150 186.900 760.950 ;
        RECT 197.100 759.150 198.900 760.950 ;
        RECT 200.400 760.050 201.600 773.400 ;
        RECT 209.550 772.950 214.050 774.450 ;
        RECT 224.400 773.400 226.200 779.400 ;
        RECT 202.950 760.950 205.050 763.050 ;
        RECT 199.950 757.950 202.050 760.050 ;
        RECT 203.100 759.150 204.900 760.950 ;
        RECT 104.700 754.200 105.600 757.950 ;
        RECT 104.700 753.000 108.000 754.200 ;
        RECT 97.950 745.950 100.050 748.050 ;
        RECT 106.200 744.600 108.000 753.000 ;
        RECT 119.550 748.050 120.450 757.950 ;
        RECT 134.400 750.600 135.600 757.950 ;
        RECT 130.500 749.400 135.600 750.600 ;
        RECT 119.550 746.550 124.050 748.050 ;
        RECT 120.000 745.950 124.050 746.550 ;
        RECT 130.500 744.600 132.300 749.400 ;
        RECT 146.550 748.050 147.450 757.950 ;
        RECT 152.700 754.200 153.600 757.950 ;
        RECT 152.700 753.000 156.000 754.200 ;
        RECT 145.950 745.950 148.050 748.050 ;
        RECT 154.200 744.600 156.000 753.000 ;
        RECT 170.550 748.050 171.450 757.950 ;
        RECT 176.400 750.600 177.600 757.950 ;
        RECT 200.400 752.700 201.600 757.950 ;
        RECT 200.400 751.800 204.600 752.700 ;
        RECT 176.400 749.400 181.500 750.600 ;
        RECT 169.950 745.950 172.050 748.050 ;
        RECT 179.700 744.600 181.500 749.400 ;
        RECT 202.800 744.600 204.600 751.800 ;
        RECT 209.550 748.050 210.450 772.950 ;
        RECT 220.950 760.950 223.050 763.050 ;
        RECT 221.100 759.150 222.900 760.950 ;
        RECT 224.850 760.050 226.050 773.400 ;
        RECT 235.950 772.950 238.050 775.050 ;
        RECT 226.950 760.950 229.050 763.050 ;
        RECT 223.950 757.950 226.050 760.050 ;
        RECT 227.100 759.150 228.900 760.950 ;
        RECT 230.100 760.050 231.900 761.850 ;
        RECT 229.950 757.950 232.050 760.050 ;
        RECT 223.950 753.750 225.150 757.950 ;
        RECT 236.550 757.050 237.450 772.950 ;
        RECT 244.800 767.400 246.600 779.400 ;
        RECT 262.800 773.400 264.600 779.400 ;
        RECT 245.400 760.050 246.600 767.400 ;
        RECT 263.700 773.100 264.600 773.400 ;
        RECT 268.800 773.400 270.600 779.400 ;
        RECT 268.800 773.100 270.300 773.400 ;
        RECT 263.700 772.200 270.300 773.100 ;
        RECT 247.950 760.950 250.050 763.050 ;
        RECT 244.950 757.950 247.050 760.050 ;
        RECT 248.100 759.150 249.900 760.950 ;
        RECT 263.700 760.050 264.600 772.200 ;
        RECT 284.400 768.300 286.200 779.400 ;
        RECT 290.400 768.300 292.200 779.400 ;
        RECT 284.400 767.400 292.200 768.300 ;
        RECT 293.400 767.400 295.200 779.400 ;
        RECT 311.400 773.400 313.200 779.400 ;
        RECT 311.700 773.100 313.200 773.400 ;
        RECT 317.400 773.400 319.200 779.400 ;
        RECT 338.400 773.400 340.200 779.400 ;
        RECT 317.400 773.100 318.300 773.400 ;
        RECT 311.700 772.200 318.300 773.100 ;
        RECT 265.950 760.950 268.050 763.050 ;
        RECT 262.950 757.950 265.050 760.050 ;
        RECT 266.100 759.150 267.900 760.950 ;
        RECT 269.100 760.050 270.900 761.850 ;
        RECT 271.950 760.950 274.050 763.050 ;
        RECT 283.950 760.950 286.050 763.050 ;
        RECT 268.950 757.950 271.050 760.050 ;
        RECT 272.100 759.150 273.900 760.950 ;
        RECT 284.100 759.150 285.900 760.950 ;
        RECT 287.100 760.050 288.900 761.850 ;
        RECT 289.950 760.950 292.050 763.050 ;
        RECT 286.950 757.950 289.050 760.050 ;
        RECT 290.100 759.150 291.900 760.950 ;
        RECT 293.400 760.050 294.600 767.400 ;
        RECT 307.950 760.950 310.050 763.050 ;
        RECT 292.950 757.950 295.050 760.050 ;
        RECT 308.100 759.150 309.900 760.950 ;
        RECT 311.100 760.050 312.900 761.850 ;
        RECT 313.950 760.950 316.050 763.050 ;
        RECT 310.950 757.950 313.050 760.050 ;
        RECT 314.100 759.150 315.900 760.950 ;
        RECT 317.400 760.050 318.300 772.200 ;
        RECT 334.950 760.950 337.050 763.050 ;
        RECT 316.950 757.950 319.050 760.050 ;
        RECT 335.100 759.150 336.900 760.950 ;
        RECT 338.850 760.050 340.050 773.400 ;
        RECT 358.800 767.400 360.600 779.400 ;
        RECT 361.800 768.300 363.600 779.400 ;
        RECT 367.800 768.300 369.600 779.400 ;
        RECT 376.950 772.950 379.050 775.050 ;
        RECT 382.800 773.400 384.600 779.400 ;
        RECT 383.700 773.100 384.600 773.400 ;
        RECT 388.800 773.400 390.600 779.400 ;
        RECT 406.800 773.400 408.600 779.400 ;
        RECT 388.800 773.100 390.300 773.400 ;
        RECT 361.800 767.400 369.600 768.300 ;
        RECT 340.950 760.950 343.050 763.050 ;
        RECT 337.950 757.950 340.050 760.050 ;
        RECT 341.100 759.150 342.900 760.950 ;
        RECT 344.100 760.050 345.900 761.850 ;
        RECT 359.400 760.050 360.600 767.400 ;
        RECT 361.950 760.950 364.050 763.050 ;
        RECT 343.950 757.950 346.050 760.050 ;
        RECT 358.950 757.950 361.050 760.050 ;
        RECT 362.100 759.150 363.900 760.950 ;
        RECT 365.100 760.050 366.900 761.850 ;
        RECT 367.950 760.950 370.050 763.050 ;
        RECT 364.950 757.950 367.050 760.050 ;
        RECT 368.100 759.150 369.900 760.950 ;
        RECT 235.950 754.950 238.050 757.050 ;
        RECT 221.400 752.700 225.150 753.750 ;
        RECT 221.400 750.600 222.600 752.700 ;
        RECT 208.950 745.950 211.050 748.050 ;
        RECT 220.800 744.600 222.600 750.600 ;
        RECT 223.800 749.700 231.600 751.050 ;
        RECT 245.400 750.600 246.600 757.950 ;
        RECT 263.700 754.200 264.600 757.950 ;
        RECT 263.700 753.000 267.000 754.200 ;
        RECT 223.800 744.600 225.600 749.700 ;
        RECT 229.800 744.600 231.600 749.700 ;
        RECT 244.800 744.600 246.600 750.600 ;
        RECT 265.200 744.600 267.000 753.000 ;
        RECT 293.400 750.600 294.600 757.950 ;
        RECT 317.400 754.200 318.300 757.950 ;
        RECT 289.500 749.400 294.600 750.600 ;
        RECT 315.000 753.000 318.300 754.200 ;
        RECT 337.950 753.750 339.150 757.950 ;
        RECT 289.500 744.600 291.300 749.400 ;
        RECT 315.000 744.600 316.800 753.000 ;
        RECT 335.400 752.700 339.150 753.750 ;
        RECT 335.400 750.600 336.600 752.700 ;
        RECT 334.800 744.600 336.600 750.600 ;
        RECT 337.800 749.700 345.600 751.050 ;
        RECT 337.800 744.600 339.600 749.700 ;
        RECT 343.800 744.600 345.600 749.700 ;
        RECT 359.400 750.600 360.600 757.950 ;
        RECT 370.950 754.950 373.050 757.050 ;
        RECT 371.550 751.050 372.450 754.950 ;
        RECT 377.550 751.050 378.450 772.950 ;
        RECT 383.700 772.200 390.300 773.100 ;
        RECT 407.700 773.100 408.600 773.400 ;
        RECT 412.800 773.400 414.600 779.400 ;
        RECT 431.400 773.400 433.200 779.400 ;
        RECT 412.800 773.100 414.300 773.400 ;
        RECT 407.700 772.200 414.300 773.100 ;
        RECT 431.700 773.100 433.200 773.400 ;
        RECT 437.400 773.400 439.200 779.400 ;
        RECT 457.800 773.400 459.600 779.400 ;
        RECT 469.950 775.950 472.050 778.050 ;
        RECT 437.400 773.100 438.300 773.400 ;
        RECT 431.700 772.200 438.300 773.100 ;
        RECT 383.700 760.050 384.600 772.200 ;
        RECT 385.950 760.950 388.050 763.050 ;
        RECT 382.950 757.950 385.050 760.050 ;
        RECT 386.100 759.150 387.900 760.950 ;
        RECT 389.100 760.050 390.900 761.850 ;
        RECT 391.950 760.950 394.050 763.050 ;
        RECT 388.950 757.950 391.050 760.050 ;
        RECT 392.100 759.150 393.900 760.950 ;
        RECT 407.700 760.050 408.600 772.200 ;
        RECT 409.950 760.950 412.050 763.050 ;
        RECT 396.000 759.450 400.050 760.050 ;
        RECT 395.550 757.950 400.050 759.450 ;
        RECT 406.950 757.950 409.050 760.050 ;
        RECT 410.100 759.150 411.900 760.950 ;
        RECT 413.100 760.050 414.900 761.850 ;
        RECT 415.950 760.950 418.050 763.050 ;
        RECT 427.950 760.950 430.050 763.050 ;
        RECT 412.950 757.950 415.050 760.050 ;
        RECT 416.100 759.150 417.900 760.950 ;
        RECT 428.100 759.150 429.900 760.950 ;
        RECT 431.100 760.050 432.900 761.850 ;
        RECT 433.950 760.950 436.050 763.050 ;
        RECT 430.950 757.950 433.050 760.050 ;
        RECT 434.100 759.150 435.900 760.950 ;
        RECT 437.400 760.050 438.300 772.200 ;
        RECT 452.100 760.050 453.900 761.850 ;
        RECT 454.950 760.950 457.050 763.050 ;
        RECT 436.950 757.950 439.050 760.050 ;
        RECT 451.950 757.950 454.050 760.050 ;
        RECT 455.100 759.150 456.900 760.950 ;
        RECT 457.950 760.050 459.150 773.400 ;
        RECT 466.950 769.950 469.050 772.050 ;
        RECT 460.950 760.950 463.050 763.050 ;
        RECT 457.950 757.950 460.050 760.050 ;
        RECT 461.100 759.150 462.900 760.950 ;
        RECT 463.950 757.950 466.050 760.050 ;
        RECT 383.700 754.200 384.600 757.950 ;
        RECT 383.700 753.000 387.000 754.200 ;
        RECT 395.550 754.050 396.450 757.950 ;
        RECT 407.700 754.200 408.600 757.950 ;
        RECT 437.400 754.200 438.300 757.950 ;
        RECT 359.400 749.400 364.500 750.600 ;
        RECT 362.700 744.600 364.500 749.400 ;
        RECT 370.950 748.950 373.050 751.050 ;
        RECT 376.950 748.950 379.050 751.050 ;
        RECT 385.200 744.600 387.000 753.000 ;
        RECT 394.950 751.950 397.050 754.050 ;
        RECT 407.700 753.000 411.000 754.200 ;
        RECT 409.200 744.600 411.000 753.000 ;
        RECT 435.000 753.000 438.300 754.200 ;
        RECT 458.850 753.750 460.050 757.950 ;
        RECT 464.550 754.050 465.450 757.950 ;
        RECT 435.000 744.600 436.800 753.000 ;
        RECT 458.850 752.700 462.600 753.750 ;
        RECT 452.400 749.700 460.200 751.050 ;
        RECT 452.400 744.600 454.200 749.700 ;
        RECT 458.400 744.600 460.200 749.700 ;
        RECT 461.400 750.600 462.600 752.700 ;
        RECT 463.800 751.950 465.900 754.050 ;
        RECT 461.400 744.600 463.200 750.600 ;
        RECT 467.550 748.050 468.450 769.950 ;
        RECT 470.550 754.050 471.450 775.950 ;
        RECT 476.400 768.300 478.200 779.400 ;
        RECT 482.400 768.300 484.200 779.400 ;
        RECT 476.400 767.400 484.200 768.300 ;
        RECT 485.400 767.400 487.200 779.400 ;
        RECT 493.950 775.950 496.050 778.050 ;
        RECT 490.950 772.950 493.050 775.050 ;
        RECT 475.950 760.950 478.050 763.050 ;
        RECT 476.100 759.150 477.900 760.950 ;
        RECT 479.100 760.050 480.900 761.850 ;
        RECT 481.950 760.950 484.050 763.050 ;
        RECT 478.950 757.950 481.050 760.050 ;
        RECT 482.100 759.150 483.900 760.950 ;
        RECT 485.400 760.050 486.600 767.400 ;
        RECT 484.950 757.950 487.050 760.050 ;
        RECT 469.950 751.950 472.050 754.050 ;
        RECT 485.400 750.600 486.600 757.950 ;
        RECT 491.550 751.050 492.450 772.950 ;
        RECT 494.550 754.050 495.450 775.950 ;
        RECT 496.950 772.950 499.050 775.050 ;
        RECT 506.400 773.400 508.200 779.400 ;
        RECT 497.550 757.050 498.450 772.950 ;
        RECT 502.950 760.950 505.050 763.050 ;
        RECT 503.100 759.150 504.900 760.950 ;
        RECT 506.850 760.050 508.050 773.400 ;
        RECT 526.800 767.400 528.600 779.400 ;
        RECT 538.950 775.950 541.050 778.050 ;
        RECT 508.950 760.950 511.050 763.050 ;
        RECT 505.950 757.950 508.050 760.050 ;
        RECT 509.100 759.150 510.900 760.950 ;
        RECT 512.100 760.050 513.900 761.850 ;
        RECT 527.400 760.050 528.600 767.400 ;
        RECT 529.950 760.950 532.050 763.050 ;
        RECT 511.950 757.950 514.050 760.050 ;
        RECT 526.950 757.950 529.050 760.050 ;
        RECT 530.100 759.150 531.900 760.950 ;
        RECT 496.950 754.950 499.050 757.050 ;
        RECT 493.950 751.950 496.050 754.050 ;
        RECT 505.950 753.750 507.150 757.950 ;
        RECT 503.400 752.700 507.150 753.750 ;
        RECT 481.500 749.400 486.600 750.600 ;
        RECT 466.950 745.950 469.050 748.050 ;
        RECT 481.500 744.600 483.300 749.400 ;
        RECT 490.950 748.950 493.050 751.050 ;
        RECT 503.400 750.600 504.600 752.700 ;
        RECT 502.800 744.600 504.600 750.600 ;
        RECT 505.800 749.700 513.600 751.050 ;
        RECT 527.400 750.600 528.600 757.950 ;
        RECT 539.550 751.050 540.450 775.950 ;
        RECT 544.800 773.400 546.600 779.400 ;
        RECT 545.700 773.100 546.600 773.400 ;
        RECT 550.800 773.400 552.600 779.400 ;
        RECT 550.800 773.100 552.300 773.400 ;
        RECT 545.700 772.200 552.300 773.100 ;
        RECT 545.700 760.050 546.600 772.200 ;
        RECT 566.400 768.300 568.200 779.400 ;
        RECT 572.400 768.300 574.200 779.400 ;
        RECT 566.400 767.400 574.200 768.300 ;
        RECT 575.400 767.400 577.200 779.400 ;
        RECT 596.400 773.400 598.200 779.400 ;
        RECT 619.800 773.400 621.600 779.400 ;
        RECT 641.400 773.400 643.200 779.400 ;
        RECT 559.950 763.950 562.050 766.050 ;
        RECT 547.950 760.950 550.050 763.050 ;
        RECT 544.950 757.950 547.050 760.050 ;
        RECT 548.100 759.150 549.900 760.950 ;
        RECT 551.100 760.050 552.900 761.850 ;
        RECT 553.950 760.950 556.050 763.050 ;
        RECT 550.950 757.950 553.050 760.050 ;
        RECT 554.100 759.150 555.900 760.950 ;
        RECT 545.700 754.200 546.600 757.950 ;
        RECT 545.700 753.000 549.000 754.200 ;
        RECT 560.550 754.050 561.450 763.950 ;
        RECT 565.950 760.950 568.050 763.050 ;
        RECT 566.100 759.150 567.900 760.950 ;
        RECT 569.100 760.050 570.900 761.850 ;
        RECT 571.950 760.950 574.050 763.050 ;
        RECT 568.950 757.950 571.050 760.050 ;
        RECT 572.100 759.150 573.900 760.950 ;
        RECT 575.400 760.050 576.600 767.400 ;
        RECT 592.950 760.950 595.050 763.050 ;
        RECT 574.950 757.950 577.050 760.050 ;
        RECT 593.100 759.150 594.900 760.950 ;
        RECT 596.850 760.050 598.050 773.400 ;
        RECT 598.950 760.950 601.050 763.050 ;
        RECT 595.950 757.950 598.050 760.050 ;
        RECT 599.100 759.150 600.900 760.950 ;
        RECT 602.100 760.050 603.900 761.850 ;
        RECT 616.950 760.950 619.050 763.050 ;
        RECT 601.950 757.950 604.050 760.050 ;
        RECT 617.100 759.150 618.900 760.950 ;
        RECT 620.400 760.050 621.600 773.400 ;
        RECT 622.950 760.950 625.050 763.050 ;
        RECT 637.950 760.950 640.050 763.050 ;
        RECT 619.950 757.950 622.050 760.050 ;
        RECT 623.100 759.150 624.900 760.950 ;
        RECT 638.100 759.150 639.900 760.950 ;
        RECT 641.850 760.050 643.050 773.400 ;
        RECT 652.950 769.950 655.050 772.050 ;
        RECT 643.950 760.950 646.050 763.050 ;
        RECT 640.950 757.950 643.050 760.050 ;
        RECT 644.100 759.150 645.900 760.950 ;
        RECT 647.100 760.050 648.900 761.850 ;
        RECT 646.950 757.950 649.050 760.050 ;
        RECT 505.800 744.600 507.600 749.700 ;
        RECT 511.800 744.600 513.600 749.700 ;
        RECT 526.800 744.600 528.600 750.600 ;
        RECT 538.950 748.950 541.050 751.050 ;
        RECT 547.200 744.600 549.000 753.000 ;
        RECT 559.950 751.950 562.050 754.050 ;
        RECT 575.400 750.600 576.600 757.950 ;
        RECT 595.950 753.750 597.150 757.950 ;
        RECT 593.400 752.700 597.150 753.750 ;
        RECT 620.400 752.700 621.600 757.950 ;
        RECT 640.950 753.750 642.150 757.950 ;
        RECT 593.400 750.600 594.600 752.700 ;
        RECT 617.400 751.800 621.600 752.700 ;
        RECT 638.400 752.700 642.150 753.750 ;
        RECT 571.500 749.400 576.600 750.600 ;
        RECT 571.500 744.600 573.300 749.400 ;
        RECT 592.800 744.600 594.600 750.600 ;
        RECT 595.800 749.700 603.600 751.050 ;
        RECT 595.800 744.600 597.600 749.700 ;
        RECT 601.800 744.600 603.600 749.700 ;
        RECT 617.400 744.600 619.200 751.800 ;
        RECT 638.400 750.600 639.600 752.700 ;
        RECT 637.800 744.600 639.600 750.600 ;
        RECT 640.800 749.700 648.600 751.050 ;
        RECT 640.800 744.600 642.600 749.700 ;
        RECT 646.800 744.600 648.600 749.700 ;
        RECT 653.550 748.050 654.450 769.950 ;
        RECT 664.500 768.600 666.300 779.400 ;
        RECT 662.700 767.400 666.300 768.600 ;
        RECT 662.700 760.050 663.600 767.400 ;
        RECT 673.950 766.950 676.050 769.050 ;
        RECT 684.900 767.400 688.200 779.400 ;
        RECT 709.800 773.400 711.600 779.400 ;
        RECT 659.100 757.050 660.900 758.850 ;
        RECT 661.950 757.950 664.050 760.050 ;
        RECT 658.950 754.950 661.050 757.050 ;
        RECT 652.950 745.950 655.050 748.050 ;
        RECT 662.700 747.600 663.600 757.950 ;
        RECT 665.100 757.050 666.900 758.850 ;
        RECT 664.950 754.950 667.050 757.050 ;
        RECT 674.550 751.050 675.450 766.950 ;
        RECT 680.100 760.050 681.900 761.850 ;
        RECT 682.950 760.950 685.050 763.050 ;
        RECT 679.950 757.950 682.050 760.050 ;
        RECT 683.100 759.150 684.900 760.950 ;
        RECT 686.100 760.050 687.300 767.400 ;
        RECT 710.400 766.050 711.600 773.400 ;
        RECT 725.400 768.300 727.200 779.400 ;
        RECT 731.400 768.300 733.200 779.400 ;
        RECT 725.400 767.400 733.200 768.300 ;
        RECT 734.400 767.400 736.200 779.400 ;
        RECT 739.950 775.950 742.050 778.050 ;
        RECT 688.950 760.950 691.050 763.050 ;
        RECT 685.950 757.950 688.050 760.050 ;
        RECT 689.100 759.150 690.900 760.950 ;
        RECT 692.100 760.050 693.900 761.850 ;
        RECT 709.950 760.950 712.050 766.050 ;
        RECT 691.950 757.950 694.050 760.050 ;
        RECT 685.950 753.300 687.300 757.950 ;
        RECT 685.950 752.100 690.600 753.300 ;
        RECT 673.950 748.950 676.050 751.050 ;
        RECT 680.400 750.000 688.200 750.900 ;
        RECT 689.700 750.600 690.600 752.100 ;
        RECT 662.400 744.600 664.200 747.600 ;
        RECT 680.400 744.600 682.200 750.000 ;
        RECT 686.400 745.500 688.200 750.000 ;
        RECT 689.400 746.400 691.200 750.600 ;
        RECT 692.400 745.500 694.200 750.600 ;
        RECT 710.400 747.600 711.600 760.950 ;
        RECT 713.100 760.050 714.900 761.850 ;
        RECT 724.950 760.950 727.050 763.050 ;
        RECT 712.950 757.950 715.050 760.050 ;
        RECT 725.100 759.150 726.900 760.950 ;
        RECT 728.100 760.050 729.900 761.850 ;
        RECT 730.950 760.950 733.050 763.050 ;
        RECT 727.950 757.950 730.050 760.050 ;
        RECT 731.100 759.150 732.900 760.950 ;
        RECT 734.400 760.050 735.600 767.400 ;
        RECT 733.950 757.950 736.050 760.050 ;
        RECT 734.400 750.600 735.600 757.950 ;
        RECT 740.550 751.050 741.450 775.950 ;
        RECT 751.800 767.400 753.600 779.400 ;
        RECT 752.400 760.050 753.600 767.400 ;
        RECT 770.400 773.400 772.200 779.400 ;
        RECT 793.800 773.400 795.600 779.400 ;
        RECT 817.800 773.400 819.600 779.400 ;
        RECT 826.950 775.950 829.050 778.050 ;
        RECT 754.950 760.950 757.050 763.050 ;
        RECT 766.950 760.950 769.050 763.050 ;
        RECT 751.950 757.950 754.050 760.050 ;
        RECT 755.100 759.150 756.900 760.950 ;
        RECT 767.100 759.150 768.900 760.950 ;
        RECT 770.400 760.050 771.600 773.400 ;
        RECT 772.950 760.950 775.050 763.050 ;
        RECT 769.950 757.950 772.050 760.050 ;
        RECT 773.100 759.150 774.900 760.950 ;
        RECT 788.100 760.050 789.900 761.850 ;
        RECT 790.950 760.950 793.050 763.050 ;
        RECT 787.950 757.950 790.050 760.050 ;
        RECT 791.100 759.150 792.900 760.950 ;
        RECT 793.950 760.050 795.150 773.400 ;
        RECT 808.950 769.950 811.050 772.050 ;
        RECT 796.950 760.950 799.050 763.050 ;
        RECT 793.950 757.950 796.050 760.050 ;
        RECT 797.100 759.150 798.900 760.950 ;
        RECT 686.400 744.600 694.200 745.500 ;
        RECT 709.800 744.600 711.600 747.600 ;
        RECT 730.500 749.400 735.600 750.600 ;
        RECT 730.500 744.600 732.300 749.400 ;
        RECT 739.950 748.950 742.050 751.050 ;
        RECT 752.400 750.600 753.600 757.950 ;
        RECT 770.400 752.700 771.600 757.950 ;
        RECT 794.850 753.750 796.050 757.950 ;
        RECT 794.850 752.700 798.600 753.750 ;
        RECT 770.400 751.800 774.600 752.700 ;
        RECT 751.800 744.600 753.600 750.600 ;
        RECT 772.800 744.600 774.600 751.800 ;
        RECT 788.400 749.700 796.200 751.050 ;
        RECT 788.400 744.600 790.200 749.700 ;
        RECT 794.400 744.600 796.200 749.700 ;
        RECT 797.400 750.600 798.600 752.700 ;
        RECT 797.400 744.600 799.200 750.600 ;
        RECT 809.550 748.050 810.450 769.950 ;
        RECT 814.950 760.950 817.050 763.050 ;
        RECT 815.100 759.150 816.900 760.950 ;
        RECT 818.400 760.050 819.600 773.400 ;
        RECT 820.950 760.950 823.050 763.050 ;
        RECT 817.950 757.950 820.050 760.050 ;
        RECT 821.100 759.150 822.900 760.950 ;
        RECT 818.400 752.700 819.600 757.950 ;
        RECT 827.550 757.050 828.450 775.950 ;
        RECT 833.400 773.400 835.200 779.400 ;
        RECT 833.400 766.500 834.600 773.400 ;
        RECT 839.700 767.400 841.500 779.400 ;
        RECT 859.800 773.400 861.600 779.400 ;
        RECT 878.400 773.400 880.200 779.400 ;
        RECT 833.400 765.600 839.400 766.500 ;
        RECT 837.150 764.700 839.400 765.600 ;
        RECT 833.100 760.050 834.900 761.850 ;
        RECT 832.950 757.950 835.050 760.050 ;
        RECT 827.100 754.950 829.200 757.050 ;
        RECT 815.400 751.800 819.600 752.700 ;
        RECT 837.150 753.300 838.050 764.700 ;
        RECT 840.300 760.050 841.500 767.400 ;
        RECT 854.100 760.050 855.900 761.850 ;
        RECT 856.950 760.950 859.050 763.050 ;
        RECT 838.950 757.950 841.500 760.050 ;
        RECT 853.950 757.950 856.050 760.050 ;
        RECT 857.100 759.150 858.900 760.950 ;
        RECT 859.950 760.050 861.150 773.400 ;
        RECT 878.400 766.500 879.600 773.400 ;
        RECT 884.700 767.400 886.500 779.400 ;
        RECT 895.950 769.950 898.050 772.050 ;
        RECT 878.400 765.600 884.400 766.500 ;
        RECT 882.150 764.700 884.400 765.600 ;
        RECT 862.950 760.950 865.050 763.050 ;
        RECT 859.950 757.950 862.050 760.050 ;
        RECT 863.100 759.150 864.900 760.950 ;
        RECT 878.100 760.050 879.900 761.850 ;
        RECT 877.950 757.950 880.050 760.050 ;
        RECT 837.150 752.400 839.400 753.300 ;
        RECT 808.950 745.950 811.050 748.050 ;
        RECT 815.400 744.600 817.200 751.800 ;
        RECT 833.400 751.500 839.400 752.400 ;
        RECT 833.400 747.600 834.600 751.500 ;
        RECT 840.300 750.600 841.500 757.950 ;
        RECT 860.850 753.750 862.050 757.950 ;
        RECT 860.850 752.700 864.600 753.750 ;
        RECT 833.400 744.600 835.200 747.600 ;
        RECT 839.700 744.600 841.500 750.600 ;
        RECT 854.400 749.700 862.200 751.050 ;
        RECT 854.400 744.600 856.200 749.700 ;
        RECT 860.400 744.600 862.200 749.700 ;
        RECT 863.400 750.600 864.600 752.700 ;
        RECT 882.150 753.300 883.050 764.700 ;
        RECT 885.300 760.050 886.500 767.400 ;
        RECT 896.550 760.050 897.450 769.950 ;
        RECT 904.500 768.600 906.300 779.400 ;
        RECT 902.700 767.400 906.300 768.600 ;
        RECT 902.700 760.050 903.600 767.400 ;
        RECT 883.950 757.950 886.500 760.050 ;
        RECT 892.950 758.550 897.450 760.050 ;
        RECT 892.950 757.950 897.000 758.550 ;
        RECT 882.150 752.400 884.400 753.300 ;
        RECT 878.400 751.500 884.400 752.400 ;
        RECT 863.400 744.600 865.200 750.600 ;
        RECT 878.400 747.600 879.600 751.500 ;
        RECT 885.300 750.600 886.500 757.950 ;
        RECT 899.100 757.050 900.900 758.850 ;
        RECT 901.950 757.950 904.050 760.050 ;
        RECT 898.950 754.950 901.050 757.050 ;
        RECT 878.400 744.600 880.200 747.600 ;
        RECT 884.700 744.600 886.500 750.600 ;
        RECT 902.700 747.600 903.600 757.950 ;
        RECT 905.100 757.050 906.900 758.850 ;
        RECT 904.950 754.950 907.050 757.050 ;
        RECT 902.400 744.600 904.200 747.600 ;
        RECT 13.800 737.400 15.600 740.400 ;
        RECT 14.400 724.050 15.600 737.400 ;
        RECT 29.400 735.300 31.200 740.400 ;
        RECT 35.400 735.300 37.200 740.400 ;
        RECT 29.400 733.950 37.200 735.300 ;
        RECT 38.400 734.400 40.200 740.400 ;
        RECT 58.500 735.600 60.300 740.400 ;
        RECT 79.800 737.400 81.600 740.400 ;
        RECT 58.500 734.400 63.600 735.600 ;
        RECT 38.400 732.300 39.600 734.400 ;
        RECT 35.850 731.250 39.600 732.300 ;
        RECT 35.850 727.050 37.050 731.250 ;
        RECT 62.400 727.050 63.600 734.400 ;
        RECT 67.950 730.950 70.050 733.050 ;
        RECT 16.950 724.950 19.050 727.050 ;
        RECT 28.950 724.950 31.050 727.050 ;
        RECT 13.950 718.950 16.050 724.050 ;
        RECT 17.100 723.150 18.900 724.950 ;
        RECT 29.100 723.150 30.900 724.950 ;
        RECT 32.100 724.050 33.900 725.850 ;
        RECT 34.950 724.950 37.050 727.050 ;
        RECT 31.950 721.950 34.050 724.050 ;
        RECT 14.400 711.600 15.600 718.950 ;
        RECT 34.950 711.600 36.150 724.950 ;
        RECT 38.100 724.050 39.900 725.850 ;
        RECT 53.100 724.050 54.900 725.850 ;
        RECT 55.950 724.950 58.050 727.050 ;
        RECT 37.950 721.950 40.050 724.050 ;
        RECT 52.950 721.950 55.050 724.050 ;
        RECT 56.100 723.150 57.900 724.950 ;
        RECT 59.100 724.050 60.900 725.850 ;
        RECT 61.950 724.950 64.050 727.050 ;
        RECT 58.950 721.950 61.050 724.050 ;
        RECT 62.400 717.600 63.600 724.950 ;
        RECT 53.400 716.700 61.200 717.600 ;
        RECT 13.800 705.600 15.600 711.600 ;
        RECT 34.800 705.600 36.600 711.600 ;
        RECT 53.400 705.600 55.200 716.700 ;
        RECT 59.400 705.600 61.200 716.700 ;
        RECT 62.400 705.600 64.200 717.600 ;
        RECT 68.550 709.050 69.450 730.950 ;
        RECT 80.400 724.050 81.600 737.400 ;
        RECT 97.800 734.400 99.600 740.400 ;
        RECT 98.400 732.300 99.600 734.400 ;
        RECT 100.800 735.300 102.600 740.400 ;
        RECT 106.800 735.300 108.600 740.400 ;
        RECT 100.800 733.950 108.600 735.300 ;
        RECT 119.400 735.300 121.200 740.400 ;
        RECT 125.400 735.300 127.200 740.400 ;
        RECT 119.400 733.950 127.200 735.300 ;
        RECT 128.400 734.400 130.200 740.400 ;
        RECT 143.400 735.300 145.200 740.400 ;
        RECT 149.400 735.300 151.200 740.400 ;
        RECT 128.400 732.300 129.600 734.400 ;
        RECT 143.400 733.950 151.200 735.300 ;
        RECT 152.400 734.400 154.200 740.400 ;
        RECT 172.500 735.600 174.300 740.400 ;
        RECT 194.400 737.400 196.200 740.400 ;
        RECT 215.400 737.400 217.200 740.400 ;
        RECT 172.500 734.400 177.600 735.600 ;
        RECT 152.400 732.300 153.600 734.400 ;
        RECT 98.400 731.250 102.150 732.300 ;
        RECT 88.950 727.950 91.050 730.050 ;
        RECT 82.950 724.950 85.050 727.050 ;
        RECT 79.950 718.950 82.050 724.050 ;
        RECT 83.100 723.150 84.900 724.950 ;
        RECT 80.400 711.600 81.600 718.950 ;
        RECT 89.550 712.050 90.450 727.950 ;
        RECT 100.950 727.050 102.150 731.250 ;
        RECT 125.850 731.250 129.600 732.300 ;
        RECT 149.850 731.250 153.600 732.300 ;
        RECT 125.850 727.050 127.050 731.250 ;
        RECT 149.850 727.050 151.050 731.250 ;
        RECT 176.400 727.050 177.600 734.400 ;
        RECT 190.950 727.950 193.050 730.050 ;
        RECT 98.100 724.050 99.900 725.850 ;
        RECT 100.950 724.950 103.050 727.050 ;
        RECT 97.950 721.950 100.050 724.050 ;
        RECT 67.950 706.950 70.050 709.050 ;
        RECT 79.800 705.600 81.600 711.600 ;
        RECT 88.950 709.950 91.050 712.050 ;
        RECT 101.850 711.600 103.050 724.950 ;
        RECT 104.100 724.050 105.900 725.850 ;
        RECT 106.950 724.950 109.050 727.050 ;
        RECT 118.950 724.950 121.050 727.050 ;
        RECT 103.950 721.950 106.050 724.050 ;
        RECT 107.100 723.150 108.900 724.950 ;
        RECT 119.100 723.150 120.900 724.950 ;
        RECT 122.100 724.050 123.900 725.850 ;
        RECT 124.950 724.950 127.050 727.050 ;
        RECT 121.950 721.950 124.050 724.050 ;
        RECT 124.950 711.600 126.150 724.950 ;
        RECT 128.100 724.050 129.900 725.850 ;
        RECT 142.950 724.950 145.050 727.050 ;
        RECT 127.950 721.950 130.050 724.050 ;
        RECT 143.100 723.150 144.900 724.950 ;
        RECT 146.100 724.050 147.900 725.850 ;
        RECT 148.950 724.950 151.050 727.050 ;
        RECT 145.950 721.950 148.050 724.050 ;
        RECT 148.950 711.600 150.150 724.950 ;
        RECT 152.100 724.050 153.900 725.850 ;
        RECT 167.100 724.050 168.900 725.850 ;
        RECT 169.950 724.950 172.050 727.050 ;
        RECT 151.950 721.950 154.050 724.050 ;
        RECT 166.950 721.950 169.050 724.050 ;
        RECT 170.100 723.150 171.900 724.950 ;
        RECT 173.100 724.050 174.900 725.850 ;
        RECT 175.950 724.950 178.050 727.050 ;
        RECT 191.100 726.150 192.900 727.950 ;
        RECT 194.700 727.050 195.600 737.400 ;
        RECT 196.950 727.950 199.050 730.050 ;
        RECT 193.950 724.950 196.050 727.050 ;
        RECT 197.100 726.150 198.900 727.950 ;
        RECT 211.950 724.950 214.050 727.050 ;
        RECT 172.950 721.950 175.050 724.050 ;
        RECT 176.400 717.600 177.600 724.950 ;
        RECT 181.950 721.950 184.050 724.050 ;
        RECT 167.400 716.700 175.200 717.600 ;
        RECT 101.400 705.600 103.200 711.600 ;
        RECT 124.800 705.600 126.600 711.600 ;
        RECT 148.800 705.600 150.600 711.600 ;
        RECT 167.400 705.600 169.200 716.700 ;
        RECT 173.400 705.600 175.200 716.700 ;
        RECT 176.400 705.600 178.200 717.600 ;
        RECT 182.550 712.050 183.450 721.950 ;
        RECT 194.700 717.600 195.600 724.950 ;
        RECT 212.100 723.150 213.900 724.950 ;
        RECT 215.400 724.050 216.600 737.400 ;
        RECT 235.800 733.200 237.600 740.400 ;
        RECT 247.950 736.950 250.050 739.050 ;
        RECT 233.400 732.300 237.600 733.200 ;
        RECT 233.400 727.050 234.600 732.300 ;
        RECT 230.100 724.050 231.900 725.850 ;
        RECT 232.950 724.950 235.050 727.050 ;
        RECT 214.950 718.950 217.050 724.050 ;
        RECT 229.950 721.950 232.050 724.050 ;
        RECT 194.700 716.400 198.300 717.600 ;
        RECT 181.800 709.950 183.900 712.050 ;
        RECT 196.500 705.600 198.300 716.400 ;
        RECT 215.400 711.600 216.600 718.950 ;
        RECT 233.400 711.600 234.600 724.950 ;
        RECT 236.100 724.050 237.900 725.850 ;
        RECT 235.950 721.950 238.050 724.050 ;
        RECT 248.550 718.050 249.450 736.950 ;
        RECT 253.800 734.400 255.600 740.400 ;
        RECT 254.400 732.300 255.600 734.400 ;
        RECT 256.800 735.300 258.600 740.400 ;
        RECT 262.800 735.300 264.600 740.400 ;
        RECT 256.800 733.950 264.600 735.300 ;
        RECT 280.800 733.200 282.600 740.400 ;
        RECT 298.800 734.400 300.600 740.400 ;
        RECT 278.400 732.300 282.600 733.200 ;
        RECT 299.400 732.300 300.600 734.400 ;
        RECT 301.800 735.300 303.600 740.400 ;
        RECT 307.800 735.300 309.600 740.400 ;
        RECT 301.800 733.950 309.600 735.300 ;
        RECT 313.800 733.950 315.900 736.050 ;
        RECT 254.400 731.250 258.150 732.300 ;
        RECT 256.950 727.050 258.150 731.250 ;
        RECT 278.400 727.050 279.600 732.300 ;
        RECT 299.400 731.250 303.150 732.300 ;
        RECT 292.950 727.950 295.050 730.050 ;
        RECT 254.100 724.050 255.900 725.850 ;
        RECT 256.950 724.950 259.050 727.050 ;
        RECT 253.950 721.950 256.050 724.050 ;
        RECT 244.950 716.550 249.450 718.050 ;
        RECT 244.950 715.950 249.000 716.550 ;
        RECT 257.850 711.600 259.050 724.950 ;
        RECT 260.100 724.050 261.900 725.850 ;
        RECT 262.950 724.950 265.050 727.050 ;
        RECT 259.950 721.950 262.050 724.050 ;
        RECT 263.100 723.150 264.900 724.950 ;
        RECT 275.100 724.050 276.900 725.850 ;
        RECT 277.950 724.950 280.050 727.050 ;
        RECT 274.950 721.950 277.050 724.050 ;
        RECT 278.400 711.600 279.600 724.950 ;
        RECT 281.100 724.050 282.900 725.850 ;
        RECT 280.950 721.950 283.050 724.050 ;
        RECT 215.400 705.600 217.200 711.600 ;
        RECT 233.400 705.600 235.200 711.600 ;
        RECT 257.400 705.600 259.200 711.600 ;
        RECT 278.400 705.600 280.200 711.600 ;
        RECT 293.550 709.050 294.450 727.950 ;
        RECT 301.950 727.050 303.150 731.250 ;
        RECT 314.550 730.050 315.450 733.950 ;
        RECT 325.800 733.200 327.600 740.400 ;
        RECT 346.800 733.200 348.600 740.400 ;
        RECT 323.400 732.300 327.600 733.200 ;
        RECT 344.400 732.300 348.600 733.200 ;
        RECT 362.400 732.600 364.200 740.400 ;
        RECT 369.900 736.200 371.700 740.400 ;
        RECT 376.950 736.950 379.050 739.050 ;
        RECT 369.900 734.400 372.600 736.200 ;
        RECT 368.100 732.600 369.900 733.500 ;
        RECT 313.950 727.950 316.050 730.050 ;
        RECT 323.400 727.050 324.600 732.300 ;
        RECT 344.400 727.050 345.600 732.300 ;
        RECT 362.400 731.700 369.900 732.600 ;
        RECT 362.100 727.050 363.900 728.850 ;
        RECT 299.100 724.050 300.900 725.850 ;
        RECT 301.950 724.950 304.050 727.050 ;
        RECT 298.950 721.950 301.050 724.050 ;
        RECT 302.850 711.600 304.050 724.950 ;
        RECT 305.100 724.050 306.900 725.850 ;
        RECT 307.950 724.950 310.050 727.050 ;
        RECT 304.950 721.950 307.050 724.050 ;
        RECT 308.100 723.150 309.900 724.950 ;
        RECT 320.100 724.050 321.900 725.850 ;
        RECT 322.950 724.950 325.050 727.050 ;
        RECT 319.950 721.950 322.050 724.050 ;
        RECT 323.400 711.600 324.600 724.950 ;
        RECT 326.100 724.050 327.900 725.850 ;
        RECT 331.950 724.950 334.050 727.050 ;
        RECT 325.950 721.950 328.050 724.050 ;
        RECT 292.950 706.950 295.050 709.050 ;
        RECT 302.400 705.600 304.200 711.600 ;
        RECT 323.400 705.600 325.200 711.600 ;
        RECT 332.550 709.050 333.450 724.950 ;
        RECT 341.100 724.050 342.900 725.850 ;
        RECT 343.950 724.950 346.050 727.050 ;
        RECT 340.950 721.950 343.050 724.050 ;
        RECT 344.400 711.600 345.600 724.950 ;
        RECT 347.100 724.050 348.900 725.850 ;
        RECT 361.950 724.950 364.050 727.050 ;
        RECT 346.950 721.950 349.050 724.050 ;
        RECT 365.400 711.600 366.300 731.700 ;
        RECT 371.700 727.050 372.600 734.400 ;
        RECT 377.550 727.050 378.450 736.950 ;
        RECT 393.000 732.000 394.800 740.400 ;
        RECT 415.500 735.600 417.300 740.400 ;
        RECT 437.400 737.400 439.200 740.400 ;
        RECT 415.500 734.400 420.600 735.600 ;
        RECT 393.000 730.800 396.300 732.000 ;
        RECT 395.400 727.050 396.300 730.800 ;
        RECT 400.950 727.950 403.050 730.050 ;
        RECT 367.950 724.950 370.050 727.050 ;
        RECT 370.950 724.950 373.050 727.050 ;
        RECT 376.950 724.950 379.050 727.050 ;
        RECT 368.100 723.150 369.900 724.950 ;
        RECT 371.700 717.600 372.600 724.950 ;
        RECT 386.100 724.050 387.900 725.850 ;
        RECT 388.950 724.950 391.050 727.050 ;
        RECT 385.950 721.950 388.050 724.050 ;
        RECT 389.100 723.150 390.900 724.950 ;
        RECT 392.100 724.050 393.900 725.850 ;
        RECT 394.950 724.950 397.050 727.050 ;
        RECT 391.950 721.950 394.050 724.050 ;
        RECT 331.950 706.950 334.050 709.050 ;
        RECT 344.400 705.600 346.200 711.600 ;
        RECT 365.400 705.600 367.200 711.600 ;
        RECT 371.700 705.600 373.500 717.600 ;
        RECT 395.400 712.800 396.300 724.950 ;
        RECT 401.550 715.050 402.450 727.950 ;
        RECT 419.400 727.050 420.600 734.400 ;
        RECT 424.950 727.950 427.050 730.050 ;
        RECT 410.100 724.050 411.900 725.850 ;
        RECT 412.950 724.950 415.050 727.050 ;
        RECT 409.950 721.950 412.050 724.050 ;
        RECT 413.100 723.150 414.900 724.950 ;
        RECT 416.100 724.050 417.900 725.850 ;
        RECT 418.950 724.950 421.050 727.050 ;
        RECT 415.950 721.950 418.050 724.050 ;
        RECT 419.400 717.600 420.600 724.950 ;
        RECT 410.400 716.700 418.200 717.600 ;
        RECT 400.950 712.950 403.050 715.050 ;
        RECT 389.700 711.900 396.300 712.800 ;
        RECT 389.700 711.600 391.200 711.900 ;
        RECT 389.400 705.600 391.200 711.600 ;
        RECT 395.400 711.600 396.300 711.900 ;
        RECT 395.400 705.600 397.200 711.600 ;
        RECT 410.400 705.600 412.200 716.700 ;
        RECT 416.400 705.600 418.200 716.700 ;
        RECT 419.400 705.600 421.200 717.600 ;
        RECT 425.550 712.050 426.450 727.950 ;
        RECT 433.950 724.950 436.050 727.050 ;
        RECT 434.100 723.150 435.900 724.950 ;
        RECT 437.400 724.050 438.600 737.400 ;
        RECT 455.400 734.400 457.200 740.400 ;
        RECT 470.400 735.300 472.200 740.400 ;
        RECT 476.400 735.300 478.200 740.400 ;
        RECT 455.400 727.050 456.600 734.400 ;
        RECT 470.400 733.950 478.200 735.300 ;
        RECT 479.400 734.400 481.200 740.400 ;
        RECT 479.400 732.300 480.600 734.400 ;
        RECT 499.800 733.200 501.600 740.400 ;
        RECT 515.400 735.300 517.200 740.400 ;
        RECT 521.400 735.300 523.200 740.400 ;
        RECT 515.400 733.950 523.200 735.300 ;
        RECT 524.400 734.400 526.200 740.400 ;
        RECT 543.300 736.200 545.100 740.400 ;
        RECT 476.850 731.250 480.600 732.300 ;
        RECT 497.400 732.300 501.600 733.200 ;
        RECT 524.400 732.300 525.600 734.400 ;
        RECT 532.950 733.950 535.050 736.050 ;
        RECT 542.400 734.400 545.100 736.200 ;
        RECT 476.850 727.050 478.050 731.250 ;
        RECT 497.400 727.050 498.600 732.300 ;
        RECT 521.850 731.250 525.600 732.300 ;
        RECT 521.850 727.050 523.050 731.250 ;
        RECT 529.950 727.950 532.050 730.050 ;
        RECT 452.100 724.050 453.900 725.850 ;
        RECT 454.950 724.950 457.050 727.050 ;
        RECT 469.950 724.950 472.050 727.050 ;
        RECT 436.950 718.950 439.050 724.050 ;
        RECT 451.950 721.950 454.050 724.050 ;
        RECT 424.950 709.950 427.050 712.050 ;
        RECT 437.400 711.600 438.600 718.950 ;
        RECT 455.400 717.600 456.600 724.950 ;
        RECT 470.100 723.150 471.900 724.950 ;
        RECT 473.100 724.050 474.900 725.850 ;
        RECT 475.950 724.950 478.050 727.050 ;
        RECT 472.950 721.950 475.050 724.050 ;
        RECT 437.400 705.600 439.200 711.600 ;
        RECT 455.400 705.600 457.200 717.600 ;
        RECT 475.950 711.600 477.150 724.950 ;
        RECT 479.100 724.050 480.900 725.850 ;
        RECT 494.100 724.050 495.900 725.850 ;
        RECT 496.950 724.950 499.050 727.050 ;
        RECT 478.950 721.950 481.050 724.050 ;
        RECT 493.950 721.950 496.050 724.050 ;
        RECT 497.400 711.600 498.600 724.950 ;
        RECT 500.100 724.050 501.900 725.850 ;
        RECT 514.950 724.950 517.050 727.050 ;
        RECT 499.950 721.950 502.050 724.050 ;
        RECT 515.100 723.150 516.900 724.950 ;
        RECT 518.100 724.050 519.900 725.850 ;
        RECT 520.950 724.950 523.050 727.050 ;
        RECT 517.950 721.950 520.050 724.050 ;
        RECT 520.950 711.600 522.150 724.950 ;
        RECT 524.100 724.050 525.900 725.850 ;
        RECT 523.950 721.950 526.050 724.050 ;
        RECT 475.800 705.600 477.600 711.600 ;
        RECT 497.400 705.600 499.200 711.600 ;
        RECT 520.800 705.600 522.600 711.600 ;
        RECT 530.550 709.050 531.450 727.950 ;
        RECT 533.550 712.050 534.450 733.950 ;
        RECT 542.400 727.050 543.300 734.400 ;
        RECT 545.100 732.600 546.900 733.500 ;
        RECT 550.800 732.600 552.600 740.400 ;
        RECT 567.300 736.200 569.100 740.400 ;
        RECT 545.100 731.700 552.600 732.600 ;
        RECT 566.400 734.400 569.100 736.200 ;
        RECT 541.950 724.950 544.050 727.050 ;
        RECT 544.950 724.950 547.050 727.050 ;
        RECT 542.400 717.600 543.300 724.950 ;
        RECT 545.100 723.150 546.900 724.950 ;
        RECT 532.950 709.950 535.050 712.050 ;
        RECT 529.950 706.950 532.050 709.050 ;
        RECT 541.500 705.600 543.300 717.600 ;
        RECT 548.700 711.600 549.600 731.700 ;
        RECT 551.100 727.050 552.900 728.850 ;
        RECT 566.400 727.050 567.300 734.400 ;
        RECT 569.100 732.600 570.900 733.500 ;
        RECT 574.800 732.600 576.600 740.400 ;
        RECT 589.800 734.400 591.600 740.400 ;
        RECT 569.100 731.700 576.600 732.600 ;
        RECT 590.400 732.300 591.600 734.400 ;
        RECT 592.800 735.300 594.600 740.400 ;
        RECT 598.800 735.300 600.600 740.400 ;
        RECT 592.800 733.950 600.600 735.300 ;
        RECT 611.400 735.300 613.200 740.400 ;
        RECT 617.400 735.300 619.200 740.400 ;
        RECT 611.400 733.950 619.200 735.300 ;
        RECT 620.400 734.400 622.200 740.400 ;
        RECT 628.950 736.950 631.050 739.050 ;
        RECT 620.400 732.300 621.600 734.400 ;
        RECT 550.950 724.950 553.050 727.050 ;
        RECT 565.950 724.950 568.050 727.050 ;
        RECT 568.950 724.950 571.050 727.050 ;
        RECT 566.400 717.600 567.300 724.950 ;
        RECT 569.100 723.150 570.900 724.950 ;
        RECT 547.800 705.600 549.600 711.600 ;
        RECT 565.500 705.600 567.300 717.600 ;
        RECT 572.700 711.600 573.600 731.700 ;
        RECT 590.400 731.250 594.150 732.300 ;
        RECT 575.100 727.050 576.900 728.850 ;
        RECT 583.950 727.950 586.050 730.050 ;
        RECT 574.950 724.950 577.050 727.050 ;
        RECT 571.800 705.600 573.600 711.600 ;
        RECT 584.550 709.050 585.450 727.950 ;
        RECT 592.950 727.050 594.150 731.250 ;
        RECT 617.850 731.250 621.600 732.300 ;
        RECT 617.850 727.050 619.050 731.250 ;
        RECT 590.100 724.050 591.900 725.850 ;
        RECT 592.950 724.950 595.050 727.050 ;
        RECT 589.950 721.950 592.050 724.050 ;
        RECT 593.850 711.600 595.050 724.950 ;
        RECT 596.100 724.050 597.900 725.850 ;
        RECT 598.950 724.950 601.050 727.050 ;
        RECT 610.950 724.950 613.050 727.050 ;
        RECT 595.950 721.950 598.050 724.050 ;
        RECT 599.100 723.150 600.900 724.950 ;
        RECT 611.100 723.150 612.900 724.950 ;
        RECT 614.100 724.050 615.900 725.850 ;
        RECT 616.950 724.950 619.050 727.050 ;
        RECT 613.950 721.950 616.050 724.050 ;
        RECT 616.950 711.600 618.150 724.950 ;
        RECT 620.100 724.050 621.900 725.850 ;
        RECT 619.950 721.950 622.050 724.050 ;
        RECT 629.550 715.050 630.450 736.950 ;
        RECT 634.950 733.950 637.050 736.050 ;
        RECT 635.550 730.050 636.450 733.950 ;
        RECT 638.400 733.200 640.200 740.400 ;
        RECT 649.950 733.950 652.050 736.050 ;
        RECT 658.800 734.400 660.600 740.400 ;
        RECT 638.400 732.300 642.600 733.200 ;
        RECT 634.950 727.950 637.050 730.050 ;
        RECT 641.400 727.050 642.600 732.300 ;
        RECT 638.100 724.050 639.900 725.850 ;
        RECT 640.950 724.950 643.050 727.050 ;
        RECT 637.950 721.950 640.050 724.050 ;
        RECT 628.950 712.950 631.050 715.050 ;
        RECT 641.400 711.600 642.600 724.950 ;
        RECT 644.100 724.050 645.900 725.850 ;
        RECT 643.950 721.950 646.050 724.050 ;
        RECT 583.950 706.950 586.050 709.050 ;
        RECT 593.400 705.600 595.200 711.600 ;
        RECT 616.800 705.600 618.600 711.600 ;
        RECT 640.800 705.600 642.600 711.600 ;
        RECT 650.550 712.050 651.450 733.950 ;
        RECT 659.400 732.300 660.600 734.400 ;
        RECT 661.800 735.300 663.600 740.400 ;
        RECT 667.800 735.300 669.600 740.400 ;
        RECT 661.800 733.950 669.600 735.300 ;
        RECT 683.400 733.200 685.200 740.400 ;
        RECT 694.950 736.950 697.050 739.050 ;
        RECT 683.400 732.300 687.600 733.200 ;
        RECT 659.400 731.250 663.150 732.300 ;
        RECT 661.950 727.050 663.150 731.250 ;
        RECT 686.400 727.050 687.600 732.300 ;
        RECT 659.100 724.050 660.900 725.850 ;
        RECT 661.950 724.950 664.050 727.050 ;
        RECT 658.950 721.950 661.050 724.050 ;
        RECT 650.550 710.550 655.050 712.050 ;
        RECT 662.850 711.600 664.050 724.950 ;
        RECT 665.100 724.050 666.900 725.850 ;
        RECT 667.950 724.950 670.050 727.050 ;
        RECT 664.950 721.950 667.050 724.050 ;
        RECT 668.100 723.150 669.900 724.950 ;
        RECT 683.100 724.050 684.900 725.850 ;
        RECT 685.950 724.950 688.050 727.050 ;
        RECT 682.950 721.950 685.050 724.050 ;
        RECT 686.400 711.600 687.600 724.950 ;
        RECT 689.100 724.050 690.900 725.850 ;
        RECT 688.950 721.950 691.050 724.050 ;
        RECT 695.550 715.050 696.450 736.950 ;
        RECT 701.400 735.300 703.200 740.400 ;
        RECT 707.400 735.300 709.200 740.400 ;
        RECT 701.400 733.950 709.200 735.300 ;
        RECT 710.400 734.400 712.200 740.400 ;
        RECT 715.800 736.950 717.900 739.050 ;
        RECT 728.400 737.400 730.200 740.400 ;
        RECT 710.400 732.300 711.600 734.400 ;
        RECT 707.850 731.250 711.600 732.300 ;
        RECT 707.850 727.050 709.050 731.250 ;
        RECT 700.950 724.950 703.050 727.050 ;
        RECT 701.100 723.150 702.900 724.950 ;
        RECT 704.100 724.050 705.900 725.850 ;
        RECT 706.950 724.950 709.050 727.050 ;
        RECT 703.950 721.950 706.050 724.050 ;
        RECT 694.950 712.950 697.050 715.050 ;
        RECT 706.950 711.600 708.150 724.950 ;
        RECT 710.100 724.050 711.900 725.850 ;
        RECT 716.550 724.050 717.450 736.950 ;
        RECT 724.950 727.950 727.050 730.050 ;
        RECT 725.100 726.150 726.900 727.950 ;
        RECT 728.700 727.050 729.600 737.400 ;
        RECT 746.400 735.300 748.200 740.400 ;
        RECT 752.400 735.300 754.200 740.400 ;
        RECT 746.400 733.950 754.200 735.300 ;
        RECT 755.400 734.400 757.200 740.400 ;
        RECT 755.400 732.300 756.600 734.400 ;
        RECT 775.800 733.200 777.600 740.400 ;
        RECT 781.950 736.950 784.050 739.050 ;
        RECT 752.850 731.250 756.600 732.300 ;
        RECT 773.400 732.300 777.600 733.200 ;
        RECT 730.950 727.950 733.050 730.050 ;
        RECT 727.950 724.950 730.050 727.050 ;
        RECT 731.100 726.150 732.900 727.950 ;
        RECT 752.850 727.050 754.050 731.250 ;
        RECT 763.950 727.950 766.050 730.050 ;
        RECT 745.950 724.950 748.050 727.050 ;
        RECT 709.950 721.950 712.050 724.050 ;
        RECT 715.950 721.950 718.050 724.050 ;
        RECT 728.700 717.600 729.600 724.950 ;
        RECT 746.100 723.150 747.900 724.950 ;
        RECT 749.100 724.050 750.900 725.850 ;
        RECT 751.950 724.950 754.050 727.050 ;
        RECT 748.950 721.950 751.050 724.050 ;
        RECT 728.700 716.400 732.300 717.600 ;
        RECT 651.000 709.950 655.050 710.550 ;
        RECT 662.400 705.600 664.200 711.600 ;
        RECT 685.800 705.600 687.600 711.600 ;
        RECT 706.800 705.600 708.600 711.600 ;
        RECT 730.500 705.600 732.300 716.400 ;
        RECT 751.950 711.600 753.150 724.950 ;
        RECT 755.100 724.050 756.900 725.850 ;
        RECT 754.950 721.950 757.050 724.050 ;
        RECT 760.950 718.950 763.050 721.050 ;
        RECT 751.800 705.600 753.600 711.600 ;
        RECT 761.550 709.050 762.450 718.950 ;
        RECT 764.550 709.050 765.450 727.950 ;
        RECT 773.400 727.050 774.600 732.300 ;
        RECT 770.100 724.050 771.900 725.850 ;
        RECT 772.950 724.950 775.050 727.050 ;
        RECT 769.950 721.950 772.050 724.050 ;
        RECT 773.400 711.600 774.600 724.950 ;
        RECT 776.100 724.050 777.900 725.850 ;
        RECT 775.950 721.950 778.050 724.050 ;
        RECT 782.550 715.050 783.450 736.950 ;
        RECT 796.800 733.200 798.600 740.400 ;
        RECT 802.950 736.950 805.050 739.050 ;
        RECT 794.400 732.300 798.600 733.200 ;
        RECT 794.400 727.050 795.600 732.300 ;
        RECT 791.100 724.050 792.900 725.850 ;
        RECT 793.950 724.950 796.050 727.050 ;
        RECT 790.950 721.950 793.050 724.050 ;
        RECT 781.800 712.950 783.900 715.050 ;
        RECT 794.400 711.600 795.600 724.950 ;
        RECT 797.100 724.050 798.900 725.850 ;
        RECT 796.950 721.950 799.050 724.050 ;
        RECT 760.800 706.950 762.900 709.050 ;
        RECT 764.100 706.950 766.200 709.050 ;
        RECT 773.400 705.600 775.200 711.600 ;
        RECT 794.400 705.600 796.200 711.600 ;
        RECT 803.550 709.050 804.450 736.950 ;
        RECT 814.800 734.400 816.600 740.400 ;
        RECT 815.400 727.050 816.600 734.400 ;
        RECT 833.400 737.400 835.200 740.400 ;
        RECT 848.400 737.400 850.200 740.400 ;
        RECT 814.950 724.950 817.050 727.050 ;
        RECT 815.400 717.600 816.600 724.950 ;
        RECT 818.100 724.050 819.900 725.850 ;
        RECT 829.950 724.950 832.050 727.050 ;
        RECT 817.950 721.950 820.050 724.050 ;
        RECT 830.100 723.150 831.900 724.950 ;
        RECT 833.400 724.050 834.600 737.400 ;
        RECT 848.400 733.500 849.600 737.400 ;
        RECT 854.700 734.400 856.500 740.400 ;
        RECT 848.400 732.600 854.400 733.500 ;
        RECT 852.150 731.700 854.400 732.600 ;
        RECT 847.950 724.950 850.050 727.050 ;
        RECT 832.950 718.950 835.050 724.050 ;
        RECT 848.100 723.150 849.900 724.950 ;
        RECT 852.150 720.300 853.050 731.700 ;
        RECT 855.300 727.050 856.500 734.400 ;
        RECT 874.800 733.200 876.600 740.400 ;
        RECT 886.950 736.950 889.050 739.050 ;
        RECT 872.400 732.300 876.600 733.200 ;
        RECT 872.400 727.050 873.600 732.300 ;
        RECT 883.950 730.950 886.050 733.050 ;
        RECT 853.950 724.950 856.500 727.050 ;
        RECT 852.150 719.400 854.400 720.300 ;
        RECT 802.950 706.950 805.050 709.050 ;
        RECT 814.800 705.600 816.600 717.600 ;
        RECT 833.400 711.600 834.600 718.950 ;
        RECT 848.400 718.500 854.400 719.400 ;
        RECT 848.400 711.600 849.600 718.500 ;
        RECT 855.300 717.600 856.500 724.950 ;
        RECT 869.100 724.050 870.900 725.850 ;
        RECT 871.950 724.950 874.050 727.050 ;
        RECT 868.950 721.950 871.050 724.050 ;
        RECT 833.400 705.600 835.200 711.600 ;
        RECT 848.400 705.600 850.200 711.600 ;
        RECT 854.700 705.600 856.500 717.600 ;
        RECT 872.400 711.600 873.600 724.950 ;
        RECT 875.100 724.050 876.900 725.850 ;
        RECT 874.950 721.950 877.050 724.050 ;
        RECT 884.550 712.050 885.450 730.950 ;
        RECT 887.550 727.050 888.450 736.950 ;
        RECT 897.000 732.000 898.800 740.400 ;
        RECT 904.950 736.950 907.050 739.050 ;
        RECT 897.000 730.800 900.300 732.000 ;
        RECT 899.400 727.050 900.300 730.800 ;
        RECT 886.950 724.950 889.050 727.050 ;
        RECT 890.100 724.050 891.900 725.850 ;
        RECT 892.950 724.950 895.050 727.050 ;
        RECT 889.950 721.950 892.050 724.050 ;
        RECT 893.100 723.150 894.900 724.950 ;
        RECT 896.100 724.050 897.900 725.850 ;
        RECT 898.950 724.950 901.050 727.050 ;
        RECT 895.950 721.950 898.050 724.050 ;
        RECT 899.400 712.800 900.300 724.950 ;
        RECT 905.550 724.050 906.450 736.950 ;
        RECT 907.950 733.950 910.050 736.050 ;
        RECT 904.800 721.950 906.900 724.050 ;
        RECT 872.400 705.600 874.200 711.600 ;
        RECT 883.950 709.950 886.050 712.050 ;
        RECT 893.700 711.900 900.300 712.800 ;
        RECT 908.550 712.050 909.450 733.950 ;
        RECT 893.700 711.600 895.200 711.900 ;
        RECT 893.400 705.600 895.200 711.600 ;
        RECT 899.400 711.600 900.300 711.900 ;
        RECT 899.400 705.600 901.200 711.600 ;
        RECT 908.100 709.950 910.200 712.050 ;
        RECT 13.800 695.400 15.600 701.400 ;
        RECT 31.800 695.400 33.600 701.400 ;
        RECT 14.400 688.050 15.600 695.400 ;
        RECT 32.700 695.100 33.600 695.400 ;
        RECT 37.800 695.400 39.600 701.400 ;
        RECT 55.800 695.400 57.600 701.400 ;
        RECT 37.800 695.100 39.300 695.400 ;
        RECT 32.700 694.200 39.300 695.100 ;
        RECT 56.700 695.100 57.600 695.400 ;
        RECT 61.800 695.400 63.600 701.400 ;
        RECT 79.800 695.400 81.600 701.400 ;
        RECT 90.000 696.450 93.900 697.050 ;
        RECT 61.800 695.100 63.300 695.400 ;
        RECT 56.700 694.200 63.300 695.100 ;
        RECT 13.950 682.950 16.050 688.050 ;
        RECT 14.400 669.600 15.600 682.950 ;
        RECT 17.100 682.050 18.900 683.850 ;
        RECT 32.700 682.050 33.600 694.200 ;
        RECT 34.950 682.950 37.050 685.050 ;
        RECT 16.950 679.950 19.050 682.050 ;
        RECT 31.950 679.950 34.050 682.050 ;
        RECT 35.100 681.150 36.900 682.950 ;
        RECT 38.100 682.050 39.900 683.850 ;
        RECT 40.950 682.950 43.050 685.050 ;
        RECT 37.950 679.950 40.050 682.050 ;
        RECT 41.100 681.150 42.900 682.950 ;
        RECT 56.700 682.050 57.600 694.200 ;
        RECT 80.400 688.050 81.600 695.400 ;
        RECT 89.550 694.950 93.900 696.450 ;
        RECT 97.800 695.400 99.600 701.400 ;
        RECT 98.700 695.100 99.600 695.400 ;
        RECT 103.800 695.400 105.600 701.400 ;
        RECT 124.800 695.400 126.600 701.400 ;
        RECT 103.800 695.100 105.300 695.400 ;
        RECT 58.950 682.950 61.050 685.050 ;
        RECT 55.950 679.950 58.050 682.050 ;
        RECT 59.100 681.150 60.900 682.950 ;
        RECT 62.100 682.050 63.900 683.850 ;
        RECT 64.950 682.950 67.050 685.050 ;
        RECT 79.950 682.950 82.050 688.050 ;
        RECT 61.950 679.950 64.050 682.050 ;
        RECT 65.100 681.150 66.900 682.950 ;
        RECT 32.700 676.200 33.600 679.950 ;
        RECT 56.700 676.200 57.600 679.950 ;
        RECT 32.700 675.000 36.000 676.200 ;
        RECT 56.700 675.000 60.000 676.200 ;
        RECT 13.800 666.600 15.600 669.600 ;
        RECT 34.200 666.600 36.000 675.000 ;
        RECT 58.200 666.600 60.000 675.000 ;
        RECT 80.400 669.600 81.600 682.950 ;
        RECT 83.100 682.050 84.900 683.850 ;
        RECT 82.950 679.950 85.050 682.050 ;
        RECT 89.550 673.050 90.450 694.950 ;
        RECT 98.700 694.200 105.300 695.100 ;
        RECT 98.700 682.050 99.600 694.200 ;
        RECT 100.950 682.950 103.050 685.050 ;
        RECT 97.950 679.950 100.050 682.050 ;
        RECT 101.100 681.150 102.900 682.950 ;
        RECT 104.100 682.050 105.900 683.850 ;
        RECT 106.950 682.950 109.050 685.050 ;
        RECT 103.950 679.950 106.050 682.050 ;
        RECT 107.100 681.150 108.900 682.950 ;
        RECT 119.100 682.050 120.900 683.850 ;
        RECT 121.950 682.950 124.050 685.050 ;
        RECT 118.950 679.950 121.050 682.050 ;
        RECT 122.100 681.150 123.900 682.950 ;
        RECT 124.950 682.050 126.150 695.400 ;
        RECT 143.400 690.600 145.200 701.400 ;
        RECT 149.400 700.500 157.200 701.400 ;
        RECT 149.400 690.600 151.200 700.500 ;
        RECT 143.400 689.700 151.200 690.600 ;
        RECT 152.400 688.500 154.200 699.600 ;
        RECT 155.400 689.400 157.200 700.500 ;
        RECT 175.800 695.400 177.600 701.400 ;
        RECT 149.100 687.600 154.200 688.500 ;
        RECT 127.950 682.950 130.050 685.050 ;
        RECT 124.950 679.950 127.050 682.050 ;
        RECT 128.100 681.150 129.900 682.950 ;
        RECT 149.100 682.050 150.000 687.600 ;
        RECT 160.950 685.950 163.050 688.050 ;
        RECT 142.950 679.950 145.050 682.050 ;
        RECT 98.700 676.200 99.600 679.950 ;
        RECT 98.700 675.000 102.000 676.200 ;
        RECT 88.950 670.950 91.050 673.050 ;
        RECT 79.800 666.600 81.600 669.600 ;
        RECT 100.200 666.600 102.000 675.000 ;
        RECT 125.850 675.750 127.050 679.950 ;
        RECT 143.100 678.150 144.900 679.950 ;
        RECT 146.100 679.050 147.900 680.850 ;
        RECT 148.950 679.950 151.050 682.050 ;
        RECT 145.950 676.950 148.050 679.050 ;
        RECT 125.850 674.700 129.600 675.750 ;
        RECT 119.400 671.700 127.200 673.050 ;
        RECT 119.400 666.600 121.200 671.700 ;
        RECT 125.400 666.600 127.200 671.700 ;
        RECT 128.400 672.600 129.600 674.700 ;
        RECT 148.950 672.600 150.000 679.950 ;
        RECT 152.100 679.050 153.900 680.850 ;
        RECT 154.950 679.950 157.050 682.050 ;
        RECT 151.950 676.950 154.050 679.050 ;
        RECT 155.100 678.150 156.900 679.950 ;
        RECT 161.550 679.050 162.450 685.950 ;
        RECT 172.950 682.950 175.050 685.050 ;
        RECT 173.100 681.150 174.900 682.950 ;
        RECT 176.400 682.050 177.600 695.400 ;
        RECT 184.950 694.950 187.050 697.050 ;
        RECT 197.400 695.400 199.200 701.400 ;
        RECT 220.800 695.400 222.600 701.400 ;
        RECT 242.400 695.400 244.200 701.400 ;
        RECT 262.800 695.400 264.600 701.400 ;
        RECT 281.400 695.400 283.200 701.400 ;
        RECT 178.950 682.950 181.050 685.050 ;
        RECT 175.950 679.950 178.050 682.050 ;
        RECT 179.100 681.150 180.900 682.950 ;
        RECT 160.950 676.950 163.050 679.050 ;
        RECT 176.400 674.700 177.600 679.950 ;
        RECT 128.400 666.600 130.200 672.600 ;
        RECT 148.200 666.600 150.000 672.600 ;
        RECT 173.400 673.800 177.600 674.700 ;
        RECT 173.400 666.600 175.200 673.800 ;
        RECT 185.550 670.050 186.450 694.950 ;
        RECT 193.950 682.950 196.050 685.050 ;
        RECT 194.100 681.150 195.900 682.950 ;
        RECT 197.850 682.050 199.050 695.400 ;
        RECT 199.950 682.950 202.050 685.050 ;
        RECT 196.950 679.950 199.050 682.050 ;
        RECT 200.100 681.150 201.900 682.950 ;
        RECT 203.100 682.050 204.900 683.850 ;
        RECT 215.100 682.050 216.900 683.850 ;
        RECT 217.950 682.950 220.050 685.050 ;
        RECT 202.950 679.950 205.050 682.050 ;
        RECT 214.950 679.950 217.050 682.050 ;
        RECT 218.100 681.150 219.900 682.950 ;
        RECT 220.950 682.050 222.150 695.400 ;
        RECT 232.950 691.950 235.050 694.050 ;
        RECT 233.550 688.050 234.450 691.950 ;
        RECT 232.950 685.950 235.050 688.050 ;
        RECT 223.950 682.950 226.050 685.050 ;
        RECT 220.950 679.950 223.050 682.050 ;
        RECT 224.100 681.150 225.900 682.950 ;
        RECT 196.950 675.750 198.150 679.950 ;
        RECT 194.400 674.700 198.150 675.750 ;
        RECT 221.850 675.750 223.050 679.950 ;
        RECT 221.850 674.700 225.600 675.750 ;
        RECT 194.400 672.600 195.600 674.700 ;
        RECT 184.950 667.950 187.050 670.050 ;
        RECT 193.800 666.600 195.600 672.600 ;
        RECT 196.800 671.700 204.600 673.050 ;
        RECT 196.800 666.600 198.600 671.700 ;
        RECT 202.800 666.600 204.600 671.700 ;
        RECT 215.400 671.700 223.200 673.050 ;
        RECT 215.400 666.600 217.200 671.700 ;
        RECT 221.400 666.600 223.200 671.700 ;
        RECT 224.400 672.600 225.600 674.700 ;
        RECT 233.550 673.050 234.450 685.950 ;
        RECT 238.950 682.950 241.050 685.050 ;
        RECT 239.100 681.150 240.900 682.950 ;
        RECT 242.400 682.050 243.600 695.400 ;
        RECT 250.950 691.950 253.050 694.050 ;
        RECT 244.950 682.950 247.050 685.050 ;
        RECT 241.950 679.950 244.050 682.050 ;
        RECT 245.100 681.150 246.900 682.950 ;
        RECT 242.400 674.700 243.600 679.950 ;
        RECT 242.400 673.800 246.600 674.700 ;
        RECT 224.400 666.600 226.200 672.600 ;
        RECT 232.950 670.950 235.050 673.050 ;
        RECT 244.800 666.600 246.600 673.800 ;
        RECT 251.550 670.050 252.450 691.950 ;
        RECT 263.400 688.050 264.600 695.400 ;
        RECT 281.700 695.100 283.200 695.400 ;
        RECT 287.400 695.400 289.200 701.400 ;
        RECT 305.400 695.400 307.200 701.400 ;
        RECT 287.400 695.100 288.300 695.400 ;
        RECT 281.700 694.200 288.300 695.100 ;
        RECT 305.700 695.100 307.200 695.400 ;
        RECT 311.400 695.400 313.200 701.400 ;
        RECT 311.400 695.100 312.300 695.400 ;
        RECT 305.700 694.200 312.300 695.100 ;
        RECT 316.950 694.950 319.050 697.050 ;
        RECT 331.800 695.400 333.600 701.400 ;
        RECT 343.800 697.950 345.900 700.050 ;
        RECT 262.950 682.950 265.050 688.050 ;
        RECT 250.950 667.950 253.050 670.050 ;
        RECT 263.400 669.600 264.600 682.950 ;
        RECT 266.100 682.050 267.900 683.850 ;
        RECT 277.950 682.950 280.050 685.050 ;
        RECT 265.950 679.950 268.050 682.050 ;
        RECT 278.100 681.150 279.900 682.950 ;
        RECT 281.100 682.050 282.900 683.850 ;
        RECT 283.950 682.950 286.050 685.050 ;
        RECT 280.950 679.950 283.050 682.050 ;
        RECT 284.100 681.150 285.900 682.950 ;
        RECT 287.400 682.050 288.300 694.200 ;
        RECT 301.950 682.950 304.050 685.050 ;
        RECT 286.950 679.950 289.050 682.050 ;
        RECT 302.100 681.150 303.900 682.950 ;
        RECT 305.100 682.050 306.900 683.850 ;
        RECT 307.950 682.950 310.050 685.050 ;
        RECT 304.950 679.950 307.050 682.050 ;
        RECT 308.100 681.150 309.900 682.950 ;
        RECT 311.400 682.050 312.300 694.200 ;
        RECT 310.950 679.950 313.050 682.050 ;
        RECT 287.400 676.200 288.300 679.950 ;
        RECT 298.950 676.950 301.050 679.050 ;
        RECT 262.800 666.600 264.600 669.600 ;
        RECT 285.000 675.000 288.300 676.200 ;
        RECT 285.000 666.600 286.800 675.000 ;
        RECT 299.550 670.050 300.450 676.950 ;
        RECT 311.400 676.200 312.300 679.950 ;
        RECT 317.550 678.450 318.450 694.950 ;
        RECT 326.100 682.050 327.900 683.850 ;
        RECT 328.950 682.950 331.050 685.050 ;
        RECT 325.950 679.950 328.050 682.050 ;
        RECT 329.100 681.150 330.900 682.950 ;
        RECT 331.950 682.050 333.150 695.400 ;
        RECT 337.800 694.950 339.900 697.050 ;
        RECT 338.550 691.050 339.450 694.950 ;
        RECT 338.550 689.550 343.050 691.050 ;
        RECT 339.000 688.950 343.050 689.550 ;
        RECT 334.950 682.950 337.050 685.050 ;
        RECT 331.950 679.950 334.050 682.050 ;
        RECT 335.100 681.150 336.900 682.950 ;
        RECT 309.000 675.000 312.300 676.200 ;
        RECT 314.550 677.550 318.450 678.450 ;
        RECT 298.950 667.950 301.050 670.050 ;
        RECT 309.000 666.600 310.800 675.000 ;
        RECT 314.550 670.050 315.450 677.550 ;
        RECT 332.850 675.750 334.050 679.950 ;
        RECT 344.550 679.050 345.450 697.950 ;
        RECT 353.400 695.400 355.200 701.400 ;
        RECT 374.400 695.400 376.200 701.400 ;
        RECT 397.800 695.400 399.600 701.400 ;
        RECT 404.550 699.000 411.450 699.450 ;
        RECT 403.950 698.550 411.450 699.000 ;
        RECT 403.950 697.050 406.050 698.550 ;
        RECT 403.800 696.000 406.050 697.050 ;
        RECT 349.950 682.950 352.050 685.050 ;
        RECT 350.100 681.150 351.900 682.950 ;
        RECT 353.400 682.050 354.600 695.400 ;
        RECT 361.950 691.950 364.050 694.050 ;
        RECT 355.950 682.950 358.050 685.050 ;
        RECT 352.950 679.950 355.050 682.050 ;
        RECT 356.100 681.150 357.900 682.950 ;
        RECT 343.950 676.950 346.050 679.050 ;
        RECT 332.850 674.700 336.600 675.750 ;
        RECT 326.400 671.700 334.200 673.050 ;
        RECT 313.800 667.950 315.900 670.050 ;
        RECT 326.400 666.600 328.200 671.700 ;
        RECT 332.400 666.600 334.200 671.700 ;
        RECT 335.400 672.600 336.600 674.700 ;
        RECT 335.400 666.600 337.200 672.600 ;
        RECT 344.550 670.050 345.450 676.950 ;
        RECT 353.400 674.700 354.600 679.950 ;
        RECT 353.400 673.800 357.600 674.700 ;
        RECT 344.550 668.550 349.050 670.050 ;
        RECT 345.000 667.950 349.050 668.550 ;
        RECT 355.800 666.600 357.600 673.800 ;
        RECT 362.550 670.050 363.450 691.950 ;
        RECT 370.950 682.950 373.050 685.050 ;
        RECT 371.100 681.150 372.900 682.950 ;
        RECT 374.400 682.050 375.600 695.400 ;
        RECT 376.950 682.950 379.050 685.050 ;
        RECT 373.950 679.950 376.050 682.050 ;
        RECT 377.100 681.150 378.900 682.950 ;
        RECT 392.100 682.050 393.900 683.850 ;
        RECT 394.950 682.950 397.050 685.050 ;
        RECT 391.950 679.950 394.050 682.050 ;
        RECT 395.100 681.150 396.900 682.950 ;
        RECT 397.950 682.050 399.150 695.400 ;
        RECT 403.800 694.950 405.900 696.000 ;
        RECT 407.100 694.950 409.200 697.050 ;
        RECT 400.950 682.950 403.050 685.050 ;
        RECT 397.950 679.950 400.050 682.050 ;
        RECT 401.100 681.150 402.900 682.950 ;
        RECT 374.400 674.700 375.600 679.950 ;
        RECT 398.850 675.750 400.050 679.950 ;
        RECT 398.850 674.700 402.600 675.750 ;
        RECT 374.400 673.800 378.600 674.700 ;
        RECT 361.950 667.950 364.050 670.050 ;
        RECT 376.800 666.600 378.600 673.800 ;
        RECT 392.400 671.700 400.200 673.050 ;
        RECT 392.400 666.600 394.200 671.700 ;
        RECT 398.400 666.600 400.200 671.700 ;
        RECT 401.400 672.600 402.600 674.700 ;
        RECT 401.400 666.600 403.200 672.600 ;
        RECT 407.550 670.050 408.450 694.950 ;
        RECT 410.550 694.050 411.450 698.550 ;
        RECT 418.800 695.400 420.600 701.400 ;
        RECT 410.100 691.950 412.200 694.050 ;
        RECT 419.400 688.050 420.600 695.400 ;
        RECT 437.400 695.400 439.200 701.400 ;
        RECT 458.400 695.400 460.200 701.400 ;
        RECT 427.950 690.450 432.000 691.050 ;
        RECT 427.950 690.000 432.450 690.450 ;
        RECT 427.950 688.950 433.050 690.000 ;
        RECT 418.950 682.950 421.050 688.050 ;
        RECT 430.950 685.950 433.050 688.950 ;
        RECT 412.950 676.950 415.050 679.050 ;
        RECT 413.550 670.050 414.450 676.950 ;
        RECT 406.950 667.950 409.050 670.050 ;
        RECT 412.950 667.950 415.050 670.050 ;
        RECT 419.400 669.600 420.600 682.950 ;
        RECT 422.100 682.050 423.900 683.850 ;
        RECT 427.950 682.950 430.050 685.050 ;
        RECT 433.950 682.950 436.050 685.050 ;
        RECT 421.950 679.950 424.050 682.050 ;
        RECT 428.550 676.050 429.450 682.950 ;
        RECT 434.100 681.150 435.900 682.950 ;
        RECT 437.400 682.050 438.600 695.400 ;
        RECT 458.700 695.100 460.200 695.400 ;
        RECT 464.400 695.400 466.200 701.400 ;
        RECT 464.400 695.100 465.300 695.400 ;
        RECT 458.700 694.200 465.300 695.100 ;
        RECT 448.950 691.950 451.050 694.050 ;
        RECT 439.950 682.950 442.050 685.050 ;
        RECT 436.950 679.950 439.050 682.050 ;
        RECT 440.100 681.150 441.900 682.950 ;
        RECT 428.550 674.550 433.050 676.050 ;
        RECT 429.000 673.950 433.050 674.550 ;
        RECT 437.400 674.700 438.600 679.950 ;
        RECT 437.400 673.800 441.600 674.700 ;
        RECT 418.800 666.600 420.600 669.600 ;
        RECT 439.800 666.600 441.600 673.800 ;
        RECT 449.550 670.050 450.450 691.950 ;
        RECT 454.950 682.950 457.050 685.050 ;
        RECT 455.100 681.150 456.900 682.950 ;
        RECT 458.100 682.050 459.900 683.850 ;
        RECT 460.950 682.950 463.050 685.050 ;
        RECT 457.950 679.950 460.050 682.050 ;
        RECT 461.100 681.150 462.900 682.950 ;
        RECT 464.400 682.050 465.300 694.200 ;
        RECT 481.800 689.400 483.600 701.400 ;
        RECT 499.800 689.400 501.600 701.400 ;
        RECT 517.800 689.400 519.600 701.400 ;
        RECT 526.950 697.950 529.050 700.050 ;
        RECT 482.400 682.050 483.600 689.400 ;
        RECT 484.950 682.950 487.050 685.050 ;
        RECT 463.950 679.950 466.050 682.050 ;
        RECT 481.950 679.950 484.050 682.050 ;
        RECT 485.100 681.150 486.900 682.950 ;
        RECT 500.400 682.050 501.600 689.400 ;
        RECT 502.950 682.950 505.050 685.050 ;
        RECT 499.950 679.950 502.050 682.050 ;
        RECT 503.100 681.150 504.900 682.950 ;
        RECT 518.400 682.050 519.600 689.400 ;
        RECT 520.950 682.950 523.050 685.050 ;
        RECT 517.950 679.950 520.050 682.050 ;
        RECT 521.100 681.150 522.900 682.950 ;
        RECT 523.950 679.950 526.050 682.050 ;
        RECT 464.400 676.200 465.300 679.950 ;
        RECT 462.000 675.000 465.300 676.200 ;
        RECT 448.950 667.950 451.050 670.050 ;
        RECT 462.000 666.600 463.800 675.000 ;
        RECT 482.400 672.600 483.600 679.950 ;
        RECT 500.400 672.600 501.600 679.950 ;
        RECT 518.400 672.600 519.600 679.950 ;
        RECT 524.550 673.050 525.450 679.950 ;
        RECT 527.550 676.050 528.450 697.950 ;
        RECT 535.800 695.400 537.600 701.400 ;
        RECT 536.700 695.100 537.600 695.400 ;
        RECT 541.800 695.400 543.600 701.400 ;
        RECT 550.950 697.950 553.050 700.050 ;
        RECT 541.800 695.100 543.300 695.400 ;
        RECT 536.700 694.200 543.300 695.100 ;
        RECT 536.700 682.050 537.600 694.200 ;
        RECT 538.950 682.950 541.050 685.050 ;
        RECT 535.950 679.950 538.050 682.050 ;
        RECT 539.100 681.150 540.900 682.950 ;
        RECT 542.100 682.050 543.900 683.850 ;
        RECT 544.950 682.950 547.050 685.050 ;
        RECT 541.950 679.950 544.050 682.050 ;
        RECT 545.100 681.150 546.900 682.950 ;
        RECT 536.700 676.200 537.600 679.950 ;
        RECT 527.100 673.950 529.200 676.050 ;
        RECT 536.700 675.000 540.000 676.200 ;
        RECT 481.800 666.600 483.600 672.600 ;
        RECT 499.800 666.600 501.600 672.600 ;
        RECT 517.800 666.600 519.600 672.600 ;
        RECT 523.800 670.950 525.900 673.050 ;
        RECT 538.200 666.600 540.000 675.000 ;
        RECT 551.550 673.050 552.450 697.950 ;
        RECT 560.400 695.400 562.200 701.400 ;
        RECT 560.700 695.100 562.200 695.400 ;
        RECT 566.400 695.400 568.200 701.400 ;
        RECT 574.950 697.950 577.050 700.050 ;
        RECT 566.400 695.100 567.300 695.400 ;
        RECT 560.700 694.200 567.300 695.100 ;
        RECT 556.950 682.950 559.050 685.050 ;
        RECT 557.100 681.150 558.900 682.950 ;
        RECT 560.100 682.050 561.900 683.850 ;
        RECT 562.950 682.950 565.050 685.050 ;
        RECT 559.950 679.950 562.050 682.050 ;
        RECT 563.100 681.150 564.900 682.950 ;
        RECT 566.400 682.050 567.300 694.200 ;
        RECT 565.950 679.950 568.050 682.050 ;
        RECT 566.400 676.200 567.300 679.950 ;
        RECT 575.550 679.050 576.450 697.950 ;
        RECT 581.400 690.300 583.200 701.400 ;
        RECT 587.400 690.300 589.200 701.400 ;
        RECT 581.400 689.400 589.200 690.300 ;
        RECT 590.400 689.400 592.200 701.400 ;
        RECT 608.400 689.400 610.200 701.400 ;
        RECT 626.400 695.400 628.200 701.400 ;
        RECT 637.950 697.950 640.050 700.050 ;
        RECT 580.950 682.950 583.050 685.050 ;
        RECT 581.100 681.150 582.900 682.950 ;
        RECT 584.100 682.050 585.900 683.850 ;
        RECT 586.950 682.950 589.050 685.050 ;
        RECT 583.950 679.950 586.050 682.050 ;
        RECT 587.100 681.150 588.900 682.950 ;
        RECT 590.400 682.050 591.600 689.400 ;
        RECT 604.950 682.950 607.050 685.050 ;
        RECT 589.950 679.950 592.050 682.050 ;
        RECT 605.100 681.150 606.900 682.950 ;
        RECT 608.400 682.050 609.600 689.400 ;
        RECT 613.950 688.950 616.050 691.050 ;
        RECT 607.950 679.950 610.050 682.050 ;
        RECT 574.950 676.950 577.050 679.050 ;
        RECT 564.000 675.000 567.300 676.200 ;
        RECT 550.950 670.950 553.050 673.050 ;
        RECT 564.000 666.600 565.800 675.000 ;
        RECT 590.400 672.600 591.600 679.950 ;
        RECT 586.500 671.400 591.600 672.600 ;
        RECT 608.400 672.600 609.600 679.950 ;
        RECT 614.550 673.050 615.450 688.950 ;
        RECT 622.950 682.950 625.050 685.050 ;
        RECT 623.100 681.150 624.900 682.950 ;
        RECT 626.400 682.050 627.600 695.400 ;
        RECT 628.950 682.950 631.050 685.050 ;
        RECT 625.950 679.950 628.050 682.050 ;
        RECT 629.100 681.150 630.900 682.950 ;
        RECT 626.400 674.700 627.600 679.950 ;
        RECT 626.400 673.800 630.600 674.700 ;
        RECT 586.500 666.600 588.300 671.400 ;
        RECT 608.400 666.600 610.200 672.600 ;
        RECT 613.950 670.950 616.050 673.050 ;
        RECT 628.800 666.600 630.600 673.800 ;
        RECT 638.550 670.050 639.450 697.950 ;
        RECT 649.800 695.400 651.600 701.400 ;
        RECT 655.800 697.950 657.900 700.050 ;
        RECT 661.950 697.950 664.050 700.050 ;
        RECT 644.100 682.050 645.900 683.850 ;
        RECT 646.950 682.950 649.050 685.050 ;
        RECT 643.950 679.950 646.050 682.050 ;
        RECT 647.100 681.150 648.900 682.950 ;
        RECT 649.950 682.050 651.150 695.400 ;
        RECT 656.550 687.450 657.450 697.950 ;
        RECT 656.550 686.550 660.450 687.450 ;
        RECT 652.950 682.950 655.050 685.050 ;
        RECT 649.950 679.950 652.050 682.050 ;
        RECT 653.100 681.150 654.900 682.950 ;
        RECT 650.850 675.750 652.050 679.950 ;
        RECT 659.550 676.050 660.450 686.550 ;
        RECT 650.850 674.700 654.600 675.750 ;
        RECT 644.400 671.700 652.200 673.050 ;
        RECT 637.950 667.950 640.050 670.050 ;
        RECT 644.400 666.600 646.200 671.700 ;
        RECT 650.400 666.600 652.200 671.700 ;
        RECT 653.400 672.600 654.600 674.700 ;
        RECT 655.950 674.550 660.450 676.050 ;
        RECT 655.950 673.950 660.000 674.550 ;
        RECT 662.550 673.050 663.450 697.950 ;
        RECT 671.400 695.400 673.200 701.400 ;
        RECT 667.950 682.950 670.050 685.050 ;
        RECT 668.100 681.150 669.900 682.950 ;
        RECT 671.400 682.050 672.600 695.400 ;
        RECT 692.700 690.600 694.500 701.400 ;
        RECT 715.800 695.400 717.600 701.400 ;
        RECT 721.950 699.450 726.000 700.050 ;
        RECT 721.950 697.950 726.450 699.450 ;
        RECT 692.700 689.400 696.300 690.600 ;
        RECT 673.950 682.950 676.050 685.050 ;
        RECT 670.950 679.950 673.050 682.050 ;
        RECT 674.100 681.150 675.900 682.950 ;
        RECT 695.400 682.050 696.300 689.400 ;
        RECT 710.100 682.050 711.900 683.850 ;
        RECT 712.950 682.950 715.050 685.050 ;
        RECT 671.400 674.700 672.600 679.950 ;
        RECT 692.100 679.050 693.900 680.850 ;
        RECT 694.950 679.950 697.050 682.050 ;
        RECT 691.950 676.950 694.050 679.050 ;
        RECT 671.400 673.800 675.600 674.700 ;
        RECT 653.400 666.600 655.200 672.600 ;
        RECT 661.950 670.950 664.050 673.050 ;
        RECT 673.800 666.600 675.600 673.800 ;
        RECT 695.400 669.600 696.300 679.950 ;
        RECT 698.100 679.050 699.900 680.850 ;
        RECT 709.950 679.950 712.050 682.050 ;
        RECT 713.100 681.150 714.900 682.950 ;
        RECT 715.950 682.050 717.150 695.400 ;
        RECT 718.950 682.950 721.050 685.050 ;
        RECT 715.950 679.950 718.050 682.050 ;
        RECT 719.100 681.150 720.900 682.950 ;
        RECT 697.950 676.950 700.050 679.050 ;
        RECT 716.850 675.750 718.050 679.950 ;
        RECT 716.850 674.700 720.600 675.750 ;
        RECT 710.400 671.700 718.200 673.050 ;
        RECT 694.800 666.600 696.600 669.600 ;
        RECT 710.400 666.600 712.200 671.700 ;
        RECT 716.400 666.600 718.200 671.700 ;
        RECT 719.400 672.600 720.600 674.700 ;
        RECT 719.400 666.600 721.200 672.600 ;
        RECT 725.550 670.050 726.450 697.950 ;
        RECT 730.950 694.950 733.050 697.050 ;
        RECT 739.800 695.400 741.600 701.400 ;
        RECT 751.950 697.950 754.050 700.050 ;
        RECT 731.550 685.050 732.450 694.950 ;
        RECT 727.950 683.550 732.450 685.050 ;
        RECT 727.950 682.950 732.000 683.550 ;
        RECT 736.950 682.950 739.050 685.050 ;
        RECT 737.100 681.150 738.900 682.950 ;
        RECT 740.400 682.050 741.600 695.400 ;
        RECT 742.950 682.950 745.050 685.050 ;
        RECT 739.950 679.950 742.050 682.050 ;
        RECT 743.100 681.150 744.900 682.950 ;
        RECT 752.550 682.050 753.450 697.950 ;
        RECT 761.400 695.400 763.200 701.400 ;
        RECT 772.950 697.950 775.050 700.050 ;
        RECT 757.950 682.950 760.050 685.050 ;
        RECT 751.950 679.950 754.050 682.050 ;
        RECT 758.100 681.150 759.900 682.950 ;
        RECT 761.850 682.050 763.050 695.400 ;
        RECT 763.950 682.950 766.050 685.050 ;
        RECT 760.950 679.950 763.050 682.050 ;
        RECT 764.100 681.150 765.900 682.950 ;
        RECT 767.100 682.050 768.900 683.850 ;
        RECT 766.950 679.950 769.050 682.050 ;
        RECT 733.950 676.950 736.050 679.050 ;
        RECT 734.550 670.050 735.450 676.950 ;
        RECT 740.400 674.700 741.600 679.950 ;
        RECT 760.950 675.750 762.150 679.950 ;
        RECT 737.400 673.800 741.600 674.700 ;
        RECT 758.400 674.700 762.150 675.750 ;
        RECT 724.950 667.950 727.050 670.050 ;
        RECT 733.950 667.950 736.050 670.050 ;
        RECT 737.400 666.600 739.200 673.800 ;
        RECT 758.400 672.600 759.600 674.700 ;
        RECT 757.800 666.600 759.600 672.600 ;
        RECT 760.800 671.700 768.600 673.050 ;
        RECT 760.800 666.600 762.600 671.700 ;
        RECT 766.800 666.600 768.600 671.700 ;
        RECT 773.550 670.050 774.450 697.950 ;
        RECT 782.400 695.400 784.200 701.400 ;
        RECT 782.700 695.100 784.200 695.400 ;
        RECT 788.400 695.400 790.200 701.400 ;
        RECT 806.400 695.400 808.200 701.400 ;
        RECT 788.400 695.100 789.300 695.400 ;
        RECT 782.700 694.200 789.300 695.100 ;
        RECT 778.950 682.950 781.050 685.050 ;
        RECT 779.100 681.150 780.900 682.950 ;
        RECT 782.100 682.050 783.900 683.850 ;
        RECT 784.950 682.950 787.050 685.050 ;
        RECT 781.950 679.950 784.050 682.050 ;
        RECT 785.100 681.150 786.900 682.950 ;
        RECT 788.400 682.050 789.300 694.200 ;
        RECT 802.950 682.950 805.050 685.050 ;
        RECT 787.950 679.950 790.050 682.050 ;
        RECT 803.100 681.150 804.900 682.950 ;
        RECT 806.400 682.050 807.600 695.400 ;
        RECT 824.400 690.300 826.200 701.400 ;
        RECT 830.400 690.300 832.200 701.400 ;
        RECT 824.400 689.400 832.200 690.300 ;
        RECT 833.400 689.400 835.200 701.400 ;
        RECT 841.950 697.950 844.050 700.050 ;
        RECT 808.950 682.950 811.050 685.050 ;
        RECT 823.950 682.950 826.050 685.050 ;
        RECT 805.950 679.950 808.050 682.050 ;
        RECT 809.100 681.150 810.900 682.950 ;
        RECT 824.100 681.150 825.900 682.950 ;
        RECT 827.100 682.050 828.900 683.850 ;
        RECT 829.950 682.950 832.050 685.050 ;
        RECT 826.950 679.950 829.050 682.050 ;
        RECT 830.100 681.150 831.900 682.950 ;
        RECT 833.400 682.050 834.600 689.400 ;
        RECT 832.950 679.950 835.050 682.050 ;
        RECT 788.400 676.200 789.300 679.950 ;
        RECT 770.100 668.550 774.450 670.050 ;
        RECT 786.000 675.000 789.300 676.200 ;
        RECT 770.100 667.950 774.000 668.550 ;
        RECT 786.000 666.600 787.800 675.000 ;
        RECT 806.400 674.700 807.600 679.950 ;
        RECT 806.400 673.800 810.600 674.700 ;
        RECT 808.800 666.600 810.600 673.800 ;
        RECT 833.400 672.600 834.600 679.950 ;
        RECT 842.550 679.050 843.450 697.950 ;
        RECT 854.400 695.400 856.200 701.400 ;
        RECT 850.950 682.950 853.050 685.050 ;
        RECT 851.100 681.150 852.900 682.950 ;
        RECT 854.850 682.050 856.050 695.400 ;
        RECT 865.950 694.950 868.050 697.050 ;
        RECT 877.800 695.400 879.600 701.400 ;
        RECT 856.950 682.950 859.050 685.050 ;
        RECT 853.950 679.950 856.050 682.050 ;
        RECT 857.100 681.150 858.900 682.950 ;
        RECT 860.100 682.050 861.900 683.850 ;
        RECT 859.950 679.950 862.050 682.050 ;
        RECT 841.950 676.950 844.050 679.050 ;
        RECT 853.950 675.750 855.150 679.950 ;
        RECT 851.400 674.700 855.150 675.750 ;
        RECT 851.400 672.600 852.600 674.700 ;
        RECT 866.550 673.050 867.450 694.950 ;
        RECT 872.100 682.050 873.900 683.850 ;
        RECT 874.950 682.950 877.050 685.050 ;
        RECT 871.950 679.950 874.050 682.050 ;
        RECT 875.100 681.150 876.900 682.950 ;
        RECT 877.950 682.050 879.150 695.400 ;
        RECT 886.950 694.950 889.050 697.050 ;
        RECT 899.400 695.400 901.200 701.400 ;
        RECT 904.950 697.950 907.050 700.050 ;
        RECT 880.950 682.950 883.050 685.050 ;
        RECT 877.950 679.950 880.050 682.050 ;
        RECT 881.100 681.150 882.900 682.950 ;
        RECT 878.850 675.750 880.050 679.950 ;
        RECT 878.850 674.700 882.600 675.750 ;
        RECT 829.500 671.400 834.600 672.600 ;
        RECT 829.500 666.600 831.300 671.400 ;
        RECT 850.800 666.600 852.600 672.600 ;
        RECT 853.800 671.700 861.600 673.050 ;
        RECT 853.800 666.600 855.600 671.700 ;
        RECT 859.800 666.600 861.600 671.700 ;
        RECT 865.950 670.950 868.050 673.050 ;
        RECT 872.400 671.700 880.200 673.050 ;
        RECT 872.400 666.600 874.200 671.700 ;
        RECT 878.400 666.600 880.200 671.700 ;
        RECT 881.400 672.600 882.600 674.700 ;
        RECT 887.550 673.050 888.450 694.950 ;
        RECT 899.400 688.050 900.600 695.400 ;
        RECT 890.100 685.950 892.200 688.050 ;
        RECT 890.550 682.050 891.450 685.950 ;
        RECT 896.100 682.050 897.900 683.850 ;
        RECT 898.950 682.950 901.050 688.050 ;
        RECT 889.950 679.950 892.050 682.050 ;
        RECT 895.950 679.950 898.050 682.050 ;
        RECT 881.400 666.600 883.200 672.600 ;
        RECT 886.950 670.950 889.050 673.050 ;
        RECT 899.400 669.600 900.600 682.950 ;
        RECT 905.550 670.050 906.450 697.950 ;
        RECT 899.400 666.600 901.200 669.600 ;
        RECT 905.550 668.550 910.050 670.050 ;
        RECT 906.000 667.950 910.050 668.550 ;
        RECT 16.200 654.000 18.000 662.400 ;
        RECT 40.500 657.600 42.300 662.400 ;
        RECT 61.800 659.400 63.600 662.400 ;
        RECT 82.800 659.400 84.600 662.400 ;
        RECT 40.500 656.400 45.600 657.600 ;
        RECT 14.700 652.800 18.000 654.000 ;
        RECT 14.700 649.050 15.600 652.800 ;
        RECT 44.400 649.050 45.600 656.400 ;
        RECT 49.950 655.950 52.050 658.050 ;
        RECT 13.950 646.950 16.050 649.050 ;
        RECT 14.700 634.800 15.600 646.950 ;
        RECT 17.100 646.050 18.900 647.850 ;
        RECT 19.950 646.950 22.050 649.050 ;
        RECT 16.950 643.950 19.050 646.050 ;
        RECT 20.100 645.150 21.900 646.950 ;
        RECT 23.100 646.050 24.900 647.850 ;
        RECT 35.100 646.050 36.900 647.850 ;
        RECT 37.950 646.950 40.050 649.050 ;
        RECT 22.950 643.950 25.050 646.050 ;
        RECT 28.950 643.950 31.050 646.050 ;
        RECT 34.950 643.950 37.050 646.050 ;
        RECT 38.100 645.150 39.900 646.950 ;
        RECT 41.100 646.050 42.900 647.850 ;
        RECT 43.950 646.950 46.050 649.050 ;
        RECT 40.950 643.950 43.050 646.050 ;
        RECT 14.700 633.900 21.300 634.800 ;
        RECT 14.700 633.600 15.600 633.900 ;
        RECT 13.800 627.600 15.600 633.600 ;
        RECT 19.800 633.600 21.300 633.900 ;
        RECT 19.800 627.600 21.600 633.600 ;
        RECT 29.550 631.050 30.450 643.950 ;
        RECT 44.400 639.600 45.600 646.950 ;
        RECT 35.400 638.700 43.200 639.600 ;
        RECT 28.800 628.950 30.900 631.050 ;
        RECT 35.400 627.600 37.200 638.700 ;
        RECT 41.400 627.600 43.200 638.700 ;
        RECT 44.400 627.600 46.200 639.600 ;
        RECT 50.550 637.050 51.450 655.950 ;
        RECT 62.400 646.050 63.600 659.400 ;
        RECT 79.950 649.950 82.050 652.050 ;
        RECT 64.950 646.950 67.050 649.050 ;
        RECT 80.100 648.150 81.900 649.950 ;
        RECT 83.400 649.050 84.300 659.400 ;
        RECT 104.700 657.600 106.500 662.400 ;
        RECT 101.400 656.400 106.500 657.600 ;
        RECT 85.950 649.950 88.050 652.050 ;
        RECT 82.950 646.950 85.050 649.050 ;
        RECT 86.100 648.150 87.900 649.950 ;
        RECT 101.400 649.050 102.600 656.400 ;
        RECT 129.000 654.000 130.800 662.400 ;
        RECT 138.150 656.400 139.950 662.400 ;
        RECT 145.950 660.300 147.750 662.400 ;
        RECT 144.000 659.400 147.750 660.300 ;
        RECT 153.750 659.400 155.550 662.400 ;
        RECT 161.550 659.400 163.350 662.400 ;
        RECT 144.000 658.500 145.050 659.400 ;
        RECT 153.750 658.500 154.800 659.400 ;
        RECT 142.950 656.400 145.050 658.500 ;
        RECT 129.000 652.800 132.300 654.000 ;
        RECT 131.400 649.050 132.300 652.800 ;
        RECT 100.950 646.950 103.050 649.050 ;
        RECT 61.950 640.950 64.050 646.050 ;
        RECT 65.100 645.150 66.900 646.950 ;
        RECT 49.950 634.950 52.050 637.050 ;
        RECT 62.400 633.600 63.600 640.950 ;
        RECT 83.400 639.600 84.300 646.950 ;
        RECT 101.400 639.600 102.600 646.950 ;
        RECT 104.100 646.050 105.900 647.850 ;
        RECT 106.950 646.950 109.050 649.050 ;
        RECT 103.950 643.950 106.050 646.050 ;
        RECT 107.100 645.150 108.900 646.950 ;
        RECT 110.100 646.050 111.900 647.850 ;
        RECT 122.100 646.050 123.900 647.850 ;
        RECT 124.950 646.950 127.050 649.050 ;
        RECT 109.950 643.950 112.050 646.050 ;
        RECT 121.950 643.950 124.050 646.050 ;
        RECT 125.100 645.150 126.900 646.950 ;
        RECT 128.100 646.050 129.900 647.850 ;
        RECT 130.950 646.950 133.050 649.050 ;
        RECT 127.950 643.950 130.050 646.050 ;
        RECT 61.800 627.600 63.600 633.600 ;
        RECT 80.700 638.400 84.300 639.600 ;
        RECT 80.700 627.600 82.500 638.400 ;
        RECT 100.800 627.600 102.600 639.600 ;
        RECT 103.800 638.700 111.600 639.600 ;
        RECT 103.800 627.600 105.600 638.700 ;
        RECT 109.800 627.600 111.600 638.700 ;
        RECT 131.400 634.800 132.300 646.950 ;
        RECT 125.700 633.900 132.300 634.800 ;
        RECT 125.700 633.600 127.200 633.900 ;
        RECT 125.400 627.600 127.200 633.600 ;
        RECT 131.400 633.600 132.300 633.900 ;
        RECT 138.150 641.700 139.050 656.400 ;
        RECT 146.550 655.800 148.350 657.600 ;
        RECT 149.850 657.450 154.800 658.500 ;
        RECT 162.300 658.500 163.350 659.400 ;
        RECT 149.850 656.700 151.650 657.450 ;
        RECT 162.300 657.300 166.050 658.500 ;
        RECT 163.950 656.400 166.050 657.300 ;
        RECT 169.650 656.400 171.450 662.400 ;
        RECT 185.400 659.400 187.200 662.400 ;
        RECT 146.850 654.000 147.900 655.800 ;
        RECT 157.050 654.000 158.850 654.600 ;
        RECT 146.850 652.800 158.850 654.000 ;
        RECT 141.000 651.600 147.900 652.800 ;
        RECT 141.000 650.850 141.900 651.600 ;
        RECT 146.100 651.000 147.900 651.600 ;
        RECT 140.100 649.050 141.900 650.850 ;
        RECT 143.100 649.800 144.900 650.400 ;
        RECT 139.950 646.950 142.050 649.050 ;
        RECT 143.100 648.600 151.050 649.800 ;
        RECT 148.950 646.950 151.050 648.600 ;
        RECT 147.450 641.700 149.250 642.000 ;
        RECT 138.150 641.100 149.250 641.700 ;
        RECT 138.150 640.500 155.850 641.100 ;
        RECT 138.150 639.600 139.050 640.500 ;
        RECT 147.450 640.200 155.850 640.500 ;
        RECT 131.400 627.600 133.200 633.600 ;
        RECT 138.150 627.600 139.950 639.600 ;
        RECT 152.250 638.700 154.050 639.300 ;
        RECT 146.550 637.500 154.050 638.700 ;
        RECT 154.950 638.100 155.850 640.200 ;
        RECT 157.950 640.200 158.850 652.800 ;
        RECT 170.250 649.050 171.450 656.400 ;
        RECT 181.950 649.950 184.050 652.050 ;
        RECT 165.150 647.250 171.450 649.050 ;
        RECT 182.100 648.150 183.900 649.950 ;
        RECT 185.700 649.050 186.600 659.400 ;
        RECT 208.800 655.200 210.600 662.400 ;
        RECT 226.800 659.400 228.600 662.400 ;
        RECT 206.400 654.300 210.600 655.200 ;
        RECT 187.950 649.950 190.050 652.050 ;
        RECT 166.950 646.950 171.450 647.250 ;
        RECT 184.950 646.950 187.050 649.050 ;
        RECT 188.100 648.150 189.900 649.950 ;
        RECT 206.400 649.050 207.600 654.300 ;
        RECT 167.250 641.400 169.050 643.200 ;
        RECT 163.950 640.200 168.150 641.400 ;
        RECT 157.950 639.300 163.050 640.200 ;
        RECT 163.950 639.300 166.050 640.200 ;
        RECT 170.250 639.600 171.450 646.950 ;
        RECT 178.950 640.950 181.050 643.050 ;
        RECT 162.150 638.400 163.050 639.300 ;
        RECT 159.450 638.100 161.250 638.400 ;
        RECT 146.550 636.600 147.750 637.500 ;
        RECT 154.950 637.200 161.250 638.100 ;
        RECT 159.450 636.600 161.250 637.200 ;
        RECT 162.150 636.600 164.850 638.400 ;
        RECT 142.950 634.500 147.750 636.600 ;
        RECT 150.450 635.550 152.250 636.300 ;
        RECT 155.250 635.550 157.050 636.300 ;
        RECT 150.450 634.500 157.050 635.550 ;
        RECT 146.550 633.600 147.750 634.500 ;
        RECT 146.550 627.600 148.350 633.600 ;
        RECT 154.350 627.600 156.150 634.500 ;
        RECT 162.150 633.600 166.050 635.700 ;
        RECT 162.150 627.600 163.950 633.600 ;
        RECT 169.650 627.600 171.450 639.600 ;
        RECT 179.550 637.050 180.450 640.950 ;
        RECT 185.700 639.600 186.600 646.950 ;
        RECT 203.100 646.050 204.900 647.850 ;
        RECT 205.950 646.950 208.050 649.050 ;
        RECT 202.950 643.950 205.050 646.050 ;
        RECT 185.700 638.400 189.300 639.600 ;
        RECT 178.950 634.950 181.050 637.050 ;
        RECT 187.500 627.600 189.300 638.400 ;
        RECT 206.400 633.600 207.600 646.950 ;
        RECT 209.100 646.050 210.900 647.850 ;
        RECT 227.400 646.050 228.600 659.400 ;
        RECT 235.950 658.950 238.050 661.050 ;
        RECT 229.950 646.950 232.050 649.050 ;
        RECT 208.950 643.950 211.050 646.050 ;
        RECT 226.950 640.950 229.050 646.050 ;
        RECT 230.100 645.150 231.900 646.950 ;
        RECT 236.550 646.050 237.450 658.950 ;
        RECT 244.800 656.400 246.600 662.400 ;
        RECT 245.400 654.300 246.600 656.400 ;
        RECT 247.800 657.300 249.600 662.400 ;
        RECT 253.800 657.300 255.600 662.400 ;
        RECT 247.800 655.950 255.600 657.300 ;
        RECT 266.400 654.600 268.200 662.400 ;
        RECT 273.900 658.200 275.700 662.400 ;
        RECT 273.900 656.400 276.600 658.200 ;
        RECT 272.100 654.600 273.900 655.500 ;
        RECT 245.400 653.250 249.150 654.300 ;
        RECT 266.400 653.700 273.900 654.600 ;
        RECT 247.950 649.050 249.150 653.250 ;
        RECT 266.100 649.050 267.900 650.850 ;
        RECT 245.100 646.050 246.900 647.850 ;
        RECT 247.950 646.950 250.050 649.050 ;
        RECT 235.950 643.950 238.050 646.050 ;
        RECT 244.950 643.950 247.050 646.050 ;
        RECT 227.400 633.600 228.600 640.950 ;
        RECT 248.850 633.600 250.050 646.950 ;
        RECT 251.100 646.050 252.900 647.850 ;
        RECT 253.950 646.950 256.050 649.050 ;
        RECT 265.950 646.950 268.050 649.050 ;
        RECT 250.950 643.950 253.050 646.050 ;
        RECT 254.100 645.150 255.900 646.950 ;
        RECT 269.400 633.600 270.300 653.700 ;
        RECT 275.700 649.050 276.600 656.400 ;
        RECT 280.950 655.950 283.050 658.050 ;
        RECT 271.950 646.950 274.050 649.050 ;
        RECT 274.950 646.950 277.050 649.050 ;
        RECT 272.100 645.150 273.900 646.950 ;
        RECT 275.700 639.600 276.600 646.950 ;
        RECT 281.550 646.050 282.450 655.950 ;
        RECT 293.400 655.200 295.200 662.400 ;
        RECT 313.800 656.400 315.600 662.400 ;
        RECT 293.400 654.300 297.600 655.200 ;
        RECT 296.400 649.050 297.600 654.300 ;
        RECT 314.400 654.300 315.600 656.400 ;
        RECT 316.800 657.300 318.600 662.400 ;
        RECT 322.800 657.300 324.600 662.400 ;
        RECT 316.800 655.950 324.600 657.300 ;
        RECT 335.400 657.300 337.200 662.400 ;
        RECT 341.400 657.300 343.200 662.400 ;
        RECT 335.400 655.950 343.200 657.300 ;
        RECT 344.400 656.400 346.200 662.400 ;
        RECT 361.800 656.400 363.600 662.400 ;
        RECT 344.400 654.300 345.600 656.400 ;
        RECT 314.400 653.250 318.150 654.300 ;
        RECT 316.950 649.050 318.150 653.250 ;
        RECT 341.850 653.250 345.600 654.300 ;
        RECT 362.400 654.300 363.600 656.400 ;
        RECT 364.800 657.300 366.600 662.400 ;
        RECT 370.800 657.300 372.600 662.400 ;
        RECT 364.800 655.950 372.600 657.300 ;
        RECT 375.150 656.400 376.950 662.400 ;
        RECT 382.950 660.300 384.750 662.400 ;
        RECT 381.000 659.400 384.750 660.300 ;
        RECT 390.750 659.400 392.550 662.400 ;
        RECT 398.550 659.400 400.350 662.400 ;
        RECT 381.000 658.500 382.050 659.400 ;
        RECT 390.750 658.500 391.800 659.400 ;
        RECT 379.950 656.400 382.050 658.500 ;
        RECT 362.400 653.250 366.150 654.300 ;
        RECT 341.850 649.050 343.050 653.250 ;
        RECT 293.100 646.050 294.900 647.850 ;
        RECT 295.950 646.950 298.050 649.050 ;
        RECT 280.950 643.950 283.050 646.050 ;
        RECT 292.950 643.950 295.050 646.050 ;
        RECT 206.400 627.600 208.200 633.600 ;
        RECT 226.800 627.600 228.600 633.600 ;
        RECT 248.400 627.600 250.200 633.600 ;
        RECT 269.400 627.600 271.200 633.600 ;
        RECT 275.700 627.600 277.500 639.600 ;
        RECT 296.400 633.600 297.600 646.950 ;
        RECT 299.100 646.050 300.900 647.850 ;
        RECT 314.100 646.050 315.900 647.850 ;
        RECT 316.950 646.950 319.050 649.050 ;
        RECT 298.950 643.950 301.050 646.050 ;
        RECT 313.950 643.950 316.050 646.050 ;
        RECT 317.850 633.600 319.050 646.950 ;
        RECT 320.100 646.050 321.900 647.850 ;
        RECT 322.950 646.950 325.050 649.050 ;
        RECT 334.950 646.950 337.050 649.050 ;
        RECT 319.950 643.950 322.050 646.050 ;
        RECT 323.100 645.150 324.900 646.950 ;
        RECT 327.000 645.450 331.050 646.050 ;
        RECT 326.550 643.950 331.050 645.450 ;
        RECT 335.100 645.150 336.900 646.950 ;
        RECT 338.100 646.050 339.900 647.850 ;
        RECT 340.950 646.950 343.050 649.050 ;
        RECT 364.950 649.050 366.150 653.250 ;
        RECT 337.950 643.950 340.050 646.050 ;
        RECT 295.800 627.600 297.600 633.600 ;
        RECT 317.400 627.600 319.200 633.600 ;
        RECT 326.550 631.050 327.450 643.950 ;
        RECT 340.950 633.600 342.150 646.950 ;
        RECT 344.100 646.050 345.900 647.850 ;
        RECT 362.100 646.050 363.900 647.850 ;
        RECT 364.950 646.950 367.050 649.050 ;
        RECT 343.950 643.950 346.050 646.050 ;
        RECT 361.950 643.950 364.050 646.050 ;
        RECT 365.850 633.600 367.050 646.950 ;
        RECT 368.100 646.050 369.900 647.850 ;
        RECT 370.950 646.950 373.050 649.050 ;
        RECT 367.950 643.950 370.050 646.050 ;
        RECT 371.100 645.150 372.900 646.950 ;
        RECT 375.150 641.700 376.050 656.400 ;
        RECT 383.550 655.800 385.350 657.600 ;
        RECT 386.850 657.450 391.800 658.500 ;
        RECT 399.300 658.500 400.350 659.400 ;
        RECT 386.850 656.700 388.650 657.450 ;
        RECT 399.300 657.300 403.050 658.500 ;
        RECT 400.950 656.400 403.050 657.300 ;
        RECT 406.650 656.400 408.450 662.400 ;
        RECT 383.850 654.000 384.900 655.800 ;
        RECT 394.050 654.000 395.850 654.600 ;
        RECT 383.850 652.800 395.850 654.000 ;
        RECT 378.000 651.600 384.900 652.800 ;
        RECT 378.000 650.850 378.900 651.600 ;
        RECT 383.100 651.000 384.900 651.600 ;
        RECT 377.100 649.050 378.900 650.850 ;
        RECT 380.100 649.800 381.900 650.400 ;
        RECT 376.950 646.950 379.050 649.050 ;
        RECT 380.100 648.600 388.050 649.800 ;
        RECT 385.950 646.950 388.050 648.600 ;
        RECT 384.450 641.700 386.250 642.000 ;
        RECT 375.150 641.100 386.250 641.700 ;
        RECT 375.150 640.500 392.850 641.100 ;
        RECT 375.150 639.600 376.050 640.500 ;
        RECT 384.450 640.200 392.850 640.500 ;
        RECT 325.950 628.950 328.050 631.050 ;
        RECT 340.800 627.600 342.600 633.600 ;
        RECT 365.400 627.600 367.200 633.600 ;
        RECT 375.150 627.600 376.950 639.600 ;
        RECT 389.250 638.700 391.050 639.300 ;
        RECT 383.550 637.500 391.050 638.700 ;
        RECT 391.950 638.100 392.850 640.200 ;
        RECT 394.950 640.200 395.850 652.800 ;
        RECT 407.250 649.050 408.450 656.400 ;
        RECT 426.000 654.000 427.800 662.400 ;
        RECT 442.950 658.950 445.050 661.050 ;
        RECT 426.000 652.800 429.300 654.000 ;
        RECT 428.400 649.050 429.300 652.800 ;
        RECT 443.550 652.050 444.450 658.950 ;
        RECT 447.300 658.200 449.100 662.400 ;
        RECT 446.400 656.400 449.100 658.200 ;
        RECT 442.950 649.950 445.050 652.050 ;
        RECT 446.400 649.050 447.300 656.400 ;
        RECT 449.100 654.600 450.900 655.500 ;
        RECT 454.800 654.600 456.600 662.400 ;
        RECT 472.800 655.200 474.600 662.400 ;
        RECT 490.800 659.400 492.600 662.400 ;
        RECT 482.100 655.950 484.200 658.050 ;
        RECT 449.100 653.700 456.600 654.600 ;
        RECT 470.400 654.300 474.600 655.200 ;
        RECT 402.150 647.250 408.450 649.050 ;
        RECT 403.950 646.950 408.450 647.250 ;
        RECT 404.250 641.400 406.050 643.200 ;
        RECT 400.950 640.200 405.150 641.400 ;
        RECT 394.950 639.300 400.050 640.200 ;
        RECT 400.950 639.300 403.050 640.200 ;
        RECT 407.250 639.600 408.450 646.950 ;
        RECT 419.100 646.050 420.900 647.850 ;
        RECT 421.950 646.950 424.050 649.050 ;
        RECT 418.950 643.950 421.050 646.050 ;
        RECT 422.100 645.150 423.900 646.950 ;
        RECT 425.100 646.050 426.900 647.850 ;
        RECT 427.950 646.950 430.050 649.050 ;
        RECT 445.950 646.950 448.050 649.050 ;
        RECT 448.950 646.950 451.050 649.050 ;
        RECT 424.950 643.950 427.050 646.050 ;
        RECT 399.150 638.400 400.050 639.300 ;
        RECT 396.450 638.100 398.250 638.400 ;
        RECT 383.550 636.600 384.750 637.500 ;
        RECT 391.950 637.200 398.250 638.100 ;
        RECT 396.450 636.600 398.250 637.200 ;
        RECT 399.150 636.600 401.850 638.400 ;
        RECT 379.950 634.500 384.750 636.600 ;
        RECT 387.450 635.550 389.250 636.300 ;
        RECT 392.250 635.550 394.050 636.300 ;
        RECT 387.450 634.500 394.050 635.550 ;
        RECT 383.550 633.600 384.750 634.500 ;
        RECT 383.550 627.600 385.350 633.600 ;
        RECT 391.350 627.600 393.150 634.500 ;
        RECT 399.150 633.600 403.050 635.700 ;
        RECT 399.150 627.600 400.950 633.600 ;
        RECT 406.650 627.600 408.450 639.600 ;
        RECT 415.950 634.950 418.050 637.050 ;
        RECT 416.550 631.050 417.450 634.950 ;
        RECT 428.400 634.800 429.300 646.950 ;
        RECT 446.400 639.600 447.300 646.950 ;
        RECT 449.100 645.150 450.900 646.950 ;
        RECT 422.700 633.900 429.300 634.800 ;
        RECT 422.700 633.600 424.200 633.900 ;
        RECT 413.100 629.550 417.450 631.050 ;
        RECT 413.100 628.950 417.000 629.550 ;
        RECT 422.400 627.600 424.200 633.600 ;
        RECT 428.400 633.600 429.300 633.900 ;
        RECT 428.400 627.600 430.200 633.600 ;
        RECT 445.500 627.600 447.300 639.600 ;
        RECT 452.700 633.600 453.600 653.700 ;
        RECT 455.100 649.050 456.900 650.850 ;
        RECT 470.400 649.050 471.600 654.300 ;
        RECT 454.950 646.950 457.050 649.050 ;
        RECT 467.100 646.050 468.900 647.850 ;
        RECT 469.950 646.950 472.050 649.050 ;
        RECT 466.950 643.950 469.050 646.050 ;
        RECT 451.800 627.600 453.600 633.600 ;
        RECT 470.400 633.600 471.600 646.950 ;
        RECT 473.100 646.050 474.900 647.850 ;
        RECT 472.950 643.950 475.050 646.050 ;
        RECT 482.550 637.050 483.450 655.950 ;
        RECT 491.400 646.050 492.600 659.400 ;
        RECT 508.800 656.400 510.600 662.400 ;
        RECT 509.400 654.300 510.600 656.400 ;
        RECT 511.800 657.300 513.600 662.400 ;
        RECT 517.800 657.300 519.600 662.400 ;
        RECT 511.800 655.950 519.600 657.300 ;
        RECT 522.150 656.400 523.950 662.400 ;
        RECT 529.950 660.300 531.750 662.400 ;
        RECT 528.000 659.400 531.750 660.300 ;
        RECT 537.750 659.400 539.550 662.400 ;
        RECT 545.550 659.400 547.350 662.400 ;
        RECT 528.000 658.500 529.050 659.400 ;
        RECT 537.750 658.500 538.800 659.400 ;
        RECT 526.950 656.400 529.050 658.500 ;
        RECT 509.400 653.250 513.150 654.300 ;
        RECT 511.950 649.050 513.150 653.250 ;
        RECT 493.950 646.950 496.050 649.050 ;
        RECT 490.950 640.950 493.050 646.050 ;
        RECT 494.100 645.150 495.900 646.950 ;
        RECT 509.100 646.050 510.900 647.850 ;
        RECT 511.950 646.950 514.050 649.050 ;
        RECT 508.950 643.950 511.050 646.050 ;
        RECT 481.950 634.950 484.050 637.050 ;
        RECT 491.400 633.600 492.600 640.950 ;
        RECT 512.850 633.600 514.050 646.950 ;
        RECT 515.100 646.050 516.900 647.850 ;
        RECT 517.950 646.950 520.050 649.050 ;
        RECT 514.950 643.950 517.050 646.050 ;
        RECT 518.100 645.150 519.900 646.950 ;
        RECT 522.150 641.700 523.050 656.400 ;
        RECT 530.550 655.800 532.350 657.600 ;
        RECT 533.850 657.450 538.800 658.500 ;
        RECT 546.300 658.500 547.350 659.400 ;
        RECT 533.850 656.700 535.650 657.450 ;
        RECT 546.300 657.300 550.050 658.500 ;
        RECT 547.950 656.400 550.050 657.300 ;
        RECT 553.650 656.400 555.450 662.400 ;
        RECT 530.850 654.000 531.900 655.800 ;
        RECT 541.050 654.000 542.850 654.600 ;
        RECT 530.850 652.800 542.850 654.000 ;
        RECT 525.000 651.600 531.900 652.800 ;
        RECT 525.000 650.850 525.900 651.600 ;
        RECT 530.100 651.000 531.900 651.600 ;
        RECT 524.100 649.050 525.900 650.850 ;
        RECT 527.100 649.800 528.900 650.400 ;
        RECT 523.950 646.950 526.050 649.050 ;
        RECT 527.100 648.600 535.050 649.800 ;
        RECT 532.950 646.950 535.050 648.600 ;
        RECT 531.450 641.700 533.250 642.000 ;
        RECT 522.150 641.100 533.250 641.700 ;
        RECT 522.150 640.500 539.850 641.100 ;
        RECT 522.150 639.600 523.050 640.500 ;
        RECT 531.450 640.200 539.850 640.500 ;
        RECT 470.400 627.600 472.200 633.600 ;
        RECT 490.800 627.600 492.600 633.600 ;
        RECT 512.400 627.600 514.200 633.600 ;
        RECT 522.150 627.600 523.950 639.600 ;
        RECT 536.250 638.700 538.050 639.300 ;
        RECT 530.550 637.500 538.050 638.700 ;
        RECT 538.950 638.100 539.850 640.200 ;
        RECT 541.950 640.200 542.850 652.800 ;
        RECT 554.250 649.050 555.450 656.400 ;
        RECT 566.400 654.600 568.200 662.400 ;
        RECT 573.900 658.200 575.700 662.400 ;
        RECT 581.100 658.950 583.200 661.050 ;
        RECT 573.900 656.400 576.600 658.200 ;
        RECT 572.100 654.600 573.900 655.500 ;
        RECT 566.400 653.700 573.900 654.600 ;
        RECT 566.100 649.050 567.900 650.850 ;
        RECT 549.150 647.250 555.450 649.050 ;
        RECT 550.950 646.950 555.450 647.250 ;
        RECT 565.950 646.950 568.050 649.050 ;
        RECT 551.250 641.400 553.050 643.200 ;
        RECT 547.950 640.200 552.150 641.400 ;
        RECT 541.950 639.300 547.050 640.200 ;
        RECT 547.950 639.300 550.050 640.200 ;
        RECT 554.250 639.600 555.450 646.950 ;
        RECT 546.150 638.400 547.050 639.300 ;
        RECT 543.450 638.100 545.250 638.400 ;
        RECT 530.550 636.600 531.750 637.500 ;
        RECT 538.950 637.200 545.250 638.100 ;
        RECT 543.450 636.600 545.250 637.200 ;
        RECT 546.150 636.600 548.850 638.400 ;
        RECT 526.950 634.500 531.750 636.600 ;
        RECT 534.450 635.550 536.250 636.300 ;
        RECT 539.250 635.550 541.050 636.300 ;
        RECT 534.450 634.500 541.050 635.550 ;
        RECT 530.550 633.600 531.750 634.500 ;
        RECT 530.550 627.600 532.350 633.600 ;
        RECT 538.350 627.600 540.150 634.500 ;
        RECT 546.150 633.600 550.050 635.700 ;
        RECT 546.150 627.600 547.950 633.600 ;
        RECT 553.650 627.600 555.450 639.600 ;
        RECT 569.400 633.600 570.300 653.700 ;
        RECT 575.700 649.050 576.600 656.400 ;
        RECT 571.950 646.950 574.050 649.050 ;
        RECT 574.950 646.950 577.050 649.050 ;
        RECT 572.100 645.150 573.900 646.950 ;
        RECT 575.700 639.600 576.600 646.950 ;
        RECT 569.400 627.600 571.200 633.600 ;
        RECT 575.700 627.600 577.500 639.600 ;
        RECT 581.550 637.050 582.450 658.950 ;
        RECT 592.800 656.400 594.600 662.400 ;
        RECT 593.400 654.300 594.600 656.400 ;
        RECT 595.800 657.300 597.600 662.400 ;
        RECT 601.800 657.300 603.600 662.400 ;
        RECT 595.800 655.950 603.600 657.300 ;
        RECT 593.400 653.250 597.150 654.300 ;
        RECT 619.200 654.000 621.000 662.400 ;
        RECT 586.950 649.950 589.050 652.050 ;
        RECT 587.550 637.050 588.450 649.950 ;
        RECT 595.950 649.050 597.150 653.250 ;
        RECT 617.700 652.800 621.000 654.000 ;
        RECT 641.400 659.400 643.200 662.400 ;
        RECT 617.700 649.050 618.600 652.800 ;
        RECT 593.100 646.050 594.900 647.850 ;
        RECT 595.950 646.950 598.050 649.050 ;
        RECT 592.950 643.950 595.050 646.050 ;
        RECT 580.950 634.950 583.050 637.050 ;
        RECT 586.950 634.950 589.050 637.050 ;
        RECT 596.850 633.600 598.050 646.950 ;
        RECT 599.100 646.050 600.900 647.850 ;
        RECT 601.950 646.950 604.050 649.050 ;
        RECT 616.950 646.950 619.050 649.050 ;
        RECT 598.950 643.950 601.050 646.050 ;
        RECT 602.100 645.150 603.900 646.950 ;
        RECT 617.700 634.800 618.600 646.950 ;
        RECT 620.100 646.050 621.900 647.850 ;
        RECT 622.950 646.950 625.050 649.050 ;
        RECT 619.950 643.950 622.050 646.050 ;
        RECT 623.100 645.150 624.900 646.950 ;
        RECT 626.100 646.050 627.900 647.850 ;
        RECT 637.950 646.950 640.050 649.050 ;
        RECT 625.950 643.950 628.050 646.050 ;
        RECT 638.100 645.150 639.900 646.950 ;
        RECT 641.400 646.050 642.600 659.400 ;
        RECT 656.400 657.300 658.200 662.400 ;
        RECT 662.400 657.300 664.200 662.400 ;
        RECT 656.400 655.950 664.200 657.300 ;
        RECT 665.400 656.400 667.200 662.400 ;
        RECT 665.400 654.300 666.600 656.400 ;
        RECT 662.850 653.250 666.600 654.300 ;
        RECT 680.400 654.600 682.200 662.400 ;
        RECT 687.900 658.200 689.700 662.400 ;
        RECT 707.400 659.400 709.200 662.400 ;
        RECT 687.900 656.400 690.600 658.200 ;
        RECT 686.100 654.600 687.900 655.500 ;
        RECT 680.400 653.700 687.900 654.600 ;
        RECT 662.850 649.050 664.050 653.250 ;
        RECT 680.100 649.050 681.900 650.850 ;
        RECT 655.950 646.950 658.050 649.050 ;
        RECT 640.950 640.950 643.050 646.050 ;
        RECT 656.100 645.150 657.900 646.950 ;
        RECT 659.100 646.050 660.900 647.850 ;
        RECT 661.950 646.950 664.050 649.050 ;
        RECT 658.950 643.950 661.050 646.050 ;
        RECT 617.700 633.900 624.300 634.800 ;
        RECT 617.700 633.600 618.600 633.900 ;
        RECT 596.400 627.600 598.200 633.600 ;
        RECT 616.800 627.600 618.600 633.600 ;
        RECT 622.800 633.600 624.300 633.900 ;
        RECT 641.400 633.600 642.600 640.950 ;
        RECT 661.950 633.600 663.150 646.950 ;
        RECT 665.100 646.050 666.900 647.850 ;
        RECT 679.950 646.950 682.050 649.050 ;
        RECT 664.950 643.950 667.050 646.050 ;
        RECT 683.400 633.600 684.300 653.700 ;
        RECT 689.700 649.050 690.600 656.400 ;
        RECT 703.950 649.950 706.050 652.050 ;
        RECT 685.950 646.950 688.050 649.050 ;
        RECT 688.950 646.950 691.050 649.050 ;
        RECT 704.100 648.150 705.900 649.950 ;
        RECT 707.700 649.050 708.600 659.400 ;
        RECT 725.400 657.300 727.200 662.400 ;
        RECT 731.400 657.300 733.200 662.400 ;
        RECT 725.400 655.950 733.200 657.300 ;
        RECT 734.400 656.400 736.200 662.400 ;
        RECT 739.950 658.950 742.050 661.050 ;
        RECT 718.950 652.950 721.050 655.050 ;
        RECT 734.400 654.300 735.600 656.400 ;
        RECT 731.850 653.250 735.600 654.300 ;
        RECT 709.950 649.950 712.050 652.050 ;
        RECT 706.950 646.950 709.050 649.050 ;
        RECT 710.100 648.150 711.900 649.950 ;
        RECT 686.100 645.150 687.900 646.950 ;
        RECT 689.700 639.600 690.600 646.950 ;
        RECT 707.700 639.600 708.600 646.950 ;
        RECT 622.800 627.600 624.600 633.600 ;
        RECT 641.400 627.600 643.200 633.600 ;
        RECT 661.800 627.600 663.600 633.600 ;
        RECT 683.400 627.600 685.200 633.600 ;
        RECT 689.700 627.600 691.500 639.600 ;
        RECT 707.700 638.400 711.300 639.600 ;
        RECT 709.500 627.600 711.300 638.400 ;
        RECT 719.550 631.050 720.450 652.950 ;
        RECT 731.850 649.050 733.050 653.250 ;
        RECT 724.950 646.950 727.050 649.050 ;
        RECT 725.100 645.150 726.900 646.950 ;
        RECT 728.100 646.050 729.900 647.850 ;
        RECT 730.950 646.950 733.050 649.050 ;
        RECT 727.950 643.950 730.050 646.050 ;
        RECT 730.950 633.600 732.150 646.950 ;
        RECT 734.100 646.050 735.900 647.850 ;
        RECT 733.950 643.950 736.050 646.050 ;
        RECT 740.550 640.050 741.450 658.950 ;
        RECT 749.400 657.300 751.200 662.400 ;
        RECT 755.400 657.300 757.200 662.400 ;
        RECT 749.400 655.950 757.200 657.300 ;
        RECT 758.400 656.400 760.200 662.400 ;
        RECT 775.800 656.400 777.600 662.400 ;
        RECT 758.400 654.300 759.600 656.400 ;
        RECT 755.850 653.250 759.600 654.300 ;
        RECT 776.400 654.300 777.600 656.400 ;
        RECT 778.800 657.300 780.600 662.400 ;
        RECT 784.800 657.300 786.600 662.400 ;
        RECT 778.800 655.950 786.600 657.300 ;
        RECT 802.800 655.200 804.600 662.400 ;
        RECT 800.400 654.300 804.600 655.200 ;
        RECT 821.400 655.200 823.200 662.400 ;
        RECT 842.400 659.400 844.200 662.400 ;
        RECT 843.300 655.200 844.200 659.400 ;
        RECT 848.400 656.400 850.200 662.400 ;
        RECT 856.950 658.950 859.050 661.050 ;
        RECT 821.400 654.300 825.600 655.200 ;
        RECT 843.300 654.300 846.600 655.200 ;
        RECT 776.400 653.250 780.150 654.300 ;
        RECT 755.850 649.050 757.050 653.250 ;
        RECT 748.950 646.950 751.050 649.050 ;
        RECT 742.950 645.450 747.000 646.050 ;
        RECT 742.950 643.950 747.450 645.450 ;
        RECT 749.100 645.150 750.900 646.950 ;
        RECT 752.100 646.050 753.900 647.850 ;
        RECT 754.950 646.950 757.050 649.050 ;
        RECT 778.950 649.050 780.150 653.250 ;
        RECT 790.950 649.950 793.050 652.050 ;
        RECT 751.950 643.950 754.050 646.050 ;
        RECT 739.950 637.950 742.050 640.050 ;
        RECT 746.550 637.050 747.450 643.950 ;
        RECT 745.950 634.950 748.050 637.050 ;
        RECT 754.950 633.600 756.150 646.950 ;
        RECT 758.100 646.050 759.900 647.850 ;
        RECT 776.100 646.050 777.900 647.850 ;
        RECT 778.950 646.950 781.050 649.050 ;
        RECT 757.950 643.950 760.050 646.050 ;
        RECT 775.950 643.950 778.050 646.050 ;
        RECT 779.850 633.600 781.050 646.950 ;
        RECT 782.100 646.050 783.900 647.850 ;
        RECT 784.950 646.950 787.050 649.050 ;
        RECT 781.950 643.950 784.050 646.050 ;
        RECT 785.100 645.150 786.900 646.950 ;
        RECT 791.550 640.050 792.450 649.950 ;
        RECT 800.400 649.050 801.600 654.300 ;
        RECT 824.400 649.050 825.600 654.300 ;
        RECT 844.800 653.400 846.600 654.300 ;
        RECT 797.100 646.050 798.900 647.850 ;
        RECT 799.950 646.950 802.050 649.050 ;
        RECT 796.950 643.950 799.050 646.050 ;
        RECT 790.950 637.950 793.050 640.050 ;
        RECT 800.400 633.600 801.600 646.950 ;
        RECT 803.100 646.050 804.900 647.850 ;
        RECT 821.100 646.050 822.900 647.850 ;
        RECT 823.950 646.950 826.050 649.050 ;
        RECT 802.950 643.950 805.050 646.050 ;
        RECT 820.950 643.950 823.050 646.050 ;
        RECT 824.400 633.600 825.600 646.950 ;
        RECT 827.100 646.050 828.900 647.850 ;
        RECT 839.100 646.050 840.900 647.850 ;
        RECT 841.950 646.950 844.050 649.050 ;
        RECT 826.950 643.950 829.050 646.050 ;
        RECT 838.950 643.950 841.050 646.050 ;
        RECT 842.100 645.150 843.900 646.950 ;
        RECT 845.700 642.900 846.600 653.400 ;
        RECT 849.000 649.050 850.050 656.400 ;
        RECT 844.800 642.300 846.600 642.900 ;
        RECT 718.950 628.950 721.050 631.050 ;
        RECT 730.800 627.600 732.600 633.600 ;
        RECT 754.800 627.600 756.600 633.600 ;
        RECT 779.400 627.600 781.200 633.600 ;
        RECT 800.400 627.600 802.200 633.600 ;
        RECT 823.800 627.600 825.600 633.600 ;
        RECT 839.400 641.100 846.600 642.300 ;
        RECT 847.950 646.950 850.050 649.050 ;
        RECT 839.400 639.600 840.600 641.100 ;
        RECT 847.950 639.600 849.300 646.950 ;
        RECT 839.400 627.600 841.200 639.600 ;
        RECT 846.900 638.100 849.300 639.600 ;
        RECT 846.900 627.600 848.700 638.100 ;
        RECT 857.550 631.050 858.450 658.950 ;
        RECT 868.200 654.000 870.000 662.400 ;
        RECT 866.700 652.800 870.000 654.000 ;
        RECT 894.000 654.000 895.800 662.400 ;
        RECT 894.000 652.800 897.300 654.000 ;
        RECT 859.950 649.950 862.050 652.050 ;
        RECT 860.550 637.050 861.450 649.950 ;
        RECT 866.700 649.050 867.600 652.800 ;
        RECT 896.400 649.050 897.300 652.800 ;
        RECT 865.950 646.950 868.050 649.050 ;
        RECT 859.950 634.950 862.050 637.050 ;
        RECT 866.700 634.800 867.600 646.950 ;
        RECT 869.100 646.050 870.900 647.850 ;
        RECT 871.950 646.950 874.050 649.050 ;
        RECT 868.950 643.950 871.050 646.050 ;
        RECT 872.100 645.150 873.900 646.950 ;
        RECT 875.100 646.050 876.900 647.850 ;
        RECT 887.100 646.050 888.900 647.850 ;
        RECT 889.950 646.950 892.050 649.050 ;
        RECT 874.950 643.950 877.050 646.050 ;
        RECT 886.950 643.950 889.050 646.050 ;
        RECT 890.100 645.150 891.900 646.950 ;
        RECT 893.100 646.050 894.900 647.850 ;
        RECT 895.950 646.950 898.050 649.050 ;
        RECT 892.950 643.950 895.050 646.050 ;
        RECT 896.400 634.800 897.300 646.950 ;
        RECT 866.700 633.900 873.300 634.800 ;
        RECT 866.700 633.600 867.600 633.900 ;
        RECT 856.950 628.950 859.050 631.050 ;
        RECT 865.800 627.600 867.600 633.600 ;
        RECT 871.800 633.600 873.300 633.900 ;
        RECT 890.700 633.900 897.300 634.800 ;
        RECT 890.700 633.600 892.200 633.900 ;
        RECT 871.800 627.600 873.600 633.600 ;
        RECT 890.400 627.600 892.200 633.600 ;
        RECT 896.400 633.600 897.300 633.900 ;
        RECT 896.400 627.600 898.200 633.600 ;
        RECT 16.800 617.400 18.600 623.400 ;
        RECT 34.800 617.400 36.600 623.400 ;
        RECT 13.950 604.950 16.050 607.050 ;
        RECT 14.100 603.150 15.900 604.950 ;
        RECT 17.400 604.050 18.600 617.400 ;
        RECT 35.700 617.100 36.600 617.400 ;
        RECT 40.800 617.400 42.600 623.400 ;
        RECT 61.800 617.400 63.600 623.400 ;
        RECT 40.800 617.100 42.300 617.400 ;
        RECT 35.700 616.200 42.300 617.100 ;
        RECT 19.950 604.950 22.050 607.050 ;
        RECT 16.950 601.950 19.050 604.050 ;
        RECT 20.100 603.150 21.900 604.950 ;
        RECT 35.700 604.050 36.600 616.200 ;
        RECT 37.950 604.950 40.050 607.050 ;
        RECT 34.950 601.950 37.050 604.050 ;
        RECT 38.100 603.150 39.900 604.950 ;
        RECT 41.100 604.050 42.900 605.850 ;
        RECT 43.950 604.950 46.050 607.050 ;
        RECT 58.950 604.950 61.050 607.050 ;
        RECT 40.950 601.950 43.050 604.050 ;
        RECT 44.100 603.150 45.900 604.950 ;
        RECT 59.100 603.150 60.900 604.950 ;
        RECT 62.400 604.050 63.600 617.400 ;
        RECT 73.950 616.950 76.050 619.050 ;
        RECT 83.400 617.400 85.200 623.400 ;
        RECT 64.950 604.950 67.050 607.050 ;
        RECT 61.950 601.950 64.050 604.050 ;
        RECT 65.100 603.150 66.900 604.950 ;
        RECT 70.950 601.950 73.050 604.050 ;
        RECT 74.550 603.450 75.450 616.950 ;
        RECT 79.950 604.950 82.050 607.050 ;
        RECT 74.550 603.000 78.450 603.450 ;
        RECT 80.100 603.150 81.900 604.950 ;
        RECT 83.850 604.050 85.050 617.400 ;
        RECT 92.550 611.400 94.350 623.400 ;
        RECT 100.050 617.400 101.850 623.400 ;
        RECT 97.950 615.300 101.850 617.400 ;
        RECT 107.850 616.500 109.650 623.400 ;
        RECT 115.650 617.400 117.450 623.400 ;
        RECT 116.250 616.500 117.450 617.400 ;
        RECT 106.950 615.450 113.550 616.500 ;
        RECT 106.950 614.700 108.750 615.450 ;
        RECT 111.750 614.700 113.550 615.450 ;
        RECT 116.250 614.400 121.050 616.500 ;
        RECT 99.150 612.600 101.850 614.400 ;
        RECT 102.750 613.800 104.550 614.400 ;
        RECT 102.750 612.900 109.050 613.800 ;
        RECT 116.250 613.500 117.450 614.400 ;
        RECT 102.750 612.600 104.550 612.900 ;
        RECT 100.950 611.700 101.850 612.600 ;
        RECT 85.950 604.950 88.050 607.050 ;
        RECT 74.550 602.550 79.050 603.000 ;
        RECT 17.400 596.700 18.600 601.950 ;
        RECT 35.700 598.200 36.600 601.950 ;
        RECT 35.700 597.000 39.000 598.200 ;
        RECT 14.400 595.800 18.600 596.700 ;
        RECT 14.400 588.600 16.200 595.800 ;
        RECT 37.200 588.600 39.000 597.000 ;
        RECT 62.400 596.700 63.600 601.950 ;
        RECT 59.400 595.800 63.600 596.700 ;
        RECT 59.400 588.600 61.200 595.800 ;
        RECT 71.550 595.050 72.450 601.950 ;
        RECT 76.950 601.050 79.050 602.550 ;
        RECT 82.950 601.950 85.050 604.050 ;
        RECT 86.100 603.150 87.900 604.950 ;
        RECT 89.100 604.050 90.900 605.850 ;
        RECT 92.550 604.050 93.750 611.400 ;
        RECT 97.950 610.800 100.050 611.700 ;
        RECT 100.950 610.800 106.050 611.700 ;
        RECT 95.850 609.600 100.050 610.800 ;
        RECT 94.950 607.800 96.750 609.600 ;
        RECT 88.950 601.950 91.050 604.050 ;
        RECT 92.550 603.750 97.050 604.050 ;
        RECT 92.550 601.950 98.850 603.750 ;
        RECT 76.950 600.000 79.200 601.050 ;
        RECT 77.100 598.950 79.200 600.000 ;
        RECT 82.950 597.750 84.150 601.950 ;
        RECT 80.400 596.700 84.150 597.750 ;
        RECT 70.950 592.950 73.050 595.050 ;
        RECT 80.400 594.600 81.600 596.700 ;
        RECT 79.800 588.600 81.600 594.600 ;
        RECT 82.800 593.700 90.600 595.050 ;
        RECT 82.800 588.600 84.600 593.700 ;
        RECT 88.800 588.600 90.600 593.700 ;
        RECT 92.550 594.600 93.750 601.950 ;
        RECT 105.150 598.200 106.050 610.800 ;
        RECT 108.150 610.800 109.050 612.900 ;
        RECT 109.950 612.300 117.450 613.500 ;
        RECT 109.950 611.700 111.750 612.300 ;
        RECT 124.050 611.400 125.850 623.400 ;
        RECT 143.400 617.400 145.200 623.400 ;
        RECT 108.150 610.500 116.550 610.800 ;
        RECT 124.950 610.500 125.850 611.400 ;
        RECT 127.950 610.950 130.050 613.050 ;
        RECT 108.150 609.900 125.850 610.500 ;
        RECT 114.750 609.300 125.850 609.900 ;
        RECT 114.750 609.000 116.550 609.300 ;
        RECT 112.950 602.400 115.050 604.050 ;
        RECT 112.950 601.200 120.900 602.400 ;
        RECT 121.950 601.950 124.050 604.050 ;
        RECT 119.100 600.600 120.900 601.200 ;
        RECT 122.100 600.150 123.900 601.950 ;
        RECT 116.100 599.400 117.900 600.000 ;
        RECT 122.100 599.400 123.000 600.150 ;
        RECT 116.100 598.200 123.000 599.400 ;
        RECT 105.150 597.000 117.150 598.200 ;
        RECT 105.150 596.400 106.950 597.000 ;
        RECT 116.100 595.200 117.150 597.000 ;
        RECT 92.550 588.600 94.350 594.600 ;
        RECT 97.950 593.700 100.050 594.600 ;
        RECT 97.950 592.500 101.700 593.700 ;
        RECT 112.350 593.550 114.150 594.300 ;
        RECT 100.650 591.600 101.700 592.500 ;
        RECT 109.200 592.500 114.150 593.550 ;
        RECT 115.650 593.400 117.450 595.200 ;
        RECT 124.950 594.600 125.850 609.300 ;
        RECT 128.550 601.050 129.450 610.950 ;
        RECT 139.950 604.950 142.050 607.050 ;
        RECT 140.100 603.150 141.900 604.950 ;
        RECT 143.850 604.050 145.050 617.400 ;
        RECT 153.150 611.400 154.950 623.400 ;
        RECT 161.550 617.400 163.350 623.400 ;
        RECT 161.550 616.500 162.750 617.400 ;
        RECT 169.350 616.500 171.150 623.400 ;
        RECT 177.150 617.400 178.950 623.400 ;
        RECT 157.950 614.400 162.750 616.500 ;
        RECT 165.450 615.450 172.050 616.500 ;
        RECT 165.450 614.700 167.250 615.450 ;
        RECT 170.250 614.700 172.050 615.450 ;
        RECT 177.150 615.300 181.050 617.400 ;
        RECT 161.550 613.500 162.750 614.400 ;
        RECT 174.450 613.800 176.250 614.400 ;
        RECT 161.550 612.300 169.050 613.500 ;
        RECT 167.250 611.700 169.050 612.300 ;
        RECT 169.950 612.900 176.250 613.800 ;
        RECT 153.150 610.500 154.050 611.400 ;
        RECT 169.950 610.800 170.850 612.900 ;
        RECT 174.450 612.600 176.250 612.900 ;
        RECT 177.150 612.600 179.850 614.400 ;
        RECT 177.150 611.700 178.050 612.600 ;
        RECT 162.450 610.500 170.850 610.800 ;
        RECT 153.150 609.900 170.850 610.500 ;
        RECT 172.950 610.800 178.050 611.700 ;
        RECT 178.950 610.800 181.050 611.700 ;
        RECT 184.650 611.400 186.450 623.400 ;
        RECT 203.400 617.400 205.200 623.400 ;
        RECT 224.400 617.400 226.200 623.400 ;
        RECT 232.800 619.950 234.900 622.050 ;
        RECT 153.150 609.300 164.250 609.900 ;
        RECT 145.950 604.950 148.050 607.050 ;
        RECT 142.950 601.950 145.050 604.050 ;
        RECT 146.100 603.150 147.900 604.950 ;
        RECT 149.100 604.050 150.900 605.850 ;
        RECT 148.950 601.950 151.050 604.050 ;
        RECT 127.950 598.950 130.050 601.050 ;
        RECT 142.950 597.750 144.150 601.950 ;
        RECT 140.400 596.700 144.150 597.750 ;
        RECT 140.400 594.600 141.600 596.700 ;
        RECT 118.950 592.500 121.050 594.600 ;
        RECT 109.200 591.600 110.250 592.500 ;
        RECT 118.950 591.600 120.000 592.500 ;
        RECT 100.650 588.600 102.450 591.600 ;
        RECT 108.450 588.600 110.250 591.600 ;
        RECT 116.250 590.700 120.000 591.600 ;
        RECT 116.250 588.600 118.050 590.700 ;
        RECT 124.050 588.600 125.850 594.600 ;
        RECT 139.800 588.600 141.600 594.600 ;
        RECT 142.800 593.700 150.600 595.050 ;
        RECT 142.800 588.600 144.600 593.700 ;
        RECT 148.800 588.600 150.600 593.700 ;
        RECT 153.150 594.600 154.050 609.300 ;
        RECT 162.450 609.000 164.250 609.300 ;
        RECT 154.950 601.950 157.050 604.050 ;
        RECT 163.950 602.400 166.050 604.050 ;
        RECT 155.100 600.150 156.900 601.950 ;
        RECT 158.100 601.200 166.050 602.400 ;
        RECT 158.100 600.600 159.900 601.200 ;
        RECT 156.000 599.400 156.900 600.150 ;
        RECT 161.100 599.400 162.900 600.000 ;
        RECT 156.000 598.200 162.900 599.400 ;
        RECT 172.950 598.200 173.850 610.800 ;
        RECT 178.950 609.600 183.150 610.800 ;
        RECT 182.250 607.800 184.050 609.600 ;
        RECT 185.250 604.050 186.450 611.400 ;
        RECT 199.950 604.950 202.050 607.050 ;
        RECT 181.950 603.750 186.450 604.050 ;
        RECT 180.150 601.950 186.450 603.750 ;
        RECT 200.100 603.150 201.900 604.950 ;
        RECT 203.850 604.050 205.050 617.400 ;
        RECT 205.950 604.950 208.050 607.050 ;
        RECT 161.850 597.000 173.850 598.200 ;
        RECT 161.850 595.200 162.900 597.000 ;
        RECT 172.050 596.400 173.850 597.000 ;
        RECT 153.150 588.600 154.950 594.600 ;
        RECT 157.950 592.500 160.050 594.600 ;
        RECT 161.550 593.400 163.350 595.200 ;
        RECT 185.250 594.600 186.450 601.950 ;
        RECT 202.950 601.950 205.050 604.050 ;
        RECT 206.100 603.150 207.900 604.950 ;
        RECT 209.100 604.050 210.900 605.850 ;
        RECT 220.950 604.950 223.050 607.050 ;
        RECT 208.950 601.950 211.050 604.050 ;
        RECT 221.100 603.150 222.900 604.950 ;
        RECT 224.400 604.050 225.600 617.400 ;
        RECT 226.950 604.950 229.050 607.050 ;
        RECT 223.950 601.950 226.050 604.050 ;
        RECT 227.100 603.150 228.900 604.950 ;
        RECT 202.950 597.750 204.150 601.950 ;
        RECT 200.400 596.700 204.150 597.750 ;
        RECT 224.400 596.700 225.600 601.950 ;
        RECT 200.400 594.600 201.600 596.700 ;
        RECT 224.400 595.800 228.600 596.700 ;
        RECT 164.850 593.550 166.650 594.300 ;
        RECT 178.950 593.700 181.050 594.600 ;
        RECT 164.850 592.500 169.800 593.550 ;
        RECT 159.000 591.600 160.050 592.500 ;
        RECT 168.750 591.600 169.800 592.500 ;
        RECT 177.300 592.500 181.050 593.700 ;
        RECT 177.300 591.600 178.350 592.500 ;
        RECT 159.000 590.700 162.750 591.600 ;
        RECT 160.950 588.600 162.750 590.700 ;
        RECT 168.750 588.600 170.550 591.600 ;
        RECT 176.550 588.600 178.350 591.600 ;
        RECT 184.650 588.600 186.450 594.600 ;
        RECT 199.800 588.600 201.600 594.600 ;
        RECT 202.800 593.700 210.600 595.050 ;
        RECT 202.800 588.600 204.600 593.700 ;
        RECT 208.800 588.600 210.600 593.700 ;
        RECT 226.800 588.600 228.600 595.800 ;
        RECT 233.550 592.050 234.450 619.950 ;
        RECT 245.400 617.400 247.200 623.400 ;
        RECT 266.400 617.400 268.200 623.400 ;
        RECT 287.400 617.400 289.200 623.400 ;
        RECT 241.950 604.950 244.050 607.050 ;
        RECT 242.100 603.150 243.900 604.950 ;
        RECT 245.400 604.050 246.600 617.400 ;
        RECT 247.950 604.950 250.050 607.050 ;
        RECT 262.950 604.950 265.050 607.050 ;
        RECT 244.950 601.950 247.050 604.050 ;
        RECT 248.100 603.150 249.900 604.950 ;
        RECT 263.100 603.150 264.900 604.950 ;
        RECT 266.400 604.050 267.600 617.400 ;
        RECT 268.950 604.950 271.050 607.050 ;
        RECT 265.950 601.950 268.050 604.050 ;
        RECT 269.100 603.150 270.900 604.950 ;
        RECT 283.950 601.950 286.050 604.050 ;
        RECT 245.400 596.700 246.600 601.950 ;
        RECT 266.400 596.700 267.600 601.950 ;
        RECT 284.100 600.150 285.900 601.950 ;
        RECT 287.400 597.300 288.300 617.400 ;
        RECT 293.700 611.400 295.500 623.400 ;
        RECT 310.800 617.400 312.600 623.400 ;
        RECT 311.700 617.100 312.600 617.400 ;
        RECT 316.800 617.400 318.600 623.400 ;
        RECT 338.400 617.400 340.200 623.400 ;
        RECT 346.950 619.950 349.050 622.050 ;
        RECT 316.800 617.100 318.300 617.400 ;
        RECT 311.700 616.200 318.300 617.100 ;
        RECT 290.100 604.050 291.900 605.850 ;
        RECT 293.700 604.050 294.600 611.400 ;
        RECT 311.700 604.050 312.600 616.200 ;
        RECT 325.800 613.950 327.900 616.050 ;
        RECT 313.950 604.950 316.050 607.050 ;
        RECT 289.950 601.950 292.050 604.050 ;
        RECT 292.950 601.950 295.050 604.050 ;
        RECT 310.950 601.950 313.050 604.050 ;
        RECT 314.100 603.150 315.900 604.950 ;
        RECT 317.100 604.050 318.900 605.850 ;
        RECT 319.950 604.950 322.050 607.050 ;
        RECT 316.950 601.950 319.050 604.050 ;
        RECT 320.100 603.150 321.900 604.950 ;
        RECT 245.400 595.800 249.600 596.700 ;
        RECT 266.400 595.800 270.600 596.700 ;
        RECT 232.950 589.950 235.050 592.050 ;
        RECT 247.800 588.600 249.600 595.800 ;
        RECT 268.800 588.600 270.600 595.800 ;
        RECT 284.400 596.400 291.900 597.300 ;
        RECT 284.400 588.600 286.200 596.400 ;
        RECT 290.100 595.500 291.900 596.400 ;
        RECT 293.700 594.600 294.600 601.950 ;
        RECT 311.700 598.200 312.600 601.950 ;
        RECT 311.700 597.000 315.000 598.200 ;
        RECT 291.900 592.800 294.600 594.600 ;
        RECT 291.900 588.600 293.700 592.800 ;
        RECT 313.200 588.600 315.000 597.000 ;
        RECT 326.550 592.050 327.450 613.950 ;
        RECT 334.950 604.950 337.050 607.050 ;
        RECT 335.100 603.150 336.900 604.950 ;
        RECT 338.850 604.050 340.050 617.400 ;
        RECT 347.550 613.050 348.450 619.950 ;
        RECT 361.800 617.400 363.600 623.400 ;
        RECT 373.950 619.950 376.050 622.050 ;
        RECT 346.950 610.950 349.050 613.050 ;
        RECT 340.950 604.950 343.050 607.050 ;
        RECT 337.950 601.950 340.050 604.050 ;
        RECT 341.100 603.150 342.900 604.950 ;
        RECT 344.100 604.050 345.900 605.850 ;
        RECT 356.100 604.050 357.900 605.850 ;
        RECT 358.950 604.950 361.050 607.050 ;
        RECT 343.950 601.950 346.050 604.050 ;
        RECT 355.950 601.950 358.050 604.050 ;
        RECT 359.100 603.150 360.900 604.950 ;
        RECT 361.950 604.050 363.150 617.400 ;
        RECT 364.950 604.950 367.050 607.050 ;
        RECT 361.950 601.950 364.050 604.050 ;
        RECT 365.100 603.150 366.900 604.950 ;
        RECT 337.950 597.750 339.150 601.950 ;
        RECT 335.400 596.700 339.150 597.750 ;
        RECT 362.850 597.750 364.050 601.950 ;
        RECT 362.850 596.700 366.600 597.750 ;
        RECT 335.400 594.600 336.600 596.700 ;
        RECT 325.950 589.950 328.050 592.050 ;
        RECT 334.800 588.600 336.600 594.600 ;
        RECT 337.800 593.700 345.600 595.050 ;
        RECT 337.800 588.600 339.600 593.700 ;
        RECT 343.800 588.600 345.600 593.700 ;
        RECT 356.400 593.700 364.200 595.050 ;
        RECT 356.400 588.600 358.200 593.700 ;
        RECT 362.400 588.600 364.200 593.700 ;
        RECT 365.400 594.600 366.600 596.700 ;
        RECT 374.550 595.050 375.450 619.950 ;
        RECT 382.800 617.400 384.600 623.400 ;
        RECT 383.700 617.100 384.600 617.400 ;
        RECT 388.800 617.400 390.600 623.400 ;
        RECT 388.800 617.100 390.300 617.400 ;
        RECT 383.700 616.200 390.300 617.100 ;
        RECT 383.700 604.050 384.600 616.200 ;
        RECT 406.800 611.400 408.600 623.400 ;
        RECT 409.800 612.300 411.600 623.400 ;
        RECT 415.800 612.300 417.600 623.400 ;
        RECT 409.800 611.400 417.600 612.300 ;
        RECT 420.150 611.400 421.950 623.400 ;
        RECT 428.550 617.400 430.350 623.400 ;
        RECT 428.550 616.500 429.750 617.400 ;
        RECT 436.350 616.500 438.150 623.400 ;
        RECT 444.150 617.400 445.950 623.400 ;
        RECT 424.950 614.400 429.750 616.500 ;
        RECT 432.450 615.450 439.050 616.500 ;
        RECT 432.450 614.700 434.250 615.450 ;
        RECT 437.250 614.700 439.050 615.450 ;
        RECT 444.150 615.300 448.050 617.400 ;
        RECT 428.550 613.500 429.750 614.400 ;
        RECT 441.450 613.800 443.250 614.400 ;
        RECT 428.550 612.300 436.050 613.500 ;
        RECT 434.250 611.700 436.050 612.300 ;
        RECT 436.950 612.900 443.250 613.800 ;
        RECT 385.950 604.950 388.050 607.050 ;
        RECT 382.950 601.950 385.050 604.050 ;
        RECT 386.100 603.150 387.900 604.950 ;
        RECT 389.100 604.050 390.900 605.850 ;
        RECT 391.950 604.950 394.050 607.050 ;
        RECT 388.950 601.950 391.050 604.050 ;
        RECT 392.100 603.150 393.900 604.950 ;
        RECT 407.400 604.050 408.600 611.400 ;
        RECT 420.150 610.500 421.050 611.400 ;
        RECT 436.950 610.800 437.850 612.900 ;
        RECT 441.450 612.600 443.250 612.900 ;
        RECT 444.150 612.600 446.850 614.400 ;
        RECT 444.150 611.700 445.050 612.600 ;
        RECT 429.450 610.500 437.850 610.800 ;
        RECT 420.150 609.900 437.850 610.500 ;
        RECT 439.950 610.800 445.050 611.700 ;
        RECT 445.950 610.800 448.050 611.700 ;
        RECT 451.650 611.400 453.450 623.400 ;
        RECT 457.950 619.950 460.050 622.050 ;
        RECT 420.150 609.300 431.250 609.900 ;
        RECT 409.950 604.950 412.050 607.050 ;
        RECT 406.950 601.950 409.050 604.050 ;
        RECT 410.100 603.150 411.900 604.950 ;
        RECT 413.100 604.050 414.900 605.850 ;
        RECT 415.950 604.950 418.050 607.050 ;
        RECT 412.950 601.950 415.050 604.050 ;
        RECT 416.100 603.150 417.900 604.950 ;
        RECT 383.700 598.200 384.600 601.950 ;
        RECT 383.700 597.000 387.000 598.200 ;
        RECT 365.400 588.600 367.200 594.600 ;
        RECT 373.950 592.950 376.050 595.050 ;
        RECT 385.200 588.600 387.000 597.000 ;
        RECT 407.400 594.600 408.600 601.950 ;
        RECT 420.150 594.600 421.050 609.300 ;
        RECT 429.450 609.000 431.250 609.300 ;
        RECT 421.950 601.950 424.050 604.050 ;
        RECT 430.950 602.400 433.050 604.050 ;
        RECT 422.100 600.150 423.900 601.950 ;
        RECT 425.100 601.200 433.050 602.400 ;
        RECT 425.100 600.600 426.900 601.200 ;
        RECT 423.000 599.400 423.900 600.150 ;
        RECT 428.100 599.400 429.900 600.000 ;
        RECT 423.000 598.200 429.900 599.400 ;
        RECT 439.950 598.200 440.850 610.800 ;
        RECT 445.950 609.600 450.150 610.800 ;
        RECT 449.250 607.800 451.050 609.600 ;
        RECT 452.250 604.050 453.450 611.400 ;
        RECT 448.950 603.750 453.450 604.050 ;
        RECT 447.150 601.950 453.450 603.750 ;
        RECT 428.850 597.000 440.850 598.200 ;
        RECT 428.850 595.200 429.900 597.000 ;
        RECT 439.050 596.400 440.850 597.000 ;
        RECT 407.400 593.400 412.500 594.600 ;
        RECT 410.700 588.600 412.500 593.400 ;
        RECT 420.150 588.600 421.950 594.600 ;
        RECT 424.950 592.500 427.050 594.600 ;
        RECT 428.550 593.400 430.350 595.200 ;
        RECT 452.250 594.600 453.450 601.950 ;
        RECT 458.550 595.050 459.450 619.950 ;
        RECT 464.400 612.300 466.200 623.400 ;
        RECT 470.400 612.300 472.200 623.400 ;
        RECT 464.400 611.400 472.200 612.300 ;
        RECT 473.400 611.400 475.200 623.400 ;
        RECT 494.400 617.400 496.200 623.400 ;
        RECT 463.950 604.950 466.050 607.050 ;
        RECT 464.100 603.150 465.900 604.950 ;
        RECT 467.100 604.050 468.900 605.850 ;
        RECT 469.950 604.950 472.050 607.050 ;
        RECT 466.950 601.950 469.050 604.050 ;
        RECT 470.100 603.150 471.900 604.950 ;
        RECT 473.400 604.050 474.600 611.400 ;
        RECT 490.950 604.950 493.050 607.050 ;
        RECT 472.950 601.950 475.050 604.050 ;
        RECT 491.100 603.150 492.900 604.950 ;
        RECT 494.850 604.050 496.050 617.400 ;
        RECT 504.150 611.400 505.950 623.400 ;
        RECT 512.550 617.400 514.350 623.400 ;
        RECT 512.550 616.500 513.750 617.400 ;
        RECT 520.350 616.500 522.150 623.400 ;
        RECT 528.150 617.400 529.950 623.400 ;
        RECT 508.950 614.400 513.750 616.500 ;
        RECT 516.450 615.450 523.050 616.500 ;
        RECT 516.450 614.700 518.250 615.450 ;
        RECT 521.250 614.700 523.050 615.450 ;
        RECT 528.150 615.300 532.050 617.400 ;
        RECT 512.550 613.500 513.750 614.400 ;
        RECT 525.450 613.800 527.250 614.400 ;
        RECT 512.550 612.300 520.050 613.500 ;
        RECT 518.250 611.700 520.050 612.300 ;
        RECT 520.950 612.900 527.250 613.800 ;
        RECT 504.150 610.500 505.050 611.400 ;
        RECT 520.950 610.800 521.850 612.900 ;
        RECT 525.450 612.600 527.250 612.900 ;
        RECT 528.150 612.600 530.850 614.400 ;
        RECT 528.150 611.700 529.050 612.600 ;
        RECT 513.450 610.500 521.850 610.800 ;
        RECT 504.150 609.900 521.850 610.500 ;
        RECT 523.950 610.800 529.050 611.700 ;
        RECT 529.950 610.800 532.050 611.700 ;
        RECT 535.650 611.400 537.450 623.400 ;
        RECT 550.800 611.400 552.600 623.400 ;
        RECT 553.800 612.300 555.600 623.400 ;
        RECT 559.800 612.300 561.600 623.400 ;
        RECT 574.800 617.400 576.600 623.400 ;
        RECT 575.700 617.100 576.600 617.400 ;
        RECT 580.800 617.400 582.600 623.400 ;
        RECT 602.400 617.400 604.200 623.400 ;
        RECT 625.800 617.400 627.600 623.400 ;
        RECT 643.800 617.400 645.600 623.400 ;
        RECT 580.800 617.100 582.300 617.400 ;
        RECT 575.700 616.200 582.300 617.100 ;
        RECT 568.950 613.950 571.050 616.050 ;
        RECT 553.800 611.400 561.600 612.300 ;
        RECT 504.150 609.300 515.250 609.900 ;
        RECT 496.950 604.950 499.050 607.050 ;
        RECT 493.950 601.950 496.050 604.050 ;
        RECT 497.100 603.150 498.900 604.950 ;
        RECT 500.100 604.050 501.900 605.850 ;
        RECT 499.950 601.950 502.050 604.050 ;
        RECT 431.850 593.550 433.650 594.300 ;
        RECT 445.950 593.700 448.050 594.600 ;
        RECT 431.850 592.500 436.800 593.550 ;
        RECT 426.000 591.600 427.050 592.500 ;
        RECT 435.750 591.600 436.800 592.500 ;
        RECT 444.300 592.500 448.050 593.700 ;
        RECT 444.300 591.600 445.350 592.500 ;
        RECT 426.000 590.700 429.750 591.600 ;
        RECT 427.950 588.600 429.750 590.700 ;
        RECT 435.750 588.600 437.550 591.600 ;
        RECT 443.550 588.600 445.350 591.600 ;
        RECT 451.650 588.600 453.450 594.600 ;
        RECT 457.950 592.950 460.050 595.050 ;
        RECT 473.400 594.600 474.600 601.950 ;
        RECT 493.950 597.750 495.150 601.950 ;
        RECT 491.400 596.700 495.150 597.750 ;
        RECT 491.400 594.600 492.600 596.700 ;
        RECT 469.500 593.400 474.600 594.600 ;
        RECT 469.500 588.600 471.300 593.400 ;
        RECT 490.800 588.600 492.600 594.600 ;
        RECT 493.800 593.700 501.600 595.050 ;
        RECT 493.800 588.600 495.600 593.700 ;
        RECT 499.800 588.600 501.600 593.700 ;
        RECT 504.150 594.600 505.050 609.300 ;
        RECT 513.450 609.000 515.250 609.300 ;
        RECT 505.950 601.950 508.050 604.050 ;
        RECT 514.950 602.400 517.050 604.050 ;
        RECT 506.100 600.150 507.900 601.950 ;
        RECT 509.100 601.200 517.050 602.400 ;
        RECT 509.100 600.600 510.900 601.200 ;
        RECT 507.000 599.400 507.900 600.150 ;
        RECT 512.100 599.400 513.900 600.000 ;
        RECT 507.000 598.200 513.900 599.400 ;
        RECT 523.950 598.200 524.850 610.800 ;
        RECT 529.950 609.600 534.150 610.800 ;
        RECT 533.250 607.800 535.050 609.600 ;
        RECT 536.250 604.050 537.450 611.400 ;
        RECT 551.400 604.050 552.600 611.400 ;
        RECT 553.950 604.950 556.050 607.050 ;
        RECT 532.950 603.750 537.450 604.050 ;
        RECT 531.150 601.950 537.450 603.750 ;
        RECT 550.950 601.950 553.050 604.050 ;
        RECT 554.100 603.150 555.900 604.950 ;
        RECT 557.100 604.050 558.900 605.850 ;
        RECT 559.950 604.950 562.050 607.050 ;
        RECT 556.950 601.950 559.050 604.050 ;
        RECT 560.100 603.150 561.900 604.950 ;
        RECT 512.850 597.000 524.850 598.200 ;
        RECT 512.850 595.200 513.900 597.000 ;
        RECT 523.050 596.400 524.850 597.000 ;
        RECT 504.150 588.600 505.950 594.600 ;
        RECT 508.950 592.500 511.050 594.600 ;
        RECT 512.550 593.400 514.350 595.200 ;
        RECT 536.250 594.600 537.450 601.950 ;
        RECT 515.850 593.550 517.650 594.300 ;
        RECT 529.950 593.700 532.050 594.600 ;
        RECT 515.850 592.500 520.800 593.550 ;
        RECT 510.000 591.600 511.050 592.500 ;
        RECT 519.750 591.600 520.800 592.500 ;
        RECT 528.300 592.500 532.050 593.700 ;
        RECT 528.300 591.600 529.350 592.500 ;
        RECT 510.000 590.700 513.750 591.600 ;
        RECT 511.950 588.600 513.750 590.700 ;
        RECT 519.750 588.600 521.550 591.600 ;
        RECT 527.550 588.600 529.350 591.600 ;
        RECT 535.650 588.600 537.450 594.600 ;
        RECT 551.400 594.600 552.600 601.950 ;
        RECT 551.400 593.400 556.500 594.600 ;
        RECT 554.700 588.600 556.500 593.400 ;
        RECT 569.550 592.050 570.450 613.950 ;
        RECT 575.700 604.050 576.600 616.200 ;
        RECT 577.950 604.950 580.050 607.050 ;
        RECT 574.950 601.950 577.050 604.050 ;
        RECT 578.100 603.150 579.900 604.950 ;
        RECT 581.100 604.050 582.900 605.850 ;
        RECT 583.950 604.950 586.050 607.050 ;
        RECT 598.950 604.950 601.050 607.050 ;
        RECT 580.950 601.950 583.050 604.050 ;
        RECT 584.100 603.150 585.900 604.950 ;
        RECT 599.100 603.150 600.900 604.950 ;
        RECT 602.850 604.050 604.050 617.400 ;
        RECT 604.950 604.950 607.050 607.050 ;
        RECT 601.950 601.950 604.050 604.050 ;
        RECT 605.100 603.150 606.900 604.950 ;
        RECT 608.100 604.050 609.900 605.850 ;
        RECT 622.950 604.950 625.050 607.050 ;
        RECT 607.950 601.950 610.050 604.050 ;
        RECT 623.100 603.150 624.900 604.950 ;
        RECT 626.400 604.050 627.600 617.400 ;
        RECT 644.700 617.100 645.600 617.400 ;
        RECT 649.800 617.400 651.600 623.400 ;
        RECT 668.400 617.400 670.200 623.400 ;
        RECT 692.400 617.400 694.200 623.400 ;
        RECT 715.800 617.400 717.600 623.400 ;
        RECT 737.400 617.400 739.200 623.400 ;
        RECT 758.400 617.400 760.200 623.400 ;
        RECT 781.800 617.400 783.600 623.400 ;
        RECT 790.800 619.950 792.900 622.050 ;
        RECT 794.100 619.950 796.200 622.050 ;
        RECT 649.800 617.100 651.300 617.400 ;
        RECT 644.700 616.200 651.300 617.100 ;
        RECT 634.950 613.950 637.050 616.050 ;
        RECT 628.950 604.950 631.050 607.050 ;
        RECT 625.950 601.950 628.050 604.050 ;
        RECT 629.100 603.150 630.900 604.950 ;
        RECT 575.700 598.200 576.600 601.950 ;
        RECT 575.700 597.000 579.000 598.200 ;
        RECT 601.950 597.750 603.150 601.950 ;
        RECT 568.950 589.950 571.050 592.050 ;
        RECT 577.200 588.600 579.000 597.000 ;
        RECT 599.400 596.700 603.150 597.750 ;
        RECT 626.400 596.700 627.600 601.950 ;
        RECT 599.400 594.600 600.600 596.700 ;
        RECT 623.400 595.800 627.600 596.700 ;
        RECT 598.800 588.600 600.600 594.600 ;
        RECT 601.800 593.700 609.600 595.050 ;
        RECT 601.800 588.600 603.600 593.700 ;
        RECT 607.800 588.600 609.600 593.700 ;
        RECT 623.400 588.600 625.200 595.800 ;
        RECT 635.550 592.050 636.450 613.950 ;
        RECT 644.700 604.050 645.600 616.200 ;
        RECT 646.950 604.950 649.050 607.050 ;
        RECT 643.950 601.950 646.050 604.050 ;
        RECT 647.100 603.150 648.900 604.950 ;
        RECT 650.100 604.050 651.900 605.850 ;
        RECT 652.950 604.950 655.050 607.050 ;
        RECT 664.950 604.950 667.050 607.050 ;
        RECT 649.950 601.950 652.050 604.050 ;
        RECT 653.100 603.150 654.900 604.950 ;
        RECT 665.100 603.150 666.900 604.950 ;
        RECT 668.400 604.050 669.600 617.400 ;
        RECT 670.950 604.950 673.050 607.050 ;
        RECT 688.950 604.950 691.050 607.050 ;
        RECT 667.950 601.950 670.050 604.050 ;
        RECT 671.100 603.150 672.900 604.950 ;
        RECT 689.100 603.150 690.900 604.950 ;
        RECT 692.850 604.050 694.050 617.400 ;
        RECT 694.950 604.950 697.050 607.050 ;
        RECT 691.950 601.950 694.050 604.050 ;
        RECT 695.100 603.150 696.900 604.950 ;
        RECT 698.100 604.050 699.900 605.850 ;
        RECT 710.100 604.050 711.900 605.850 ;
        RECT 712.950 604.950 715.050 607.050 ;
        RECT 697.950 601.950 700.050 604.050 ;
        RECT 709.950 601.950 712.050 604.050 ;
        RECT 713.100 603.150 714.900 604.950 ;
        RECT 715.950 604.050 717.150 617.400 ;
        RECT 718.950 604.950 721.050 607.050 ;
        RECT 733.950 604.950 736.050 607.050 ;
        RECT 715.950 601.950 718.050 604.050 ;
        RECT 719.100 603.150 720.900 604.950 ;
        RECT 734.100 603.150 735.900 604.950 ;
        RECT 737.400 604.050 738.600 617.400 ;
        RECT 739.950 604.950 742.050 607.050 ;
        RECT 754.950 604.950 757.050 607.050 ;
        RECT 736.950 601.950 739.050 604.050 ;
        RECT 740.100 603.150 741.900 604.950 ;
        RECT 755.100 603.150 756.900 604.950 ;
        RECT 758.400 604.050 759.600 617.400 ;
        RECT 760.950 604.950 763.050 607.050 ;
        RECT 757.950 601.950 760.050 604.050 ;
        RECT 761.100 603.150 762.900 604.950 ;
        RECT 776.100 604.050 777.900 605.850 ;
        RECT 778.950 604.950 781.050 607.050 ;
        RECT 775.950 601.950 778.050 604.050 ;
        RECT 779.100 603.150 780.900 604.950 ;
        RECT 781.950 604.050 783.150 617.400 ;
        RECT 791.550 613.050 792.450 619.950 ;
        RECT 790.950 610.950 793.050 613.050 ;
        RECT 784.950 604.950 787.050 607.050 ;
        RECT 781.950 601.950 784.050 604.050 ;
        RECT 785.100 603.150 786.900 604.950 ;
        RECT 644.700 598.200 645.600 601.950 ;
        RECT 644.700 597.000 648.000 598.200 ;
        RECT 634.950 589.950 637.050 592.050 ;
        RECT 646.200 588.600 648.000 597.000 ;
        RECT 668.400 596.700 669.600 601.950 ;
        RECT 691.950 597.750 693.150 601.950 ;
        RECT 689.400 596.700 693.150 597.750 ;
        RECT 716.850 597.750 718.050 601.950 ;
        RECT 716.850 596.700 720.600 597.750 ;
        RECT 668.400 595.800 672.600 596.700 ;
        RECT 670.800 588.600 672.600 595.800 ;
        RECT 689.400 594.600 690.600 596.700 ;
        RECT 688.800 588.600 690.600 594.600 ;
        RECT 691.800 593.700 699.600 595.050 ;
        RECT 691.800 588.600 693.600 593.700 ;
        RECT 697.800 588.600 699.600 593.700 ;
        RECT 710.400 593.700 718.200 595.050 ;
        RECT 710.400 588.600 712.200 593.700 ;
        RECT 716.400 588.600 718.200 593.700 ;
        RECT 719.400 594.600 720.600 596.700 ;
        RECT 737.400 596.700 738.600 601.950 ;
        RECT 758.400 596.700 759.600 601.950 ;
        RECT 782.850 597.750 784.050 601.950 ;
        RECT 790.950 598.950 793.050 601.050 ;
        RECT 782.850 596.700 786.600 597.750 ;
        RECT 737.400 595.800 741.600 596.700 ;
        RECT 758.400 595.800 762.600 596.700 ;
        RECT 719.400 588.600 721.200 594.600 ;
        RECT 739.800 588.600 741.600 595.800 ;
        RECT 760.800 588.600 762.600 595.800 ;
        RECT 776.400 593.700 784.200 595.050 ;
        RECT 776.400 588.600 778.200 593.700 ;
        RECT 782.400 588.600 784.200 593.700 ;
        RECT 785.400 594.600 786.600 596.700 ;
        RECT 785.400 588.600 787.200 594.600 ;
        RECT 791.550 592.050 792.450 598.950 ;
        RECT 794.550 595.050 795.450 619.950 ;
        RECT 805.800 617.400 807.600 623.400 ;
        RECT 829.800 617.400 831.600 623.400 ;
        RECT 800.100 604.050 801.900 605.850 ;
        RECT 802.950 604.950 805.050 607.050 ;
        RECT 799.950 601.950 802.050 604.050 ;
        RECT 803.100 603.150 804.900 604.950 ;
        RECT 805.950 604.050 807.150 617.400 ;
        RECT 817.950 613.950 820.050 616.050 ;
        RECT 808.950 604.950 811.050 607.050 ;
        RECT 805.950 601.950 808.050 604.050 ;
        RECT 809.100 603.150 810.900 604.950 ;
        RECT 806.850 597.750 808.050 601.950 ;
        RECT 806.850 596.700 810.600 597.750 ;
        RECT 793.950 592.950 796.050 595.050 ;
        RECT 800.400 593.700 808.200 595.050 ;
        RECT 790.950 589.950 793.050 592.050 ;
        RECT 800.400 588.600 802.200 593.700 ;
        RECT 806.400 588.600 808.200 593.700 ;
        RECT 809.400 594.600 810.600 596.700 ;
        RECT 818.550 595.050 819.450 613.950 ;
        RECT 824.100 604.050 825.900 605.850 ;
        RECT 826.950 604.950 829.050 607.050 ;
        RECT 823.950 601.950 826.050 604.050 ;
        RECT 827.100 603.150 828.900 604.950 ;
        RECT 829.950 604.050 831.150 617.400 ;
        RECT 838.950 616.950 841.050 619.050 ;
        RECT 851.400 617.400 853.200 623.400 ;
        RECT 832.950 604.950 835.050 607.050 ;
        RECT 829.950 601.950 832.050 604.050 ;
        RECT 833.100 603.150 834.900 604.950 ;
        RECT 830.850 597.750 832.050 601.950 ;
        RECT 830.850 596.700 834.600 597.750 ;
        RECT 809.400 588.600 811.200 594.600 ;
        RECT 817.950 592.950 820.050 595.050 ;
        RECT 824.400 593.700 832.200 595.050 ;
        RECT 824.400 588.600 826.200 593.700 ;
        RECT 830.400 588.600 832.200 593.700 ;
        RECT 833.400 594.600 834.600 596.700 ;
        RECT 833.400 588.600 835.200 594.600 ;
        RECT 839.550 592.050 840.450 616.950 ;
        RECT 847.950 604.950 850.050 607.050 ;
        RECT 848.100 603.150 849.900 604.950 ;
        RECT 851.400 604.050 852.600 617.400 ;
        RECT 865.950 613.950 868.050 616.050 ;
        RECT 853.950 604.950 856.050 607.050 ;
        RECT 850.950 601.950 853.050 604.050 ;
        RECT 854.100 603.150 855.900 604.950 ;
        RECT 851.400 596.700 852.600 601.950 ;
        RECT 866.550 601.050 867.450 613.950 ;
        RECT 871.800 611.400 873.600 623.400 ;
        RECT 874.800 612.300 876.600 623.400 ;
        RECT 880.800 612.300 882.600 623.400 ;
        RECT 886.950 619.950 889.050 622.050 ;
        RECT 874.800 611.400 882.600 612.300 ;
        RECT 872.400 604.050 873.600 611.400 ;
        RECT 874.950 604.950 877.050 607.050 ;
        RECT 871.950 601.950 874.050 604.050 ;
        RECT 875.100 603.150 876.900 604.950 ;
        RECT 878.100 604.050 879.900 605.850 ;
        RECT 880.950 604.950 883.050 607.050 ;
        RECT 877.950 601.950 880.050 604.050 ;
        RECT 881.100 603.150 882.900 604.950 ;
        RECT 865.800 598.950 867.900 601.050 ;
        RECT 851.400 595.800 855.600 596.700 ;
        RECT 838.950 589.950 841.050 592.050 ;
        RECT 853.800 588.600 855.600 595.800 ;
        RECT 872.400 594.600 873.600 601.950 ;
        RECT 872.400 593.400 877.500 594.600 ;
        RECT 875.700 588.600 877.500 593.400 ;
        RECT 887.550 592.050 888.450 619.950 ;
        RECT 896.400 617.400 898.200 623.400 ;
        RECT 896.700 617.100 898.200 617.400 ;
        RECT 902.400 617.400 904.200 623.400 ;
        RECT 902.400 617.100 903.300 617.400 ;
        RECT 896.700 616.200 903.300 617.100 ;
        RECT 892.950 604.950 895.050 607.050 ;
        RECT 893.100 603.150 894.900 604.950 ;
        RECT 896.100 604.050 897.900 605.850 ;
        RECT 898.950 604.950 901.050 607.050 ;
        RECT 895.950 601.950 898.050 604.050 ;
        RECT 899.100 603.150 900.900 604.950 ;
        RECT 902.400 604.050 903.300 616.200 ;
        RECT 901.950 601.950 904.050 604.050 ;
        RECT 902.400 598.200 903.300 601.950 ;
        RECT 900.000 597.000 903.300 598.200 ;
        RECT 886.950 589.950 889.050 592.050 ;
        RECT 900.000 588.600 901.800 597.000 ;
        RECT 1.800 580.950 3.900 583.050 ;
        RECT 2.550 577.050 3.450 580.950 ;
        RECT 14.400 577.200 16.200 584.400 ;
        RECT 1.950 574.950 4.050 577.050 ;
        RECT 14.400 576.300 18.600 577.200 ;
        RECT 17.400 571.050 18.600 576.300 ;
        RECT 39.000 576.000 40.800 584.400 ;
        RECT 59.400 577.200 61.200 584.400 ;
        RECT 80.400 577.200 82.200 584.400 ;
        RECT 91.950 580.950 94.050 583.050 ;
        RECT 59.400 576.300 63.600 577.200 ;
        RECT 80.400 576.300 84.600 577.200 ;
        RECT 39.000 574.800 42.300 576.000 ;
        RECT 41.400 571.050 42.300 574.800 ;
        RECT 46.950 571.950 49.050 574.050 ;
        RECT 14.100 568.050 15.900 569.850 ;
        RECT 16.950 568.950 19.050 571.050 ;
        RECT 13.950 565.950 16.050 568.050 ;
        RECT 17.400 555.600 18.600 568.950 ;
        RECT 20.100 568.050 21.900 569.850 ;
        RECT 32.100 568.050 33.900 569.850 ;
        RECT 34.950 568.950 37.050 571.050 ;
        RECT 19.950 565.950 22.050 568.050 ;
        RECT 31.950 565.950 34.050 568.050 ;
        RECT 35.100 567.150 36.900 568.950 ;
        RECT 38.100 568.050 39.900 569.850 ;
        RECT 40.950 568.950 43.050 571.050 ;
        RECT 37.950 565.950 40.050 568.050 ;
        RECT 41.400 556.800 42.300 568.950 ;
        RECT 47.550 559.050 48.450 571.950 ;
        RECT 62.400 571.050 63.600 576.300 ;
        RECT 83.400 571.050 84.600 576.300 ;
        RECT 59.100 568.050 60.900 569.850 ;
        RECT 61.950 568.950 64.050 571.050 ;
        RECT 58.950 565.950 61.050 568.050 ;
        RECT 46.950 556.950 49.050 559.050 ;
        RECT 35.700 555.900 42.300 556.800 ;
        RECT 35.700 555.600 37.200 555.900 ;
        RECT 16.800 549.600 18.600 555.600 ;
        RECT 35.400 549.600 37.200 555.600 ;
        RECT 41.400 555.600 42.300 555.900 ;
        RECT 62.400 555.600 63.600 568.950 ;
        RECT 65.100 568.050 66.900 569.850 ;
        RECT 80.100 568.050 81.900 569.850 ;
        RECT 82.950 568.950 85.050 571.050 ;
        RECT 64.950 565.950 67.050 568.050 ;
        RECT 79.950 565.950 82.050 568.050 ;
        RECT 83.400 555.600 84.600 568.950 ;
        RECT 86.100 568.050 87.900 569.850 ;
        RECT 85.950 565.950 88.050 568.050 ;
        RECT 41.400 549.600 43.200 555.600 ;
        RECT 61.800 549.600 63.600 555.600 ;
        RECT 82.800 549.600 84.600 555.600 ;
        RECT 92.550 553.050 93.450 580.950 ;
        RECT 104.700 579.600 106.500 584.400 ;
        RECT 101.400 578.400 106.500 579.600 ;
        RECT 101.400 571.050 102.600 578.400 ;
        RECT 127.200 576.000 129.000 584.400 ;
        RECT 151.800 577.200 153.600 584.400 ;
        RECT 169.800 581.400 171.600 584.400 ;
        RECT 125.700 574.800 129.000 576.000 ;
        RECT 149.400 576.300 153.600 577.200 ;
        RECT 120.000 573.450 124.200 574.050 ;
        RECT 119.550 571.950 124.200 573.450 ;
        RECT 100.950 568.950 103.050 571.050 ;
        RECT 101.400 561.600 102.600 568.950 ;
        RECT 104.100 568.050 105.900 569.850 ;
        RECT 106.950 568.950 109.050 571.050 ;
        RECT 103.950 565.950 106.050 568.050 ;
        RECT 107.100 567.150 108.900 568.950 ;
        RECT 110.100 568.050 111.900 569.850 ;
        RECT 109.950 565.950 112.050 568.050 ;
        RECT 116.100 562.950 118.200 565.050 ;
        RECT 91.950 550.950 94.050 553.050 ;
        RECT 100.800 549.600 102.600 561.600 ;
        RECT 103.800 560.700 111.600 561.600 ;
        RECT 103.800 549.600 105.600 560.700 ;
        RECT 109.800 549.600 111.600 560.700 ;
        RECT 116.550 556.050 117.450 562.950 ;
        RECT 115.800 553.950 117.900 556.050 ;
        RECT 119.550 553.050 120.450 571.950 ;
        RECT 125.700 571.050 126.600 574.800 ;
        RECT 149.400 571.050 150.600 576.300 ;
        RECT 124.950 568.950 127.050 571.050 ;
        RECT 125.700 556.800 126.600 568.950 ;
        RECT 128.100 568.050 129.900 569.850 ;
        RECT 130.950 568.950 133.050 571.050 ;
        RECT 127.950 565.950 130.050 568.050 ;
        RECT 131.100 567.150 132.900 568.950 ;
        RECT 134.100 568.050 135.900 569.850 ;
        RECT 146.100 568.050 147.900 569.850 ;
        RECT 148.950 568.950 151.050 571.050 ;
        RECT 133.950 565.950 136.050 568.050 ;
        RECT 145.950 565.950 148.050 568.050 ;
        RECT 125.700 555.900 132.300 556.800 ;
        RECT 125.700 555.600 126.600 555.900 ;
        RECT 118.950 550.950 121.050 553.050 ;
        RECT 124.800 549.600 126.600 555.600 ;
        RECT 130.800 555.600 132.300 555.900 ;
        RECT 149.400 555.600 150.600 568.950 ;
        RECT 152.100 568.050 153.900 569.850 ;
        RECT 170.400 568.050 171.600 581.400 ;
        RECT 188.400 581.400 190.200 584.400 ;
        RECT 172.950 568.950 175.050 571.050 ;
        RECT 184.950 568.950 187.050 571.050 ;
        RECT 151.950 565.950 154.050 568.050 ;
        RECT 169.950 562.950 172.050 568.050 ;
        RECT 173.100 567.150 174.900 568.950 ;
        RECT 185.100 567.150 186.900 568.950 ;
        RECT 188.400 568.050 189.600 581.400 ;
        RECT 208.200 576.000 210.000 584.400 ;
        RECT 232.200 576.000 234.000 584.400 ;
        RECT 256.800 577.200 258.600 584.400 ;
        RECT 278.700 579.600 280.500 584.400 ;
        RECT 206.700 574.800 210.000 576.000 ;
        RECT 230.700 574.800 234.000 576.000 ;
        RECT 254.400 576.300 258.600 577.200 ;
        RECT 275.400 578.400 280.500 579.600 ;
        RECT 199.950 571.950 202.050 574.050 ;
        RECT 187.950 562.950 190.050 568.050 ;
        RECT 170.400 555.600 171.600 562.950 ;
        RECT 130.800 549.600 132.600 555.600 ;
        RECT 149.400 549.600 151.200 555.600 ;
        RECT 169.800 549.600 171.600 555.600 ;
        RECT 188.400 555.600 189.600 562.950 ;
        RECT 200.550 556.050 201.450 571.950 ;
        RECT 206.700 571.050 207.600 574.800 ;
        RECT 230.700 571.050 231.600 574.800 ;
        RECT 254.400 571.050 255.600 576.300 ;
        RECT 275.400 571.050 276.600 578.400 ;
        RECT 301.200 576.000 303.000 584.400 ;
        RECT 322.800 581.400 324.600 584.400 ;
        RECT 299.700 574.800 303.000 576.000 ;
        RECT 299.700 571.050 300.600 574.800 ;
        RECT 205.950 568.950 208.050 571.050 ;
        RECT 206.700 556.800 207.600 568.950 ;
        RECT 209.100 568.050 210.900 569.850 ;
        RECT 211.950 568.950 214.050 571.050 ;
        RECT 208.950 565.950 211.050 568.050 ;
        RECT 212.100 567.150 213.900 568.950 ;
        RECT 215.100 568.050 216.900 569.850 ;
        RECT 229.950 568.950 232.050 571.050 ;
        RECT 214.950 565.950 217.050 568.050 ;
        RECT 230.700 556.800 231.600 568.950 ;
        RECT 233.100 568.050 234.900 569.850 ;
        RECT 235.950 568.950 238.050 571.050 ;
        RECT 232.950 565.950 235.050 568.050 ;
        RECT 236.100 567.150 237.900 568.950 ;
        RECT 239.100 568.050 240.900 569.850 ;
        RECT 251.100 568.050 252.900 569.850 ;
        RECT 253.950 568.950 256.050 571.050 ;
        RECT 238.950 565.950 241.050 568.050 ;
        RECT 250.950 565.950 253.050 568.050 ;
        RECT 188.400 549.600 190.200 555.600 ;
        RECT 199.950 553.950 202.050 556.050 ;
        RECT 206.700 555.900 213.300 556.800 ;
        RECT 206.700 555.600 207.600 555.900 ;
        RECT 205.800 549.600 207.600 555.600 ;
        RECT 211.800 555.600 213.300 555.900 ;
        RECT 230.700 555.900 237.300 556.800 ;
        RECT 230.700 555.600 231.600 555.900 ;
        RECT 211.800 549.600 213.600 555.600 ;
        RECT 229.800 549.600 231.600 555.600 ;
        RECT 235.800 555.600 237.300 555.900 ;
        RECT 254.400 555.600 255.600 568.950 ;
        RECT 257.100 568.050 258.900 569.850 ;
        RECT 274.950 568.950 277.050 571.050 ;
        RECT 256.950 565.950 259.050 568.050 ;
        RECT 275.400 561.600 276.600 568.950 ;
        RECT 278.100 568.050 279.900 569.850 ;
        RECT 280.950 568.950 283.050 571.050 ;
        RECT 277.950 565.950 280.050 568.050 ;
        RECT 281.100 567.150 282.900 568.950 ;
        RECT 284.100 568.050 285.900 569.850 ;
        RECT 298.950 568.950 301.050 571.050 ;
        RECT 283.950 565.950 286.050 568.050 ;
        RECT 235.800 549.600 237.600 555.600 ;
        RECT 254.400 549.600 256.200 555.600 ;
        RECT 274.800 549.600 276.600 561.600 ;
        RECT 277.800 560.700 285.600 561.600 ;
        RECT 277.800 549.600 279.600 560.700 ;
        RECT 283.800 549.600 285.600 560.700 ;
        RECT 299.700 556.800 300.600 568.950 ;
        RECT 302.100 568.050 303.900 569.850 ;
        RECT 304.950 568.950 307.050 571.050 ;
        RECT 301.950 565.950 304.050 568.050 ;
        RECT 305.100 567.150 306.900 568.950 ;
        RECT 308.100 568.050 309.900 569.850 ;
        RECT 323.400 568.050 324.600 581.400 ;
        RECT 344.700 579.600 346.500 584.400 ;
        RECT 341.400 578.400 346.500 579.600 ;
        RECT 341.400 571.050 342.600 578.400 ;
        RECT 367.200 576.000 369.000 584.400 ;
        RECT 379.950 577.950 382.050 580.050 ;
        RECT 365.700 574.800 369.000 576.000 ;
        RECT 355.950 571.950 358.050 574.050 ;
        RECT 325.950 568.950 328.050 571.050 ;
        RECT 340.950 568.950 343.050 571.050 ;
        RECT 307.950 565.950 310.050 568.050 ;
        RECT 322.950 562.950 325.050 568.050 ;
        RECT 326.100 567.150 327.900 568.950 ;
        RECT 299.700 555.900 306.300 556.800 ;
        RECT 299.700 555.600 300.600 555.900 ;
        RECT 298.800 549.600 300.600 555.600 ;
        RECT 304.800 555.600 306.300 555.900 ;
        RECT 323.400 555.600 324.600 562.950 ;
        RECT 341.400 561.600 342.600 568.950 ;
        RECT 344.100 568.050 345.900 569.850 ;
        RECT 346.950 568.950 349.050 571.050 ;
        RECT 343.950 565.950 346.050 568.050 ;
        RECT 347.100 567.150 348.900 568.950 ;
        RECT 350.100 568.050 351.900 569.850 ;
        RECT 349.950 565.950 352.050 568.050 ;
        RECT 304.800 549.600 306.600 555.600 ;
        RECT 322.800 549.600 324.600 555.600 ;
        RECT 340.800 549.600 342.600 561.600 ;
        RECT 343.800 560.700 351.600 561.600 ;
        RECT 343.800 549.600 345.600 560.700 ;
        RECT 349.800 549.600 351.600 560.700 ;
        RECT 356.550 553.050 357.450 571.950 ;
        RECT 365.700 571.050 366.600 574.800 ;
        RECT 364.950 568.950 367.050 571.050 ;
        RECT 365.700 556.800 366.600 568.950 ;
        RECT 368.100 568.050 369.900 569.850 ;
        RECT 370.950 568.950 373.050 571.050 ;
        RECT 367.950 565.950 370.050 568.050 ;
        RECT 371.100 567.150 372.900 568.950 ;
        RECT 374.100 568.050 375.900 569.850 ;
        RECT 373.950 565.950 376.050 568.050 ;
        RECT 380.550 559.050 381.450 577.950 ;
        RECT 389.400 577.200 391.200 584.400 ;
        RECT 412.800 577.200 414.600 584.400 ;
        RECT 430.800 578.400 432.600 584.400 ;
        RECT 389.400 576.300 393.600 577.200 ;
        RECT 392.400 571.050 393.600 576.300 ;
        RECT 410.400 576.300 414.600 577.200 ;
        RECT 431.400 576.300 432.600 578.400 ;
        RECT 433.800 579.300 435.600 584.400 ;
        RECT 439.800 579.300 441.600 584.400 ;
        RECT 433.800 577.950 441.600 579.300 ;
        RECT 455.400 577.200 457.200 584.400 ;
        RECT 475.800 578.400 477.600 584.400 ;
        RECT 455.400 576.300 459.600 577.200 ;
        RECT 400.950 571.950 403.050 574.050 ;
        RECT 389.100 568.050 390.900 569.850 ;
        RECT 391.950 568.950 394.050 571.050 ;
        RECT 388.950 565.950 391.050 568.050 ;
        RECT 379.950 556.950 382.050 559.050 ;
        RECT 365.700 555.900 372.300 556.800 ;
        RECT 365.700 555.600 366.600 555.900 ;
        RECT 355.950 550.950 358.050 553.050 ;
        RECT 364.800 549.600 366.600 555.600 ;
        RECT 370.800 555.600 372.300 555.900 ;
        RECT 392.400 555.600 393.600 568.950 ;
        RECT 395.100 568.050 396.900 569.850 ;
        RECT 394.950 565.950 397.050 568.050 ;
        RECT 401.550 556.050 402.450 571.950 ;
        RECT 410.400 571.050 411.600 576.300 ;
        RECT 431.400 575.250 435.150 576.300 ;
        RECT 433.950 571.050 435.150 575.250 ;
        RECT 458.400 571.050 459.600 576.300 ;
        RECT 476.400 576.300 477.600 578.400 ;
        RECT 478.800 579.300 480.600 584.400 ;
        RECT 484.800 579.300 486.600 584.400 ;
        RECT 478.800 577.950 486.600 579.300 ;
        RECT 497.400 579.300 499.200 584.400 ;
        RECT 503.400 579.300 505.200 584.400 ;
        RECT 497.400 577.950 505.200 579.300 ;
        RECT 506.400 578.400 508.200 584.400 ;
        RECT 527.700 579.600 529.500 584.400 ;
        RECT 524.400 578.400 529.500 579.600 ;
        RECT 506.400 576.300 507.600 578.400 ;
        RECT 476.400 575.250 480.150 576.300 ;
        RECT 478.950 571.050 480.150 575.250 ;
        RECT 503.850 575.250 507.600 576.300 ;
        RECT 503.850 571.050 505.050 575.250 ;
        RECT 511.800 571.950 513.900 574.050 ;
        RECT 407.100 568.050 408.900 569.850 ;
        RECT 409.950 568.950 412.050 571.050 ;
        RECT 406.950 565.950 409.050 568.050 ;
        RECT 370.800 549.600 372.600 555.600 ;
        RECT 391.800 549.600 393.600 555.600 ;
        RECT 400.950 553.950 403.050 556.050 ;
        RECT 410.400 555.600 411.600 568.950 ;
        RECT 413.100 568.050 414.900 569.850 ;
        RECT 431.100 568.050 432.900 569.850 ;
        RECT 433.950 568.950 436.050 571.050 ;
        RECT 412.950 565.950 415.050 568.050 ;
        RECT 430.950 565.950 433.050 568.050 ;
        RECT 434.850 555.600 436.050 568.950 ;
        RECT 437.100 568.050 438.900 569.850 ;
        RECT 439.950 568.950 442.050 571.050 ;
        RECT 436.950 565.950 439.050 568.050 ;
        RECT 440.100 567.150 441.900 568.950 ;
        RECT 455.100 568.050 456.900 569.850 ;
        RECT 457.950 568.950 460.050 571.050 ;
        RECT 454.950 565.950 457.050 568.050 ;
        RECT 458.400 555.600 459.600 568.950 ;
        RECT 461.100 568.050 462.900 569.850 ;
        RECT 476.100 568.050 477.900 569.850 ;
        RECT 478.950 568.950 481.050 571.050 ;
        RECT 460.950 565.950 463.050 568.050 ;
        RECT 475.950 565.950 478.050 568.050 ;
        RECT 466.950 562.950 469.050 565.050 ;
        RECT 410.400 549.600 412.200 555.600 ;
        RECT 434.400 549.600 436.200 555.600 ;
        RECT 457.800 549.600 459.600 555.600 ;
        RECT 467.550 553.050 468.450 562.950 ;
        RECT 479.850 555.600 481.050 568.950 ;
        RECT 482.100 568.050 483.900 569.850 ;
        RECT 484.950 568.950 487.050 571.050 ;
        RECT 496.950 568.950 499.050 571.050 ;
        RECT 481.950 565.950 484.050 568.050 ;
        RECT 485.100 567.150 486.900 568.950 ;
        RECT 497.100 567.150 498.900 568.950 ;
        RECT 500.100 568.050 501.900 569.850 ;
        RECT 502.950 568.950 505.050 571.050 ;
        RECT 499.950 565.950 502.050 568.050 ;
        RECT 502.950 555.600 504.150 568.950 ;
        RECT 506.100 568.050 507.900 569.850 ;
        RECT 505.950 565.950 508.050 568.050 ;
        RECT 467.100 550.950 469.200 553.050 ;
        RECT 479.400 549.600 481.200 555.600 ;
        RECT 502.800 549.600 504.600 555.600 ;
        RECT 512.550 553.050 513.450 571.950 ;
        RECT 524.400 571.050 525.600 578.400 ;
        RECT 550.200 576.000 552.000 584.400 ;
        RECT 571.800 581.400 573.600 584.400 ;
        RECT 562.950 577.950 565.050 580.050 ;
        RECT 548.700 574.800 552.000 576.000 ;
        RECT 548.700 571.050 549.600 574.800 ;
        RECT 523.950 568.950 526.050 571.050 ;
        RECT 524.400 561.600 525.600 568.950 ;
        RECT 527.100 568.050 528.900 569.850 ;
        RECT 529.950 568.950 532.050 571.050 ;
        RECT 526.950 565.950 529.050 568.050 ;
        RECT 530.100 567.150 531.900 568.950 ;
        RECT 533.100 568.050 534.900 569.850 ;
        RECT 547.950 568.950 550.050 571.050 ;
        RECT 532.950 565.950 535.050 568.050 ;
        RECT 511.950 550.950 514.050 553.050 ;
        RECT 523.800 549.600 525.600 561.600 ;
        RECT 526.800 560.700 534.600 561.600 ;
        RECT 526.800 549.600 528.600 560.700 ;
        RECT 532.800 549.600 534.600 560.700 ;
        RECT 548.700 556.800 549.600 568.950 ;
        RECT 551.100 568.050 552.900 569.850 ;
        RECT 553.950 568.950 556.050 571.050 ;
        RECT 550.950 565.950 553.050 568.050 ;
        RECT 554.100 567.150 555.900 568.950 ;
        RECT 557.100 568.050 558.900 569.850 ;
        RECT 556.950 565.950 559.050 568.050 ;
        RECT 563.550 559.050 564.450 577.950 ;
        RECT 572.400 568.050 573.600 581.400 ;
        RECT 592.500 579.600 594.300 584.400 ;
        RECT 615.300 580.200 617.100 584.400 ;
        RECT 592.500 578.400 597.600 579.600 ;
        RECT 580.950 571.950 583.050 574.050 ;
        RECT 574.950 568.950 577.050 571.050 ;
        RECT 571.950 562.950 574.050 568.050 ;
        RECT 575.100 567.150 576.900 568.950 ;
        RECT 577.950 562.950 580.050 565.050 ;
        RECT 562.950 556.950 565.050 559.050 ;
        RECT 548.700 555.900 555.300 556.800 ;
        RECT 548.700 555.600 549.600 555.900 ;
        RECT 547.800 549.600 549.600 555.600 ;
        RECT 553.800 555.600 555.300 555.900 ;
        RECT 572.400 555.600 573.600 562.950 ;
        RECT 553.800 549.600 555.600 555.600 ;
        RECT 571.800 549.600 573.600 555.600 ;
        RECT 578.550 553.050 579.450 562.950 ;
        RECT 581.550 562.050 582.450 571.950 ;
        RECT 596.400 571.050 597.600 578.400 ;
        RECT 614.400 578.400 617.100 580.200 ;
        RECT 614.400 571.050 615.300 578.400 ;
        RECT 617.100 576.600 618.900 577.500 ;
        RECT 622.800 576.600 624.600 584.400 ;
        RECT 625.950 580.950 628.050 583.050 ;
        RECT 626.550 577.050 627.450 580.950 ;
        RECT 640.800 577.200 642.600 584.400 ;
        RECT 658.800 578.400 660.600 584.400 ;
        RECT 617.100 575.700 624.600 576.600 ;
        RECT 587.100 568.050 588.900 569.850 ;
        RECT 589.950 568.950 592.050 571.050 ;
        RECT 586.950 565.950 589.050 568.050 ;
        RECT 590.100 567.150 591.900 568.950 ;
        RECT 593.100 568.050 594.900 569.850 ;
        RECT 595.950 568.950 598.050 571.050 ;
        RECT 613.950 568.950 616.050 571.050 ;
        RECT 616.950 568.950 619.050 571.050 ;
        RECT 592.950 565.950 595.050 568.050 ;
        RECT 580.950 559.950 583.050 562.050 ;
        RECT 596.400 561.600 597.600 568.950 ;
        RECT 614.400 561.600 615.300 568.950 ;
        RECT 617.100 567.150 618.900 568.950 ;
        RECT 587.400 560.700 595.200 561.600 ;
        RECT 578.100 550.950 580.200 553.050 ;
        RECT 587.400 549.600 589.200 560.700 ;
        RECT 593.400 549.600 595.200 560.700 ;
        RECT 596.400 549.600 598.200 561.600 ;
        RECT 613.500 549.600 615.300 561.600 ;
        RECT 620.700 555.600 621.600 575.700 ;
        RECT 625.950 574.950 628.050 577.050 ;
        RECT 638.400 576.300 642.600 577.200 ;
        RECT 659.400 576.300 660.600 578.400 ;
        RECT 661.800 579.300 663.600 584.400 ;
        RECT 667.800 579.300 669.600 584.400 ;
        RECT 661.800 577.950 669.600 579.300 ;
        RECT 623.100 571.050 624.900 572.850 ;
        RECT 638.400 571.050 639.600 576.300 ;
        RECT 659.400 575.250 663.150 576.300 ;
        RECT 685.200 576.000 687.000 584.400 ;
        RECT 710.700 579.600 712.500 584.400 ;
        RECT 721.800 580.950 723.900 583.050 ;
        RECT 725.100 580.950 727.200 583.050 ;
        RECT 661.950 571.050 663.150 575.250 ;
        RECT 683.700 574.800 687.000 576.000 ;
        RECT 707.400 578.400 712.500 579.600 ;
        RECT 683.700 571.050 684.600 574.800 ;
        RECT 707.400 571.050 708.600 578.400 ;
        RECT 622.950 568.950 625.050 571.050 ;
        RECT 635.100 568.050 636.900 569.850 ;
        RECT 637.950 568.950 640.050 571.050 ;
        RECT 634.950 565.950 637.050 568.050 ;
        RECT 619.800 549.600 621.600 555.600 ;
        RECT 638.400 555.600 639.600 568.950 ;
        RECT 641.100 568.050 642.900 569.850 ;
        RECT 659.100 568.050 660.900 569.850 ;
        RECT 661.950 568.950 664.050 571.050 ;
        RECT 640.950 565.950 643.050 568.050 ;
        RECT 658.950 565.950 661.050 568.050 ;
        RECT 662.850 555.600 664.050 568.950 ;
        RECT 665.100 568.050 666.900 569.850 ;
        RECT 667.950 568.950 670.050 571.050 ;
        RECT 682.950 568.950 685.050 571.050 ;
        RECT 664.950 565.950 667.050 568.050 ;
        RECT 668.100 567.150 669.900 568.950 ;
        RECT 683.700 556.800 684.600 568.950 ;
        RECT 686.100 568.050 687.900 569.850 ;
        RECT 688.950 568.950 691.050 571.050 ;
        RECT 685.950 565.950 688.050 568.050 ;
        RECT 689.100 567.150 690.900 568.950 ;
        RECT 692.100 568.050 693.900 569.850 ;
        RECT 706.950 568.950 709.050 571.050 ;
        RECT 691.950 565.950 694.050 568.050 ;
        RECT 707.400 561.600 708.600 568.950 ;
        RECT 710.100 568.050 711.900 569.850 ;
        RECT 712.950 568.950 715.050 571.050 ;
        RECT 709.950 565.950 712.050 568.050 ;
        RECT 713.100 567.150 714.900 568.950 ;
        RECT 716.100 568.050 717.900 569.850 ;
        RECT 715.950 565.950 718.050 568.050 ;
        RECT 683.700 555.900 690.300 556.800 ;
        RECT 683.700 555.600 684.600 555.900 ;
        RECT 638.400 549.600 640.200 555.600 ;
        RECT 662.400 549.600 664.200 555.600 ;
        RECT 682.800 549.600 684.600 555.600 ;
        RECT 688.800 555.600 690.300 555.900 ;
        RECT 688.800 549.600 690.600 555.600 ;
        RECT 706.800 549.600 708.600 561.600 ;
        RECT 709.800 560.700 717.600 561.600 ;
        RECT 709.800 549.600 711.600 560.700 ;
        RECT 715.800 549.600 717.600 560.700 ;
        RECT 722.550 559.050 723.450 580.950 ;
        RECT 725.550 577.050 726.450 580.950 ;
        RECT 724.950 574.950 727.050 577.050 ;
        RECT 735.000 576.000 736.800 584.400 ;
        RECT 755.400 581.400 757.200 584.400 ;
        RECT 776.400 581.400 778.200 584.400 ;
        RECT 735.000 574.800 738.300 576.000 ;
        RECT 737.400 571.050 738.300 574.800 ;
        RECT 751.950 571.950 754.050 574.050 ;
        RECT 728.100 568.050 729.900 569.850 ;
        RECT 730.950 568.950 733.050 571.050 ;
        RECT 727.950 565.950 730.050 568.050 ;
        RECT 731.100 567.150 732.900 568.950 ;
        RECT 734.100 568.050 735.900 569.850 ;
        RECT 736.950 568.950 739.050 571.050 ;
        RECT 752.100 570.150 753.900 571.950 ;
        RECT 755.700 571.050 756.600 581.400 ;
        RECT 757.950 571.950 760.050 574.050 ;
        RECT 754.950 568.950 757.050 571.050 ;
        RECT 758.100 570.150 759.900 571.950 ;
        RECT 772.950 568.950 775.050 571.050 ;
        RECT 733.950 565.950 736.050 568.050 ;
        RECT 721.950 556.950 724.050 559.050 ;
        RECT 737.400 556.800 738.300 568.950 ;
        RECT 755.700 561.600 756.600 568.950 ;
        RECT 773.100 567.150 774.900 568.950 ;
        RECT 776.400 568.050 777.600 581.400 ;
        RECT 782.100 577.950 784.200 580.050 ;
        RECT 775.950 562.950 778.050 568.050 ;
        RECT 755.700 560.400 759.300 561.600 ;
        RECT 731.700 555.900 738.300 556.800 ;
        RECT 731.700 555.600 733.200 555.900 ;
        RECT 731.400 549.600 733.200 555.600 ;
        RECT 737.400 555.600 738.300 555.900 ;
        RECT 737.400 549.600 739.200 555.600 ;
        RECT 757.500 549.600 759.300 560.400 ;
        RECT 776.400 555.600 777.600 562.950 ;
        RECT 776.400 549.600 778.200 555.600 ;
        RECT 782.550 553.050 783.450 577.950 ;
        RECT 796.200 576.000 798.000 584.400 ;
        RECT 794.700 574.800 798.000 576.000 ;
        RECT 822.000 576.000 823.800 584.400 ;
        RECT 841.800 581.400 843.600 584.400 ;
        RECT 822.000 574.800 825.300 576.000 ;
        RECT 794.700 571.050 795.600 574.800 ;
        RECT 824.400 571.050 825.300 574.800 ;
        RECT 793.950 568.950 796.050 571.050 ;
        RECT 794.700 556.800 795.600 568.950 ;
        RECT 797.100 568.050 798.900 569.850 ;
        RECT 799.950 568.950 802.050 571.050 ;
        RECT 796.950 565.950 799.050 568.050 ;
        RECT 800.100 567.150 801.900 568.950 ;
        RECT 803.100 568.050 804.900 569.850 ;
        RECT 815.100 568.050 816.900 569.850 ;
        RECT 817.950 568.950 820.050 571.050 ;
        RECT 802.950 565.950 805.050 568.050 ;
        RECT 814.950 565.950 817.050 568.050 ;
        RECT 818.100 567.150 819.900 568.950 ;
        RECT 821.100 568.050 822.900 569.850 ;
        RECT 823.950 568.950 826.050 571.050 ;
        RECT 820.950 565.950 823.050 568.050 ;
        RECT 824.400 556.800 825.300 568.950 ;
        RECT 842.400 568.050 843.600 581.400 ;
        RECT 859.800 578.400 861.600 584.400 ;
        RECT 860.400 576.300 861.600 578.400 ;
        RECT 862.800 579.300 864.600 584.400 ;
        RECT 868.800 579.300 870.600 584.400 ;
        RECT 862.800 577.950 870.600 579.300 ;
        RECT 884.400 581.400 886.200 584.400 ;
        RECT 899.400 581.400 901.200 584.400 ;
        RECT 860.400 575.250 864.150 576.300 ;
        RECT 862.950 571.050 864.150 575.250 ;
        RECT 844.950 568.950 847.050 571.050 ;
        RECT 841.950 562.950 844.050 568.050 ;
        RECT 845.100 567.150 846.900 568.950 ;
        RECT 860.100 568.050 861.900 569.850 ;
        RECT 862.950 568.950 865.050 571.050 ;
        RECT 859.950 565.950 862.050 568.050 ;
        RECT 794.700 555.900 801.300 556.800 ;
        RECT 794.700 555.600 795.600 555.900 ;
        RECT 781.950 550.950 784.050 553.050 ;
        RECT 793.800 549.600 795.600 555.600 ;
        RECT 799.800 555.600 801.300 555.900 ;
        RECT 818.700 555.900 825.300 556.800 ;
        RECT 818.700 555.600 820.200 555.900 ;
        RECT 799.800 549.600 801.600 555.600 ;
        RECT 818.400 549.600 820.200 555.600 ;
        RECT 824.400 555.600 825.300 555.900 ;
        RECT 842.400 555.600 843.600 562.950 ;
        RECT 863.850 555.600 865.050 568.950 ;
        RECT 866.100 568.050 867.900 569.850 ;
        RECT 868.950 568.950 871.050 571.050 ;
        RECT 880.950 568.950 883.050 571.050 ;
        RECT 865.950 565.950 868.050 568.050 ;
        RECT 869.100 567.150 870.900 568.950 ;
        RECT 881.100 567.150 882.900 568.950 ;
        RECT 884.400 568.050 885.600 581.400 ;
        RECT 899.400 577.500 900.600 581.400 ;
        RECT 905.700 578.400 907.500 584.400 ;
        RECT 899.400 576.600 905.400 577.500 ;
        RECT 903.150 575.700 905.400 576.600 ;
        RECT 898.950 568.950 901.050 571.050 ;
        RECT 883.950 562.950 886.050 568.050 ;
        RECT 899.100 567.150 900.900 568.950 ;
        RECT 903.150 564.300 904.050 575.700 ;
        RECT 906.300 571.050 907.500 578.400 ;
        RECT 904.950 568.950 907.500 571.050 ;
        RECT 903.150 563.400 905.400 564.300 ;
        RECT 884.400 555.600 885.600 562.950 ;
        RECT 899.400 562.500 905.400 563.400 ;
        RECT 899.400 555.600 900.600 562.500 ;
        RECT 906.300 561.600 907.500 568.950 ;
        RECT 824.400 549.600 826.200 555.600 ;
        RECT 841.800 549.600 843.600 555.600 ;
        RECT 863.400 549.600 865.200 555.600 ;
        RECT 884.400 549.600 886.200 555.600 ;
        RECT 899.400 549.600 901.200 555.600 ;
        RECT 905.700 549.600 907.500 561.600 ;
        RECT 13.800 539.400 15.600 545.400 ;
        RECT 14.400 532.050 15.600 539.400 ;
        RECT 29.400 534.300 31.200 545.400 ;
        RECT 35.400 534.300 37.200 545.400 ;
        RECT 29.400 533.400 37.200 534.300 ;
        RECT 38.400 533.400 40.200 545.400 ;
        RECT 43.950 538.950 46.050 541.050 ;
        RECT 55.800 539.400 57.600 545.400 ;
        RECT 74.400 539.400 76.200 545.400 ;
        RECT 13.950 526.950 16.050 532.050 ;
        RECT 14.400 513.600 15.600 526.950 ;
        RECT 17.100 526.050 18.900 527.850 ;
        RECT 28.950 526.950 31.050 529.050 ;
        RECT 16.950 523.950 19.050 526.050 ;
        RECT 29.100 525.150 30.900 526.950 ;
        RECT 32.100 526.050 33.900 527.850 ;
        RECT 34.950 526.950 37.050 529.050 ;
        RECT 31.950 523.950 34.050 526.050 ;
        RECT 35.100 525.150 36.900 526.950 ;
        RECT 38.400 526.050 39.600 533.400 ;
        RECT 37.950 523.950 40.050 526.050 ;
        RECT 38.400 516.600 39.600 523.950 ;
        RECT 13.800 510.600 15.600 513.600 ;
        RECT 34.500 515.400 39.600 516.600 ;
        RECT 34.500 510.600 36.300 515.400 ;
        RECT 44.550 514.050 45.450 538.950 ;
        RECT 56.400 532.050 57.600 539.400 ;
        RECT 74.700 539.100 76.200 539.400 ;
        RECT 80.400 539.400 82.200 545.400 ;
        RECT 100.800 539.400 102.600 545.400 ;
        RECT 119.400 539.400 121.200 545.400 ;
        RECT 80.400 539.100 81.300 539.400 ;
        RECT 74.700 538.200 81.300 539.100 ;
        RECT 55.950 526.950 58.050 532.050 ;
        RECT 43.950 511.950 46.050 514.050 ;
        RECT 56.400 513.600 57.600 526.950 ;
        RECT 59.100 526.050 60.900 527.850 ;
        RECT 70.950 526.950 73.050 529.050 ;
        RECT 58.950 523.950 61.050 526.050 ;
        RECT 71.100 525.150 72.900 526.950 ;
        RECT 74.100 526.050 75.900 527.850 ;
        RECT 76.950 526.950 79.050 529.050 ;
        RECT 73.950 523.950 76.050 526.050 ;
        RECT 77.100 525.150 78.900 526.950 ;
        RECT 80.400 526.050 81.300 538.200 ;
        RECT 85.950 535.950 88.050 538.050 ;
        RECT 79.950 523.950 82.050 526.050 ;
        RECT 80.400 520.200 81.300 523.950 ;
        RECT 86.550 523.050 87.450 535.950 ;
        RECT 95.100 526.050 96.900 527.850 ;
        RECT 97.950 526.950 100.050 529.050 ;
        RECT 94.950 523.950 97.050 526.050 ;
        RECT 98.100 525.150 99.900 526.950 ;
        RECT 100.950 526.050 102.150 539.400 ;
        RECT 119.400 532.500 120.600 539.400 ;
        RECT 125.700 533.400 127.500 545.400 ;
        RECT 119.400 531.600 125.400 532.500 ;
        RECT 123.150 530.700 125.400 531.600 ;
        RECT 103.950 526.950 106.050 529.050 ;
        RECT 100.950 523.950 103.050 526.050 ;
        RECT 104.100 525.150 105.900 526.950 ;
        RECT 119.100 526.050 120.900 527.850 ;
        RECT 118.950 523.950 121.050 526.050 ;
        RECT 85.950 520.950 88.050 523.050 ;
        RECT 55.800 510.600 57.600 513.600 ;
        RECT 78.000 519.000 81.300 520.200 ;
        RECT 78.000 510.600 79.800 519.000 ;
        RECT 86.550 517.050 87.450 520.950 ;
        RECT 101.850 519.750 103.050 523.950 ;
        RECT 101.850 518.700 105.600 519.750 ;
        RECT 85.950 514.950 88.050 517.050 ;
        RECT 95.400 515.700 103.200 517.050 ;
        RECT 95.400 510.600 97.200 515.700 ;
        RECT 101.400 510.600 103.200 515.700 ;
        RECT 104.400 516.600 105.600 518.700 ;
        RECT 123.150 519.300 124.050 530.700 ;
        RECT 126.300 526.050 127.500 533.400 ;
        RECT 124.950 523.950 127.500 526.050 ;
        RECT 123.150 518.400 125.400 519.300 ;
        RECT 119.400 517.500 125.400 518.400 ;
        RECT 104.400 510.600 106.200 516.600 ;
        RECT 119.400 513.600 120.600 517.500 ;
        RECT 126.300 516.600 127.500 523.950 ;
        RECT 119.400 510.600 121.200 513.600 ;
        RECT 125.700 510.600 127.500 516.600 ;
        RECT 132.150 533.400 133.950 545.400 ;
        RECT 140.550 539.400 142.350 545.400 ;
        RECT 140.550 538.500 141.750 539.400 ;
        RECT 148.350 538.500 150.150 545.400 ;
        RECT 156.150 539.400 157.950 545.400 ;
        RECT 136.950 536.400 141.750 538.500 ;
        RECT 144.450 537.450 151.050 538.500 ;
        RECT 144.450 536.700 146.250 537.450 ;
        RECT 149.250 536.700 151.050 537.450 ;
        RECT 156.150 537.300 160.050 539.400 ;
        RECT 140.550 535.500 141.750 536.400 ;
        RECT 153.450 535.800 155.250 536.400 ;
        RECT 140.550 534.300 148.050 535.500 ;
        RECT 146.250 533.700 148.050 534.300 ;
        RECT 148.950 534.900 155.250 535.800 ;
        RECT 132.150 532.500 133.050 533.400 ;
        RECT 148.950 532.800 149.850 534.900 ;
        RECT 153.450 534.600 155.250 534.900 ;
        RECT 156.150 534.600 158.850 536.400 ;
        RECT 156.150 533.700 157.050 534.600 ;
        RECT 141.450 532.500 149.850 532.800 ;
        RECT 132.150 531.900 149.850 532.500 ;
        RECT 151.950 532.800 157.050 533.700 ;
        RECT 157.950 532.800 160.050 533.700 ;
        RECT 163.650 533.400 165.450 545.400 ;
        RECT 181.800 539.400 183.600 545.400 ;
        RECT 205.800 539.400 207.600 545.400 ;
        RECT 227.400 539.400 229.200 545.400 ;
        RECT 251.400 539.400 253.200 545.400 ;
        RECT 132.150 531.300 143.250 531.900 ;
        RECT 132.150 516.600 133.050 531.300 ;
        RECT 141.450 531.000 143.250 531.300 ;
        RECT 133.950 523.950 136.050 526.050 ;
        RECT 142.950 524.400 145.050 526.050 ;
        RECT 134.100 522.150 135.900 523.950 ;
        RECT 137.100 523.200 145.050 524.400 ;
        RECT 137.100 522.600 138.900 523.200 ;
        RECT 135.000 521.400 135.900 522.150 ;
        RECT 140.100 521.400 141.900 522.000 ;
        RECT 135.000 520.200 141.900 521.400 ;
        RECT 151.950 520.200 152.850 532.800 ;
        RECT 157.950 531.600 162.150 532.800 ;
        RECT 161.250 529.800 163.050 531.600 ;
        RECT 164.250 526.050 165.450 533.400 ;
        RECT 176.100 526.050 177.900 527.850 ;
        RECT 178.950 526.950 181.050 529.050 ;
        RECT 160.950 525.750 165.450 526.050 ;
        RECT 159.150 523.950 165.450 525.750 ;
        RECT 175.950 523.950 178.050 526.050 ;
        RECT 179.100 525.150 180.900 526.950 ;
        RECT 181.950 526.050 183.150 539.400 ;
        RECT 184.950 526.950 187.050 529.050 ;
        RECT 202.950 526.950 205.050 529.050 ;
        RECT 181.950 523.950 184.050 526.050 ;
        RECT 185.100 525.150 186.900 526.950 ;
        RECT 203.100 525.150 204.900 526.950 ;
        RECT 206.400 526.050 207.600 539.400 ;
        RECT 208.950 526.950 211.050 529.050 ;
        RECT 223.950 526.950 226.050 529.050 ;
        RECT 205.950 523.950 208.050 526.050 ;
        RECT 209.100 525.150 210.900 526.950 ;
        RECT 224.100 525.150 225.900 526.950 ;
        RECT 227.850 526.050 229.050 539.400 ;
        RECT 229.950 526.950 232.050 529.050 ;
        RECT 226.950 523.950 229.050 526.050 ;
        RECT 230.100 525.150 231.900 526.950 ;
        RECT 233.100 526.050 234.900 527.850 ;
        RECT 247.950 526.950 250.050 529.050 ;
        RECT 232.950 523.950 235.050 526.050 ;
        RECT 248.100 525.150 249.900 526.950 ;
        RECT 251.850 526.050 253.050 539.400 ;
        RECT 271.800 533.400 273.600 545.400 ;
        RECT 274.800 534.300 276.600 545.400 ;
        RECT 280.800 534.300 282.600 545.400 ;
        RECT 295.800 539.400 297.600 545.400 ;
        RECT 274.800 533.400 282.600 534.300 ;
        RECT 296.700 539.100 297.600 539.400 ;
        RECT 301.800 539.400 303.600 545.400 ;
        RECT 320.400 539.400 322.200 545.400 ;
        RECT 301.800 539.100 303.300 539.400 ;
        RECT 296.700 538.200 303.300 539.100 ;
        RECT 320.700 539.100 322.200 539.400 ;
        RECT 326.400 539.400 328.200 545.400 ;
        RECT 346.800 539.400 348.600 545.400 ;
        RECT 326.400 539.100 327.300 539.400 ;
        RECT 320.700 538.200 327.300 539.100 ;
        RECT 253.950 526.950 256.050 529.050 ;
        RECT 250.950 523.950 253.050 526.050 ;
        RECT 254.100 525.150 255.900 526.950 ;
        RECT 257.100 526.050 258.900 527.850 ;
        RECT 272.400 526.050 273.600 533.400 ;
        RECT 274.950 526.950 277.050 529.050 ;
        RECT 256.950 523.950 259.050 526.050 ;
        RECT 271.950 523.950 274.050 526.050 ;
        RECT 275.100 525.150 276.900 526.950 ;
        RECT 278.100 526.050 279.900 527.850 ;
        RECT 280.950 526.950 283.050 529.050 ;
        RECT 277.950 523.950 280.050 526.050 ;
        RECT 281.100 525.150 282.900 526.950 ;
        RECT 296.700 526.050 297.600 538.200 ;
        RECT 298.950 526.950 301.050 529.050 ;
        RECT 295.950 523.950 298.050 526.050 ;
        RECT 299.100 525.150 300.900 526.950 ;
        RECT 302.100 526.050 303.900 527.850 ;
        RECT 304.950 526.950 307.050 529.050 ;
        RECT 316.950 526.950 319.050 529.050 ;
        RECT 301.950 523.950 304.050 526.050 ;
        RECT 305.100 525.150 306.900 526.950 ;
        RECT 317.100 525.150 318.900 526.950 ;
        RECT 320.100 526.050 321.900 527.850 ;
        RECT 322.950 526.950 325.050 529.050 ;
        RECT 319.950 523.950 322.050 526.050 ;
        RECT 323.100 525.150 324.900 526.950 ;
        RECT 326.400 526.050 327.300 538.200 ;
        RECT 341.100 526.050 342.900 527.850 ;
        RECT 343.950 526.950 346.050 529.050 ;
        RECT 325.950 523.950 328.050 526.050 ;
        RECT 340.950 523.950 343.050 526.050 ;
        RECT 344.100 525.150 345.900 526.950 ;
        RECT 346.950 526.050 348.150 539.400 ;
        RECT 365.400 534.600 367.200 545.400 ;
        RECT 371.400 544.500 379.200 545.400 ;
        RECT 371.400 534.600 373.200 544.500 ;
        RECT 365.400 533.700 373.200 534.600 ;
        RECT 374.400 532.500 376.200 543.600 ;
        RECT 377.400 533.400 379.200 544.500 ;
        RECT 394.500 533.400 396.300 545.400 ;
        RECT 400.800 539.400 402.600 545.400 ;
        RECT 415.800 539.400 417.600 545.400 ;
        RECT 371.100 531.600 376.200 532.500 ;
        RECT 349.950 526.950 352.050 529.050 ;
        RECT 346.950 523.950 349.050 526.050 ;
        RECT 350.100 525.150 351.900 526.950 ;
        RECT 371.100 526.050 372.000 531.600 ;
        RECT 394.500 526.050 395.700 533.400 ;
        RECT 401.400 532.500 402.600 539.400 ;
        RECT 396.600 531.600 402.600 532.500 ;
        RECT 416.700 539.100 417.600 539.400 ;
        RECT 421.800 539.400 423.600 545.400 ;
        RECT 439.800 539.400 441.600 545.400 ;
        RECT 421.800 539.100 423.300 539.400 ;
        RECT 416.700 538.200 423.300 539.100 ;
        RECT 440.700 539.100 441.600 539.400 ;
        RECT 445.800 539.400 447.600 545.400 ;
        RECT 457.950 541.950 460.050 544.050 ;
        RECT 445.800 539.100 447.300 539.400 ;
        RECT 440.700 538.200 447.300 539.100 ;
        RECT 396.600 530.700 398.850 531.600 ;
        RECT 364.950 523.950 367.050 526.050 ;
        RECT 140.850 519.000 152.850 520.200 ;
        RECT 140.850 517.200 141.900 519.000 ;
        RECT 151.050 518.400 152.850 519.000 ;
        RECT 132.150 510.600 133.950 516.600 ;
        RECT 136.950 514.500 139.050 516.600 ;
        RECT 140.550 515.400 142.350 517.200 ;
        RECT 164.250 516.600 165.450 523.950 ;
        RECT 182.850 519.750 184.050 523.950 ;
        RECT 182.850 518.700 186.600 519.750 ;
        RECT 206.400 518.700 207.600 523.950 ;
        RECT 226.950 519.750 228.150 523.950 ;
        RECT 250.950 519.750 252.150 523.950 ;
        RECT 143.850 515.550 145.650 516.300 ;
        RECT 157.950 515.700 160.050 516.600 ;
        RECT 143.850 514.500 148.800 515.550 ;
        RECT 138.000 513.600 139.050 514.500 ;
        RECT 147.750 513.600 148.800 514.500 ;
        RECT 156.300 514.500 160.050 515.700 ;
        RECT 156.300 513.600 157.350 514.500 ;
        RECT 138.000 512.700 141.750 513.600 ;
        RECT 139.950 510.600 141.750 512.700 ;
        RECT 147.750 510.600 149.550 513.600 ;
        RECT 155.550 510.600 157.350 513.600 ;
        RECT 163.650 510.600 165.450 516.600 ;
        RECT 176.400 515.700 184.200 517.050 ;
        RECT 176.400 510.600 178.200 515.700 ;
        RECT 182.400 510.600 184.200 515.700 ;
        RECT 185.400 516.600 186.600 518.700 ;
        RECT 203.400 517.800 207.600 518.700 ;
        RECT 224.400 518.700 228.150 519.750 ;
        RECT 248.400 518.700 252.150 519.750 ;
        RECT 185.400 510.600 187.200 516.600 ;
        RECT 203.400 510.600 205.200 517.800 ;
        RECT 224.400 516.600 225.600 518.700 ;
        RECT 223.800 510.600 225.600 516.600 ;
        RECT 226.800 515.700 234.600 517.050 ;
        RECT 248.400 516.600 249.600 518.700 ;
        RECT 226.800 510.600 228.600 515.700 ;
        RECT 232.800 510.600 234.600 515.700 ;
        RECT 247.800 510.600 249.600 516.600 ;
        RECT 250.800 515.700 258.600 517.050 ;
        RECT 250.800 510.600 252.600 515.700 ;
        RECT 256.800 510.600 258.600 515.700 ;
        RECT 272.400 516.600 273.600 523.950 ;
        RECT 296.700 520.200 297.600 523.950 ;
        RECT 326.400 520.200 327.300 523.950 ;
        RECT 296.700 519.000 300.000 520.200 ;
        RECT 272.400 515.400 277.500 516.600 ;
        RECT 275.700 510.600 277.500 515.400 ;
        RECT 298.200 510.600 300.000 519.000 ;
        RECT 324.000 519.000 327.300 520.200 ;
        RECT 347.850 519.750 349.050 523.950 ;
        RECT 361.950 520.950 364.050 523.050 ;
        RECT 365.100 522.150 366.900 523.950 ;
        RECT 368.100 523.050 369.900 524.850 ;
        RECT 370.950 523.950 373.050 526.050 ;
        RECT 367.950 520.950 370.050 523.050 ;
        RECT 324.000 510.600 325.800 519.000 ;
        RECT 347.850 518.700 351.600 519.750 ;
        RECT 341.400 515.700 349.200 517.050 ;
        RECT 341.400 510.600 343.200 515.700 ;
        RECT 347.400 510.600 349.200 515.700 ;
        RECT 350.400 516.600 351.600 518.700 ;
        RECT 350.400 510.600 352.200 516.600 ;
        RECT 362.550 514.050 363.450 520.950 ;
        RECT 370.950 516.600 372.000 523.950 ;
        RECT 374.100 523.050 375.900 524.850 ;
        RECT 376.950 523.950 379.050 526.050 ;
        RECT 394.500 523.950 397.050 526.050 ;
        RECT 373.950 520.950 376.050 523.050 ;
        RECT 377.100 522.150 378.900 523.950 ;
        RECT 362.100 511.950 364.200 514.050 ;
        RECT 370.200 510.600 372.000 516.600 ;
        RECT 394.500 516.600 395.700 523.950 ;
        RECT 397.950 519.300 398.850 530.700 ;
        RECT 401.100 526.050 402.900 527.850 ;
        RECT 416.700 526.050 417.600 538.200 ;
        RECT 418.950 526.950 421.050 529.050 ;
        RECT 400.950 523.950 403.050 526.050 ;
        RECT 415.950 523.950 418.050 526.050 ;
        RECT 419.100 525.150 420.900 526.950 ;
        RECT 422.100 526.050 423.900 527.850 ;
        RECT 424.950 526.950 427.050 529.050 ;
        RECT 421.950 523.950 424.050 526.050 ;
        RECT 425.100 525.150 426.900 526.950 ;
        RECT 440.700 526.050 441.600 538.200 ;
        RECT 442.950 526.950 445.050 529.050 ;
        RECT 439.950 523.950 442.050 526.050 ;
        RECT 443.100 525.150 444.900 526.950 ;
        RECT 446.100 526.050 447.900 527.850 ;
        RECT 448.950 526.950 451.050 529.050 ;
        RECT 445.950 523.950 448.050 526.050 ;
        RECT 449.100 525.150 450.900 526.950 ;
        RECT 396.600 518.400 398.850 519.300 ;
        RECT 416.700 520.200 417.600 523.950 ;
        RECT 440.700 520.200 441.600 523.950 ;
        RECT 416.700 519.000 420.000 520.200 ;
        RECT 440.700 519.000 444.000 520.200 ;
        RECT 396.600 517.500 402.600 518.400 ;
        RECT 394.500 510.600 396.300 516.600 ;
        RECT 401.400 513.600 402.600 517.500 ;
        RECT 400.800 510.600 402.600 513.600 ;
        RECT 418.200 510.600 420.000 519.000 ;
        RECT 442.200 510.600 444.000 519.000 ;
        RECT 458.550 514.050 459.450 541.950 ;
        RECT 463.800 539.400 465.600 545.400 ;
        RECT 464.700 539.100 465.600 539.400 ;
        RECT 469.800 539.400 471.600 545.400 ;
        RECT 487.800 539.400 489.600 545.400 ;
        RECT 469.800 539.100 471.300 539.400 ;
        RECT 464.700 538.200 471.300 539.100 ;
        RECT 488.700 539.100 489.600 539.400 ;
        RECT 493.800 539.400 495.600 545.400 ;
        RECT 502.950 541.950 505.050 544.050 ;
        RECT 493.800 539.100 495.300 539.400 ;
        RECT 488.700 538.200 495.300 539.100 ;
        RECT 464.700 526.050 465.600 538.200 ;
        RECT 466.950 526.950 469.050 529.050 ;
        RECT 463.950 523.950 466.050 526.050 ;
        RECT 467.100 525.150 468.900 526.950 ;
        RECT 470.100 526.050 471.900 527.850 ;
        RECT 472.950 526.950 475.050 529.050 ;
        RECT 469.950 523.950 472.050 526.050 ;
        RECT 473.100 525.150 474.900 526.950 ;
        RECT 488.700 526.050 489.600 538.200 ;
        RECT 490.950 526.950 493.050 529.050 ;
        RECT 487.950 523.950 490.050 526.050 ;
        RECT 491.100 525.150 492.900 526.950 ;
        RECT 494.100 526.050 495.900 527.850 ;
        RECT 496.950 526.950 499.050 529.050 ;
        RECT 493.950 523.950 496.050 526.050 ;
        RECT 497.100 525.150 498.900 526.950 ;
        RECT 464.700 520.200 465.600 523.950 ;
        RECT 488.700 520.200 489.600 523.950 ;
        RECT 464.700 519.000 468.000 520.200 ;
        RECT 488.700 519.000 492.000 520.200 ;
        RECT 458.100 511.950 460.200 514.050 ;
        RECT 466.200 510.600 468.000 519.000 ;
        RECT 490.200 510.600 492.000 519.000 ;
        RECT 503.550 517.050 504.450 541.950 ;
        RECT 509.400 534.300 511.200 545.400 ;
        RECT 515.400 534.300 517.200 545.400 ;
        RECT 509.400 533.400 517.200 534.300 ;
        RECT 518.400 533.400 520.200 545.400 ;
        RECT 539.400 539.400 541.200 545.400 ;
        RECT 508.950 526.950 511.050 529.050 ;
        RECT 509.100 525.150 510.900 526.950 ;
        RECT 512.100 526.050 513.900 527.850 ;
        RECT 514.950 526.950 517.050 529.050 ;
        RECT 511.950 523.950 514.050 526.050 ;
        RECT 515.100 525.150 516.900 526.950 ;
        RECT 518.400 526.050 519.600 533.400 ;
        RECT 535.950 526.950 538.050 529.050 ;
        RECT 517.950 523.950 520.050 526.050 ;
        RECT 536.100 525.150 537.900 526.950 ;
        RECT 539.850 526.050 541.050 539.400 ;
        RECT 559.800 533.400 561.600 545.400 ;
        RECT 562.800 534.300 564.600 545.400 ;
        RECT 568.800 534.300 570.600 545.400 ;
        RECT 584.400 539.400 586.200 545.400 ;
        RECT 584.700 539.100 586.200 539.400 ;
        RECT 590.400 539.400 592.200 545.400 ;
        RECT 608.400 539.400 610.200 545.400 ;
        RECT 590.400 539.100 591.300 539.400 ;
        RECT 584.700 538.200 591.300 539.100 ;
        RECT 562.800 533.400 570.600 534.300 ;
        RECT 541.950 526.950 544.050 529.050 ;
        RECT 538.950 523.950 541.050 526.050 ;
        RECT 542.100 525.150 543.900 526.950 ;
        RECT 545.100 526.050 546.900 527.850 ;
        RECT 560.400 526.050 561.600 533.400 ;
        RECT 562.950 526.950 565.050 529.050 ;
        RECT 544.950 523.950 547.050 526.050 ;
        RECT 559.950 523.950 562.050 526.050 ;
        RECT 563.100 525.150 564.900 526.950 ;
        RECT 566.100 526.050 567.900 527.850 ;
        RECT 568.950 526.950 571.050 529.050 ;
        RECT 580.950 526.950 583.050 529.050 ;
        RECT 565.950 523.950 568.050 526.050 ;
        RECT 569.100 525.150 570.900 526.950 ;
        RECT 581.100 525.150 582.900 526.950 ;
        RECT 584.100 526.050 585.900 527.850 ;
        RECT 586.950 526.950 589.050 529.050 ;
        RECT 583.950 523.950 586.050 526.050 ;
        RECT 587.100 525.150 588.900 526.950 ;
        RECT 590.400 526.050 591.300 538.200 ;
        RECT 608.400 532.050 609.600 539.400 ;
        RECT 625.800 533.400 627.600 545.400 ;
        RECT 628.800 534.300 630.600 545.400 ;
        RECT 634.800 534.300 636.600 545.400 ;
        RECT 640.950 541.950 643.050 544.050 ;
        RECT 628.800 533.400 636.600 534.300 ;
        RECT 605.100 526.050 606.900 527.850 ;
        RECT 607.950 526.950 610.050 532.050 ;
        RECT 589.950 523.950 592.050 526.050 ;
        RECT 604.950 523.950 607.050 526.050 ;
        RECT 502.950 514.950 505.050 517.050 ;
        RECT 518.400 516.600 519.600 523.950 ;
        RECT 538.950 519.750 540.150 523.950 ;
        RECT 536.400 518.700 540.150 519.750 ;
        RECT 536.400 516.600 537.600 518.700 ;
        RECT 514.500 515.400 519.600 516.600 ;
        RECT 514.500 510.600 516.300 515.400 ;
        RECT 535.800 510.600 537.600 516.600 ;
        RECT 538.800 515.700 546.600 517.050 ;
        RECT 538.800 510.600 540.600 515.700 ;
        RECT 544.800 510.600 546.600 515.700 ;
        RECT 560.400 516.600 561.600 523.950 ;
        RECT 590.400 520.200 591.300 523.950 ;
        RECT 588.000 519.000 591.300 520.200 ;
        RECT 560.400 515.400 565.500 516.600 ;
        RECT 563.700 510.600 565.500 515.400 ;
        RECT 588.000 510.600 589.800 519.000 ;
        RECT 608.400 513.600 609.600 526.950 ;
        RECT 626.400 526.050 627.600 533.400 ;
        RECT 628.950 526.950 631.050 529.050 ;
        RECT 625.950 523.950 628.050 526.050 ;
        RECT 629.100 525.150 630.900 526.950 ;
        RECT 632.100 526.050 633.900 527.850 ;
        RECT 634.950 526.950 637.050 529.050 ;
        RECT 631.950 523.950 634.050 526.050 ;
        RECT 635.100 525.150 636.900 526.950 ;
        RECT 626.400 516.600 627.600 523.950 ;
        RECT 641.550 520.050 642.450 541.950 ;
        RECT 649.800 539.400 651.600 545.400 ;
        RECT 650.700 539.100 651.600 539.400 ;
        RECT 655.800 539.400 657.600 545.400 ;
        RECT 664.950 541.950 667.050 544.050 ;
        RECT 655.800 539.100 657.300 539.400 ;
        RECT 650.700 538.200 657.300 539.100 ;
        RECT 650.700 526.050 651.600 538.200 ;
        RECT 652.950 526.950 655.050 529.050 ;
        RECT 649.950 523.950 652.050 526.050 ;
        RECT 653.100 525.150 654.900 526.950 ;
        RECT 656.100 526.050 657.900 527.850 ;
        RECT 658.950 526.950 661.050 529.050 ;
        RECT 655.950 523.950 658.050 526.050 ;
        RECT 659.100 525.150 660.900 526.950 ;
        RECT 650.700 520.200 651.600 523.950 ;
        RECT 640.950 517.950 643.050 520.050 ;
        RECT 650.700 519.000 654.000 520.200 ;
        RECT 665.550 520.050 666.450 541.950 ;
        RECT 673.800 539.400 675.600 545.400 ;
        RECT 674.700 539.100 675.600 539.400 ;
        RECT 679.800 539.400 681.600 545.400 ;
        RECT 700.800 539.400 702.600 545.400 ;
        RECT 722.400 539.400 724.200 545.400 ;
        RECT 742.800 544.500 750.600 545.400 ;
        RECT 679.800 539.100 681.300 539.400 ;
        RECT 674.700 538.200 681.300 539.100 ;
        RECT 674.700 526.050 675.600 538.200 ;
        RECT 676.950 526.950 679.050 529.050 ;
        RECT 673.950 523.950 676.050 526.050 ;
        RECT 677.100 525.150 678.900 526.950 ;
        RECT 680.100 526.050 681.900 527.850 ;
        RECT 682.950 526.950 685.050 529.050 ;
        RECT 679.950 523.950 682.050 526.050 ;
        RECT 683.100 525.150 684.900 526.950 ;
        RECT 695.100 526.050 696.900 527.850 ;
        RECT 697.950 526.950 700.050 529.050 ;
        RECT 694.950 523.950 697.050 526.050 ;
        RECT 698.100 525.150 699.900 526.950 ;
        RECT 700.950 526.050 702.150 539.400 ;
        RECT 703.950 526.950 706.050 529.050 ;
        RECT 718.950 526.950 721.050 529.050 ;
        RECT 700.950 523.950 703.050 526.050 ;
        RECT 704.100 525.150 705.900 526.950 ;
        RECT 719.100 525.150 720.900 526.950 ;
        RECT 722.400 526.050 723.600 539.400 ;
        RECT 742.800 533.400 744.600 544.500 ;
        RECT 745.800 532.500 747.600 543.600 ;
        RECT 748.800 534.600 750.600 544.500 ;
        RECT 754.800 534.600 756.600 545.400 ;
        RECT 769.800 539.400 771.600 545.400 ;
        RECT 748.800 533.700 756.600 534.600 ;
        RECT 770.700 539.100 771.600 539.400 ;
        RECT 775.800 539.400 777.600 545.400 ;
        RECT 793.800 539.400 795.600 545.400 ;
        RECT 802.950 541.950 805.050 544.050 ;
        RECT 775.800 539.100 777.300 539.400 ;
        RECT 770.700 538.200 777.300 539.100 ;
        RECT 745.800 531.600 750.900 532.500 ;
        RECT 724.950 526.950 727.050 529.050 ;
        RECT 721.950 523.950 724.050 526.050 ;
        RECT 725.100 525.150 726.900 526.950 ;
        RECT 750.000 526.050 750.900 531.600 ;
        RECT 770.700 526.050 771.600 538.200 ;
        RECT 794.400 532.050 795.600 539.400 ;
        RECT 772.950 526.950 775.050 529.050 ;
        RECT 742.950 523.950 745.050 526.050 ;
        RECT 674.700 520.200 675.600 523.950 ;
        RECT 626.400 515.400 631.500 516.600 ;
        RECT 608.400 510.600 610.200 513.600 ;
        RECT 629.700 510.600 631.500 515.400 ;
        RECT 652.200 510.600 654.000 519.000 ;
        RECT 664.950 517.950 667.050 520.050 ;
        RECT 674.700 519.000 678.000 520.200 ;
        RECT 676.200 510.600 678.000 519.000 ;
        RECT 701.850 519.750 703.050 523.950 ;
        RECT 701.850 518.700 705.600 519.750 ;
        RECT 695.400 515.700 703.200 517.050 ;
        RECT 695.400 510.600 697.200 515.700 ;
        RECT 701.400 510.600 703.200 515.700 ;
        RECT 704.400 516.600 705.600 518.700 ;
        RECT 722.400 518.700 723.600 523.950 ;
        RECT 743.100 522.150 744.900 523.950 ;
        RECT 746.100 523.050 747.900 524.850 ;
        RECT 748.950 523.950 751.050 526.050 ;
        RECT 745.950 520.950 748.050 523.050 ;
        RECT 722.400 517.800 726.600 518.700 ;
        RECT 704.400 510.600 706.200 516.600 ;
        RECT 724.800 510.600 726.600 517.800 ;
        RECT 750.000 516.600 751.050 523.950 ;
        RECT 752.100 523.050 753.900 524.850 ;
        RECT 754.950 523.950 757.050 526.050 ;
        RECT 769.950 523.950 772.050 526.050 ;
        RECT 773.100 525.150 774.900 526.950 ;
        RECT 776.100 526.050 777.900 527.850 ;
        RECT 778.950 526.950 781.050 529.050 ;
        RECT 793.950 526.950 796.050 532.050 ;
        RECT 775.950 523.950 778.050 526.050 ;
        RECT 779.100 525.150 780.900 526.950 ;
        RECT 751.950 520.950 754.050 523.050 ;
        RECT 755.100 522.150 756.900 523.950 ;
        RECT 770.700 520.200 771.600 523.950 ;
        RECT 770.700 519.000 774.000 520.200 ;
        RECT 750.000 510.600 751.800 516.600 ;
        RECT 772.200 510.600 774.000 519.000 ;
        RECT 794.400 513.600 795.600 526.950 ;
        RECT 797.100 526.050 798.900 527.850 ;
        RECT 796.950 523.950 799.050 526.050 ;
        RECT 803.550 514.050 804.450 541.950 ;
        RECT 812.400 539.400 814.200 545.400 ;
        RECT 812.700 539.100 814.200 539.400 ;
        RECT 818.400 539.400 820.200 545.400 ;
        RECT 835.800 539.400 837.600 545.400 ;
        RECT 853.800 539.400 855.600 545.400 ;
        RECT 818.400 539.100 819.300 539.400 ;
        RECT 812.700 538.200 819.300 539.100 ;
        RECT 808.950 526.950 811.050 529.050 ;
        RECT 809.100 525.150 810.900 526.950 ;
        RECT 812.100 526.050 813.900 527.850 ;
        RECT 814.950 526.950 817.050 529.050 ;
        RECT 811.950 523.950 814.050 526.050 ;
        RECT 815.100 525.150 816.900 526.950 ;
        RECT 818.400 526.050 819.300 538.200 ;
        RECT 836.400 532.050 837.600 539.400 ;
        RECT 854.700 539.100 855.600 539.400 ;
        RECT 859.800 539.400 861.600 545.400 ;
        RECT 859.800 539.100 861.300 539.400 ;
        RECT 854.700 538.200 861.300 539.100 ;
        RECT 835.950 526.950 838.050 532.050 ;
        RECT 817.950 523.950 820.050 526.050 ;
        RECT 818.400 520.200 819.300 523.950 ;
        RECT 816.000 519.000 819.300 520.200 ;
        RECT 793.800 510.600 795.600 513.600 ;
        RECT 802.950 511.950 805.050 514.050 ;
        RECT 816.000 510.600 817.800 519.000 ;
        RECT 836.400 513.600 837.600 526.950 ;
        RECT 839.100 526.050 840.900 527.850 ;
        RECT 854.700 526.050 855.600 538.200 ;
        RECT 875.400 534.300 877.200 545.400 ;
        RECT 881.400 534.300 883.200 545.400 ;
        RECT 875.400 533.400 883.200 534.300 ;
        RECT 884.400 533.400 886.200 545.400 ;
        RECT 902.400 539.400 904.200 545.400 ;
        RECT 856.950 526.950 859.050 529.050 ;
        RECT 838.950 523.950 841.050 526.050 ;
        RECT 853.950 523.950 856.050 526.050 ;
        RECT 857.100 525.150 858.900 526.950 ;
        RECT 860.100 526.050 861.900 527.850 ;
        RECT 862.950 526.950 865.050 529.050 ;
        RECT 874.950 526.950 877.050 529.050 ;
        RECT 859.950 523.950 862.050 526.050 ;
        RECT 863.100 525.150 864.900 526.950 ;
        RECT 875.100 525.150 876.900 526.950 ;
        RECT 878.100 526.050 879.900 527.850 ;
        RECT 880.950 526.950 883.050 529.050 ;
        RECT 877.950 523.950 880.050 526.050 ;
        RECT 881.100 525.150 882.900 526.950 ;
        RECT 884.400 526.050 885.600 533.400 ;
        RECT 892.950 532.950 895.050 535.050 ;
        RECT 883.950 523.950 886.050 526.050 ;
        RECT 854.700 520.200 855.600 523.950 ;
        RECT 854.700 519.000 858.000 520.200 ;
        RECT 835.800 510.600 837.600 513.600 ;
        RECT 856.200 510.600 858.000 519.000 ;
        RECT 884.400 516.600 885.600 523.950 ;
        RECT 893.550 517.050 894.450 532.950 ;
        RECT 902.400 532.050 903.600 539.400 ;
        RECT 899.100 526.050 900.900 527.850 ;
        RECT 901.950 526.950 904.050 532.050 ;
        RECT 898.950 523.950 901.050 526.050 ;
        RECT 880.500 515.400 885.600 516.600 ;
        RECT 880.500 510.600 882.300 515.400 ;
        RECT 892.950 514.950 895.050 517.050 ;
        RECT 902.400 513.600 903.600 526.950 ;
        RECT 902.400 510.600 904.200 513.600 ;
        RECT 17.700 501.600 19.500 506.400 ;
        RECT 14.400 500.400 19.500 501.600 ;
        RECT 14.400 493.050 15.600 500.400 ;
        RECT 42.000 498.000 43.800 506.400 ;
        RECT 52.950 502.950 55.050 505.050 ;
        RECT 62.400 503.400 64.200 506.400 ;
        RECT 42.000 496.800 45.300 498.000 ;
        RECT 44.400 493.050 45.300 496.800 ;
        RECT 13.950 490.950 16.050 493.050 ;
        RECT 14.400 483.600 15.600 490.950 ;
        RECT 17.100 490.050 18.900 491.850 ;
        RECT 19.950 490.950 22.050 493.050 ;
        RECT 16.950 487.950 19.050 490.050 ;
        RECT 20.100 489.150 21.900 490.950 ;
        RECT 23.100 490.050 24.900 491.850 ;
        RECT 35.100 490.050 36.900 491.850 ;
        RECT 37.950 490.950 40.050 493.050 ;
        RECT 22.950 487.950 25.050 490.050 ;
        RECT 34.950 487.950 37.050 490.050 ;
        RECT 38.100 489.150 39.900 490.950 ;
        RECT 41.100 490.050 42.900 491.850 ;
        RECT 43.950 490.950 46.050 493.050 ;
        RECT 40.950 487.950 43.050 490.050 ;
        RECT 13.800 471.600 15.600 483.600 ;
        RECT 16.800 482.700 24.600 483.600 ;
        RECT 16.800 471.600 18.600 482.700 ;
        RECT 22.800 471.600 24.600 482.700 ;
        RECT 44.400 478.800 45.300 490.950 ;
        RECT 38.700 477.900 45.300 478.800 ;
        RECT 38.700 477.600 40.200 477.900 ;
        RECT 38.400 471.600 40.200 477.600 ;
        RECT 44.400 477.600 45.300 477.900 ;
        RECT 44.400 471.600 46.200 477.600 ;
        RECT 53.550 475.050 54.450 502.950 ;
        RECT 58.950 490.950 61.050 493.050 ;
        RECT 59.100 489.150 60.900 490.950 ;
        RECT 62.400 490.050 63.600 503.400 ;
        RECT 80.400 499.200 82.200 506.400 ;
        RECT 94.950 502.950 97.050 505.050 ;
        RECT 80.400 498.300 84.600 499.200 ;
        RECT 83.400 493.050 84.600 498.300 ;
        RECT 80.100 490.050 81.900 491.850 ;
        RECT 82.950 490.950 85.050 493.050 ;
        RECT 61.950 484.950 64.050 490.050 ;
        RECT 79.950 487.950 82.050 490.050 ;
        RECT 49.950 473.550 54.450 475.050 ;
        RECT 62.400 477.600 63.600 484.950 ;
        RECT 83.400 477.600 84.600 490.950 ;
        RECT 86.100 490.050 87.900 491.850 ;
        RECT 85.950 487.950 88.050 490.050 ;
        RECT 95.550 481.050 96.450 502.950 ;
        RECT 108.000 500.400 109.800 506.400 ;
        RECT 101.100 493.050 102.900 494.850 ;
        RECT 103.950 493.950 106.050 496.050 ;
        RECT 100.950 490.950 103.050 493.050 ;
        RECT 104.100 492.150 105.900 493.950 ;
        RECT 108.000 493.050 109.050 500.400 ;
        RECT 127.800 499.200 129.600 506.400 ;
        RECT 130.950 502.950 133.050 505.050 ;
        RECT 146.400 503.400 148.200 506.400 ;
        RECT 125.400 498.300 129.600 499.200 ;
        RECT 109.950 493.950 112.050 496.050 ;
        RECT 106.950 490.950 109.050 493.050 ;
        RECT 110.100 492.150 111.900 493.950 ;
        RECT 113.100 493.050 114.900 494.850 ;
        RECT 125.400 493.050 126.600 498.300 ;
        RECT 131.550 496.050 132.450 502.950 ;
        RECT 147.300 499.200 148.200 503.400 ;
        RECT 152.400 500.400 154.200 506.400 ;
        RECT 147.300 498.300 150.600 499.200 ;
        RECT 148.800 497.400 150.600 498.300 ;
        RECT 130.950 493.950 133.050 496.050 ;
        RECT 112.950 490.950 115.050 493.050 ;
        RECT 108.000 485.400 108.900 490.950 ;
        RECT 122.100 490.050 123.900 491.850 ;
        RECT 124.950 490.950 127.050 493.050 ;
        RECT 121.950 487.950 124.050 490.050 ;
        RECT 103.800 484.500 108.900 485.400 ;
        RECT 94.950 478.950 97.050 481.050 ;
        RECT 49.950 472.950 54.000 473.550 ;
        RECT 62.400 471.600 64.200 477.600 ;
        RECT 82.800 471.600 84.600 477.600 ;
        RECT 100.800 472.500 102.600 483.600 ;
        RECT 103.800 473.400 105.600 484.500 ;
        RECT 106.800 482.400 114.600 483.300 ;
        RECT 106.800 472.500 108.600 482.400 ;
        RECT 100.800 471.600 108.600 472.500 ;
        RECT 112.800 471.600 114.600 482.400 ;
        RECT 125.400 477.600 126.600 490.950 ;
        RECT 128.100 490.050 129.900 491.850 ;
        RECT 143.100 490.050 144.900 491.850 ;
        RECT 145.950 490.950 148.050 493.050 ;
        RECT 127.950 487.950 130.050 490.050 ;
        RECT 142.950 487.950 145.050 490.050 ;
        RECT 146.100 489.150 147.900 490.950 ;
        RECT 149.700 486.900 150.600 497.400 ;
        RECT 153.000 493.050 154.050 500.400 ;
        RECT 172.800 499.500 174.600 506.400 ;
        RECT 178.800 499.500 180.600 506.400 ;
        RECT 184.800 499.500 186.600 506.400 ;
        RECT 190.800 499.500 192.600 506.400 ;
        RECT 208.800 503.400 210.600 506.400 ;
        RECT 171.900 498.300 174.600 499.500 ;
        RECT 176.700 498.300 180.600 499.500 ;
        RECT 182.700 498.300 186.600 499.500 ;
        RECT 188.700 498.300 192.600 499.500 ;
        RECT 171.900 493.050 172.800 498.300 ;
        RECT 176.700 497.400 177.900 498.300 ;
        RECT 182.700 497.400 183.900 498.300 ;
        RECT 188.700 497.400 189.900 498.300 ;
        RECT 173.700 496.200 177.900 497.400 ;
        RECT 173.700 495.600 175.500 496.200 ;
        RECT 148.800 486.300 150.600 486.900 ;
        RECT 143.400 485.100 150.600 486.300 ;
        RECT 151.950 490.950 154.050 493.050 ;
        RECT 169.950 490.950 172.800 493.050 ;
        RECT 143.400 483.600 144.600 485.100 ;
        RECT 151.950 483.600 153.300 490.950 ;
        RECT 171.900 485.700 172.800 490.950 ;
        RECT 176.700 485.700 177.900 496.200 ;
        RECT 179.700 496.200 183.900 497.400 ;
        RECT 179.700 495.600 181.500 496.200 ;
        RECT 182.700 485.700 183.900 496.200 ;
        RECT 185.700 496.200 189.900 497.400 ;
        RECT 185.700 495.600 187.500 496.200 ;
        RECT 188.700 485.700 189.900 496.200 ;
        RECT 191.100 493.050 192.900 494.850 ;
        RECT 190.950 490.950 193.050 493.050 ;
        RECT 209.400 490.050 210.600 503.400 ;
        RECT 216.150 500.400 217.950 506.400 ;
        RECT 223.950 504.300 225.750 506.400 ;
        RECT 222.000 503.400 225.750 504.300 ;
        RECT 231.750 503.400 233.550 506.400 ;
        RECT 239.550 503.400 241.350 506.400 ;
        RECT 222.000 502.500 223.050 503.400 ;
        RECT 231.750 502.500 232.800 503.400 ;
        RECT 220.950 500.400 223.050 502.500 ;
        RECT 211.950 490.950 214.050 493.050 ;
        RECT 171.900 484.500 174.600 485.700 ;
        RECT 176.700 484.500 180.600 485.700 ;
        RECT 182.700 484.500 186.600 485.700 ;
        RECT 188.700 484.500 192.600 485.700 ;
        RECT 208.950 484.950 211.050 490.050 ;
        RECT 212.100 489.150 213.900 490.950 ;
        RECT 216.150 485.700 217.050 500.400 ;
        RECT 224.550 499.800 226.350 501.600 ;
        RECT 227.850 501.450 232.800 502.500 ;
        RECT 240.300 502.500 241.350 503.400 ;
        RECT 227.850 500.700 229.650 501.450 ;
        RECT 240.300 501.300 244.050 502.500 ;
        RECT 241.950 500.400 244.050 501.300 ;
        RECT 247.650 500.400 249.450 506.400 ;
        RECT 224.850 498.000 225.900 499.800 ;
        RECT 235.050 498.000 236.850 498.600 ;
        RECT 224.850 496.800 236.850 498.000 ;
        RECT 219.000 495.600 225.900 496.800 ;
        RECT 219.000 494.850 219.900 495.600 ;
        RECT 224.100 495.000 225.900 495.600 ;
        RECT 218.100 493.050 219.900 494.850 ;
        RECT 221.100 493.800 222.900 494.400 ;
        RECT 217.950 490.950 220.050 493.050 ;
        RECT 221.100 492.600 229.050 493.800 ;
        RECT 226.950 490.950 229.050 492.600 ;
        RECT 225.450 485.700 227.250 486.000 ;
        RECT 216.150 485.100 227.250 485.700 ;
        RECT 125.400 471.600 127.200 477.600 ;
        RECT 143.400 471.600 145.200 483.600 ;
        RECT 150.900 482.100 153.300 483.600 ;
        RECT 150.900 471.600 152.700 482.100 ;
        RECT 172.800 471.600 174.600 484.500 ;
        RECT 178.800 471.600 180.600 484.500 ;
        RECT 184.800 471.600 186.600 484.500 ;
        RECT 190.800 471.600 192.600 484.500 ;
        RECT 209.400 477.600 210.600 484.950 ;
        RECT 208.800 471.600 210.600 477.600 ;
        RECT 216.150 484.500 233.850 485.100 ;
        RECT 216.150 483.600 217.050 484.500 ;
        RECT 225.450 484.200 233.850 484.500 ;
        RECT 216.150 471.600 217.950 483.600 ;
        RECT 230.250 482.700 232.050 483.300 ;
        RECT 224.550 481.500 232.050 482.700 ;
        RECT 232.950 482.100 233.850 484.200 ;
        RECT 235.950 484.200 236.850 496.800 ;
        RECT 248.250 493.050 249.450 500.400 ;
        RECT 263.400 503.400 265.200 506.400 ;
        RECT 280.800 503.400 282.600 506.400 ;
        RECT 243.150 491.250 249.450 493.050 ;
        RECT 244.950 490.950 249.450 491.250 ;
        RECT 259.950 490.950 262.050 493.050 ;
        RECT 245.250 485.400 247.050 487.200 ;
        RECT 241.950 484.200 246.150 485.400 ;
        RECT 235.950 483.300 241.050 484.200 ;
        RECT 241.950 483.300 244.050 484.200 ;
        RECT 248.250 483.600 249.450 490.950 ;
        RECT 260.100 489.150 261.900 490.950 ;
        RECT 263.400 490.050 264.600 503.400 ;
        RECT 281.400 490.050 282.600 503.400 ;
        RECT 287.550 500.400 289.350 506.400 ;
        RECT 295.650 503.400 297.450 506.400 ;
        RECT 303.450 503.400 305.250 506.400 ;
        RECT 311.250 504.300 313.050 506.400 ;
        RECT 311.250 503.400 315.000 504.300 ;
        RECT 295.650 502.500 296.700 503.400 ;
        RECT 292.950 501.300 296.700 502.500 ;
        RECT 304.200 502.500 305.250 503.400 ;
        RECT 313.950 502.500 315.000 503.400 ;
        RECT 304.200 501.450 309.150 502.500 ;
        RECT 292.950 500.400 295.050 501.300 ;
        RECT 307.350 500.700 309.150 501.450 ;
        RECT 287.550 493.050 288.750 500.400 ;
        RECT 310.650 499.800 312.450 501.600 ;
        RECT 313.950 500.400 316.050 502.500 ;
        RECT 319.050 500.400 320.850 506.400 ;
        RECT 336.300 502.200 338.100 506.400 ;
        RECT 300.150 498.000 301.950 498.600 ;
        RECT 311.100 498.000 312.150 499.800 ;
        RECT 300.150 496.800 312.150 498.000 ;
        RECT 283.950 490.950 286.050 493.050 ;
        RECT 287.550 491.250 293.850 493.050 ;
        RECT 287.550 490.950 292.050 491.250 ;
        RECT 262.950 484.950 265.050 490.050 ;
        RECT 280.950 484.950 283.050 490.050 ;
        RECT 284.100 489.150 285.900 490.950 ;
        RECT 240.150 482.400 241.050 483.300 ;
        RECT 237.450 482.100 239.250 482.400 ;
        RECT 224.550 480.600 225.750 481.500 ;
        RECT 232.950 481.200 239.250 482.100 ;
        RECT 237.450 480.600 239.250 481.200 ;
        RECT 240.150 480.600 242.850 482.400 ;
        RECT 220.950 478.500 225.750 480.600 ;
        RECT 228.450 479.550 230.250 480.300 ;
        RECT 233.250 479.550 235.050 480.300 ;
        RECT 228.450 478.500 235.050 479.550 ;
        RECT 224.550 477.600 225.750 478.500 ;
        RECT 224.550 471.600 226.350 477.600 ;
        RECT 232.350 471.600 234.150 478.500 ;
        RECT 240.150 477.600 244.050 479.700 ;
        RECT 240.150 471.600 241.950 477.600 ;
        RECT 247.650 471.600 249.450 483.600 ;
        RECT 263.400 477.600 264.600 484.950 ;
        RECT 281.400 477.600 282.600 484.950 ;
        RECT 263.400 471.600 265.200 477.600 ;
        RECT 280.800 471.600 282.600 477.600 ;
        RECT 287.550 483.600 288.750 490.950 ;
        RECT 289.950 485.400 291.750 487.200 ;
        RECT 290.850 484.200 295.050 485.400 ;
        RECT 300.150 484.200 301.050 496.800 ;
        RECT 311.100 495.600 318.000 496.800 ;
        RECT 311.100 495.000 312.900 495.600 ;
        RECT 317.100 494.850 318.000 495.600 ;
        RECT 314.100 493.800 315.900 494.400 ;
        RECT 307.950 492.600 315.900 493.800 ;
        RECT 317.100 493.050 318.900 494.850 ;
        RECT 307.950 490.950 310.050 492.600 ;
        RECT 316.950 490.950 319.050 493.050 ;
        RECT 309.750 485.700 311.550 486.000 ;
        RECT 319.950 485.700 320.850 500.400 ;
        RECT 335.400 500.400 338.100 502.200 ;
        RECT 335.400 493.050 336.300 500.400 ;
        RECT 338.100 498.600 339.900 499.500 ;
        RECT 343.800 498.600 345.600 506.400 ;
        RECT 338.100 497.700 345.600 498.600 ;
        RECT 363.000 498.000 364.800 506.400 ;
        RECT 385.800 503.400 387.600 506.400 ;
        RECT 334.950 490.950 337.050 493.050 ;
        RECT 337.950 490.950 340.050 493.050 ;
        RECT 309.750 485.100 320.850 485.700 ;
        RECT 287.550 471.600 289.350 483.600 ;
        RECT 292.950 483.300 295.050 484.200 ;
        RECT 295.950 483.300 301.050 484.200 ;
        RECT 303.150 484.500 320.850 485.100 ;
        RECT 303.150 484.200 311.550 484.500 ;
        RECT 295.950 482.400 296.850 483.300 ;
        RECT 294.150 480.600 296.850 482.400 ;
        RECT 297.750 482.100 299.550 482.400 ;
        RECT 303.150 482.100 304.050 484.200 ;
        RECT 319.950 483.600 320.850 484.500 ;
        RECT 335.400 483.600 336.300 490.950 ;
        RECT 338.100 489.150 339.900 490.950 ;
        RECT 297.750 481.200 304.050 482.100 ;
        RECT 304.950 482.700 306.750 483.300 ;
        RECT 304.950 481.500 312.450 482.700 ;
        RECT 297.750 480.600 299.550 481.200 ;
        RECT 311.250 480.600 312.450 481.500 ;
        RECT 292.950 477.600 296.850 479.700 ;
        RECT 301.950 479.550 303.750 480.300 ;
        RECT 306.750 479.550 308.550 480.300 ;
        RECT 301.950 478.500 308.550 479.550 ;
        RECT 311.250 478.500 316.050 480.600 ;
        RECT 295.050 471.600 296.850 477.600 ;
        RECT 302.850 471.600 304.650 478.500 ;
        RECT 311.250 477.600 312.450 478.500 ;
        RECT 310.650 471.600 312.450 477.600 ;
        RECT 319.050 471.600 320.850 483.600 ;
        RECT 334.500 471.600 336.300 483.600 ;
        RECT 341.700 477.600 342.600 497.700 ;
        RECT 363.000 496.800 366.300 498.000 ;
        RECT 344.100 493.050 345.900 494.850 ;
        RECT 365.400 493.050 366.300 496.800 ;
        RECT 382.950 493.950 385.050 496.050 ;
        RECT 343.950 490.950 346.050 493.050 ;
        RECT 356.100 490.050 357.900 491.850 ;
        RECT 358.950 490.950 361.050 493.050 ;
        RECT 355.950 487.950 358.050 490.050 ;
        RECT 359.100 489.150 360.900 490.950 ;
        RECT 362.100 490.050 363.900 491.850 ;
        RECT 364.950 490.950 367.050 493.050 ;
        RECT 383.100 492.150 384.900 493.950 ;
        RECT 386.400 493.050 387.300 503.400 ;
        RECT 394.950 502.950 397.050 505.050 ;
        RECT 395.550 496.050 396.450 502.950 ;
        RECT 407.700 501.600 409.500 506.400 ;
        RECT 404.400 500.400 409.500 501.600 ;
        RECT 388.950 493.950 391.050 496.050 ;
        RECT 394.950 493.950 397.050 496.050 ;
        RECT 385.950 490.950 388.050 493.050 ;
        RECT 389.100 492.150 390.900 493.950 ;
        RECT 404.400 493.050 405.600 500.400 ;
        RECT 432.000 498.000 433.800 506.400 ;
        RECT 451.800 503.400 453.600 506.400 ;
        RECT 432.000 496.800 435.300 498.000 ;
        RECT 434.400 493.050 435.300 496.800 ;
        RECT 403.950 490.950 406.050 493.050 ;
        RECT 361.950 487.950 364.050 490.050 ;
        RECT 365.400 478.800 366.300 490.950 ;
        RECT 386.400 483.600 387.300 490.950 ;
        RECT 404.400 483.600 405.600 490.950 ;
        RECT 407.100 490.050 408.900 491.850 ;
        RECT 409.950 490.950 412.050 493.050 ;
        RECT 406.950 487.950 409.050 490.050 ;
        RECT 410.100 489.150 411.900 490.950 ;
        RECT 413.100 490.050 414.900 491.850 ;
        RECT 425.100 490.050 426.900 491.850 ;
        RECT 427.950 490.950 430.050 493.050 ;
        RECT 412.950 487.950 415.050 490.050 ;
        RECT 424.950 487.950 427.050 490.050 ;
        RECT 428.100 489.150 429.900 490.950 ;
        RECT 431.100 490.050 432.900 491.850 ;
        RECT 433.950 490.950 436.050 493.050 ;
        RECT 430.950 487.950 433.050 490.050 ;
        RECT 359.700 477.900 366.300 478.800 ;
        RECT 359.700 477.600 361.200 477.900 ;
        RECT 340.800 471.600 342.600 477.600 ;
        RECT 359.400 471.600 361.200 477.600 ;
        RECT 365.400 477.600 366.300 477.900 ;
        RECT 383.700 482.400 387.300 483.600 ;
        RECT 365.400 471.600 367.200 477.600 ;
        RECT 383.700 471.600 385.500 482.400 ;
        RECT 403.800 471.600 405.600 483.600 ;
        RECT 406.800 482.700 414.600 483.600 ;
        RECT 406.800 471.600 408.600 482.700 ;
        RECT 412.800 471.600 414.600 482.700 ;
        RECT 434.400 478.800 435.300 490.950 ;
        RECT 452.400 490.050 453.600 503.400 ;
        RECT 460.950 502.950 463.050 505.050 ;
        RECT 454.950 490.950 457.050 493.050 ;
        RECT 451.950 484.950 454.050 490.050 ;
        RECT 455.100 489.150 456.900 490.950 ;
        RECT 457.950 484.950 460.050 487.050 ;
        RECT 428.700 477.900 435.300 478.800 ;
        RECT 428.700 477.600 430.200 477.900 ;
        RECT 428.400 471.600 430.200 477.600 ;
        RECT 434.400 477.600 435.300 477.900 ;
        RECT 452.400 477.600 453.600 484.950 ;
        RECT 458.550 478.050 459.450 484.950 ;
        RECT 461.550 481.050 462.450 502.950 ;
        RECT 474.000 498.000 475.800 506.400 ;
        RECT 484.950 502.950 487.050 505.050 ;
        RECT 474.000 496.800 477.300 498.000 ;
        RECT 476.400 493.050 477.300 496.800 ;
        RECT 467.100 490.050 468.900 491.850 ;
        RECT 469.950 490.950 472.050 493.050 ;
        RECT 466.950 487.950 469.050 490.050 ;
        RECT 470.100 489.150 471.900 490.950 ;
        RECT 473.100 490.050 474.900 491.850 ;
        RECT 475.950 490.950 478.050 493.050 ;
        RECT 472.950 487.950 475.050 490.050 ;
        RECT 460.950 478.950 463.050 481.050 ;
        RECT 476.400 478.800 477.300 490.950 ;
        RECT 485.550 481.050 486.450 502.950 ;
        RECT 496.200 498.000 498.000 506.400 ;
        RECT 520.200 498.000 522.000 506.400 ;
        RECT 494.700 496.800 498.000 498.000 ;
        RECT 518.700 496.800 522.000 498.000 ;
        RECT 542.400 503.400 544.200 506.400 ;
        RECT 488.100 493.950 490.200 496.050 ;
        RECT 484.950 478.950 487.050 481.050 ;
        RECT 434.400 471.600 436.200 477.600 ;
        RECT 451.800 471.600 453.600 477.600 ;
        RECT 457.950 475.950 460.050 478.050 ;
        RECT 470.700 477.900 477.300 478.800 ;
        RECT 488.550 478.050 489.450 493.950 ;
        RECT 494.700 493.050 495.600 496.800 ;
        RECT 518.700 493.050 519.600 496.800 ;
        RECT 493.950 490.950 496.050 493.050 ;
        RECT 494.700 478.800 495.600 490.950 ;
        RECT 497.100 490.050 498.900 491.850 ;
        RECT 499.950 490.950 502.050 493.050 ;
        RECT 496.950 487.950 499.050 490.050 ;
        RECT 500.100 489.150 501.900 490.950 ;
        RECT 503.100 490.050 504.900 491.850 ;
        RECT 517.950 490.950 520.050 493.050 ;
        RECT 502.950 487.950 505.050 490.050 ;
        RECT 518.700 478.800 519.600 490.950 ;
        RECT 521.100 490.050 522.900 491.850 ;
        RECT 523.950 490.950 526.050 493.050 ;
        RECT 520.950 487.950 523.050 490.050 ;
        RECT 524.100 489.150 525.900 490.950 ;
        RECT 527.100 490.050 528.900 491.850 ;
        RECT 538.950 490.950 541.050 493.050 ;
        RECT 526.950 487.950 529.050 490.050 ;
        RECT 539.100 489.150 540.900 490.950 ;
        RECT 542.400 490.050 543.600 503.400 ;
        RECT 557.400 501.300 559.200 506.400 ;
        RECT 563.400 501.300 565.200 506.400 ;
        RECT 557.400 499.950 565.200 501.300 ;
        RECT 566.400 500.400 568.200 506.400 ;
        RECT 571.950 502.950 574.050 505.050 ;
        RECT 583.800 503.400 585.600 506.400 ;
        RECT 566.400 498.300 567.600 500.400 ;
        RECT 563.850 497.250 567.600 498.300 ;
        RECT 563.850 493.050 565.050 497.250 ;
        RECT 556.950 490.950 559.050 493.050 ;
        RECT 541.950 484.950 544.050 490.050 ;
        RECT 557.100 489.150 558.900 490.950 ;
        RECT 560.100 490.050 561.900 491.850 ;
        RECT 562.950 490.950 565.050 493.050 ;
        RECT 559.950 487.950 562.050 490.050 ;
        RECT 470.700 477.600 472.200 477.900 ;
        RECT 470.400 471.600 472.200 477.600 ;
        RECT 476.400 477.600 477.300 477.900 ;
        RECT 476.400 471.600 478.200 477.600 ;
        RECT 487.950 475.950 490.050 478.050 ;
        RECT 494.700 477.900 501.300 478.800 ;
        RECT 494.700 477.600 495.600 477.900 ;
        RECT 493.800 471.600 495.600 477.600 ;
        RECT 499.800 477.600 501.300 477.900 ;
        RECT 518.700 477.900 525.300 478.800 ;
        RECT 518.700 477.600 519.600 477.900 ;
        RECT 499.800 471.600 501.600 477.600 ;
        RECT 517.800 471.600 519.600 477.600 ;
        RECT 523.800 477.600 525.300 477.900 ;
        RECT 542.400 477.600 543.600 484.950 ;
        RECT 562.950 477.600 564.150 490.950 ;
        RECT 566.100 490.050 567.900 491.850 ;
        RECT 565.950 487.950 568.050 490.050 ;
        RECT 572.550 487.050 573.450 502.950 ;
        RECT 584.400 490.050 585.600 503.400 ;
        RECT 606.000 498.000 607.800 506.400 ;
        RECT 626.400 499.200 628.200 506.400 ;
        RECT 649.800 503.400 651.600 506.400 ;
        RECT 626.400 498.300 630.600 499.200 ;
        RECT 606.000 496.800 609.300 498.000 ;
        RECT 608.400 493.050 609.300 496.800 ;
        RECT 616.950 493.950 619.050 496.050 ;
        RECT 586.950 490.950 589.050 493.050 ;
        RECT 571.950 484.950 574.050 487.050 ;
        RECT 583.950 484.950 586.050 490.050 ;
        RECT 587.100 489.150 588.900 490.950 ;
        RECT 599.100 490.050 600.900 491.850 ;
        RECT 601.950 490.950 604.050 493.050 ;
        RECT 598.950 487.950 601.050 490.050 ;
        RECT 602.100 489.150 603.900 490.950 ;
        RECT 605.100 490.050 606.900 491.850 ;
        RECT 607.950 490.950 610.050 493.050 ;
        RECT 604.950 487.950 607.050 490.050 ;
        RECT 584.400 477.600 585.600 484.950 ;
        RECT 608.400 478.800 609.300 490.950 ;
        RECT 617.550 481.050 618.450 493.950 ;
        RECT 629.400 493.050 630.600 498.300 ;
        RECT 646.950 493.950 649.050 496.050 ;
        RECT 626.100 490.050 627.900 491.850 ;
        RECT 628.950 490.950 631.050 493.050 ;
        RECT 647.100 492.150 648.900 493.950 ;
        RECT 650.400 493.050 651.300 503.400 ;
        RECT 668.400 499.200 670.200 506.400 ;
        RECT 686.400 501.300 688.200 506.400 ;
        RECT 692.400 501.300 694.200 506.400 ;
        RECT 686.400 499.950 694.200 501.300 ;
        RECT 695.400 500.400 697.200 506.400 ;
        RECT 668.400 498.300 672.600 499.200 ;
        RECT 695.400 498.300 696.600 500.400 ;
        RECT 652.950 493.950 655.050 496.050 ;
        RECT 625.950 487.950 628.050 490.050 ;
        RECT 616.950 478.950 619.050 481.050 ;
        RECT 602.700 477.900 609.300 478.800 ;
        RECT 602.700 477.600 604.200 477.900 ;
        RECT 523.800 471.600 525.600 477.600 ;
        RECT 542.400 471.600 544.200 477.600 ;
        RECT 562.800 471.600 564.600 477.600 ;
        RECT 583.800 471.600 585.600 477.600 ;
        RECT 602.400 471.600 604.200 477.600 ;
        RECT 608.400 477.600 609.300 477.900 ;
        RECT 629.400 477.600 630.600 490.950 ;
        RECT 632.100 490.050 633.900 491.850 ;
        RECT 649.950 490.950 652.050 493.050 ;
        RECT 653.100 492.150 654.900 493.950 ;
        RECT 671.400 493.050 672.600 498.300 ;
        RECT 692.850 497.250 696.600 498.300 ;
        RECT 715.200 498.000 717.000 506.400 ;
        RECT 737.400 503.400 739.200 506.400 ;
        RECT 692.850 493.050 694.050 497.250 ;
        RECT 713.700 496.800 717.000 498.000 ;
        RECT 704.100 493.950 706.200 496.050 ;
        RECT 631.950 487.950 634.050 490.050 ;
        RECT 650.400 483.600 651.300 490.950 ;
        RECT 668.100 490.050 669.900 491.850 ;
        RECT 670.950 490.950 673.050 493.050 ;
        RECT 667.950 487.950 670.050 490.050 ;
        RECT 608.400 471.600 610.200 477.600 ;
        RECT 628.800 471.600 630.600 477.600 ;
        RECT 647.700 482.400 651.300 483.600 ;
        RECT 647.700 471.600 649.500 482.400 ;
        RECT 671.400 477.600 672.600 490.950 ;
        RECT 674.100 490.050 675.900 491.850 ;
        RECT 685.950 490.950 688.050 493.050 ;
        RECT 673.950 487.950 676.050 490.050 ;
        RECT 686.100 489.150 687.900 490.950 ;
        RECT 689.100 490.050 690.900 491.850 ;
        RECT 691.950 490.950 694.050 493.050 ;
        RECT 688.950 487.950 691.050 490.050 ;
        RECT 691.950 477.600 693.150 490.950 ;
        RECT 695.100 490.050 696.900 491.850 ;
        RECT 694.950 487.950 697.050 490.050 ;
        RECT 704.550 481.050 705.450 493.950 ;
        RECT 713.700 493.050 714.600 496.800 ;
        RECT 733.950 493.950 736.050 496.050 ;
        RECT 712.950 490.950 715.050 493.050 ;
        RECT 703.950 478.950 706.050 481.050 ;
        RECT 713.700 478.800 714.600 490.950 ;
        RECT 716.100 490.050 717.900 491.850 ;
        RECT 718.950 490.950 721.050 493.050 ;
        RECT 734.100 492.150 735.900 493.950 ;
        RECT 737.700 493.050 738.600 503.400 ;
        RECT 761.700 501.600 763.500 506.400 ;
        RECT 758.400 500.400 763.500 501.600 ;
        RECT 739.950 493.950 742.050 496.050 ;
        RECT 715.950 487.950 718.050 490.050 ;
        RECT 719.100 489.150 720.900 490.950 ;
        RECT 722.100 490.050 723.900 491.850 ;
        RECT 736.950 490.950 739.050 493.050 ;
        RECT 740.100 492.150 741.900 493.950 ;
        RECT 758.400 493.050 759.600 500.400 ;
        RECT 782.400 499.200 784.200 506.400 ;
        RECT 782.400 498.300 786.600 499.200 ;
        RECT 785.400 493.050 786.600 498.300 ;
        RECT 800.400 498.600 802.200 506.400 ;
        RECT 807.900 502.200 809.700 506.400 ;
        RECT 820.950 502.950 823.050 505.050 ;
        RECT 807.900 500.400 810.600 502.200 ;
        RECT 806.100 498.600 807.900 499.500 ;
        RECT 800.400 497.700 807.900 498.600 ;
        RECT 800.100 493.050 801.900 494.850 ;
        RECT 757.950 490.950 760.050 493.050 ;
        RECT 721.950 487.950 724.050 490.050 ;
        RECT 737.700 483.600 738.600 490.950 ;
        RECT 758.400 483.600 759.600 490.950 ;
        RECT 761.100 490.050 762.900 491.850 ;
        RECT 763.950 490.950 766.050 493.050 ;
        RECT 760.950 487.950 763.050 490.050 ;
        RECT 764.100 489.150 765.900 490.950 ;
        RECT 767.100 490.050 768.900 491.850 ;
        RECT 782.100 490.050 783.900 491.850 ;
        RECT 784.950 490.950 787.050 493.050 ;
        RECT 766.950 487.950 769.050 490.050 ;
        RECT 781.950 487.950 784.050 490.050 ;
        RECT 737.700 482.400 741.300 483.600 ;
        RECT 713.700 477.900 720.300 478.800 ;
        RECT 713.700 477.600 714.600 477.900 ;
        RECT 670.800 471.600 672.600 477.600 ;
        RECT 691.800 471.600 693.600 477.600 ;
        RECT 712.800 471.600 714.600 477.600 ;
        RECT 718.800 477.600 720.300 477.900 ;
        RECT 718.800 471.600 720.600 477.600 ;
        RECT 739.500 471.600 741.300 482.400 ;
        RECT 757.800 471.600 759.600 483.600 ;
        RECT 760.800 482.700 768.600 483.600 ;
        RECT 760.800 471.600 762.600 482.700 ;
        RECT 766.800 471.600 768.600 482.700 ;
        RECT 785.400 477.600 786.600 490.950 ;
        RECT 788.100 490.050 789.900 491.850 ;
        RECT 799.950 490.950 802.050 493.050 ;
        RECT 787.950 487.950 790.050 490.050 ;
        RECT 784.800 471.600 786.600 477.600 ;
        RECT 803.400 477.600 804.300 497.700 ;
        RECT 809.700 493.050 810.600 500.400 ;
        RECT 805.950 490.950 808.050 493.050 ;
        RECT 808.950 490.950 811.050 493.050 ;
        RECT 806.100 489.150 807.900 490.950 ;
        RECT 809.700 483.600 810.600 490.950 ;
        RECT 803.400 471.600 805.200 477.600 ;
        RECT 809.700 471.600 811.500 483.600 ;
        RECT 821.550 475.050 822.450 502.950 ;
        RECT 829.200 498.000 831.000 506.400 ;
        RECT 841.950 502.950 844.050 505.050 ;
        RECT 827.700 496.800 831.000 498.000 ;
        RECT 827.700 493.050 828.600 496.800 ;
        RECT 826.950 490.950 829.050 493.050 ;
        RECT 827.700 478.800 828.600 490.950 ;
        RECT 830.100 490.050 831.900 491.850 ;
        RECT 832.950 490.950 835.050 493.050 ;
        RECT 829.950 487.950 832.050 490.050 ;
        RECT 833.100 489.150 834.900 490.950 ;
        RECT 836.100 490.050 837.900 491.850 ;
        RECT 835.950 487.950 838.050 490.050 ;
        RECT 827.700 477.900 834.300 478.800 ;
        RECT 842.550 478.050 843.450 502.950 ;
        RECT 851.400 499.200 853.200 506.400 ;
        RECT 851.400 498.300 855.600 499.200 ;
        RECT 854.400 493.050 855.600 498.300 ;
        RECT 874.200 498.000 876.000 506.400 ;
        RECT 883.950 502.950 886.050 505.050 ;
        RECT 872.700 496.800 876.000 498.000 ;
        RECT 862.800 493.950 864.900 496.050 ;
        RECT 851.100 490.050 852.900 491.850 ;
        RECT 853.950 490.950 856.050 493.050 ;
        RECT 850.950 487.950 853.050 490.050 ;
        RECT 827.700 477.600 828.600 477.900 ;
        RECT 820.950 472.950 823.050 475.050 ;
        RECT 826.800 471.600 828.600 477.600 ;
        RECT 832.800 477.600 834.300 477.900 ;
        RECT 832.800 471.600 834.600 477.600 ;
        RECT 841.950 475.950 844.050 478.050 ;
        RECT 854.400 477.600 855.600 490.950 ;
        RECT 857.100 490.050 858.900 491.850 ;
        RECT 856.950 487.950 859.050 490.050 ;
        RECT 863.550 481.050 864.450 493.950 ;
        RECT 872.700 493.050 873.600 496.800 ;
        RECT 884.550 496.050 885.450 502.950 ;
        RECT 898.800 499.200 900.600 506.400 ;
        RECT 896.400 498.300 900.600 499.200 ;
        RECT 883.950 493.950 886.050 496.050 ;
        RECT 896.400 493.050 897.600 498.300 ;
        RECT 871.950 490.950 874.050 493.050 ;
        RECT 862.950 478.950 865.050 481.050 ;
        RECT 872.700 478.800 873.600 490.950 ;
        RECT 875.100 490.050 876.900 491.850 ;
        RECT 877.950 490.950 880.050 493.050 ;
        RECT 874.950 487.950 877.050 490.050 ;
        RECT 878.100 489.150 879.900 490.950 ;
        RECT 881.100 490.050 882.900 491.850 ;
        RECT 893.100 490.050 894.900 491.850 ;
        RECT 895.950 490.950 898.050 493.050 ;
        RECT 880.950 487.950 883.050 490.050 ;
        RECT 892.950 487.950 895.050 490.050 ;
        RECT 872.700 477.900 879.300 478.800 ;
        RECT 872.700 477.600 873.600 477.900 ;
        RECT 853.800 471.600 855.600 477.600 ;
        RECT 871.800 471.600 873.600 477.600 ;
        RECT 877.800 477.600 879.300 477.900 ;
        RECT 896.400 477.600 897.600 490.950 ;
        RECT 899.100 490.050 900.900 491.850 ;
        RECT 898.950 487.950 901.050 490.050 ;
        RECT 877.800 471.600 879.600 477.600 ;
        RECT 896.400 471.600 898.200 477.600 ;
        RECT 19.800 455.400 23.100 467.400 ;
        RECT 41.400 461.400 43.200 467.400 ;
        RECT 64.800 461.400 66.600 467.400 ;
        RECT 85.800 461.400 87.600 467.400 ;
        RECT 107.400 461.400 109.200 467.400 ;
        RECT 14.100 448.050 15.900 449.850 ;
        RECT 16.950 448.950 19.050 451.050 ;
        RECT 13.950 445.950 16.050 448.050 ;
        RECT 17.100 447.150 18.900 448.950 ;
        RECT 20.700 448.050 21.900 455.400 ;
        RECT 31.950 454.950 34.050 457.050 ;
        RECT 22.950 448.950 25.050 451.050 ;
        RECT 19.950 445.950 22.050 448.050 ;
        RECT 23.100 447.150 24.900 448.950 ;
        RECT 26.100 448.050 27.900 449.850 ;
        RECT 25.950 445.950 28.050 448.050 ;
        RECT 20.700 441.300 22.050 445.950 ;
        RECT 32.550 445.050 33.450 454.950 ;
        RECT 37.950 448.950 40.050 451.050 ;
        RECT 38.100 447.150 39.900 448.950 ;
        RECT 41.400 448.050 42.600 461.400 ;
        RECT 43.950 448.950 46.050 451.050 ;
        RECT 61.950 448.950 64.050 451.050 ;
        RECT 40.950 445.950 43.050 448.050 ;
        RECT 44.100 447.150 45.900 448.950 ;
        RECT 62.100 447.150 63.900 448.950 ;
        RECT 65.400 448.050 66.600 461.400 ;
        RECT 67.950 448.950 70.050 451.050 ;
        RECT 82.950 448.950 85.050 451.050 ;
        RECT 64.950 445.950 67.050 448.050 ;
        RECT 68.100 447.150 69.900 448.950 ;
        RECT 83.100 447.150 84.900 448.950 ;
        RECT 86.400 448.050 87.600 461.400 ;
        RECT 88.950 448.950 91.050 451.050 ;
        RECT 103.950 448.950 106.050 451.050 ;
        RECT 85.950 445.950 88.050 448.050 ;
        RECT 89.100 447.150 90.900 448.950 ;
        RECT 104.100 447.150 105.900 448.950 ;
        RECT 107.850 448.050 109.050 461.400 ;
        RECT 128.700 456.600 130.500 467.400 ;
        RECT 149.400 461.400 151.200 467.400 ;
        RECT 169.800 461.400 171.600 467.400 ;
        RECT 190.800 461.400 192.600 467.400 ;
        RECT 128.700 455.400 132.300 456.600 ;
        RECT 109.950 448.950 112.050 451.050 ;
        RECT 106.950 445.950 109.050 448.050 ;
        RECT 110.100 447.150 111.900 448.950 ;
        RECT 113.100 448.050 114.900 449.850 ;
        RECT 131.400 448.050 132.300 455.400 ;
        RECT 149.400 454.050 150.600 461.400 ;
        RECT 146.100 448.050 147.900 449.850 ;
        RECT 148.950 448.950 151.050 454.050 ;
        RECT 112.950 445.950 115.050 448.050 ;
        RECT 31.950 442.950 34.050 445.050 ;
        RECT 17.400 440.100 22.050 441.300 ;
        RECT 41.400 440.700 42.600 445.950 ;
        RECT 65.400 440.700 66.600 445.950 ;
        RECT 86.400 440.700 87.600 445.950 ;
        RECT 106.950 441.750 108.150 445.950 ;
        RECT 128.100 445.050 129.900 446.850 ;
        RECT 130.950 445.950 133.050 448.050 ;
        RECT 127.950 442.950 130.050 445.050 ;
        RECT 17.400 438.600 18.300 440.100 ;
        RECT 41.400 439.800 45.600 440.700 ;
        RECT 13.800 433.500 15.600 438.600 ;
        RECT 16.800 434.400 18.600 438.600 ;
        RECT 19.800 438.000 27.600 438.900 ;
        RECT 19.800 433.500 21.600 438.000 ;
        RECT 13.800 432.600 21.600 433.500 ;
        RECT 25.800 432.600 27.600 438.000 ;
        RECT 43.800 432.600 45.600 439.800 ;
        RECT 62.400 439.800 66.600 440.700 ;
        RECT 83.400 439.800 87.600 440.700 ;
        RECT 104.400 440.700 108.150 441.750 ;
        RECT 62.400 432.600 64.200 439.800 ;
        RECT 83.400 432.600 85.200 439.800 ;
        RECT 104.400 438.600 105.600 440.700 ;
        RECT 103.800 432.600 105.600 438.600 ;
        RECT 106.800 437.700 114.600 439.050 ;
        RECT 106.800 432.600 108.600 437.700 ;
        RECT 112.800 432.600 114.600 437.700 ;
        RECT 131.400 435.600 132.300 445.950 ;
        RECT 134.100 445.050 135.900 446.850 ;
        RECT 145.950 445.950 148.050 448.050 ;
        RECT 133.950 442.950 136.050 445.050 ;
        RECT 149.400 435.600 150.600 448.950 ;
        RECT 164.100 448.050 165.900 449.850 ;
        RECT 166.950 448.950 169.050 451.050 ;
        RECT 163.950 445.950 166.050 448.050 ;
        RECT 167.100 447.150 168.900 448.950 ;
        RECT 169.950 448.050 171.150 461.400 ;
        RECT 191.700 461.100 192.600 461.400 ;
        RECT 196.800 461.400 198.600 467.400 ;
        RECT 218.400 461.400 220.200 467.400 ;
        RECT 196.800 461.100 198.300 461.400 ;
        RECT 191.700 460.200 198.300 461.100 ;
        RECT 172.950 448.950 175.050 451.050 ;
        RECT 169.950 445.950 172.050 448.050 ;
        RECT 173.100 447.150 174.900 448.950 ;
        RECT 191.700 448.050 192.600 460.200 ;
        RECT 193.950 448.950 196.050 451.050 ;
        RECT 190.950 445.950 193.050 448.050 ;
        RECT 194.100 447.150 195.900 448.950 ;
        RECT 197.100 448.050 198.900 449.850 ;
        RECT 199.950 448.950 202.050 451.050 ;
        RECT 214.950 448.950 217.050 451.050 ;
        RECT 196.950 445.950 199.050 448.050 ;
        RECT 200.100 447.150 201.900 448.950 ;
        RECT 215.100 447.150 216.900 448.950 ;
        RECT 218.850 448.050 220.050 461.400 ;
        RECT 238.500 455.400 240.300 467.400 ;
        RECT 244.800 461.400 246.600 467.400 ;
        RECT 220.950 448.950 223.050 451.050 ;
        RECT 217.950 445.950 220.050 448.050 ;
        RECT 221.100 447.150 222.900 448.950 ;
        RECT 224.100 448.050 225.900 449.850 ;
        RECT 238.500 448.050 239.700 455.400 ;
        RECT 245.400 454.500 246.600 461.400 ;
        RECT 261.900 455.400 265.200 467.400 ;
        RECT 289.500 456.600 291.300 467.400 ;
        RECT 310.800 461.400 312.600 467.400 ;
        RECT 331.800 461.400 333.600 467.400 ;
        RECT 356.400 461.400 358.200 467.400 ;
        RECT 377.400 461.400 379.200 467.400 ;
        RECT 287.700 455.400 291.300 456.600 ;
        RECT 240.600 453.600 246.600 454.500 ;
        RECT 240.600 452.700 242.850 453.600 ;
        RECT 223.950 445.950 226.050 448.050 ;
        RECT 238.500 445.950 241.050 448.050 ;
        RECT 170.850 441.750 172.050 445.950 ;
        RECT 191.700 442.200 192.600 445.950 ;
        RECT 170.850 440.700 174.600 441.750 ;
        RECT 191.700 441.000 195.000 442.200 ;
        RECT 217.950 441.750 219.150 445.950 ;
        RECT 164.400 437.700 172.200 439.050 ;
        RECT 130.800 432.600 132.600 435.600 ;
        RECT 149.400 432.600 151.200 435.600 ;
        RECT 164.400 432.600 166.200 437.700 ;
        RECT 170.400 432.600 172.200 437.700 ;
        RECT 173.400 438.600 174.600 440.700 ;
        RECT 173.400 432.600 175.200 438.600 ;
        RECT 193.200 432.600 195.000 441.000 ;
        RECT 215.400 440.700 219.150 441.750 ;
        RECT 215.400 438.600 216.600 440.700 ;
        RECT 214.800 432.600 216.600 438.600 ;
        RECT 217.800 437.700 225.600 439.050 ;
        RECT 217.800 432.600 219.600 437.700 ;
        RECT 223.800 432.600 225.600 437.700 ;
        RECT 238.500 438.600 239.700 445.950 ;
        RECT 241.950 441.300 242.850 452.700 ;
        RECT 245.100 448.050 246.900 449.850 ;
        RECT 257.100 448.050 258.900 449.850 ;
        RECT 259.950 448.950 262.050 451.050 ;
        RECT 244.950 445.950 247.050 448.050 ;
        RECT 256.950 445.950 259.050 448.050 ;
        RECT 260.100 447.150 261.900 448.950 ;
        RECT 263.100 448.050 264.300 455.400 ;
        RECT 265.950 448.950 268.050 451.050 ;
        RECT 262.950 445.950 265.050 448.050 ;
        RECT 266.100 447.150 267.900 448.950 ;
        RECT 269.100 448.050 270.900 449.850 ;
        RECT 287.700 448.050 288.600 455.400 ;
        RECT 307.950 448.950 310.050 451.050 ;
        RECT 268.950 445.950 271.050 448.050 ;
        RECT 240.600 440.400 242.850 441.300 ;
        RECT 262.950 441.300 264.300 445.950 ;
        RECT 284.100 445.050 285.900 446.850 ;
        RECT 286.950 445.950 289.050 448.050 ;
        RECT 308.100 447.150 309.900 448.950 ;
        RECT 311.400 448.050 312.600 461.400 ;
        RECT 313.950 448.950 316.050 451.050 ;
        RECT 283.950 442.950 286.050 445.050 ;
        RECT 240.600 439.500 246.600 440.400 ;
        RECT 262.950 440.100 267.600 441.300 ;
        RECT 238.500 432.600 240.300 438.600 ;
        RECT 245.400 435.600 246.600 439.500 ;
        RECT 244.800 432.600 246.600 435.600 ;
        RECT 257.400 438.000 265.200 438.900 ;
        RECT 266.700 438.600 267.600 440.100 ;
        RECT 257.400 432.600 259.200 438.000 ;
        RECT 263.400 433.500 265.200 438.000 ;
        RECT 266.400 434.400 268.200 438.600 ;
        RECT 269.400 433.500 271.200 438.600 ;
        RECT 287.700 435.600 288.600 445.950 ;
        RECT 290.100 445.050 291.900 446.850 ;
        RECT 310.950 445.950 313.050 448.050 ;
        RECT 314.100 447.150 315.900 448.950 ;
        RECT 326.100 448.050 327.900 449.850 ;
        RECT 328.950 448.950 331.050 451.050 ;
        RECT 325.950 445.950 328.050 448.050 ;
        RECT 329.100 447.150 330.900 448.950 ;
        RECT 331.950 448.050 333.150 461.400 ;
        RECT 334.950 448.950 337.050 451.050 ;
        RECT 352.950 448.950 355.050 451.050 ;
        RECT 331.950 445.950 334.050 448.050 ;
        RECT 335.100 447.150 336.900 448.950 ;
        RECT 353.100 447.150 354.900 448.950 ;
        RECT 356.850 448.050 358.050 461.400 ;
        RECT 377.400 454.050 378.600 461.400 ;
        RECT 385.950 460.950 388.050 463.050 ;
        RECT 397.800 461.400 399.600 467.400 ;
        RECT 358.950 448.950 361.050 451.050 ;
        RECT 289.950 442.950 292.050 445.050 ;
        RECT 311.400 440.700 312.600 445.950 ;
        RECT 332.850 441.750 334.050 445.950 ;
        RECT 355.950 445.950 358.050 448.050 ;
        RECT 359.100 447.150 360.900 448.950 ;
        RECT 362.100 448.050 363.900 449.850 ;
        RECT 374.100 448.050 375.900 449.850 ;
        RECT 376.950 448.950 379.050 454.050 ;
        RECT 361.950 445.950 364.050 448.050 ;
        RECT 373.950 445.950 376.050 448.050 ;
        RECT 355.950 441.750 357.150 445.950 ;
        RECT 332.850 440.700 336.600 441.750 ;
        RECT 308.400 439.800 312.600 440.700 ;
        RECT 263.400 432.600 271.200 433.500 ;
        RECT 287.400 432.600 289.200 435.600 ;
        RECT 308.400 432.600 310.200 439.800 ;
        RECT 326.400 437.700 334.200 439.050 ;
        RECT 326.400 432.600 328.200 437.700 ;
        RECT 332.400 432.600 334.200 437.700 ;
        RECT 335.400 438.600 336.600 440.700 ;
        RECT 353.400 440.700 357.150 441.750 ;
        RECT 353.400 438.600 354.600 440.700 ;
        RECT 335.400 432.600 337.200 438.600 ;
        RECT 352.800 432.600 354.600 438.600 ;
        RECT 355.800 437.700 363.600 439.050 ;
        RECT 355.800 432.600 357.600 437.700 ;
        RECT 361.800 432.600 363.600 437.700 ;
        RECT 377.400 435.600 378.600 448.950 ;
        RECT 386.550 439.050 387.450 460.950 ;
        RECT 392.100 448.050 393.900 449.850 ;
        RECT 394.950 448.950 397.050 451.050 ;
        RECT 391.950 445.950 394.050 448.050 ;
        RECT 395.100 447.150 396.900 448.950 ;
        RECT 397.950 448.050 399.150 461.400 ;
        RECT 415.800 455.400 417.600 467.400 ;
        RECT 418.800 456.300 420.600 467.400 ;
        RECT 424.800 456.300 426.600 467.400 ;
        RECT 430.950 460.950 433.050 463.050 ;
        RECT 440.400 461.400 442.200 467.400 ;
        RECT 440.700 461.100 442.200 461.400 ;
        RECT 446.400 461.400 448.200 467.400 ;
        RECT 466.800 461.400 468.600 467.400 ;
        RECT 446.400 461.100 447.300 461.400 ;
        RECT 418.800 455.400 426.600 456.300 ;
        RECT 400.950 448.950 403.050 451.050 ;
        RECT 397.950 445.950 400.050 448.050 ;
        RECT 401.100 447.150 402.900 448.950 ;
        RECT 416.400 448.050 417.600 455.400 ;
        RECT 418.950 448.950 421.050 451.050 ;
        RECT 415.950 445.950 418.050 448.050 ;
        RECT 419.100 447.150 420.900 448.950 ;
        RECT 422.100 448.050 423.900 449.850 ;
        RECT 424.950 448.950 427.050 451.050 ;
        RECT 421.950 445.950 424.050 448.050 ;
        RECT 425.100 447.150 426.900 448.950 ;
        RECT 398.850 441.750 400.050 445.950 ;
        RECT 398.850 440.700 402.600 441.750 ;
        RECT 385.950 436.950 388.050 439.050 ;
        RECT 392.400 437.700 400.200 439.050 ;
        RECT 377.400 432.600 379.200 435.600 ;
        RECT 392.400 432.600 394.200 437.700 ;
        RECT 398.400 432.600 400.200 437.700 ;
        RECT 401.400 438.600 402.600 440.700 ;
        RECT 416.400 438.600 417.600 445.950 ;
        RECT 431.550 439.050 432.450 460.950 ;
        RECT 440.700 460.200 447.300 461.100 ;
        RECT 436.950 448.950 439.050 451.050 ;
        RECT 437.100 447.150 438.900 448.950 ;
        RECT 440.100 448.050 441.900 449.850 ;
        RECT 442.950 448.950 445.050 451.050 ;
        RECT 439.950 445.950 442.050 448.050 ;
        RECT 443.100 447.150 444.900 448.950 ;
        RECT 446.400 448.050 447.300 460.200 ;
        RECT 463.950 448.950 466.050 451.050 ;
        RECT 445.950 445.950 448.050 448.050 ;
        RECT 464.100 447.150 465.900 448.950 ;
        RECT 467.400 448.050 468.600 461.400 ;
        RECT 485.400 461.400 487.200 467.400 ;
        RECT 506.400 461.400 508.200 467.400 ;
        RECT 475.950 457.950 478.050 460.050 ;
        RECT 469.950 448.950 472.050 451.050 ;
        RECT 466.950 445.950 469.050 448.050 ;
        RECT 470.100 447.150 471.900 448.950 ;
        RECT 446.400 442.200 447.300 445.950 ;
        RECT 444.000 441.000 447.300 442.200 ;
        RECT 401.400 432.600 403.200 438.600 ;
        RECT 416.400 437.400 421.500 438.600 ;
        RECT 419.700 432.600 421.500 437.400 ;
        RECT 431.100 436.950 433.200 439.050 ;
        RECT 444.000 432.600 445.800 441.000 ;
        RECT 467.400 440.700 468.600 445.950 ;
        RECT 476.550 445.050 477.450 457.950 ;
        RECT 481.950 448.950 484.050 451.050 ;
        RECT 482.100 447.150 483.900 448.950 ;
        RECT 485.400 448.050 486.600 461.400 ;
        RECT 487.950 448.950 490.050 451.050 ;
        RECT 502.950 448.950 505.050 451.050 ;
        RECT 484.950 445.950 487.050 448.050 ;
        RECT 488.100 447.150 489.900 448.950 ;
        RECT 503.100 447.150 504.900 448.950 ;
        RECT 506.400 448.050 507.600 461.400 ;
        RECT 524.400 456.300 526.200 467.400 ;
        RECT 530.400 456.300 532.200 467.400 ;
        RECT 524.400 455.400 532.200 456.300 ;
        RECT 533.400 455.400 535.200 467.400 ;
        RECT 553.800 461.400 555.600 467.400 ;
        RECT 574.800 461.400 576.600 467.400 ;
        RECT 598.800 461.400 600.600 467.400 ;
        RECT 620.400 461.400 622.200 467.400 ;
        RECT 508.950 448.950 511.050 451.050 ;
        RECT 523.950 448.950 526.050 451.050 ;
        RECT 505.950 445.950 508.050 448.050 ;
        RECT 509.100 447.150 510.900 448.950 ;
        RECT 524.100 447.150 525.900 448.950 ;
        RECT 527.100 448.050 528.900 449.850 ;
        RECT 529.950 448.950 532.050 451.050 ;
        RECT 526.950 445.950 529.050 448.050 ;
        RECT 530.100 447.150 531.900 448.950 ;
        RECT 533.400 448.050 534.600 455.400 ;
        RECT 550.950 448.950 553.050 451.050 ;
        RECT 532.950 445.950 535.050 448.050 ;
        RECT 551.100 447.150 552.900 448.950 ;
        RECT 554.400 448.050 555.600 461.400 ;
        RECT 556.950 448.950 559.050 451.050 ;
        RECT 553.950 445.950 556.050 448.050 ;
        RECT 557.100 447.150 558.900 448.950 ;
        RECT 569.100 448.050 570.900 449.850 ;
        RECT 571.950 448.950 574.050 451.050 ;
        RECT 568.950 445.950 571.050 448.050 ;
        RECT 572.100 447.150 573.900 448.950 ;
        RECT 574.950 448.050 576.150 461.400 ;
        RECT 577.950 448.950 580.050 451.050 ;
        RECT 574.950 445.950 577.050 448.050 ;
        RECT 578.100 447.150 579.900 448.950 ;
        RECT 593.100 448.050 594.900 449.850 ;
        RECT 595.950 448.950 598.050 451.050 ;
        RECT 592.950 445.950 595.050 448.050 ;
        RECT 596.100 447.150 597.900 448.950 ;
        RECT 598.950 448.050 600.150 461.400 ;
        RECT 620.400 454.050 621.600 461.400 ;
        RECT 637.800 455.400 639.600 467.400 ;
        RECT 640.800 456.300 642.600 467.400 ;
        RECT 646.800 456.300 648.600 467.400 ;
        RECT 662.400 461.400 664.200 467.400 ;
        RECT 662.700 461.100 664.200 461.400 ;
        RECT 668.400 461.400 670.200 467.400 ;
        RECT 668.400 461.100 669.300 461.400 ;
        RECT 662.700 460.200 669.300 461.100 ;
        RECT 640.800 455.400 648.600 456.300 ;
        RECT 601.950 448.950 604.050 451.050 ;
        RECT 598.950 445.950 601.050 448.050 ;
        RECT 602.100 447.150 603.900 448.950 ;
        RECT 617.100 448.050 618.900 449.850 ;
        RECT 619.950 448.950 622.050 454.050 ;
        RECT 616.950 445.950 619.050 448.050 ;
        RECT 475.800 442.950 477.900 445.050 ;
        RECT 464.400 439.800 468.600 440.700 ;
        RECT 485.400 440.700 486.600 445.950 ;
        RECT 506.400 440.700 507.600 445.950 ;
        RECT 485.400 439.800 489.600 440.700 ;
        RECT 506.400 439.800 510.600 440.700 ;
        RECT 464.400 432.600 466.200 439.800 ;
        RECT 487.800 432.600 489.600 439.800 ;
        RECT 508.800 432.600 510.600 439.800 ;
        RECT 533.400 438.600 534.600 445.950 ;
        RECT 554.400 440.700 555.600 445.950 ;
        RECT 575.850 441.750 577.050 445.950 ;
        RECT 599.850 441.750 601.050 445.950 ;
        RECT 575.850 440.700 579.600 441.750 ;
        RECT 599.850 440.700 603.600 441.750 ;
        RECT 529.500 437.400 534.600 438.600 ;
        RECT 551.400 439.800 555.600 440.700 ;
        RECT 529.500 432.600 531.300 437.400 ;
        RECT 551.400 432.600 553.200 439.800 ;
        RECT 569.400 437.700 577.200 439.050 ;
        RECT 569.400 432.600 571.200 437.700 ;
        RECT 575.400 432.600 577.200 437.700 ;
        RECT 578.400 438.600 579.600 440.700 ;
        RECT 578.400 432.600 580.200 438.600 ;
        RECT 593.400 437.700 601.200 439.050 ;
        RECT 593.400 432.600 595.200 437.700 ;
        RECT 599.400 432.600 601.200 437.700 ;
        RECT 602.400 438.600 603.600 440.700 ;
        RECT 602.400 432.600 604.200 438.600 ;
        RECT 620.400 435.600 621.600 448.950 ;
        RECT 638.400 448.050 639.600 455.400 ;
        RECT 640.950 448.950 643.050 451.050 ;
        RECT 637.950 445.950 640.050 448.050 ;
        RECT 641.100 447.150 642.900 448.950 ;
        RECT 644.100 448.050 645.900 449.850 ;
        RECT 646.950 448.950 649.050 451.050 ;
        RECT 658.950 448.950 661.050 451.050 ;
        RECT 643.950 445.950 646.050 448.050 ;
        RECT 647.100 447.150 648.900 448.950 ;
        RECT 659.100 447.150 660.900 448.950 ;
        RECT 662.100 448.050 663.900 449.850 ;
        RECT 664.950 448.950 667.050 451.050 ;
        RECT 661.950 445.950 664.050 448.050 ;
        RECT 665.100 447.150 666.900 448.950 ;
        RECT 668.400 448.050 669.300 460.200 ;
        RECT 685.500 455.400 687.300 467.400 ;
        RECT 691.800 461.400 693.600 467.400 ;
        RECT 685.500 448.050 686.700 455.400 ;
        RECT 692.400 454.500 693.600 461.400 ;
        RECT 687.600 453.600 693.600 454.500 ;
        RECT 707.400 461.400 709.200 467.400 ;
        RECT 724.800 461.400 726.600 467.400 ;
        RECT 707.400 454.050 708.600 461.400 ;
        RECT 725.700 461.100 726.600 461.400 ;
        RECT 730.800 461.400 732.600 467.400 ;
        RECT 749.400 461.400 751.200 467.400 ;
        RECT 773.400 461.400 775.200 467.400 ;
        RECT 794.400 461.400 796.200 467.400 ;
        RECT 802.950 463.950 805.050 466.050 ;
        RECT 730.800 461.100 732.300 461.400 ;
        RECT 725.700 460.200 732.300 461.100 ;
        RECT 687.600 452.700 689.850 453.600 ;
        RECT 667.950 445.950 670.050 448.050 ;
        RECT 685.500 445.950 688.050 448.050 ;
        RECT 638.400 438.600 639.600 445.950 ;
        RECT 668.400 442.200 669.300 445.950 ;
        RECT 666.000 441.000 669.300 442.200 ;
        RECT 638.400 437.400 643.500 438.600 ;
        RECT 620.400 432.600 622.200 435.600 ;
        RECT 641.700 432.600 643.500 437.400 ;
        RECT 666.000 432.600 667.800 441.000 ;
        RECT 685.500 438.600 686.700 445.950 ;
        RECT 688.950 441.300 689.850 452.700 ;
        RECT 692.100 448.050 693.900 449.850 ;
        RECT 704.100 448.050 705.900 449.850 ;
        RECT 706.950 448.950 709.050 454.050 ;
        RECT 691.950 445.950 694.050 448.050 ;
        RECT 703.950 445.950 706.050 448.050 ;
        RECT 687.600 440.400 689.850 441.300 ;
        RECT 687.600 439.500 693.600 440.400 ;
        RECT 685.500 432.600 687.300 438.600 ;
        RECT 692.400 435.600 693.600 439.500 ;
        RECT 691.800 432.600 693.600 435.600 ;
        RECT 707.400 435.600 708.600 448.950 ;
        RECT 725.700 448.050 726.600 460.200 ;
        RECT 727.950 448.950 730.050 451.050 ;
        RECT 724.950 445.950 727.050 448.050 ;
        RECT 728.100 447.150 729.900 448.950 ;
        RECT 731.100 448.050 732.900 449.850 ;
        RECT 733.950 448.950 736.050 451.050 ;
        RECT 745.950 448.950 748.050 451.050 ;
        RECT 730.950 445.950 733.050 448.050 ;
        RECT 734.100 447.150 735.900 448.950 ;
        RECT 746.100 447.150 747.900 448.950 ;
        RECT 749.400 448.050 750.600 461.400 ;
        RECT 751.950 448.950 754.050 451.050 ;
        RECT 769.950 448.950 772.050 451.050 ;
        RECT 748.950 445.950 751.050 448.050 ;
        RECT 752.100 447.150 753.900 448.950 ;
        RECT 770.100 447.150 771.900 448.950 ;
        RECT 773.850 448.050 775.050 461.400 ;
        RECT 794.400 454.050 795.600 461.400 ;
        RECT 775.950 448.950 778.050 451.050 ;
        RECT 772.950 445.950 775.050 448.050 ;
        RECT 776.100 447.150 777.900 448.950 ;
        RECT 779.100 448.050 780.900 449.850 ;
        RECT 791.100 448.050 792.900 449.850 ;
        RECT 793.950 448.950 796.050 454.050 ;
        RECT 799.950 451.950 802.050 454.050 ;
        RECT 778.950 445.950 781.050 448.050 ;
        RECT 790.950 445.950 793.050 448.050 ;
        RECT 725.700 442.200 726.600 445.950 ;
        RECT 725.700 441.000 729.000 442.200 ;
        RECT 707.400 432.600 709.200 435.600 ;
        RECT 727.200 432.600 729.000 441.000 ;
        RECT 749.400 440.700 750.600 445.950 ;
        RECT 772.950 441.750 774.150 445.950 ;
        RECT 770.400 440.700 774.150 441.750 ;
        RECT 749.400 439.800 753.600 440.700 ;
        RECT 751.800 432.600 753.600 439.800 ;
        RECT 770.400 438.600 771.600 440.700 ;
        RECT 769.800 432.600 771.600 438.600 ;
        RECT 772.800 437.700 780.600 439.050 ;
        RECT 772.800 432.600 774.600 437.700 ;
        RECT 778.800 432.600 780.600 437.700 ;
        RECT 794.400 435.600 795.600 448.950 ;
        RECT 800.550 439.050 801.450 451.950 ;
        RECT 799.800 436.950 801.900 439.050 ;
        RECT 803.550 436.050 804.450 463.950 ;
        RECT 811.800 461.400 813.600 467.400 ;
        RECT 812.700 461.100 813.600 461.400 ;
        RECT 817.800 461.400 819.600 467.400 ;
        RECT 836.400 461.400 838.200 467.400 ;
        RECT 854.400 461.400 856.200 467.400 ;
        RECT 817.800 461.100 819.300 461.400 ;
        RECT 812.700 460.200 819.300 461.100 ;
        RECT 812.700 448.050 813.600 460.200 ;
        RECT 836.400 454.050 837.600 461.400 ;
        RECT 814.950 448.950 817.050 451.050 ;
        RECT 811.950 445.950 814.050 448.050 ;
        RECT 815.100 447.150 816.900 448.950 ;
        RECT 818.100 448.050 819.900 449.850 ;
        RECT 820.950 448.950 823.050 451.050 ;
        RECT 817.950 445.950 820.050 448.050 ;
        RECT 821.100 447.150 822.900 448.950 ;
        RECT 833.100 448.050 834.900 449.850 ;
        RECT 835.950 448.950 838.050 454.050 ;
        RECT 850.950 448.950 853.050 451.050 ;
        RECT 832.950 445.950 835.050 448.050 ;
        RECT 812.700 442.200 813.600 445.950 ;
        RECT 812.700 441.000 816.000 442.200 ;
        RECT 794.400 432.600 796.200 435.600 ;
        RECT 803.100 433.950 805.200 436.050 ;
        RECT 814.200 432.600 816.000 441.000 ;
        RECT 836.400 435.600 837.600 448.950 ;
        RECT 851.100 447.150 852.900 448.950 ;
        RECT 854.400 448.050 855.600 461.400 ;
        RECT 872.400 455.400 874.200 467.400 ;
        RECT 879.900 456.900 881.700 467.400 ;
        RECT 899.400 461.400 901.200 467.400 ;
        RECT 879.900 455.400 882.300 456.900 ;
        RECT 872.400 453.900 873.600 455.400 ;
        RECT 872.400 452.700 879.600 453.900 ;
        RECT 877.800 452.100 879.600 452.700 ;
        RECT 856.950 448.950 859.050 451.050 ;
        RECT 871.950 448.950 874.050 451.050 ;
        RECT 853.950 445.950 856.050 448.050 ;
        RECT 857.100 447.150 858.900 448.950 ;
        RECT 872.100 447.150 873.900 448.950 ;
        RECT 875.100 448.050 876.900 449.850 ;
        RECT 874.950 445.950 877.050 448.050 ;
        RECT 854.400 440.700 855.600 445.950 ;
        RECT 878.700 441.600 879.600 452.100 ;
        RECT 880.950 448.050 882.300 455.400 ;
        RECT 895.950 448.950 898.050 451.050 ;
        RECT 880.950 445.950 883.050 448.050 ;
        RECT 896.100 447.150 897.900 448.950 ;
        RECT 899.400 448.050 900.600 461.400 ;
        RECT 901.950 448.950 904.050 451.050 ;
        RECT 898.950 445.950 901.050 448.050 ;
        RECT 902.100 447.150 903.900 448.950 ;
        RECT 877.800 440.700 879.600 441.600 ;
        RECT 854.400 439.800 858.600 440.700 ;
        RECT 836.400 432.600 838.200 435.600 ;
        RECT 856.800 432.600 858.600 439.800 ;
        RECT 876.300 439.800 879.600 440.700 ;
        RECT 876.300 435.600 877.200 439.800 ;
        RECT 882.000 438.600 883.050 445.950 ;
        RECT 892.950 442.950 895.050 445.050 ;
        RECT 875.400 432.600 877.200 435.600 ;
        RECT 881.400 432.600 883.200 438.600 ;
        RECT 893.550 436.050 894.450 442.950 ;
        RECT 899.400 440.700 900.600 445.950 ;
        RECT 899.400 439.800 903.600 440.700 ;
        RECT 892.950 433.950 895.050 436.050 ;
        RECT 901.800 432.600 903.600 439.800 ;
        RECT 3.150 422.400 4.950 428.400 ;
        RECT 10.950 426.300 12.750 428.400 ;
        RECT 9.000 425.400 12.750 426.300 ;
        RECT 18.750 425.400 20.550 428.400 ;
        RECT 26.550 425.400 28.350 428.400 ;
        RECT 9.000 424.500 10.050 425.400 ;
        RECT 18.750 424.500 19.800 425.400 ;
        RECT 7.950 422.400 10.050 424.500 ;
        RECT 3.150 407.700 4.050 422.400 ;
        RECT 11.550 421.800 13.350 423.600 ;
        RECT 14.850 423.450 19.800 424.500 ;
        RECT 27.300 424.500 28.350 425.400 ;
        RECT 14.850 422.700 16.650 423.450 ;
        RECT 27.300 423.300 31.050 424.500 ;
        RECT 28.950 422.400 31.050 423.300 ;
        RECT 34.650 422.400 36.450 428.400 ;
        RECT 49.800 427.500 57.600 428.400 ;
        RECT 11.850 420.000 12.900 421.800 ;
        RECT 22.050 420.000 23.850 420.600 ;
        RECT 11.850 418.800 23.850 420.000 ;
        RECT 6.000 417.600 12.900 418.800 ;
        RECT 6.000 416.850 6.900 417.600 ;
        RECT 11.100 417.000 12.900 417.600 ;
        RECT 5.100 415.050 6.900 416.850 ;
        RECT 8.100 415.800 9.900 416.400 ;
        RECT 4.950 412.950 7.050 415.050 ;
        RECT 8.100 414.600 16.050 415.800 ;
        RECT 13.950 412.950 16.050 414.600 ;
        RECT 12.450 407.700 14.250 408.000 ;
        RECT 3.150 407.100 14.250 407.700 ;
        RECT 3.150 406.500 20.850 407.100 ;
        RECT 3.150 405.600 4.050 406.500 ;
        RECT 12.450 406.200 20.850 406.500 ;
        RECT 3.150 393.600 4.950 405.600 ;
        RECT 17.250 404.700 19.050 405.300 ;
        RECT 11.550 403.500 19.050 404.700 ;
        RECT 19.950 404.100 20.850 406.200 ;
        RECT 22.950 406.200 23.850 418.800 ;
        RECT 35.250 415.050 36.450 422.400 ;
        RECT 43.950 421.950 46.050 424.050 ;
        RECT 49.800 422.400 51.600 427.500 ;
        RECT 52.800 422.400 54.600 426.600 ;
        RECT 55.800 423.000 57.600 427.500 ;
        RECT 61.800 423.000 63.600 428.400 ;
        RECT 30.150 413.250 36.450 415.050 ;
        RECT 31.950 412.950 36.450 413.250 ;
        RECT 32.250 407.400 34.050 409.200 ;
        RECT 28.950 406.200 33.150 407.400 ;
        RECT 22.950 405.300 28.050 406.200 ;
        RECT 28.950 405.300 31.050 406.200 ;
        RECT 35.250 405.600 36.450 412.950 ;
        RECT 27.150 404.400 28.050 405.300 ;
        RECT 24.450 404.100 26.250 404.400 ;
        RECT 11.550 402.600 12.750 403.500 ;
        RECT 19.950 403.200 26.250 404.100 ;
        RECT 24.450 402.600 26.250 403.200 ;
        RECT 27.150 402.600 29.850 404.400 ;
        RECT 7.950 400.500 12.750 402.600 ;
        RECT 15.450 401.550 17.250 402.300 ;
        RECT 20.250 401.550 22.050 402.300 ;
        RECT 15.450 400.500 22.050 401.550 ;
        RECT 11.550 399.600 12.750 400.500 ;
        RECT 11.550 393.600 13.350 399.600 ;
        RECT 19.350 393.600 21.150 400.500 ;
        RECT 27.150 399.600 31.050 401.700 ;
        RECT 27.150 393.600 28.950 399.600 ;
        RECT 34.650 393.600 36.450 405.600 ;
        RECT 44.550 403.050 45.450 421.950 ;
        RECT 53.400 420.900 54.300 422.400 ;
        RECT 55.800 422.100 63.600 423.000 ;
        RECT 66.150 422.400 67.950 428.400 ;
        RECT 73.950 426.300 75.750 428.400 ;
        RECT 72.000 425.400 75.750 426.300 ;
        RECT 81.750 425.400 83.550 428.400 ;
        RECT 89.550 425.400 91.350 428.400 ;
        RECT 72.000 424.500 73.050 425.400 ;
        RECT 81.750 424.500 82.800 425.400 ;
        RECT 70.950 422.400 73.050 424.500 ;
        RECT 53.400 419.700 58.050 420.900 ;
        RECT 56.700 415.050 58.050 419.700 ;
        RECT 49.950 412.950 52.050 415.050 ;
        RECT 50.100 411.150 51.900 412.950 ;
        RECT 53.100 412.050 54.900 413.850 ;
        RECT 55.950 412.950 58.050 415.050 ;
        RECT 52.950 409.950 55.050 412.050 ;
        RECT 56.700 405.600 57.900 412.950 ;
        RECT 59.100 412.050 60.900 413.850 ;
        RECT 61.950 412.950 64.050 415.050 ;
        RECT 58.950 409.950 61.050 412.050 ;
        RECT 62.100 411.150 63.900 412.950 ;
        RECT 66.150 407.700 67.050 422.400 ;
        RECT 74.550 421.800 76.350 423.600 ;
        RECT 77.850 423.450 82.800 424.500 ;
        RECT 90.300 424.500 91.350 425.400 ;
        RECT 77.850 422.700 79.650 423.450 ;
        RECT 90.300 423.300 94.050 424.500 ;
        RECT 91.950 422.400 94.050 423.300 ;
        RECT 97.650 422.400 99.450 428.400 ;
        RECT 112.800 425.400 114.600 428.400 ;
        RECT 133.800 425.400 135.600 428.400 ;
        RECT 74.850 420.000 75.900 421.800 ;
        RECT 85.050 420.000 86.850 420.600 ;
        RECT 74.850 418.800 86.850 420.000 ;
        RECT 69.000 417.600 75.900 418.800 ;
        RECT 69.000 416.850 69.900 417.600 ;
        RECT 74.100 417.000 75.900 417.600 ;
        RECT 68.100 415.050 69.900 416.850 ;
        RECT 71.100 415.800 72.900 416.400 ;
        RECT 67.950 412.950 70.050 415.050 ;
        RECT 71.100 414.600 79.050 415.800 ;
        RECT 76.950 412.950 79.050 414.600 ;
        RECT 75.450 407.700 77.250 408.000 ;
        RECT 66.150 407.100 77.250 407.700 ;
        RECT 66.150 406.500 83.850 407.100 ;
        RECT 66.150 405.600 67.050 406.500 ;
        RECT 75.450 406.200 83.850 406.500 ;
        RECT 43.950 400.950 46.050 403.050 ;
        RECT 55.800 393.600 59.100 405.600 ;
        RECT 66.150 393.600 67.950 405.600 ;
        RECT 80.250 404.700 82.050 405.300 ;
        RECT 74.550 403.500 82.050 404.700 ;
        RECT 82.950 404.100 83.850 406.200 ;
        RECT 85.950 406.200 86.850 418.800 ;
        RECT 98.250 415.050 99.450 422.400 ;
        RECT 93.150 413.250 99.450 415.050 ;
        RECT 94.950 412.950 99.450 413.250 ;
        RECT 95.250 407.400 97.050 409.200 ;
        RECT 91.950 406.200 96.150 407.400 ;
        RECT 85.950 405.300 91.050 406.200 ;
        RECT 91.950 405.300 94.050 406.200 ;
        RECT 98.250 405.600 99.450 412.950 ;
        RECT 113.400 412.050 114.600 425.400 ;
        RECT 130.950 415.950 133.050 418.050 ;
        RECT 115.950 412.950 118.050 415.050 ;
        RECT 131.100 414.150 132.900 415.950 ;
        RECT 134.400 415.050 135.300 425.400 ;
        RECT 140.550 422.400 142.350 428.400 ;
        RECT 148.650 425.400 150.450 428.400 ;
        RECT 156.450 425.400 158.250 428.400 ;
        RECT 164.250 426.300 166.050 428.400 ;
        RECT 164.250 425.400 168.000 426.300 ;
        RECT 148.650 424.500 149.700 425.400 ;
        RECT 145.950 423.300 149.700 424.500 ;
        RECT 157.200 424.500 158.250 425.400 ;
        RECT 166.950 424.500 168.000 425.400 ;
        RECT 157.200 423.450 162.150 424.500 ;
        RECT 145.950 422.400 148.050 423.300 ;
        RECT 160.350 422.700 162.150 423.450 ;
        RECT 136.950 415.950 139.050 418.050 ;
        RECT 133.950 412.950 136.050 415.050 ;
        RECT 137.100 414.150 138.900 415.950 ;
        RECT 140.550 415.050 141.750 422.400 ;
        RECT 163.650 421.800 165.450 423.600 ;
        RECT 166.950 422.400 169.050 424.500 ;
        RECT 172.050 422.400 173.850 428.400 ;
        RECT 153.150 420.000 154.950 420.600 ;
        RECT 164.100 420.000 165.150 421.800 ;
        RECT 153.150 418.800 165.150 420.000 ;
        RECT 140.550 413.250 146.850 415.050 ;
        RECT 140.550 412.950 145.050 413.250 ;
        RECT 112.950 406.950 115.050 412.050 ;
        RECT 116.100 411.150 117.900 412.950 ;
        RECT 90.150 404.400 91.050 405.300 ;
        RECT 87.450 404.100 89.250 404.400 ;
        RECT 74.550 402.600 75.750 403.500 ;
        RECT 82.950 403.200 89.250 404.100 ;
        RECT 87.450 402.600 89.250 403.200 ;
        RECT 90.150 402.600 92.850 404.400 ;
        RECT 70.950 400.500 75.750 402.600 ;
        RECT 78.450 401.550 80.250 402.300 ;
        RECT 83.250 401.550 85.050 402.300 ;
        RECT 78.450 400.500 85.050 401.550 ;
        RECT 74.550 399.600 75.750 400.500 ;
        RECT 74.550 393.600 76.350 399.600 ;
        RECT 82.350 393.600 84.150 400.500 ;
        RECT 90.150 399.600 94.050 401.700 ;
        RECT 90.150 393.600 91.950 399.600 ;
        RECT 97.650 393.600 99.450 405.600 ;
        RECT 113.400 399.600 114.600 406.950 ;
        RECT 134.400 405.600 135.300 412.950 ;
        RECT 112.800 393.600 114.600 399.600 ;
        RECT 131.700 404.400 135.300 405.600 ;
        RECT 140.550 405.600 141.750 412.950 ;
        RECT 142.950 407.400 144.750 409.200 ;
        RECT 143.850 406.200 148.050 407.400 ;
        RECT 153.150 406.200 154.050 418.800 ;
        RECT 164.100 417.600 171.000 418.800 ;
        RECT 164.100 417.000 165.900 417.600 ;
        RECT 170.100 416.850 171.000 417.600 ;
        RECT 167.100 415.800 168.900 416.400 ;
        RECT 160.950 414.600 168.900 415.800 ;
        RECT 170.100 415.050 171.900 416.850 ;
        RECT 160.950 412.950 163.050 414.600 ;
        RECT 169.950 412.950 172.050 415.050 ;
        RECT 162.750 407.700 164.550 408.000 ;
        RECT 172.950 407.700 173.850 422.400 ;
        RECT 162.750 407.100 173.850 407.700 ;
        RECT 131.700 393.600 133.500 404.400 ;
        RECT 140.550 393.600 142.350 405.600 ;
        RECT 145.950 405.300 148.050 406.200 ;
        RECT 148.950 405.300 154.050 406.200 ;
        RECT 156.150 406.500 173.850 407.100 ;
        RECT 156.150 406.200 164.550 406.500 ;
        RECT 148.950 404.400 149.850 405.300 ;
        RECT 147.150 402.600 149.850 404.400 ;
        RECT 150.750 404.100 152.550 404.400 ;
        RECT 156.150 404.100 157.050 406.200 ;
        RECT 172.950 405.600 173.850 406.500 ;
        RECT 150.750 403.200 157.050 404.100 ;
        RECT 157.950 404.700 159.750 405.300 ;
        RECT 157.950 403.500 165.450 404.700 ;
        RECT 150.750 402.600 152.550 403.200 ;
        RECT 164.250 402.600 165.450 403.500 ;
        RECT 145.950 399.600 149.850 401.700 ;
        RECT 154.950 401.550 156.750 402.300 ;
        RECT 159.750 401.550 161.550 402.300 ;
        RECT 154.950 400.500 161.550 401.550 ;
        RECT 164.250 400.500 169.050 402.600 ;
        RECT 148.050 393.600 149.850 399.600 ;
        RECT 155.850 393.600 157.650 400.500 ;
        RECT 164.250 399.600 165.450 400.500 ;
        RECT 163.650 393.600 165.450 399.600 ;
        RECT 172.050 393.600 173.850 405.600 ;
        RECT 176.550 422.400 178.350 428.400 ;
        RECT 184.650 425.400 186.450 428.400 ;
        RECT 192.450 425.400 194.250 428.400 ;
        RECT 200.250 426.300 202.050 428.400 ;
        RECT 200.250 425.400 204.000 426.300 ;
        RECT 184.650 424.500 185.700 425.400 ;
        RECT 181.950 423.300 185.700 424.500 ;
        RECT 193.200 424.500 194.250 425.400 ;
        RECT 202.950 424.500 204.000 425.400 ;
        RECT 193.200 423.450 198.150 424.500 ;
        RECT 181.950 422.400 184.050 423.300 ;
        RECT 196.350 422.700 198.150 423.450 ;
        RECT 176.550 415.050 177.750 422.400 ;
        RECT 199.650 421.800 201.450 423.600 ;
        RECT 202.950 422.400 205.050 424.500 ;
        RECT 208.050 422.400 209.850 428.400 ;
        RECT 189.150 420.000 190.950 420.600 ;
        RECT 200.100 420.000 201.150 421.800 ;
        RECT 189.150 418.800 201.150 420.000 ;
        RECT 176.550 413.250 182.850 415.050 ;
        RECT 176.550 412.950 181.050 413.250 ;
        RECT 176.550 405.600 177.750 412.950 ;
        RECT 178.950 407.400 180.750 409.200 ;
        RECT 179.850 406.200 184.050 407.400 ;
        RECT 189.150 406.200 190.050 418.800 ;
        RECT 200.100 417.600 207.000 418.800 ;
        RECT 200.100 417.000 201.900 417.600 ;
        RECT 206.100 416.850 207.000 417.600 ;
        RECT 203.100 415.800 204.900 416.400 ;
        RECT 196.950 414.600 204.900 415.800 ;
        RECT 206.100 415.050 207.900 416.850 ;
        RECT 196.950 412.950 199.050 414.600 ;
        RECT 205.950 412.950 208.050 415.050 ;
        RECT 198.750 407.700 200.550 408.000 ;
        RECT 208.950 407.700 209.850 422.400 ;
        RECT 198.750 407.100 209.850 407.700 ;
        RECT 176.550 393.600 178.350 405.600 ;
        RECT 181.950 405.300 184.050 406.200 ;
        RECT 184.950 405.300 190.050 406.200 ;
        RECT 192.150 406.500 209.850 407.100 ;
        RECT 192.150 406.200 200.550 406.500 ;
        RECT 184.950 404.400 185.850 405.300 ;
        RECT 183.150 402.600 185.850 404.400 ;
        RECT 186.750 404.100 188.550 404.400 ;
        RECT 192.150 404.100 193.050 406.200 ;
        RECT 208.950 405.600 209.850 406.500 ;
        RECT 186.750 403.200 193.050 404.100 ;
        RECT 193.950 404.700 195.750 405.300 ;
        RECT 193.950 403.500 201.450 404.700 ;
        RECT 186.750 402.600 188.550 403.200 ;
        RECT 200.250 402.600 201.450 403.500 ;
        RECT 181.950 399.600 185.850 401.700 ;
        RECT 190.950 401.550 192.750 402.300 ;
        RECT 195.750 401.550 197.550 402.300 ;
        RECT 190.950 400.500 197.550 401.550 ;
        RECT 200.250 400.500 205.050 402.600 ;
        RECT 184.050 393.600 185.850 399.600 ;
        RECT 191.850 393.600 193.650 400.500 ;
        RECT 200.250 399.600 201.450 400.500 ;
        RECT 199.650 393.600 201.450 399.600 ;
        RECT 208.050 393.600 209.850 405.600 ;
        RECT 213.150 422.400 214.950 428.400 ;
        RECT 220.950 426.300 222.750 428.400 ;
        RECT 219.000 425.400 222.750 426.300 ;
        RECT 228.750 425.400 230.550 428.400 ;
        RECT 236.550 425.400 238.350 428.400 ;
        RECT 219.000 424.500 220.050 425.400 ;
        RECT 228.750 424.500 229.800 425.400 ;
        RECT 217.950 422.400 220.050 424.500 ;
        RECT 213.150 407.700 214.050 422.400 ;
        RECT 221.550 421.800 223.350 423.600 ;
        RECT 224.850 423.450 229.800 424.500 ;
        RECT 237.300 424.500 238.350 425.400 ;
        RECT 224.850 422.700 226.650 423.450 ;
        RECT 237.300 423.300 241.050 424.500 ;
        RECT 238.950 422.400 241.050 423.300 ;
        RECT 244.650 422.400 246.450 428.400 ;
        RECT 221.850 420.000 222.900 421.800 ;
        RECT 232.050 420.000 233.850 420.600 ;
        RECT 221.850 418.800 233.850 420.000 ;
        RECT 216.000 417.600 222.900 418.800 ;
        RECT 216.000 416.850 216.900 417.600 ;
        RECT 221.100 417.000 222.900 417.600 ;
        RECT 215.100 415.050 216.900 416.850 ;
        RECT 218.100 415.800 219.900 416.400 ;
        RECT 214.950 412.950 217.050 415.050 ;
        RECT 218.100 414.600 226.050 415.800 ;
        RECT 223.950 412.950 226.050 414.600 ;
        RECT 222.450 407.700 224.250 408.000 ;
        RECT 213.150 407.100 224.250 407.700 ;
        RECT 213.150 406.500 230.850 407.100 ;
        RECT 213.150 405.600 214.050 406.500 ;
        RECT 222.450 406.200 230.850 406.500 ;
        RECT 213.150 393.600 214.950 405.600 ;
        RECT 227.250 404.700 229.050 405.300 ;
        RECT 221.550 403.500 229.050 404.700 ;
        RECT 229.950 404.100 230.850 406.200 ;
        RECT 232.950 406.200 233.850 418.800 ;
        RECT 245.250 415.050 246.450 422.400 ;
        RECT 260.400 425.400 262.200 428.400 ;
        RECT 278.400 425.400 280.200 428.400 ;
        RECT 301.800 425.400 303.600 428.400 ;
        RECT 320.400 425.400 322.200 428.400 ;
        RECT 335.400 425.400 337.200 428.400 ;
        RECT 240.150 413.250 246.450 415.050 ;
        RECT 241.950 412.950 246.450 413.250 ;
        RECT 256.950 412.950 259.050 415.050 ;
        RECT 242.250 407.400 244.050 409.200 ;
        RECT 238.950 406.200 243.150 407.400 ;
        RECT 232.950 405.300 238.050 406.200 ;
        RECT 238.950 405.300 241.050 406.200 ;
        RECT 245.250 405.600 246.450 412.950 ;
        RECT 257.100 411.150 258.900 412.950 ;
        RECT 260.400 412.050 261.600 425.400 ;
        RECT 265.950 418.950 268.050 421.050 ;
        RECT 259.950 406.950 262.050 412.050 ;
        RECT 237.150 404.400 238.050 405.300 ;
        RECT 234.450 404.100 236.250 404.400 ;
        RECT 221.550 402.600 222.750 403.500 ;
        RECT 229.950 403.200 236.250 404.100 ;
        RECT 234.450 402.600 236.250 403.200 ;
        RECT 237.150 402.600 239.850 404.400 ;
        RECT 217.950 400.500 222.750 402.600 ;
        RECT 225.450 401.550 227.250 402.300 ;
        RECT 230.250 401.550 232.050 402.300 ;
        RECT 225.450 400.500 232.050 401.550 ;
        RECT 221.550 399.600 222.750 400.500 ;
        RECT 221.550 393.600 223.350 399.600 ;
        RECT 229.350 393.600 231.150 400.500 ;
        RECT 237.150 399.600 241.050 401.700 ;
        RECT 237.150 393.600 238.950 399.600 ;
        RECT 244.650 393.600 246.450 405.600 ;
        RECT 247.950 400.950 250.050 403.050 ;
        RECT 248.550 397.050 249.450 400.950 ;
        RECT 260.400 399.600 261.600 406.950 ;
        RECT 266.550 400.050 267.450 418.950 ;
        RECT 274.950 415.950 277.050 418.050 ;
        RECT 275.100 414.150 276.900 415.950 ;
        RECT 278.700 415.050 279.600 425.400 ;
        RECT 280.950 415.950 283.050 418.050 ;
        RECT 298.950 415.950 301.050 418.050 ;
        RECT 277.950 412.950 280.050 415.050 ;
        RECT 281.100 414.150 282.900 415.950 ;
        RECT 299.100 414.150 300.900 415.950 ;
        RECT 302.400 415.050 303.300 425.400 ;
        RECT 310.950 418.950 313.050 421.050 ;
        RECT 304.950 415.950 307.050 418.050 ;
        RECT 301.950 412.950 304.050 415.050 ;
        RECT 305.100 414.150 306.900 415.950 ;
        RECT 278.700 405.600 279.600 412.950 ;
        RECT 302.400 405.600 303.300 412.950 ;
        RECT 278.700 404.400 282.300 405.600 ;
        RECT 247.950 394.950 250.050 397.050 ;
        RECT 260.400 393.600 262.200 399.600 ;
        RECT 265.950 397.950 268.050 400.050 ;
        RECT 280.500 393.600 282.300 404.400 ;
        RECT 299.700 404.400 303.300 405.600 ;
        RECT 299.700 393.600 301.500 404.400 ;
        RECT 311.550 397.050 312.450 418.950 ;
        RECT 316.950 412.950 319.050 415.050 ;
        RECT 317.100 411.150 318.900 412.950 ;
        RECT 320.400 412.050 321.600 425.400 ;
        RECT 335.400 421.500 336.600 425.400 ;
        RECT 341.700 422.400 343.500 428.400 ;
        RECT 335.400 420.600 341.400 421.500 ;
        RECT 339.150 419.700 341.400 420.600 ;
        RECT 334.950 412.950 337.050 415.050 ;
        RECT 319.950 406.950 322.050 412.050 ;
        RECT 335.100 411.150 336.900 412.950 ;
        RECT 339.150 408.300 340.050 419.700 ;
        RECT 342.300 415.050 343.500 422.400 ;
        RECT 359.400 421.200 361.200 428.400 ;
        RECT 382.800 421.200 384.600 428.400 ;
        RECT 403.800 425.400 405.600 428.400 ;
        RECT 359.400 420.300 363.600 421.200 ;
        RECT 362.400 415.050 363.600 420.300 ;
        RECT 380.400 420.300 384.600 421.200 ;
        RECT 380.400 415.050 381.600 420.300 ;
        RECT 400.950 415.950 403.050 418.050 ;
        RECT 340.950 412.950 343.500 415.050 ;
        RECT 339.150 407.400 341.400 408.300 ;
        RECT 320.400 399.600 321.600 406.950 ;
        RECT 335.400 406.500 341.400 407.400 ;
        RECT 335.400 399.600 336.600 406.500 ;
        RECT 342.300 405.600 343.500 412.950 ;
        RECT 359.100 412.050 360.900 413.850 ;
        RECT 361.950 412.950 364.050 415.050 ;
        RECT 358.950 409.950 361.050 412.050 ;
        RECT 310.950 394.950 313.050 397.050 ;
        RECT 320.400 393.600 322.200 399.600 ;
        RECT 335.400 393.600 337.200 399.600 ;
        RECT 341.700 393.600 343.500 405.600 ;
        RECT 362.400 399.600 363.600 412.950 ;
        RECT 365.100 412.050 366.900 413.850 ;
        RECT 377.100 412.050 378.900 413.850 ;
        RECT 379.950 412.950 382.050 415.050 ;
        RECT 401.100 414.150 402.900 415.950 ;
        RECT 404.400 415.050 405.300 425.400 ;
        RECT 419.400 423.300 421.200 428.400 ;
        RECT 425.400 423.300 427.200 428.400 ;
        RECT 419.400 421.950 427.200 423.300 ;
        RECT 428.400 422.400 430.200 428.400 ;
        RECT 443.400 425.400 445.200 428.400 ;
        RECT 428.400 420.300 429.600 422.400 ;
        RECT 443.400 421.500 444.600 425.400 ;
        RECT 449.700 422.400 451.500 428.400 ;
        RECT 443.400 420.600 449.400 421.500 ;
        RECT 425.850 419.250 429.600 420.300 ;
        RECT 447.150 419.700 449.400 420.600 ;
        RECT 406.950 415.950 409.050 418.050 ;
        RECT 364.950 409.950 367.050 412.050 ;
        RECT 376.950 409.950 379.050 412.050 ;
        RECT 361.800 393.600 363.600 399.600 ;
        RECT 380.400 399.600 381.600 412.950 ;
        RECT 383.100 412.050 384.900 413.850 ;
        RECT 403.950 412.950 406.050 415.050 ;
        RECT 407.100 414.150 408.900 415.950 ;
        RECT 425.850 415.050 427.050 419.250 ;
        RECT 418.950 412.950 421.050 415.050 ;
        RECT 382.950 409.950 385.050 412.050 ;
        RECT 404.400 405.600 405.300 412.950 ;
        RECT 419.100 411.150 420.900 412.950 ;
        RECT 422.100 412.050 423.900 413.850 ;
        RECT 424.950 412.950 427.050 415.050 ;
        RECT 421.950 409.950 424.050 412.050 ;
        RECT 401.700 404.400 405.300 405.600 ;
        RECT 380.400 393.600 382.200 399.600 ;
        RECT 401.700 393.600 403.500 404.400 ;
        RECT 424.950 399.600 426.150 412.950 ;
        RECT 428.100 412.050 429.900 413.850 ;
        RECT 442.950 412.950 445.050 415.050 ;
        RECT 427.950 409.950 430.050 412.050 ;
        RECT 443.100 411.150 444.900 412.950 ;
        RECT 447.150 408.300 448.050 419.700 ;
        RECT 450.300 415.050 451.500 422.400 ;
        RECT 448.950 412.950 451.500 415.050 ;
        RECT 447.150 407.400 449.400 408.300 ;
        RECT 443.400 406.500 449.400 407.400 ;
        RECT 443.400 399.600 444.600 406.500 ;
        RECT 450.300 405.600 451.500 412.950 ;
        RECT 424.800 393.600 426.600 399.600 ;
        RECT 443.400 393.600 445.200 399.600 ;
        RECT 449.700 393.600 451.500 405.600 ;
        RECT 466.500 422.400 468.300 428.400 ;
        RECT 472.800 425.400 474.600 428.400 ;
        RECT 466.500 415.050 467.700 422.400 ;
        RECT 473.400 421.500 474.600 425.400 ;
        RECT 485.400 423.300 487.200 428.400 ;
        RECT 491.400 423.300 493.200 428.400 ;
        RECT 485.400 421.950 493.200 423.300 ;
        RECT 494.400 422.400 496.200 428.400 ;
        RECT 468.600 420.600 474.600 421.500 ;
        RECT 468.600 419.700 470.850 420.600 ;
        RECT 494.400 420.300 495.600 422.400 ;
        RECT 466.500 412.950 469.050 415.050 ;
        RECT 466.500 405.600 467.700 412.950 ;
        RECT 469.950 408.300 470.850 419.700 ;
        RECT 491.850 419.250 495.600 420.300 ;
        RECT 514.200 420.000 516.000 428.400 ;
        RECT 538.200 420.000 540.000 428.400 ;
        RECT 560.400 421.200 562.200 428.400 ;
        RECT 560.400 420.300 564.600 421.200 ;
        RECT 491.850 415.050 493.050 419.250 ;
        RECT 512.700 418.800 516.000 420.000 ;
        RECT 536.700 418.800 540.000 420.000 ;
        RECT 505.950 415.950 508.050 418.050 ;
        RECT 472.950 412.950 475.050 415.050 ;
        RECT 484.950 412.950 487.050 415.050 ;
        RECT 473.100 411.150 474.900 412.950 ;
        RECT 485.100 411.150 486.900 412.950 ;
        RECT 488.100 412.050 489.900 413.850 ;
        RECT 490.950 412.950 493.050 415.050 ;
        RECT 487.950 409.950 490.050 412.050 ;
        RECT 468.600 407.400 470.850 408.300 ;
        RECT 468.600 406.500 474.600 407.400 ;
        RECT 466.500 393.600 468.300 405.600 ;
        RECT 473.400 399.600 474.600 406.500 ;
        RECT 490.950 399.600 492.150 412.950 ;
        RECT 494.100 412.050 495.900 413.850 ;
        RECT 493.950 409.950 496.050 412.050 ;
        RECT 506.550 400.050 507.450 415.950 ;
        RECT 512.700 415.050 513.600 418.800 ;
        RECT 536.700 415.050 537.600 418.800 ;
        RECT 563.400 415.050 564.600 420.300 ;
        RECT 583.200 420.000 585.000 428.400 ;
        RECT 601.800 425.400 603.600 428.400 ;
        RECT 619.800 425.400 621.600 428.400 ;
        RECT 581.700 418.800 585.000 420.000 ;
        RECT 581.700 415.050 582.600 418.800 ;
        RECT 511.950 412.950 514.050 415.050 ;
        RECT 512.700 400.800 513.600 412.950 ;
        RECT 515.100 412.050 516.900 413.850 ;
        RECT 517.950 412.950 520.050 415.050 ;
        RECT 514.950 409.950 517.050 412.050 ;
        RECT 518.100 411.150 519.900 412.950 ;
        RECT 521.100 412.050 522.900 413.850 ;
        RECT 535.950 412.950 538.050 415.050 ;
        RECT 520.950 409.950 523.050 412.050 ;
        RECT 536.700 400.800 537.600 412.950 ;
        RECT 539.100 412.050 540.900 413.850 ;
        RECT 541.950 412.950 544.050 415.050 ;
        RECT 538.950 409.950 541.050 412.050 ;
        RECT 542.100 411.150 543.900 412.950 ;
        RECT 545.100 412.050 546.900 413.850 ;
        RECT 560.100 412.050 561.900 413.850 ;
        RECT 562.950 412.950 565.050 415.050 ;
        RECT 544.950 409.950 547.050 412.050 ;
        RECT 559.950 409.950 562.050 412.050 ;
        RECT 472.800 393.600 474.600 399.600 ;
        RECT 490.800 393.600 492.600 399.600 ;
        RECT 505.950 397.950 508.050 400.050 ;
        RECT 512.700 399.900 519.300 400.800 ;
        RECT 512.700 399.600 513.600 399.900 ;
        RECT 511.800 393.600 513.600 399.600 ;
        RECT 517.800 399.600 519.300 399.900 ;
        RECT 536.700 399.900 543.300 400.800 ;
        RECT 536.700 399.600 537.600 399.900 ;
        RECT 517.800 393.600 519.600 399.600 ;
        RECT 535.800 393.600 537.600 399.600 ;
        RECT 541.800 399.600 543.300 399.900 ;
        RECT 563.400 399.600 564.600 412.950 ;
        RECT 566.100 412.050 567.900 413.850 ;
        RECT 580.950 412.950 583.050 415.050 ;
        RECT 565.950 409.950 568.050 412.050 ;
        RECT 581.700 400.800 582.600 412.950 ;
        RECT 584.100 412.050 585.900 413.850 ;
        RECT 586.950 412.950 589.050 415.050 ;
        RECT 583.950 409.950 586.050 412.050 ;
        RECT 587.100 411.150 588.900 412.950 ;
        RECT 590.100 412.050 591.900 413.850 ;
        RECT 602.400 412.050 603.600 425.400 ;
        RECT 604.950 412.950 607.050 415.050 ;
        RECT 589.950 409.950 592.050 412.050 ;
        RECT 601.950 406.950 604.050 412.050 ;
        RECT 605.100 411.150 606.900 412.950 ;
        RECT 620.400 412.050 621.600 425.400 ;
        RECT 635.400 423.300 637.200 428.400 ;
        RECT 641.400 423.300 643.200 428.400 ;
        RECT 635.400 421.950 643.200 423.300 ;
        RECT 644.400 422.400 646.200 428.400 ;
        RECT 662.400 425.400 664.200 428.400 ;
        RECT 679.800 425.400 681.600 428.400 ;
        RECT 700.800 425.400 702.600 428.400 ;
        RECT 644.400 420.300 645.600 422.400 ;
        RECT 641.850 419.250 645.600 420.300 ;
        RECT 641.850 415.050 643.050 419.250 ;
        RECT 622.950 412.950 625.050 415.050 ;
        RECT 634.950 412.950 637.050 415.050 ;
        RECT 619.950 406.950 622.050 412.050 ;
        RECT 623.100 411.150 624.900 412.950 ;
        RECT 635.100 411.150 636.900 412.950 ;
        RECT 638.100 412.050 639.900 413.850 ;
        RECT 640.950 412.950 643.050 415.050 ;
        RECT 637.950 409.950 640.050 412.050 ;
        RECT 581.700 399.900 588.300 400.800 ;
        RECT 581.700 399.600 582.600 399.900 ;
        RECT 541.800 393.600 543.600 399.600 ;
        RECT 562.800 393.600 564.600 399.600 ;
        RECT 580.800 393.600 582.600 399.600 ;
        RECT 586.800 399.600 588.300 399.900 ;
        RECT 602.400 399.600 603.600 406.950 ;
        RECT 620.400 399.600 621.600 406.950 ;
        RECT 640.950 399.600 642.150 412.950 ;
        RECT 644.100 412.050 645.900 413.850 ;
        RECT 658.950 412.950 661.050 415.050 ;
        RECT 643.950 409.950 646.050 412.050 ;
        RECT 659.100 411.150 660.900 412.950 ;
        RECT 662.400 412.050 663.600 425.400 ;
        RECT 680.400 412.050 681.600 425.400 ;
        RECT 697.950 415.950 700.050 418.050 ;
        RECT 682.950 412.950 685.050 415.050 ;
        RECT 698.100 414.150 699.900 415.950 ;
        RECT 701.400 415.050 702.300 425.400 ;
        RECT 716.400 423.300 718.200 428.400 ;
        RECT 722.400 423.300 724.200 428.400 ;
        RECT 716.400 421.950 724.200 423.300 ;
        RECT 725.400 422.400 727.200 428.400 ;
        RECT 742.800 425.400 744.600 428.400 ;
        RECT 763.800 425.400 765.600 428.400 ;
        RECT 784.800 425.400 786.600 428.400 ;
        RECT 725.400 420.300 726.600 422.400 ;
        RECT 722.850 419.250 726.600 420.300 ;
        RECT 703.950 415.950 706.050 418.050 ;
        RECT 709.950 415.950 712.050 418.050 ;
        RECT 700.950 412.950 703.050 415.050 ;
        RECT 704.100 414.150 705.900 415.950 ;
        RECT 661.950 406.950 664.050 412.050 ;
        RECT 679.950 406.950 682.050 412.050 ;
        RECT 683.100 411.150 684.900 412.950 ;
        RECT 662.400 399.600 663.600 406.950 ;
        RECT 680.400 399.600 681.600 406.950 ;
        RECT 701.400 405.600 702.300 412.950 ;
        RECT 710.550 406.050 711.450 415.950 ;
        RECT 722.850 415.050 724.050 419.250 ;
        RECT 730.950 415.950 733.050 418.050 ;
        RECT 715.950 412.950 718.050 415.050 ;
        RECT 716.100 411.150 717.900 412.950 ;
        RECT 719.100 412.050 720.900 413.850 ;
        RECT 721.950 412.950 724.050 415.050 ;
        RECT 718.950 409.950 721.050 412.050 ;
        RECT 586.800 393.600 588.600 399.600 ;
        RECT 601.800 393.600 603.600 399.600 ;
        RECT 619.800 393.600 621.600 399.600 ;
        RECT 640.800 393.600 642.600 399.600 ;
        RECT 662.400 393.600 664.200 399.600 ;
        RECT 679.800 393.600 681.600 399.600 ;
        RECT 698.700 404.400 702.300 405.600 ;
        RECT 698.700 393.600 700.500 404.400 ;
        RECT 709.950 403.950 712.050 406.050 ;
        RECT 721.950 399.600 723.150 412.950 ;
        RECT 725.100 412.050 726.900 413.850 ;
        RECT 724.950 409.950 727.050 412.050 ;
        RECT 721.800 393.600 723.600 399.600 ;
        RECT 731.550 397.050 732.450 415.950 ;
        RECT 743.400 412.050 744.600 425.400 ;
        RECT 760.950 415.950 763.050 418.050 ;
        RECT 745.950 412.950 748.050 415.050 ;
        RECT 761.100 414.150 762.900 415.950 ;
        RECT 764.400 415.050 765.300 425.400 ;
        RECT 766.950 415.950 769.050 418.050 ;
        RECT 781.950 415.950 784.050 418.050 ;
        RECT 763.950 412.950 766.050 415.050 ;
        RECT 767.100 414.150 768.900 415.950 ;
        RECT 782.100 414.150 783.900 415.950 ;
        RECT 785.400 415.050 786.300 425.400 ;
        RECT 800.400 423.300 802.200 428.400 ;
        RECT 806.400 423.300 808.200 428.400 ;
        RECT 800.400 421.950 808.200 423.300 ;
        RECT 809.400 422.400 811.200 428.400 ;
        RECT 827.400 425.400 829.200 428.400 ;
        RECT 848.400 425.400 850.200 428.400 ;
        RECT 809.400 420.300 810.600 422.400 ;
        RECT 806.850 419.250 810.600 420.300 ;
        RECT 787.950 415.950 790.050 418.050 ;
        RECT 784.950 412.950 787.050 415.050 ;
        RECT 788.100 414.150 789.900 415.950 ;
        RECT 806.850 415.050 808.050 419.250 ;
        RECT 814.950 415.950 817.050 418.050 ;
        RECT 823.950 415.950 826.050 418.050 ;
        RECT 799.950 412.950 802.050 415.050 ;
        RECT 742.950 406.950 745.050 412.050 ;
        RECT 746.100 411.150 747.900 412.950 ;
        RECT 743.400 399.600 744.600 406.950 ;
        RECT 764.400 405.600 765.300 412.950 ;
        RECT 785.400 405.600 786.300 412.950 ;
        RECT 800.100 411.150 801.900 412.950 ;
        RECT 803.100 412.050 804.900 413.850 ;
        RECT 805.950 412.950 808.050 415.050 ;
        RECT 802.950 409.950 805.050 412.050 ;
        RECT 730.950 394.950 733.050 397.050 ;
        RECT 742.800 393.600 744.600 399.600 ;
        RECT 761.700 404.400 765.300 405.600 ;
        RECT 782.700 404.400 786.300 405.600 ;
        RECT 761.700 393.600 763.500 404.400 ;
        RECT 782.700 393.600 784.500 404.400 ;
        RECT 805.950 399.600 807.150 412.950 ;
        RECT 809.100 412.050 810.900 413.850 ;
        RECT 808.950 409.950 811.050 412.050 ;
        RECT 805.800 393.600 807.600 399.600 ;
        RECT 815.550 397.050 816.450 415.950 ;
        RECT 824.100 414.150 825.900 415.950 ;
        RECT 827.700 415.050 828.600 425.400 ;
        RECT 829.950 415.950 832.050 418.050 ;
        RECT 844.950 415.950 847.050 418.050 ;
        RECT 826.950 412.950 829.050 415.050 ;
        RECT 830.100 414.150 831.900 415.950 ;
        RECT 845.100 414.150 846.900 415.950 ;
        RECT 848.700 415.050 849.600 425.400 ;
        RECT 870.300 424.200 872.100 428.400 ;
        RECT 869.400 422.400 872.100 424.200 ;
        RECT 850.950 415.950 853.050 418.050 ;
        RECT 847.950 412.950 850.050 415.050 ;
        RECT 851.100 414.150 852.900 415.950 ;
        RECT 869.400 415.050 870.300 422.400 ;
        RECT 872.100 420.600 873.900 421.500 ;
        RECT 877.800 420.600 879.600 428.400 ;
        RECT 893.400 425.400 895.200 428.400 ;
        RECT 872.100 419.700 879.600 420.600 ;
        RECT 868.950 412.950 871.050 415.050 ;
        RECT 871.950 412.950 874.050 415.050 ;
        RECT 827.700 405.600 828.600 412.950 ;
        RECT 848.700 405.600 849.600 412.950 ;
        RECT 869.400 405.600 870.300 412.950 ;
        RECT 872.100 411.150 873.900 412.950 ;
        RECT 827.700 404.400 831.300 405.600 ;
        RECT 848.700 404.400 852.300 405.600 ;
        RECT 814.950 394.950 817.050 397.050 ;
        RECT 829.500 393.600 831.300 404.400 ;
        RECT 850.500 393.600 852.300 404.400 ;
        RECT 868.500 393.600 870.300 405.600 ;
        RECT 875.700 399.600 876.600 419.700 ;
        RECT 878.100 415.050 879.900 416.850 ;
        RECT 889.950 415.950 892.050 418.050 ;
        RECT 877.950 412.950 880.050 415.050 ;
        RECT 890.100 414.150 891.900 415.950 ;
        RECT 893.700 415.050 894.600 425.400 ;
        RECT 895.950 415.950 898.050 418.050 ;
        RECT 892.950 412.950 895.050 415.050 ;
        RECT 896.100 414.150 897.900 415.950 ;
        RECT 893.700 405.600 894.600 412.950 ;
        RECT 893.700 404.400 897.300 405.600 ;
        RECT 874.800 393.600 876.600 399.600 ;
        RECT 895.500 393.600 897.300 404.400 ;
        RECT 2.550 377.400 4.350 389.400 ;
        RECT 10.050 383.400 11.850 389.400 ;
        RECT 7.950 381.300 11.850 383.400 ;
        RECT 17.850 382.500 19.650 389.400 ;
        RECT 25.650 383.400 27.450 389.400 ;
        RECT 26.250 382.500 27.450 383.400 ;
        RECT 16.950 381.450 23.550 382.500 ;
        RECT 16.950 380.700 18.750 381.450 ;
        RECT 21.750 380.700 23.550 381.450 ;
        RECT 26.250 380.400 31.050 382.500 ;
        RECT 9.150 378.600 11.850 380.400 ;
        RECT 12.750 379.800 14.550 380.400 ;
        RECT 12.750 378.900 19.050 379.800 ;
        RECT 26.250 379.500 27.450 380.400 ;
        RECT 12.750 378.600 14.550 378.900 ;
        RECT 10.950 377.700 11.850 378.600 ;
        RECT 2.550 370.050 3.750 377.400 ;
        RECT 7.950 376.800 10.050 377.700 ;
        RECT 10.950 376.800 16.050 377.700 ;
        RECT 5.850 375.600 10.050 376.800 ;
        RECT 4.950 373.800 6.750 375.600 ;
        RECT 2.550 369.750 7.050 370.050 ;
        RECT 2.550 367.950 8.850 369.750 ;
        RECT 2.550 360.600 3.750 367.950 ;
        RECT 15.150 364.200 16.050 376.800 ;
        RECT 18.150 376.800 19.050 378.900 ;
        RECT 19.950 378.300 27.450 379.500 ;
        RECT 19.950 377.700 21.750 378.300 ;
        RECT 34.050 377.400 35.850 389.400 ;
        RECT 18.150 376.500 26.550 376.800 ;
        RECT 34.950 376.500 35.850 377.400 ;
        RECT 18.150 375.900 35.850 376.500 ;
        RECT 24.750 375.300 35.850 375.900 ;
        RECT 24.750 375.000 26.550 375.300 ;
        RECT 22.950 368.400 25.050 370.050 ;
        RECT 22.950 367.200 30.900 368.400 ;
        RECT 31.950 367.950 34.050 370.050 ;
        RECT 29.100 366.600 30.900 367.200 ;
        RECT 32.100 366.150 33.900 367.950 ;
        RECT 26.100 365.400 27.900 366.000 ;
        RECT 32.100 365.400 33.000 366.150 ;
        RECT 26.100 364.200 33.000 365.400 ;
        RECT 15.150 363.000 27.150 364.200 ;
        RECT 15.150 362.400 16.950 363.000 ;
        RECT 26.100 361.200 27.150 363.000 ;
        RECT 2.550 354.600 4.350 360.600 ;
        RECT 7.950 359.700 10.050 360.600 ;
        RECT 7.950 358.500 11.700 359.700 ;
        RECT 22.350 359.550 24.150 360.300 ;
        RECT 10.650 357.600 11.700 358.500 ;
        RECT 19.200 358.500 24.150 359.550 ;
        RECT 25.650 359.400 27.450 361.200 ;
        RECT 34.950 360.600 35.850 375.300 ;
        RECT 28.950 358.500 31.050 360.600 ;
        RECT 19.200 357.600 20.250 358.500 ;
        RECT 28.950 357.600 30.000 358.500 ;
        RECT 10.650 354.600 12.450 357.600 ;
        RECT 18.450 354.600 20.250 357.600 ;
        RECT 26.250 356.700 30.000 357.600 ;
        RECT 26.250 354.600 28.050 356.700 ;
        RECT 34.050 354.600 35.850 360.600 ;
        RECT 39.150 377.400 40.950 389.400 ;
        RECT 47.550 383.400 49.350 389.400 ;
        RECT 47.550 382.500 48.750 383.400 ;
        RECT 55.350 382.500 57.150 389.400 ;
        RECT 63.150 383.400 64.950 389.400 ;
        RECT 43.950 380.400 48.750 382.500 ;
        RECT 51.450 381.450 58.050 382.500 ;
        RECT 51.450 380.700 53.250 381.450 ;
        RECT 56.250 380.700 58.050 381.450 ;
        RECT 63.150 381.300 67.050 383.400 ;
        RECT 47.550 379.500 48.750 380.400 ;
        RECT 60.450 379.800 62.250 380.400 ;
        RECT 47.550 378.300 55.050 379.500 ;
        RECT 53.250 377.700 55.050 378.300 ;
        RECT 55.950 378.900 62.250 379.800 ;
        RECT 39.150 376.500 40.050 377.400 ;
        RECT 55.950 376.800 56.850 378.900 ;
        RECT 60.450 378.600 62.250 378.900 ;
        RECT 63.150 378.600 65.850 380.400 ;
        RECT 63.150 377.700 64.050 378.600 ;
        RECT 48.450 376.500 56.850 376.800 ;
        RECT 39.150 375.900 56.850 376.500 ;
        RECT 58.950 376.800 64.050 377.700 ;
        RECT 64.950 376.800 67.050 377.700 ;
        RECT 70.650 377.400 72.450 389.400 ;
        RECT 85.800 383.400 87.600 389.400 ;
        RECT 39.150 375.300 50.250 375.900 ;
        RECT 39.150 360.600 40.050 375.300 ;
        RECT 48.450 375.000 50.250 375.300 ;
        RECT 40.950 367.950 43.050 370.050 ;
        RECT 49.950 368.400 52.050 370.050 ;
        RECT 41.100 366.150 42.900 367.950 ;
        RECT 44.100 367.200 52.050 368.400 ;
        RECT 44.100 366.600 45.900 367.200 ;
        RECT 42.000 365.400 42.900 366.150 ;
        RECT 47.100 365.400 48.900 366.000 ;
        RECT 42.000 364.200 48.900 365.400 ;
        RECT 58.950 364.200 59.850 376.800 ;
        RECT 64.950 375.600 69.150 376.800 ;
        RECT 68.250 373.800 70.050 375.600 ;
        RECT 71.250 370.050 72.450 377.400 ;
        RECT 86.400 376.050 87.600 383.400 ;
        RECT 103.800 377.400 105.600 389.400 ;
        RECT 106.800 378.300 108.600 389.400 ;
        RECT 112.800 378.300 114.600 389.400 ;
        RECT 106.800 377.400 114.600 378.300 ;
        RECT 128.700 378.600 130.500 389.400 ;
        RECT 128.700 377.400 132.300 378.600 ;
        RECT 85.950 370.950 88.050 376.050 ;
        RECT 67.950 369.750 72.450 370.050 ;
        RECT 66.150 367.950 72.450 369.750 ;
        RECT 47.850 363.000 59.850 364.200 ;
        RECT 47.850 361.200 48.900 363.000 ;
        RECT 58.050 362.400 59.850 363.000 ;
        RECT 39.150 354.600 40.950 360.600 ;
        RECT 43.950 358.500 46.050 360.600 ;
        RECT 47.550 359.400 49.350 361.200 ;
        RECT 71.250 360.600 72.450 367.950 ;
        RECT 50.850 359.550 52.650 360.300 ;
        RECT 64.950 359.700 67.050 360.600 ;
        RECT 50.850 358.500 55.800 359.550 ;
        RECT 45.000 357.600 46.050 358.500 ;
        RECT 54.750 357.600 55.800 358.500 ;
        RECT 63.300 358.500 67.050 359.700 ;
        RECT 63.300 357.600 64.350 358.500 ;
        RECT 45.000 356.700 48.750 357.600 ;
        RECT 46.950 354.600 48.750 356.700 ;
        RECT 54.750 354.600 56.550 357.600 ;
        RECT 62.550 354.600 64.350 357.600 ;
        RECT 70.650 354.600 72.450 360.600 ;
        RECT 86.400 357.600 87.600 370.950 ;
        RECT 89.100 370.050 90.900 371.850 ;
        RECT 104.400 370.050 105.600 377.400 ;
        RECT 106.950 370.950 109.050 373.050 ;
        RECT 88.950 367.950 91.050 370.050 ;
        RECT 103.950 367.950 106.050 370.050 ;
        RECT 107.100 369.150 108.900 370.950 ;
        RECT 110.100 370.050 111.900 371.850 ;
        RECT 112.950 370.950 115.050 373.050 ;
        RECT 109.950 367.950 112.050 370.050 ;
        RECT 113.100 369.150 114.900 370.950 ;
        RECT 131.400 370.050 132.300 377.400 ;
        RECT 146.400 377.400 148.200 389.400 ;
        RECT 153.900 378.900 155.700 389.400 ;
        RECT 173.400 383.400 175.200 389.400 ;
        RECT 184.950 385.950 187.050 388.050 ;
        RECT 153.900 377.400 156.300 378.900 ;
        RECT 146.400 375.900 147.600 377.400 ;
        RECT 146.400 374.700 153.600 375.900 ;
        RECT 151.800 374.100 153.600 374.700 ;
        RECT 145.950 370.950 148.050 373.050 ;
        RECT 104.400 360.600 105.600 367.950 ;
        RECT 128.100 367.050 129.900 368.850 ;
        RECT 130.950 367.950 133.050 370.050 ;
        RECT 146.100 369.150 147.900 370.950 ;
        RECT 149.100 370.050 150.900 371.850 ;
        RECT 127.950 364.950 130.050 367.050 ;
        RECT 104.400 359.400 109.500 360.600 ;
        RECT 85.800 354.600 87.600 357.600 ;
        RECT 107.700 354.600 109.500 359.400 ;
        RECT 131.400 357.600 132.300 367.950 ;
        RECT 134.100 367.050 135.900 368.850 ;
        RECT 148.950 367.950 151.050 370.050 ;
        RECT 133.950 364.950 136.050 367.050 ;
        RECT 152.700 363.600 153.600 374.100 ;
        RECT 154.950 370.050 156.300 377.400 ;
        RECT 169.950 370.950 172.050 373.050 ;
        RECT 154.950 367.950 157.050 370.050 ;
        RECT 170.100 369.150 171.900 370.950 ;
        RECT 173.400 370.050 174.600 383.400 ;
        RECT 181.950 373.950 184.050 376.050 ;
        RECT 175.950 370.950 178.050 373.050 ;
        RECT 172.950 367.950 175.050 370.050 ;
        RECT 176.100 369.150 177.900 370.950 ;
        RECT 151.800 362.700 153.600 363.600 ;
        RECT 150.300 361.800 153.600 362.700 ;
        RECT 150.300 357.600 151.200 361.800 ;
        RECT 156.000 360.600 157.050 367.950 ;
        RECT 173.400 362.700 174.600 367.950 ;
        RECT 182.550 367.050 183.450 373.950 ;
        RECT 185.550 370.050 186.450 385.950 ;
        RECT 194.400 383.400 196.200 389.400 ;
        RECT 218.400 383.400 220.200 389.400 ;
        RECT 229.950 385.950 232.050 388.050 ;
        RECT 190.950 370.950 193.050 373.050 ;
        RECT 184.950 367.950 187.050 370.050 ;
        RECT 191.100 369.150 192.900 370.950 ;
        RECT 194.400 370.050 195.600 383.400 ;
        RECT 202.950 379.950 205.050 382.050 ;
        RECT 196.950 370.950 199.050 373.050 ;
        RECT 193.950 367.950 196.050 370.050 ;
        RECT 197.100 369.150 198.900 370.950 ;
        RECT 181.800 364.950 183.900 367.050 ;
        RECT 194.400 362.700 195.600 367.950 ;
        RECT 173.400 361.800 177.600 362.700 ;
        RECT 194.400 361.800 198.600 362.700 ;
        RECT 130.800 354.600 132.600 357.600 ;
        RECT 149.400 354.600 151.200 357.600 ;
        RECT 155.400 354.600 157.200 360.600 ;
        RECT 175.800 354.600 177.600 361.800 ;
        RECT 196.800 354.600 198.600 361.800 ;
        RECT 203.550 358.050 204.450 379.950 ;
        RECT 214.950 370.950 217.050 373.050 ;
        RECT 215.100 369.150 216.900 370.950 ;
        RECT 218.850 370.050 220.050 383.400 ;
        RECT 220.950 370.950 223.050 373.050 ;
        RECT 217.950 367.950 220.050 370.050 ;
        RECT 221.100 369.150 222.900 370.950 ;
        RECT 224.100 370.050 225.900 371.850 ;
        RECT 223.950 367.950 226.050 370.050 ;
        RECT 217.950 363.750 219.150 367.950 ;
        RECT 215.400 362.700 219.150 363.750 ;
        RECT 215.400 360.600 216.600 362.700 ;
        RECT 202.950 355.950 205.050 358.050 ;
        RECT 214.800 354.600 216.600 360.600 ;
        RECT 217.800 359.700 225.600 361.050 ;
        RECT 217.800 354.600 219.600 359.700 ;
        RECT 223.800 354.600 225.600 359.700 ;
        RECT 230.550 358.050 231.450 385.950 ;
        RECT 241.500 378.600 243.300 389.400 ;
        RECT 239.700 377.400 243.300 378.600 ;
        RECT 260.700 378.600 262.500 389.400 ;
        RECT 283.800 383.400 285.600 389.400 ;
        RECT 304.800 383.400 306.600 389.400 ;
        RECT 326.400 383.400 328.200 389.400 ;
        RECT 349.800 383.400 351.600 389.400 ;
        RECT 260.700 377.400 264.300 378.600 ;
        RECT 239.700 370.050 240.600 377.400 ;
        RECT 263.400 370.050 264.300 377.400 ;
        RECT 280.950 370.950 283.050 373.050 ;
        RECT 236.100 367.050 237.900 368.850 ;
        RECT 238.950 367.950 241.050 370.050 ;
        RECT 235.950 364.950 238.050 367.050 ;
        RECT 230.550 356.550 235.050 358.050 ;
        RECT 239.700 357.600 240.600 367.950 ;
        RECT 242.100 367.050 243.900 368.850 ;
        RECT 260.100 367.050 261.900 368.850 ;
        RECT 262.950 367.950 265.050 370.050 ;
        RECT 281.100 369.150 282.900 370.950 ;
        RECT 284.400 370.050 285.600 383.400 ;
        RECT 292.950 373.950 295.050 376.050 ;
        RECT 286.950 370.950 289.050 373.050 ;
        RECT 241.950 364.950 244.050 367.050 ;
        RECT 259.950 364.950 262.050 367.050 ;
        RECT 263.400 357.600 264.300 367.950 ;
        RECT 266.100 367.050 267.900 368.850 ;
        RECT 283.950 367.950 286.050 370.050 ;
        RECT 287.100 369.150 288.900 370.950 ;
        RECT 265.950 364.950 268.050 367.050 ;
        RECT 284.400 362.700 285.600 367.950 ;
        RECT 281.400 361.800 285.600 362.700 ;
        RECT 231.000 355.950 235.050 356.550 ;
        RECT 239.400 354.600 241.200 357.600 ;
        RECT 262.800 354.600 264.600 357.600 ;
        RECT 281.400 354.600 283.200 361.800 ;
        RECT 293.550 358.050 294.450 373.950 ;
        RECT 299.100 370.050 300.900 371.850 ;
        RECT 301.950 370.950 304.050 373.050 ;
        RECT 298.950 367.950 301.050 370.050 ;
        RECT 302.100 369.150 303.900 370.950 ;
        RECT 304.950 370.050 306.150 383.400 ;
        RECT 316.950 379.950 319.050 382.050 ;
        RECT 307.950 370.950 310.050 373.050 ;
        RECT 304.950 367.950 307.050 370.050 ;
        RECT 308.100 369.150 309.900 370.950 ;
        RECT 305.850 363.750 307.050 367.950 ;
        RECT 317.550 367.050 318.450 379.950 ;
        RECT 322.950 370.950 325.050 373.050 ;
        RECT 323.100 369.150 324.900 370.950 ;
        RECT 326.400 370.050 327.600 383.400 ;
        RECT 328.950 370.950 331.050 373.050 ;
        RECT 346.950 370.950 349.050 373.050 ;
        RECT 325.950 367.950 328.050 370.050 ;
        RECT 329.100 369.150 330.900 370.950 ;
        RECT 347.100 369.150 348.900 370.950 ;
        RECT 350.400 370.050 351.600 383.400 ;
        RECT 368.700 378.600 370.500 389.400 ;
        RECT 368.700 377.400 372.300 378.600 ;
        RECT 388.800 377.400 390.600 389.400 ;
        RECT 391.800 378.300 393.600 389.400 ;
        RECT 397.800 378.300 399.600 389.400 ;
        RECT 391.800 377.400 399.600 378.300 ;
        RECT 401.550 377.400 403.350 389.400 ;
        RECT 409.050 383.400 410.850 389.400 ;
        RECT 406.950 381.300 410.850 383.400 ;
        RECT 416.850 382.500 418.650 389.400 ;
        RECT 424.650 383.400 426.450 389.400 ;
        RECT 425.250 382.500 426.450 383.400 ;
        RECT 415.950 381.450 422.550 382.500 ;
        RECT 415.950 380.700 417.750 381.450 ;
        RECT 420.750 380.700 422.550 381.450 ;
        RECT 425.250 380.400 430.050 382.500 ;
        RECT 408.150 378.600 410.850 380.400 ;
        RECT 411.750 379.800 413.550 380.400 ;
        RECT 411.750 378.900 418.050 379.800 ;
        RECT 425.250 379.500 426.450 380.400 ;
        RECT 411.750 378.600 413.550 378.900 ;
        RECT 409.950 377.700 410.850 378.600 ;
        RECT 352.950 370.950 355.050 373.050 ;
        RECT 349.950 367.950 352.050 370.050 ;
        RECT 353.100 369.150 354.900 370.950 ;
        RECT 371.400 370.050 372.300 377.400 ;
        RECT 389.400 370.050 390.600 377.400 ;
        RECT 391.950 370.950 394.050 373.050 ;
        RECT 316.950 364.950 319.050 367.050 ;
        RECT 305.850 362.700 309.600 363.750 ;
        RECT 299.400 359.700 307.200 361.050 ;
        RECT 292.950 355.950 295.050 358.050 ;
        RECT 299.400 354.600 301.200 359.700 ;
        RECT 305.400 354.600 307.200 359.700 ;
        RECT 308.400 360.600 309.600 362.700 ;
        RECT 326.400 362.700 327.600 367.950 ;
        RECT 350.400 362.700 351.600 367.950 ;
        RECT 368.100 367.050 369.900 368.850 ;
        RECT 370.950 367.950 373.050 370.050 ;
        RECT 367.950 364.950 370.050 367.050 ;
        RECT 326.400 361.800 330.600 362.700 ;
        RECT 308.400 354.600 310.200 360.600 ;
        RECT 328.800 354.600 330.600 361.800 ;
        RECT 347.400 361.800 351.600 362.700 ;
        RECT 347.400 354.600 349.200 361.800 ;
        RECT 371.400 357.600 372.300 367.950 ;
        RECT 374.100 367.050 375.900 368.850 ;
        RECT 388.950 367.950 391.050 370.050 ;
        RECT 392.100 369.150 393.900 370.950 ;
        RECT 395.100 370.050 396.900 371.850 ;
        RECT 397.950 370.950 400.050 373.050 ;
        RECT 394.950 367.950 397.050 370.050 ;
        RECT 398.100 369.150 399.900 370.950 ;
        RECT 401.550 370.050 402.750 377.400 ;
        RECT 406.950 376.800 409.050 377.700 ;
        RECT 409.950 376.800 415.050 377.700 ;
        RECT 404.850 375.600 409.050 376.800 ;
        RECT 403.950 373.800 405.750 375.600 ;
        RECT 401.550 369.750 406.050 370.050 ;
        RECT 401.550 367.950 407.850 369.750 ;
        RECT 373.950 364.950 376.050 367.050 ;
        RECT 389.400 360.600 390.600 367.950 ;
        RECT 401.550 360.600 402.750 367.950 ;
        RECT 414.150 364.200 415.050 376.800 ;
        RECT 417.150 376.800 418.050 378.900 ;
        RECT 418.950 378.300 426.450 379.500 ;
        RECT 418.950 377.700 420.750 378.300 ;
        RECT 433.050 377.400 434.850 389.400 ;
        RECT 451.800 383.400 453.600 389.400 ;
        RECT 417.150 376.500 425.550 376.800 ;
        RECT 433.950 376.500 434.850 377.400 ;
        RECT 417.150 375.900 434.850 376.500 ;
        RECT 423.750 375.300 434.850 375.900 ;
        RECT 423.750 375.000 425.550 375.300 ;
        RECT 421.950 368.400 424.050 370.050 ;
        RECT 421.950 367.200 429.900 368.400 ;
        RECT 430.950 367.950 433.050 370.050 ;
        RECT 428.100 366.600 429.900 367.200 ;
        RECT 431.100 366.150 432.900 367.950 ;
        RECT 425.100 365.400 426.900 366.000 ;
        RECT 431.100 365.400 432.000 366.150 ;
        RECT 425.100 364.200 432.000 365.400 ;
        RECT 414.150 363.000 426.150 364.200 ;
        RECT 414.150 362.400 415.950 363.000 ;
        RECT 425.100 361.200 426.150 363.000 ;
        RECT 389.400 359.400 394.500 360.600 ;
        RECT 370.800 354.600 372.600 357.600 ;
        RECT 392.700 354.600 394.500 359.400 ;
        RECT 401.550 354.600 403.350 360.600 ;
        RECT 406.950 359.700 409.050 360.600 ;
        RECT 406.950 358.500 410.700 359.700 ;
        RECT 421.350 359.550 423.150 360.300 ;
        RECT 409.650 357.600 410.700 358.500 ;
        RECT 418.200 358.500 423.150 359.550 ;
        RECT 424.650 359.400 426.450 361.200 ;
        RECT 433.950 360.600 434.850 375.300 ;
        RECT 446.100 370.050 447.900 371.850 ;
        RECT 448.950 370.950 451.050 373.050 ;
        RECT 445.950 367.950 448.050 370.050 ;
        RECT 449.100 369.150 450.900 370.950 ;
        RECT 451.950 370.050 453.150 383.400 ;
        RECT 470.400 378.300 472.200 389.400 ;
        RECT 476.400 378.300 478.200 389.400 ;
        RECT 470.400 377.400 478.200 378.300 ;
        RECT 479.400 377.400 481.200 389.400 ;
        RECT 486.150 377.400 487.950 389.400 ;
        RECT 494.550 383.400 496.350 389.400 ;
        RECT 494.550 382.500 495.750 383.400 ;
        RECT 502.350 382.500 504.150 389.400 ;
        RECT 510.150 383.400 511.950 389.400 ;
        RECT 490.950 380.400 495.750 382.500 ;
        RECT 498.450 381.450 505.050 382.500 ;
        RECT 498.450 380.700 500.250 381.450 ;
        RECT 503.250 380.700 505.050 381.450 ;
        RECT 510.150 381.300 514.050 383.400 ;
        RECT 494.550 379.500 495.750 380.400 ;
        RECT 507.450 379.800 509.250 380.400 ;
        RECT 494.550 378.300 502.050 379.500 ;
        RECT 500.250 377.700 502.050 378.300 ;
        RECT 502.950 378.900 509.250 379.800 ;
        RECT 454.950 370.950 457.050 373.050 ;
        RECT 469.950 370.950 472.050 373.050 ;
        RECT 451.950 367.950 454.050 370.050 ;
        RECT 455.100 369.150 456.900 370.950 ;
        RECT 470.100 369.150 471.900 370.950 ;
        RECT 473.100 370.050 474.900 371.850 ;
        RECT 475.950 370.950 478.050 373.050 ;
        RECT 472.950 367.950 475.050 370.050 ;
        RECT 476.100 369.150 477.900 370.950 ;
        RECT 479.400 370.050 480.600 377.400 ;
        RECT 486.150 376.500 487.050 377.400 ;
        RECT 502.950 376.800 503.850 378.900 ;
        RECT 507.450 378.600 509.250 378.900 ;
        RECT 510.150 378.600 512.850 380.400 ;
        RECT 510.150 377.700 511.050 378.600 ;
        RECT 495.450 376.500 503.850 376.800 ;
        RECT 486.150 375.900 503.850 376.500 ;
        RECT 505.950 376.800 511.050 377.700 ;
        RECT 511.950 376.800 514.050 377.700 ;
        RECT 517.650 377.400 519.450 389.400 ;
        RECT 520.950 385.950 523.050 388.050 ;
        RECT 486.150 375.300 497.250 375.900 ;
        RECT 478.950 367.950 481.050 370.050 ;
        RECT 452.850 363.750 454.050 367.950 ;
        RECT 452.850 362.700 456.600 363.750 ;
        RECT 427.950 358.500 430.050 360.600 ;
        RECT 418.200 357.600 419.250 358.500 ;
        RECT 427.950 357.600 429.000 358.500 ;
        RECT 409.650 354.600 411.450 357.600 ;
        RECT 417.450 354.600 419.250 357.600 ;
        RECT 425.250 356.700 429.000 357.600 ;
        RECT 425.250 354.600 427.050 356.700 ;
        RECT 433.050 354.600 434.850 360.600 ;
        RECT 446.400 359.700 454.200 361.050 ;
        RECT 446.400 354.600 448.200 359.700 ;
        RECT 452.400 354.600 454.200 359.700 ;
        RECT 455.400 360.600 456.600 362.700 ;
        RECT 479.400 360.600 480.600 367.950 ;
        RECT 455.400 354.600 457.200 360.600 ;
        RECT 475.500 359.400 480.600 360.600 ;
        RECT 486.150 360.600 487.050 375.300 ;
        RECT 495.450 375.000 497.250 375.300 ;
        RECT 487.950 367.950 490.050 370.050 ;
        RECT 496.950 368.400 499.050 370.050 ;
        RECT 488.100 366.150 489.900 367.950 ;
        RECT 491.100 367.200 499.050 368.400 ;
        RECT 491.100 366.600 492.900 367.200 ;
        RECT 489.000 365.400 489.900 366.150 ;
        RECT 494.100 365.400 495.900 366.000 ;
        RECT 489.000 364.200 495.900 365.400 ;
        RECT 505.950 364.200 506.850 376.800 ;
        RECT 511.950 375.600 516.150 376.800 ;
        RECT 515.250 373.800 517.050 375.600 ;
        RECT 518.250 370.050 519.450 377.400 ;
        RECT 521.550 373.050 522.450 385.950 ;
        RECT 535.500 378.600 537.300 389.400 ;
        RECT 556.800 383.400 558.600 389.400 ;
        RECT 578.400 383.400 580.200 389.400 ;
        RECT 599.400 383.400 601.200 389.400 ;
        RECT 533.700 377.400 537.300 378.600 ;
        RECT 520.950 370.950 523.050 373.050 ;
        RECT 533.700 370.050 534.600 377.400 ;
        RECT 553.950 370.950 556.050 373.050 ;
        RECT 514.950 369.750 519.450 370.050 ;
        RECT 513.150 367.950 519.450 369.750 ;
        RECT 494.850 363.000 506.850 364.200 ;
        RECT 494.850 361.200 495.900 363.000 ;
        RECT 505.050 362.400 506.850 363.000 ;
        RECT 475.500 354.600 477.300 359.400 ;
        RECT 486.150 354.600 487.950 360.600 ;
        RECT 490.950 358.500 493.050 360.600 ;
        RECT 494.550 359.400 496.350 361.200 ;
        RECT 518.250 360.600 519.450 367.950 ;
        RECT 530.100 367.050 531.900 368.850 ;
        RECT 532.950 367.950 535.050 370.050 ;
        RECT 554.100 369.150 555.900 370.950 ;
        RECT 557.400 370.050 558.600 383.400 ;
        RECT 559.950 370.950 562.050 373.050 ;
        RECT 574.950 370.950 577.050 373.050 ;
        RECT 529.950 364.950 532.050 367.050 ;
        RECT 497.850 359.550 499.650 360.300 ;
        RECT 511.950 359.700 514.050 360.600 ;
        RECT 497.850 358.500 502.800 359.550 ;
        RECT 492.000 357.600 493.050 358.500 ;
        RECT 501.750 357.600 502.800 358.500 ;
        RECT 510.300 358.500 514.050 359.700 ;
        RECT 510.300 357.600 511.350 358.500 ;
        RECT 492.000 356.700 495.750 357.600 ;
        RECT 493.950 354.600 495.750 356.700 ;
        RECT 501.750 354.600 503.550 357.600 ;
        RECT 509.550 354.600 511.350 357.600 ;
        RECT 517.650 354.600 519.450 360.600 ;
        RECT 533.700 357.600 534.600 367.950 ;
        RECT 536.100 367.050 537.900 368.850 ;
        RECT 556.950 367.950 559.050 370.050 ;
        RECT 560.100 369.150 561.900 370.950 ;
        RECT 575.100 369.150 576.900 370.950 ;
        RECT 578.850 370.050 580.050 383.400 ;
        RECT 599.400 376.050 600.600 383.400 ;
        RECT 605.550 377.400 607.350 389.400 ;
        RECT 613.050 383.400 614.850 389.400 ;
        RECT 610.950 381.300 614.850 383.400 ;
        RECT 620.850 382.500 622.650 389.400 ;
        RECT 628.650 383.400 630.450 389.400 ;
        RECT 629.250 382.500 630.450 383.400 ;
        RECT 619.950 381.450 626.550 382.500 ;
        RECT 619.950 380.700 621.750 381.450 ;
        RECT 624.750 380.700 626.550 381.450 ;
        RECT 629.250 380.400 634.050 382.500 ;
        RECT 612.150 378.600 614.850 380.400 ;
        RECT 615.750 379.800 617.550 380.400 ;
        RECT 615.750 378.900 622.050 379.800 ;
        RECT 629.250 379.500 630.450 380.400 ;
        RECT 615.750 378.600 617.550 378.900 ;
        RECT 613.950 377.700 614.850 378.600 ;
        RECT 580.950 370.950 583.050 373.050 ;
        RECT 577.950 367.950 580.050 370.050 ;
        RECT 581.100 369.150 582.900 370.950 ;
        RECT 584.100 370.050 585.900 371.850 ;
        RECT 596.100 370.050 597.900 371.850 ;
        RECT 598.950 370.950 601.050 376.050 ;
        RECT 583.950 367.950 586.050 370.050 ;
        RECT 595.950 367.950 598.050 370.050 ;
        RECT 535.950 364.950 538.050 367.050 ;
        RECT 557.400 362.700 558.600 367.950 ;
        RECT 577.950 363.750 579.150 367.950 ;
        RECT 554.400 361.800 558.600 362.700 ;
        RECT 575.400 362.700 579.150 363.750 ;
        RECT 533.400 354.600 535.200 357.600 ;
        RECT 554.400 354.600 556.200 361.800 ;
        RECT 575.400 360.600 576.600 362.700 ;
        RECT 574.800 354.600 576.600 360.600 ;
        RECT 577.800 359.700 585.600 361.050 ;
        RECT 577.800 354.600 579.600 359.700 ;
        RECT 583.800 354.600 585.600 359.700 ;
        RECT 599.400 357.600 600.600 370.950 ;
        RECT 605.550 370.050 606.750 377.400 ;
        RECT 610.950 376.800 613.050 377.700 ;
        RECT 613.950 376.800 619.050 377.700 ;
        RECT 608.850 375.600 613.050 376.800 ;
        RECT 607.950 373.800 609.750 375.600 ;
        RECT 605.550 369.750 610.050 370.050 ;
        RECT 605.550 367.950 611.850 369.750 ;
        RECT 605.550 360.600 606.750 367.950 ;
        RECT 618.150 364.200 619.050 376.800 ;
        RECT 621.150 376.800 622.050 378.900 ;
        RECT 622.950 378.300 630.450 379.500 ;
        RECT 622.950 377.700 624.750 378.300 ;
        RECT 637.050 377.400 638.850 389.400 ;
        RECT 621.150 376.500 629.550 376.800 ;
        RECT 637.950 376.500 638.850 377.400 ;
        RECT 640.950 376.950 643.050 379.050 ;
        RECT 654.900 377.400 658.200 389.400 ;
        RECT 682.500 378.600 684.300 389.400 ;
        RECT 680.700 377.400 684.300 378.600 ;
        RECT 621.150 375.900 638.850 376.500 ;
        RECT 627.750 375.300 638.850 375.900 ;
        RECT 627.750 375.000 629.550 375.300 ;
        RECT 625.950 368.400 628.050 370.050 ;
        RECT 625.950 367.200 633.900 368.400 ;
        RECT 634.950 367.950 637.050 370.050 ;
        RECT 632.100 366.600 633.900 367.200 ;
        RECT 635.100 366.150 636.900 367.950 ;
        RECT 629.100 365.400 630.900 366.000 ;
        RECT 635.100 365.400 636.000 366.150 ;
        RECT 629.100 364.200 636.000 365.400 ;
        RECT 618.150 363.000 630.150 364.200 ;
        RECT 618.150 362.400 619.950 363.000 ;
        RECT 629.100 361.200 630.150 363.000 ;
        RECT 599.400 354.600 601.200 357.600 ;
        RECT 605.550 354.600 607.350 360.600 ;
        RECT 610.950 359.700 613.050 360.600 ;
        RECT 610.950 358.500 614.700 359.700 ;
        RECT 625.350 359.550 627.150 360.300 ;
        RECT 613.650 357.600 614.700 358.500 ;
        RECT 622.200 358.500 627.150 359.550 ;
        RECT 628.650 359.400 630.450 361.200 ;
        RECT 637.950 360.600 638.850 375.300 ;
        RECT 641.550 361.050 642.450 376.950 ;
        RECT 650.100 370.050 651.900 371.850 ;
        RECT 652.950 370.950 655.050 373.050 ;
        RECT 649.950 367.950 652.050 370.050 ;
        RECT 653.100 369.150 654.900 370.950 ;
        RECT 656.100 370.050 657.300 377.400 ;
        RECT 658.950 370.950 661.050 373.050 ;
        RECT 655.950 367.950 658.050 370.050 ;
        RECT 659.100 369.150 660.900 370.950 ;
        RECT 662.100 370.050 663.900 371.850 ;
        RECT 680.700 370.050 681.600 377.400 ;
        RECT 691.950 376.950 694.050 379.050 ;
        RECT 698.400 378.300 700.200 389.400 ;
        RECT 704.400 378.300 706.200 389.400 ;
        RECT 698.400 377.400 706.200 378.300 ;
        RECT 707.400 377.400 709.200 389.400 ;
        RECT 722.400 378.300 724.200 389.400 ;
        RECT 728.400 378.300 730.200 389.400 ;
        RECT 722.400 377.400 730.200 378.300 ;
        RECT 731.400 377.400 733.200 389.400 ;
        RECT 738.150 377.400 739.950 389.400 ;
        RECT 746.550 383.400 748.350 389.400 ;
        RECT 746.550 382.500 747.750 383.400 ;
        RECT 754.350 382.500 756.150 389.400 ;
        RECT 762.150 383.400 763.950 389.400 ;
        RECT 742.950 380.400 747.750 382.500 ;
        RECT 750.450 381.450 757.050 382.500 ;
        RECT 750.450 380.700 752.250 381.450 ;
        RECT 755.250 380.700 757.050 381.450 ;
        RECT 762.150 381.300 766.050 383.400 ;
        RECT 746.550 379.500 747.750 380.400 ;
        RECT 759.450 379.800 761.250 380.400 ;
        RECT 746.550 378.300 754.050 379.500 ;
        RECT 752.250 377.700 754.050 378.300 ;
        RECT 754.950 378.900 761.250 379.800 ;
        RECT 661.950 367.950 664.050 370.050 ;
        RECT 655.950 363.300 657.300 367.950 ;
        RECT 677.100 367.050 678.900 368.850 ;
        RECT 679.950 367.950 682.050 370.050 ;
        RECT 676.950 364.950 679.050 367.050 ;
        RECT 655.950 362.100 660.600 363.300 ;
        RECT 631.950 358.500 634.050 360.600 ;
        RECT 622.200 357.600 623.250 358.500 ;
        RECT 631.950 357.600 633.000 358.500 ;
        RECT 613.650 354.600 615.450 357.600 ;
        RECT 621.450 354.600 623.250 357.600 ;
        RECT 629.250 356.700 633.000 357.600 ;
        RECT 629.250 354.600 631.050 356.700 ;
        RECT 637.050 354.600 638.850 360.600 ;
        RECT 640.950 358.950 643.050 361.050 ;
        RECT 650.400 360.000 658.200 360.900 ;
        RECT 659.700 360.600 660.600 362.100 ;
        RECT 650.400 354.600 652.200 360.000 ;
        RECT 656.400 355.500 658.200 360.000 ;
        RECT 659.400 356.400 661.200 360.600 ;
        RECT 662.400 355.500 664.200 360.600 ;
        RECT 680.700 357.600 681.600 367.950 ;
        RECT 683.100 367.050 684.900 368.850 ;
        RECT 682.950 364.950 685.050 367.050 ;
        RECT 692.550 361.050 693.450 376.950 ;
        RECT 697.950 370.950 700.050 373.050 ;
        RECT 698.100 369.150 699.900 370.950 ;
        RECT 701.100 370.050 702.900 371.850 ;
        RECT 703.950 370.950 706.050 373.050 ;
        RECT 700.950 367.950 703.050 370.050 ;
        RECT 704.100 369.150 705.900 370.950 ;
        RECT 707.400 370.050 708.600 377.400 ;
        RECT 721.950 370.950 724.050 373.050 ;
        RECT 706.950 367.950 709.050 370.050 ;
        RECT 722.100 369.150 723.900 370.950 ;
        RECT 725.100 370.050 726.900 371.850 ;
        RECT 727.950 370.950 730.050 373.050 ;
        RECT 724.950 367.950 727.050 370.050 ;
        RECT 728.100 369.150 729.900 370.950 ;
        RECT 731.400 370.050 732.600 377.400 ;
        RECT 738.150 376.500 739.050 377.400 ;
        RECT 754.950 376.800 755.850 378.900 ;
        RECT 759.450 378.600 761.250 378.900 ;
        RECT 762.150 378.600 764.850 380.400 ;
        RECT 762.150 377.700 763.050 378.600 ;
        RECT 747.450 376.500 755.850 376.800 ;
        RECT 738.150 375.900 755.850 376.500 ;
        RECT 757.950 376.800 763.050 377.700 ;
        RECT 763.950 376.800 766.050 377.700 ;
        RECT 769.650 377.400 771.450 389.400 ;
        RECT 782.400 378.600 784.200 389.400 ;
        RECT 788.400 388.500 796.200 389.400 ;
        RECT 788.400 378.600 790.200 388.500 ;
        RECT 782.400 377.700 790.200 378.600 ;
        RECT 738.150 375.300 749.250 375.900 ;
        RECT 730.950 367.950 733.050 370.050 ;
        RECT 691.950 358.950 694.050 361.050 ;
        RECT 707.400 360.600 708.600 367.950 ;
        RECT 731.400 360.600 732.600 367.950 ;
        RECT 703.500 359.400 708.600 360.600 ;
        RECT 727.500 359.400 732.600 360.600 ;
        RECT 738.150 360.600 739.050 375.300 ;
        RECT 747.450 375.000 749.250 375.300 ;
        RECT 739.950 367.950 742.050 370.050 ;
        RECT 748.950 368.400 751.050 370.050 ;
        RECT 740.100 366.150 741.900 367.950 ;
        RECT 743.100 367.200 751.050 368.400 ;
        RECT 743.100 366.600 744.900 367.200 ;
        RECT 741.000 365.400 741.900 366.150 ;
        RECT 746.100 365.400 747.900 366.000 ;
        RECT 741.000 364.200 747.900 365.400 ;
        RECT 757.950 364.200 758.850 376.800 ;
        RECT 763.950 375.600 768.150 376.800 ;
        RECT 767.250 373.800 769.050 375.600 ;
        RECT 770.250 370.050 771.450 377.400 ;
        RECT 791.400 376.500 793.200 387.600 ;
        RECT 794.400 377.400 796.200 388.500 ;
        RECT 812.400 383.400 814.200 389.400 ;
        RECT 826.950 385.950 829.050 388.050 ;
        RECT 788.100 375.600 793.200 376.500 ;
        RECT 788.100 370.050 789.000 375.600 ;
        RECT 808.950 370.950 811.050 373.050 ;
        RECT 766.950 369.750 771.450 370.050 ;
        RECT 765.150 367.950 771.450 369.750 ;
        RECT 781.950 367.950 784.050 370.050 ;
        RECT 746.850 363.000 758.850 364.200 ;
        RECT 746.850 361.200 747.900 363.000 ;
        RECT 757.050 362.400 758.850 363.000 ;
        RECT 656.400 354.600 664.200 355.500 ;
        RECT 680.400 354.600 682.200 357.600 ;
        RECT 703.500 354.600 705.300 359.400 ;
        RECT 727.500 354.600 729.300 359.400 ;
        RECT 738.150 354.600 739.950 360.600 ;
        RECT 742.950 358.500 745.050 360.600 ;
        RECT 746.550 359.400 748.350 361.200 ;
        RECT 770.250 360.600 771.450 367.950 ;
        RECT 782.100 366.150 783.900 367.950 ;
        RECT 785.100 367.050 786.900 368.850 ;
        RECT 787.950 367.950 790.050 370.050 ;
        RECT 784.950 364.950 787.050 367.050 ;
        RECT 787.950 360.600 789.000 367.950 ;
        RECT 791.100 367.050 792.900 368.850 ;
        RECT 793.950 367.950 796.050 370.050 ;
        RECT 809.100 369.150 810.900 370.950 ;
        RECT 812.400 370.050 813.600 383.400 ;
        RECT 814.950 370.950 817.050 373.050 ;
        RECT 811.950 367.950 814.050 370.050 ;
        RECT 815.100 369.150 816.900 370.950 ;
        RECT 790.950 364.950 793.050 367.050 ;
        RECT 794.100 366.150 795.900 367.950 ;
        RECT 812.400 362.700 813.600 367.950 ;
        RECT 812.400 361.800 816.600 362.700 ;
        RECT 749.850 359.550 751.650 360.300 ;
        RECT 763.950 359.700 766.050 360.600 ;
        RECT 749.850 358.500 754.800 359.550 ;
        RECT 744.000 357.600 745.050 358.500 ;
        RECT 753.750 357.600 754.800 358.500 ;
        RECT 762.300 358.500 766.050 359.700 ;
        RECT 762.300 357.600 763.350 358.500 ;
        RECT 744.000 356.700 747.750 357.600 ;
        RECT 745.950 354.600 747.750 356.700 ;
        RECT 753.750 354.600 755.550 357.600 ;
        RECT 761.550 354.600 763.350 357.600 ;
        RECT 769.650 354.600 771.450 360.600 ;
        RECT 787.200 354.600 789.000 360.600 ;
        RECT 814.800 354.600 816.600 361.800 ;
        RECT 827.550 358.050 828.450 385.950 ;
        RECT 834.300 378.900 836.100 389.400 ;
        RECT 833.700 377.400 836.100 378.900 ;
        RECT 841.800 377.400 843.600 389.400 ;
        RECT 859.800 383.400 861.600 389.400 ;
        RECT 833.700 370.050 835.050 377.400 ;
        RECT 842.400 375.900 843.600 377.400 ;
        RECT 832.950 367.950 835.050 370.050 ;
        RECT 836.400 374.700 843.600 375.900 ;
        RECT 836.400 374.100 838.200 374.700 ;
        RECT 832.950 360.600 834.000 367.950 ;
        RECT 836.400 363.600 837.300 374.100 ;
        RECT 839.100 370.050 840.900 371.850 ;
        RECT 841.950 370.950 844.050 373.050 ;
        RECT 838.950 367.950 841.050 370.050 ;
        RECT 842.100 369.150 843.900 370.950 ;
        RECT 854.100 370.050 855.900 371.850 ;
        RECT 856.950 370.950 859.050 373.050 ;
        RECT 853.950 367.950 856.050 370.050 ;
        RECT 857.100 369.150 858.900 370.950 ;
        RECT 859.950 370.050 861.150 383.400 ;
        RECT 870.150 377.400 871.950 389.400 ;
        RECT 878.550 383.400 880.350 389.400 ;
        RECT 878.550 382.500 879.750 383.400 ;
        RECT 886.350 382.500 888.150 389.400 ;
        RECT 894.150 383.400 895.950 389.400 ;
        RECT 874.950 380.400 879.750 382.500 ;
        RECT 882.450 381.450 889.050 382.500 ;
        RECT 882.450 380.700 884.250 381.450 ;
        RECT 887.250 380.700 889.050 381.450 ;
        RECT 894.150 381.300 898.050 383.400 ;
        RECT 878.550 379.500 879.750 380.400 ;
        RECT 891.450 379.800 893.250 380.400 ;
        RECT 878.550 378.300 886.050 379.500 ;
        RECT 884.250 377.700 886.050 378.300 ;
        RECT 886.950 378.900 893.250 379.800 ;
        RECT 870.150 376.500 871.050 377.400 ;
        RECT 886.950 376.800 887.850 378.900 ;
        RECT 891.450 378.600 893.250 378.900 ;
        RECT 894.150 378.600 896.850 380.400 ;
        RECT 894.150 377.700 895.050 378.600 ;
        RECT 879.450 376.500 887.850 376.800 ;
        RECT 870.150 375.900 887.850 376.500 ;
        RECT 889.950 376.800 895.050 377.700 ;
        RECT 895.950 376.800 898.050 377.700 ;
        RECT 901.650 377.400 903.450 389.400 ;
        RECT 870.150 375.300 881.250 375.900 ;
        RECT 862.950 370.950 865.050 373.050 ;
        RECT 859.950 367.950 862.050 370.050 ;
        RECT 863.100 369.150 864.900 370.950 ;
        RECT 860.850 363.750 862.050 367.950 ;
        RECT 836.400 362.700 838.200 363.600 ;
        RECT 860.850 362.700 864.600 363.750 ;
        RECT 836.400 361.800 839.700 362.700 ;
        RECT 826.950 355.950 829.050 358.050 ;
        RECT 832.800 354.600 834.600 360.600 ;
        RECT 838.800 357.600 839.700 361.800 ;
        RECT 854.400 359.700 862.200 361.050 ;
        RECT 838.800 354.600 840.600 357.600 ;
        RECT 854.400 354.600 856.200 359.700 ;
        RECT 860.400 354.600 862.200 359.700 ;
        RECT 863.400 360.600 864.600 362.700 ;
        RECT 870.150 360.600 871.050 375.300 ;
        RECT 879.450 375.000 881.250 375.300 ;
        RECT 871.950 367.950 874.050 370.050 ;
        RECT 880.950 368.400 883.050 370.050 ;
        RECT 872.100 366.150 873.900 367.950 ;
        RECT 875.100 367.200 883.050 368.400 ;
        RECT 875.100 366.600 876.900 367.200 ;
        RECT 873.000 365.400 873.900 366.150 ;
        RECT 878.100 365.400 879.900 366.000 ;
        RECT 873.000 364.200 879.900 365.400 ;
        RECT 889.950 364.200 890.850 376.800 ;
        RECT 895.950 375.600 900.150 376.800 ;
        RECT 899.250 373.800 901.050 375.600 ;
        RECT 902.250 370.050 903.450 377.400 ;
        RECT 898.950 369.750 903.450 370.050 ;
        RECT 897.150 367.950 903.450 369.750 ;
        RECT 878.850 363.000 890.850 364.200 ;
        RECT 878.850 361.200 879.900 363.000 ;
        RECT 889.050 362.400 890.850 363.000 ;
        RECT 863.400 354.600 865.200 360.600 ;
        RECT 870.150 354.600 871.950 360.600 ;
        RECT 874.950 358.500 877.050 360.600 ;
        RECT 878.550 359.400 880.350 361.200 ;
        RECT 902.250 360.600 903.450 367.950 ;
        RECT 881.850 359.550 883.650 360.300 ;
        RECT 895.950 359.700 898.050 360.600 ;
        RECT 881.850 358.500 886.800 359.550 ;
        RECT 876.000 357.600 877.050 358.500 ;
        RECT 885.750 357.600 886.800 358.500 ;
        RECT 894.300 358.500 898.050 359.700 ;
        RECT 894.300 357.600 895.350 358.500 ;
        RECT 876.000 356.700 879.750 357.600 ;
        RECT 877.950 354.600 879.750 356.700 ;
        RECT 885.750 354.600 887.550 357.600 ;
        RECT 893.550 354.600 895.350 357.600 ;
        RECT 901.650 354.600 903.450 360.600 ;
        RECT 14.400 347.400 16.200 350.400 ;
        RECT 31.800 347.400 33.600 350.400 ;
        RECT 49.800 347.400 51.600 350.400 ;
        RECT 70.800 347.400 72.600 350.400 ;
        RECT 91.800 347.400 93.600 350.400 ;
        RECT 109.800 347.400 111.600 350.400 ;
        RECT 10.950 334.950 13.050 337.050 ;
        RECT 11.100 333.150 12.900 334.950 ;
        RECT 14.400 334.050 15.600 347.400 ;
        RECT 32.400 334.050 33.600 347.400 ;
        RECT 34.950 334.950 37.050 337.050 ;
        RECT 13.950 328.950 16.050 334.050 ;
        RECT 31.950 328.950 34.050 334.050 ;
        RECT 35.100 333.150 36.900 334.950 ;
        RECT 50.400 334.050 51.600 347.400 ;
        RECT 67.950 337.950 70.050 340.050 ;
        RECT 52.950 334.950 55.050 337.050 ;
        RECT 68.100 336.150 69.900 337.950 ;
        RECT 71.400 337.050 72.300 347.400 ;
        RECT 82.950 340.950 85.050 343.050 ;
        RECT 73.950 337.950 76.050 340.050 ;
        RECT 70.950 334.950 73.050 337.050 ;
        RECT 74.100 336.150 75.900 337.950 ;
        RECT 49.950 328.950 52.050 334.050 ;
        RECT 53.100 333.150 54.900 334.950 ;
        RECT 14.400 321.600 15.600 328.950 ;
        RECT 32.400 321.600 33.600 328.950 ;
        RECT 50.400 321.600 51.600 328.950 ;
        RECT 71.400 327.600 72.300 334.950 ;
        RECT 14.400 315.600 16.200 321.600 ;
        RECT 31.800 315.600 33.600 321.600 ;
        RECT 49.800 315.600 51.600 321.600 ;
        RECT 68.700 326.400 72.300 327.600 ;
        RECT 68.700 315.600 70.500 326.400 ;
        RECT 83.550 325.050 84.450 340.950 ;
        RECT 88.950 337.950 91.050 340.050 ;
        RECT 89.100 336.150 90.900 337.950 ;
        RECT 92.400 337.050 93.300 347.400 ;
        RECT 94.950 337.950 97.050 340.050 ;
        RECT 91.950 334.950 94.050 337.050 ;
        RECT 95.100 336.150 96.900 337.950 ;
        RECT 92.400 327.600 93.300 334.950 ;
        RECT 110.400 334.050 111.600 347.400 ;
        RECT 116.550 344.400 118.350 350.400 ;
        RECT 124.650 347.400 126.450 350.400 ;
        RECT 132.450 347.400 134.250 350.400 ;
        RECT 140.250 348.300 142.050 350.400 ;
        RECT 140.250 347.400 144.000 348.300 ;
        RECT 124.650 346.500 125.700 347.400 ;
        RECT 121.950 345.300 125.700 346.500 ;
        RECT 133.200 346.500 134.250 347.400 ;
        RECT 142.950 346.500 144.000 347.400 ;
        RECT 133.200 345.450 138.150 346.500 ;
        RECT 121.950 344.400 124.050 345.300 ;
        RECT 136.350 344.700 138.150 345.450 ;
        RECT 116.550 337.050 117.750 344.400 ;
        RECT 139.650 343.800 141.450 345.600 ;
        RECT 142.950 344.400 145.050 346.500 ;
        RECT 148.050 344.400 149.850 350.400 ;
        RECT 163.800 344.400 165.600 350.400 ;
        RECT 129.150 342.000 130.950 342.600 ;
        RECT 140.100 342.000 141.150 343.800 ;
        RECT 129.150 340.800 141.150 342.000 ;
        RECT 112.950 334.950 115.050 337.050 ;
        RECT 116.550 335.250 122.850 337.050 ;
        RECT 116.550 334.950 121.050 335.250 ;
        RECT 109.950 328.950 112.050 334.050 ;
        RECT 113.100 333.150 114.900 334.950 ;
        RECT 89.700 326.400 93.300 327.600 ;
        RECT 82.950 322.950 85.050 325.050 ;
        RECT 89.700 315.600 91.500 326.400 ;
        RECT 110.400 321.600 111.600 328.950 ;
        RECT 109.800 315.600 111.600 321.600 ;
        RECT 116.550 327.600 117.750 334.950 ;
        RECT 118.950 329.400 120.750 331.200 ;
        RECT 119.850 328.200 124.050 329.400 ;
        RECT 129.150 328.200 130.050 340.800 ;
        RECT 140.100 339.600 147.000 340.800 ;
        RECT 140.100 339.000 141.900 339.600 ;
        RECT 146.100 338.850 147.000 339.600 ;
        RECT 143.100 337.800 144.900 338.400 ;
        RECT 136.950 336.600 144.900 337.800 ;
        RECT 146.100 337.050 147.900 338.850 ;
        RECT 136.950 334.950 139.050 336.600 ;
        RECT 145.950 334.950 148.050 337.050 ;
        RECT 138.750 329.700 140.550 330.000 ;
        RECT 148.950 329.700 149.850 344.400 ;
        RECT 164.400 342.300 165.600 344.400 ;
        RECT 166.800 345.300 168.600 350.400 ;
        RECT 172.800 345.300 174.600 350.400 ;
        RECT 166.800 343.950 174.600 345.300 ;
        RECT 177.150 344.400 178.950 350.400 ;
        RECT 184.950 348.300 186.750 350.400 ;
        RECT 183.000 347.400 186.750 348.300 ;
        RECT 192.750 347.400 194.550 350.400 ;
        RECT 200.550 347.400 202.350 350.400 ;
        RECT 183.000 346.500 184.050 347.400 ;
        RECT 192.750 346.500 193.800 347.400 ;
        RECT 181.950 344.400 184.050 346.500 ;
        RECT 164.400 341.250 168.150 342.300 ;
        RECT 166.950 337.050 168.150 341.250 ;
        RECT 164.100 334.050 165.900 335.850 ;
        RECT 166.950 334.950 169.050 337.050 ;
        RECT 163.950 331.950 166.050 334.050 ;
        RECT 138.750 329.100 149.850 329.700 ;
        RECT 116.550 315.600 118.350 327.600 ;
        RECT 121.950 327.300 124.050 328.200 ;
        RECT 124.950 327.300 130.050 328.200 ;
        RECT 132.150 328.500 149.850 329.100 ;
        RECT 132.150 328.200 140.550 328.500 ;
        RECT 124.950 326.400 125.850 327.300 ;
        RECT 123.150 324.600 125.850 326.400 ;
        RECT 126.750 326.100 128.550 326.400 ;
        RECT 132.150 326.100 133.050 328.200 ;
        RECT 148.950 327.600 149.850 328.500 ;
        RECT 126.750 325.200 133.050 326.100 ;
        RECT 133.950 326.700 135.750 327.300 ;
        RECT 133.950 325.500 141.450 326.700 ;
        RECT 126.750 324.600 128.550 325.200 ;
        RECT 140.250 324.600 141.450 325.500 ;
        RECT 121.950 321.600 125.850 323.700 ;
        RECT 130.950 323.550 132.750 324.300 ;
        RECT 135.750 323.550 137.550 324.300 ;
        RECT 130.950 322.500 137.550 323.550 ;
        RECT 140.250 322.500 145.050 324.600 ;
        RECT 124.050 315.600 125.850 321.600 ;
        RECT 131.850 315.600 133.650 322.500 ;
        RECT 140.250 321.600 141.450 322.500 ;
        RECT 139.650 315.600 141.450 321.600 ;
        RECT 148.050 315.600 149.850 327.600 ;
        RECT 167.850 321.600 169.050 334.950 ;
        RECT 170.100 334.050 171.900 335.850 ;
        RECT 172.950 334.950 175.050 337.050 ;
        RECT 169.950 331.950 172.050 334.050 ;
        RECT 173.100 333.150 174.900 334.950 ;
        RECT 177.150 329.700 178.050 344.400 ;
        RECT 185.550 343.800 187.350 345.600 ;
        RECT 188.850 345.450 193.800 346.500 ;
        RECT 201.300 346.500 202.350 347.400 ;
        RECT 188.850 344.700 190.650 345.450 ;
        RECT 201.300 345.300 205.050 346.500 ;
        RECT 202.950 344.400 205.050 345.300 ;
        RECT 208.650 344.400 210.450 350.400 ;
        RECT 185.850 342.000 186.900 343.800 ;
        RECT 196.050 342.000 197.850 342.600 ;
        RECT 185.850 340.800 197.850 342.000 ;
        RECT 180.000 339.600 186.900 340.800 ;
        RECT 180.000 338.850 180.900 339.600 ;
        RECT 185.100 339.000 186.900 339.600 ;
        RECT 179.100 337.050 180.900 338.850 ;
        RECT 182.100 337.800 183.900 338.400 ;
        RECT 178.950 334.950 181.050 337.050 ;
        RECT 182.100 336.600 190.050 337.800 ;
        RECT 187.950 334.950 190.050 336.600 ;
        RECT 186.450 329.700 188.250 330.000 ;
        RECT 177.150 329.100 188.250 329.700 ;
        RECT 177.150 328.500 194.850 329.100 ;
        RECT 177.150 327.600 178.050 328.500 ;
        RECT 186.450 328.200 194.850 328.500 ;
        RECT 167.400 315.600 169.200 321.600 ;
        RECT 177.150 315.600 178.950 327.600 ;
        RECT 191.250 326.700 193.050 327.300 ;
        RECT 185.550 325.500 193.050 326.700 ;
        RECT 193.950 326.100 194.850 328.200 ;
        RECT 196.950 328.200 197.850 340.800 ;
        RECT 209.250 337.050 210.450 344.400 ;
        RECT 224.400 347.400 226.200 350.400 ;
        RECT 204.150 335.250 210.450 337.050 ;
        RECT 205.950 334.950 210.450 335.250 ;
        RECT 220.950 334.950 223.050 337.050 ;
        RECT 206.250 329.400 208.050 331.200 ;
        RECT 202.950 328.200 207.150 329.400 ;
        RECT 196.950 327.300 202.050 328.200 ;
        RECT 202.950 327.300 205.050 328.200 ;
        RECT 209.250 327.600 210.450 334.950 ;
        RECT 221.100 333.150 222.900 334.950 ;
        RECT 224.400 334.050 225.600 347.400 ;
        RECT 239.400 345.300 241.200 350.400 ;
        RECT 245.400 345.300 247.200 350.400 ;
        RECT 239.400 343.950 247.200 345.300 ;
        RECT 248.400 344.400 250.200 350.400 ;
        RECT 263.400 347.400 265.200 350.400 ;
        RECT 248.400 342.300 249.600 344.400 ;
        RECT 263.400 343.500 264.600 347.400 ;
        RECT 269.700 344.400 271.500 350.400 ;
        RECT 263.400 342.600 269.400 343.500 ;
        RECT 245.850 341.250 249.600 342.300 ;
        RECT 267.150 341.700 269.400 342.600 ;
        RECT 245.850 337.050 247.050 341.250 ;
        RECT 238.950 334.950 241.050 337.050 ;
        RECT 223.950 328.950 226.050 334.050 ;
        RECT 239.100 333.150 240.900 334.950 ;
        RECT 242.100 334.050 243.900 335.850 ;
        RECT 244.950 334.950 247.050 337.050 ;
        RECT 241.950 331.950 244.050 334.050 ;
        RECT 201.150 326.400 202.050 327.300 ;
        RECT 198.450 326.100 200.250 326.400 ;
        RECT 185.550 324.600 186.750 325.500 ;
        RECT 193.950 325.200 200.250 326.100 ;
        RECT 198.450 324.600 200.250 325.200 ;
        RECT 201.150 324.600 203.850 326.400 ;
        RECT 181.950 322.500 186.750 324.600 ;
        RECT 189.450 323.550 191.250 324.300 ;
        RECT 194.250 323.550 196.050 324.300 ;
        RECT 189.450 322.500 196.050 323.550 ;
        RECT 185.550 321.600 186.750 322.500 ;
        RECT 185.550 315.600 187.350 321.600 ;
        RECT 193.350 315.600 195.150 322.500 ;
        RECT 201.150 321.600 205.050 323.700 ;
        RECT 201.150 315.600 202.950 321.600 ;
        RECT 208.650 315.600 210.450 327.600 ;
        RECT 224.400 321.600 225.600 328.950 ;
        RECT 244.950 321.600 246.150 334.950 ;
        RECT 248.100 334.050 249.900 335.850 ;
        RECT 262.950 334.950 265.050 337.050 ;
        RECT 247.950 331.950 250.050 334.050 ;
        RECT 263.100 333.150 264.900 334.950 ;
        RECT 267.150 330.300 268.050 341.700 ;
        RECT 270.300 337.050 271.500 344.400 ;
        RECT 289.800 343.200 291.600 350.400 ;
        RECT 287.400 342.300 291.600 343.200 ;
        RECT 307.500 344.400 309.300 350.400 ;
        RECT 313.800 347.400 315.600 350.400 ;
        RECT 287.400 337.050 288.600 342.300 ;
        RECT 307.500 337.050 308.700 344.400 ;
        RECT 314.400 343.500 315.600 347.400 ;
        RECT 309.600 342.600 315.600 343.500 ;
        RECT 328.500 344.400 330.300 350.400 ;
        RECT 334.800 347.400 336.600 350.400 ;
        RECT 352.800 347.400 354.600 350.400 ;
        RECT 309.600 341.700 311.850 342.600 ;
        RECT 268.950 334.950 271.500 337.050 ;
        RECT 267.150 329.400 269.400 330.300 ;
        RECT 263.400 328.500 269.400 329.400 ;
        RECT 263.400 321.600 264.600 328.500 ;
        RECT 270.300 327.600 271.500 334.950 ;
        RECT 284.100 334.050 285.900 335.850 ;
        RECT 286.950 334.950 289.050 337.050 ;
        RECT 283.950 331.950 286.050 334.050 ;
        RECT 224.400 315.600 226.200 321.600 ;
        RECT 244.800 315.600 246.600 321.600 ;
        RECT 263.400 315.600 265.200 321.600 ;
        RECT 269.700 315.600 271.500 327.600 ;
        RECT 287.400 321.600 288.600 334.950 ;
        RECT 290.100 334.050 291.900 335.850 ;
        RECT 307.500 334.950 310.050 337.050 ;
        RECT 289.950 331.950 292.050 334.050 ;
        RECT 307.500 327.600 308.700 334.950 ;
        RECT 310.950 330.300 311.850 341.700 ;
        RECT 328.500 337.050 329.700 344.400 ;
        RECT 335.400 343.500 336.600 347.400 ;
        RECT 330.600 342.600 336.600 343.500 ;
        RECT 330.600 341.700 332.850 342.600 ;
        RECT 313.950 334.950 316.050 337.050 ;
        RECT 328.500 334.950 331.050 337.050 ;
        RECT 314.100 333.150 315.900 334.950 ;
        RECT 309.600 329.400 311.850 330.300 ;
        RECT 309.600 328.500 315.600 329.400 ;
        RECT 287.400 315.600 289.200 321.600 ;
        RECT 307.500 315.600 309.300 327.600 ;
        RECT 314.400 321.600 315.600 328.500 ;
        RECT 313.800 315.600 315.600 321.600 ;
        RECT 328.500 327.600 329.700 334.950 ;
        RECT 331.950 330.300 332.850 341.700 ;
        RECT 349.950 337.950 352.050 340.050 ;
        RECT 334.950 334.950 337.050 337.050 ;
        RECT 350.100 336.150 351.900 337.950 ;
        RECT 353.400 337.050 354.300 347.400 ;
        RECT 359.550 344.400 361.350 350.400 ;
        RECT 367.650 347.400 369.450 350.400 ;
        RECT 375.450 347.400 377.250 350.400 ;
        RECT 383.250 348.300 385.050 350.400 ;
        RECT 383.250 347.400 387.000 348.300 ;
        RECT 367.650 346.500 368.700 347.400 ;
        RECT 364.950 345.300 368.700 346.500 ;
        RECT 376.200 346.500 377.250 347.400 ;
        RECT 385.950 346.500 387.000 347.400 ;
        RECT 376.200 345.450 381.150 346.500 ;
        RECT 364.950 344.400 367.050 345.300 ;
        RECT 379.350 344.700 381.150 345.450 ;
        RECT 355.950 337.950 358.050 340.050 ;
        RECT 352.950 334.950 355.050 337.050 ;
        RECT 356.100 336.150 357.900 337.950 ;
        RECT 359.550 337.050 360.750 344.400 ;
        RECT 382.650 343.800 384.450 345.600 ;
        RECT 385.950 344.400 388.050 346.500 ;
        RECT 391.050 344.400 392.850 350.400 ;
        RECT 409.800 347.400 411.600 350.400 ;
        RECT 372.150 342.000 373.950 342.600 ;
        RECT 383.100 342.000 384.150 343.800 ;
        RECT 372.150 340.800 384.150 342.000 ;
        RECT 359.550 335.250 365.850 337.050 ;
        RECT 359.550 334.950 364.050 335.250 ;
        RECT 335.100 333.150 336.900 334.950 ;
        RECT 330.600 329.400 332.850 330.300 ;
        RECT 330.600 328.500 336.600 329.400 ;
        RECT 328.500 315.600 330.300 327.600 ;
        RECT 335.400 321.600 336.600 328.500 ;
        RECT 353.400 327.600 354.300 334.950 ;
        RECT 334.800 315.600 336.600 321.600 ;
        RECT 350.700 326.400 354.300 327.600 ;
        RECT 359.550 327.600 360.750 334.950 ;
        RECT 361.950 329.400 363.750 331.200 ;
        RECT 362.850 328.200 367.050 329.400 ;
        RECT 372.150 328.200 373.050 340.800 ;
        RECT 383.100 339.600 390.000 340.800 ;
        RECT 383.100 339.000 384.900 339.600 ;
        RECT 389.100 338.850 390.000 339.600 ;
        RECT 386.100 337.800 387.900 338.400 ;
        RECT 379.950 336.600 387.900 337.800 ;
        RECT 389.100 337.050 390.900 338.850 ;
        RECT 379.950 334.950 382.050 336.600 ;
        RECT 388.950 334.950 391.050 337.050 ;
        RECT 381.750 329.700 383.550 330.000 ;
        RECT 391.950 329.700 392.850 344.400 ;
        RECT 406.950 337.950 409.050 340.050 ;
        RECT 407.100 336.150 408.900 337.950 ;
        RECT 410.400 337.050 411.300 347.400 ;
        RECT 431.700 345.600 433.500 350.400 ;
        RECT 428.400 344.400 433.500 345.600 ;
        RECT 441.150 344.400 442.950 350.400 ;
        RECT 448.950 348.300 450.750 350.400 ;
        RECT 447.000 347.400 450.750 348.300 ;
        RECT 456.750 347.400 458.550 350.400 ;
        RECT 464.550 347.400 466.350 350.400 ;
        RECT 447.000 346.500 448.050 347.400 ;
        RECT 456.750 346.500 457.800 347.400 ;
        RECT 445.950 344.400 448.050 346.500 ;
        RECT 412.950 337.950 415.050 340.050 ;
        RECT 409.950 334.950 412.050 337.050 ;
        RECT 413.100 336.150 414.900 337.950 ;
        RECT 428.400 337.050 429.600 344.400 ;
        RECT 427.950 334.950 430.050 337.050 ;
        RECT 381.750 329.100 392.850 329.700 ;
        RECT 350.700 315.600 352.500 326.400 ;
        RECT 359.550 315.600 361.350 327.600 ;
        RECT 364.950 327.300 367.050 328.200 ;
        RECT 367.950 327.300 373.050 328.200 ;
        RECT 375.150 328.500 392.850 329.100 ;
        RECT 375.150 328.200 383.550 328.500 ;
        RECT 367.950 326.400 368.850 327.300 ;
        RECT 366.150 324.600 368.850 326.400 ;
        RECT 369.750 326.100 371.550 326.400 ;
        RECT 375.150 326.100 376.050 328.200 ;
        RECT 391.950 327.600 392.850 328.500 ;
        RECT 410.400 327.600 411.300 334.950 ;
        RECT 428.400 327.600 429.600 334.950 ;
        RECT 431.100 334.050 432.900 335.850 ;
        RECT 433.950 334.950 436.050 337.050 ;
        RECT 430.950 331.950 433.050 334.050 ;
        RECT 434.100 333.150 435.900 334.950 ;
        RECT 437.100 334.050 438.900 335.850 ;
        RECT 436.950 331.950 439.050 334.050 ;
        RECT 441.150 329.700 442.050 344.400 ;
        RECT 449.550 343.800 451.350 345.600 ;
        RECT 452.850 345.450 457.800 346.500 ;
        RECT 465.300 346.500 466.350 347.400 ;
        RECT 452.850 344.700 454.650 345.450 ;
        RECT 465.300 345.300 469.050 346.500 ;
        RECT 466.950 344.400 469.050 345.300 ;
        RECT 472.650 344.400 474.450 350.400 ;
        RECT 490.500 345.600 492.300 350.400 ;
        RECT 514.800 347.400 516.600 350.400 ;
        RECT 490.500 344.400 495.600 345.600 ;
        RECT 449.850 342.000 450.900 343.800 ;
        RECT 460.050 342.000 461.850 342.600 ;
        RECT 449.850 340.800 461.850 342.000 ;
        RECT 444.000 339.600 450.900 340.800 ;
        RECT 444.000 338.850 444.900 339.600 ;
        RECT 449.100 339.000 450.900 339.600 ;
        RECT 443.100 337.050 444.900 338.850 ;
        RECT 446.100 337.800 447.900 338.400 ;
        RECT 442.950 334.950 445.050 337.050 ;
        RECT 446.100 336.600 454.050 337.800 ;
        RECT 451.950 334.950 454.050 336.600 ;
        RECT 450.450 329.700 452.250 330.000 ;
        RECT 441.150 329.100 452.250 329.700 ;
        RECT 441.150 328.500 458.850 329.100 ;
        RECT 441.150 327.600 442.050 328.500 ;
        RECT 450.450 328.200 458.850 328.500 ;
        RECT 369.750 325.200 376.050 326.100 ;
        RECT 376.950 326.700 378.750 327.300 ;
        RECT 376.950 325.500 384.450 326.700 ;
        RECT 369.750 324.600 371.550 325.200 ;
        RECT 383.250 324.600 384.450 325.500 ;
        RECT 364.950 321.600 368.850 323.700 ;
        RECT 373.950 323.550 375.750 324.300 ;
        RECT 378.750 323.550 380.550 324.300 ;
        RECT 373.950 322.500 380.550 323.550 ;
        RECT 383.250 322.500 388.050 324.600 ;
        RECT 367.050 315.600 368.850 321.600 ;
        RECT 374.850 315.600 376.650 322.500 ;
        RECT 383.250 321.600 384.450 322.500 ;
        RECT 382.650 315.600 384.450 321.600 ;
        RECT 391.050 315.600 392.850 327.600 ;
        RECT 407.700 326.400 411.300 327.600 ;
        RECT 407.700 315.600 409.500 326.400 ;
        RECT 427.800 315.600 429.600 327.600 ;
        RECT 430.800 326.700 438.600 327.600 ;
        RECT 430.800 315.600 432.600 326.700 ;
        RECT 436.800 315.600 438.600 326.700 ;
        RECT 441.150 315.600 442.950 327.600 ;
        RECT 455.250 326.700 457.050 327.300 ;
        RECT 449.550 325.500 457.050 326.700 ;
        RECT 457.950 326.100 458.850 328.200 ;
        RECT 460.950 328.200 461.850 340.800 ;
        RECT 473.250 337.050 474.450 344.400 ;
        RECT 494.400 337.050 495.600 344.400 ;
        RECT 505.950 337.950 508.050 340.050 ;
        RECT 511.950 337.950 514.050 340.050 ;
        RECT 468.150 335.250 474.450 337.050 ;
        RECT 469.950 334.950 474.450 335.250 ;
        RECT 470.250 329.400 472.050 331.200 ;
        RECT 466.950 328.200 471.150 329.400 ;
        RECT 460.950 327.300 466.050 328.200 ;
        RECT 466.950 327.300 469.050 328.200 ;
        RECT 473.250 327.600 474.450 334.950 ;
        RECT 485.100 334.050 486.900 335.850 ;
        RECT 487.950 334.950 490.050 337.050 ;
        RECT 484.950 331.950 487.050 334.050 ;
        RECT 488.100 333.150 489.900 334.950 ;
        RECT 491.100 334.050 492.900 335.850 ;
        RECT 493.950 334.950 496.050 337.050 ;
        RECT 490.950 331.950 493.050 334.050 ;
        RECT 494.400 327.600 495.600 334.950 ;
        RECT 506.550 328.050 507.450 337.950 ;
        RECT 512.100 336.150 513.900 337.950 ;
        RECT 515.400 337.050 516.300 347.400 ;
        RECT 521.550 344.400 523.350 350.400 ;
        RECT 529.650 347.400 531.450 350.400 ;
        RECT 537.450 347.400 539.250 350.400 ;
        RECT 545.250 348.300 547.050 350.400 ;
        RECT 545.250 347.400 549.000 348.300 ;
        RECT 529.650 346.500 530.700 347.400 ;
        RECT 526.950 345.300 530.700 346.500 ;
        RECT 538.200 346.500 539.250 347.400 ;
        RECT 547.950 346.500 549.000 347.400 ;
        RECT 538.200 345.450 543.150 346.500 ;
        RECT 526.950 344.400 529.050 345.300 ;
        RECT 541.350 344.700 543.150 345.450 ;
        RECT 517.950 337.950 520.050 340.050 ;
        RECT 514.950 334.950 517.050 337.050 ;
        RECT 518.100 336.150 519.900 337.950 ;
        RECT 521.550 337.050 522.750 344.400 ;
        RECT 544.650 343.800 546.450 345.600 ;
        RECT 547.950 344.400 550.050 346.500 ;
        RECT 553.050 344.400 554.850 350.400 ;
        RECT 534.150 342.000 535.950 342.600 ;
        RECT 545.100 342.000 546.150 343.800 ;
        RECT 534.150 340.800 546.150 342.000 ;
        RECT 521.550 335.250 527.850 337.050 ;
        RECT 521.550 334.950 526.050 335.250 ;
        RECT 465.150 326.400 466.050 327.300 ;
        RECT 462.450 326.100 464.250 326.400 ;
        RECT 449.550 324.600 450.750 325.500 ;
        RECT 457.950 325.200 464.250 326.100 ;
        RECT 462.450 324.600 464.250 325.200 ;
        RECT 465.150 324.600 467.850 326.400 ;
        RECT 445.950 322.500 450.750 324.600 ;
        RECT 453.450 323.550 455.250 324.300 ;
        RECT 458.250 323.550 460.050 324.300 ;
        RECT 453.450 322.500 460.050 323.550 ;
        RECT 449.550 321.600 450.750 322.500 ;
        RECT 449.550 315.600 451.350 321.600 ;
        RECT 457.350 315.600 459.150 322.500 ;
        RECT 465.150 321.600 469.050 323.700 ;
        RECT 465.150 315.600 466.950 321.600 ;
        RECT 472.650 315.600 474.450 327.600 ;
        RECT 485.400 326.700 493.200 327.600 ;
        RECT 485.400 315.600 487.200 326.700 ;
        RECT 491.400 315.600 493.200 326.700 ;
        RECT 494.400 315.600 496.200 327.600 ;
        RECT 505.950 325.950 508.050 328.050 ;
        RECT 515.400 327.600 516.300 334.950 ;
        RECT 512.700 326.400 516.300 327.600 ;
        RECT 521.550 327.600 522.750 334.950 ;
        RECT 523.950 329.400 525.750 331.200 ;
        RECT 524.850 328.200 529.050 329.400 ;
        RECT 534.150 328.200 535.050 340.800 ;
        RECT 545.100 339.600 552.000 340.800 ;
        RECT 545.100 339.000 546.900 339.600 ;
        RECT 551.100 338.850 552.000 339.600 ;
        RECT 548.100 337.800 549.900 338.400 ;
        RECT 541.950 336.600 549.900 337.800 ;
        RECT 551.100 337.050 552.900 338.850 ;
        RECT 541.950 334.950 544.050 336.600 ;
        RECT 550.950 334.950 553.050 337.050 ;
        RECT 543.750 329.700 545.550 330.000 ;
        RECT 553.950 329.700 554.850 344.400 ;
        RECT 543.750 329.100 554.850 329.700 ;
        RECT 512.700 315.600 514.500 326.400 ;
        RECT 521.550 315.600 523.350 327.600 ;
        RECT 526.950 327.300 529.050 328.200 ;
        RECT 529.950 327.300 535.050 328.200 ;
        RECT 537.150 328.500 554.850 329.100 ;
        RECT 537.150 328.200 545.550 328.500 ;
        RECT 529.950 326.400 530.850 327.300 ;
        RECT 528.150 324.600 530.850 326.400 ;
        RECT 531.750 326.100 533.550 326.400 ;
        RECT 537.150 326.100 538.050 328.200 ;
        RECT 553.950 327.600 554.850 328.500 ;
        RECT 531.750 325.200 538.050 326.100 ;
        RECT 538.950 326.700 540.750 327.300 ;
        RECT 538.950 325.500 546.450 326.700 ;
        RECT 531.750 324.600 533.550 325.200 ;
        RECT 545.250 324.600 546.450 325.500 ;
        RECT 526.950 321.600 530.850 323.700 ;
        RECT 535.950 323.550 537.750 324.300 ;
        RECT 540.750 323.550 542.550 324.300 ;
        RECT 535.950 322.500 542.550 323.550 ;
        RECT 545.250 322.500 550.050 324.600 ;
        RECT 529.050 315.600 530.850 321.600 ;
        RECT 536.850 315.600 538.650 322.500 ;
        RECT 545.250 321.600 546.450 322.500 ;
        RECT 544.650 315.600 546.450 321.600 ;
        RECT 553.050 315.600 554.850 327.600 ;
        RECT 558.150 344.400 559.950 350.400 ;
        RECT 565.950 348.300 567.750 350.400 ;
        RECT 564.000 347.400 567.750 348.300 ;
        RECT 573.750 347.400 575.550 350.400 ;
        RECT 581.550 347.400 583.350 350.400 ;
        RECT 564.000 346.500 565.050 347.400 ;
        RECT 573.750 346.500 574.800 347.400 ;
        RECT 562.950 344.400 565.050 346.500 ;
        RECT 558.150 329.700 559.050 344.400 ;
        RECT 566.550 343.800 568.350 345.600 ;
        RECT 569.850 345.450 574.800 346.500 ;
        RECT 582.300 346.500 583.350 347.400 ;
        RECT 569.850 344.700 571.650 345.450 ;
        RECT 582.300 345.300 586.050 346.500 ;
        RECT 583.950 344.400 586.050 345.300 ;
        RECT 589.650 344.400 591.450 350.400 ;
        RECT 605.400 347.400 607.200 350.400 ;
        RECT 566.850 342.000 567.900 343.800 ;
        RECT 577.050 342.000 578.850 342.600 ;
        RECT 566.850 340.800 578.850 342.000 ;
        RECT 561.000 339.600 567.900 340.800 ;
        RECT 561.000 338.850 561.900 339.600 ;
        RECT 566.100 339.000 567.900 339.600 ;
        RECT 560.100 337.050 561.900 338.850 ;
        RECT 563.100 337.800 564.900 338.400 ;
        RECT 559.950 334.950 562.050 337.050 ;
        RECT 563.100 336.600 571.050 337.800 ;
        RECT 568.950 334.950 571.050 336.600 ;
        RECT 567.450 329.700 569.250 330.000 ;
        RECT 558.150 329.100 569.250 329.700 ;
        RECT 558.150 328.500 575.850 329.100 ;
        RECT 558.150 327.600 559.050 328.500 ;
        RECT 567.450 328.200 575.850 328.500 ;
        RECT 558.150 315.600 559.950 327.600 ;
        RECT 572.250 326.700 574.050 327.300 ;
        RECT 566.550 325.500 574.050 326.700 ;
        RECT 574.950 326.100 575.850 328.200 ;
        RECT 577.950 328.200 578.850 340.800 ;
        RECT 590.250 337.050 591.450 344.400 ;
        RECT 601.950 337.950 604.050 340.050 ;
        RECT 585.150 335.250 591.450 337.050 ;
        RECT 602.100 336.150 603.900 337.950 ;
        RECT 605.700 337.050 606.600 347.400 ;
        RECT 613.950 346.950 616.050 349.050 ;
        RECT 626.400 347.400 628.200 350.400 ;
        RECT 644.400 347.400 646.200 350.400 ;
        RECT 614.550 340.050 615.450 346.950 ;
        RECT 607.950 337.950 610.050 340.050 ;
        RECT 613.950 337.950 616.050 340.050 ;
        RECT 586.950 334.950 591.450 335.250 ;
        RECT 604.950 334.950 607.050 337.050 ;
        RECT 608.100 336.150 609.900 337.950 ;
        RECT 622.950 334.950 625.050 337.050 ;
        RECT 587.250 329.400 589.050 331.200 ;
        RECT 583.950 328.200 588.150 329.400 ;
        RECT 577.950 327.300 583.050 328.200 ;
        RECT 583.950 327.300 586.050 328.200 ;
        RECT 590.250 327.600 591.450 334.950 ;
        RECT 582.150 326.400 583.050 327.300 ;
        RECT 579.450 326.100 581.250 326.400 ;
        RECT 566.550 324.600 567.750 325.500 ;
        RECT 574.950 325.200 581.250 326.100 ;
        RECT 579.450 324.600 581.250 325.200 ;
        RECT 582.150 324.600 584.850 326.400 ;
        RECT 562.950 322.500 567.750 324.600 ;
        RECT 570.450 323.550 572.250 324.300 ;
        RECT 575.250 323.550 577.050 324.300 ;
        RECT 570.450 322.500 577.050 323.550 ;
        RECT 566.550 321.600 567.750 322.500 ;
        RECT 566.550 315.600 568.350 321.600 ;
        RECT 574.350 315.600 576.150 322.500 ;
        RECT 582.150 321.600 586.050 323.700 ;
        RECT 582.150 315.600 583.950 321.600 ;
        RECT 589.650 315.600 591.450 327.600 ;
        RECT 605.700 327.600 606.600 334.950 ;
        RECT 623.100 333.150 624.900 334.950 ;
        RECT 626.400 334.050 627.600 347.400 ;
        RECT 640.950 337.950 643.050 340.050 ;
        RECT 641.100 336.150 642.900 337.950 ;
        RECT 644.700 337.050 645.600 347.400 ;
        RECT 667.500 345.600 669.300 350.400 ;
        RECT 667.500 344.400 672.600 345.600 ;
        RECT 691.200 344.400 693.000 350.400 ;
        RECT 716.400 347.400 718.200 350.400 ;
        RECT 646.950 337.950 649.050 340.050 ;
        RECT 643.950 334.950 646.050 337.050 ;
        RECT 647.100 336.150 648.900 337.950 ;
        RECT 671.400 337.050 672.600 344.400 ;
        RECT 686.100 337.050 687.900 338.850 ;
        RECT 688.950 337.950 691.050 340.050 ;
        RECT 625.950 328.950 628.050 334.050 ;
        RECT 605.700 326.400 609.300 327.600 ;
        RECT 607.500 315.600 609.300 326.400 ;
        RECT 626.400 321.600 627.600 328.950 ;
        RECT 644.700 327.600 645.600 334.950 ;
        RECT 662.100 334.050 663.900 335.850 ;
        RECT 664.950 334.950 667.050 337.050 ;
        RECT 661.950 331.950 664.050 334.050 ;
        RECT 665.100 333.150 666.900 334.950 ;
        RECT 668.100 334.050 669.900 335.850 ;
        RECT 670.950 334.950 673.050 337.050 ;
        RECT 685.950 334.950 688.050 337.050 ;
        RECT 689.100 336.150 690.900 337.950 ;
        RECT 691.950 337.050 693.000 344.400 ;
        RECT 717.300 343.200 718.200 347.400 ;
        RECT 722.400 344.400 724.200 350.400 ;
        RECT 729.150 344.400 730.950 350.400 ;
        RECT 736.950 348.300 738.750 350.400 ;
        RECT 735.000 347.400 738.750 348.300 ;
        RECT 744.750 347.400 746.550 350.400 ;
        RECT 752.550 347.400 754.350 350.400 ;
        RECT 735.000 346.500 736.050 347.400 ;
        RECT 744.750 346.500 745.800 347.400 ;
        RECT 733.950 344.400 736.050 346.500 ;
        RECT 717.300 342.300 720.600 343.200 ;
        RECT 718.800 341.400 720.600 342.300 ;
        RECT 694.950 337.950 697.050 340.050 ;
        RECT 691.950 334.950 694.050 337.050 ;
        RECT 695.100 336.150 696.900 337.950 ;
        RECT 698.100 337.050 699.900 338.850 ;
        RECT 697.950 334.950 700.050 337.050 ;
        RECT 667.950 331.950 670.050 334.050 ;
        RECT 671.400 327.600 672.600 334.950 ;
        RECT 692.100 329.400 693.000 334.950 ;
        RECT 713.100 334.050 714.900 335.850 ;
        RECT 715.950 334.950 718.050 337.050 ;
        RECT 712.950 331.950 715.050 334.050 ;
        RECT 716.100 333.150 717.900 334.950 ;
        RECT 719.700 330.900 720.600 341.400 ;
        RECT 723.000 337.050 724.050 344.400 ;
        RECT 718.800 330.300 720.600 330.900 ;
        RECT 692.100 328.500 697.200 329.400 ;
        RECT 644.700 326.400 648.300 327.600 ;
        RECT 626.400 315.600 628.200 321.600 ;
        RECT 646.500 315.600 648.300 326.400 ;
        RECT 662.400 326.700 670.200 327.600 ;
        RECT 662.400 315.600 664.200 326.700 ;
        RECT 668.400 315.600 670.200 326.700 ;
        RECT 671.400 315.600 673.200 327.600 ;
        RECT 686.400 326.400 694.200 327.300 ;
        RECT 686.400 315.600 688.200 326.400 ;
        RECT 692.400 316.500 694.200 326.400 ;
        RECT 695.400 317.400 697.200 328.500 ;
        RECT 713.400 329.100 720.600 330.300 ;
        RECT 721.950 334.950 724.050 337.050 ;
        RECT 713.400 327.600 714.600 329.100 ;
        RECT 721.950 327.600 723.300 334.950 ;
        RECT 698.400 316.500 700.200 327.600 ;
        RECT 692.400 315.600 700.200 316.500 ;
        RECT 713.400 315.600 715.200 327.600 ;
        RECT 720.900 326.100 723.300 327.600 ;
        RECT 729.150 329.700 730.050 344.400 ;
        RECT 737.550 343.800 739.350 345.600 ;
        RECT 740.850 345.450 745.800 346.500 ;
        RECT 753.300 346.500 754.350 347.400 ;
        RECT 740.850 344.700 742.650 345.450 ;
        RECT 753.300 345.300 757.050 346.500 ;
        RECT 754.950 344.400 757.050 345.300 ;
        RECT 760.650 344.400 762.450 350.400 ;
        RECT 737.850 342.000 738.900 343.800 ;
        RECT 748.050 342.000 749.850 342.600 ;
        RECT 737.850 340.800 749.850 342.000 ;
        RECT 732.000 339.600 738.900 340.800 ;
        RECT 732.000 338.850 732.900 339.600 ;
        RECT 737.100 339.000 738.900 339.600 ;
        RECT 731.100 337.050 732.900 338.850 ;
        RECT 734.100 337.800 735.900 338.400 ;
        RECT 730.950 334.950 733.050 337.050 ;
        RECT 734.100 336.600 742.050 337.800 ;
        RECT 739.950 334.950 742.050 336.600 ;
        RECT 738.450 329.700 740.250 330.000 ;
        RECT 729.150 329.100 740.250 329.700 ;
        RECT 729.150 328.500 746.850 329.100 ;
        RECT 729.150 327.600 730.050 328.500 ;
        RECT 738.450 328.200 746.850 328.500 ;
        RECT 720.900 315.600 722.700 326.100 ;
        RECT 729.150 315.600 730.950 327.600 ;
        RECT 743.250 326.700 745.050 327.300 ;
        RECT 737.550 325.500 745.050 326.700 ;
        RECT 745.950 326.100 746.850 328.200 ;
        RECT 748.950 328.200 749.850 340.800 ;
        RECT 761.250 337.050 762.450 344.400 ;
        RECT 776.400 347.400 778.200 350.400 ;
        RECT 796.800 347.400 798.600 350.400 ;
        RECT 815.400 347.400 817.200 350.400 ;
        RECT 756.150 335.250 762.450 337.050 ;
        RECT 757.950 334.950 762.450 335.250 ;
        RECT 772.950 334.950 775.050 337.050 ;
        RECT 758.250 329.400 760.050 331.200 ;
        RECT 754.950 328.200 759.150 329.400 ;
        RECT 748.950 327.300 754.050 328.200 ;
        RECT 754.950 327.300 757.050 328.200 ;
        RECT 761.250 327.600 762.450 334.950 ;
        RECT 773.100 333.150 774.900 334.950 ;
        RECT 776.400 334.050 777.600 347.400 ;
        RECT 778.950 343.950 781.050 346.050 ;
        RECT 779.550 337.050 780.450 343.950 ;
        RECT 793.950 337.950 796.050 340.050 ;
        RECT 778.950 334.950 781.050 337.050 ;
        RECT 794.100 336.150 795.900 337.950 ;
        RECT 797.400 337.050 798.300 347.400 ;
        RECT 799.950 337.950 802.050 340.050 ;
        RECT 796.950 334.950 799.050 337.050 ;
        RECT 800.100 336.150 801.900 337.950 ;
        RECT 811.950 334.950 814.050 337.050 ;
        RECT 775.950 328.950 778.050 334.050 ;
        RECT 753.150 326.400 754.050 327.300 ;
        RECT 750.450 326.100 752.250 326.400 ;
        RECT 737.550 324.600 738.750 325.500 ;
        RECT 745.950 325.200 752.250 326.100 ;
        RECT 750.450 324.600 752.250 325.200 ;
        RECT 753.150 324.600 755.850 326.400 ;
        RECT 733.950 322.500 738.750 324.600 ;
        RECT 741.450 323.550 743.250 324.300 ;
        RECT 746.250 323.550 748.050 324.300 ;
        RECT 741.450 322.500 748.050 323.550 ;
        RECT 737.550 321.600 738.750 322.500 ;
        RECT 737.550 315.600 739.350 321.600 ;
        RECT 745.350 315.600 747.150 322.500 ;
        RECT 753.150 321.600 757.050 323.700 ;
        RECT 753.150 315.600 754.950 321.600 ;
        RECT 760.650 315.600 762.450 327.600 ;
        RECT 776.400 321.600 777.600 328.950 ;
        RECT 797.400 327.600 798.300 334.950 ;
        RECT 812.100 333.150 813.900 334.950 ;
        RECT 815.400 334.050 816.600 347.400 ;
        RECT 833.400 343.200 835.200 350.400 ;
        RECT 854.400 347.400 856.200 350.400 ;
        RECT 871.800 349.500 879.600 350.400 ;
        RECT 833.400 342.300 837.600 343.200 ;
        RECT 836.400 337.050 837.600 342.300 ;
        RECT 833.100 334.050 834.900 335.850 ;
        RECT 835.950 334.950 838.050 337.050 ;
        RECT 814.950 328.950 817.050 334.050 ;
        RECT 832.950 331.950 835.050 334.050 ;
        RECT 794.700 326.400 798.300 327.600 ;
        RECT 776.400 315.600 778.200 321.600 ;
        RECT 794.700 315.600 796.500 326.400 ;
        RECT 815.400 321.600 816.600 328.950 ;
        RECT 836.400 321.600 837.600 334.950 ;
        RECT 839.100 334.050 840.900 335.850 ;
        RECT 850.950 334.950 853.050 337.050 ;
        RECT 838.950 331.950 841.050 334.050 ;
        RECT 851.100 333.150 852.900 334.950 ;
        RECT 854.400 334.050 855.600 347.400 ;
        RECT 871.800 344.400 873.600 349.500 ;
        RECT 874.800 344.400 876.600 348.600 ;
        RECT 877.800 345.000 879.600 349.500 ;
        RECT 883.800 345.000 885.600 350.400 ;
        RECT 898.800 347.400 900.600 350.400 ;
        RECT 875.400 342.900 876.300 344.400 ;
        RECT 877.800 344.100 885.600 345.000 ;
        RECT 875.400 341.700 880.050 342.900 ;
        RECT 878.700 337.050 880.050 341.700 ;
        RECT 889.950 337.950 892.050 340.050 ;
        RECT 871.950 334.950 874.050 337.050 ;
        RECT 853.950 328.950 856.050 334.050 ;
        RECT 872.100 333.150 873.900 334.950 ;
        RECT 875.100 334.050 876.900 335.850 ;
        RECT 877.950 334.950 880.050 337.050 ;
        RECT 874.950 331.950 877.050 334.050 ;
        RECT 815.400 315.600 817.200 321.600 ;
        RECT 835.800 315.600 837.600 321.600 ;
        RECT 854.400 321.600 855.600 328.950 ;
        RECT 878.700 327.600 879.900 334.950 ;
        RECT 881.100 334.050 882.900 335.850 ;
        RECT 883.950 334.950 886.050 337.050 ;
        RECT 880.950 331.950 883.050 334.050 ;
        RECT 884.100 333.150 885.900 334.950 ;
        RECT 854.400 315.600 856.200 321.600 ;
        RECT 877.800 315.600 881.100 327.600 ;
        RECT 890.550 319.050 891.450 337.950 ;
        RECT 899.400 334.050 900.600 347.400 ;
        RECT 901.950 334.950 904.050 337.050 ;
        RECT 898.950 328.950 901.050 334.050 ;
        RECT 902.100 333.150 903.900 334.950 ;
        RECT 899.400 321.600 900.600 328.950 ;
        RECT 889.950 316.950 892.050 319.050 ;
        RECT 898.800 315.600 900.600 321.600 ;
        RECT 14.700 300.600 16.500 311.400 ;
        RECT 34.800 305.400 36.600 311.400 ;
        RECT 35.700 305.100 36.600 305.400 ;
        RECT 40.800 305.400 42.600 311.400 ;
        RECT 62.400 305.400 64.200 311.400 ;
        RECT 82.800 305.400 84.600 311.400 ;
        RECT 103.800 305.400 105.600 311.400 ;
        RECT 125.400 305.400 127.200 311.400 ;
        RECT 146.400 305.400 148.200 311.400 ;
        RECT 40.800 305.100 42.300 305.400 ;
        RECT 35.700 304.200 42.300 305.100 ;
        RECT 14.700 299.400 18.300 300.600 ;
        RECT 17.400 292.050 18.300 299.400 ;
        RECT 35.700 292.050 36.600 304.200 ;
        RECT 37.950 292.950 40.050 295.050 ;
        RECT 14.100 289.050 15.900 290.850 ;
        RECT 16.950 289.950 19.050 292.050 ;
        RECT 13.950 286.950 16.050 289.050 ;
        RECT 17.400 279.600 18.300 289.950 ;
        RECT 20.100 289.050 21.900 290.850 ;
        RECT 34.950 289.950 37.050 292.050 ;
        RECT 38.100 291.150 39.900 292.950 ;
        RECT 41.100 292.050 42.900 293.850 ;
        RECT 43.950 292.950 46.050 295.050 ;
        RECT 58.950 292.950 61.050 295.050 ;
        RECT 40.950 289.950 43.050 292.050 ;
        RECT 44.100 291.150 45.900 292.950 ;
        RECT 59.100 291.150 60.900 292.950 ;
        RECT 62.850 292.050 64.050 305.400 ;
        RECT 83.400 298.050 84.600 305.400 ;
        RECT 64.950 292.950 67.050 295.050 ;
        RECT 61.950 289.950 64.050 292.050 ;
        RECT 65.100 291.150 66.900 292.950 ;
        RECT 68.100 292.050 69.900 293.850 ;
        RECT 82.950 292.950 85.050 298.050 ;
        RECT 67.950 289.950 70.050 292.050 ;
        RECT 19.950 286.950 22.050 289.050 ;
        RECT 35.700 286.200 36.600 289.950 ;
        RECT 35.700 285.000 39.000 286.200 ;
        RECT 61.950 285.750 63.150 289.950 ;
        RECT 16.800 276.600 18.600 279.600 ;
        RECT 37.200 276.600 39.000 285.000 ;
        RECT 59.400 284.700 63.150 285.750 ;
        RECT 59.400 282.600 60.600 284.700 ;
        RECT 58.800 276.600 60.600 282.600 ;
        RECT 61.800 281.700 69.600 283.050 ;
        RECT 61.800 276.600 63.600 281.700 ;
        RECT 67.800 276.600 69.600 281.700 ;
        RECT 83.400 279.600 84.600 292.950 ;
        RECT 86.100 292.050 87.900 293.850 ;
        RECT 98.100 292.050 99.900 293.850 ;
        RECT 100.950 292.950 103.050 295.050 ;
        RECT 85.950 289.950 88.050 292.050 ;
        RECT 97.950 289.950 100.050 292.050 ;
        RECT 101.100 291.150 102.900 292.950 ;
        RECT 103.950 292.050 105.150 305.400 ;
        RECT 106.950 292.950 109.050 295.050 ;
        RECT 121.950 292.950 124.050 295.050 ;
        RECT 103.950 289.950 106.050 292.050 ;
        RECT 107.100 291.150 108.900 292.950 ;
        RECT 122.100 291.150 123.900 292.950 ;
        RECT 125.400 292.050 126.600 305.400 ;
        RECT 146.400 298.050 147.600 305.400 ;
        RECT 152.550 299.400 154.350 311.400 ;
        RECT 160.050 305.400 161.850 311.400 ;
        RECT 157.950 303.300 161.850 305.400 ;
        RECT 167.850 304.500 169.650 311.400 ;
        RECT 175.650 305.400 177.450 311.400 ;
        RECT 176.250 304.500 177.450 305.400 ;
        RECT 166.950 303.450 173.550 304.500 ;
        RECT 166.950 302.700 168.750 303.450 ;
        RECT 171.750 302.700 173.550 303.450 ;
        RECT 176.250 302.400 181.050 304.500 ;
        RECT 159.150 300.600 161.850 302.400 ;
        RECT 162.750 301.800 164.550 302.400 ;
        RECT 162.750 300.900 169.050 301.800 ;
        RECT 176.250 301.500 177.450 302.400 ;
        RECT 162.750 300.600 164.550 300.900 ;
        RECT 160.950 299.700 161.850 300.600 ;
        RECT 127.950 292.950 130.050 295.050 ;
        RECT 124.950 289.950 127.050 292.050 ;
        RECT 128.100 291.150 129.900 292.950 ;
        RECT 143.100 292.050 144.900 293.850 ;
        RECT 145.950 292.950 148.050 298.050 ;
        RECT 142.950 289.950 145.050 292.050 ;
        RECT 104.850 285.750 106.050 289.950 ;
        RECT 104.850 284.700 108.600 285.750 ;
        RECT 82.800 276.600 84.600 279.600 ;
        RECT 98.400 281.700 106.200 283.050 ;
        RECT 98.400 276.600 100.200 281.700 ;
        RECT 104.400 276.600 106.200 281.700 ;
        RECT 107.400 282.600 108.600 284.700 ;
        RECT 125.400 284.700 126.600 289.950 ;
        RECT 125.400 283.800 129.600 284.700 ;
        RECT 107.400 276.600 109.200 282.600 ;
        RECT 127.800 276.600 129.600 283.800 ;
        RECT 146.400 279.600 147.600 292.950 ;
        RECT 152.550 292.050 153.750 299.400 ;
        RECT 157.950 298.800 160.050 299.700 ;
        RECT 160.950 298.800 166.050 299.700 ;
        RECT 155.850 297.600 160.050 298.800 ;
        RECT 154.950 295.800 156.750 297.600 ;
        RECT 152.550 291.750 157.050 292.050 ;
        RECT 152.550 289.950 158.850 291.750 ;
        RECT 152.550 282.600 153.750 289.950 ;
        RECT 165.150 286.200 166.050 298.800 ;
        RECT 168.150 298.800 169.050 300.900 ;
        RECT 169.950 300.300 177.450 301.500 ;
        RECT 169.950 299.700 171.750 300.300 ;
        RECT 184.050 299.400 185.850 311.400 ;
        RECT 202.800 305.400 204.600 311.400 ;
        RECT 168.150 298.500 176.550 298.800 ;
        RECT 184.950 298.500 185.850 299.400 ;
        RECT 168.150 297.900 185.850 298.500 ;
        RECT 174.750 297.300 185.850 297.900 ;
        RECT 174.750 297.000 176.550 297.300 ;
        RECT 172.950 290.400 175.050 292.050 ;
        RECT 172.950 289.200 180.900 290.400 ;
        RECT 181.950 289.950 184.050 292.050 ;
        RECT 179.100 288.600 180.900 289.200 ;
        RECT 182.100 288.150 183.900 289.950 ;
        RECT 176.100 287.400 177.900 288.000 ;
        RECT 182.100 287.400 183.000 288.150 ;
        RECT 176.100 286.200 183.000 287.400 ;
        RECT 165.150 285.000 177.150 286.200 ;
        RECT 165.150 284.400 166.950 285.000 ;
        RECT 176.100 283.200 177.150 285.000 ;
        RECT 146.400 276.600 148.200 279.600 ;
        RECT 152.550 276.600 154.350 282.600 ;
        RECT 157.950 281.700 160.050 282.600 ;
        RECT 157.950 280.500 161.700 281.700 ;
        RECT 172.350 281.550 174.150 282.300 ;
        RECT 160.650 279.600 161.700 280.500 ;
        RECT 169.200 280.500 174.150 281.550 ;
        RECT 175.650 281.400 177.450 283.200 ;
        RECT 184.950 282.600 185.850 297.300 ;
        RECT 197.100 292.050 198.900 293.850 ;
        RECT 199.950 292.950 202.050 295.050 ;
        RECT 196.950 289.950 199.050 292.050 ;
        RECT 200.100 291.150 201.900 292.950 ;
        RECT 202.950 292.050 204.150 305.400 ;
        RECT 211.950 304.950 214.050 307.050 ;
        RECT 224.400 305.400 226.200 311.400 ;
        RECT 205.950 292.950 208.050 295.050 ;
        RECT 202.950 289.950 205.050 292.050 ;
        RECT 206.100 291.150 207.900 292.950 ;
        RECT 203.850 285.750 205.050 289.950 ;
        RECT 203.850 284.700 207.600 285.750 ;
        RECT 178.950 280.500 181.050 282.600 ;
        RECT 169.200 279.600 170.250 280.500 ;
        RECT 178.950 279.600 180.000 280.500 ;
        RECT 160.650 276.600 162.450 279.600 ;
        RECT 168.450 276.600 170.250 279.600 ;
        RECT 176.250 278.700 180.000 279.600 ;
        RECT 176.250 276.600 178.050 278.700 ;
        RECT 184.050 276.600 185.850 282.600 ;
        RECT 197.400 281.700 205.200 283.050 ;
        RECT 197.400 276.600 199.200 281.700 ;
        RECT 203.400 276.600 205.200 281.700 ;
        RECT 206.400 282.600 207.600 284.700 ;
        RECT 206.400 276.600 208.200 282.600 ;
        RECT 212.550 280.050 213.450 304.950 ;
        RECT 220.950 292.950 223.050 295.050 ;
        RECT 221.100 291.150 222.900 292.950 ;
        RECT 224.400 292.050 225.600 305.400 ;
        RECT 245.700 300.600 247.500 311.400 ;
        RECT 245.700 299.400 249.300 300.600 ;
        RECT 226.950 292.950 229.050 295.050 ;
        RECT 223.950 289.950 226.050 292.050 ;
        RECT 227.100 291.150 228.900 292.950 ;
        RECT 248.400 292.050 249.300 299.400 ;
        RECT 254.550 299.400 256.350 311.400 ;
        RECT 262.050 305.400 263.850 311.400 ;
        RECT 259.950 303.300 263.850 305.400 ;
        RECT 269.850 304.500 271.650 311.400 ;
        RECT 277.650 305.400 279.450 311.400 ;
        RECT 278.250 304.500 279.450 305.400 ;
        RECT 268.950 303.450 275.550 304.500 ;
        RECT 268.950 302.700 270.750 303.450 ;
        RECT 273.750 302.700 275.550 303.450 ;
        RECT 278.250 302.400 283.050 304.500 ;
        RECT 261.150 300.600 263.850 302.400 ;
        RECT 264.750 301.800 266.550 302.400 ;
        RECT 264.750 300.900 271.050 301.800 ;
        RECT 278.250 301.500 279.450 302.400 ;
        RECT 264.750 300.600 266.550 300.900 ;
        RECT 262.950 299.700 263.850 300.600 ;
        RECT 254.550 292.050 255.750 299.400 ;
        RECT 259.950 298.800 262.050 299.700 ;
        RECT 262.950 298.800 268.050 299.700 ;
        RECT 257.850 297.600 262.050 298.800 ;
        RECT 256.950 295.800 258.750 297.600 ;
        RECT 224.400 284.700 225.600 289.950 ;
        RECT 245.100 289.050 246.900 290.850 ;
        RECT 247.950 289.950 250.050 292.050 ;
        RECT 254.550 291.750 259.050 292.050 ;
        RECT 244.950 286.950 247.050 289.050 ;
        RECT 224.400 283.800 228.600 284.700 ;
        RECT 211.950 277.950 214.050 280.050 ;
        RECT 226.800 276.600 228.600 283.800 ;
        RECT 248.400 279.600 249.300 289.950 ;
        RECT 251.100 289.050 252.900 290.850 ;
        RECT 254.550 289.950 260.850 291.750 ;
        RECT 250.950 286.950 253.050 289.050 ;
        RECT 254.550 282.600 255.750 289.950 ;
        RECT 267.150 286.200 268.050 298.800 ;
        RECT 270.150 298.800 271.050 300.900 ;
        RECT 271.950 300.300 279.450 301.500 ;
        RECT 271.950 299.700 273.750 300.300 ;
        RECT 286.050 299.400 287.850 311.400 ;
        RECT 301.800 299.400 303.600 311.400 ;
        RECT 304.800 300.300 306.600 311.400 ;
        RECT 310.800 300.300 312.600 311.400 ;
        RECT 304.800 299.400 312.600 300.300 ;
        RECT 270.150 298.500 278.550 298.800 ;
        RECT 286.950 298.500 287.850 299.400 ;
        RECT 270.150 297.900 287.850 298.500 ;
        RECT 276.750 297.300 287.850 297.900 ;
        RECT 276.750 297.000 278.550 297.300 ;
        RECT 274.950 290.400 277.050 292.050 ;
        RECT 274.950 289.200 282.900 290.400 ;
        RECT 283.950 289.950 286.050 292.050 ;
        RECT 281.100 288.600 282.900 289.200 ;
        RECT 284.100 288.150 285.900 289.950 ;
        RECT 278.100 287.400 279.900 288.000 ;
        RECT 284.100 287.400 285.000 288.150 ;
        RECT 278.100 286.200 285.000 287.400 ;
        RECT 267.150 285.000 279.150 286.200 ;
        RECT 267.150 284.400 268.950 285.000 ;
        RECT 278.100 283.200 279.150 285.000 ;
        RECT 247.800 276.600 249.600 279.600 ;
        RECT 254.550 276.600 256.350 282.600 ;
        RECT 259.950 281.700 262.050 282.600 ;
        RECT 259.950 280.500 263.700 281.700 ;
        RECT 274.350 281.550 276.150 282.300 ;
        RECT 262.650 279.600 263.700 280.500 ;
        RECT 271.200 280.500 276.150 281.550 ;
        RECT 277.650 281.400 279.450 283.200 ;
        RECT 286.950 282.600 287.850 297.300 ;
        RECT 302.400 292.050 303.600 299.400 ;
        RECT 328.800 298.500 330.600 311.400 ;
        RECT 334.800 298.500 336.600 311.400 ;
        RECT 340.800 298.500 342.600 311.400 ;
        RECT 346.800 298.500 348.600 311.400 ;
        RECT 362.400 300.300 364.200 311.400 ;
        RECT 368.400 300.300 370.200 311.400 ;
        RECT 362.400 299.400 370.200 300.300 ;
        RECT 371.400 299.400 373.200 311.400 ;
        RECT 378.150 299.400 379.950 311.400 ;
        RECT 386.550 305.400 388.350 311.400 ;
        RECT 386.550 304.500 387.750 305.400 ;
        RECT 394.350 304.500 396.150 311.400 ;
        RECT 402.150 305.400 403.950 311.400 ;
        RECT 382.950 302.400 387.750 304.500 ;
        RECT 390.450 303.450 397.050 304.500 ;
        RECT 390.450 302.700 392.250 303.450 ;
        RECT 395.250 302.700 397.050 303.450 ;
        RECT 402.150 303.300 406.050 305.400 ;
        RECT 386.550 301.500 387.750 302.400 ;
        RECT 399.450 301.800 401.250 302.400 ;
        RECT 386.550 300.300 394.050 301.500 ;
        RECT 392.250 299.700 394.050 300.300 ;
        RECT 394.950 300.900 401.250 301.800 ;
        RECT 327.900 297.300 330.600 298.500 ;
        RECT 332.700 297.300 336.600 298.500 ;
        RECT 338.700 297.300 342.600 298.500 ;
        RECT 344.700 297.300 348.600 298.500 ;
        RECT 304.950 292.950 307.050 295.050 ;
        RECT 301.950 289.950 304.050 292.050 ;
        RECT 305.100 291.150 306.900 292.950 ;
        RECT 308.100 292.050 309.900 293.850 ;
        RECT 310.950 292.950 313.050 295.050 ;
        RECT 307.950 289.950 310.050 292.050 ;
        RECT 311.100 291.150 312.900 292.950 ;
        RECT 327.900 292.050 328.800 297.300 ;
        RECT 325.950 289.950 328.800 292.050 ;
        RECT 280.950 280.500 283.050 282.600 ;
        RECT 271.200 279.600 272.250 280.500 ;
        RECT 280.950 279.600 282.000 280.500 ;
        RECT 262.650 276.600 264.450 279.600 ;
        RECT 270.450 276.600 272.250 279.600 ;
        RECT 278.250 278.700 282.000 279.600 ;
        RECT 278.250 276.600 280.050 278.700 ;
        RECT 286.050 276.600 287.850 282.600 ;
        RECT 302.400 282.600 303.600 289.950 ;
        RECT 327.900 284.700 328.800 289.950 ;
        RECT 329.700 286.800 331.500 287.400 ;
        RECT 332.700 286.800 333.900 297.300 ;
        RECT 329.700 285.600 333.900 286.800 ;
        RECT 335.700 286.800 337.500 287.400 ;
        RECT 338.700 286.800 339.900 297.300 ;
        RECT 335.700 285.600 339.900 286.800 ;
        RECT 341.700 286.800 343.500 287.400 ;
        RECT 344.700 286.800 345.900 297.300 ;
        RECT 361.950 292.950 364.050 295.050 ;
        RECT 346.950 289.950 349.050 292.050 ;
        RECT 362.100 291.150 363.900 292.950 ;
        RECT 365.100 292.050 366.900 293.850 ;
        RECT 367.950 292.950 370.050 295.050 ;
        RECT 364.950 289.950 367.050 292.050 ;
        RECT 368.100 291.150 369.900 292.950 ;
        RECT 371.400 292.050 372.600 299.400 ;
        RECT 378.150 298.500 379.050 299.400 ;
        RECT 394.950 298.800 395.850 300.900 ;
        RECT 399.450 300.600 401.250 300.900 ;
        RECT 402.150 300.600 404.850 302.400 ;
        RECT 402.150 299.700 403.050 300.600 ;
        RECT 387.450 298.500 395.850 298.800 ;
        RECT 378.150 297.900 395.850 298.500 ;
        RECT 397.950 298.800 403.050 299.700 ;
        RECT 403.950 298.800 406.050 299.700 ;
        RECT 409.650 299.400 411.450 311.400 ;
        RECT 378.150 297.300 389.250 297.900 ;
        RECT 370.950 289.950 373.050 292.050 ;
        RECT 347.100 288.150 348.900 289.950 ;
        RECT 341.700 285.600 345.900 286.800 ;
        RECT 332.700 284.700 333.900 285.600 ;
        RECT 338.700 284.700 339.900 285.600 ;
        RECT 344.700 284.700 345.900 285.600 ;
        RECT 327.900 283.500 330.600 284.700 ;
        RECT 332.700 283.500 336.600 284.700 ;
        RECT 338.700 283.500 342.600 284.700 ;
        RECT 344.700 283.500 348.600 284.700 ;
        RECT 302.400 281.400 307.500 282.600 ;
        RECT 305.700 276.600 307.500 281.400 ;
        RECT 328.800 276.600 330.600 283.500 ;
        RECT 334.800 276.600 336.600 283.500 ;
        RECT 340.800 276.600 342.600 283.500 ;
        RECT 346.800 276.600 348.600 283.500 ;
        RECT 371.400 282.600 372.600 289.950 ;
        RECT 367.500 281.400 372.600 282.600 ;
        RECT 378.150 282.600 379.050 297.300 ;
        RECT 387.450 297.000 389.250 297.300 ;
        RECT 379.950 289.950 382.050 292.050 ;
        RECT 388.950 290.400 391.050 292.050 ;
        RECT 380.100 288.150 381.900 289.950 ;
        RECT 383.100 289.200 391.050 290.400 ;
        RECT 383.100 288.600 384.900 289.200 ;
        RECT 381.000 287.400 381.900 288.150 ;
        RECT 386.100 287.400 387.900 288.000 ;
        RECT 381.000 286.200 387.900 287.400 ;
        RECT 397.950 286.200 398.850 298.800 ;
        RECT 403.950 297.600 408.150 298.800 ;
        RECT 407.250 295.800 409.050 297.600 ;
        RECT 410.250 292.050 411.450 299.400 ;
        RECT 406.950 291.750 411.450 292.050 ;
        RECT 405.150 289.950 411.450 291.750 ;
        RECT 386.850 285.000 398.850 286.200 ;
        RECT 386.850 283.200 387.900 285.000 ;
        RECT 397.050 284.400 398.850 285.000 ;
        RECT 367.500 276.600 369.300 281.400 ;
        RECT 378.150 276.600 379.950 282.600 ;
        RECT 382.950 280.500 385.050 282.600 ;
        RECT 386.550 281.400 388.350 283.200 ;
        RECT 410.250 282.600 411.450 289.950 ;
        RECT 389.850 281.550 391.650 282.300 ;
        RECT 403.950 281.700 406.050 282.600 ;
        RECT 389.850 280.500 394.800 281.550 ;
        RECT 384.000 279.600 385.050 280.500 ;
        RECT 393.750 279.600 394.800 280.500 ;
        RECT 402.300 280.500 406.050 281.700 ;
        RECT 402.300 279.600 403.350 280.500 ;
        RECT 384.000 278.700 387.750 279.600 ;
        RECT 385.950 276.600 387.750 278.700 ;
        RECT 393.750 276.600 395.550 279.600 ;
        RECT 401.550 276.600 403.350 279.600 ;
        RECT 409.650 276.600 411.450 282.600 ;
        RECT 413.550 299.400 415.350 311.400 ;
        RECT 421.050 305.400 422.850 311.400 ;
        RECT 418.950 303.300 422.850 305.400 ;
        RECT 428.850 304.500 430.650 311.400 ;
        RECT 436.650 305.400 438.450 311.400 ;
        RECT 437.250 304.500 438.450 305.400 ;
        RECT 427.950 303.450 434.550 304.500 ;
        RECT 427.950 302.700 429.750 303.450 ;
        RECT 432.750 302.700 434.550 303.450 ;
        RECT 437.250 302.400 442.050 304.500 ;
        RECT 420.150 300.600 422.850 302.400 ;
        RECT 423.750 301.800 425.550 302.400 ;
        RECT 423.750 300.900 430.050 301.800 ;
        RECT 437.250 301.500 438.450 302.400 ;
        RECT 423.750 300.600 425.550 300.900 ;
        RECT 421.950 299.700 422.850 300.600 ;
        RECT 413.550 292.050 414.750 299.400 ;
        RECT 418.950 298.800 421.050 299.700 ;
        RECT 421.950 298.800 427.050 299.700 ;
        RECT 416.850 297.600 421.050 298.800 ;
        RECT 415.950 295.800 417.750 297.600 ;
        RECT 413.550 291.750 418.050 292.050 ;
        RECT 413.550 289.950 419.850 291.750 ;
        RECT 413.550 282.600 414.750 289.950 ;
        RECT 426.150 286.200 427.050 298.800 ;
        RECT 429.150 298.800 430.050 300.900 ;
        RECT 430.950 300.300 438.450 301.500 ;
        RECT 430.950 299.700 432.750 300.300 ;
        RECT 445.050 299.400 446.850 311.400 ;
        RECT 460.800 305.400 462.600 311.400 ;
        RECT 429.150 298.500 437.550 298.800 ;
        RECT 445.950 298.500 446.850 299.400 ;
        RECT 429.150 297.900 446.850 298.500 ;
        RECT 461.400 298.050 462.600 305.400 ;
        RECT 467.550 299.400 469.350 311.400 ;
        RECT 475.050 305.400 476.850 311.400 ;
        RECT 472.950 303.300 476.850 305.400 ;
        RECT 482.850 304.500 484.650 311.400 ;
        RECT 490.650 305.400 492.450 311.400 ;
        RECT 491.250 304.500 492.450 305.400 ;
        RECT 481.950 303.450 488.550 304.500 ;
        RECT 481.950 302.700 483.750 303.450 ;
        RECT 486.750 302.700 488.550 303.450 ;
        RECT 491.250 302.400 496.050 304.500 ;
        RECT 474.150 300.600 476.850 302.400 ;
        RECT 477.750 301.800 479.550 302.400 ;
        RECT 477.750 300.900 484.050 301.800 ;
        RECT 491.250 301.500 492.450 302.400 ;
        RECT 477.750 300.600 479.550 300.900 ;
        RECT 475.950 299.700 476.850 300.600 ;
        RECT 435.750 297.300 446.850 297.900 ;
        RECT 435.750 297.000 437.550 297.300 ;
        RECT 433.950 290.400 436.050 292.050 ;
        RECT 433.950 289.200 441.900 290.400 ;
        RECT 442.950 289.950 445.050 292.050 ;
        RECT 440.100 288.600 441.900 289.200 ;
        RECT 443.100 288.150 444.900 289.950 ;
        RECT 437.100 287.400 438.900 288.000 ;
        RECT 443.100 287.400 444.000 288.150 ;
        RECT 437.100 286.200 444.000 287.400 ;
        RECT 426.150 285.000 438.150 286.200 ;
        RECT 426.150 284.400 427.950 285.000 ;
        RECT 437.100 283.200 438.150 285.000 ;
        RECT 413.550 276.600 415.350 282.600 ;
        RECT 418.950 281.700 421.050 282.600 ;
        RECT 418.950 280.500 422.700 281.700 ;
        RECT 433.350 281.550 435.150 282.300 ;
        RECT 421.650 279.600 422.700 280.500 ;
        RECT 430.200 280.500 435.150 281.550 ;
        RECT 436.650 281.400 438.450 283.200 ;
        RECT 445.950 282.600 446.850 297.300 ;
        RECT 460.950 292.950 463.050 298.050 ;
        RECT 439.950 280.500 442.050 282.600 ;
        RECT 430.200 279.600 431.250 280.500 ;
        RECT 439.950 279.600 441.000 280.500 ;
        RECT 421.650 276.600 423.450 279.600 ;
        RECT 429.450 276.600 431.250 279.600 ;
        RECT 437.250 278.700 441.000 279.600 ;
        RECT 437.250 276.600 439.050 278.700 ;
        RECT 445.050 276.600 446.850 282.600 ;
        RECT 461.400 279.600 462.600 292.950 ;
        RECT 464.100 292.050 465.900 293.850 ;
        RECT 467.550 292.050 468.750 299.400 ;
        RECT 472.950 298.800 475.050 299.700 ;
        RECT 475.950 298.800 481.050 299.700 ;
        RECT 470.850 297.600 475.050 298.800 ;
        RECT 469.950 295.800 471.750 297.600 ;
        RECT 463.950 289.950 466.050 292.050 ;
        RECT 467.550 291.750 472.050 292.050 ;
        RECT 467.550 289.950 473.850 291.750 ;
        RECT 460.800 276.600 462.600 279.600 ;
        RECT 467.550 282.600 468.750 289.950 ;
        RECT 480.150 286.200 481.050 298.800 ;
        RECT 483.150 298.800 484.050 300.900 ;
        RECT 484.950 300.300 492.450 301.500 ;
        RECT 484.950 299.700 486.750 300.300 ;
        RECT 499.050 299.400 500.850 311.400 ;
        RECT 483.150 298.500 491.550 298.800 ;
        RECT 499.950 298.500 500.850 299.400 ;
        RECT 483.150 297.900 500.850 298.500 ;
        RECT 489.750 297.300 500.850 297.900 ;
        RECT 489.750 297.000 491.550 297.300 ;
        RECT 487.950 290.400 490.050 292.050 ;
        RECT 487.950 289.200 495.900 290.400 ;
        RECT 496.950 289.950 499.050 292.050 ;
        RECT 494.100 288.600 495.900 289.200 ;
        RECT 497.100 288.150 498.900 289.950 ;
        RECT 491.100 287.400 492.900 288.000 ;
        RECT 497.100 287.400 498.000 288.150 ;
        RECT 491.100 286.200 498.000 287.400 ;
        RECT 480.150 285.000 492.150 286.200 ;
        RECT 480.150 284.400 481.950 285.000 ;
        RECT 491.100 283.200 492.150 285.000 ;
        RECT 467.550 276.600 469.350 282.600 ;
        RECT 472.950 281.700 475.050 282.600 ;
        RECT 472.950 280.500 476.700 281.700 ;
        RECT 487.350 281.550 489.150 282.300 ;
        RECT 475.650 279.600 476.700 280.500 ;
        RECT 484.200 280.500 489.150 281.550 ;
        RECT 490.650 281.400 492.450 283.200 ;
        RECT 499.950 282.600 500.850 297.300 ;
        RECT 515.400 305.400 517.200 311.400 ;
        RECT 511.950 292.950 514.050 295.050 ;
        RECT 512.100 291.150 513.900 292.950 ;
        RECT 515.400 292.050 516.600 305.400 ;
        RECT 524.550 299.400 526.350 311.400 ;
        RECT 532.050 305.400 533.850 311.400 ;
        RECT 529.950 303.300 533.850 305.400 ;
        RECT 539.850 304.500 541.650 311.400 ;
        RECT 547.650 305.400 549.450 311.400 ;
        RECT 548.250 304.500 549.450 305.400 ;
        RECT 538.950 303.450 545.550 304.500 ;
        RECT 538.950 302.700 540.750 303.450 ;
        RECT 543.750 302.700 545.550 303.450 ;
        RECT 548.250 302.400 553.050 304.500 ;
        RECT 531.150 300.600 533.850 302.400 ;
        RECT 534.750 301.800 536.550 302.400 ;
        RECT 534.750 300.900 541.050 301.800 ;
        RECT 548.250 301.500 549.450 302.400 ;
        RECT 534.750 300.600 536.550 300.900 ;
        RECT 532.950 299.700 533.850 300.600 ;
        RECT 517.950 292.950 520.050 295.050 ;
        RECT 514.950 289.950 517.050 292.050 ;
        RECT 518.100 291.150 519.900 292.950 ;
        RECT 524.550 292.050 525.750 299.400 ;
        RECT 529.950 298.800 532.050 299.700 ;
        RECT 532.950 298.800 538.050 299.700 ;
        RECT 527.850 297.600 532.050 298.800 ;
        RECT 526.950 295.800 528.750 297.600 ;
        RECT 524.550 291.750 529.050 292.050 ;
        RECT 524.550 289.950 530.850 291.750 ;
        RECT 515.400 284.700 516.600 289.950 ;
        RECT 515.400 283.800 519.600 284.700 ;
        RECT 493.950 280.500 496.050 282.600 ;
        RECT 484.200 279.600 485.250 280.500 ;
        RECT 493.950 279.600 495.000 280.500 ;
        RECT 475.650 276.600 477.450 279.600 ;
        RECT 483.450 276.600 485.250 279.600 ;
        RECT 491.250 278.700 495.000 279.600 ;
        RECT 491.250 276.600 493.050 278.700 ;
        RECT 499.050 276.600 500.850 282.600 ;
        RECT 517.800 276.600 519.600 283.800 ;
        RECT 524.550 282.600 525.750 289.950 ;
        RECT 537.150 286.200 538.050 298.800 ;
        RECT 540.150 298.800 541.050 300.900 ;
        RECT 541.950 300.300 549.450 301.500 ;
        RECT 541.950 299.700 543.750 300.300 ;
        RECT 556.050 299.400 557.850 311.400 ;
        RECT 540.150 298.500 548.550 298.800 ;
        RECT 556.950 298.500 557.850 299.400 ;
        RECT 574.800 298.500 576.600 311.400 ;
        RECT 580.800 298.500 582.600 311.400 ;
        RECT 586.800 298.500 588.600 311.400 ;
        RECT 592.800 298.500 594.600 311.400 ;
        RECT 613.800 305.400 615.600 311.400 ;
        RECT 540.150 297.900 557.850 298.500 ;
        RECT 546.750 297.300 557.850 297.900 ;
        RECT 546.750 297.000 548.550 297.300 ;
        RECT 544.950 290.400 547.050 292.050 ;
        RECT 544.950 289.200 552.900 290.400 ;
        RECT 553.950 289.950 556.050 292.050 ;
        RECT 551.100 288.600 552.900 289.200 ;
        RECT 554.100 288.150 555.900 289.950 ;
        RECT 548.100 287.400 549.900 288.000 ;
        RECT 554.100 287.400 555.000 288.150 ;
        RECT 548.100 286.200 555.000 287.400 ;
        RECT 537.150 285.000 549.150 286.200 ;
        RECT 537.150 284.400 538.950 285.000 ;
        RECT 548.100 283.200 549.150 285.000 ;
        RECT 524.550 276.600 526.350 282.600 ;
        RECT 529.950 281.700 532.050 282.600 ;
        RECT 529.950 280.500 533.700 281.700 ;
        RECT 544.350 281.550 546.150 282.300 ;
        RECT 532.650 279.600 533.700 280.500 ;
        RECT 541.200 280.500 546.150 281.550 ;
        RECT 547.650 281.400 549.450 283.200 ;
        RECT 556.950 282.600 557.850 297.300 ;
        RECT 573.900 297.300 576.600 298.500 ;
        RECT 578.700 297.300 582.600 298.500 ;
        RECT 584.700 297.300 588.600 298.500 ;
        RECT 590.700 297.300 594.600 298.500 ;
        RECT 573.900 292.050 574.800 297.300 ;
        RECT 571.950 289.950 574.800 292.050 ;
        RECT 573.900 284.700 574.800 289.950 ;
        RECT 575.700 286.800 577.500 287.400 ;
        RECT 578.700 286.800 579.900 297.300 ;
        RECT 575.700 285.600 579.900 286.800 ;
        RECT 581.700 286.800 583.500 287.400 ;
        RECT 584.700 286.800 585.900 297.300 ;
        RECT 581.700 285.600 585.900 286.800 ;
        RECT 587.700 286.800 589.500 287.400 ;
        RECT 590.700 286.800 591.900 297.300 ;
        RECT 608.100 292.050 609.900 293.850 ;
        RECT 610.950 292.950 613.050 295.050 ;
        RECT 592.950 289.950 595.050 292.050 ;
        RECT 607.950 289.950 610.050 292.050 ;
        RECT 611.100 291.150 612.900 292.950 ;
        RECT 613.950 292.050 615.150 305.400 ;
        RECT 624.150 299.400 625.950 311.400 ;
        RECT 632.550 305.400 634.350 311.400 ;
        RECT 632.550 304.500 633.750 305.400 ;
        RECT 640.350 304.500 642.150 311.400 ;
        RECT 648.150 305.400 649.950 311.400 ;
        RECT 628.950 302.400 633.750 304.500 ;
        RECT 636.450 303.450 643.050 304.500 ;
        RECT 636.450 302.700 638.250 303.450 ;
        RECT 641.250 302.700 643.050 303.450 ;
        RECT 648.150 303.300 652.050 305.400 ;
        RECT 632.550 301.500 633.750 302.400 ;
        RECT 645.450 301.800 647.250 302.400 ;
        RECT 632.550 300.300 640.050 301.500 ;
        RECT 638.250 299.700 640.050 300.300 ;
        RECT 640.950 300.900 647.250 301.800 ;
        RECT 624.150 298.500 625.050 299.400 ;
        RECT 640.950 298.800 641.850 300.900 ;
        RECT 645.450 300.600 647.250 300.900 ;
        RECT 648.150 300.600 650.850 302.400 ;
        RECT 648.150 299.700 649.050 300.600 ;
        RECT 633.450 298.500 641.850 298.800 ;
        RECT 624.150 297.900 641.850 298.500 ;
        RECT 643.950 298.800 649.050 299.700 ;
        RECT 649.950 298.800 652.050 299.700 ;
        RECT 655.650 299.400 657.450 311.400 ;
        RECT 624.150 297.300 635.250 297.900 ;
        RECT 616.950 292.950 619.050 295.050 ;
        RECT 613.950 289.950 616.050 292.050 ;
        RECT 617.100 291.150 618.900 292.950 ;
        RECT 593.100 288.150 594.900 289.950 ;
        RECT 587.700 285.600 591.900 286.800 ;
        RECT 578.700 284.700 579.900 285.600 ;
        RECT 584.700 284.700 585.900 285.600 ;
        RECT 590.700 284.700 591.900 285.600 ;
        RECT 614.850 285.750 616.050 289.950 ;
        RECT 614.850 284.700 618.600 285.750 ;
        RECT 573.900 283.500 576.600 284.700 ;
        RECT 578.700 283.500 582.600 284.700 ;
        RECT 584.700 283.500 588.600 284.700 ;
        RECT 590.700 283.500 594.600 284.700 ;
        RECT 550.950 280.500 553.050 282.600 ;
        RECT 541.200 279.600 542.250 280.500 ;
        RECT 550.950 279.600 552.000 280.500 ;
        RECT 532.650 276.600 534.450 279.600 ;
        RECT 540.450 276.600 542.250 279.600 ;
        RECT 548.250 278.700 552.000 279.600 ;
        RECT 548.250 276.600 550.050 278.700 ;
        RECT 556.050 276.600 557.850 282.600 ;
        RECT 574.800 276.600 576.600 283.500 ;
        RECT 580.800 276.600 582.600 283.500 ;
        RECT 586.800 276.600 588.600 283.500 ;
        RECT 592.800 276.600 594.600 283.500 ;
        RECT 608.400 281.700 616.200 283.050 ;
        RECT 608.400 276.600 610.200 281.700 ;
        RECT 614.400 276.600 616.200 281.700 ;
        RECT 617.400 282.600 618.600 284.700 ;
        RECT 624.150 282.600 625.050 297.300 ;
        RECT 633.450 297.000 635.250 297.300 ;
        RECT 625.950 289.950 628.050 292.050 ;
        RECT 634.950 290.400 637.050 292.050 ;
        RECT 626.100 288.150 627.900 289.950 ;
        RECT 629.100 289.200 637.050 290.400 ;
        RECT 629.100 288.600 630.900 289.200 ;
        RECT 627.000 287.400 627.900 288.150 ;
        RECT 632.100 287.400 633.900 288.000 ;
        RECT 627.000 286.200 633.900 287.400 ;
        RECT 643.950 286.200 644.850 298.800 ;
        RECT 649.950 297.600 654.150 298.800 ;
        RECT 653.250 295.800 655.050 297.600 ;
        RECT 656.250 292.050 657.450 299.400 ;
        RECT 671.400 305.400 673.200 311.400 ;
        RECT 667.950 292.950 670.050 295.050 ;
        RECT 652.950 291.750 657.450 292.050 ;
        RECT 651.150 289.950 657.450 291.750 ;
        RECT 668.100 291.150 669.900 292.950 ;
        RECT 671.400 292.050 672.600 305.400 ;
        RECT 680.550 299.400 682.350 311.400 ;
        RECT 688.050 305.400 689.850 311.400 ;
        RECT 685.950 303.300 689.850 305.400 ;
        RECT 695.850 304.500 697.650 311.400 ;
        RECT 703.650 305.400 705.450 311.400 ;
        RECT 704.250 304.500 705.450 305.400 ;
        RECT 694.950 303.450 701.550 304.500 ;
        RECT 694.950 302.700 696.750 303.450 ;
        RECT 699.750 302.700 701.550 303.450 ;
        RECT 704.250 302.400 709.050 304.500 ;
        RECT 687.150 300.600 689.850 302.400 ;
        RECT 690.750 301.800 692.550 302.400 ;
        RECT 690.750 300.900 697.050 301.800 ;
        RECT 704.250 301.500 705.450 302.400 ;
        RECT 690.750 300.600 692.550 300.900 ;
        RECT 688.950 299.700 689.850 300.600 ;
        RECT 673.950 292.950 676.050 295.050 ;
        RECT 670.950 289.950 673.050 292.050 ;
        RECT 674.100 291.150 675.900 292.950 ;
        RECT 680.550 292.050 681.750 299.400 ;
        RECT 685.950 298.800 688.050 299.700 ;
        RECT 688.950 298.800 694.050 299.700 ;
        RECT 683.850 297.600 688.050 298.800 ;
        RECT 682.950 295.800 684.750 297.600 ;
        RECT 680.550 291.750 685.050 292.050 ;
        RECT 680.550 289.950 686.850 291.750 ;
        RECT 632.850 285.000 644.850 286.200 ;
        RECT 632.850 283.200 633.900 285.000 ;
        RECT 643.050 284.400 644.850 285.000 ;
        RECT 617.400 276.600 619.200 282.600 ;
        RECT 624.150 276.600 625.950 282.600 ;
        RECT 628.950 280.500 631.050 282.600 ;
        RECT 632.550 281.400 634.350 283.200 ;
        RECT 656.250 282.600 657.450 289.950 ;
        RECT 671.400 284.700 672.600 289.950 ;
        RECT 671.400 283.800 675.600 284.700 ;
        RECT 635.850 281.550 637.650 282.300 ;
        RECT 649.950 281.700 652.050 282.600 ;
        RECT 635.850 280.500 640.800 281.550 ;
        RECT 630.000 279.600 631.050 280.500 ;
        RECT 639.750 279.600 640.800 280.500 ;
        RECT 648.300 280.500 652.050 281.700 ;
        RECT 648.300 279.600 649.350 280.500 ;
        RECT 630.000 278.700 633.750 279.600 ;
        RECT 631.950 276.600 633.750 278.700 ;
        RECT 639.750 276.600 641.550 279.600 ;
        RECT 647.550 276.600 649.350 279.600 ;
        RECT 655.650 276.600 657.450 282.600 ;
        RECT 673.800 276.600 675.600 283.800 ;
        RECT 680.550 282.600 681.750 289.950 ;
        RECT 693.150 286.200 694.050 298.800 ;
        RECT 696.150 298.800 697.050 300.900 ;
        RECT 697.950 300.300 705.450 301.500 ;
        RECT 697.950 299.700 699.750 300.300 ;
        RECT 712.050 299.400 713.850 311.400 ;
        RECT 696.150 298.500 704.550 298.800 ;
        RECT 712.950 298.500 713.850 299.400 ;
        RECT 696.150 297.900 713.850 298.500 ;
        RECT 702.750 297.300 713.850 297.900 ;
        RECT 702.750 297.000 704.550 297.300 ;
        RECT 700.950 290.400 703.050 292.050 ;
        RECT 700.950 289.200 708.900 290.400 ;
        RECT 709.950 289.950 712.050 292.050 ;
        RECT 707.100 288.600 708.900 289.200 ;
        RECT 710.100 288.150 711.900 289.950 ;
        RECT 704.100 287.400 705.900 288.000 ;
        RECT 710.100 287.400 711.000 288.150 ;
        RECT 704.100 286.200 711.000 287.400 ;
        RECT 693.150 285.000 705.150 286.200 ;
        RECT 693.150 284.400 694.950 285.000 ;
        RECT 704.100 283.200 705.150 285.000 ;
        RECT 680.550 276.600 682.350 282.600 ;
        RECT 685.950 281.700 688.050 282.600 ;
        RECT 685.950 280.500 689.700 281.700 ;
        RECT 700.350 281.550 702.150 282.300 ;
        RECT 688.650 279.600 689.700 280.500 ;
        RECT 697.200 280.500 702.150 281.550 ;
        RECT 703.650 281.400 705.450 283.200 ;
        RECT 712.950 282.600 713.850 297.300 ;
        RECT 728.400 305.400 730.200 311.400 ;
        RECT 724.950 292.950 727.050 295.050 ;
        RECT 725.100 291.150 726.900 292.950 ;
        RECT 728.400 292.050 729.600 305.400 ;
        RECT 738.150 299.400 739.950 311.400 ;
        RECT 746.550 305.400 748.350 311.400 ;
        RECT 746.550 304.500 747.750 305.400 ;
        RECT 754.350 304.500 756.150 311.400 ;
        RECT 762.150 305.400 763.950 311.400 ;
        RECT 742.950 302.400 747.750 304.500 ;
        RECT 750.450 303.450 757.050 304.500 ;
        RECT 750.450 302.700 752.250 303.450 ;
        RECT 755.250 302.700 757.050 303.450 ;
        RECT 762.150 303.300 766.050 305.400 ;
        RECT 746.550 301.500 747.750 302.400 ;
        RECT 759.450 301.800 761.250 302.400 ;
        RECT 746.550 300.300 754.050 301.500 ;
        RECT 752.250 299.700 754.050 300.300 ;
        RECT 754.950 300.900 761.250 301.800 ;
        RECT 738.150 298.500 739.050 299.400 ;
        RECT 754.950 298.800 755.850 300.900 ;
        RECT 759.450 300.600 761.250 300.900 ;
        RECT 762.150 300.600 764.850 302.400 ;
        RECT 762.150 299.700 763.050 300.600 ;
        RECT 747.450 298.500 755.850 298.800 ;
        RECT 738.150 297.900 755.850 298.500 ;
        RECT 757.950 298.800 763.050 299.700 ;
        RECT 763.950 298.800 766.050 299.700 ;
        RECT 769.650 299.400 771.450 311.400 ;
        RECT 788.400 305.400 790.200 311.400 ;
        RECT 738.150 297.300 749.250 297.900 ;
        RECT 730.950 292.950 733.050 295.050 ;
        RECT 727.950 289.950 730.050 292.050 ;
        RECT 731.100 291.150 732.900 292.950 ;
        RECT 728.400 284.700 729.600 289.950 ;
        RECT 728.400 283.800 732.600 284.700 ;
        RECT 706.950 280.500 709.050 282.600 ;
        RECT 697.200 279.600 698.250 280.500 ;
        RECT 706.950 279.600 708.000 280.500 ;
        RECT 688.650 276.600 690.450 279.600 ;
        RECT 696.450 276.600 698.250 279.600 ;
        RECT 704.250 278.700 708.000 279.600 ;
        RECT 704.250 276.600 706.050 278.700 ;
        RECT 712.050 276.600 713.850 282.600 ;
        RECT 730.800 276.600 732.600 283.800 ;
        RECT 738.150 282.600 739.050 297.300 ;
        RECT 747.450 297.000 749.250 297.300 ;
        RECT 739.950 289.950 742.050 292.050 ;
        RECT 748.950 290.400 751.050 292.050 ;
        RECT 740.100 288.150 741.900 289.950 ;
        RECT 743.100 289.200 751.050 290.400 ;
        RECT 743.100 288.600 744.900 289.200 ;
        RECT 741.000 287.400 741.900 288.150 ;
        RECT 746.100 287.400 747.900 288.000 ;
        RECT 741.000 286.200 747.900 287.400 ;
        RECT 757.950 286.200 758.850 298.800 ;
        RECT 763.950 297.600 768.150 298.800 ;
        RECT 767.250 295.800 769.050 297.600 ;
        RECT 770.250 292.050 771.450 299.400 ;
        RECT 784.950 292.950 787.050 295.050 ;
        RECT 766.950 291.750 771.450 292.050 ;
        RECT 765.150 289.950 771.450 291.750 ;
        RECT 785.100 291.150 786.900 292.950 ;
        RECT 788.850 292.050 790.050 305.400 ;
        RECT 809.700 300.600 811.500 311.400 ;
        RECT 809.700 299.400 813.300 300.600 ;
        RECT 790.950 292.950 793.050 295.050 ;
        RECT 746.850 285.000 758.850 286.200 ;
        RECT 746.850 283.200 747.900 285.000 ;
        RECT 757.050 284.400 758.850 285.000 ;
        RECT 738.150 276.600 739.950 282.600 ;
        RECT 742.950 280.500 745.050 282.600 ;
        RECT 746.550 281.400 748.350 283.200 ;
        RECT 770.250 282.600 771.450 289.950 ;
        RECT 787.950 289.950 790.050 292.050 ;
        RECT 791.100 291.150 792.900 292.950 ;
        RECT 794.100 292.050 795.900 293.850 ;
        RECT 812.400 292.050 813.300 299.400 ;
        RECT 819.150 299.400 820.950 311.400 ;
        RECT 827.550 305.400 829.350 311.400 ;
        RECT 827.550 304.500 828.750 305.400 ;
        RECT 835.350 304.500 837.150 311.400 ;
        RECT 843.150 305.400 844.950 311.400 ;
        RECT 823.950 302.400 828.750 304.500 ;
        RECT 831.450 303.450 838.050 304.500 ;
        RECT 831.450 302.700 833.250 303.450 ;
        RECT 836.250 302.700 838.050 303.450 ;
        RECT 843.150 303.300 847.050 305.400 ;
        RECT 827.550 301.500 828.750 302.400 ;
        RECT 840.450 301.800 842.250 302.400 ;
        RECT 827.550 300.300 835.050 301.500 ;
        RECT 833.250 299.700 835.050 300.300 ;
        RECT 835.950 300.900 842.250 301.800 ;
        RECT 819.150 298.500 820.050 299.400 ;
        RECT 835.950 298.800 836.850 300.900 ;
        RECT 840.450 300.600 842.250 300.900 ;
        RECT 843.150 300.600 845.850 302.400 ;
        RECT 843.150 299.700 844.050 300.600 ;
        RECT 828.450 298.500 836.850 298.800 ;
        RECT 819.150 297.900 836.850 298.500 ;
        RECT 838.950 298.800 844.050 299.700 ;
        RECT 844.950 298.800 847.050 299.700 ;
        RECT 850.650 299.400 852.450 311.400 ;
        RECT 819.150 297.300 830.250 297.900 ;
        RECT 793.950 289.950 796.050 292.050 ;
        RECT 787.950 285.750 789.150 289.950 ;
        RECT 809.100 289.050 810.900 290.850 ;
        RECT 811.950 289.950 814.050 292.050 ;
        RECT 808.950 286.950 811.050 289.050 ;
        RECT 785.400 284.700 789.150 285.750 ;
        RECT 785.400 282.600 786.600 284.700 ;
        RECT 749.850 281.550 751.650 282.300 ;
        RECT 763.950 281.700 766.050 282.600 ;
        RECT 749.850 280.500 754.800 281.550 ;
        RECT 744.000 279.600 745.050 280.500 ;
        RECT 753.750 279.600 754.800 280.500 ;
        RECT 762.300 280.500 766.050 281.700 ;
        RECT 762.300 279.600 763.350 280.500 ;
        RECT 744.000 278.700 747.750 279.600 ;
        RECT 745.950 276.600 747.750 278.700 ;
        RECT 753.750 276.600 755.550 279.600 ;
        RECT 761.550 276.600 763.350 279.600 ;
        RECT 769.650 276.600 771.450 282.600 ;
        RECT 784.800 276.600 786.600 282.600 ;
        RECT 787.800 281.700 795.600 283.050 ;
        RECT 787.800 276.600 789.600 281.700 ;
        RECT 793.800 276.600 795.600 281.700 ;
        RECT 812.400 279.600 813.300 289.950 ;
        RECT 815.100 289.050 816.900 290.850 ;
        RECT 814.950 286.950 817.050 289.050 ;
        RECT 819.150 282.600 820.050 297.300 ;
        RECT 828.450 297.000 830.250 297.300 ;
        RECT 820.950 289.950 823.050 292.050 ;
        RECT 829.950 290.400 832.050 292.050 ;
        RECT 821.100 288.150 822.900 289.950 ;
        RECT 824.100 289.200 832.050 290.400 ;
        RECT 824.100 288.600 825.900 289.200 ;
        RECT 822.000 287.400 822.900 288.150 ;
        RECT 827.100 287.400 828.900 288.000 ;
        RECT 822.000 286.200 828.900 287.400 ;
        RECT 838.950 286.200 839.850 298.800 ;
        RECT 844.950 297.600 849.150 298.800 ;
        RECT 848.250 295.800 850.050 297.600 ;
        RECT 851.250 292.050 852.450 299.400 ;
        RECT 866.400 298.500 868.200 311.400 ;
        RECT 872.400 298.500 874.200 311.400 ;
        RECT 878.400 298.500 880.200 311.400 ;
        RECT 884.400 298.500 886.200 311.400 ;
        RECT 866.400 297.300 870.300 298.500 ;
        RECT 872.400 297.300 876.300 298.500 ;
        RECT 878.400 297.300 882.300 298.500 ;
        RECT 884.400 297.300 887.100 298.500 ;
        RECT 847.950 291.750 852.450 292.050 ;
        RECT 846.150 289.950 852.450 291.750 ;
        RECT 865.950 289.950 868.050 292.050 ;
        RECT 827.850 285.000 839.850 286.200 ;
        RECT 827.850 283.200 828.900 285.000 ;
        RECT 838.050 284.400 839.850 285.000 ;
        RECT 811.800 276.600 813.600 279.600 ;
        RECT 819.150 276.600 820.950 282.600 ;
        RECT 823.950 280.500 826.050 282.600 ;
        RECT 827.550 281.400 829.350 283.200 ;
        RECT 851.250 282.600 852.450 289.950 ;
        RECT 866.100 288.150 867.900 289.950 ;
        RECT 869.100 286.800 870.300 297.300 ;
        RECT 871.500 286.800 873.300 287.400 ;
        RECT 869.100 285.600 873.300 286.800 ;
        RECT 875.100 286.800 876.300 297.300 ;
        RECT 877.500 286.800 879.300 287.400 ;
        RECT 875.100 285.600 879.300 286.800 ;
        RECT 881.100 286.800 882.300 297.300 ;
        RECT 886.200 292.050 887.100 297.300 ;
        RECT 886.200 289.950 889.050 292.050 ;
        RECT 883.500 286.800 885.300 287.400 ;
        RECT 881.100 285.600 885.300 286.800 ;
        RECT 869.100 284.700 870.300 285.600 ;
        RECT 875.100 284.700 876.300 285.600 ;
        RECT 881.100 284.700 882.300 285.600 ;
        RECT 886.200 284.700 887.100 289.950 ;
        RECT 830.850 281.550 832.650 282.300 ;
        RECT 844.950 281.700 847.050 282.600 ;
        RECT 830.850 280.500 835.800 281.550 ;
        RECT 825.000 279.600 826.050 280.500 ;
        RECT 834.750 279.600 835.800 280.500 ;
        RECT 843.300 280.500 847.050 281.700 ;
        RECT 843.300 279.600 844.350 280.500 ;
        RECT 825.000 278.700 828.750 279.600 ;
        RECT 826.950 276.600 828.750 278.700 ;
        RECT 834.750 276.600 836.550 279.600 ;
        RECT 842.550 276.600 844.350 279.600 ;
        RECT 850.650 276.600 852.450 282.600 ;
        RECT 866.400 283.500 870.300 284.700 ;
        RECT 872.400 283.500 876.300 284.700 ;
        RECT 878.400 283.500 882.300 284.700 ;
        RECT 884.400 283.500 887.100 284.700 ;
        RECT 866.400 276.600 868.200 283.500 ;
        RECT 872.400 276.600 874.200 283.500 ;
        RECT 878.400 276.600 880.200 283.500 ;
        RECT 884.400 276.600 886.200 283.500 ;
        RECT 16.800 269.400 18.600 272.400 ;
        RECT 13.950 259.950 16.050 262.050 ;
        RECT 14.100 258.150 15.900 259.950 ;
        RECT 17.400 259.050 18.300 269.400 ;
        RECT 28.950 268.950 31.050 271.050 ;
        RECT 34.800 269.400 36.600 272.400 ;
        RECT 19.950 259.950 22.050 262.050 ;
        RECT 16.950 256.950 19.050 259.050 ;
        RECT 20.100 258.150 21.900 259.950 ;
        RECT 17.400 249.600 18.300 256.950 ;
        RECT 14.700 248.400 18.300 249.600 ;
        RECT 14.700 237.600 16.500 248.400 ;
        RECT 29.550 247.050 30.450 268.950 ;
        RECT 35.400 256.050 36.600 269.400 ;
        RECT 41.550 266.400 43.350 272.400 ;
        RECT 49.650 269.400 51.450 272.400 ;
        RECT 57.450 269.400 59.250 272.400 ;
        RECT 65.250 270.300 67.050 272.400 ;
        RECT 65.250 269.400 69.000 270.300 ;
        RECT 49.650 268.500 50.700 269.400 ;
        RECT 46.950 267.300 50.700 268.500 ;
        RECT 58.200 268.500 59.250 269.400 ;
        RECT 67.950 268.500 69.000 269.400 ;
        RECT 58.200 267.450 63.150 268.500 ;
        RECT 46.950 266.400 49.050 267.300 ;
        RECT 61.350 266.700 63.150 267.450 ;
        RECT 41.550 259.050 42.750 266.400 ;
        RECT 64.650 265.800 66.450 267.600 ;
        RECT 67.950 266.400 70.050 268.500 ;
        RECT 73.050 266.400 74.850 272.400 ;
        RECT 54.150 264.000 55.950 264.600 ;
        RECT 65.100 264.000 66.150 265.800 ;
        RECT 54.150 262.800 66.150 264.000 ;
        RECT 37.950 256.950 40.050 259.050 ;
        RECT 41.550 257.250 47.850 259.050 ;
        RECT 41.550 256.950 46.050 257.250 ;
        RECT 34.950 250.950 37.050 256.050 ;
        RECT 38.100 255.150 39.900 256.950 ;
        RECT 28.950 244.950 31.050 247.050 ;
        RECT 35.400 243.600 36.600 250.950 ;
        RECT 34.800 237.600 36.600 243.600 ;
        RECT 41.550 249.600 42.750 256.950 ;
        RECT 43.950 251.400 45.750 253.200 ;
        RECT 44.850 250.200 49.050 251.400 ;
        RECT 54.150 250.200 55.050 262.800 ;
        RECT 65.100 261.600 72.000 262.800 ;
        RECT 65.100 261.000 66.900 261.600 ;
        RECT 71.100 260.850 72.000 261.600 ;
        RECT 68.100 259.800 69.900 260.400 ;
        RECT 61.950 258.600 69.900 259.800 ;
        RECT 71.100 259.050 72.900 260.850 ;
        RECT 61.950 256.950 64.050 258.600 ;
        RECT 70.950 256.950 73.050 259.050 ;
        RECT 63.750 251.700 65.550 252.000 ;
        RECT 73.950 251.700 74.850 266.400 ;
        RECT 86.400 267.300 88.200 272.400 ;
        RECT 92.400 267.300 94.200 272.400 ;
        RECT 86.400 265.950 94.200 267.300 ;
        RECT 95.400 266.400 97.200 272.400 ;
        RECT 115.800 269.400 117.600 272.400 ;
        RECT 133.800 269.400 135.600 272.400 ;
        RECT 95.400 264.300 96.600 266.400 ;
        RECT 92.850 263.250 96.600 264.300 ;
        RECT 92.850 259.050 94.050 263.250 ;
        RECT 112.950 259.950 115.050 262.050 ;
        RECT 85.950 256.950 88.050 259.050 ;
        RECT 86.100 255.150 87.900 256.950 ;
        RECT 89.100 256.050 90.900 257.850 ;
        RECT 91.950 256.950 94.050 259.050 ;
        RECT 113.100 258.150 114.900 259.950 ;
        RECT 116.400 259.050 117.300 269.400 ;
        RECT 118.950 259.950 121.050 262.050 ;
        RECT 88.950 253.950 91.050 256.050 ;
        RECT 63.750 251.100 74.850 251.700 ;
        RECT 41.550 237.600 43.350 249.600 ;
        RECT 46.950 249.300 49.050 250.200 ;
        RECT 49.950 249.300 55.050 250.200 ;
        RECT 57.150 250.500 74.850 251.100 ;
        RECT 57.150 250.200 65.550 250.500 ;
        RECT 49.950 248.400 50.850 249.300 ;
        RECT 48.150 246.600 50.850 248.400 ;
        RECT 51.750 248.100 53.550 248.400 ;
        RECT 57.150 248.100 58.050 250.200 ;
        RECT 73.950 249.600 74.850 250.500 ;
        RECT 51.750 247.200 58.050 248.100 ;
        RECT 58.950 248.700 60.750 249.300 ;
        RECT 58.950 247.500 66.450 248.700 ;
        RECT 51.750 246.600 53.550 247.200 ;
        RECT 65.250 246.600 66.450 247.500 ;
        RECT 46.950 243.600 50.850 245.700 ;
        RECT 55.950 245.550 57.750 246.300 ;
        RECT 60.750 245.550 62.550 246.300 ;
        RECT 55.950 244.500 62.550 245.550 ;
        RECT 65.250 244.500 70.050 246.600 ;
        RECT 49.050 237.600 50.850 243.600 ;
        RECT 56.850 237.600 58.650 244.500 ;
        RECT 65.250 243.600 66.450 244.500 ;
        RECT 64.650 237.600 66.450 243.600 ;
        RECT 73.050 237.600 74.850 249.600 ;
        RECT 91.950 243.600 93.150 256.950 ;
        RECT 95.100 256.050 96.900 257.850 ;
        RECT 115.950 256.950 118.050 259.050 ;
        RECT 119.100 258.150 120.900 259.950 ;
        RECT 94.950 253.950 97.050 256.050 ;
        RECT 116.400 249.600 117.300 256.950 ;
        RECT 134.400 256.050 135.600 269.400 ;
        RECT 140.550 266.400 142.350 272.400 ;
        RECT 148.650 269.400 150.450 272.400 ;
        RECT 156.450 269.400 158.250 272.400 ;
        RECT 164.250 270.300 166.050 272.400 ;
        RECT 164.250 269.400 168.000 270.300 ;
        RECT 148.650 268.500 149.700 269.400 ;
        RECT 145.950 267.300 149.700 268.500 ;
        RECT 157.200 268.500 158.250 269.400 ;
        RECT 166.950 268.500 168.000 269.400 ;
        RECT 157.200 267.450 162.150 268.500 ;
        RECT 145.950 266.400 148.050 267.300 ;
        RECT 160.350 266.700 162.150 267.450 ;
        RECT 140.550 259.050 141.750 266.400 ;
        RECT 163.650 265.800 165.450 267.600 ;
        RECT 166.950 266.400 169.050 268.500 ;
        RECT 172.050 266.400 173.850 272.400 ;
        RECT 153.150 264.000 154.950 264.600 ;
        RECT 164.100 264.000 165.150 265.800 ;
        RECT 153.150 262.800 165.150 264.000 ;
        RECT 136.950 256.950 139.050 259.050 ;
        RECT 140.550 257.250 146.850 259.050 ;
        RECT 140.550 256.950 145.050 257.250 ;
        RECT 133.950 250.950 136.050 256.050 ;
        RECT 137.100 255.150 138.900 256.950 ;
        RECT 113.700 248.400 117.300 249.600 ;
        RECT 91.800 237.600 93.600 243.600 ;
        RECT 113.700 237.600 115.500 248.400 ;
        RECT 134.400 243.600 135.600 250.950 ;
        RECT 133.800 237.600 135.600 243.600 ;
        RECT 140.550 249.600 141.750 256.950 ;
        RECT 142.950 251.400 144.750 253.200 ;
        RECT 143.850 250.200 148.050 251.400 ;
        RECT 153.150 250.200 154.050 262.800 ;
        RECT 164.100 261.600 171.000 262.800 ;
        RECT 164.100 261.000 165.900 261.600 ;
        RECT 170.100 260.850 171.000 261.600 ;
        RECT 167.100 259.800 168.900 260.400 ;
        RECT 160.950 258.600 168.900 259.800 ;
        RECT 170.100 259.050 171.900 260.850 ;
        RECT 160.950 256.950 163.050 258.600 ;
        RECT 169.950 256.950 172.050 259.050 ;
        RECT 162.750 251.700 164.550 252.000 ;
        RECT 172.950 251.700 173.850 266.400 ;
        RECT 185.400 267.300 187.200 272.400 ;
        RECT 191.400 267.300 193.200 272.400 ;
        RECT 185.400 265.950 193.200 267.300 ;
        RECT 194.400 266.400 196.200 272.400 ;
        RECT 212.400 269.400 214.200 272.400 ;
        RECT 194.400 264.300 195.600 266.400 ;
        RECT 191.850 263.250 195.600 264.300 ;
        RECT 191.850 259.050 193.050 263.250 ;
        RECT 184.950 256.950 187.050 259.050 ;
        RECT 185.100 255.150 186.900 256.950 ;
        RECT 188.100 256.050 189.900 257.850 ;
        RECT 190.950 256.950 193.050 259.050 ;
        RECT 187.950 253.950 190.050 256.050 ;
        RECT 162.750 251.100 173.850 251.700 ;
        RECT 140.550 237.600 142.350 249.600 ;
        RECT 145.950 249.300 148.050 250.200 ;
        RECT 148.950 249.300 154.050 250.200 ;
        RECT 156.150 250.500 173.850 251.100 ;
        RECT 156.150 250.200 164.550 250.500 ;
        RECT 148.950 248.400 149.850 249.300 ;
        RECT 147.150 246.600 149.850 248.400 ;
        RECT 150.750 248.100 152.550 248.400 ;
        RECT 156.150 248.100 157.050 250.200 ;
        RECT 172.950 249.600 173.850 250.500 ;
        RECT 150.750 247.200 157.050 248.100 ;
        RECT 157.950 248.700 159.750 249.300 ;
        RECT 157.950 247.500 165.450 248.700 ;
        RECT 150.750 246.600 152.550 247.200 ;
        RECT 164.250 246.600 165.450 247.500 ;
        RECT 145.950 243.600 149.850 245.700 ;
        RECT 154.950 245.550 156.750 246.300 ;
        RECT 159.750 245.550 161.550 246.300 ;
        RECT 154.950 244.500 161.550 245.550 ;
        RECT 164.250 244.500 169.050 246.600 ;
        RECT 148.050 237.600 149.850 243.600 ;
        RECT 155.850 237.600 157.650 244.500 ;
        RECT 164.250 243.600 165.450 244.500 ;
        RECT 163.650 237.600 165.450 243.600 ;
        RECT 172.050 237.600 173.850 249.600 ;
        RECT 190.950 243.600 192.150 256.950 ;
        RECT 194.100 256.050 195.900 257.850 ;
        RECT 208.950 256.950 211.050 259.050 ;
        RECT 193.950 253.950 196.050 256.050 ;
        RECT 209.100 255.150 210.900 256.950 ;
        RECT 212.400 256.050 213.600 269.400 ;
        RECT 230.400 265.200 232.200 272.400 ;
        RECT 253.800 265.200 255.600 272.400 ;
        RECT 271.800 266.400 273.600 272.400 ;
        RECT 230.400 264.300 234.600 265.200 ;
        RECT 233.400 259.050 234.600 264.300 ;
        RECT 251.400 264.300 255.600 265.200 ;
        RECT 272.400 264.300 273.600 266.400 ;
        RECT 274.800 267.300 276.600 272.400 ;
        RECT 280.800 267.300 282.600 272.400 ;
        RECT 274.800 265.950 282.600 267.300 ;
        RECT 284.550 266.400 286.350 272.400 ;
        RECT 292.650 269.400 294.450 272.400 ;
        RECT 300.450 269.400 302.250 272.400 ;
        RECT 308.250 270.300 310.050 272.400 ;
        RECT 308.250 269.400 312.000 270.300 ;
        RECT 292.650 268.500 293.700 269.400 ;
        RECT 289.950 267.300 293.700 268.500 ;
        RECT 301.200 268.500 302.250 269.400 ;
        RECT 310.950 268.500 312.000 269.400 ;
        RECT 301.200 267.450 306.150 268.500 ;
        RECT 289.950 266.400 292.050 267.300 ;
        RECT 304.350 266.700 306.150 267.450 ;
        RECT 241.950 259.950 244.050 262.050 ;
        RECT 230.100 256.050 231.900 257.850 ;
        RECT 232.950 256.950 235.050 259.050 ;
        RECT 196.950 250.950 199.050 253.050 ;
        RECT 211.950 250.950 214.050 256.050 ;
        RECT 229.950 253.950 232.050 256.050 ;
        RECT 197.550 247.050 198.450 250.950 ;
        RECT 197.100 244.950 199.200 247.050 ;
        RECT 212.400 243.600 213.600 250.950 ;
        RECT 233.400 243.600 234.600 256.950 ;
        RECT 236.100 256.050 237.900 257.850 ;
        RECT 235.950 253.950 238.050 256.050 ;
        RECT 242.550 247.050 243.450 259.950 ;
        RECT 251.400 259.050 252.600 264.300 ;
        RECT 272.400 263.250 276.150 264.300 ;
        RECT 274.950 259.050 276.150 263.250 ;
        RECT 284.550 259.050 285.750 266.400 ;
        RECT 307.650 265.800 309.450 267.600 ;
        RECT 310.950 266.400 313.050 268.500 ;
        RECT 316.050 266.400 317.850 272.400 ;
        RECT 331.800 266.400 333.600 272.400 ;
        RECT 297.150 264.000 298.950 264.600 ;
        RECT 308.100 264.000 309.150 265.800 ;
        RECT 297.150 262.800 309.150 264.000 ;
        RECT 248.100 256.050 249.900 257.850 ;
        RECT 250.950 256.950 253.050 259.050 ;
        RECT 247.950 253.950 250.050 256.050 ;
        RECT 241.950 244.950 244.050 247.050 ;
        RECT 190.800 237.600 192.600 243.600 ;
        RECT 212.400 237.600 214.200 243.600 ;
        RECT 232.800 237.600 234.600 243.600 ;
        RECT 251.400 243.600 252.600 256.950 ;
        RECT 254.100 256.050 255.900 257.850 ;
        RECT 272.100 256.050 273.900 257.850 ;
        RECT 274.950 256.950 277.050 259.050 ;
        RECT 253.950 253.950 256.050 256.050 ;
        RECT 271.950 253.950 274.050 256.050 ;
        RECT 275.850 243.600 277.050 256.950 ;
        RECT 278.100 256.050 279.900 257.850 ;
        RECT 280.950 256.950 283.050 259.050 ;
        RECT 284.550 257.250 290.850 259.050 ;
        RECT 284.550 256.950 289.050 257.250 ;
        RECT 277.950 253.950 280.050 256.050 ;
        RECT 281.100 255.150 282.900 256.950 ;
        RECT 284.550 249.600 285.750 256.950 ;
        RECT 286.950 251.400 288.750 253.200 ;
        RECT 287.850 250.200 292.050 251.400 ;
        RECT 297.150 250.200 298.050 262.800 ;
        RECT 308.100 261.600 315.000 262.800 ;
        RECT 308.100 261.000 309.900 261.600 ;
        RECT 314.100 260.850 315.000 261.600 ;
        RECT 311.100 259.800 312.900 260.400 ;
        RECT 304.950 258.600 312.900 259.800 ;
        RECT 314.100 259.050 315.900 260.850 ;
        RECT 304.950 256.950 307.050 258.600 ;
        RECT 313.950 256.950 316.050 259.050 ;
        RECT 306.750 251.700 308.550 252.000 ;
        RECT 316.950 251.700 317.850 266.400 ;
        RECT 332.400 264.300 333.600 266.400 ;
        RECT 334.800 267.300 336.600 272.400 ;
        RECT 340.800 267.300 342.600 272.400 ;
        RECT 334.800 265.950 342.600 267.300 ;
        RECT 353.400 267.300 355.200 272.400 ;
        RECT 359.400 267.300 361.200 272.400 ;
        RECT 353.400 265.950 361.200 267.300 ;
        RECT 362.400 266.400 364.200 272.400 ;
        RECT 379.800 266.400 381.600 272.400 ;
        RECT 362.400 264.300 363.600 266.400 ;
        RECT 332.400 263.250 336.150 264.300 ;
        RECT 334.950 259.050 336.150 263.250 ;
        RECT 359.850 263.250 363.600 264.300 ;
        RECT 380.400 264.300 381.600 266.400 ;
        RECT 382.800 267.300 384.600 272.400 ;
        RECT 388.800 267.300 390.600 272.400 ;
        RECT 382.800 265.950 390.600 267.300 ;
        RECT 404.400 269.400 406.200 272.400 ;
        RECT 380.400 263.250 384.150 264.300 ;
        RECT 359.850 259.050 361.050 263.250 ;
        RECT 332.100 256.050 333.900 257.850 ;
        RECT 334.950 256.950 337.050 259.050 ;
        RECT 331.950 253.950 334.050 256.050 ;
        RECT 306.750 251.100 317.850 251.700 ;
        RECT 251.400 237.600 253.200 243.600 ;
        RECT 275.400 237.600 277.200 243.600 ;
        RECT 284.550 237.600 286.350 249.600 ;
        RECT 289.950 249.300 292.050 250.200 ;
        RECT 292.950 249.300 298.050 250.200 ;
        RECT 300.150 250.500 317.850 251.100 ;
        RECT 300.150 250.200 308.550 250.500 ;
        RECT 292.950 248.400 293.850 249.300 ;
        RECT 291.150 246.600 293.850 248.400 ;
        RECT 294.750 248.100 296.550 248.400 ;
        RECT 300.150 248.100 301.050 250.200 ;
        RECT 316.950 249.600 317.850 250.500 ;
        RECT 294.750 247.200 301.050 248.100 ;
        RECT 301.950 248.700 303.750 249.300 ;
        RECT 301.950 247.500 309.450 248.700 ;
        RECT 294.750 246.600 296.550 247.200 ;
        RECT 308.250 246.600 309.450 247.500 ;
        RECT 289.950 243.600 293.850 245.700 ;
        RECT 298.950 245.550 300.750 246.300 ;
        RECT 303.750 245.550 305.550 246.300 ;
        RECT 298.950 244.500 305.550 245.550 ;
        RECT 308.250 244.500 313.050 246.600 ;
        RECT 292.050 237.600 293.850 243.600 ;
        RECT 299.850 237.600 301.650 244.500 ;
        RECT 308.250 243.600 309.450 244.500 ;
        RECT 307.650 237.600 309.450 243.600 ;
        RECT 316.050 237.600 317.850 249.600 ;
        RECT 335.850 243.600 337.050 256.950 ;
        RECT 338.100 256.050 339.900 257.850 ;
        RECT 340.950 256.950 343.050 259.050 ;
        RECT 352.950 256.950 355.050 259.050 ;
        RECT 337.950 253.950 340.050 256.050 ;
        RECT 341.100 255.150 342.900 256.950 ;
        RECT 353.100 255.150 354.900 256.950 ;
        RECT 356.100 256.050 357.900 257.850 ;
        RECT 358.950 256.950 361.050 259.050 ;
        RECT 382.950 259.050 384.150 263.250 ;
        RECT 355.950 253.950 358.050 256.050 ;
        RECT 358.950 243.600 360.150 256.950 ;
        RECT 362.100 256.050 363.900 257.850 ;
        RECT 380.100 256.050 381.900 257.850 ;
        RECT 382.950 256.950 385.050 259.050 ;
        RECT 361.950 253.950 364.050 256.050 ;
        RECT 379.950 253.950 382.050 256.050 ;
        RECT 383.850 243.600 385.050 256.950 ;
        RECT 386.100 256.050 387.900 257.850 ;
        RECT 388.950 256.950 391.050 259.050 ;
        RECT 400.950 256.950 403.050 259.050 ;
        RECT 385.950 253.950 388.050 256.050 ;
        RECT 389.100 255.150 390.900 256.950 ;
        RECT 401.100 255.150 402.900 256.950 ;
        RECT 404.400 256.050 405.600 269.400 ;
        RECT 421.800 266.400 423.600 272.400 ;
        RECT 442.800 269.400 444.600 272.400 ;
        RECT 463.800 269.400 465.600 272.400 ;
        RECT 482.400 269.400 484.200 272.400 ;
        RECT 422.400 259.050 423.600 266.400 ;
        RECT 439.950 259.950 442.050 262.050 ;
        RECT 421.950 256.950 424.050 259.050 ;
        RECT 440.100 258.150 441.900 259.950 ;
        RECT 443.400 259.050 444.300 269.400 ;
        RECT 454.950 262.950 457.050 265.050 ;
        RECT 445.950 259.950 448.050 262.050 ;
        RECT 403.950 250.950 406.050 256.050 ;
        RECT 404.400 243.600 405.600 250.950 ;
        RECT 422.400 249.600 423.600 256.950 ;
        RECT 425.100 256.050 426.900 257.850 ;
        RECT 442.950 256.950 445.050 259.050 ;
        RECT 446.100 258.150 447.900 259.950 ;
        RECT 424.950 253.950 427.050 256.050 ;
        RECT 443.400 249.600 444.300 256.950 ;
        RECT 448.950 253.950 451.050 256.050 ;
        RECT 335.400 237.600 337.200 243.600 ;
        RECT 358.800 237.600 360.600 243.600 ;
        RECT 383.400 237.600 385.200 243.600 ;
        RECT 404.400 237.600 406.200 243.600 ;
        RECT 421.800 237.600 423.600 249.600 ;
        RECT 440.700 248.400 444.300 249.600 ;
        RECT 440.700 237.600 442.500 248.400 ;
        RECT 449.550 241.050 450.450 253.950 ;
        RECT 455.550 244.050 456.450 262.950 ;
        RECT 460.950 259.950 463.050 262.050 ;
        RECT 461.100 258.150 462.900 259.950 ;
        RECT 464.400 259.050 465.300 269.400 ;
        RECT 466.950 259.950 469.050 262.050 ;
        RECT 463.950 256.950 466.050 259.050 ;
        RECT 467.100 258.150 468.900 259.950 ;
        RECT 478.950 256.950 481.050 259.050 ;
        RECT 464.400 249.600 465.300 256.950 ;
        RECT 479.100 255.150 480.900 256.950 ;
        RECT 482.400 256.050 483.600 269.400 ;
        RECT 497.400 267.300 499.200 272.400 ;
        RECT 503.400 267.300 505.200 272.400 ;
        RECT 497.400 265.950 505.200 267.300 ;
        RECT 506.400 266.400 508.200 272.400 ;
        RECT 514.950 268.950 517.050 271.050 ;
        RECT 521.400 269.400 523.200 272.400 ;
        RECT 506.400 264.300 507.600 266.400 ;
        RECT 503.850 263.250 507.600 264.300 ;
        RECT 503.850 259.050 505.050 263.250 ;
        RECT 496.950 256.950 499.050 259.050 ;
        RECT 481.950 250.950 484.050 256.050 ;
        RECT 497.100 255.150 498.900 256.950 ;
        RECT 500.100 256.050 501.900 257.850 ;
        RECT 502.950 256.950 505.050 259.050 ;
        RECT 499.950 253.950 502.050 256.050 ;
        RECT 461.700 248.400 465.300 249.600 ;
        RECT 455.100 241.950 457.200 244.050 ;
        RECT 448.950 238.950 451.050 241.050 ;
        RECT 461.700 237.600 463.500 248.400 ;
        RECT 482.400 243.600 483.600 250.950 ;
        RECT 502.950 243.600 504.150 256.950 ;
        RECT 506.100 256.050 507.900 257.850 ;
        RECT 511.950 256.950 514.050 259.050 ;
        RECT 505.950 253.950 508.050 256.050 ;
        RECT 512.550 250.050 513.450 256.950 ;
        RECT 511.950 247.950 514.050 250.050 ;
        RECT 515.550 244.050 516.450 268.950 ;
        RECT 521.400 265.500 522.600 269.400 ;
        RECT 527.700 266.400 529.500 272.400 ;
        RECT 521.400 264.600 527.400 265.500 ;
        RECT 525.150 263.700 527.400 264.600 ;
        RECT 520.950 256.950 523.050 259.050 ;
        RECT 521.100 255.150 522.900 256.950 ;
        RECT 525.150 252.300 526.050 263.700 ;
        RECT 528.300 259.050 529.500 266.400 ;
        RECT 526.950 256.950 529.500 259.050 ;
        RECT 525.150 251.400 527.400 252.300 ;
        RECT 521.400 250.500 527.400 251.400 ;
        RECT 482.400 237.600 484.200 243.600 ;
        RECT 502.800 237.600 504.600 243.600 ;
        RECT 514.950 241.950 517.050 244.050 ;
        RECT 521.400 243.600 522.600 250.500 ;
        RECT 528.300 249.600 529.500 256.950 ;
        RECT 521.400 237.600 523.200 243.600 ;
        RECT 527.700 237.600 529.500 249.600 ;
        RECT 534.150 266.400 535.950 272.400 ;
        RECT 541.950 270.300 543.750 272.400 ;
        RECT 540.000 269.400 543.750 270.300 ;
        RECT 549.750 269.400 551.550 272.400 ;
        RECT 557.550 269.400 559.350 272.400 ;
        RECT 540.000 268.500 541.050 269.400 ;
        RECT 549.750 268.500 550.800 269.400 ;
        RECT 538.950 266.400 541.050 268.500 ;
        RECT 534.150 251.700 535.050 266.400 ;
        RECT 542.550 265.800 544.350 267.600 ;
        RECT 545.850 267.450 550.800 268.500 ;
        RECT 558.300 268.500 559.350 269.400 ;
        RECT 545.850 266.700 547.650 267.450 ;
        RECT 558.300 267.300 562.050 268.500 ;
        RECT 559.950 266.400 562.050 267.300 ;
        RECT 565.650 266.400 567.450 272.400 ;
        RECT 542.850 264.000 543.900 265.800 ;
        RECT 553.050 264.000 554.850 264.600 ;
        RECT 542.850 262.800 554.850 264.000 ;
        RECT 537.000 261.600 543.900 262.800 ;
        RECT 537.000 260.850 537.900 261.600 ;
        RECT 542.100 261.000 543.900 261.600 ;
        RECT 536.100 259.050 537.900 260.850 ;
        RECT 539.100 259.800 540.900 260.400 ;
        RECT 535.950 256.950 538.050 259.050 ;
        RECT 539.100 258.600 547.050 259.800 ;
        RECT 544.950 256.950 547.050 258.600 ;
        RECT 543.450 251.700 545.250 252.000 ;
        RECT 534.150 251.100 545.250 251.700 ;
        RECT 534.150 250.500 551.850 251.100 ;
        RECT 534.150 249.600 535.050 250.500 ;
        RECT 543.450 250.200 551.850 250.500 ;
        RECT 534.150 237.600 535.950 249.600 ;
        RECT 548.250 248.700 550.050 249.300 ;
        RECT 542.550 247.500 550.050 248.700 ;
        RECT 550.950 248.100 551.850 250.200 ;
        RECT 553.950 250.200 554.850 262.800 ;
        RECT 566.250 259.050 567.450 266.400 ;
        RECT 578.400 267.300 580.200 272.400 ;
        RECT 584.400 267.300 586.200 272.400 ;
        RECT 578.400 265.950 586.200 267.300 ;
        RECT 587.400 266.400 589.200 272.400 ;
        RECT 587.400 264.300 588.600 266.400 ;
        RECT 607.800 265.200 609.600 272.400 ;
        RECT 626.400 269.400 628.200 272.400 ;
        RECT 584.850 263.250 588.600 264.300 ;
        RECT 605.400 264.300 609.600 265.200 ;
        RECT 584.850 259.050 586.050 263.250 ;
        RECT 605.400 259.050 606.600 264.300 ;
        RECT 622.950 259.950 625.050 262.050 ;
        RECT 561.150 257.250 567.450 259.050 ;
        RECT 562.950 256.950 567.450 257.250 ;
        RECT 577.950 256.950 580.050 259.050 ;
        RECT 563.250 251.400 565.050 253.200 ;
        RECT 559.950 250.200 564.150 251.400 ;
        RECT 553.950 249.300 559.050 250.200 ;
        RECT 559.950 249.300 562.050 250.200 ;
        RECT 566.250 249.600 567.450 256.950 ;
        RECT 578.100 255.150 579.900 256.950 ;
        RECT 581.100 256.050 582.900 257.850 ;
        RECT 583.950 256.950 586.050 259.050 ;
        RECT 580.950 253.950 583.050 256.050 ;
        RECT 558.150 248.400 559.050 249.300 ;
        RECT 555.450 248.100 557.250 248.400 ;
        RECT 542.550 246.600 543.750 247.500 ;
        RECT 550.950 247.200 557.250 248.100 ;
        RECT 555.450 246.600 557.250 247.200 ;
        RECT 558.150 246.600 560.850 248.400 ;
        RECT 538.950 244.500 543.750 246.600 ;
        RECT 546.450 245.550 548.250 246.300 ;
        RECT 551.250 245.550 553.050 246.300 ;
        RECT 546.450 244.500 553.050 245.550 ;
        RECT 542.550 243.600 543.750 244.500 ;
        RECT 542.550 237.600 544.350 243.600 ;
        RECT 550.350 237.600 552.150 244.500 ;
        RECT 558.150 243.600 562.050 245.700 ;
        RECT 558.150 237.600 559.950 243.600 ;
        RECT 565.650 237.600 567.450 249.600 ;
        RECT 583.950 243.600 585.150 256.950 ;
        RECT 587.100 256.050 588.900 257.850 ;
        RECT 602.100 256.050 603.900 257.850 ;
        RECT 604.950 256.950 607.050 259.050 ;
        RECT 623.100 258.150 624.900 259.950 ;
        RECT 626.700 259.050 627.600 269.400 ;
        RECT 647.400 265.500 649.200 272.400 ;
        RECT 653.400 265.500 655.200 272.400 ;
        RECT 659.400 265.500 661.200 272.400 ;
        RECT 665.400 265.500 667.200 272.400 ;
        RECT 686.400 269.400 688.200 272.400 ;
        RECT 647.400 264.300 651.300 265.500 ;
        RECT 653.400 264.300 657.300 265.500 ;
        RECT 659.400 264.300 663.300 265.500 ;
        RECT 665.400 264.300 668.100 265.500 ;
        RECT 650.100 263.400 651.300 264.300 ;
        RECT 656.100 263.400 657.300 264.300 ;
        RECT 662.100 263.400 663.300 264.300 ;
        RECT 650.100 262.200 654.300 263.400 ;
        RECT 628.950 259.950 631.050 262.050 ;
        RECT 586.950 253.950 589.050 256.050 ;
        RECT 601.950 253.950 604.050 256.050 ;
        RECT 605.400 243.600 606.600 256.950 ;
        RECT 608.100 256.050 609.900 257.850 ;
        RECT 625.950 256.950 628.050 259.050 ;
        RECT 629.100 258.150 630.900 259.950 ;
        RECT 647.100 259.050 648.900 260.850 ;
        RECT 646.950 256.950 649.050 259.050 ;
        RECT 607.950 253.950 610.050 256.050 ;
        RECT 626.700 249.600 627.600 256.950 ;
        RECT 650.100 251.700 651.300 262.200 ;
        RECT 652.500 261.600 654.300 262.200 ;
        RECT 656.100 262.200 660.300 263.400 ;
        RECT 656.100 251.700 657.300 262.200 ;
        RECT 658.500 261.600 660.300 262.200 ;
        RECT 662.100 262.200 666.300 263.400 ;
        RECT 662.100 251.700 663.300 262.200 ;
        RECT 664.500 261.600 666.300 262.200 ;
        RECT 667.200 259.050 668.100 264.300 ;
        RECT 667.200 256.950 670.050 259.050 ;
        RECT 682.950 256.950 685.050 259.050 ;
        RECT 667.200 251.700 668.100 256.950 ;
        RECT 679.950 253.950 682.050 256.050 ;
        RECT 683.100 255.150 684.900 256.950 ;
        RECT 686.400 256.050 687.600 269.400 ;
        RECT 701.400 267.300 703.200 272.400 ;
        RECT 707.400 267.300 709.200 272.400 ;
        RECT 701.400 265.950 709.200 267.300 ;
        RECT 710.400 266.400 712.200 272.400 ;
        RECT 715.950 268.950 718.050 271.050 ;
        RECT 710.400 264.300 711.600 266.400 ;
        RECT 707.850 263.250 711.600 264.300 ;
        RECT 707.850 259.050 709.050 263.250 ;
        RECT 700.950 256.950 703.050 259.050 ;
        RECT 647.400 250.500 651.300 251.700 ;
        RECT 653.400 250.500 657.300 251.700 ;
        RECT 659.400 250.500 663.300 251.700 ;
        RECT 665.400 250.500 668.100 251.700 ;
        RECT 626.700 248.400 630.300 249.600 ;
        RECT 583.800 237.600 585.600 243.600 ;
        RECT 605.400 237.600 607.200 243.600 ;
        RECT 628.500 237.600 630.300 248.400 ;
        RECT 647.400 237.600 649.200 250.500 ;
        RECT 653.400 237.600 655.200 250.500 ;
        RECT 659.400 237.600 661.200 250.500 ;
        RECT 665.400 237.600 667.200 250.500 ;
        RECT 680.550 241.050 681.450 253.950 ;
        RECT 685.950 250.950 688.050 256.050 ;
        RECT 701.100 255.150 702.900 256.950 ;
        RECT 704.100 256.050 705.900 257.850 ;
        RECT 706.950 256.950 709.050 259.050 ;
        RECT 703.950 253.950 706.050 256.050 ;
        RECT 686.400 243.600 687.600 250.950 ;
        RECT 706.950 243.600 708.150 256.950 ;
        RECT 710.100 256.050 711.900 257.850 ;
        RECT 709.950 253.950 712.050 256.050 ;
        RECT 716.550 247.050 717.450 268.950 ;
        RECT 728.400 265.200 730.200 272.400 ;
        RECT 749.400 265.200 751.200 272.400 ;
        RECT 770.400 265.200 772.200 272.400 ;
        RECT 788.400 267.300 790.200 272.400 ;
        RECT 794.400 267.300 796.200 272.400 ;
        RECT 788.400 265.950 796.200 267.300 ;
        RECT 797.400 266.400 799.200 272.400 ;
        RECT 728.400 264.300 732.600 265.200 ;
        RECT 749.400 264.300 753.600 265.200 ;
        RECT 770.400 264.300 774.600 265.200 ;
        RECT 797.400 264.300 798.600 266.400 ;
        RECT 802.950 265.950 805.050 268.050 ;
        RECT 814.800 266.400 816.600 272.400 ;
        RECT 731.400 259.050 732.600 264.300 ;
        RECT 752.400 259.050 753.600 264.300 ;
        RECT 773.400 259.050 774.600 264.300 ;
        RECT 794.850 263.250 798.600 264.300 ;
        RECT 794.850 259.050 796.050 263.250 ;
        RECT 728.100 256.050 729.900 257.850 ;
        RECT 730.950 256.950 733.050 259.050 ;
        RECT 727.950 253.950 730.050 256.050 ;
        RECT 715.950 244.950 718.050 247.050 ;
        RECT 679.950 238.950 682.050 241.050 ;
        RECT 686.400 237.600 688.200 243.600 ;
        RECT 706.800 237.600 708.600 243.600 ;
        RECT 712.950 243.450 715.050 244.050 ;
        RECT 718.950 243.450 721.050 244.050 ;
        RECT 731.400 243.600 732.600 256.950 ;
        RECT 734.100 256.050 735.900 257.850 ;
        RECT 749.100 256.050 750.900 257.850 ;
        RECT 751.950 256.950 754.050 259.050 ;
        RECT 733.950 253.950 736.050 256.050 ;
        RECT 748.950 253.950 751.050 256.050 ;
        RECT 752.400 243.600 753.600 256.950 ;
        RECT 755.100 256.050 756.900 257.850 ;
        RECT 770.100 256.050 771.900 257.850 ;
        RECT 772.950 256.950 775.050 259.050 ;
        RECT 754.950 253.950 757.050 256.050 ;
        RECT 769.950 253.950 772.050 256.050 ;
        RECT 773.400 243.600 774.600 256.950 ;
        RECT 776.100 256.050 777.900 257.850 ;
        RECT 787.950 256.950 790.050 259.050 ;
        RECT 775.950 253.950 778.050 256.050 ;
        RECT 788.100 255.150 789.900 256.950 ;
        RECT 791.100 256.050 792.900 257.850 ;
        RECT 793.950 256.950 796.050 259.050 ;
        RECT 790.950 253.950 793.050 256.050 ;
        RECT 793.950 243.600 795.150 256.950 ;
        RECT 797.100 256.050 798.900 257.850 ;
        RECT 796.950 253.950 799.050 256.050 ;
        RECT 803.550 247.050 804.450 265.950 ;
        RECT 815.400 264.300 816.600 266.400 ;
        RECT 817.800 267.300 819.600 272.400 ;
        RECT 823.800 267.300 825.600 272.400 ;
        RECT 838.800 269.400 840.600 272.400 ;
        RECT 857.400 269.400 859.200 272.400 ;
        RECT 878.400 269.400 880.200 272.400 ;
        RECT 896.400 269.400 898.200 272.400 ;
        RECT 817.800 265.950 825.600 267.300 ;
        RECT 815.400 263.250 819.150 264.300 ;
        RECT 817.950 259.050 819.150 263.250 ;
        RECT 815.100 256.050 816.900 257.850 ;
        RECT 817.950 256.950 820.050 259.050 ;
        RECT 814.950 253.950 817.050 256.050 ;
        RECT 802.950 244.950 805.050 247.050 ;
        RECT 818.850 243.600 820.050 256.950 ;
        RECT 821.100 256.050 822.900 257.850 ;
        RECT 823.950 256.950 826.050 259.050 ;
        RECT 820.950 253.950 823.050 256.050 ;
        RECT 824.100 255.150 825.900 256.950 ;
        RECT 839.400 256.050 840.600 269.400 ;
        RECT 847.950 262.950 850.050 265.050 ;
        RECT 841.950 256.950 844.050 259.050 ;
        RECT 838.950 250.950 841.050 256.050 ;
        RECT 842.100 255.150 843.900 256.950 ;
        RECT 839.400 243.600 840.600 250.950 ;
        RECT 848.550 247.050 849.450 262.950 ;
        RECT 853.950 259.950 856.050 262.050 ;
        RECT 854.100 258.150 855.900 259.950 ;
        RECT 857.700 259.050 858.600 269.400 ;
        RECT 859.950 259.950 862.050 262.050 ;
        RECT 874.950 259.950 877.050 262.050 ;
        RECT 856.950 256.950 859.050 259.050 ;
        RECT 860.100 258.150 861.900 259.950 ;
        RECT 875.100 258.150 876.900 259.950 ;
        RECT 878.700 259.050 879.600 269.400 ;
        RECT 896.400 265.500 897.600 269.400 ;
        RECT 902.700 266.400 904.500 272.400 ;
        RECT 896.400 264.600 902.400 265.500 ;
        RECT 900.150 263.700 902.400 264.600 ;
        RECT 880.950 259.950 883.050 262.050 ;
        RECT 877.950 256.950 880.050 259.050 ;
        RECT 881.100 258.150 882.900 259.950 ;
        RECT 895.950 256.950 898.050 259.050 ;
        RECT 857.700 249.600 858.600 256.950 ;
        RECT 878.700 249.600 879.600 256.950 ;
        RECT 896.100 255.150 897.900 256.950 ;
        RECT 900.150 252.300 901.050 263.700 ;
        RECT 903.300 259.050 904.500 266.400 ;
        RECT 901.950 256.950 904.500 259.050 ;
        RECT 900.150 251.400 902.400 252.300 ;
        RECT 896.400 250.500 902.400 251.400 ;
        RECT 857.700 248.400 861.300 249.600 ;
        RECT 878.700 248.400 882.300 249.600 ;
        RECT 847.950 244.950 850.050 247.050 ;
        RECT 712.950 242.550 721.050 243.450 ;
        RECT 712.950 241.950 715.050 242.550 ;
        RECT 718.950 241.950 721.050 242.550 ;
        RECT 730.800 237.600 732.600 243.600 ;
        RECT 751.800 237.600 753.600 243.600 ;
        RECT 772.800 237.600 774.600 243.600 ;
        RECT 793.800 237.600 795.600 243.600 ;
        RECT 818.400 237.600 820.200 243.600 ;
        RECT 838.800 237.600 840.600 243.600 ;
        RECT 859.500 237.600 861.300 248.400 ;
        RECT 880.500 237.600 882.300 248.400 ;
        RECT 896.400 243.600 897.600 250.500 ;
        RECT 903.300 249.600 904.500 256.950 ;
        RECT 896.400 237.600 898.200 243.600 ;
        RECT 902.700 237.600 904.500 249.600 ;
        RECT 16.800 227.400 18.600 233.400 ;
        RECT 38.400 227.400 40.200 233.400 ;
        RECT 13.950 214.950 16.050 217.050 ;
        RECT 14.100 213.150 15.900 214.950 ;
        RECT 17.400 214.050 18.600 227.400 ;
        RECT 19.950 214.950 22.050 217.050 ;
        RECT 34.950 214.950 37.050 217.050 ;
        RECT 16.950 211.950 19.050 214.050 ;
        RECT 20.100 213.150 21.900 214.950 ;
        RECT 35.100 213.150 36.900 214.950 ;
        RECT 38.850 214.050 40.050 227.400 ;
        RECT 59.700 222.600 61.500 233.400 ;
        RECT 70.950 223.950 73.050 226.050 ;
        RECT 59.700 221.400 63.300 222.600 ;
        RECT 40.950 214.950 43.050 217.050 ;
        RECT 37.950 211.950 40.050 214.050 ;
        RECT 41.100 213.150 42.900 214.950 ;
        RECT 44.100 214.050 45.900 215.850 ;
        RECT 62.400 214.050 63.300 221.400 ;
        RECT 71.550 217.050 72.450 223.950 ;
        RECT 80.700 222.600 82.500 233.400 ;
        RECT 80.700 221.400 84.300 222.600 ;
        RECT 70.950 214.950 73.050 217.050 ;
        RECT 83.400 214.050 84.300 221.400 ;
        RECT 89.550 221.400 91.350 233.400 ;
        RECT 97.050 227.400 98.850 233.400 ;
        RECT 94.950 225.300 98.850 227.400 ;
        RECT 104.850 226.500 106.650 233.400 ;
        RECT 112.650 227.400 114.450 233.400 ;
        RECT 113.250 226.500 114.450 227.400 ;
        RECT 103.950 225.450 110.550 226.500 ;
        RECT 103.950 224.700 105.750 225.450 ;
        RECT 108.750 224.700 110.550 225.450 ;
        RECT 113.250 224.400 118.050 226.500 ;
        RECT 96.150 222.600 98.850 224.400 ;
        RECT 99.750 223.800 101.550 224.400 ;
        RECT 99.750 222.900 106.050 223.800 ;
        RECT 113.250 223.500 114.450 224.400 ;
        RECT 99.750 222.600 101.550 222.900 ;
        RECT 97.950 221.700 98.850 222.600 ;
        RECT 89.550 214.050 90.750 221.400 ;
        RECT 94.950 220.800 97.050 221.700 ;
        RECT 97.950 220.800 103.050 221.700 ;
        RECT 92.850 219.600 97.050 220.800 ;
        RECT 91.950 217.800 93.750 219.600 ;
        RECT 43.950 211.950 46.050 214.050 ;
        RECT 17.400 206.700 18.600 211.950 ;
        RECT 37.950 207.750 39.150 211.950 ;
        RECT 59.100 211.050 60.900 212.850 ;
        RECT 61.950 211.950 64.050 214.050 ;
        RECT 58.950 208.950 61.050 211.050 ;
        RECT 14.400 205.800 18.600 206.700 ;
        RECT 35.400 206.700 39.150 207.750 ;
        RECT 14.400 198.600 16.200 205.800 ;
        RECT 35.400 204.600 36.600 206.700 ;
        RECT 34.800 198.600 36.600 204.600 ;
        RECT 37.800 203.700 45.600 205.050 ;
        RECT 37.800 198.600 39.600 203.700 ;
        RECT 43.800 198.600 45.600 203.700 ;
        RECT 62.400 201.600 63.300 211.950 ;
        RECT 65.100 211.050 66.900 212.850 ;
        RECT 80.100 211.050 81.900 212.850 ;
        RECT 82.950 211.950 85.050 214.050 ;
        RECT 89.550 213.750 94.050 214.050 ;
        RECT 64.950 208.950 67.050 211.050 ;
        RECT 79.950 208.950 82.050 211.050 ;
        RECT 83.400 201.600 84.300 211.950 ;
        RECT 86.100 211.050 87.900 212.850 ;
        RECT 89.550 211.950 95.850 213.750 ;
        RECT 85.950 208.950 88.050 211.050 ;
        RECT 89.550 204.600 90.750 211.950 ;
        RECT 102.150 208.200 103.050 220.800 ;
        RECT 105.150 220.800 106.050 222.900 ;
        RECT 106.950 222.300 114.450 223.500 ;
        RECT 106.950 221.700 108.750 222.300 ;
        RECT 121.050 221.400 122.850 233.400 ;
        RECT 139.800 227.400 141.600 233.400 ;
        RECT 161.400 227.400 163.200 233.400 ;
        RECT 105.150 220.500 113.550 220.800 ;
        RECT 121.950 220.500 122.850 221.400 ;
        RECT 105.150 219.900 122.850 220.500 ;
        RECT 111.750 219.300 122.850 219.900 ;
        RECT 111.750 219.000 113.550 219.300 ;
        RECT 109.950 212.400 112.050 214.050 ;
        RECT 109.950 211.200 117.900 212.400 ;
        RECT 118.950 211.950 121.050 214.050 ;
        RECT 116.100 210.600 117.900 211.200 ;
        RECT 119.100 210.150 120.900 211.950 ;
        RECT 113.100 209.400 114.900 210.000 ;
        RECT 119.100 209.400 120.000 210.150 ;
        RECT 113.100 208.200 120.000 209.400 ;
        RECT 102.150 207.000 114.150 208.200 ;
        RECT 102.150 206.400 103.950 207.000 ;
        RECT 113.100 205.200 114.150 207.000 ;
        RECT 61.800 198.600 63.600 201.600 ;
        RECT 82.800 198.600 84.600 201.600 ;
        RECT 89.550 198.600 91.350 204.600 ;
        RECT 94.950 203.700 97.050 204.600 ;
        RECT 94.950 202.500 98.700 203.700 ;
        RECT 109.350 203.550 111.150 204.300 ;
        RECT 97.650 201.600 98.700 202.500 ;
        RECT 106.200 202.500 111.150 203.550 ;
        RECT 112.650 203.400 114.450 205.200 ;
        RECT 121.950 204.600 122.850 219.300 ;
        RECT 134.100 214.050 135.900 215.850 ;
        RECT 136.950 214.950 139.050 217.050 ;
        RECT 133.950 211.950 136.050 214.050 ;
        RECT 137.100 213.150 138.900 214.950 ;
        RECT 139.950 214.050 141.150 227.400 ;
        RECT 142.950 214.950 145.050 217.050 ;
        RECT 157.950 214.950 160.050 217.050 ;
        RECT 139.950 211.950 142.050 214.050 ;
        RECT 143.100 213.150 144.900 214.950 ;
        RECT 158.100 213.150 159.900 214.950 ;
        RECT 161.400 214.050 162.600 227.400 ;
        RECT 170.550 221.400 172.350 233.400 ;
        RECT 178.050 227.400 179.850 233.400 ;
        RECT 175.950 225.300 179.850 227.400 ;
        RECT 185.850 226.500 187.650 233.400 ;
        RECT 193.650 227.400 195.450 233.400 ;
        RECT 194.250 226.500 195.450 227.400 ;
        RECT 184.950 225.450 191.550 226.500 ;
        RECT 184.950 224.700 186.750 225.450 ;
        RECT 189.750 224.700 191.550 225.450 ;
        RECT 194.250 224.400 199.050 226.500 ;
        RECT 177.150 222.600 179.850 224.400 ;
        RECT 180.750 223.800 182.550 224.400 ;
        RECT 180.750 222.900 187.050 223.800 ;
        RECT 194.250 223.500 195.450 224.400 ;
        RECT 180.750 222.600 182.550 222.900 ;
        RECT 178.950 221.700 179.850 222.600 ;
        RECT 163.950 214.950 166.050 217.050 ;
        RECT 160.950 211.950 163.050 214.050 ;
        RECT 164.100 213.150 165.900 214.950 ;
        RECT 170.550 214.050 171.750 221.400 ;
        RECT 175.950 220.800 178.050 221.700 ;
        RECT 178.950 220.800 184.050 221.700 ;
        RECT 173.850 219.600 178.050 220.800 ;
        RECT 172.950 217.800 174.750 219.600 ;
        RECT 170.550 213.750 175.050 214.050 ;
        RECT 170.550 211.950 176.850 213.750 ;
        RECT 140.850 207.750 142.050 211.950 ;
        RECT 140.850 206.700 144.600 207.750 ;
        RECT 115.950 202.500 118.050 204.600 ;
        RECT 106.200 201.600 107.250 202.500 ;
        RECT 115.950 201.600 117.000 202.500 ;
        RECT 97.650 198.600 99.450 201.600 ;
        RECT 105.450 198.600 107.250 201.600 ;
        RECT 113.250 200.700 117.000 201.600 ;
        RECT 113.250 198.600 115.050 200.700 ;
        RECT 121.050 198.600 122.850 204.600 ;
        RECT 134.400 203.700 142.200 205.050 ;
        RECT 134.400 198.600 136.200 203.700 ;
        RECT 140.400 198.600 142.200 203.700 ;
        RECT 143.400 204.600 144.600 206.700 ;
        RECT 161.400 206.700 162.600 211.950 ;
        RECT 161.400 205.800 165.600 206.700 ;
        RECT 143.400 198.600 145.200 204.600 ;
        RECT 163.800 198.600 165.600 205.800 ;
        RECT 170.550 204.600 171.750 211.950 ;
        RECT 183.150 208.200 184.050 220.800 ;
        RECT 186.150 220.800 187.050 222.900 ;
        RECT 187.950 222.300 195.450 223.500 ;
        RECT 187.950 221.700 189.750 222.300 ;
        RECT 202.050 221.400 203.850 233.400 ;
        RECT 221.400 227.400 223.200 233.400 ;
        RECT 245.400 227.400 247.200 233.400 ;
        RECT 268.800 227.400 270.600 233.400 ;
        RECT 186.150 220.500 194.550 220.800 ;
        RECT 202.950 220.500 203.850 221.400 ;
        RECT 186.150 219.900 203.850 220.500 ;
        RECT 192.750 219.300 203.850 219.900 ;
        RECT 192.750 219.000 194.550 219.300 ;
        RECT 190.950 212.400 193.050 214.050 ;
        RECT 190.950 211.200 198.900 212.400 ;
        RECT 199.950 211.950 202.050 214.050 ;
        RECT 197.100 210.600 198.900 211.200 ;
        RECT 200.100 210.150 201.900 211.950 ;
        RECT 194.100 209.400 195.900 210.000 ;
        RECT 200.100 209.400 201.000 210.150 ;
        RECT 194.100 208.200 201.000 209.400 ;
        RECT 183.150 207.000 195.150 208.200 ;
        RECT 183.150 206.400 184.950 207.000 ;
        RECT 194.100 205.200 195.150 207.000 ;
        RECT 170.550 198.600 172.350 204.600 ;
        RECT 175.950 203.700 178.050 204.600 ;
        RECT 175.950 202.500 179.700 203.700 ;
        RECT 190.350 203.550 192.150 204.300 ;
        RECT 178.650 201.600 179.700 202.500 ;
        RECT 187.200 202.500 192.150 203.550 ;
        RECT 193.650 203.400 195.450 205.200 ;
        RECT 202.950 204.600 203.850 219.300 ;
        RECT 217.950 214.950 220.050 217.050 ;
        RECT 218.100 213.150 219.900 214.950 ;
        RECT 221.850 214.050 223.050 227.400 ;
        RECT 223.950 214.950 226.050 217.050 ;
        RECT 220.950 211.950 223.050 214.050 ;
        RECT 224.100 213.150 225.900 214.950 ;
        RECT 227.100 214.050 228.900 215.850 ;
        RECT 241.950 214.950 244.050 217.050 ;
        RECT 226.950 211.950 229.050 214.050 ;
        RECT 242.100 213.150 243.900 214.950 ;
        RECT 245.850 214.050 247.050 227.400 ;
        RECT 247.950 214.950 250.050 217.050 ;
        RECT 244.950 211.950 247.050 214.050 ;
        RECT 248.100 213.150 249.900 214.950 ;
        RECT 251.100 214.050 252.900 215.850 ;
        RECT 263.100 214.050 264.900 215.850 ;
        RECT 265.950 214.950 268.050 217.050 ;
        RECT 250.950 211.950 253.050 214.050 ;
        RECT 262.950 211.950 265.050 214.050 ;
        RECT 266.100 213.150 267.900 214.950 ;
        RECT 268.950 214.050 270.150 227.400 ;
        RECT 290.700 222.600 292.500 233.400 ;
        RECT 314.400 227.400 316.200 233.400 ;
        RECT 334.800 227.400 336.600 233.400 ;
        RECT 290.700 221.400 294.300 222.600 ;
        RECT 271.950 214.950 274.050 217.050 ;
        RECT 268.950 211.950 271.050 214.050 ;
        RECT 272.100 213.150 273.900 214.950 ;
        RECT 293.400 214.050 294.300 221.400 ;
        RECT 310.950 214.950 313.050 217.050 ;
        RECT 220.950 207.750 222.150 211.950 ;
        RECT 244.950 207.750 246.150 211.950 ;
        RECT 218.400 206.700 222.150 207.750 ;
        RECT 242.400 206.700 246.150 207.750 ;
        RECT 269.850 207.750 271.050 211.950 ;
        RECT 290.100 211.050 291.900 212.850 ;
        RECT 292.950 211.950 295.050 214.050 ;
        RECT 311.100 213.150 312.900 214.950 ;
        RECT 314.850 214.050 316.050 227.400 ;
        RECT 335.400 220.050 336.600 227.400 ;
        RECT 350.400 227.400 352.200 233.400 ;
        RECT 316.950 214.950 319.050 217.050 ;
        RECT 289.950 208.950 292.050 211.050 ;
        RECT 269.850 206.700 273.600 207.750 ;
        RECT 218.400 204.600 219.600 206.700 ;
        RECT 196.950 202.500 199.050 204.600 ;
        RECT 187.200 201.600 188.250 202.500 ;
        RECT 196.950 201.600 198.000 202.500 ;
        RECT 178.650 198.600 180.450 201.600 ;
        RECT 186.450 198.600 188.250 201.600 ;
        RECT 194.250 200.700 198.000 201.600 ;
        RECT 194.250 198.600 196.050 200.700 ;
        RECT 202.050 198.600 203.850 204.600 ;
        RECT 217.800 198.600 219.600 204.600 ;
        RECT 220.800 203.700 228.600 205.050 ;
        RECT 242.400 204.600 243.600 206.700 ;
        RECT 220.800 198.600 222.600 203.700 ;
        RECT 226.800 198.600 228.600 203.700 ;
        RECT 241.800 198.600 243.600 204.600 ;
        RECT 244.800 203.700 252.600 205.050 ;
        RECT 244.800 198.600 246.600 203.700 ;
        RECT 250.800 198.600 252.600 203.700 ;
        RECT 263.400 203.700 271.200 205.050 ;
        RECT 263.400 198.600 265.200 203.700 ;
        RECT 269.400 198.600 271.200 203.700 ;
        RECT 272.400 204.600 273.600 206.700 ;
        RECT 272.400 198.600 274.200 204.600 ;
        RECT 293.400 201.600 294.300 211.950 ;
        RECT 296.100 211.050 297.900 212.850 ;
        RECT 313.950 211.950 316.050 214.050 ;
        RECT 317.100 213.150 318.900 214.950 ;
        RECT 320.100 214.050 321.900 215.850 ;
        RECT 334.950 214.950 337.050 220.050 ;
        RECT 319.950 211.950 322.050 214.050 ;
        RECT 295.950 208.950 298.050 211.050 ;
        RECT 313.950 207.750 315.150 211.950 ;
        RECT 311.400 206.700 315.150 207.750 ;
        RECT 311.400 204.600 312.600 206.700 ;
        RECT 292.800 198.600 294.600 201.600 ;
        RECT 310.800 198.600 312.600 204.600 ;
        RECT 313.800 203.700 321.600 205.050 ;
        RECT 313.800 198.600 315.600 203.700 ;
        RECT 319.800 198.600 321.600 203.700 ;
        RECT 335.400 201.600 336.600 214.950 ;
        RECT 338.100 214.050 339.900 215.850 ;
        RECT 346.950 214.950 349.050 217.050 ;
        RECT 337.950 211.950 340.050 214.050 ;
        RECT 347.100 213.150 348.900 214.950 ;
        RECT 350.400 214.050 351.600 227.400 ;
        RECT 359.550 221.400 361.350 233.400 ;
        RECT 367.050 227.400 368.850 233.400 ;
        RECT 364.950 225.300 368.850 227.400 ;
        RECT 374.850 226.500 376.650 233.400 ;
        RECT 382.650 227.400 384.450 233.400 ;
        RECT 383.250 226.500 384.450 227.400 ;
        RECT 373.950 225.450 380.550 226.500 ;
        RECT 373.950 224.700 375.750 225.450 ;
        RECT 378.750 224.700 380.550 225.450 ;
        RECT 383.250 224.400 388.050 226.500 ;
        RECT 366.150 222.600 368.850 224.400 ;
        RECT 369.750 223.800 371.550 224.400 ;
        RECT 369.750 222.900 376.050 223.800 ;
        RECT 383.250 223.500 384.450 224.400 ;
        RECT 369.750 222.600 371.550 222.900 ;
        RECT 367.950 221.700 368.850 222.600 ;
        RECT 352.950 214.950 355.050 217.050 ;
        RECT 349.950 211.950 352.050 214.050 ;
        RECT 353.100 213.150 354.900 214.950 ;
        RECT 359.550 214.050 360.750 221.400 ;
        RECT 364.950 220.800 367.050 221.700 ;
        RECT 367.950 220.800 373.050 221.700 ;
        RECT 362.850 219.600 367.050 220.800 ;
        RECT 361.950 217.800 363.750 219.600 ;
        RECT 359.550 213.750 364.050 214.050 ;
        RECT 359.550 211.950 365.850 213.750 ;
        RECT 350.400 206.700 351.600 211.950 ;
        RECT 350.400 205.800 354.600 206.700 ;
        RECT 334.800 198.600 336.600 201.600 ;
        RECT 352.800 198.600 354.600 205.800 ;
        RECT 359.550 204.600 360.750 211.950 ;
        RECT 372.150 208.200 373.050 220.800 ;
        RECT 375.150 220.800 376.050 222.900 ;
        RECT 376.950 222.300 384.450 223.500 ;
        RECT 376.950 221.700 378.750 222.300 ;
        RECT 391.050 221.400 392.850 233.400 ;
        RECT 375.150 220.500 383.550 220.800 ;
        RECT 391.950 220.500 392.850 221.400 ;
        RECT 394.950 220.950 397.050 223.050 ;
        RECT 406.800 221.400 408.600 233.400 ;
        RECT 409.800 222.300 411.600 233.400 ;
        RECT 415.800 222.300 417.600 233.400 ;
        RECT 421.950 226.950 424.050 229.050 ;
        RECT 409.800 221.400 417.600 222.300 ;
        RECT 375.150 219.900 392.850 220.500 ;
        RECT 381.750 219.300 392.850 219.900 ;
        RECT 381.750 219.000 383.550 219.300 ;
        RECT 379.950 212.400 382.050 214.050 ;
        RECT 379.950 211.200 387.900 212.400 ;
        RECT 388.950 211.950 391.050 214.050 ;
        RECT 386.100 210.600 387.900 211.200 ;
        RECT 389.100 210.150 390.900 211.950 ;
        RECT 383.100 209.400 384.900 210.000 ;
        RECT 389.100 209.400 390.000 210.150 ;
        RECT 383.100 208.200 390.000 209.400 ;
        RECT 372.150 207.000 384.150 208.200 ;
        RECT 372.150 206.400 373.950 207.000 ;
        RECT 383.100 205.200 384.150 207.000 ;
        RECT 359.550 198.600 361.350 204.600 ;
        RECT 364.950 203.700 367.050 204.600 ;
        RECT 364.950 202.500 368.700 203.700 ;
        RECT 379.350 203.550 381.150 204.300 ;
        RECT 367.650 201.600 368.700 202.500 ;
        RECT 376.200 202.500 381.150 203.550 ;
        RECT 382.650 203.400 384.450 205.200 ;
        RECT 391.950 204.600 392.850 219.300 ;
        RECT 385.950 202.500 388.050 204.600 ;
        RECT 376.200 201.600 377.250 202.500 ;
        RECT 385.950 201.600 387.000 202.500 ;
        RECT 367.650 198.600 369.450 201.600 ;
        RECT 375.450 198.600 377.250 201.600 ;
        RECT 383.250 200.700 387.000 201.600 ;
        RECT 383.250 198.600 385.050 200.700 ;
        RECT 391.050 198.600 392.850 204.600 ;
        RECT 395.550 202.050 396.450 220.950 ;
        RECT 407.400 214.050 408.600 221.400 ;
        RECT 409.950 214.950 412.050 217.050 ;
        RECT 406.950 211.950 409.050 214.050 ;
        RECT 410.100 213.150 411.900 214.950 ;
        RECT 413.100 214.050 414.900 215.850 ;
        RECT 415.950 214.950 418.050 217.050 ;
        RECT 412.950 211.950 415.050 214.050 ;
        RECT 416.100 213.150 417.900 214.950 ;
        RECT 407.400 204.600 408.600 211.950 ;
        RECT 422.550 208.050 423.450 226.950 ;
        RECT 433.500 222.600 435.300 233.400 ;
        RECT 442.950 229.950 445.050 232.050 ;
        RECT 431.700 221.400 435.300 222.600 ;
        RECT 431.700 214.050 432.600 221.400 ;
        RECT 428.100 211.050 429.900 212.850 ;
        RECT 430.950 211.950 433.050 214.050 ;
        RECT 427.950 208.950 430.050 211.050 ;
        RECT 421.950 205.950 424.050 208.050 ;
        RECT 407.400 203.400 412.500 204.600 ;
        RECT 394.950 199.950 397.050 202.050 ;
        RECT 410.700 198.600 412.500 203.400 ;
        RECT 431.700 201.600 432.600 211.950 ;
        RECT 434.100 211.050 435.900 212.850 ;
        RECT 433.950 208.950 436.050 211.050 ;
        RECT 443.550 205.050 444.450 229.950 ;
        RECT 449.400 222.300 451.200 233.400 ;
        RECT 455.400 222.300 457.200 233.400 ;
        RECT 449.400 221.400 457.200 222.300 ;
        RECT 458.400 221.400 460.200 233.400 ;
        RECT 465.150 221.400 466.950 233.400 ;
        RECT 473.550 227.400 475.350 233.400 ;
        RECT 473.550 226.500 474.750 227.400 ;
        RECT 481.350 226.500 483.150 233.400 ;
        RECT 489.150 227.400 490.950 233.400 ;
        RECT 469.950 224.400 474.750 226.500 ;
        RECT 477.450 225.450 484.050 226.500 ;
        RECT 477.450 224.700 479.250 225.450 ;
        RECT 482.250 224.700 484.050 225.450 ;
        RECT 489.150 225.300 493.050 227.400 ;
        RECT 473.550 223.500 474.750 224.400 ;
        RECT 486.450 223.800 488.250 224.400 ;
        RECT 473.550 222.300 481.050 223.500 ;
        RECT 479.250 221.700 481.050 222.300 ;
        RECT 481.950 222.900 488.250 223.800 ;
        RECT 448.950 214.950 451.050 217.050 ;
        RECT 449.100 213.150 450.900 214.950 ;
        RECT 452.100 214.050 453.900 215.850 ;
        RECT 454.950 214.950 457.050 217.050 ;
        RECT 451.950 211.950 454.050 214.050 ;
        RECT 455.100 213.150 456.900 214.950 ;
        RECT 458.400 214.050 459.600 221.400 ;
        RECT 465.150 220.500 466.050 221.400 ;
        RECT 481.950 220.800 482.850 222.900 ;
        RECT 486.450 222.600 488.250 222.900 ;
        RECT 489.150 222.600 491.850 224.400 ;
        RECT 489.150 221.700 490.050 222.600 ;
        RECT 474.450 220.500 482.850 220.800 ;
        RECT 465.150 219.900 482.850 220.500 ;
        RECT 484.950 220.800 490.050 221.700 ;
        RECT 490.950 220.800 493.050 221.700 ;
        RECT 496.650 221.400 498.450 233.400 ;
        RECT 514.500 222.600 516.300 233.400 ;
        RECT 535.800 227.400 537.600 233.400 ;
        RECT 557.400 227.400 559.200 233.400 ;
        RECT 465.150 219.300 476.250 219.900 ;
        RECT 457.950 211.950 460.050 214.050 ;
        RECT 442.950 202.950 445.050 205.050 ;
        RECT 458.400 204.600 459.600 211.950 ;
        RECT 454.500 203.400 459.600 204.600 ;
        RECT 465.150 204.600 466.050 219.300 ;
        RECT 474.450 219.000 476.250 219.300 ;
        RECT 466.950 211.950 469.050 214.050 ;
        RECT 475.950 212.400 478.050 214.050 ;
        RECT 467.100 210.150 468.900 211.950 ;
        RECT 470.100 211.200 478.050 212.400 ;
        RECT 470.100 210.600 471.900 211.200 ;
        RECT 468.000 209.400 468.900 210.150 ;
        RECT 473.100 209.400 474.900 210.000 ;
        RECT 468.000 208.200 474.900 209.400 ;
        RECT 484.950 208.200 485.850 220.800 ;
        RECT 490.950 219.600 495.150 220.800 ;
        RECT 494.250 217.800 496.050 219.600 ;
        RECT 497.250 214.050 498.450 221.400 ;
        RECT 512.700 221.400 516.300 222.600 ;
        RECT 512.700 214.050 513.600 221.400 ;
        RECT 532.950 214.950 535.050 217.050 ;
        RECT 493.950 213.750 498.450 214.050 ;
        RECT 492.150 211.950 498.450 213.750 ;
        RECT 473.850 207.000 485.850 208.200 ;
        RECT 473.850 205.200 474.900 207.000 ;
        RECT 484.050 206.400 485.850 207.000 ;
        RECT 431.400 198.600 433.200 201.600 ;
        RECT 454.500 198.600 456.300 203.400 ;
        RECT 465.150 198.600 466.950 204.600 ;
        RECT 469.950 202.500 472.050 204.600 ;
        RECT 473.550 203.400 475.350 205.200 ;
        RECT 497.250 204.600 498.450 211.950 ;
        RECT 509.100 211.050 510.900 212.850 ;
        RECT 511.950 211.950 514.050 214.050 ;
        RECT 533.100 213.150 534.900 214.950 ;
        RECT 536.400 214.050 537.600 227.400 ;
        RECT 538.950 214.950 541.050 217.050 ;
        RECT 553.950 214.950 556.050 217.050 ;
        RECT 508.950 208.950 511.050 211.050 ;
        RECT 476.850 203.550 478.650 204.300 ;
        RECT 490.950 203.700 493.050 204.600 ;
        RECT 476.850 202.500 481.800 203.550 ;
        RECT 471.000 201.600 472.050 202.500 ;
        RECT 480.750 201.600 481.800 202.500 ;
        RECT 489.300 202.500 493.050 203.700 ;
        RECT 489.300 201.600 490.350 202.500 ;
        RECT 471.000 200.700 474.750 201.600 ;
        RECT 472.950 198.600 474.750 200.700 ;
        RECT 480.750 198.600 482.550 201.600 ;
        RECT 488.550 198.600 490.350 201.600 ;
        RECT 496.650 198.600 498.450 204.600 ;
        RECT 512.700 201.600 513.600 211.950 ;
        RECT 515.100 211.050 516.900 212.850 ;
        RECT 535.950 211.950 538.050 214.050 ;
        RECT 539.100 213.150 540.900 214.950 ;
        RECT 554.100 213.150 555.900 214.950 ;
        RECT 557.850 214.050 559.050 227.400 ;
        RECT 567.150 221.400 568.950 233.400 ;
        RECT 575.550 227.400 577.350 233.400 ;
        RECT 575.550 226.500 576.750 227.400 ;
        RECT 583.350 226.500 585.150 233.400 ;
        RECT 591.150 227.400 592.950 233.400 ;
        RECT 571.950 224.400 576.750 226.500 ;
        RECT 579.450 225.450 586.050 226.500 ;
        RECT 579.450 224.700 581.250 225.450 ;
        RECT 584.250 224.700 586.050 225.450 ;
        RECT 591.150 225.300 595.050 227.400 ;
        RECT 575.550 223.500 576.750 224.400 ;
        RECT 588.450 223.800 590.250 224.400 ;
        RECT 575.550 222.300 583.050 223.500 ;
        RECT 581.250 221.700 583.050 222.300 ;
        RECT 583.950 222.900 590.250 223.800 ;
        RECT 567.150 220.500 568.050 221.400 ;
        RECT 583.950 220.800 584.850 222.900 ;
        RECT 588.450 222.600 590.250 222.900 ;
        RECT 591.150 222.600 593.850 224.400 ;
        RECT 591.150 221.700 592.050 222.600 ;
        RECT 576.450 220.500 584.850 220.800 ;
        RECT 567.150 219.900 584.850 220.500 ;
        RECT 586.950 220.800 592.050 221.700 ;
        RECT 592.950 220.800 595.050 221.700 ;
        RECT 598.650 221.400 600.450 233.400 ;
        RECT 567.150 219.300 578.250 219.900 ;
        RECT 559.950 214.950 562.050 217.050 ;
        RECT 556.950 211.950 559.050 214.050 ;
        RECT 560.100 213.150 561.900 214.950 ;
        RECT 563.100 214.050 564.900 215.850 ;
        RECT 562.950 211.950 565.050 214.050 ;
        RECT 514.950 208.950 517.050 211.050 ;
        RECT 536.400 206.700 537.600 211.950 ;
        RECT 556.950 207.750 558.150 211.950 ;
        RECT 533.400 205.800 537.600 206.700 ;
        RECT 554.400 206.700 558.150 207.750 ;
        RECT 512.400 198.600 514.200 201.600 ;
        RECT 533.400 198.600 535.200 205.800 ;
        RECT 554.400 204.600 555.600 206.700 ;
        RECT 553.800 198.600 555.600 204.600 ;
        RECT 556.800 203.700 564.600 205.050 ;
        RECT 556.800 198.600 558.600 203.700 ;
        RECT 562.800 198.600 564.600 203.700 ;
        RECT 567.150 204.600 568.050 219.300 ;
        RECT 576.450 219.000 578.250 219.300 ;
        RECT 568.950 211.950 571.050 214.050 ;
        RECT 577.950 212.400 580.050 214.050 ;
        RECT 569.100 210.150 570.900 211.950 ;
        RECT 572.100 211.200 580.050 212.400 ;
        RECT 572.100 210.600 573.900 211.200 ;
        RECT 570.000 209.400 570.900 210.150 ;
        RECT 575.100 209.400 576.900 210.000 ;
        RECT 570.000 208.200 576.900 209.400 ;
        RECT 586.950 208.200 587.850 220.800 ;
        RECT 592.950 219.600 597.150 220.800 ;
        RECT 596.250 217.800 598.050 219.600 ;
        RECT 599.250 214.050 600.450 221.400 ;
        RECT 614.400 227.400 616.200 233.400 ;
        RECT 634.800 227.400 636.600 233.400 ;
        RECT 659.400 227.400 661.200 233.400 ;
        RECT 614.400 220.050 615.600 227.400 ;
        RECT 611.100 214.050 612.900 215.850 ;
        RECT 613.950 214.950 616.050 220.050 ;
        RECT 595.950 213.750 600.450 214.050 ;
        RECT 594.150 211.950 600.450 213.750 ;
        RECT 610.950 211.950 613.050 214.050 ;
        RECT 575.850 207.000 587.850 208.200 ;
        RECT 575.850 205.200 576.900 207.000 ;
        RECT 586.050 206.400 587.850 207.000 ;
        RECT 567.150 198.600 568.950 204.600 ;
        RECT 571.950 202.500 574.050 204.600 ;
        RECT 575.550 203.400 577.350 205.200 ;
        RECT 599.250 204.600 600.450 211.950 ;
        RECT 578.850 203.550 580.650 204.300 ;
        RECT 592.950 203.700 595.050 204.600 ;
        RECT 578.850 202.500 583.800 203.550 ;
        RECT 573.000 201.600 574.050 202.500 ;
        RECT 582.750 201.600 583.800 202.500 ;
        RECT 591.300 202.500 595.050 203.700 ;
        RECT 591.300 201.600 592.350 202.500 ;
        RECT 573.000 200.700 576.750 201.600 ;
        RECT 574.950 198.600 576.750 200.700 ;
        RECT 582.750 198.600 584.550 201.600 ;
        RECT 590.550 198.600 592.350 201.600 ;
        RECT 598.650 198.600 600.450 204.600 ;
        RECT 614.400 201.600 615.600 214.950 ;
        RECT 629.100 214.050 630.900 215.850 ;
        RECT 631.950 214.950 634.050 217.050 ;
        RECT 628.950 211.950 631.050 214.050 ;
        RECT 632.100 213.150 633.900 214.950 ;
        RECT 634.950 214.050 636.150 227.400 ;
        RECT 637.950 214.950 640.050 217.050 ;
        RECT 655.950 214.950 658.050 217.050 ;
        RECT 634.950 211.950 637.050 214.050 ;
        RECT 638.100 213.150 639.900 214.950 ;
        RECT 656.100 213.150 657.900 214.950 ;
        RECT 659.850 214.050 661.050 227.400 ;
        RECT 682.500 222.600 684.300 233.400 ;
        RECT 703.500 222.600 705.300 233.400 ;
        RECT 724.800 227.400 726.600 233.400 ;
        RECT 748.800 227.400 750.600 233.400 ;
        RECT 680.700 221.400 684.300 222.600 ;
        RECT 701.700 221.400 705.300 222.600 ;
        RECT 661.950 214.950 664.050 217.050 ;
        RECT 635.850 207.750 637.050 211.950 ;
        RECT 658.950 211.950 661.050 214.050 ;
        RECT 662.100 213.150 663.900 214.950 ;
        RECT 665.100 214.050 666.900 215.850 ;
        RECT 680.700 214.050 681.600 221.400 ;
        RECT 688.950 214.950 691.050 217.050 ;
        RECT 664.950 211.950 667.050 214.050 ;
        RECT 658.950 207.750 660.150 211.950 ;
        RECT 677.100 211.050 678.900 212.850 ;
        RECT 679.950 211.950 682.050 214.050 ;
        RECT 676.950 208.950 679.050 211.050 ;
        RECT 635.850 206.700 639.600 207.750 ;
        RECT 629.400 203.700 637.200 205.050 ;
        RECT 614.400 198.600 616.200 201.600 ;
        RECT 629.400 198.600 631.200 203.700 ;
        RECT 635.400 198.600 637.200 203.700 ;
        RECT 638.400 204.600 639.600 206.700 ;
        RECT 656.400 206.700 660.150 207.750 ;
        RECT 656.400 204.600 657.600 206.700 ;
        RECT 638.400 198.600 640.200 204.600 ;
        RECT 655.800 198.600 657.600 204.600 ;
        RECT 658.800 203.700 666.600 205.050 ;
        RECT 658.800 198.600 660.600 203.700 ;
        RECT 664.800 198.600 666.600 203.700 ;
        RECT 680.700 201.600 681.600 211.950 ;
        RECT 683.100 211.050 684.900 212.850 ;
        RECT 682.950 208.950 685.050 211.050 ;
        RECT 689.550 202.050 690.450 214.950 ;
        RECT 701.700 214.050 702.600 221.400 ;
        RECT 719.100 214.050 720.900 215.850 ;
        RECT 721.950 214.950 724.050 217.050 ;
        RECT 698.100 211.050 699.900 212.850 ;
        RECT 700.950 211.950 703.050 214.050 ;
        RECT 697.950 208.950 700.050 211.050 ;
        RECT 680.400 198.600 682.200 201.600 ;
        RECT 688.950 199.950 691.050 202.050 ;
        RECT 701.700 201.600 702.600 211.950 ;
        RECT 704.100 211.050 705.900 212.850 ;
        RECT 718.950 211.950 721.050 214.050 ;
        RECT 722.100 213.150 723.900 214.950 ;
        RECT 724.950 214.050 726.150 227.400 ;
        RECT 727.950 214.950 730.050 217.050 ;
        RECT 745.950 214.950 748.050 217.050 ;
        RECT 724.950 211.950 727.050 214.050 ;
        RECT 728.100 213.150 729.900 214.950 ;
        RECT 746.100 213.150 747.900 214.950 ;
        RECT 749.400 214.050 750.600 227.400 ;
        RECT 767.400 227.400 769.200 233.400 ;
        RECT 751.950 214.950 754.050 217.050 ;
        RECT 763.950 214.950 766.050 217.050 ;
        RECT 748.950 211.950 751.050 214.050 ;
        RECT 752.100 213.150 753.900 214.950 ;
        RECT 764.100 213.150 765.900 214.950 ;
        RECT 767.400 214.050 768.600 227.400 ;
        RECT 776.550 221.400 778.350 233.400 ;
        RECT 784.050 227.400 785.850 233.400 ;
        RECT 781.950 225.300 785.850 227.400 ;
        RECT 791.850 226.500 793.650 233.400 ;
        RECT 799.650 227.400 801.450 233.400 ;
        RECT 800.250 226.500 801.450 227.400 ;
        RECT 790.950 225.450 797.550 226.500 ;
        RECT 790.950 224.700 792.750 225.450 ;
        RECT 795.750 224.700 797.550 225.450 ;
        RECT 800.250 224.400 805.050 226.500 ;
        RECT 783.150 222.600 785.850 224.400 ;
        RECT 786.750 223.800 788.550 224.400 ;
        RECT 786.750 222.900 793.050 223.800 ;
        RECT 800.250 223.500 801.450 224.400 ;
        RECT 786.750 222.600 788.550 222.900 ;
        RECT 784.950 221.700 785.850 222.600 ;
        RECT 769.950 214.950 772.050 217.050 ;
        RECT 766.950 211.950 769.050 214.050 ;
        RECT 770.100 213.150 771.900 214.950 ;
        RECT 776.550 214.050 777.750 221.400 ;
        RECT 781.950 220.800 784.050 221.700 ;
        RECT 784.950 220.800 790.050 221.700 ;
        RECT 779.850 219.600 784.050 220.800 ;
        RECT 778.950 217.800 780.750 219.600 ;
        RECT 776.550 213.750 781.050 214.050 ;
        RECT 776.550 211.950 782.850 213.750 ;
        RECT 703.950 208.950 706.050 211.050 ;
        RECT 725.850 207.750 727.050 211.950 ;
        RECT 725.850 206.700 729.600 207.750 ;
        RECT 749.400 206.700 750.600 211.950 ;
        RECT 719.400 203.700 727.200 205.050 ;
        RECT 701.400 198.600 703.200 201.600 ;
        RECT 719.400 198.600 721.200 203.700 ;
        RECT 725.400 198.600 727.200 203.700 ;
        RECT 728.400 204.600 729.600 206.700 ;
        RECT 746.400 205.800 750.600 206.700 ;
        RECT 767.400 206.700 768.600 211.950 ;
        RECT 767.400 205.800 771.600 206.700 ;
        RECT 728.400 198.600 730.200 204.600 ;
        RECT 746.400 198.600 748.200 205.800 ;
        RECT 769.800 198.600 771.600 205.800 ;
        RECT 776.550 204.600 777.750 211.950 ;
        RECT 789.150 208.200 790.050 220.800 ;
        RECT 792.150 220.800 793.050 222.900 ;
        RECT 793.950 222.300 801.450 223.500 ;
        RECT 793.950 221.700 795.750 222.300 ;
        RECT 808.050 221.400 809.850 233.400 ;
        RECT 792.150 220.500 800.550 220.800 ;
        RECT 808.950 220.500 809.850 221.400 ;
        RECT 792.150 219.900 809.850 220.500 ;
        RECT 798.750 219.300 809.850 219.900 ;
        RECT 798.750 219.000 800.550 219.300 ;
        RECT 796.950 212.400 799.050 214.050 ;
        RECT 796.950 211.200 804.900 212.400 ;
        RECT 805.950 211.950 808.050 214.050 ;
        RECT 803.100 210.600 804.900 211.200 ;
        RECT 806.100 210.150 807.900 211.950 ;
        RECT 800.100 209.400 801.900 210.000 ;
        RECT 806.100 209.400 807.000 210.150 ;
        RECT 800.100 208.200 807.000 209.400 ;
        RECT 789.150 207.000 801.150 208.200 ;
        RECT 789.150 206.400 790.950 207.000 ;
        RECT 800.100 205.200 801.150 207.000 ;
        RECT 776.550 198.600 778.350 204.600 ;
        RECT 781.950 203.700 784.050 204.600 ;
        RECT 781.950 202.500 785.700 203.700 ;
        RECT 796.350 203.550 798.150 204.300 ;
        RECT 784.650 201.600 785.700 202.500 ;
        RECT 793.200 202.500 798.150 203.550 ;
        RECT 799.650 203.400 801.450 205.200 ;
        RECT 808.950 204.600 809.850 219.300 ;
        RECT 802.950 202.500 805.050 204.600 ;
        RECT 793.200 201.600 794.250 202.500 ;
        RECT 802.950 201.600 804.000 202.500 ;
        RECT 784.650 198.600 786.450 201.600 ;
        RECT 792.450 198.600 794.250 201.600 ;
        RECT 800.250 200.700 804.000 201.600 ;
        RECT 800.250 198.600 802.050 200.700 ;
        RECT 808.050 198.600 809.850 204.600 ;
        RECT 812.550 221.400 814.350 233.400 ;
        RECT 820.050 227.400 821.850 233.400 ;
        RECT 817.950 225.300 821.850 227.400 ;
        RECT 827.850 226.500 829.650 233.400 ;
        RECT 835.650 227.400 837.450 233.400 ;
        RECT 836.250 226.500 837.450 227.400 ;
        RECT 826.950 225.450 833.550 226.500 ;
        RECT 826.950 224.700 828.750 225.450 ;
        RECT 831.750 224.700 833.550 225.450 ;
        RECT 836.250 224.400 841.050 226.500 ;
        RECT 819.150 222.600 821.850 224.400 ;
        RECT 822.750 223.800 824.550 224.400 ;
        RECT 822.750 222.900 829.050 223.800 ;
        RECT 836.250 223.500 837.450 224.400 ;
        RECT 822.750 222.600 824.550 222.900 ;
        RECT 820.950 221.700 821.850 222.600 ;
        RECT 812.550 214.050 813.750 221.400 ;
        RECT 817.950 220.800 820.050 221.700 ;
        RECT 820.950 220.800 826.050 221.700 ;
        RECT 815.850 219.600 820.050 220.800 ;
        RECT 814.950 217.800 816.750 219.600 ;
        RECT 812.550 213.750 817.050 214.050 ;
        RECT 812.550 211.950 818.850 213.750 ;
        RECT 812.550 204.600 813.750 211.950 ;
        RECT 825.150 208.200 826.050 220.800 ;
        RECT 828.150 220.800 829.050 222.900 ;
        RECT 829.950 222.300 837.450 223.500 ;
        RECT 829.950 221.700 831.750 222.300 ;
        RECT 844.050 221.400 845.850 233.400 ;
        RECT 828.150 220.500 836.550 220.800 ;
        RECT 844.950 220.500 845.850 221.400 ;
        RECT 828.150 219.900 845.850 220.500 ;
        RECT 834.750 219.300 845.850 219.900 ;
        RECT 834.750 219.000 836.550 219.300 ;
        RECT 832.950 212.400 835.050 214.050 ;
        RECT 832.950 211.200 840.900 212.400 ;
        RECT 841.950 211.950 844.050 214.050 ;
        RECT 839.100 210.600 840.900 211.200 ;
        RECT 842.100 210.150 843.900 211.950 ;
        RECT 836.100 209.400 837.900 210.000 ;
        RECT 842.100 209.400 843.000 210.150 ;
        RECT 836.100 208.200 843.000 209.400 ;
        RECT 825.150 207.000 837.150 208.200 ;
        RECT 825.150 206.400 826.950 207.000 ;
        RECT 836.100 205.200 837.150 207.000 ;
        RECT 812.550 198.600 814.350 204.600 ;
        RECT 817.950 203.700 820.050 204.600 ;
        RECT 817.950 202.500 821.700 203.700 ;
        RECT 832.350 203.550 834.150 204.300 ;
        RECT 820.650 201.600 821.700 202.500 ;
        RECT 829.200 202.500 834.150 203.550 ;
        RECT 835.650 203.400 837.450 205.200 ;
        RECT 844.950 204.600 845.850 219.300 ;
        RECT 838.950 202.500 841.050 204.600 ;
        RECT 829.200 201.600 830.250 202.500 ;
        RECT 838.950 201.600 840.000 202.500 ;
        RECT 820.650 198.600 822.450 201.600 ;
        RECT 828.450 198.600 830.250 201.600 ;
        RECT 836.250 200.700 840.000 201.600 ;
        RECT 836.250 198.600 838.050 200.700 ;
        RECT 844.050 198.600 845.850 204.600 ;
        RECT 849.150 221.400 850.950 233.400 ;
        RECT 857.550 227.400 859.350 233.400 ;
        RECT 857.550 226.500 858.750 227.400 ;
        RECT 865.350 226.500 867.150 233.400 ;
        RECT 873.150 227.400 874.950 233.400 ;
        RECT 853.950 224.400 858.750 226.500 ;
        RECT 861.450 225.450 868.050 226.500 ;
        RECT 861.450 224.700 863.250 225.450 ;
        RECT 866.250 224.700 868.050 225.450 ;
        RECT 873.150 225.300 877.050 227.400 ;
        RECT 857.550 223.500 858.750 224.400 ;
        RECT 870.450 223.800 872.250 224.400 ;
        RECT 857.550 222.300 865.050 223.500 ;
        RECT 863.250 221.700 865.050 222.300 ;
        RECT 865.950 222.900 872.250 223.800 ;
        RECT 849.150 220.500 850.050 221.400 ;
        RECT 865.950 220.800 866.850 222.900 ;
        RECT 870.450 222.600 872.250 222.900 ;
        RECT 873.150 222.600 875.850 224.400 ;
        RECT 873.150 221.700 874.050 222.600 ;
        RECT 858.450 220.500 866.850 220.800 ;
        RECT 849.150 219.900 866.850 220.500 ;
        RECT 868.950 220.800 874.050 221.700 ;
        RECT 874.950 220.800 877.050 221.700 ;
        RECT 880.650 221.400 882.450 233.400 ;
        RECT 883.950 229.950 886.050 232.050 ;
        RECT 849.150 219.300 860.250 219.900 ;
        RECT 849.150 204.600 850.050 219.300 ;
        RECT 858.450 219.000 860.250 219.300 ;
        RECT 850.950 211.950 853.050 214.050 ;
        RECT 859.950 212.400 862.050 214.050 ;
        RECT 851.100 210.150 852.900 211.950 ;
        RECT 854.100 211.200 862.050 212.400 ;
        RECT 854.100 210.600 855.900 211.200 ;
        RECT 852.000 209.400 852.900 210.150 ;
        RECT 857.100 209.400 858.900 210.000 ;
        RECT 852.000 208.200 858.900 209.400 ;
        RECT 868.950 208.200 869.850 220.800 ;
        RECT 874.950 219.600 879.150 220.800 ;
        RECT 878.250 217.800 880.050 219.600 ;
        RECT 881.250 214.050 882.450 221.400 ;
        RECT 877.950 213.750 882.450 214.050 ;
        RECT 876.150 211.950 882.450 213.750 ;
        RECT 857.850 207.000 869.850 208.200 ;
        RECT 857.850 205.200 858.900 207.000 ;
        RECT 868.050 206.400 869.850 207.000 ;
        RECT 849.150 198.600 850.950 204.600 ;
        RECT 853.950 202.500 856.050 204.600 ;
        RECT 857.550 203.400 859.350 205.200 ;
        RECT 881.250 204.600 882.450 211.950 ;
        RECT 860.850 203.550 862.650 204.300 ;
        RECT 874.950 203.700 877.050 204.600 ;
        RECT 860.850 202.500 865.800 203.550 ;
        RECT 855.000 201.600 856.050 202.500 ;
        RECT 864.750 201.600 865.800 202.500 ;
        RECT 873.300 202.500 877.050 203.700 ;
        RECT 873.300 201.600 874.350 202.500 ;
        RECT 855.000 200.700 858.750 201.600 ;
        RECT 856.950 198.600 858.750 200.700 ;
        RECT 864.750 198.600 866.550 201.600 ;
        RECT 872.550 198.600 874.350 201.600 ;
        RECT 880.650 198.600 882.450 204.600 ;
        RECT 884.550 202.050 885.450 229.950 ;
        RECT 895.800 221.400 897.600 233.400 ;
        RECT 898.800 222.300 900.600 233.400 ;
        RECT 904.800 222.300 906.600 233.400 ;
        RECT 898.800 221.400 906.600 222.300 ;
        RECT 896.400 214.050 897.600 221.400 ;
        RECT 898.950 214.950 901.050 217.050 ;
        RECT 895.950 211.950 898.050 214.050 ;
        RECT 899.100 213.150 900.900 214.950 ;
        RECT 902.100 214.050 903.900 215.850 ;
        RECT 904.950 214.950 907.050 217.050 ;
        RECT 901.950 211.950 904.050 214.050 ;
        RECT 905.100 213.150 906.900 214.950 ;
        RECT 896.400 204.600 897.600 211.950 ;
        RECT 896.400 203.400 901.500 204.600 ;
        RECT 883.950 199.950 886.050 202.050 ;
        RECT 899.700 198.600 901.500 203.400 ;
        RECT 16.800 191.400 18.600 194.400 ;
        RECT 13.950 181.950 16.050 184.050 ;
        RECT 14.100 180.150 15.900 181.950 ;
        RECT 17.400 181.050 18.300 191.400 ;
        RECT 32.400 189.300 34.200 194.400 ;
        RECT 38.400 189.300 40.200 194.400 ;
        RECT 32.400 187.950 40.200 189.300 ;
        RECT 41.400 188.400 43.200 194.400 ;
        RECT 59.400 191.400 61.200 194.400 ;
        RECT 41.400 186.300 42.600 188.400 ;
        RECT 38.850 185.250 42.600 186.300 ;
        RECT 19.950 181.950 22.050 184.050 ;
        RECT 16.950 178.950 19.050 181.050 ;
        RECT 20.100 180.150 21.900 181.950 ;
        RECT 38.850 181.050 40.050 185.250 ;
        RECT 31.950 178.950 34.050 181.050 ;
        RECT 17.400 171.600 18.300 178.950 ;
        RECT 32.100 177.150 33.900 178.950 ;
        RECT 35.100 178.050 36.900 179.850 ;
        RECT 37.950 178.950 40.050 181.050 ;
        RECT 34.950 175.950 37.050 178.050 ;
        RECT 14.700 170.400 18.300 171.600 ;
        RECT 14.700 159.600 16.500 170.400 ;
        RECT 37.950 165.600 39.150 178.950 ;
        RECT 41.100 178.050 42.900 179.850 ;
        RECT 55.950 178.950 58.050 181.050 ;
        RECT 40.950 175.950 43.050 178.050 ;
        RECT 56.100 177.150 57.900 178.950 ;
        RECT 59.400 178.050 60.600 191.400 ;
        RECT 79.800 187.200 81.600 194.400 ;
        RECT 98.400 191.400 100.200 194.400 ;
        RECT 119.400 191.400 121.200 194.400 ;
        RECT 137.400 191.400 139.200 194.400 ;
        RECT 77.400 186.300 81.600 187.200 ;
        RECT 77.400 181.050 78.600 186.300 ;
        RECT 88.950 181.950 91.050 184.050 ;
        RECT 94.950 181.950 97.050 184.050 ;
        RECT 74.100 178.050 75.900 179.850 ;
        RECT 76.950 178.950 79.050 181.050 ;
        RECT 58.950 172.950 61.050 178.050 ;
        RECT 73.950 175.950 76.050 178.050 ;
        RECT 59.400 165.600 60.600 172.950 ;
        RECT 77.400 165.600 78.600 178.950 ;
        RECT 80.100 178.050 81.900 179.850 ;
        RECT 79.950 175.950 82.050 178.050 ;
        RECT 37.800 159.600 39.600 165.600 ;
        RECT 59.400 159.600 61.200 165.600 ;
        RECT 77.400 159.600 79.200 165.600 ;
        RECT 89.550 163.050 90.450 181.950 ;
        RECT 95.100 180.150 96.900 181.950 ;
        RECT 98.700 181.050 99.600 191.400 ;
        RECT 100.950 181.950 103.050 184.050 ;
        RECT 97.950 178.950 100.050 181.050 ;
        RECT 101.100 180.150 102.900 181.950 ;
        RECT 115.950 178.950 118.050 181.050 ;
        RECT 98.700 171.600 99.600 178.950 ;
        RECT 116.100 177.150 117.900 178.950 ;
        RECT 119.400 178.050 120.600 191.400 ;
        RECT 133.950 178.950 136.050 181.050 ;
        RECT 118.950 172.950 121.050 178.050 ;
        RECT 134.100 177.150 135.900 178.950 ;
        RECT 137.400 178.050 138.600 191.400 ;
        RECT 143.550 188.400 145.350 194.400 ;
        RECT 151.650 191.400 153.450 194.400 ;
        RECT 159.450 191.400 161.250 194.400 ;
        RECT 167.250 192.300 169.050 194.400 ;
        RECT 167.250 191.400 171.000 192.300 ;
        RECT 151.650 190.500 152.700 191.400 ;
        RECT 148.950 189.300 152.700 190.500 ;
        RECT 160.200 190.500 161.250 191.400 ;
        RECT 169.950 190.500 171.000 191.400 ;
        RECT 160.200 189.450 165.150 190.500 ;
        RECT 148.950 188.400 151.050 189.300 ;
        RECT 163.350 188.700 165.150 189.450 ;
        RECT 143.550 181.050 144.750 188.400 ;
        RECT 166.650 187.800 168.450 189.600 ;
        RECT 169.950 188.400 172.050 190.500 ;
        RECT 175.050 188.400 176.850 194.400 ;
        RECT 156.150 186.000 157.950 186.600 ;
        RECT 167.100 186.000 168.150 187.800 ;
        RECT 156.150 184.800 168.150 186.000 ;
        RECT 143.550 179.250 149.850 181.050 ;
        RECT 143.550 178.950 148.050 179.250 ;
        RECT 136.950 172.950 139.050 178.050 ;
        RECT 98.700 170.400 102.300 171.600 ;
        RECT 88.950 160.950 91.050 163.050 ;
        RECT 100.500 159.600 102.300 170.400 ;
        RECT 119.400 165.600 120.600 172.950 ;
        RECT 137.400 165.600 138.600 172.950 ;
        RECT 143.550 171.600 144.750 178.950 ;
        RECT 145.950 173.400 147.750 175.200 ;
        RECT 146.850 172.200 151.050 173.400 ;
        RECT 156.150 172.200 157.050 184.800 ;
        RECT 167.100 183.600 174.000 184.800 ;
        RECT 167.100 183.000 168.900 183.600 ;
        RECT 173.100 182.850 174.000 183.600 ;
        RECT 170.100 181.800 171.900 182.400 ;
        RECT 163.950 180.600 171.900 181.800 ;
        RECT 173.100 181.050 174.900 182.850 ;
        RECT 163.950 178.950 166.050 180.600 ;
        RECT 172.950 178.950 175.050 181.050 ;
        RECT 165.750 173.700 167.550 174.000 ;
        RECT 175.950 173.700 176.850 188.400 ;
        RECT 188.400 189.300 190.200 194.400 ;
        RECT 194.400 189.300 196.200 194.400 ;
        RECT 188.400 187.950 196.200 189.300 ;
        RECT 197.400 188.400 199.200 194.400 ;
        RECT 197.400 186.300 198.600 188.400 ;
        RECT 217.800 187.500 219.600 194.400 ;
        RECT 223.800 187.500 225.600 194.400 ;
        RECT 229.800 187.500 231.600 194.400 ;
        RECT 235.800 187.500 237.600 194.400 ;
        RECT 194.850 185.250 198.600 186.300 ;
        RECT 216.900 186.300 219.600 187.500 ;
        RECT 221.700 186.300 225.600 187.500 ;
        RECT 227.700 186.300 231.600 187.500 ;
        RECT 233.700 186.300 237.600 187.500 ;
        RECT 254.400 187.200 256.200 194.400 ;
        RECT 274.500 188.400 276.300 194.400 ;
        RECT 280.800 191.400 282.600 194.400 ;
        RECT 254.400 186.300 258.600 187.200 ;
        RECT 194.850 181.050 196.050 185.250 ;
        RECT 216.900 181.050 217.800 186.300 ;
        RECT 221.700 185.400 222.900 186.300 ;
        RECT 227.700 185.400 228.900 186.300 ;
        RECT 233.700 185.400 234.900 186.300 ;
        RECT 218.700 184.200 222.900 185.400 ;
        RECT 218.700 183.600 220.500 184.200 ;
        RECT 187.950 178.950 190.050 181.050 ;
        RECT 188.100 177.150 189.900 178.950 ;
        RECT 191.100 178.050 192.900 179.850 ;
        RECT 193.950 178.950 196.050 181.050 ;
        RECT 190.950 175.950 193.050 178.050 ;
        RECT 165.750 173.100 176.850 173.700 ;
        RECT 119.400 159.600 121.200 165.600 ;
        RECT 137.400 159.600 139.200 165.600 ;
        RECT 143.550 159.600 145.350 171.600 ;
        RECT 148.950 171.300 151.050 172.200 ;
        RECT 151.950 171.300 157.050 172.200 ;
        RECT 159.150 172.500 176.850 173.100 ;
        RECT 159.150 172.200 167.550 172.500 ;
        RECT 151.950 170.400 152.850 171.300 ;
        RECT 150.150 168.600 152.850 170.400 ;
        RECT 153.750 170.100 155.550 170.400 ;
        RECT 159.150 170.100 160.050 172.200 ;
        RECT 175.950 171.600 176.850 172.500 ;
        RECT 153.750 169.200 160.050 170.100 ;
        RECT 160.950 170.700 162.750 171.300 ;
        RECT 160.950 169.500 168.450 170.700 ;
        RECT 153.750 168.600 155.550 169.200 ;
        RECT 167.250 168.600 168.450 169.500 ;
        RECT 148.950 165.600 152.850 167.700 ;
        RECT 157.950 167.550 159.750 168.300 ;
        RECT 162.750 167.550 164.550 168.300 ;
        RECT 157.950 166.500 164.550 167.550 ;
        RECT 167.250 166.500 172.050 168.600 ;
        RECT 151.050 159.600 152.850 165.600 ;
        RECT 158.850 159.600 160.650 166.500 ;
        RECT 167.250 165.600 168.450 166.500 ;
        RECT 166.650 159.600 168.450 165.600 ;
        RECT 175.050 159.600 176.850 171.600 ;
        RECT 193.950 165.600 195.150 178.950 ;
        RECT 197.100 178.050 198.900 179.850 ;
        RECT 214.950 178.950 217.800 181.050 ;
        RECT 196.950 175.950 199.050 178.050 ;
        RECT 216.900 173.700 217.800 178.950 ;
        RECT 221.700 173.700 222.900 184.200 ;
        RECT 224.700 184.200 228.900 185.400 ;
        RECT 224.700 183.600 226.500 184.200 ;
        RECT 227.700 173.700 228.900 184.200 ;
        RECT 230.700 184.200 234.900 185.400 ;
        RECT 230.700 183.600 232.500 184.200 ;
        RECT 233.700 173.700 234.900 184.200 ;
        RECT 236.100 181.050 237.900 182.850 ;
        RECT 257.400 181.050 258.600 186.300 ;
        RECT 274.500 181.050 275.700 188.400 ;
        RECT 281.400 187.500 282.600 191.400 ;
        RECT 276.600 186.600 282.600 187.500 ;
        RECT 284.550 188.400 286.350 194.400 ;
        RECT 292.650 191.400 294.450 194.400 ;
        RECT 300.450 191.400 302.250 194.400 ;
        RECT 308.250 192.300 310.050 194.400 ;
        RECT 308.250 191.400 312.000 192.300 ;
        RECT 292.650 190.500 293.700 191.400 ;
        RECT 289.950 189.300 293.700 190.500 ;
        RECT 301.200 190.500 302.250 191.400 ;
        RECT 310.950 190.500 312.000 191.400 ;
        RECT 301.200 189.450 306.150 190.500 ;
        RECT 289.950 188.400 292.050 189.300 ;
        RECT 304.350 188.700 306.150 189.450 ;
        RECT 276.600 185.700 278.850 186.600 ;
        RECT 235.950 178.950 238.050 181.050 ;
        RECT 254.100 178.050 255.900 179.850 ;
        RECT 256.950 178.950 259.050 181.050 ;
        RECT 253.950 175.950 256.050 178.050 ;
        RECT 216.900 172.500 219.600 173.700 ;
        RECT 221.700 172.500 225.600 173.700 ;
        RECT 227.700 172.500 231.600 173.700 ;
        RECT 233.700 172.500 237.600 173.700 ;
        RECT 193.800 159.600 195.600 165.600 ;
        RECT 217.800 159.600 219.600 172.500 ;
        RECT 223.800 159.600 225.600 172.500 ;
        RECT 229.800 159.600 231.600 172.500 ;
        RECT 235.800 159.600 237.600 172.500 ;
        RECT 257.400 165.600 258.600 178.950 ;
        RECT 260.100 178.050 261.900 179.850 ;
        RECT 274.500 178.950 277.050 181.050 ;
        RECT 259.950 175.950 262.050 178.050 ;
        RECT 256.800 159.600 258.600 165.600 ;
        RECT 274.500 171.600 275.700 178.950 ;
        RECT 277.950 174.300 278.850 185.700 ;
        RECT 284.550 181.050 285.750 188.400 ;
        RECT 307.650 187.800 309.450 189.600 ;
        RECT 310.950 188.400 313.050 190.500 ;
        RECT 316.050 188.400 317.850 194.400 ;
        RECT 319.950 190.950 322.050 193.050 ;
        RECT 297.150 186.000 298.950 186.600 ;
        RECT 308.100 186.000 309.150 187.800 ;
        RECT 297.150 184.800 309.150 186.000 ;
        RECT 280.950 178.950 283.050 181.050 ;
        RECT 284.550 179.250 290.850 181.050 ;
        RECT 284.550 178.950 289.050 179.250 ;
        RECT 281.100 177.150 282.900 178.950 ;
        RECT 276.600 173.400 278.850 174.300 ;
        RECT 276.600 172.500 282.600 173.400 ;
        RECT 274.500 159.600 276.300 171.600 ;
        RECT 281.400 165.600 282.600 172.500 ;
        RECT 280.800 159.600 282.600 165.600 ;
        RECT 284.550 171.600 285.750 178.950 ;
        RECT 286.950 173.400 288.750 175.200 ;
        RECT 287.850 172.200 292.050 173.400 ;
        RECT 297.150 172.200 298.050 184.800 ;
        RECT 308.100 183.600 315.000 184.800 ;
        RECT 308.100 183.000 309.900 183.600 ;
        RECT 314.100 182.850 315.000 183.600 ;
        RECT 311.100 181.800 312.900 182.400 ;
        RECT 304.950 180.600 312.900 181.800 ;
        RECT 314.100 181.050 315.900 182.850 ;
        RECT 304.950 178.950 307.050 180.600 ;
        RECT 313.950 178.950 316.050 181.050 ;
        RECT 306.750 173.700 308.550 174.000 ;
        RECT 316.950 173.700 317.850 188.400 ;
        RECT 306.750 173.100 317.850 173.700 ;
        RECT 284.550 159.600 286.350 171.600 ;
        RECT 289.950 171.300 292.050 172.200 ;
        RECT 292.950 171.300 298.050 172.200 ;
        RECT 300.150 172.500 317.850 173.100 ;
        RECT 300.150 172.200 308.550 172.500 ;
        RECT 292.950 170.400 293.850 171.300 ;
        RECT 291.150 168.600 293.850 170.400 ;
        RECT 294.750 170.100 296.550 170.400 ;
        RECT 300.150 170.100 301.050 172.200 ;
        RECT 316.950 171.600 317.850 172.500 ;
        RECT 294.750 169.200 301.050 170.100 ;
        RECT 301.950 170.700 303.750 171.300 ;
        RECT 301.950 169.500 309.450 170.700 ;
        RECT 294.750 168.600 296.550 169.200 ;
        RECT 308.250 168.600 309.450 169.500 ;
        RECT 289.950 165.600 293.850 167.700 ;
        RECT 298.950 167.550 300.750 168.300 ;
        RECT 303.750 167.550 305.550 168.300 ;
        RECT 298.950 166.500 305.550 167.550 ;
        RECT 308.250 166.500 313.050 168.600 ;
        RECT 292.050 159.600 293.850 165.600 ;
        RECT 299.850 159.600 301.650 166.500 ;
        RECT 308.250 165.600 309.450 166.500 ;
        RECT 307.650 159.600 309.450 165.600 ;
        RECT 316.050 159.600 317.850 171.600 ;
        RECT 320.550 163.050 321.450 190.950 ;
        RECT 329.400 189.300 331.200 194.400 ;
        RECT 335.400 189.300 337.200 194.400 ;
        RECT 329.400 187.950 337.200 189.300 ;
        RECT 338.400 188.400 340.200 194.400 ;
        RECT 338.400 186.300 339.600 188.400 ;
        RECT 358.800 187.200 360.600 194.400 ;
        RECT 367.950 190.950 370.050 193.050 ;
        RECT 335.850 185.250 339.600 186.300 ;
        RECT 356.400 186.300 360.600 187.200 ;
        RECT 335.850 181.050 337.050 185.250 ;
        RECT 356.400 181.050 357.600 186.300 ;
        RECT 328.950 178.950 331.050 181.050 ;
        RECT 329.100 177.150 330.900 178.950 ;
        RECT 332.100 178.050 333.900 179.850 ;
        RECT 334.950 178.950 337.050 181.050 ;
        RECT 331.950 175.950 334.050 178.050 ;
        RECT 334.950 165.600 336.150 178.950 ;
        RECT 338.100 178.050 339.900 179.850 ;
        RECT 353.100 178.050 354.900 179.850 ;
        RECT 355.950 178.950 358.050 181.050 ;
        RECT 337.950 175.950 340.050 178.050 ;
        RECT 352.950 175.950 355.050 178.050 ;
        RECT 356.400 165.600 357.600 178.950 ;
        RECT 359.100 178.050 360.900 179.850 ;
        RECT 358.950 175.950 361.050 178.050 ;
        RECT 364.950 175.950 367.050 178.050 ;
        RECT 365.550 166.050 366.450 175.950 ;
        RECT 319.950 160.950 322.050 163.050 ;
        RECT 334.800 159.600 336.600 165.600 ;
        RECT 356.400 159.600 358.200 165.600 ;
        RECT 364.950 163.950 367.050 166.050 ;
        RECT 368.550 163.050 369.450 190.950 ;
        RECT 379.800 187.500 381.600 194.400 ;
        RECT 385.800 187.500 387.600 194.400 ;
        RECT 391.800 187.500 393.600 194.400 ;
        RECT 397.800 187.500 399.600 194.400 ;
        RECT 378.900 186.300 381.600 187.500 ;
        RECT 383.700 186.300 387.600 187.500 ;
        RECT 389.700 186.300 393.600 187.500 ;
        RECT 395.700 186.300 399.600 187.500 ;
        RECT 418.800 187.200 420.600 194.400 ;
        RECT 427.950 190.950 430.050 193.050 ;
        RECT 437.400 191.400 439.200 194.400 ;
        RECT 416.400 186.300 420.600 187.200 ;
        RECT 378.900 181.050 379.800 186.300 ;
        RECT 383.700 185.400 384.900 186.300 ;
        RECT 389.700 185.400 390.900 186.300 ;
        RECT 395.700 185.400 396.900 186.300 ;
        RECT 380.700 184.200 384.900 185.400 ;
        RECT 380.700 183.600 382.500 184.200 ;
        RECT 376.950 178.950 379.800 181.050 ;
        RECT 378.900 173.700 379.800 178.950 ;
        RECT 383.700 173.700 384.900 184.200 ;
        RECT 386.700 184.200 390.900 185.400 ;
        RECT 386.700 183.600 388.500 184.200 ;
        RECT 389.700 173.700 390.900 184.200 ;
        RECT 392.700 184.200 396.900 185.400 ;
        RECT 392.700 183.600 394.500 184.200 ;
        RECT 395.700 173.700 396.900 184.200 ;
        RECT 398.100 181.050 399.900 182.850 ;
        RECT 416.400 181.050 417.600 186.300 ;
        RECT 428.550 184.050 429.450 190.950 ;
        RECT 427.950 181.950 430.050 184.050 ;
        RECT 397.950 178.950 400.050 181.050 ;
        RECT 413.100 178.050 414.900 179.850 ;
        RECT 415.950 178.950 418.050 181.050 ;
        RECT 412.950 175.950 415.050 178.050 ;
        RECT 378.900 172.500 381.600 173.700 ;
        RECT 383.700 172.500 387.600 173.700 ;
        RECT 389.700 172.500 393.600 173.700 ;
        RECT 395.700 172.500 399.600 173.700 ;
        RECT 367.950 160.950 370.050 163.050 ;
        RECT 379.800 159.600 381.600 172.500 ;
        RECT 385.800 159.600 387.600 172.500 ;
        RECT 391.800 159.600 393.600 172.500 ;
        RECT 397.800 159.600 399.600 172.500 ;
        RECT 416.400 165.600 417.600 178.950 ;
        RECT 419.100 178.050 420.900 179.850 ;
        RECT 433.950 178.950 436.050 181.050 ;
        RECT 418.950 175.950 421.050 178.050 ;
        RECT 434.100 177.150 435.900 178.950 ;
        RECT 437.400 178.050 438.600 191.400 ;
        RECT 455.400 187.500 457.200 194.400 ;
        RECT 461.400 187.500 463.200 194.400 ;
        RECT 467.400 187.500 469.200 194.400 ;
        RECT 473.400 187.500 475.200 194.400 ;
        RECT 455.400 186.300 459.300 187.500 ;
        RECT 461.400 186.300 465.300 187.500 ;
        RECT 467.400 186.300 471.300 187.500 ;
        RECT 473.400 186.300 476.100 187.500 ;
        RECT 494.400 187.200 496.200 194.400 ;
        RECT 517.800 187.200 519.600 194.400 ;
        RECT 494.400 186.300 498.600 187.200 ;
        RECT 458.100 185.400 459.300 186.300 ;
        RECT 464.100 185.400 465.300 186.300 ;
        RECT 470.100 185.400 471.300 186.300 ;
        RECT 458.100 184.200 462.300 185.400 ;
        RECT 455.100 181.050 456.900 182.850 ;
        RECT 454.950 178.950 457.050 181.050 ;
        RECT 436.950 172.950 439.050 178.050 ;
        RECT 458.100 173.700 459.300 184.200 ;
        RECT 460.500 183.600 462.300 184.200 ;
        RECT 464.100 184.200 468.300 185.400 ;
        RECT 464.100 173.700 465.300 184.200 ;
        RECT 466.500 183.600 468.300 184.200 ;
        RECT 470.100 184.200 474.300 185.400 ;
        RECT 470.100 173.700 471.300 184.200 ;
        RECT 472.500 183.600 474.300 184.200 ;
        RECT 475.200 181.050 476.100 186.300 ;
        RECT 497.400 181.050 498.600 186.300 ;
        RECT 515.400 186.300 519.600 187.200 ;
        RECT 524.550 188.400 526.350 194.400 ;
        RECT 532.650 191.400 534.450 194.400 ;
        RECT 540.450 191.400 542.250 194.400 ;
        RECT 548.250 192.300 550.050 194.400 ;
        RECT 548.250 191.400 552.000 192.300 ;
        RECT 532.650 190.500 533.700 191.400 ;
        RECT 529.950 189.300 533.700 190.500 ;
        RECT 541.200 190.500 542.250 191.400 ;
        RECT 550.950 190.500 552.000 191.400 ;
        RECT 541.200 189.450 546.150 190.500 ;
        RECT 529.950 188.400 532.050 189.300 ;
        RECT 544.350 188.700 546.150 189.450 ;
        RECT 505.950 181.950 508.050 184.050 ;
        RECT 475.200 178.950 478.050 181.050 ;
        RECT 475.200 173.700 476.100 178.950 ;
        RECT 494.100 178.050 495.900 179.850 ;
        RECT 496.950 178.950 499.050 181.050 ;
        RECT 493.950 175.950 496.050 178.050 ;
        RECT 437.400 165.600 438.600 172.950 ;
        RECT 455.400 172.500 459.300 173.700 ;
        RECT 461.400 172.500 465.300 173.700 ;
        RECT 467.400 172.500 471.300 173.700 ;
        RECT 473.400 172.500 476.100 173.700 ;
        RECT 416.400 159.600 418.200 165.600 ;
        RECT 437.400 159.600 439.200 165.600 ;
        RECT 455.400 159.600 457.200 172.500 ;
        RECT 461.400 159.600 463.200 172.500 ;
        RECT 467.400 159.600 469.200 172.500 ;
        RECT 473.400 159.600 475.200 172.500 ;
        RECT 497.400 165.600 498.600 178.950 ;
        RECT 500.100 178.050 501.900 179.850 ;
        RECT 499.950 175.950 502.050 178.050 ;
        RECT 506.550 166.050 507.450 181.950 ;
        RECT 515.400 181.050 516.600 186.300 ;
        RECT 524.550 181.050 525.750 188.400 ;
        RECT 547.650 187.800 549.450 189.600 ;
        RECT 550.950 188.400 553.050 190.500 ;
        RECT 556.050 188.400 557.850 194.400 ;
        RECT 571.800 191.400 573.600 194.400 ;
        RECT 537.150 186.000 538.950 186.600 ;
        RECT 548.100 186.000 549.150 187.800 ;
        RECT 537.150 184.800 549.150 186.000 ;
        RECT 512.100 178.050 513.900 179.850 ;
        RECT 514.950 178.950 517.050 181.050 ;
        RECT 511.950 175.950 514.050 178.050 ;
        RECT 496.800 159.600 498.600 165.600 ;
        RECT 505.950 163.950 508.050 166.050 ;
        RECT 515.400 165.600 516.600 178.950 ;
        RECT 518.100 178.050 519.900 179.850 ;
        RECT 524.550 179.250 530.850 181.050 ;
        RECT 524.550 178.950 529.050 179.250 ;
        RECT 517.950 175.950 520.050 178.050 ;
        RECT 524.550 171.600 525.750 178.950 ;
        RECT 526.950 173.400 528.750 175.200 ;
        RECT 527.850 172.200 532.050 173.400 ;
        RECT 537.150 172.200 538.050 184.800 ;
        RECT 548.100 183.600 555.000 184.800 ;
        RECT 548.100 183.000 549.900 183.600 ;
        RECT 554.100 182.850 555.000 183.600 ;
        RECT 551.100 181.800 552.900 182.400 ;
        RECT 544.950 180.600 552.900 181.800 ;
        RECT 554.100 181.050 555.900 182.850 ;
        RECT 544.950 178.950 547.050 180.600 ;
        RECT 553.950 178.950 556.050 181.050 ;
        RECT 546.750 173.700 548.550 174.000 ;
        RECT 556.950 173.700 557.850 188.400 ;
        RECT 572.400 178.050 573.600 191.400 ;
        RECT 593.700 189.600 595.500 194.400 ;
        RECT 616.800 191.400 618.600 194.400 ;
        RECT 590.400 188.400 595.500 189.600 ;
        RECT 590.400 181.050 591.600 188.400 ;
        RECT 613.950 181.950 616.050 184.050 ;
        RECT 574.950 178.950 577.050 181.050 ;
        RECT 589.950 178.950 592.050 181.050 ;
        RECT 546.750 173.100 557.850 173.700 ;
        RECT 515.400 159.600 517.200 165.600 ;
        RECT 524.550 159.600 526.350 171.600 ;
        RECT 529.950 171.300 532.050 172.200 ;
        RECT 532.950 171.300 538.050 172.200 ;
        RECT 540.150 172.500 557.850 173.100 ;
        RECT 571.950 172.950 574.050 178.050 ;
        RECT 575.100 177.150 576.900 178.950 ;
        RECT 540.150 172.200 548.550 172.500 ;
        RECT 532.950 170.400 533.850 171.300 ;
        RECT 531.150 168.600 533.850 170.400 ;
        RECT 534.750 170.100 536.550 170.400 ;
        RECT 540.150 170.100 541.050 172.200 ;
        RECT 556.950 171.600 557.850 172.500 ;
        RECT 534.750 169.200 541.050 170.100 ;
        RECT 541.950 170.700 543.750 171.300 ;
        RECT 541.950 169.500 549.450 170.700 ;
        RECT 534.750 168.600 536.550 169.200 ;
        RECT 548.250 168.600 549.450 169.500 ;
        RECT 529.950 165.600 533.850 167.700 ;
        RECT 538.950 167.550 540.750 168.300 ;
        RECT 543.750 167.550 545.550 168.300 ;
        RECT 538.950 166.500 545.550 167.550 ;
        RECT 548.250 166.500 553.050 168.600 ;
        RECT 532.050 159.600 533.850 165.600 ;
        RECT 539.850 159.600 541.650 166.500 ;
        RECT 548.250 165.600 549.450 166.500 ;
        RECT 547.650 159.600 549.450 165.600 ;
        RECT 556.050 159.600 557.850 171.600 ;
        RECT 572.400 165.600 573.600 172.950 ;
        RECT 590.400 171.600 591.600 178.950 ;
        RECT 593.100 178.050 594.900 179.850 ;
        RECT 595.950 178.950 598.050 181.050 ;
        RECT 614.100 180.150 615.900 181.950 ;
        RECT 617.400 181.050 618.300 191.400 ;
        RECT 636.300 190.200 638.100 194.400 ;
        RECT 635.400 188.400 638.100 190.200 ;
        RECT 619.950 181.950 622.050 184.050 ;
        RECT 592.950 175.950 595.050 178.050 ;
        RECT 596.100 177.150 597.900 178.950 ;
        RECT 599.100 178.050 600.900 179.850 ;
        RECT 616.950 178.950 619.050 181.050 ;
        RECT 620.100 180.150 621.900 181.950 ;
        RECT 635.400 181.050 636.300 188.400 ;
        RECT 638.100 186.600 639.900 187.500 ;
        RECT 643.800 186.600 645.600 194.400 ;
        RECT 661.500 189.600 663.300 194.400 ;
        RECT 683.400 191.400 685.200 194.400 ;
        RECT 706.800 191.400 708.600 194.400 ;
        RECT 661.500 188.400 666.600 189.600 ;
        RECT 638.100 185.700 645.600 186.600 ;
        RECT 634.950 178.950 637.050 181.050 ;
        RECT 637.950 178.950 640.050 181.050 ;
        RECT 598.950 175.950 601.050 178.050 ;
        RECT 617.400 171.600 618.300 178.950 ;
        RECT 623.100 175.950 625.200 178.050 ;
        RECT 571.800 159.600 573.600 165.600 ;
        RECT 589.800 159.600 591.600 171.600 ;
        RECT 592.800 170.700 600.600 171.600 ;
        RECT 592.800 159.600 594.600 170.700 ;
        RECT 598.800 159.600 600.600 170.700 ;
        RECT 614.700 170.400 618.300 171.600 ;
        RECT 614.700 159.600 616.500 170.400 ;
        RECT 623.550 166.050 624.450 175.950 ;
        RECT 635.400 171.600 636.300 178.950 ;
        RECT 638.100 177.150 639.900 178.950 ;
        RECT 622.950 163.950 625.050 166.050 ;
        RECT 634.500 159.600 636.300 171.600 ;
        RECT 641.700 165.600 642.600 185.700 ;
        RECT 644.100 181.050 645.900 182.850 ;
        RECT 665.400 181.050 666.600 188.400 ;
        RECT 679.950 181.950 682.050 184.050 ;
        RECT 643.950 178.950 646.050 181.050 ;
        RECT 656.100 178.050 657.900 179.850 ;
        RECT 658.950 178.950 661.050 181.050 ;
        RECT 655.950 175.950 658.050 178.050 ;
        RECT 659.100 177.150 660.900 178.950 ;
        RECT 662.100 178.050 663.900 179.850 ;
        RECT 664.950 178.950 667.050 181.050 ;
        RECT 680.100 180.150 681.900 181.950 ;
        RECT 683.700 181.050 684.600 191.400 ;
        RECT 685.950 181.950 688.050 184.050 ;
        RECT 703.950 181.950 706.050 184.050 ;
        RECT 682.950 178.950 685.050 181.050 ;
        RECT 686.100 180.150 687.900 181.950 ;
        RECT 704.100 180.150 705.900 181.950 ;
        RECT 707.400 181.050 708.300 191.400 ;
        RECT 722.400 186.600 724.200 194.400 ;
        RECT 729.900 190.200 731.700 194.400 ;
        RECT 748.800 191.400 750.600 194.400 ;
        RECT 729.900 188.400 732.600 190.200 ;
        RECT 728.100 186.600 729.900 187.500 ;
        RECT 722.400 185.700 729.900 186.600 ;
        RECT 709.950 181.950 712.050 184.050 ;
        RECT 706.950 178.950 709.050 181.050 ;
        RECT 710.100 180.150 711.900 181.950 ;
        RECT 722.100 181.050 723.900 182.850 ;
        RECT 721.950 178.950 724.050 181.050 ;
        RECT 661.950 175.950 664.050 178.050 ;
        RECT 665.400 171.600 666.600 178.950 ;
        RECT 683.700 171.600 684.600 178.950 ;
        RECT 707.400 171.600 708.300 178.950 ;
        RECT 640.800 159.600 642.600 165.600 ;
        RECT 656.400 170.700 664.200 171.600 ;
        RECT 656.400 159.600 658.200 170.700 ;
        RECT 662.400 159.600 664.200 170.700 ;
        RECT 665.400 159.600 667.200 171.600 ;
        RECT 683.700 170.400 687.300 171.600 ;
        RECT 685.500 159.600 687.300 170.400 ;
        RECT 704.700 170.400 708.300 171.600 ;
        RECT 704.700 159.600 706.500 170.400 ;
        RECT 725.400 165.600 726.300 185.700 ;
        RECT 731.700 181.050 732.600 188.400 ;
        RECT 727.950 178.950 730.050 181.050 ;
        RECT 730.950 178.950 733.050 181.050 ;
        RECT 728.100 177.150 729.900 178.950 ;
        RECT 731.700 171.600 732.600 178.950 ;
        RECT 749.400 178.050 750.600 191.400 ;
        RECT 766.800 188.400 768.600 194.400 ;
        RECT 767.400 186.300 768.600 188.400 ;
        RECT 769.800 189.300 771.600 194.400 ;
        RECT 775.800 189.300 777.600 194.400 ;
        RECT 791.400 191.400 793.200 194.400 ;
        RECT 769.800 187.950 777.600 189.300 ;
        RECT 781.950 187.950 784.050 190.050 ;
        RECT 767.400 185.250 771.150 186.300 ;
        RECT 769.950 181.050 771.150 185.250 ;
        RECT 751.950 178.950 754.050 181.050 ;
        RECT 748.950 172.950 751.050 178.050 ;
        RECT 752.100 177.150 753.900 178.950 ;
        RECT 767.100 178.050 768.900 179.850 ;
        RECT 769.950 178.950 772.050 181.050 ;
        RECT 766.950 175.950 769.050 178.050 ;
        RECT 725.400 159.600 727.200 165.600 ;
        RECT 731.700 159.600 733.500 171.600 ;
        RECT 749.400 165.600 750.600 172.950 ;
        RECT 770.850 165.600 772.050 178.950 ;
        RECT 773.100 178.050 774.900 179.850 ;
        RECT 775.950 178.950 778.050 181.050 ;
        RECT 772.950 175.950 775.050 178.050 ;
        RECT 776.100 177.150 777.900 178.950 ;
        RECT 782.550 169.050 783.450 187.950 ;
        RECT 787.950 181.950 790.050 184.050 ;
        RECT 788.100 180.150 789.900 181.950 ;
        RECT 791.700 181.050 792.600 191.400 ;
        RECT 814.200 186.000 816.000 194.400 ;
        RECT 812.700 184.800 816.000 186.000 ;
        RECT 836.400 191.400 838.200 194.400 ;
        RECT 854.400 191.400 856.200 194.400 ;
        RECT 874.800 191.400 876.600 194.400 ;
        RECT 892.800 191.400 894.600 194.400 ;
        RECT 793.950 181.950 796.050 184.050 ;
        RECT 790.950 178.950 793.050 181.050 ;
        RECT 794.100 180.150 795.900 181.950 ;
        RECT 812.700 181.050 813.600 184.800 ;
        RECT 811.950 178.950 814.050 181.050 ;
        RECT 791.700 171.600 792.600 178.950 ;
        RECT 791.700 170.400 795.300 171.600 ;
        RECT 781.950 166.950 784.050 169.050 ;
        RECT 748.800 159.600 750.600 165.600 ;
        RECT 770.400 159.600 772.200 165.600 ;
        RECT 793.500 159.600 795.300 170.400 ;
        RECT 812.700 166.800 813.600 178.950 ;
        RECT 815.100 178.050 816.900 179.850 ;
        RECT 817.950 178.950 820.050 181.050 ;
        RECT 814.950 175.950 817.050 178.050 ;
        RECT 818.100 177.150 819.900 178.950 ;
        RECT 821.100 178.050 822.900 179.850 ;
        RECT 832.950 178.950 835.050 181.050 ;
        RECT 820.950 175.950 823.050 178.050 ;
        RECT 833.100 177.150 834.900 178.950 ;
        RECT 836.400 178.050 837.600 191.400 ;
        RECT 850.950 178.950 853.050 181.050 ;
        RECT 835.950 172.950 838.050 178.050 ;
        RECT 851.100 177.150 852.900 178.950 ;
        RECT 854.400 178.050 855.600 191.400 ;
        RECT 871.950 181.950 874.050 184.050 ;
        RECT 872.100 180.150 873.900 181.950 ;
        RECT 875.400 181.050 876.300 191.400 ;
        RECT 877.950 181.950 880.050 184.050 ;
        RECT 874.950 178.950 877.050 181.050 ;
        RECT 878.100 180.150 879.900 181.950 ;
        RECT 853.950 172.950 856.050 178.050 ;
        RECT 812.700 165.900 819.300 166.800 ;
        RECT 812.700 165.600 813.600 165.900 ;
        RECT 811.800 159.600 813.600 165.600 ;
        RECT 817.800 165.600 819.300 165.900 ;
        RECT 836.400 165.600 837.600 172.950 ;
        RECT 854.400 165.600 855.600 172.950 ;
        RECT 875.400 171.600 876.300 178.950 ;
        RECT 893.400 178.050 894.600 191.400 ;
        RECT 895.950 178.950 898.050 181.050 ;
        RECT 892.950 172.950 895.050 178.050 ;
        RECT 896.100 177.150 897.900 178.950 ;
        RECT 872.700 170.400 876.300 171.600 ;
        RECT 817.800 159.600 819.600 165.600 ;
        RECT 836.400 159.600 838.200 165.600 ;
        RECT 854.400 159.600 856.200 165.600 ;
        RECT 872.700 159.600 874.500 170.400 ;
        RECT 893.400 165.600 894.600 172.950 ;
        RECT 892.800 159.600 894.600 165.600 ;
        RECT 13.800 143.400 15.600 155.400 ;
        RECT 16.800 144.300 18.600 155.400 ;
        RECT 22.800 144.300 24.600 155.400 ;
        RECT 16.800 143.400 24.600 144.300 ;
        RECT 38.400 149.400 40.200 155.400 ;
        RECT 46.950 151.950 49.050 154.050 ;
        RECT 14.400 136.050 15.600 143.400 ;
        RECT 16.950 136.950 19.050 139.050 ;
        RECT 13.950 133.950 16.050 136.050 ;
        RECT 17.100 135.150 18.900 136.950 ;
        RECT 20.100 136.050 21.900 137.850 ;
        RECT 22.950 136.950 25.050 139.050 ;
        RECT 34.950 136.950 37.050 139.050 ;
        RECT 19.950 133.950 22.050 136.050 ;
        RECT 23.100 135.150 24.900 136.950 ;
        RECT 35.100 135.150 36.900 136.950 ;
        RECT 38.400 136.050 39.600 149.400 ;
        RECT 40.950 136.950 43.050 139.050 ;
        RECT 37.950 133.950 40.050 136.050 ;
        RECT 41.100 135.150 42.900 136.950 ;
        RECT 14.400 126.600 15.600 133.950 ;
        RECT 38.400 128.700 39.600 133.950 ;
        RECT 47.550 133.050 48.450 151.950 ;
        RECT 59.400 149.400 61.200 155.400 ;
        RECT 59.700 149.100 61.200 149.400 ;
        RECT 65.400 149.400 67.200 155.400 ;
        RECT 65.400 149.100 66.300 149.400 ;
        RECT 59.700 148.200 66.300 149.100 ;
        RECT 50.100 145.950 52.200 148.050 ;
        RECT 46.950 130.950 49.050 133.050 ;
        RECT 38.400 127.800 42.600 128.700 ;
        RECT 14.400 125.400 19.500 126.600 ;
        RECT 17.700 120.600 19.500 125.400 ;
        RECT 40.800 120.600 42.600 127.800 ;
        RECT 50.550 127.050 51.450 145.950 ;
        RECT 55.950 136.950 58.050 139.050 ;
        RECT 56.100 135.150 57.900 136.950 ;
        RECT 59.100 136.050 60.900 137.850 ;
        RECT 61.950 136.950 64.050 139.050 ;
        RECT 58.950 133.950 61.050 136.050 ;
        RECT 62.100 135.150 63.900 136.950 ;
        RECT 65.400 136.050 66.300 148.200 ;
        RECT 73.950 145.950 76.050 148.050 ;
        RECT 64.950 133.950 67.050 136.050 ;
        RECT 65.400 130.200 66.300 133.950 ;
        RECT 74.550 133.050 75.450 145.950 ;
        RECT 80.400 144.300 82.200 155.400 ;
        RECT 86.400 144.300 88.200 155.400 ;
        RECT 80.400 143.400 88.200 144.300 ;
        RECT 89.400 143.400 91.200 155.400 ;
        RECT 94.950 148.950 97.050 151.050 ;
        RECT 107.400 149.400 109.200 155.400 ;
        RECT 79.950 136.950 82.050 139.050 ;
        RECT 80.100 135.150 81.900 136.950 ;
        RECT 83.100 136.050 84.900 137.850 ;
        RECT 85.950 136.950 88.050 139.050 ;
        RECT 82.950 133.950 85.050 136.050 ;
        RECT 86.100 135.150 87.900 136.950 ;
        RECT 89.400 136.050 90.600 143.400 ;
        RECT 88.950 133.950 91.050 136.050 ;
        RECT 73.950 130.950 76.050 133.050 ;
        RECT 63.000 129.000 66.300 130.200 ;
        RECT 49.950 124.950 52.050 127.050 ;
        RECT 63.000 120.600 64.800 129.000 ;
        RECT 89.400 126.600 90.600 133.950 ;
        RECT 85.500 125.400 90.600 126.600 ;
        RECT 85.500 120.600 87.300 125.400 ;
        RECT 95.550 124.050 96.450 148.950 ;
        RECT 103.950 133.950 106.050 136.050 ;
        RECT 104.100 132.150 105.900 133.950 ;
        RECT 107.400 129.300 108.300 149.400 ;
        RECT 113.700 143.400 115.500 155.400 ;
        RECT 124.950 151.950 127.050 154.050 ;
        RECT 110.100 136.050 111.900 137.850 ;
        RECT 113.700 136.050 114.600 143.400 ;
        RECT 125.550 139.050 126.450 151.950 ;
        RECT 133.500 144.600 135.300 155.400 ;
        RECT 131.700 143.400 135.300 144.600 ;
        RECT 152.700 144.600 154.500 155.400 ;
        RECT 173.400 149.400 175.200 155.400 ;
        RECT 193.800 149.400 195.600 155.400 ;
        RECT 217.800 149.400 219.600 155.400 ;
        RECT 152.700 143.400 156.300 144.600 ;
        RECT 124.950 136.950 127.050 139.050 ;
        RECT 131.700 136.050 132.600 143.400 ;
        RECT 155.400 136.050 156.300 143.400 ;
        RECT 173.400 142.050 174.600 149.400 ;
        RECT 170.100 136.050 171.900 137.850 ;
        RECT 172.950 136.950 175.050 142.050 ;
        RECT 109.950 133.950 112.050 136.050 ;
        RECT 112.950 133.950 115.050 136.050 ;
        RECT 104.400 128.400 111.900 129.300 ;
        RECT 94.950 121.950 97.050 124.050 ;
        RECT 104.400 120.600 106.200 128.400 ;
        RECT 110.100 127.500 111.900 128.400 ;
        RECT 113.700 126.600 114.600 133.950 ;
        RECT 128.100 133.050 129.900 134.850 ;
        RECT 130.950 133.950 133.050 136.050 ;
        RECT 127.950 130.950 130.050 133.050 ;
        RECT 111.900 124.800 114.600 126.600 ;
        RECT 111.900 120.600 113.700 124.800 ;
        RECT 131.700 123.600 132.600 133.950 ;
        RECT 134.100 133.050 135.900 134.850 ;
        RECT 152.100 133.050 153.900 134.850 ;
        RECT 154.950 133.950 157.050 136.050 ;
        RECT 133.950 130.950 136.050 133.050 ;
        RECT 151.950 130.950 154.050 133.050 ;
        RECT 155.400 123.600 156.300 133.950 ;
        RECT 158.100 133.050 159.900 134.850 ;
        RECT 169.950 133.950 172.050 136.050 ;
        RECT 157.950 130.950 160.050 133.050 ;
        RECT 173.400 123.600 174.600 136.950 ;
        RECT 188.100 136.050 189.900 137.850 ;
        RECT 190.950 136.950 193.050 139.050 ;
        RECT 187.950 133.950 190.050 136.050 ;
        RECT 191.100 135.150 192.900 136.950 ;
        RECT 193.950 136.050 195.150 149.400 ;
        RECT 196.950 136.950 199.050 139.050 ;
        RECT 193.950 133.950 196.050 136.050 ;
        RECT 197.100 135.150 198.900 136.950 ;
        RECT 212.100 136.050 213.900 137.850 ;
        RECT 214.950 136.950 217.050 139.050 ;
        RECT 211.950 133.950 214.050 136.050 ;
        RECT 215.100 135.150 216.900 136.950 ;
        RECT 217.950 136.050 219.150 149.400 ;
        RECT 228.150 143.400 229.950 155.400 ;
        RECT 236.550 149.400 238.350 155.400 ;
        RECT 236.550 148.500 237.750 149.400 ;
        RECT 244.350 148.500 246.150 155.400 ;
        RECT 252.150 149.400 253.950 155.400 ;
        RECT 232.950 146.400 237.750 148.500 ;
        RECT 240.450 147.450 247.050 148.500 ;
        RECT 240.450 146.700 242.250 147.450 ;
        RECT 245.250 146.700 247.050 147.450 ;
        RECT 252.150 147.300 256.050 149.400 ;
        RECT 236.550 145.500 237.750 146.400 ;
        RECT 249.450 145.800 251.250 146.400 ;
        RECT 236.550 144.300 244.050 145.500 ;
        RECT 242.250 143.700 244.050 144.300 ;
        RECT 244.950 144.900 251.250 145.800 ;
        RECT 228.150 142.500 229.050 143.400 ;
        RECT 244.950 142.800 245.850 144.900 ;
        RECT 249.450 144.600 251.250 144.900 ;
        RECT 252.150 144.600 254.850 146.400 ;
        RECT 252.150 143.700 253.050 144.600 ;
        RECT 237.450 142.500 245.850 142.800 ;
        RECT 228.150 141.900 245.850 142.500 ;
        RECT 247.950 142.800 253.050 143.700 ;
        RECT 253.950 142.800 256.050 143.700 ;
        RECT 259.650 143.400 261.450 155.400 ;
        RECT 228.150 141.300 239.250 141.900 ;
        RECT 220.950 136.950 223.050 139.050 ;
        RECT 217.950 133.950 220.050 136.050 ;
        RECT 221.100 135.150 222.900 136.950 ;
        RECT 194.850 129.750 196.050 133.950 ;
        RECT 218.850 129.750 220.050 133.950 ;
        RECT 194.850 128.700 198.600 129.750 ;
        RECT 218.850 128.700 222.600 129.750 ;
        RECT 188.400 125.700 196.200 127.050 ;
        RECT 131.400 120.600 133.200 123.600 ;
        RECT 154.800 120.600 156.600 123.600 ;
        RECT 173.400 120.600 175.200 123.600 ;
        RECT 188.400 120.600 190.200 125.700 ;
        RECT 194.400 120.600 196.200 125.700 ;
        RECT 197.400 126.600 198.600 128.700 ;
        RECT 197.400 120.600 199.200 126.600 ;
        RECT 212.400 125.700 220.200 127.050 ;
        RECT 212.400 120.600 214.200 125.700 ;
        RECT 218.400 120.600 220.200 125.700 ;
        RECT 221.400 126.600 222.600 128.700 ;
        RECT 228.150 126.600 229.050 141.300 ;
        RECT 237.450 141.000 239.250 141.300 ;
        RECT 229.950 133.950 232.050 136.050 ;
        RECT 238.950 134.400 241.050 136.050 ;
        RECT 230.100 132.150 231.900 133.950 ;
        RECT 233.100 133.200 241.050 134.400 ;
        RECT 233.100 132.600 234.900 133.200 ;
        RECT 231.000 131.400 231.900 132.150 ;
        RECT 236.100 131.400 237.900 132.000 ;
        RECT 231.000 130.200 237.900 131.400 ;
        RECT 247.950 130.200 248.850 142.800 ;
        RECT 253.950 141.600 258.150 142.800 ;
        RECT 257.250 139.800 259.050 141.600 ;
        RECT 260.250 136.050 261.450 143.400 ;
        RECT 256.950 135.750 261.450 136.050 ;
        RECT 255.150 133.950 261.450 135.750 ;
        RECT 236.850 129.000 248.850 130.200 ;
        RECT 236.850 127.200 237.900 129.000 ;
        RECT 247.050 128.400 248.850 129.000 ;
        RECT 221.400 120.600 223.200 126.600 ;
        RECT 228.150 120.600 229.950 126.600 ;
        RECT 232.950 124.500 235.050 126.600 ;
        RECT 236.550 125.400 238.350 127.200 ;
        RECT 260.250 126.600 261.450 133.950 ;
        RECT 239.850 125.550 241.650 126.300 ;
        RECT 253.950 125.700 256.050 126.600 ;
        RECT 239.850 124.500 244.800 125.550 ;
        RECT 234.000 123.600 235.050 124.500 ;
        RECT 243.750 123.600 244.800 124.500 ;
        RECT 252.300 124.500 256.050 125.700 ;
        RECT 252.300 123.600 253.350 124.500 ;
        RECT 234.000 122.700 237.750 123.600 ;
        RECT 235.950 120.600 237.750 122.700 ;
        RECT 243.750 120.600 245.550 123.600 ;
        RECT 251.550 120.600 253.350 123.600 ;
        RECT 259.650 120.600 261.450 126.600 ;
        RECT 264.150 143.400 265.950 155.400 ;
        RECT 272.550 149.400 274.350 155.400 ;
        RECT 272.550 148.500 273.750 149.400 ;
        RECT 280.350 148.500 282.150 155.400 ;
        RECT 288.150 149.400 289.950 155.400 ;
        RECT 268.950 146.400 273.750 148.500 ;
        RECT 276.450 147.450 283.050 148.500 ;
        RECT 276.450 146.700 278.250 147.450 ;
        RECT 281.250 146.700 283.050 147.450 ;
        RECT 288.150 147.300 292.050 149.400 ;
        RECT 272.550 145.500 273.750 146.400 ;
        RECT 285.450 145.800 287.250 146.400 ;
        RECT 272.550 144.300 280.050 145.500 ;
        RECT 278.250 143.700 280.050 144.300 ;
        RECT 280.950 144.900 287.250 145.800 ;
        RECT 264.150 142.500 265.050 143.400 ;
        RECT 280.950 142.800 281.850 144.900 ;
        RECT 285.450 144.600 287.250 144.900 ;
        RECT 288.150 144.600 290.850 146.400 ;
        RECT 288.150 143.700 289.050 144.600 ;
        RECT 273.450 142.500 281.850 142.800 ;
        RECT 264.150 141.900 281.850 142.500 ;
        RECT 283.950 142.800 289.050 143.700 ;
        RECT 289.950 142.800 292.050 143.700 ;
        RECT 295.650 143.400 297.450 155.400 ;
        RECT 264.150 141.300 275.250 141.900 ;
        RECT 264.150 126.600 265.050 141.300 ;
        RECT 273.450 141.000 275.250 141.300 ;
        RECT 265.950 133.950 268.050 136.050 ;
        RECT 274.950 134.400 277.050 136.050 ;
        RECT 266.100 132.150 267.900 133.950 ;
        RECT 269.100 133.200 277.050 134.400 ;
        RECT 269.100 132.600 270.900 133.200 ;
        RECT 267.000 131.400 267.900 132.150 ;
        RECT 272.100 131.400 273.900 132.000 ;
        RECT 267.000 130.200 273.900 131.400 ;
        RECT 283.950 130.200 284.850 142.800 ;
        RECT 289.950 141.600 294.150 142.800 ;
        RECT 293.250 139.800 295.050 141.600 ;
        RECT 296.250 136.050 297.450 143.400 ;
        RECT 292.950 135.750 297.450 136.050 ;
        RECT 291.150 133.950 297.450 135.750 ;
        RECT 272.850 129.000 284.850 130.200 ;
        RECT 272.850 127.200 273.900 129.000 ;
        RECT 283.050 128.400 284.850 129.000 ;
        RECT 264.150 120.600 265.950 126.600 ;
        RECT 268.950 124.500 271.050 126.600 ;
        RECT 272.550 125.400 274.350 127.200 ;
        RECT 296.250 126.600 297.450 133.950 ;
        RECT 275.850 125.550 277.650 126.300 ;
        RECT 289.950 125.700 292.050 126.600 ;
        RECT 275.850 124.500 280.800 125.550 ;
        RECT 270.000 123.600 271.050 124.500 ;
        RECT 279.750 123.600 280.800 124.500 ;
        RECT 288.300 124.500 292.050 125.700 ;
        RECT 288.300 123.600 289.350 124.500 ;
        RECT 270.000 122.700 273.750 123.600 ;
        RECT 271.950 120.600 273.750 122.700 ;
        RECT 279.750 120.600 281.550 123.600 ;
        RECT 287.550 120.600 289.350 123.600 ;
        RECT 295.650 120.600 297.450 126.600 ;
        RECT 300.150 143.400 301.950 155.400 ;
        RECT 308.550 149.400 310.350 155.400 ;
        RECT 308.550 148.500 309.750 149.400 ;
        RECT 316.350 148.500 318.150 155.400 ;
        RECT 324.150 149.400 325.950 155.400 ;
        RECT 304.950 146.400 309.750 148.500 ;
        RECT 312.450 147.450 319.050 148.500 ;
        RECT 312.450 146.700 314.250 147.450 ;
        RECT 317.250 146.700 319.050 147.450 ;
        RECT 324.150 147.300 328.050 149.400 ;
        RECT 308.550 145.500 309.750 146.400 ;
        RECT 321.450 145.800 323.250 146.400 ;
        RECT 308.550 144.300 316.050 145.500 ;
        RECT 314.250 143.700 316.050 144.300 ;
        RECT 316.950 144.900 323.250 145.800 ;
        RECT 300.150 142.500 301.050 143.400 ;
        RECT 316.950 142.800 317.850 144.900 ;
        RECT 321.450 144.600 323.250 144.900 ;
        RECT 324.150 144.600 326.850 146.400 ;
        RECT 324.150 143.700 325.050 144.600 ;
        RECT 309.450 142.500 317.850 142.800 ;
        RECT 300.150 141.900 317.850 142.500 ;
        RECT 319.950 142.800 325.050 143.700 ;
        RECT 325.950 142.800 328.050 143.700 ;
        RECT 331.650 143.400 333.450 155.400 ;
        RECT 350.400 149.400 352.200 155.400 ;
        RECT 371.400 149.400 373.200 155.400 ;
        RECT 388.800 149.400 390.600 155.400 ;
        RECT 300.150 141.300 311.250 141.900 ;
        RECT 300.150 126.600 301.050 141.300 ;
        RECT 309.450 141.000 311.250 141.300 ;
        RECT 301.950 133.950 304.050 136.050 ;
        RECT 310.950 134.400 313.050 136.050 ;
        RECT 302.100 132.150 303.900 133.950 ;
        RECT 305.100 133.200 313.050 134.400 ;
        RECT 305.100 132.600 306.900 133.200 ;
        RECT 303.000 131.400 303.900 132.150 ;
        RECT 308.100 131.400 309.900 132.000 ;
        RECT 303.000 130.200 309.900 131.400 ;
        RECT 319.950 130.200 320.850 142.800 ;
        RECT 325.950 141.600 330.150 142.800 ;
        RECT 329.250 139.800 331.050 141.600 ;
        RECT 332.250 136.050 333.450 143.400 ;
        RECT 346.950 136.950 349.050 139.050 ;
        RECT 328.950 135.750 333.450 136.050 ;
        RECT 327.150 133.950 333.450 135.750 ;
        RECT 347.100 135.150 348.900 136.950 ;
        RECT 350.850 136.050 352.050 149.400 ;
        RECT 371.400 142.050 372.600 149.400 ;
        RECT 389.400 142.050 390.600 149.400 ;
        RECT 407.700 144.600 409.500 155.400 ;
        RECT 430.500 144.600 432.300 155.400 ;
        RECT 439.950 145.950 442.050 148.050 ;
        RECT 407.700 143.400 411.300 144.600 ;
        RECT 352.950 136.950 355.050 139.050 ;
        RECT 308.850 129.000 320.850 130.200 ;
        RECT 308.850 127.200 309.900 129.000 ;
        RECT 319.050 128.400 320.850 129.000 ;
        RECT 300.150 120.600 301.950 126.600 ;
        RECT 304.950 124.500 307.050 126.600 ;
        RECT 308.550 125.400 310.350 127.200 ;
        RECT 332.250 126.600 333.450 133.950 ;
        RECT 349.950 133.950 352.050 136.050 ;
        RECT 353.100 135.150 354.900 136.950 ;
        RECT 356.100 136.050 357.900 137.850 ;
        RECT 368.100 136.050 369.900 137.850 ;
        RECT 370.950 136.950 373.050 142.050 ;
        RECT 388.950 136.950 391.050 142.050 ;
        RECT 355.950 133.950 358.050 136.050 ;
        RECT 367.950 133.950 370.050 136.050 ;
        RECT 349.950 129.750 351.150 133.950 ;
        RECT 347.400 128.700 351.150 129.750 ;
        RECT 347.400 126.600 348.600 128.700 ;
        RECT 311.850 125.550 313.650 126.300 ;
        RECT 325.950 125.700 328.050 126.600 ;
        RECT 311.850 124.500 316.800 125.550 ;
        RECT 306.000 123.600 307.050 124.500 ;
        RECT 315.750 123.600 316.800 124.500 ;
        RECT 324.300 124.500 328.050 125.700 ;
        RECT 324.300 123.600 325.350 124.500 ;
        RECT 306.000 122.700 309.750 123.600 ;
        RECT 307.950 120.600 309.750 122.700 ;
        RECT 315.750 120.600 317.550 123.600 ;
        RECT 323.550 120.600 325.350 123.600 ;
        RECT 331.650 120.600 333.450 126.600 ;
        RECT 346.800 120.600 348.600 126.600 ;
        RECT 349.800 125.700 357.600 127.050 ;
        RECT 349.800 120.600 351.600 125.700 ;
        RECT 355.800 120.600 357.600 125.700 ;
        RECT 371.400 123.600 372.600 136.950 ;
        RECT 389.400 123.600 390.600 136.950 ;
        RECT 392.100 136.050 393.900 137.850 ;
        RECT 410.400 136.050 411.300 143.400 ;
        RECT 428.700 143.400 432.300 144.600 ;
        RECT 428.700 136.050 429.600 143.400 ;
        RECT 436.950 142.950 439.050 145.050 ;
        RECT 391.950 133.950 394.050 136.050 ;
        RECT 407.100 133.050 408.900 134.850 ;
        RECT 409.950 133.950 412.050 136.050 ;
        RECT 406.950 130.950 409.050 133.050 ;
        RECT 410.400 123.600 411.300 133.950 ;
        RECT 413.100 133.050 414.900 134.850 ;
        RECT 425.100 133.050 426.900 134.850 ;
        RECT 427.950 133.950 430.050 136.050 ;
        RECT 412.950 130.950 415.050 133.050 ;
        RECT 424.950 130.950 427.050 133.050 ;
        RECT 428.700 123.600 429.600 133.950 ;
        RECT 431.100 133.050 432.900 134.850 ;
        RECT 430.950 130.950 433.050 133.050 ;
        RECT 437.550 127.050 438.450 142.950 ;
        RECT 440.550 139.050 441.450 145.950 ;
        RECT 446.400 144.300 448.200 155.400 ;
        RECT 452.400 144.300 454.200 155.400 ;
        RECT 446.400 143.400 454.200 144.300 ;
        RECT 455.400 143.400 457.200 155.400 ;
        RECT 466.950 148.950 469.050 151.050 ;
        RECT 476.400 149.400 478.200 155.400 ;
        RECT 439.950 136.950 442.050 139.050 ;
        RECT 445.950 136.950 448.050 139.050 ;
        RECT 446.100 135.150 447.900 136.950 ;
        RECT 449.100 136.050 450.900 137.850 ;
        RECT 451.950 136.950 454.050 139.050 ;
        RECT 448.950 133.950 451.050 136.050 ;
        RECT 452.100 135.150 453.900 136.950 ;
        RECT 455.400 136.050 456.600 143.400 ;
        RECT 454.950 133.950 457.050 136.050 ;
        RECT 436.950 124.950 439.050 127.050 ;
        RECT 455.400 126.600 456.600 133.950 ;
        RECT 467.550 133.050 468.450 148.950 ;
        RECT 472.950 136.950 475.050 139.050 ;
        RECT 473.100 135.150 474.900 136.950 ;
        RECT 476.850 136.050 478.050 149.400 ;
        RECT 487.950 145.950 490.050 148.050 ;
        RECT 478.950 136.950 481.050 139.050 ;
        RECT 475.950 133.950 478.050 136.050 ;
        RECT 479.100 135.150 480.900 136.950 ;
        RECT 482.100 136.050 483.900 137.850 ;
        RECT 481.950 133.950 484.050 136.050 ;
        RECT 466.800 130.950 468.900 133.050 ;
        RECT 475.950 129.750 477.150 133.950 ;
        RECT 473.400 128.700 477.150 129.750 ;
        RECT 473.400 126.600 474.600 128.700 ;
        RECT 451.500 125.400 456.600 126.600 ;
        RECT 371.400 120.600 373.200 123.600 ;
        RECT 388.800 120.600 390.600 123.600 ;
        RECT 409.800 120.600 411.600 123.600 ;
        RECT 428.400 120.600 430.200 123.600 ;
        RECT 451.500 120.600 453.300 125.400 ;
        RECT 472.800 120.600 474.600 126.600 ;
        RECT 475.800 125.700 483.600 127.050 ;
        RECT 475.800 120.600 477.600 125.700 ;
        RECT 481.800 120.600 483.600 125.700 ;
        RECT 488.550 124.050 489.450 145.950 ;
        RECT 499.500 144.600 501.300 155.400 ;
        RECT 497.700 143.400 501.300 144.600 ;
        RECT 518.400 149.400 520.200 155.400 ;
        RECT 541.800 149.400 543.600 155.400 ;
        RECT 563.400 149.400 565.200 155.400 ;
        RECT 586.800 149.400 588.600 155.400 ;
        RECT 604.800 149.400 606.600 155.400 ;
        RECT 625.800 149.400 627.600 155.400 ;
        RECT 649.800 149.400 651.600 155.400 ;
        RECT 497.700 136.050 498.600 143.400 ;
        RECT 514.950 136.950 517.050 139.050 ;
        RECT 494.100 133.050 495.900 134.850 ;
        RECT 496.950 133.950 499.050 136.050 ;
        RECT 515.100 135.150 516.900 136.950 ;
        RECT 518.400 136.050 519.600 149.400 ;
        RECT 520.950 136.950 523.050 139.050 ;
        RECT 538.950 136.950 541.050 139.050 ;
        RECT 493.950 130.950 496.050 133.050 ;
        RECT 487.950 121.950 490.050 124.050 ;
        RECT 497.700 123.600 498.600 133.950 ;
        RECT 500.100 133.050 501.900 134.850 ;
        RECT 517.950 133.950 520.050 136.050 ;
        RECT 521.100 135.150 522.900 136.950 ;
        RECT 539.100 135.150 540.900 136.950 ;
        RECT 542.400 136.050 543.600 149.400 ;
        RECT 544.950 136.950 547.050 139.050 ;
        RECT 559.950 136.950 562.050 139.050 ;
        RECT 541.950 133.950 544.050 136.050 ;
        RECT 545.100 135.150 546.900 136.950 ;
        RECT 560.100 135.150 561.900 136.950 ;
        RECT 563.850 136.050 565.050 149.400 ;
        RECT 565.950 136.950 568.050 139.050 ;
        RECT 562.950 133.950 565.050 136.050 ;
        RECT 566.100 135.150 567.900 136.950 ;
        RECT 569.100 136.050 570.900 137.850 ;
        RECT 583.950 136.950 586.050 139.050 ;
        RECT 568.950 133.950 571.050 136.050 ;
        RECT 584.100 135.150 585.900 136.950 ;
        RECT 587.400 136.050 588.600 149.400 ;
        RECT 605.400 142.050 606.600 149.400 ;
        RECT 589.950 136.950 592.050 139.050 ;
        RECT 604.950 136.950 607.050 142.050 ;
        RECT 586.950 133.950 589.050 136.050 ;
        RECT 590.100 135.150 591.900 136.950 ;
        RECT 499.950 130.950 502.050 133.050 ;
        RECT 518.400 128.700 519.600 133.950 ;
        RECT 542.400 128.700 543.600 133.950 ;
        RECT 562.950 129.750 564.150 133.950 ;
        RECT 518.400 127.800 522.600 128.700 ;
        RECT 497.400 120.600 499.200 123.600 ;
        RECT 520.800 120.600 522.600 127.800 ;
        RECT 539.400 127.800 543.600 128.700 ;
        RECT 560.400 128.700 564.150 129.750 ;
        RECT 587.400 128.700 588.600 133.950 ;
        RECT 539.400 120.600 541.200 127.800 ;
        RECT 560.400 126.600 561.600 128.700 ;
        RECT 584.400 127.800 588.600 128.700 ;
        RECT 559.800 120.600 561.600 126.600 ;
        RECT 562.800 125.700 570.600 127.050 ;
        RECT 562.800 120.600 564.600 125.700 ;
        RECT 568.800 120.600 570.600 125.700 ;
        RECT 584.400 120.600 586.200 127.800 ;
        RECT 605.400 123.600 606.600 136.950 ;
        RECT 608.100 136.050 609.900 137.850 ;
        RECT 620.100 136.050 621.900 137.850 ;
        RECT 622.950 136.950 625.050 139.050 ;
        RECT 607.950 133.950 610.050 136.050 ;
        RECT 619.950 133.950 622.050 136.050 ;
        RECT 623.100 135.150 624.900 136.950 ;
        RECT 625.950 136.050 627.150 149.400 ;
        RECT 628.950 136.950 631.050 139.050 ;
        RECT 646.950 136.950 649.050 139.050 ;
        RECT 625.950 133.950 628.050 136.050 ;
        RECT 629.100 135.150 630.900 136.950 ;
        RECT 647.100 135.150 648.900 136.950 ;
        RECT 650.400 136.050 651.600 149.400 ;
        RECT 656.550 143.400 658.350 155.400 ;
        RECT 664.050 149.400 665.850 155.400 ;
        RECT 661.950 147.300 665.850 149.400 ;
        RECT 671.850 148.500 673.650 155.400 ;
        RECT 679.650 149.400 681.450 155.400 ;
        RECT 680.250 148.500 681.450 149.400 ;
        RECT 670.950 147.450 677.550 148.500 ;
        RECT 670.950 146.700 672.750 147.450 ;
        RECT 675.750 146.700 677.550 147.450 ;
        RECT 680.250 146.400 685.050 148.500 ;
        RECT 663.150 144.600 665.850 146.400 ;
        RECT 666.750 145.800 668.550 146.400 ;
        RECT 666.750 144.900 673.050 145.800 ;
        RECT 680.250 145.500 681.450 146.400 ;
        RECT 666.750 144.600 668.550 144.900 ;
        RECT 664.950 143.700 665.850 144.600 ;
        RECT 652.950 136.950 655.050 139.050 ;
        RECT 649.950 133.950 652.050 136.050 ;
        RECT 653.100 135.150 654.900 136.950 ;
        RECT 656.550 136.050 657.750 143.400 ;
        RECT 661.950 142.800 664.050 143.700 ;
        RECT 664.950 142.800 670.050 143.700 ;
        RECT 659.850 141.600 664.050 142.800 ;
        RECT 658.950 139.800 660.750 141.600 ;
        RECT 656.550 135.750 661.050 136.050 ;
        RECT 656.550 133.950 662.850 135.750 ;
        RECT 626.850 129.750 628.050 133.950 ;
        RECT 626.850 128.700 630.600 129.750 ;
        RECT 650.400 128.700 651.600 133.950 ;
        RECT 604.800 120.600 606.600 123.600 ;
        RECT 620.400 125.700 628.200 127.050 ;
        RECT 620.400 120.600 622.200 125.700 ;
        RECT 626.400 120.600 628.200 125.700 ;
        RECT 629.400 126.600 630.600 128.700 ;
        RECT 647.400 127.800 651.600 128.700 ;
        RECT 629.400 120.600 631.200 126.600 ;
        RECT 647.400 120.600 649.200 127.800 ;
        RECT 656.550 126.600 657.750 133.950 ;
        RECT 669.150 130.200 670.050 142.800 ;
        RECT 672.150 142.800 673.050 144.900 ;
        RECT 673.950 144.300 681.450 145.500 ;
        RECT 673.950 143.700 675.750 144.300 ;
        RECT 688.050 143.400 689.850 155.400 ;
        RECT 672.150 142.500 680.550 142.800 ;
        RECT 688.950 142.500 689.850 143.400 ;
        RECT 672.150 141.900 689.850 142.500 ;
        RECT 678.750 141.300 689.850 141.900 ;
        RECT 678.750 141.000 680.550 141.300 ;
        RECT 676.950 134.400 679.050 136.050 ;
        RECT 676.950 133.200 684.900 134.400 ;
        RECT 685.950 133.950 688.050 136.050 ;
        RECT 683.100 132.600 684.900 133.200 ;
        RECT 686.100 132.150 687.900 133.950 ;
        RECT 680.100 131.400 681.900 132.000 ;
        RECT 686.100 131.400 687.000 132.150 ;
        RECT 680.100 130.200 687.000 131.400 ;
        RECT 669.150 129.000 681.150 130.200 ;
        RECT 669.150 128.400 670.950 129.000 ;
        RECT 680.100 127.200 681.150 129.000 ;
        RECT 656.550 120.600 658.350 126.600 ;
        RECT 661.950 125.700 664.050 126.600 ;
        RECT 661.950 124.500 665.700 125.700 ;
        RECT 676.350 125.550 678.150 126.300 ;
        RECT 664.650 123.600 665.700 124.500 ;
        RECT 673.200 124.500 678.150 125.550 ;
        RECT 679.650 125.400 681.450 127.200 ;
        RECT 688.950 126.600 689.850 141.300 ;
        RECT 682.950 124.500 685.050 126.600 ;
        RECT 673.200 123.600 674.250 124.500 ;
        RECT 682.950 123.600 684.000 124.500 ;
        RECT 664.650 120.600 666.450 123.600 ;
        RECT 672.450 120.600 674.250 123.600 ;
        RECT 680.250 122.700 684.000 123.600 ;
        RECT 680.250 120.600 682.050 122.700 ;
        RECT 688.050 120.600 689.850 126.600 ;
        RECT 703.500 143.400 705.300 155.400 ;
        RECT 709.800 149.400 711.600 155.400 ;
        RECT 727.800 149.400 729.600 155.400 ;
        RECT 751.800 149.400 753.600 155.400 ;
        RECT 773.400 149.400 775.200 155.400 ;
        RECT 797.400 149.400 799.200 155.400 ;
        RECT 820.800 149.400 822.600 155.400 ;
        RECT 845.400 149.400 847.200 155.400 ;
        RECT 866.400 149.400 868.200 155.400 ;
        RECT 886.800 149.400 888.600 155.400 ;
        RECT 703.500 136.050 704.700 143.400 ;
        RECT 710.400 142.500 711.600 149.400 ;
        RECT 705.600 141.600 711.600 142.500 ;
        RECT 705.600 140.700 707.850 141.600 ;
        RECT 703.500 133.950 706.050 136.050 ;
        RECT 703.500 126.600 704.700 133.950 ;
        RECT 706.950 129.300 707.850 140.700 ;
        RECT 710.100 136.050 711.900 137.850 ;
        RECT 722.100 136.050 723.900 137.850 ;
        RECT 724.950 136.950 727.050 139.050 ;
        RECT 709.950 133.950 712.050 136.050 ;
        RECT 721.950 133.950 724.050 136.050 ;
        RECT 725.100 135.150 726.900 136.950 ;
        RECT 727.950 136.050 729.150 149.400 ;
        RECT 730.950 136.950 733.050 139.050 ;
        RECT 748.950 136.950 751.050 139.050 ;
        RECT 727.950 133.950 730.050 136.050 ;
        RECT 731.100 135.150 732.900 136.950 ;
        RECT 749.100 135.150 750.900 136.950 ;
        RECT 752.400 136.050 753.600 149.400 ;
        RECT 754.950 136.950 757.050 139.050 ;
        RECT 769.950 136.950 772.050 139.050 ;
        RECT 751.950 133.950 754.050 136.050 ;
        RECT 755.100 135.150 756.900 136.950 ;
        RECT 770.100 135.150 771.900 136.950 ;
        RECT 773.850 136.050 775.050 149.400 ;
        RECT 784.950 142.950 787.050 145.050 ;
        RECT 775.950 136.950 778.050 139.050 ;
        RECT 772.950 133.950 775.050 136.050 ;
        RECT 776.100 135.150 777.900 136.950 ;
        RECT 779.100 136.050 780.900 137.850 ;
        RECT 778.950 133.950 781.050 136.050 ;
        RECT 705.600 128.400 707.850 129.300 ;
        RECT 728.850 129.750 730.050 133.950 ;
        RECT 728.850 128.700 732.600 129.750 ;
        RECT 752.400 128.700 753.600 133.950 ;
        RECT 772.950 129.750 774.150 133.950 ;
        RECT 785.550 133.050 786.450 142.950 ;
        RECT 793.950 136.950 796.050 139.050 ;
        RECT 794.100 135.150 795.900 136.950 ;
        RECT 797.850 136.050 799.050 149.400 ;
        RECT 799.950 136.950 802.050 139.050 ;
        RECT 796.950 133.950 799.050 136.050 ;
        RECT 800.100 135.150 801.900 136.950 ;
        RECT 803.100 136.050 804.900 137.850 ;
        RECT 815.100 136.050 816.900 137.850 ;
        RECT 817.950 136.950 820.050 139.050 ;
        RECT 802.950 133.950 805.050 136.050 ;
        RECT 814.950 133.950 817.050 136.050 ;
        RECT 818.100 135.150 819.900 136.950 ;
        RECT 820.950 136.050 822.150 149.400 ;
        RECT 823.950 136.950 826.050 139.050 ;
        RECT 841.950 136.950 844.050 139.050 ;
        RECT 820.950 133.950 823.050 136.050 ;
        RECT 824.100 135.150 825.900 136.950 ;
        RECT 842.100 135.150 843.900 136.950 ;
        RECT 845.850 136.050 847.050 149.400 ;
        RECT 866.400 142.050 867.600 149.400 ;
        RECT 847.950 136.950 850.050 139.050 ;
        RECT 784.950 130.950 787.050 133.050 ;
        RECT 796.950 129.750 798.150 133.950 ;
        RECT 705.600 127.500 711.600 128.400 ;
        RECT 703.500 120.600 705.300 126.600 ;
        RECT 710.400 123.600 711.600 127.500 ;
        RECT 709.800 120.600 711.600 123.600 ;
        RECT 722.400 125.700 730.200 127.050 ;
        RECT 722.400 120.600 724.200 125.700 ;
        RECT 728.400 120.600 730.200 125.700 ;
        RECT 731.400 126.600 732.600 128.700 ;
        RECT 749.400 127.800 753.600 128.700 ;
        RECT 770.400 128.700 774.150 129.750 ;
        RECT 794.400 128.700 798.150 129.750 ;
        RECT 821.850 129.750 823.050 133.950 ;
        RECT 844.950 133.950 847.050 136.050 ;
        RECT 848.100 135.150 849.900 136.950 ;
        RECT 851.100 136.050 852.900 137.850 ;
        RECT 863.100 136.050 864.900 137.850 ;
        RECT 865.950 136.950 868.050 142.050 ;
        RECT 850.950 133.950 853.050 136.050 ;
        RECT 862.950 133.950 865.050 136.050 ;
        RECT 844.950 129.750 846.150 133.950 ;
        RECT 821.850 128.700 825.600 129.750 ;
        RECT 731.400 120.600 733.200 126.600 ;
        RECT 749.400 120.600 751.200 127.800 ;
        RECT 770.400 126.600 771.600 128.700 ;
        RECT 769.800 120.600 771.600 126.600 ;
        RECT 772.800 125.700 780.600 127.050 ;
        RECT 794.400 126.600 795.600 128.700 ;
        RECT 772.800 120.600 774.600 125.700 ;
        RECT 778.800 120.600 780.600 125.700 ;
        RECT 793.800 120.600 795.600 126.600 ;
        RECT 796.800 125.700 804.600 127.050 ;
        RECT 796.800 120.600 798.600 125.700 ;
        RECT 802.800 120.600 804.600 125.700 ;
        RECT 815.400 125.700 823.200 127.050 ;
        RECT 815.400 120.600 817.200 125.700 ;
        RECT 821.400 120.600 823.200 125.700 ;
        RECT 824.400 126.600 825.600 128.700 ;
        RECT 842.400 128.700 846.150 129.750 ;
        RECT 842.400 126.600 843.600 128.700 ;
        RECT 824.400 120.600 826.200 126.600 ;
        RECT 841.800 120.600 843.600 126.600 ;
        RECT 844.800 125.700 852.600 127.050 ;
        RECT 844.800 120.600 846.600 125.700 ;
        RECT 850.800 120.600 852.600 125.700 ;
        RECT 866.400 123.600 867.600 136.950 ;
        RECT 881.100 136.050 882.900 137.850 ;
        RECT 883.950 136.950 886.050 139.050 ;
        RECT 880.950 133.950 883.050 136.050 ;
        RECT 884.100 135.150 885.900 136.950 ;
        RECT 886.950 136.050 888.150 149.400 ;
        RECT 889.950 136.950 892.050 139.050 ;
        RECT 886.950 133.950 889.050 136.050 ;
        RECT 890.100 135.150 891.900 136.950 ;
        RECT 887.850 129.750 889.050 133.950 ;
        RECT 887.850 128.700 891.600 129.750 ;
        RECT 881.400 125.700 889.200 127.050 ;
        RECT 866.400 120.600 868.200 123.600 ;
        RECT 881.400 120.600 883.200 125.700 ;
        RECT 887.400 120.600 889.200 125.700 ;
        RECT 890.400 126.600 891.600 128.700 ;
        RECT 890.400 120.600 892.200 126.600 ;
        RECT 11.400 108.600 13.200 116.400 ;
        RECT 18.900 112.200 20.700 116.400 ;
        RECT 18.900 110.400 21.600 112.200 ;
        RECT 40.500 111.600 42.300 116.400 ;
        RECT 64.800 113.400 66.600 116.400 ;
        RECT 40.500 110.400 45.600 111.600 ;
        RECT 17.100 108.600 18.900 109.500 ;
        RECT 11.400 107.700 18.900 108.600 ;
        RECT 11.100 103.050 12.900 104.850 ;
        RECT 10.950 100.950 13.050 103.050 ;
        RECT 14.400 87.600 15.300 107.700 ;
        RECT 20.700 103.050 21.600 110.400 ;
        RECT 44.400 103.050 45.600 110.400 ;
        RECT 61.950 103.950 64.050 106.050 ;
        RECT 16.950 100.950 19.050 103.050 ;
        RECT 19.950 100.950 22.050 103.050 ;
        RECT 17.100 99.150 18.900 100.950 ;
        RECT 20.700 93.600 21.600 100.950 ;
        RECT 35.100 100.050 36.900 101.850 ;
        RECT 37.950 100.950 40.050 103.050 ;
        RECT 34.950 97.950 37.050 100.050 ;
        RECT 38.100 99.150 39.900 100.950 ;
        RECT 41.100 100.050 42.900 101.850 ;
        RECT 43.950 100.950 46.050 103.050 ;
        RECT 62.100 102.150 63.900 103.950 ;
        RECT 65.400 103.050 66.300 113.400 ;
        RECT 82.800 110.400 84.600 116.400 ;
        RECT 83.400 108.300 84.600 110.400 ;
        RECT 85.800 111.300 87.600 116.400 ;
        RECT 91.800 111.300 93.600 116.400 ;
        RECT 98.100 112.950 100.200 115.050 ;
        RECT 106.800 113.400 108.600 116.400 ;
        RECT 85.800 109.950 93.600 111.300 ;
        RECT 83.400 107.250 87.150 108.300 ;
        RECT 67.950 103.950 70.050 106.050 ;
        RECT 64.950 100.950 67.050 103.050 ;
        RECT 68.100 102.150 69.900 103.950 ;
        RECT 85.950 103.050 87.150 107.250 ;
        RECT 40.950 97.950 43.050 100.050 ;
        RECT 44.400 93.600 45.600 100.950 ;
        RECT 65.400 93.600 66.300 100.950 ;
        RECT 83.100 100.050 84.900 101.850 ;
        RECT 85.950 100.950 88.050 103.050 ;
        RECT 82.950 97.950 85.050 100.050 ;
        RECT 14.400 81.600 16.200 87.600 ;
        RECT 20.700 81.600 22.500 93.600 ;
        RECT 35.400 92.700 43.200 93.600 ;
        RECT 35.400 81.600 37.200 92.700 ;
        RECT 41.400 81.600 43.200 92.700 ;
        RECT 44.400 81.600 46.200 93.600 ;
        RECT 62.700 92.400 66.300 93.600 ;
        RECT 62.700 81.600 64.500 92.400 ;
        RECT 86.850 87.600 88.050 100.950 ;
        RECT 89.100 100.050 90.900 101.850 ;
        RECT 91.950 100.950 94.050 103.050 ;
        RECT 88.950 97.950 91.050 100.050 ;
        RECT 92.100 99.150 93.900 100.950 ;
        RECT 86.400 81.600 88.200 87.600 ;
        RECT 98.550 85.050 99.450 112.950 ;
        RECT 107.400 100.050 108.600 113.400 ;
        RECT 124.800 110.400 126.600 116.400 ;
        RECT 125.400 108.300 126.600 110.400 ;
        RECT 127.800 111.300 129.600 116.400 ;
        RECT 133.800 111.300 135.600 116.400 ;
        RECT 149.400 113.400 151.200 116.400 ;
        RECT 127.800 109.950 135.600 111.300 ;
        RECT 125.400 107.250 129.150 108.300 ;
        RECT 118.950 103.950 121.050 106.050 ;
        RECT 109.950 100.950 112.050 103.050 ;
        RECT 106.950 94.950 109.050 100.050 ;
        RECT 110.100 99.150 111.900 100.950 ;
        RECT 107.400 87.600 108.600 94.950 ;
        RECT 119.550 91.050 120.450 103.950 ;
        RECT 127.950 103.050 129.150 107.250 ;
        RECT 145.950 103.950 148.050 106.050 ;
        RECT 125.100 100.050 126.900 101.850 ;
        RECT 127.950 100.950 130.050 103.050 ;
        RECT 124.950 97.950 127.050 100.050 ;
        RECT 118.950 88.950 121.050 91.050 ;
        RECT 128.850 87.600 130.050 100.950 ;
        RECT 131.100 100.050 132.900 101.850 ;
        RECT 133.950 100.950 136.050 103.050 ;
        RECT 146.100 102.150 147.900 103.950 ;
        RECT 149.700 103.050 150.600 113.400 ;
        RECT 158.550 110.400 160.350 116.400 ;
        RECT 166.650 113.400 168.450 116.400 ;
        RECT 174.450 113.400 176.250 116.400 ;
        RECT 182.250 114.300 184.050 116.400 ;
        RECT 182.250 113.400 186.000 114.300 ;
        RECT 166.650 112.500 167.700 113.400 ;
        RECT 163.950 111.300 167.700 112.500 ;
        RECT 175.200 112.500 176.250 113.400 ;
        RECT 184.950 112.500 186.000 113.400 ;
        RECT 175.200 111.450 180.150 112.500 ;
        RECT 163.950 110.400 166.050 111.300 ;
        RECT 178.350 110.700 180.150 111.450 ;
        RECT 151.950 103.950 154.050 106.050 ;
        RECT 148.950 100.950 151.050 103.050 ;
        RECT 152.100 102.150 153.900 103.950 ;
        RECT 158.550 103.050 159.750 110.400 ;
        RECT 181.650 109.800 183.450 111.600 ;
        RECT 184.950 110.400 187.050 112.500 ;
        RECT 190.050 110.400 191.850 116.400 ;
        RECT 206.400 113.400 208.200 116.400 ;
        RECT 171.150 108.000 172.950 108.600 ;
        RECT 182.100 108.000 183.150 109.800 ;
        RECT 171.150 106.800 183.150 108.000 ;
        RECT 158.550 101.250 164.850 103.050 ;
        RECT 158.550 100.950 163.050 101.250 ;
        RECT 130.950 97.950 133.050 100.050 ;
        RECT 134.100 99.150 135.900 100.950 ;
        RECT 149.700 93.600 150.600 100.950 ;
        RECT 158.550 93.600 159.750 100.950 ;
        RECT 160.950 95.400 162.750 97.200 ;
        RECT 161.850 94.200 166.050 95.400 ;
        RECT 171.150 94.200 172.050 106.800 ;
        RECT 182.100 105.600 189.000 106.800 ;
        RECT 182.100 105.000 183.900 105.600 ;
        RECT 188.100 104.850 189.000 105.600 ;
        RECT 185.100 103.800 186.900 104.400 ;
        RECT 178.950 102.600 186.900 103.800 ;
        RECT 188.100 103.050 189.900 104.850 ;
        RECT 178.950 100.950 181.050 102.600 ;
        RECT 187.950 100.950 190.050 103.050 ;
        RECT 180.750 95.700 182.550 96.000 ;
        RECT 190.950 95.700 191.850 110.400 ;
        RECT 202.950 103.950 205.050 106.050 ;
        RECT 203.100 102.150 204.900 103.950 ;
        RECT 206.700 103.050 207.600 113.400 ;
        RECT 227.400 109.200 229.200 116.400 ;
        RECT 238.950 112.950 241.050 115.050 ;
        RECT 227.400 108.300 231.600 109.200 ;
        RECT 208.950 103.950 211.050 106.050 ;
        RECT 205.950 100.950 208.050 103.050 ;
        RECT 209.100 102.150 210.900 103.950 ;
        RECT 230.400 103.050 231.600 108.300 ;
        RECT 193.950 97.950 196.050 100.050 ;
        RECT 180.750 95.100 191.850 95.700 ;
        RECT 149.700 92.400 153.300 93.600 ;
        RECT 97.950 82.950 100.050 85.050 ;
        RECT 106.800 81.600 108.600 87.600 ;
        RECT 128.400 81.600 130.200 87.600 ;
        RECT 151.500 81.600 153.300 92.400 ;
        RECT 158.550 81.600 160.350 93.600 ;
        RECT 163.950 93.300 166.050 94.200 ;
        RECT 166.950 93.300 172.050 94.200 ;
        RECT 174.150 94.500 191.850 95.100 ;
        RECT 174.150 94.200 182.550 94.500 ;
        RECT 166.950 92.400 167.850 93.300 ;
        RECT 165.150 90.600 167.850 92.400 ;
        RECT 168.750 92.100 170.550 92.400 ;
        RECT 174.150 92.100 175.050 94.200 ;
        RECT 190.950 93.600 191.850 94.500 ;
        RECT 168.750 91.200 175.050 92.100 ;
        RECT 175.950 92.700 177.750 93.300 ;
        RECT 175.950 91.500 183.450 92.700 ;
        RECT 168.750 90.600 170.550 91.200 ;
        RECT 182.250 90.600 183.450 91.500 ;
        RECT 163.950 87.600 167.850 89.700 ;
        RECT 172.950 89.550 174.750 90.300 ;
        RECT 177.750 89.550 179.550 90.300 ;
        RECT 172.950 88.500 179.550 89.550 ;
        RECT 182.250 88.500 187.050 90.600 ;
        RECT 166.050 81.600 167.850 87.600 ;
        RECT 173.850 81.600 175.650 88.500 ;
        RECT 182.250 87.600 183.450 88.500 ;
        RECT 181.650 81.600 183.450 87.600 ;
        RECT 190.050 81.600 191.850 93.600 ;
        RECT 194.550 85.050 195.450 97.950 ;
        RECT 206.700 93.600 207.600 100.950 ;
        RECT 227.100 100.050 228.900 101.850 ;
        RECT 229.950 100.950 232.050 103.050 ;
        RECT 226.950 97.950 229.050 100.050 ;
        RECT 206.700 92.400 210.300 93.600 ;
        RECT 193.950 82.950 196.050 85.050 ;
        RECT 208.500 81.600 210.300 92.400 ;
        RECT 230.400 87.600 231.600 100.950 ;
        RECT 233.100 100.050 234.900 101.850 ;
        RECT 232.950 97.950 235.050 100.050 ;
        RECT 239.550 97.050 240.450 112.950 ;
        RECT 245.400 111.300 247.200 116.400 ;
        RECT 251.400 111.300 253.200 116.400 ;
        RECT 245.400 109.950 253.200 111.300 ;
        RECT 254.400 110.400 256.200 116.400 ;
        RECT 254.400 108.300 255.600 110.400 ;
        RECT 274.800 109.200 276.600 116.400 ;
        RECT 251.850 107.250 255.600 108.300 ;
        RECT 272.400 108.300 276.600 109.200 ;
        RECT 300.000 110.400 301.800 116.400 ;
        RECT 319.500 110.400 321.300 116.400 ;
        RECT 325.800 113.400 327.600 116.400 ;
        RECT 251.850 103.050 253.050 107.250 ;
        RECT 272.400 103.050 273.600 108.300 ;
        RECT 293.100 103.050 294.900 104.850 ;
        RECT 295.950 103.950 298.050 106.050 ;
        RECT 244.950 100.950 247.050 103.050 ;
        RECT 245.100 99.150 246.900 100.950 ;
        RECT 248.100 100.050 249.900 101.850 ;
        RECT 250.950 100.950 253.050 103.050 ;
        RECT 247.950 97.950 250.050 100.050 ;
        RECT 238.950 94.950 241.050 97.050 ;
        RECT 250.950 87.600 252.150 100.950 ;
        RECT 254.100 100.050 255.900 101.850 ;
        RECT 269.100 100.050 270.900 101.850 ;
        RECT 271.950 100.950 274.050 103.050 ;
        RECT 253.950 97.950 256.050 100.050 ;
        RECT 268.950 97.950 271.050 100.050 ;
        RECT 272.400 87.600 273.600 100.950 ;
        RECT 275.100 100.050 276.900 101.850 ;
        RECT 292.950 100.950 295.050 103.050 ;
        RECT 296.100 102.150 297.900 103.950 ;
        RECT 300.000 103.050 301.050 110.400 ;
        RECT 301.950 103.950 304.050 106.050 ;
        RECT 298.950 100.950 301.050 103.050 ;
        RECT 302.100 102.150 303.900 103.950 ;
        RECT 305.100 103.050 306.900 104.850 ;
        RECT 319.500 103.050 320.700 110.400 ;
        RECT 326.400 109.500 327.600 113.400 ;
        RECT 343.800 110.400 345.600 116.400 ;
        RECT 349.800 110.400 351.600 116.400 ;
        RECT 367.800 113.400 369.600 116.400 ;
        RECT 321.600 108.600 327.600 109.500 ;
        RECT 344.400 109.500 345.600 110.400 ;
        RECT 350.400 109.500 351.600 110.400 ;
        RECT 321.600 107.700 323.850 108.600 ;
        RECT 304.950 100.950 307.050 103.050 ;
        RECT 319.500 100.950 322.050 103.050 ;
        RECT 274.950 97.950 277.050 100.050 ;
        RECT 300.000 95.400 300.900 100.950 ;
        RECT 295.800 94.500 300.900 95.400 ;
        RECT 229.800 81.600 231.600 87.600 ;
        RECT 250.800 81.600 252.600 87.600 ;
        RECT 272.400 81.600 274.200 87.600 ;
        RECT 292.800 82.500 294.600 93.600 ;
        RECT 295.800 83.400 297.600 94.500 ;
        RECT 319.500 93.600 320.700 100.950 ;
        RECT 322.950 96.300 323.850 107.700 ;
        RECT 344.400 108.300 351.600 109.500 ;
        RECT 344.400 103.050 345.600 108.300 ;
        RECT 325.950 100.950 328.050 103.050 ;
        RECT 343.950 100.950 346.050 103.050 ;
        RECT 349.950 100.950 352.050 103.050 ;
        RECT 326.100 99.150 327.900 100.950 ;
        RECT 321.600 95.400 323.850 96.300 ;
        RECT 344.400 95.400 345.600 100.950 ;
        RECT 350.100 99.150 351.900 100.950 ;
        RECT 368.400 100.050 369.600 113.400 ;
        RECT 385.800 110.400 387.600 116.400 ;
        RECT 386.400 108.300 387.600 110.400 ;
        RECT 388.800 111.300 390.600 116.400 ;
        RECT 394.800 111.300 396.600 116.400 ;
        RECT 412.800 113.400 414.600 116.400 ;
        RECT 431.400 113.400 433.200 116.400 ;
        RECT 388.800 109.950 396.600 111.300 ;
        RECT 386.400 107.250 390.150 108.300 ;
        RECT 388.950 103.050 390.150 107.250 ;
        RECT 409.950 103.950 412.050 106.050 ;
        RECT 370.950 100.950 373.050 103.050 ;
        RECT 321.600 94.500 327.600 95.400 ;
        RECT 298.800 92.400 306.600 93.300 ;
        RECT 298.800 82.500 300.600 92.400 ;
        RECT 292.800 81.600 300.600 82.500 ;
        RECT 304.800 81.600 306.600 92.400 ;
        RECT 319.500 81.600 321.300 93.600 ;
        RECT 326.400 87.600 327.600 94.500 ;
        RECT 344.400 94.500 351.600 95.400 ;
        RECT 367.950 94.950 370.050 100.050 ;
        RECT 371.100 99.150 372.900 100.950 ;
        RECT 386.100 100.050 387.900 101.850 ;
        RECT 388.950 100.950 391.050 103.050 ;
        RECT 385.950 97.950 388.050 100.050 ;
        RECT 344.400 93.600 345.600 94.500 ;
        RECT 325.800 81.600 327.600 87.600 ;
        RECT 343.800 81.600 345.600 93.600 ;
        RECT 349.800 81.600 351.600 94.500 ;
        RECT 368.400 87.600 369.600 94.950 ;
        RECT 382.800 88.950 384.900 91.050 ;
        RECT 367.800 81.600 369.600 87.600 ;
        RECT 383.550 85.050 384.450 88.950 ;
        RECT 389.850 87.600 391.050 100.950 ;
        RECT 392.100 100.050 393.900 101.850 ;
        RECT 394.950 100.950 397.050 103.050 ;
        RECT 410.100 102.150 411.900 103.950 ;
        RECT 413.400 103.050 414.300 113.400 ;
        RECT 415.950 103.950 418.050 106.050 ;
        RECT 412.950 100.950 415.050 103.050 ;
        RECT 416.100 102.150 417.900 103.950 ;
        RECT 427.950 100.950 430.050 103.050 ;
        RECT 391.950 97.950 394.050 100.050 ;
        RECT 395.100 99.150 396.900 100.950 ;
        RECT 413.400 93.600 414.300 100.950 ;
        RECT 428.100 99.150 429.900 100.950 ;
        RECT 431.400 100.050 432.600 113.400 ;
        RECT 439.950 109.950 442.050 112.050 ;
        RECT 430.950 94.950 433.050 100.050 ;
        RECT 440.550 97.050 441.450 109.950 ;
        RECT 446.400 108.600 448.200 116.400 ;
        RECT 453.900 112.200 455.700 116.400 ;
        RECT 465.000 114.450 469.050 115.050 ;
        RECT 464.550 112.950 469.050 114.450 ;
        RECT 453.900 110.400 456.600 112.200 ;
        RECT 452.100 108.600 453.900 109.500 ;
        RECT 446.400 107.700 453.900 108.600 ;
        RECT 446.100 103.050 447.900 104.850 ;
        RECT 445.950 100.950 448.050 103.050 ;
        RECT 439.950 94.950 442.050 97.050 ;
        RECT 410.700 92.400 414.300 93.600 ;
        RECT 383.100 82.950 385.200 85.050 ;
        RECT 389.400 81.600 391.200 87.600 ;
        RECT 410.700 81.600 412.500 92.400 ;
        RECT 431.400 87.600 432.600 94.950 ;
        RECT 449.400 87.600 450.300 107.700 ;
        RECT 455.700 103.050 456.600 110.400 ;
        RECT 451.950 100.950 454.050 103.050 ;
        RECT 454.950 100.950 457.050 103.050 ;
        RECT 452.100 99.150 453.900 100.950 ;
        RECT 455.700 93.600 456.600 100.950 ;
        RECT 431.400 81.600 433.200 87.600 ;
        RECT 449.400 81.600 451.200 87.600 ;
        RECT 455.700 81.600 457.500 93.600 ;
        RECT 464.550 88.050 465.450 112.950 ;
        RECT 470.400 111.300 472.200 116.400 ;
        RECT 476.400 111.300 478.200 116.400 ;
        RECT 470.400 109.950 478.200 111.300 ;
        RECT 479.400 110.400 481.200 116.400 ;
        RECT 479.400 108.300 480.600 110.400 ;
        RECT 497.400 109.200 499.200 116.400 ;
        RECT 507.150 110.400 508.950 116.400 ;
        RECT 514.950 114.300 516.750 116.400 ;
        RECT 513.000 113.400 516.750 114.300 ;
        RECT 522.750 113.400 524.550 116.400 ;
        RECT 530.550 113.400 532.350 116.400 ;
        RECT 513.000 112.500 514.050 113.400 ;
        RECT 522.750 112.500 523.800 113.400 ;
        RECT 511.950 110.400 514.050 112.500 ;
        RECT 476.850 107.250 480.600 108.300 ;
        RECT 476.850 103.050 478.050 107.250 ;
        RECT 490.950 106.950 493.050 109.050 ;
        RECT 497.400 108.300 501.600 109.200 ;
        RECT 469.950 100.950 472.050 103.050 ;
        RECT 470.100 99.150 471.900 100.950 ;
        RECT 473.100 100.050 474.900 101.850 ;
        RECT 475.950 100.950 478.050 103.050 ;
        RECT 472.950 97.950 475.050 100.050 ;
        RECT 464.100 85.950 466.200 88.050 ;
        RECT 475.950 87.600 477.150 100.950 ;
        RECT 479.100 100.050 480.900 101.850 ;
        RECT 478.950 97.950 481.050 100.050 ;
        RECT 475.800 81.600 477.600 87.600 ;
        RECT 491.550 85.050 492.450 106.950 ;
        RECT 500.400 103.050 501.600 108.300 ;
        RECT 497.100 100.050 498.900 101.850 ;
        RECT 499.950 100.950 502.050 103.050 ;
        RECT 496.950 97.950 499.050 100.050 ;
        RECT 500.400 87.600 501.600 100.950 ;
        RECT 503.100 100.050 504.900 101.850 ;
        RECT 502.950 97.950 505.050 100.050 ;
        RECT 490.800 82.950 492.900 85.050 ;
        RECT 499.800 81.600 501.600 87.600 ;
        RECT 507.150 95.700 508.050 110.400 ;
        RECT 515.550 109.800 517.350 111.600 ;
        RECT 518.850 111.450 523.800 112.500 ;
        RECT 531.300 112.500 532.350 113.400 ;
        RECT 518.850 110.700 520.650 111.450 ;
        RECT 531.300 111.300 535.050 112.500 ;
        RECT 532.950 110.400 535.050 111.300 ;
        RECT 538.650 110.400 540.450 116.400 ;
        RECT 515.850 108.000 516.900 109.800 ;
        RECT 526.050 108.000 527.850 108.600 ;
        RECT 515.850 106.800 527.850 108.000 ;
        RECT 510.000 105.600 516.900 106.800 ;
        RECT 510.000 104.850 510.900 105.600 ;
        RECT 515.100 105.000 516.900 105.600 ;
        RECT 509.100 103.050 510.900 104.850 ;
        RECT 512.100 103.800 513.900 104.400 ;
        RECT 508.950 100.950 511.050 103.050 ;
        RECT 512.100 102.600 520.050 103.800 ;
        RECT 517.950 100.950 520.050 102.600 ;
        RECT 516.450 95.700 518.250 96.000 ;
        RECT 507.150 95.100 518.250 95.700 ;
        RECT 507.150 94.500 524.850 95.100 ;
        RECT 507.150 93.600 508.050 94.500 ;
        RECT 516.450 94.200 524.850 94.500 ;
        RECT 507.150 81.600 508.950 93.600 ;
        RECT 521.250 92.700 523.050 93.300 ;
        RECT 515.550 91.500 523.050 92.700 ;
        RECT 523.950 92.100 524.850 94.200 ;
        RECT 526.950 94.200 527.850 106.800 ;
        RECT 539.250 103.050 540.450 110.400 ;
        RECT 544.950 109.950 547.050 112.050 ;
        RECT 551.400 111.300 553.200 116.400 ;
        RECT 557.400 111.300 559.200 116.400 ;
        RECT 551.400 109.950 559.200 111.300 ;
        RECT 560.400 110.400 562.200 116.400 ;
        RECT 567.150 110.400 568.950 116.400 ;
        RECT 574.950 114.300 576.750 116.400 ;
        RECT 573.000 113.400 576.750 114.300 ;
        RECT 582.750 113.400 584.550 116.400 ;
        RECT 590.550 113.400 592.350 116.400 ;
        RECT 573.000 112.500 574.050 113.400 ;
        RECT 582.750 112.500 583.800 113.400 ;
        RECT 571.950 110.400 574.050 112.500 ;
        RECT 534.150 101.250 540.450 103.050 ;
        RECT 535.950 100.950 540.450 101.250 ;
        RECT 536.250 95.400 538.050 97.200 ;
        RECT 532.950 94.200 537.150 95.400 ;
        RECT 526.950 93.300 532.050 94.200 ;
        RECT 532.950 93.300 535.050 94.200 ;
        RECT 539.250 93.600 540.450 100.950 ;
        RECT 531.150 92.400 532.050 93.300 ;
        RECT 528.450 92.100 530.250 92.400 ;
        RECT 515.550 90.600 516.750 91.500 ;
        RECT 523.950 91.200 530.250 92.100 ;
        RECT 528.450 90.600 530.250 91.200 ;
        RECT 531.150 90.600 533.850 92.400 ;
        RECT 511.950 88.500 516.750 90.600 ;
        RECT 519.450 89.550 521.250 90.300 ;
        RECT 524.250 89.550 526.050 90.300 ;
        RECT 519.450 88.500 526.050 89.550 ;
        RECT 515.550 87.600 516.750 88.500 ;
        RECT 515.550 81.600 517.350 87.600 ;
        RECT 523.350 81.600 525.150 88.500 ;
        RECT 531.150 87.600 535.050 89.700 ;
        RECT 531.150 81.600 532.950 87.600 ;
        RECT 538.650 81.600 540.450 93.600 ;
        RECT 545.550 85.050 546.450 109.950 ;
        RECT 560.400 108.300 561.600 110.400 ;
        RECT 557.850 107.250 561.600 108.300 ;
        RECT 557.850 103.050 559.050 107.250 ;
        RECT 550.950 100.950 553.050 103.050 ;
        RECT 551.100 99.150 552.900 100.950 ;
        RECT 554.100 100.050 555.900 101.850 ;
        RECT 556.950 100.950 559.050 103.050 ;
        RECT 553.950 97.950 556.050 100.050 ;
        RECT 556.950 87.600 558.150 100.950 ;
        RECT 560.100 100.050 561.900 101.850 ;
        RECT 559.950 97.950 562.050 100.050 ;
        RECT 567.150 95.700 568.050 110.400 ;
        RECT 575.550 109.800 577.350 111.600 ;
        RECT 578.850 111.450 583.800 112.500 ;
        RECT 591.300 112.500 592.350 113.400 ;
        RECT 578.850 110.700 580.650 111.450 ;
        RECT 591.300 111.300 595.050 112.500 ;
        RECT 592.950 110.400 595.050 111.300 ;
        RECT 598.650 110.400 600.450 116.400 ;
        RECT 604.800 112.950 606.900 115.050 ;
        RECT 614.400 113.400 616.200 116.400 ;
        RECT 575.850 108.000 576.900 109.800 ;
        RECT 586.050 108.000 587.850 108.600 ;
        RECT 575.850 106.800 587.850 108.000 ;
        RECT 570.000 105.600 576.900 106.800 ;
        RECT 570.000 104.850 570.900 105.600 ;
        RECT 575.100 105.000 576.900 105.600 ;
        RECT 569.100 103.050 570.900 104.850 ;
        RECT 572.100 103.800 573.900 104.400 ;
        RECT 568.950 100.950 571.050 103.050 ;
        RECT 572.100 102.600 580.050 103.800 ;
        RECT 577.950 100.950 580.050 102.600 ;
        RECT 576.450 95.700 578.250 96.000 ;
        RECT 567.150 95.100 578.250 95.700 ;
        RECT 567.150 94.500 584.850 95.100 ;
        RECT 567.150 93.600 568.050 94.500 ;
        RECT 576.450 94.200 584.850 94.500 ;
        RECT 544.950 82.950 547.050 85.050 ;
        RECT 556.800 81.600 558.600 87.600 ;
        RECT 567.150 81.600 568.950 93.600 ;
        RECT 581.250 92.700 583.050 93.300 ;
        RECT 575.550 91.500 583.050 92.700 ;
        RECT 583.950 92.100 584.850 94.200 ;
        RECT 586.950 94.200 587.850 106.800 ;
        RECT 599.250 103.050 600.450 110.400 ;
        RECT 594.150 101.250 600.450 103.050 ;
        RECT 595.950 100.950 600.450 101.250 ;
        RECT 596.250 95.400 598.050 97.200 ;
        RECT 592.950 94.200 597.150 95.400 ;
        RECT 586.950 93.300 592.050 94.200 ;
        RECT 592.950 93.300 595.050 94.200 ;
        RECT 599.250 93.600 600.450 100.950 ;
        RECT 591.150 92.400 592.050 93.300 ;
        RECT 588.450 92.100 590.250 92.400 ;
        RECT 575.550 90.600 576.750 91.500 ;
        RECT 583.950 91.200 590.250 92.100 ;
        RECT 588.450 90.600 590.250 91.200 ;
        RECT 591.150 90.600 593.850 92.400 ;
        RECT 571.950 88.500 576.750 90.600 ;
        RECT 579.450 89.550 581.250 90.300 ;
        RECT 584.250 89.550 586.050 90.300 ;
        RECT 579.450 88.500 586.050 89.550 ;
        RECT 575.550 87.600 576.750 88.500 ;
        RECT 575.550 81.600 577.350 87.600 ;
        RECT 583.350 81.600 585.150 88.500 ;
        RECT 591.150 87.600 595.050 89.700 ;
        RECT 591.150 81.600 592.950 87.600 ;
        RECT 598.650 81.600 600.450 93.600 ;
        RECT 605.550 88.050 606.450 112.950 ;
        RECT 610.950 103.950 613.050 106.050 ;
        RECT 611.100 102.150 612.900 103.950 ;
        RECT 614.700 103.050 615.600 113.400 ;
        RECT 639.000 108.000 640.800 116.400 ;
        RECT 646.950 112.950 649.050 115.050 ;
        RECT 639.000 106.800 642.300 108.000 ;
        RECT 616.950 103.950 619.050 106.050 ;
        RECT 613.950 100.950 616.050 103.050 ;
        RECT 617.100 102.150 618.900 103.950 ;
        RECT 641.400 103.050 642.300 106.800 ;
        RECT 614.700 93.600 615.600 100.950 ;
        RECT 632.100 100.050 633.900 101.850 ;
        RECT 634.950 100.950 637.050 103.050 ;
        RECT 631.950 97.950 634.050 100.050 ;
        RECT 635.100 99.150 636.900 100.950 ;
        RECT 638.100 100.050 639.900 101.850 ;
        RECT 640.950 100.950 643.050 103.050 ;
        RECT 637.950 97.950 640.050 100.050 ;
        RECT 614.700 92.400 618.300 93.600 ;
        RECT 604.950 85.950 607.050 88.050 ;
        RECT 616.500 81.600 618.300 92.400 ;
        RECT 641.400 88.800 642.300 100.950 ;
        RECT 647.550 91.050 648.450 112.950 ;
        RECT 649.950 109.950 652.050 112.050 ;
        RECT 656.400 111.300 658.200 116.400 ;
        RECT 662.400 111.300 664.200 116.400 ;
        RECT 656.400 109.950 664.200 111.300 ;
        RECT 665.400 110.400 667.200 116.400 ;
        RECT 685.800 113.400 687.600 116.400 ;
        RECT 704.400 113.400 706.200 116.400 ;
        RECT 646.950 88.950 649.050 91.050 ;
        RECT 635.700 87.900 642.300 88.800 ;
        RECT 650.550 88.050 651.450 109.950 ;
        RECT 665.400 108.300 666.600 110.400 ;
        RECT 662.850 107.250 666.600 108.300 ;
        RECT 662.850 103.050 664.050 107.250 ;
        RECT 682.950 103.950 685.050 106.050 ;
        RECT 655.950 100.950 658.050 103.050 ;
        RECT 656.100 99.150 657.900 100.950 ;
        RECT 659.100 100.050 660.900 101.850 ;
        RECT 661.950 100.950 664.050 103.050 ;
        RECT 683.100 102.150 684.900 103.950 ;
        RECT 686.400 103.050 687.300 113.400 ;
        RECT 705.300 109.200 706.200 113.400 ;
        RECT 710.400 110.400 712.200 116.400 ;
        RECT 705.300 108.300 708.600 109.200 ;
        RECT 706.800 107.400 708.600 108.300 ;
        RECT 688.950 103.950 691.050 106.050 ;
        RECT 658.950 97.950 661.050 100.050 ;
        RECT 652.950 94.950 655.050 97.050 ;
        RECT 635.700 87.600 637.200 87.900 ;
        RECT 635.400 81.600 637.200 87.600 ;
        RECT 641.400 87.600 642.300 87.900 ;
        RECT 641.400 81.600 643.200 87.600 ;
        RECT 649.800 85.950 651.900 88.050 ;
        RECT 653.550 85.050 654.450 94.950 ;
        RECT 661.950 87.600 663.150 100.950 ;
        RECT 665.100 100.050 666.900 101.850 ;
        RECT 685.950 100.950 688.050 103.050 ;
        RECT 689.100 102.150 690.900 103.950 ;
        RECT 664.950 97.950 667.050 100.050 ;
        RECT 686.400 93.600 687.300 100.950 ;
        RECT 701.100 100.050 702.900 101.850 ;
        RECT 703.950 100.950 706.050 103.050 ;
        RECT 700.950 97.950 703.050 100.050 ;
        RECT 704.100 99.150 705.900 100.950 ;
        RECT 707.700 96.900 708.600 107.400 ;
        RECT 711.000 103.050 712.050 110.400 ;
        RECT 721.950 109.950 724.050 112.050 ;
        RECT 727.800 110.400 729.600 116.400 ;
        RECT 706.800 96.300 708.600 96.900 ;
        RECT 683.700 92.400 687.300 93.600 ;
        RECT 701.400 95.100 708.600 96.300 ;
        RECT 709.950 100.950 712.050 103.050 ;
        RECT 701.400 93.600 702.600 95.100 ;
        RECT 709.950 93.600 711.300 100.950 ;
        RECT 652.950 82.950 655.050 85.050 ;
        RECT 661.800 81.600 663.600 87.600 ;
        RECT 683.700 81.600 685.500 92.400 ;
        RECT 701.400 81.600 703.200 93.600 ;
        RECT 708.900 92.100 711.300 93.600 ;
        RECT 708.900 81.600 710.700 92.100 ;
        RECT 722.550 91.050 723.450 109.950 ;
        RECT 728.400 108.300 729.600 110.400 ;
        RECT 730.800 111.300 732.600 116.400 ;
        RECT 736.800 111.300 738.600 116.400 ;
        RECT 730.800 109.950 738.600 111.300 ;
        RECT 749.400 113.400 751.200 116.400 ;
        RECT 749.400 109.500 750.600 113.400 ;
        RECT 755.700 110.400 757.500 116.400 ;
        RECT 749.400 108.600 755.400 109.500 ;
        RECT 728.400 107.250 732.150 108.300 ;
        RECT 730.950 103.050 732.150 107.250 ;
        RECT 753.150 107.700 755.400 108.600 ;
        RECT 728.100 100.050 729.900 101.850 ;
        RECT 730.950 100.950 733.050 103.050 ;
        RECT 727.950 97.950 730.050 100.050 ;
        RECT 721.950 88.950 724.050 91.050 ;
        RECT 731.850 87.600 733.050 100.950 ;
        RECT 734.100 100.050 735.900 101.850 ;
        RECT 736.950 100.950 739.050 103.050 ;
        RECT 748.950 100.950 751.050 103.050 ;
        RECT 733.950 97.950 736.050 100.050 ;
        RECT 737.100 99.150 738.900 100.950 ;
        RECT 749.100 99.150 750.900 100.950 ;
        RECT 753.150 96.300 754.050 107.700 ;
        RECT 756.300 103.050 757.500 110.400 ;
        RECT 754.950 100.950 757.500 103.050 ;
        RECT 753.150 95.400 755.400 96.300 ;
        RECT 749.400 94.500 755.400 95.400 ;
        RECT 749.400 87.600 750.600 94.500 ;
        RECT 756.300 93.600 757.500 100.950 ;
        RECT 731.400 81.600 733.200 87.600 ;
        RECT 749.400 81.600 751.200 87.600 ;
        RECT 755.700 81.600 757.500 93.600 ;
        RECT 761.550 110.400 763.350 116.400 ;
        RECT 769.650 113.400 771.450 116.400 ;
        RECT 777.450 113.400 779.250 116.400 ;
        RECT 785.250 114.300 787.050 116.400 ;
        RECT 785.250 113.400 789.000 114.300 ;
        RECT 769.650 112.500 770.700 113.400 ;
        RECT 766.950 111.300 770.700 112.500 ;
        RECT 778.200 112.500 779.250 113.400 ;
        RECT 787.950 112.500 789.000 113.400 ;
        RECT 778.200 111.450 783.150 112.500 ;
        RECT 766.950 110.400 769.050 111.300 ;
        RECT 781.350 110.700 783.150 111.450 ;
        RECT 761.550 103.050 762.750 110.400 ;
        RECT 784.650 109.800 786.450 111.600 ;
        RECT 787.950 110.400 790.050 112.500 ;
        RECT 793.050 110.400 794.850 116.400 ;
        RECT 774.150 108.000 775.950 108.600 ;
        RECT 785.100 108.000 786.150 109.800 ;
        RECT 774.150 106.800 786.150 108.000 ;
        RECT 761.550 101.250 767.850 103.050 ;
        RECT 761.550 100.950 766.050 101.250 ;
        RECT 761.550 93.600 762.750 100.950 ;
        RECT 763.950 95.400 765.750 97.200 ;
        RECT 764.850 94.200 769.050 95.400 ;
        RECT 774.150 94.200 775.050 106.800 ;
        RECT 785.100 105.600 792.000 106.800 ;
        RECT 785.100 105.000 786.900 105.600 ;
        RECT 791.100 104.850 792.000 105.600 ;
        RECT 788.100 103.800 789.900 104.400 ;
        RECT 781.950 102.600 789.900 103.800 ;
        RECT 791.100 103.050 792.900 104.850 ;
        RECT 781.950 100.950 784.050 102.600 ;
        RECT 790.950 100.950 793.050 103.050 ;
        RECT 783.750 95.700 785.550 96.000 ;
        RECT 793.950 95.700 794.850 110.400 ;
        RECT 811.800 109.200 813.600 116.400 ;
        RECT 833.700 111.600 835.500 116.400 ;
        RECT 856.800 113.400 858.600 116.400 ;
        RECT 809.400 108.300 813.600 109.200 ;
        RECT 830.400 110.400 835.500 111.600 ;
        RECT 809.400 103.050 810.600 108.300 ;
        RECT 830.400 103.050 831.600 110.400 ;
        RECT 853.950 103.950 856.050 106.050 ;
        RECT 806.100 100.050 807.900 101.850 ;
        RECT 808.950 100.950 811.050 103.050 ;
        RECT 805.950 97.950 808.050 100.050 ;
        RECT 783.750 95.100 794.850 95.700 ;
        RECT 761.550 81.600 763.350 93.600 ;
        RECT 766.950 93.300 769.050 94.200 ;
        RECT 769.950 93.300 775.050 94.200 ;
        RECT 777.150 94.500 794.850 95.100 ;
        RECT 777.150 94.200 785.550 94.500 ;
        RECT 769.950 92.400 770.850 93.300 ;
        RECT 768.150 90.600 770.850 92.400 ;
        RECT 771.750 92.100 773.550 92.400 ;
        RECT 777.150 92.100 778.050 94.200 ;
        RECT 793.950 93.600 794.850 94.500 ;
        RECT 771.750 91.200 778.050 92.100 ;
        RECT 778.950 92.700 780.750 93.300 ;
        RECT 778.950 91.500 786.450 92.700 ;
        RECT 771.750 90.600 773.550 91.200 ;
        RECT 785.250 90.600 786.450 91.500 ;
        RECT 766.950 87.600 770.850 89.700 ;
        RECT 775.950 89.550 777.750 90.300 ;
        RECT 780.750 89.550 782.550 90.300 ;
        RECT 775.950 88.500 782.550 89.550 ;
        RECT 785.250 88.500 790.050 90.600 ;
        RECT 769.050 81.600 770.850 87.600 ;
        RECT 776.850 81.600 778.650 88.500 ;
        RECT 785.250 87.600 786.450 88.500 ;
        RECT 784.650 81.600 786.450 87.600 ;
        RECT 793.050 81.600 794.850 93.600 ;
        RECT 809.400 87.600 810.600 100.950 ;
        RECT 812.100 100.050 813.900 101.850 ;
        RECT 829.950 100.950 832.050 103.050 ;
        RECT 811.950 97.950 814.050 100.050 ;
        RECT 830.400 93.600 831.600 100.950 ;
        RECT 833.100 100.050 834.900 101.850 ;
        RECT 835.950 100.950 838.050 103.050 ;
        RECT 854.100 102.150 855.900 103.950 ;
        RECT 857.400 103.050 858.300 113.400 ;
        RECT 874.800 110.400 876.600 116.400 ;
        RECT 875.400 108.300 876.600 110.400 ;
        RECT 877.800 111.300 879.600 116.400 ;
        RECT 883.800 111.300 885.600 116.400 ;
        RECT 899.400 113.400 901.200 116.400 ;
        RECT 877.800 109.950 885.600 111.300 ;
        RECT 875.400 107.250 879.150 108.300 ;
        RECT 859.950 103.950 862.050 106.050 ;
        RECT 832.950 97.950 835.050 100.050 ;
        RECT 836.100 99.150 837.900 100.950 ;
        RECT 839.100 100.050 840.900 101.850 ;
        RECT 856.950 100.950 859.050 103.050 ;
        RECT 860.100 102.150 861.900 103.950 ;
        RECT 877.950 103.050 879.150 107.250 ;
        RECT 895.950 103.950 898.050 106.050 ;
        RECT 838.950 97.950 841.050 100.050 ;
        RECT 857.400 93.600 858.300 100.950 ;
        RECT 875.100 100.050 876.900 101.850 ;
        RECT 877.950 100.950 880.050 103.050 ;
        RECT 874.950 97.950 877.050 100.050 ;
        RECT 809.400 81.600 811.200 87.600 ;
        RECT 829.800 81.600 831.600 93.600 ;
        RECT 832.800 92.700 840.600 93.600 ;
        RECT 832.800 81.600 834.600 92.700 ;
        RECT 838.800 81.600 840.600 92.700 ;
        RECT 854.700 92.400 858.300 93.600 ;
        RECT 854.700 81.600 856.500 92.400 ;
        RECT 878.850 87.600 880.050 100.950 ;
        RECT 881.100 100.050 882.900 101.850 ;
        RECT 883.950 100.950 886.050 103.050 ;
        RECT 896.100 102.150 897.900 103.950 ;
        RECT 899.700 103.050 900.600 113.400 ;
        RECT 901.950 103.950 904.050 106.050 ;
        RECT 898.950 100.950 901.050 103.050 ;
        RECT 902.100 102.150 903.900 103.950 ;
        RECT 880.950 97.950 883.050 100.050 ;
        RECT 884.100 99.150 885.900 100.950 ;
        RECT 886.950 94.950 889.050 97.050 ;
        RECT 878.400 81.600 880.200 87.600 ;
        RECT 887.550 85.050 888.450 94.950 ;
        RECT 899.700 93.600 900.600 100.950 ;
        RECT 899.700 92.400 903.300 93.600 ;
        RECT 886.950 82.950 889.050 85.050 ;
        RECT 901.500 81.600 903.300 92.400 ;
        RECT 14.700 66.600 16.500 77.400 ;
        RECT 37.800 71.400 39.600 77.400 ;
        RECT 59.400 71.400 61.200 77.400 ;
        RECT 14.700 65.400 18.300 66.600 ;
        RECT 17.400 58.050 18.300 65.400 ;
        RECT 32.100 58.050 33.900 59.850 ;
        RECT 34.950 58.950 37.050 61.050 ;
        RECT 14.100 55.050 15.900 56.850 ;
        RECT 16.950 55.950 19.050 58.050 ;
        RECT 13.950 52.950 16.050 55.050 ;
        RECT 17.400 45.600 18.300 55.950 ;
        RECT 20.100 55.050 21.900 56.850 ;
        RECT 31.950 55.950 34.050 58.050 ;
        RECT 35.100 57.150 36.900 58.950 ;
        RECT 37.950 58.050 39.150 71.400 ;
        RECT 40.950 58.950 43.050 61.050 ;
        RECT 37.950 55.950 40.050 58.050 ;
        RECT 41.100 57.150 42.900 58.950 ;
        RECT 55.950 55.950 58.050 58.050 ;
        RECT 19.950 52.950 22.050 55.050 ;
        RECT 38.850 51.750 40.050 55.950 ;
        RECT 56.100 54.150 57.900 55.950 ;
        RECT 38.850 50.700 42.600 51.750 ;
        RECT 59.400 51.300 60.300 71.400 ;
        RECT 65.700 65.400 67.500 77.400 ;
        RECT 82.800 71.400 84.600 77.400 ;
        RECT 91.950 73.950 94.050 76.050 ;
        RECT 62.100 58.050 63.900 59.850 ;
        RECT 65.700 58.050 66.600 65.400 ;
        RECT 83.400 64.050 84.600 71.400 ;
        RECT 82.950 58.950 85.050 64.050 ;
        RECT 61.950 55.950 64.050 58.050 ;
        RECT 64.950 55.950 67.050 58.050 ;
        RECT 32.400 47.700 40.200 49.050 ;
        RECT 16.800 42.600 18.600 45.600 ;
        RECT 32.400 42.600 34.200 47.700 ;
        RECT 38.400 42.600 40.200 47.700 ;
        RECT 41.400 48.600 42.600 50.700 ;
        RECT 56.400 50.400 63.900 51.300 ;
        RECT 41.400 42.600 43.200 48.600 ;
        RECT 56.400 42.600 58.200 50.400 ;
        RECT 62.100 49.500 63.900 50.400 ;
        RECT 65.700 48.600 66.600 55.950 ;
        RECT 63.900 46.800 66.600 48.600 ;
        RECT 63.900 42.600 65.700 46.800 ;
        RECT 83.400 45.600 84.600 58.950 ;
        RECT 86.100 58.050 87.900 59.850 ;
        RECT 85.950 55.950 88.050 58.050 ;
        RECT 92.550 49.050 93.450 73.950 ;
        RECT 100.500 65.400 102.300 77.400 ;
        RECT 106.800 71.400 108.600 77.400 ;
        RECT 124.800 71.400 126.600 77.400 ;
        RECT 145.800 71.400 147.600 77.400 ;
        RECT 101.400 58.050 102.300 65.400 ;
        RECT 104.100 58.050 105.900 59.850 ;
        RECT 100.950 55.950 103.050 58.050 ;
        RECT 103.950 55.950 106.050 58.050 ;
        RECT 91.950 46.950 94.050 49.050 ;
        RECT 101.400 48.600 102.300 55.950 ;
        RECT 107.700 51.300 108.600 71.400 ;
        RECT 125.400 64.050 126.600 71.400 ;
        RECT 115.950 61.950 118.050 64.050 ;
        RECT 109.950 55.950 112.050 58.050 ;
        RECT 110.100 54.150 111.900 55.950 ;
        RECT 104.100 50.400 111.600 51.300 ;
        RECT 104.100 49.500 105.900 50.400 ;
        RECT 101.400 46.800 104.100 48.600 ;
        RECT 82.800 42.600 84.600 45.600 ;
        RECT 102.300 42.600 104.100 46.800 ;
        RECT 109.800 42.600 111.600 50.400 ;
        RECT 116.550 46.050 117.450 61.950 ;
        RECT 124.950 58.950 127.050 64.050 ;
        RECT 115.950 43.950 118.050 46.050 ;
        RECT 125.400 45.600 126.600 58.950 ;
        RECT 128.100 58.050 129.900 59.850 ;
        RECT 142.950 58.950 145.050 61.050 ;
        RECT 127.950 55.950 130.050 58.050 ;
        RECT 143.100 57.150 144.900 58.950 ;
        RECT 146.400 58.050 147.600 71.400 ;
        RECT 154.950 70.950 157.050 73.050 ;
        RECT 148.950 58.950 151.050 61.050 ;
        RECT 145.950 55.950 148.050 58.050 ;
        RECT 149.100 57.150 150.900 58.950 ;
        RECT 146.400 50.700 147.600 55.950 ;
        RECT 155.550 55.050 156.450 70.950 ;
        RECT 161.400 65.400 163.200 77.400 ;
        RECT 168.900 66.900 170.700 77.400 ;
        RECT 188.400 71.400 190.200 77.400 ;
        RECT 211.800 71.400 213.600 77.400 ;
        RECT 168.900 65.400 171.300 66.900 ;
        RECT 161.400 63.900 162.600 65.400 ;
        RECT 161.400 62.700 168.600 63.900 ;
        RECT 166.800 62.100 168.600 62.700 ;
        RECT 160.950 58.950 163.050 61.050 ;
        RECT 161.100 57.150 162.900 58.950 ;
        RECT 164.100 58.050 165.900 59.850 ;
        RECT 163.950 55.950 166.050 58.050 ;
        RECT 154.950 52.950 157.050 55.050 ;
        RECT 167.700 51.600 168.600 62.100 ;
        RECT 169.950 58.050 171.300 65.400 ;
        RECT 184.950 58.950 187.050 61.050 ;
        RECT 169.950 55.950 172.050 58.050 ;
        RECT 185.100 57.150 186.900 58.950 ;
        RECT 188.400 58.050 189.600 71.400 ;
        RECT 190.950 58.950 193.050 61.050 ;
        RECT 187.950 55.950 190.050 58.050 ;
        RECT 191.100 57.150 192.900 58.950 ;
        RECT 206.100 58.050 207.900 59.850 ;
        RECT 208.950 58.950 211.050 61.050 ;
        RECT 205.950 55.950 208.050 58.050 ;
        RECT 209.100 57.150 210.900 58.950 ;
        RECT 211.950 58.050 213.150 71.400 ;
        RECT 222.150 65.400 223.950 77.400 ;
        RECT 230.550 71.400 232.350 77.400 ;
        RECT 230.550 70.500 231.750 71.400 ;
        RECT 238.350 70.500 240.150 77.400 ;
        RECT 246.150 71.400 247.950 77.400 ;
        RECT 226.950 68.400 231.750 70.500 ;
        RECT 234.450 69.450 241.050 70.500 ;
        RECT 234.450 68.700 236.250 69.450 ;
        RECT 239.250 68.700 241.050 69.450 ;
        RECT 246.150 69.300 250.050 71.400 ;
        RECT 230.550 67.500 231.750 68.400 ;
        RECT 243.450 67.800 245.250 68.400 ;
        RECT 230.550 66.300 238.050 67.500 ;
        RECT 236.250 65.700 238.050 66.300 ;
        RECT 238.950 66.900 245.250 67.800 ;
        RECT 222.150 64.500 223.050 65.400 ;
        RECT 238.950 64.800 239.850 66.900 ;
        RECT 243.450 66.600 245.250 66.900 ;
        RECT 246.150 66.600 248.850 68.400 ;
        RECT 246.150 65.700 247.050 66.600 ;
        RECT 231.450 64.500 239.850 64.800 ;
        RECT 222.150 63.900 239.850 64.500 ;
        RECT 241.950 64.800 247.050 65.700 ;
        RECT 247.950 64.800 250.050 65.700 ;
        RECT 253.650 65.400 255.450 77.400 ;
        RECT 222.150 63.300 233.250 63.900 ;
        RECT 214.950 58.950 217.050 61.050 ;
        RECT 211.950 55.950 214.050 58.050 ;
        RECT 215.100 57.150 216.900 58.950 ;
        RECT 166.800 50.700 168.600 51.600 ;
        RECT 124.800 42.600 126.600 45.600 ;
        RECT 143.400 49.800 147.600 50.700 ;
        RECT 165.300 49.800 168.600 50.700 ;
        RECT 143.400 42.600 145.200 49.800 ;
        RECT 165.300 45.600 166.200 49.800 ;
        RECT 171.000 48.600 172.050 55.950 ;
        RECT 188.400 50.700 189.600 55.950 ;
        RECT 212.850 51.750 214.050 55.950 ;
        RECT 212.850 50.700 216.600 51.750 ;
        RECT 188.400 49.800 192.600 50.700 ;
        RECT 164.400 42.600 166.200 45.600 ;
        RECT 170.400 42.600 172.200 48.600 ;
        RECT 190.800 42.600 192.600 49.800 ;
        RECT 206.400 47.700 214.200 49.050 ;
        RECT 206.400 42.600 208.200 47.700 ;
        RECT 212.400 42.600 214.200 47.700 ;
        RECT 215.400 48.600 216.600 50.700 ;
        RECT 222.150 48.600 223.050 63.300 ;
        RECT 231.450 63.000 233.250 63.300 ;
        RECT 223.950 55.950 226.050 58.050 ;
        RECT 232.950 56.400 235.050 58.050 ;
        RECT 224.100 54.150 225.900 55.950 ;
        RECT 227.100 55.200 235.050 56.400 ;
        RECT 227.100 54.600 228.900 55.200 ;
        RECT 225.000 53.400 225.900 54.150 ;
        RECT 230.100 53.400 231.900 54.000 ;
        RECT 225.000 52.200 231.900 53.400 ;
        RECT 241.950 52.200 242.850 64.800 ;
        RECT 247.950 63.600 252.150 64.800 ;
        RECT 251.250 61.800 253.050 63.600 ;
        RECT 254.250 58.050 255.450 65.400 ;
        RECT 269.400 71.400 271.200 77.400 ;
        RECT 256.950 61.950 259.050 64.050 ;
        RECT 250.950 57.750 255.450 58.050 ;
        RECT 249.150 55.950 255.450 57.750 ;
        RECT 230.850 51.000 242.850 52.200 ;
        RECT 230.850 49.200 231.900 51.000 ;
        RECT 241.050 50.400 242.850 51.000 ;
        RECT 215.400 42.600 217.200 48.600 ;
        RECT 222.150 42.600 223.950 48.600 ;
        RECT 226.950 46.500 229.050 48.600 ;
        RECT 230.550 47.400 232.350 49.200 ;
        RECT 254.250 48.600 255.450 55.950 ;
        RECT 257.550 49.050 258.450 61.950 ;
        RECT 265.950 58.950 268.050 61.050 ;
        RECT 266.100 57.150 267.900 58.950 ;
        RECT 269.400 58.050 270.600 71.400 ;
        RECT 279.150 65.400 280.950 77.400 ;
        RECT 287.550 71.400 289.350 77.400 ;
        RECT 287.550 70.500 288.750 71.400 ;
        RECT 295.350 70.500 297.150 77.400 ;
        RECT 303.150 71.400 304.950 77.400 ;
        RECT 283.950 68.400 288.750 70.500 ;
        RECT 291.450 69.450 298.050 70.500 ;
        RECT 291.450 68.700 293.250 69.450 ;
        RECT 296.250 68.700 298.050 69.450 ;
        RECT 303.150 69.300 307.050 71.400 ;
        RECT 287.550 67.500 288.750 68.400 ;
        RECT 300.450 67.800 302.250 68.400 ;
        RECT 287.550 66.300 295.050 67.500 ;
        RECT 293.250 65.700 295.050 66.300 ;
        RECT 295.950 66.900 302.250 67.800 ;
        RECT 279.150 64.500 280.050 65.400 ;
        RECT 295.950 64.800 296.850 66.900 ;
        RECT 300.450 66.600 302.250 66.900 ;
        RECT 303.150 66.600 305.850 68.400 ;
        RECT 303.150 65.700 304.050 66.600 ;
        RECT 288.450 64.500 296.850 64.800 ;
        RECT 279.150 63.900 296.850 64.500 ;
        RECT 298.950 64.800 304.050 65.700 ;
        RECT 304.950 64.800 307.050 65.700 ;
        RECT 310.650 65.400 312.450 77.400 ;
        RECT 323.400 66.600 325.200 77.400 ;
        RECT 329.400 76.500 337.200 77.400 ;
        RECT 329.400 66.600 331.200 76.500 ;
        RECT 323.400 65.700 331.200 66.600 ;
        RECT 279.150 63.300 290.250 63.900 ;
        RECT 271.950 58.950 274.050 61.050 ;
        RECT 268.950 55.950 271.050 58.050 ;
        RECT 272.100 57.150 273.900 58.950 ;
        RECT 269.400 50.700 270.600 55.950 ;
        RECT 269.400 49.800 273.600 50.700 ;
        RECT 233.850 47.550 235.650 48.300 ;
        RECT 247.950 47.700 250.050 48.600 ;
        RECT 233.850 46.500 238.800 47.550 ;
        RECT 228.000 45.600 229.050 46.500 ;
        RECT 237.750 45.600 238.800 46.500 ;
        RECT 246.300 46.500 250.050 47.700 ;
        RECT 246.300 45.600 247.350 46.500 ;
        RECT 228.000 44.700 231.750 45.600 ;
        RECT 229.950 42.600 231.750 44.700 ;
        RECT 237.750 42.600 239.550 45.600 ;
        RECT 245.550 42.600 247.350 45.600 ;
        RECT 253.650 42.600 255.450 48.600 ;
        RECT 256.950 46.950 259.050 49.050 ;
        RECT 271.800 42.600 273.600 49.800 ;
        RECT 279.150 48.600 280.050 63.300 ;
        RECT 288.450 63.000 290.250 63.300 ;
        RECT 280.950 55.950 283.050 58.050 ;
        RECT 289.950 56.400 292.050 58.050 ;
        RECT 281.100 54.150 282.900 55.950 ;
        RECT 284.100 55.200 292.050 56.400 ;
        RECT 284.100 54.600 285.900 55.200 ;
        RECT 282.000 53.400 282.900 54.150 ;
        RECT 287.100 53.400 288.900 54.000 ;
        RECT 282.000 52.200 288.900 53.400 ;
        RECT 298.950 52.200 299.850 64.800 ;
        RECT 304.950 63.600 309.150 64.800 ;
        RECT 308.250 61.800 310.050 63.600 ;
        RECT 311.250 58.050 312.450 65.400 ;
        RECT 332.400 64.500 334.200 75.600 ;
        RECT 335.400 65.400 337.200 76.500 ;
        RECT 350.400 71.400 352.200 77.400 ;
        RECT 329.100 63.600 334.200 64.500 ;
        RECT 350.400 64.500 351.600 71.400 ;
        RECT 356.700 65.400 358.500 77.400 ;
        RECT 350.400 63.600 356.400 64.500 ;
        RECT 329.100 58.050 330.000 63.600 ;
        RECT 354.150 62.700 356.400 63.600 ;
        RECT 350.100 58.050 351.900 59.850 ;
        RECT 307.950 57.750 312.450 58.050 ;
        RECT 306.150 55.950 312.450 57.750 ;
        RECT 322.950 55.950 325.050 58.050 ;
        RECT 287.850 51.000 299.850 52.200 ;
        RECT 287.850 49.200 288.900 51.000 ;
        RECT 298.050 50.400 299.850 51.000 ;
        RECT 279.150 42.600 280.950 48.600 ;
        RECT 283.950 46.500 286.050 48.600 ;
        RECT 287.550 47.400 289.350 49.200 ;
        RECT 311.250 48.600 312.450 55.950 ;
        RECT 323.100 54.150 324.900 55.950 ;
        RECT 326.100 55.050 327.900 56.850 ;
        RECT 328.950 55.950 331.050 58.050 ;
        RECT 325.950 52.950 328.050 55.050 ;
        RECT 328.950 48.600 330.000 55.950 ;
        RECT 332.100 55.050 333.900 56.850 ;
        RECT 334.950 55.950 337.050 58.050 ;
        RECT 349.950 55.950 352.050 58.050 ;
        RECT 331.950 52.950 334.050 55.050 ;
        RECT 335.100 54.150 336.900 55.950 ;
        RECT 354.150 51.300 355.050 62.700 ;
        RECT 357.300 58.050 358.500 65.400 ;
        RECT 371.400 71.400 373.200 77.400 ;
        RECT 371.400 64.500 372.600 71.400 ;
        RECT 377.700 65.400 379.500 77.400 ;
        RECT 371.400 63.600 377.400 64.500 ;
        RECT 375.150 62.700 377.400 63.600 ;
        RECT 371.100 58.050 372.900 59.850 ;
        RECT 355.950 55.950 358.500 58.050 ;
        RECT 370.950 55.950 373.050 58.050 ;
        RECT 354.150 50.400 356.400 51.300 ;
        RECT 290.850 47.550 292.650 48.300 ;
        RECT 304.950 47.700 307.050 48.600 ;
        RECT 290.850 46.500 295.800 47.550 ;
        RECT 285.000 45.600 286.050 46.500 ;
        RECT 294.750 45.600 295.800 46.500 ;
        RECT 303.300 46.500 307.050 47.700 ;
        RECT 303.300 45.600 304.350 46.500 ;
        RECT 285.000 44.700 288.750 45.600 ;
        RECT 286.950 42.600 288.750 44.700 ;
        RECT 294.750 42.600 296.550 45.600 ;
        RECT 302.550 42.600 304.350 45.600 ;
        RECT 310.650 42.600 312.450 48.600 ;
        RECT 328.200 42.600 330.000 48.600 ;
        RECT 350.400 49.500 356.400 50.400 ;
        RECT 350.400 45.600 351.600 49.500 ;
        RECT 357.300 48.600 358.500 55.950 ;
        RECT 375.150 51.300 376.050 62.700 ;
        RECT 378.300 58.050 379.500 65.400 ;
        RECT 385.950 64.950 388.050 67.050 ;
        RECT 392.400 66.300 394.200 77.400 ;
        RECT 398.400 66.300 400.200 77.400 ;
        RECT 392.400 65.400 400.200 66.300 ;
        RECT 401.400 65.400 403.200 77.400 ;
        RECT 416.400 65.400 418.200 77.400 ;
        RECT 423.900 66.900 425.700 77.400 ;
        RECT 423.900 65.400 426.300 66.900 ;
        RECT 376.950 55.950 379.500 58.050 ;
        RECT 375.150 50.400 377.400 51.300 ;
        RECT 350.400 42.600 352.200 45.600 ;
        RECT 356.700 42.600 358.500 48.600 ;
        RECT 371.400 49.500 377.400 50.400 ;
        RECT 371.400 45.600 372.600 49.500 ;
        RECT 378.300 48.600 379.500 55.950 ;
        RECT 386.550 49.050 387.450 64.950 ;
        RECT 391.950 58.950 394.050 61.050 ;
        RECT 392.100 57.150 393.900 58.950 ;
        RECT 395.100 58.050 396.900 59.850 ;
        RECT 397.950 58.950 400.050 61.050 ;
        RECT 394.950 55.950 397.050 58.050 ;
        RECT 398.100 57.150 399.900 58.950 ;
        RECT 401.400 58.050 402.600 65.400 ;
        RECT 409.950 61.950 412.050 64.050 ;
        RECT 416.400 63.900 417.600 65.400 ;
        RECT 416.400 62.700 423.600 63.900 ;
        RECT 421.800 62.100 423.600 62.700 ;
        RECT 400.950 55.950 403.050 58.050 ;
        RECT 371.400 42.600 373.200 45.600 ;
        RECT 377.700 42.600 379.500 48.600 ;
        RECT 385.950 46.950 388.050 49.050 ;
        RECT 401.400 48.600 402.600 55.950 ;
        RECT 410.550 49.050 411.450 61.950 ;
        RECT 415.950 58.950 418.050 61.050 ;
        RECT 416.100 57.150 417.900 58.950 ;
        RECT 419.100 58.050 420.900 59.850 ;
        RECT 418.950 55.950 421.050 58.050 ;
        RECT 422.700 51.600 423.600 62.100 ;
        RECT 424.950 58.050 426.300 65.400 ;
        RECT 432.150 65.400 433.950 77.400 ;
        RECT 440.550 71.400 442.350 77.400 ;
        RECT 440.550 70.500 441.750 71.400 ;
        RECT 448.350 70.500 450.150 77.400 ;
        RECT 456.150 71.400 457.950 77.400 ;
        RECT 436.950 68.400 441.750 70.500 ;
        RECT 444.450 69.450 451.050 70.500 ;
        RECT 444.450 68.700 446.250 69.450 ;
        RECT 449.250 68.700 451.050 69.450 ;
        RECT 456.150 69.300 460.050 71.400 ;
        RECT 440.550 67.500 441.750 68.400 ;
        RECT 453.450 67.800 455.250 68.400 ;
        RECT 440.550 66.300 448.050 67.500 ;
        RECT 446.250 65.700 448.050 66.300 ;
        RECT 448.950 66.900 455.250 67.800 ;
        RECT 432.150 64.500 433.050 65.400 ;
        RECT 448.950 64.800 449.850 66.900 ;
        RECT 453.450 66.600 455.250 66.900 ;
        RECT 456.150 66.600 458.850 68.400 ;
        RECT 456.150 65.700 457.050 66.600 ;
        RECT 441.450 64.500 449.850 64.800 ;
        RECT 432.150 63.900 449.850 64.500 ;
        RECT 451.950 64.800 457.050 65.700 ;
        RECT 457.950 64.800 460.050 65.700 ;
        RECT 463.650 65.400 465.450 77.400 ;
        RECT 481.500 66.600 483.300 77.400 ;
        RECT 499.800 71.400 501.600 77.400 ;
        RECT 517.800 71.400 519.600 77.400 ;
        RECT 432.150 63.300 443.250 63.900 ;
        RECT 424.950 55.950 427.050 58.050 ;
        RECT 421.800 50.700 423.600 51.600 ;
        RECT 420.300 49.800 423.600 50.700 ;
        RECT 397.500 47.400 402.600 48.600 ;
        RECT 397.500 42.600 399.300 47.400 ;
        RECT 409.950 46.950 412.050 49.050 ;
        RECT 420.300 45.600 421.200 49.800 ;
        RECT 426.000 48.600 427.050 55.950 ;
        RECT 432.150 48.600 433.050 63.300 ;
        RECT 441.450 63.000 443.250 63.300 ;
        RECT 433.950 55.950 436.050 58.050 ;
        RECT 442.950 56.400 445.050 58.050 ;
        RECT 434.100 54.150 435.900 55.950 ;
        RECT 437.100 55.200 445.050 56.400 ;
        RECT 437.100 54.600 438.900 55.200 ;
        RECT 435.000 53.400 435.900 54.150 ;
        RECT 440.100 53.400 441.900 54.000 ;
        RECT 435.000 52.200 441.900 53.400 ;
        RECT 451.950 52.200 452.850 64.800 ;
        RECT 457.950 63.600 462.150 64.800 ;
        RECT 461.250 61.800 463.050 63.600 ;
        RECT 464.250 58.050 465.450 65.400 ;
        RECT 479.700 65.400 483.300 66.600 ;
        RECT 479.700 58.050 480.600 65.400 ;
        RECT 500.400 64.050 501.600 71.400 ;
        RECT 518.400 64.050 519.600 71.400 ;
        RECT 523.950 67.950 526.050 70.050 ;
        RECT 499.950 58.950 502.050 64.050 ;
        RECT 460.950 57.750 465.450 58.050 ;
        RECT 459.150 55.950 465.450 57.750 ;
        RECT 440.850 51.000 452.850 52.200 ;
        RECT 440.850 49.200 441.900 51.000 ;
        RECT 451.050 50.400 452.850 51.000 ;
        RECT 419.400 42.600 421.200 45.600 ;
        RECT 425.400 42.600 427.200 48.600 ;
        RECT 432.150 42.600 433.950 48.600 ;
        RECT 436.950 46.500 439.050 48.600 ;
        RECT 440.550 47.400 442.350 49.200 ;
        RECT 464.250 48.600 465.450 55.950 ;
        RECT 476.100 55.050 477.900 56.850 ;
        RECT 478.950 55.950 481.050 58.050 ;
        RECT 475.950 52.950 478.050 55.050 ;
        RECT 443.850 47.550 445.650 48.300 ;
        RECT 457.950 47.700 460.050 48.600 ;
        RECT 443.850 46.500 448.800 47.550 ;
        RECT 438.000 45.600 439.050 46.500 ;
        RECT 447.750 45.600 448.800 46.500 ;
        RECT 456.300 46.500 460.050 47.700 ;
        RECT 456.300 45.600 457.350 46.500 ;
        RECT 438.000 44.700 441.750 45.600 ;
        RECT 439.950 42.600 441.750 44.700 ;
        RECT 447.750 42.600 449.550 45.600 ;
        RECT 455.550 42.600 457.350 45.600 ;
        RECT 463.650 42.600 465.450 48.600 ;
        RECT 479.700 45.600 480.600 55.950 ;
        RECT 482.100 55.050 483.900 56.850 ;
        RECT 481.950 52.950 484.050 55.050 ;
        RECT 500.400 45.600 501.600 58.950 ;
        RECT 503.100 58.050 504.900 59.850 ;
        RECT 517.950 58.950 520.050 64.050 ;
        RECT 524.550 61.050 525.450 67.950 ;
        RECT 536.700 66.600 538.500 77.400 ;
        RECT 557.400 71.400 559.200 77.400 ;
        RECT 536.700 65.400 540.300 66.600 ;
        RECT 502.950 55.950 505.050 58.050 ;
        RECT 518.400 45.600 519.600 58.950 ;
        RECT 521.100 58.050 522.900 59.850 ;
        RECT 523.950 58.950 526.050 61.050 ;
        RECT 539.400 58.050 540.300 65.400 ;
        RECT 557.400 64.050 558.600 71.400 ;
        RECT 564.150 65.400 565.950 77.400 ;
        RECT 572.550 71.400 574.350 77.400 ;
        RECT 572.550 70.500 573.750 71.400 ;
        RECT 580.350 70.500 582.150 77.400 ;
        RECT 588.150 71.400 589.950 77.400 ;
        RECT 568.950 68.400 573.750 70.500 ;
        RECT 576.450 69.450 583.050 70.500 ;
        RECT 576.450 68.700 578.250 69.450 ;
        RECT 581.250 68.700 583.050 69.450 ;
        RECT 588.150 69.300 592.050 71.400 ;
        RECT 572.550 67.500 573.750 68.400 ;
        RECT 585.450 67.800 587.250 68.400 ;
        RECT 572.550 66.300 580.050 67.500 ;
        RECT 578.250 65.700 580.050 66.300 ;
        RECT 580.950 66.900 587.250 67.800 ;
        RECT 564.150 64.500 565.050 65.400 ;
        RECT 580.950 64.800 581.850 66.900 ;
        RECT 585.450 66.600 587.250 66.900 ;
        RECT 588.150 66.600 590.850 68.400 ;
        RECT 588.150 65.700 589.050 66.600 ;
        RECT 573.450 64.500 581.850 64.800 ;
        RECT 554.100 58.050 555.900 59.850 ;
        RECT 556.950 58.950 559.050 64.050 ;
        RECT 564.150 63.900 581.850 64.500 ;
        RECT 583.950 64.800 589.050 65.700 ;
        RECT 589.950 64.800 592.050 65.700 ;
        RECT 595.650 65.400 597.450 77.400 ;
        RECT 614.400 71.400 616.200 77.400 ;
        RECT 564.150 63.300 575.250 63.900 ;
        RECT 520.950 55.950 523.050 58.050 ;
        RECT 536.100 55.050 537.900 56.850 ;
        RECT 538.950 55.950 541.050 58.050 ;
        RECT 535.950 52.950 538.050 55.050 ;
        RECT 539.400 45.600 540.300 55.950 ;
        RECT 542.100 55.050 543.900 56.850 ;
        RECT 553.950 55.950 556.050 58.050 ;
        RECT 541.950 52.950 544.050 55.050 ;
        RECT 557.400 45.600 558.600 58.950 ;
        RECT 564.150 48.600 565.050 63.300 ;
        RECT 573.450 63.000 575.250 63.300 ;
        RECT 565.950 55.950 568.050 58.050 ;
        RECT 574.950 56.400 577.050 58.050 ;
        RECT 566.100 54.150 567.900 55.950 ;
        RECT 569.100 55.200 577.050 56.400 ;
        RECT 569.100 54.600 570.900 55.200 ;
        RECT 567.000 53.400 567.900 54.150 ;
        RECT 572.100 53.400 573.900 54.000 ;
        RECT 567.000 52.200 573.900 53.400 ;
        RECT 583.950 52.200 584.850 64.800 ;
        RECT 589.950 63.600 594.150 64.800 ;
        RECT 593.250 61.800 595.050 63.600 ;
        RECT 596.250 58.050 597.450 65.400 ;
        RECT 610.950 58.950 613.050 61.050 ;
        RECT 592.950 57.750 597.450 58.050 ;
        RECT 591.150 55.950 597.450 57.750 ;
        RECT 611.100 57.150 612.900 58.950 ;
        RECT 614.850 58.050 616.050 71.400 ;
        RECT 637.500 66.600 639.300 77.400 ;
        RECT 659.400 71.400 661.200 77.400 ;
        RECT 635.700 65.400 639.300 66.600 ;
        RECT 616.950 58.950 619.050 61.050 ;
        RECT 572.850 51.000 584.850 52.200 ;
        RECT 572.850 49.200 573.900 51.000 ;
        RECT 583.050 50.400 584.850 51.000 ;
        RECT 479.400 42.600 481.200 45.600 ;
        RECT 499.800 42.600 501.600 45.600 ;
        RECT 517.800 42.600 519.600 45.600 ;
        RECT 538.800 42.600 540.600 45.600 ;
        RECT 557.400 42.600 559.200 45.600 ;
        RECT 564.150 42.600 565.950 48.600 ;
        RECT 568.950 46.500 571.050 48.600 ;
        RECT 572.550 47.400 574.350 49.200 ;
        RECT 596.250 48.600 597.450 55.950 ;
        RECT 613.950 55.950 616.050 58.050 ;
        RECT 617.100 57.150 618.900 58.950 ;
        RECT 620.100 58.050 621.900 59.850 ;
        RECT 635.700 58.050 636.600 65.400 ;
        RECT 655.950 58.950 658.050 61.050 ;
        RECT 619.950 55.950 622.050 58.050 ;
        RECT 613.950 51.750 615.150 55.950 ;
        RECT 632.100 55.050 633.900 56.850 ;
        RECT 634.950 55.950 637.050 58.050 ;
        RECT 656.100 57.150 657.900 58.950 ;
        RECT 659.850 58.050 661.050 71.400 ;
        RECT 669.150 65.400 670.950 77.400 ;
        RECT 677.550 71.400 679.350 77.400 ;
        RECT 677.550 70.500 678.750 71.400 ;
        RECT 685.350 70.500 687.150 77.400 ;
        RECT 693.150 71.400 694.950 77.400 ;
        RECT 673.950 68.400 678.750 70.500 ;
        RECT 681.450 69.450 688.050 70.500 ;
        RECT 681.450 68.700 683.250 69.450 ;
        RECT 686.250 68.700 688.050 69.450 ;
        RECT 693.150 69.300 697.050 71.400 ;
        RECT 677.550 67.500 678.750 68.400 ;
        RECT 690.450 67.800 692.250 68.400 ;
        RECT 677.550 66.300 685.050 67.500 ;
        RECT 683.250 65.700 685.050 66.300 ;
        RECT 685.950 66.900 692.250 67.800 ;
        RECT 669.150 64.500 670.050 65.400 ;
        RECT 685.950 64.800 686.850 66.900 ;
        RECT 690.450 66.600 692.250 66.900 ;
        RECT 693.150 66.600 695.850 68.400 ;
        RECT 693.150 65.700 694.050 66.600 ;
        RECT 678.450 64.500 686.850 64.800 ;
        RECT 669.150 63.900 686.850 64.500 ;
        RECT 688.950 64.800 694.050 65.700 ;
        RECT 694.950 64.800 697.050 65.700 ;
        RECT 700.650 65.400 702.450 77.400 ;
        RECT 669.150 63.300 680.250 63.900 ;
        RECT 661.950 58.950 664.050 61.050 ;
        RECT 631.950 52.950 634.050 55.050 ;
        RECT 611.400 50.700 615.150 51.750 ;
        RECT 611.400 48.600 612.600 50.700 ;
        RECT 575.850 47.550 577.650 48.300 ;
        RECT 589.950 47.700 592.050 48.600 ;
        RECT 575.850 46.500 580.800 47.550 ;
        RECT 570.000 45.600 571.050 46.500 ;
        RECT 579.750 45.600 580.800 46.500 ;
        RECT 588.300 46.500 592.050 47.700 ;
        RECT 588.300 45.600 589.350 46.500 ;
        RECT 570.000 44.700 573.750 45.600 ;
        RECT 571.950 42.600 573.750 44.700 ;
        RECT 579.750 42.600 581.550 45.600 ;
        RECT 587.550 42.600 589.350 45.600 ;
        RECT 595.650 42.600 597.450 48.600 ;
        RECT 610.800 42.600 612.600 48.600 ;
        RECT 613.800 47.700 621.600 49.050 ;
        RECT 613.800 42.600 615.600 47.700 ;
        RECT 619.800 42.600 621.600 47.700 ;
        RECT 635.700 45.600 636.600 55.950 ;
        RECT 638.100 55.050 639.900 56.850 ;
        RECT 658.950 55.950 661.050 58.050 ;
        RECT 662.100 57.150 663.900 58.950 ;
        RECT 665.100 58.050 666.900 59.850 ;
        RECT 664.950 55.950 667.050 58.050 ;
        RECT 637.950 52.950 640.050 55.050 ;
        RECT 658.950 51.750 660.150 55.950 ;
        RECT 656.400 50.700 660.150 51.750 ;
        RECT 656.400 48.600 657.600 50.700 ;
        RECT 635.400 42.600 637.200 45.600 ;
        RECT 655.800 42.600 657.600 48.600 ;
        RECT 658.800 47.700 666.600 49.050 ;
        RECT 658.800 42.600 660.600 47.700 ;
        RECT 664.800 42.600 666.600 47.700 ;
        RECT 669.150 48.600 670.050 63.300 ;
        RECT 678.450 63.000 680.250 63.300 ;
        RECT 670.950 55.950 673.050 58.050 ;
        RECT 679.950 56.400 682.050 58.050 ;
        RECT 671.100 54.150 672.900 55.950 ;
        RECT 674.100 55.200 682.050 56.400 ;
        RECT 674.100 54.600 675.900 55.200 ;
        RECT 672.000 53.400 672.900 54.150 ;
        RECT 677.100 53.400 678.900 54.000 ;
        RECT 672.000 52.200 678.900 53.400 ;
        RECT 688.950 52.200 689.850 64.800 ;
        RECT 694.950 63.600 699.150 64.800 ;
        RECT 698.250 61.800 700.050 63.600 ;
        RECT 701.250 58.050 702.450 65.400 ;
        RECT 716.400 71.400 718.200 77.400 ;
        RECT 716.400 64.050 717.600 71.400 ;
        RECT 736.500 66.600 738.300 77.400 ;
        RECT 734.700 65.400 738.300 66.600 ;
        RECT 752.400 71.400 754.200 77.400 ;
        RECT 713.100 58.050 714.900 59.850 ;
        RECT 715.950 58.950 718.050 64.050 ;
        RECT 697.950 57.750 702.450 58.050 ;
        RECT 696.150 55.950 702.450 57.750 ;
        RECT 712.950 55.950 715.050 58.050 ;
        RECT 677.850 51.000 689.850 52.200 ;
        RECT 677.850 49.200 678.900 51.000 ;
        RECT 688.050 50.400 689.850 51.000 ;
        RECT 669.150 42.600 670.950 48.600 ;
        RECT 673.950 46.500 676.050 48.600 ;
        RECT 677.550 47.400 679.350 49.200 ;
        RECT 701.250 48.600 702.450 55.950 ;
        RECT 680.850 47.550 682.650 48.300 ;
        RECT 694.950 47.700 697.050 48.600 ;
        RECT 680.850 46.500 685.800 47.550 ;
        RECT 675.000 45.600 676.050 46.500 ;
        RECT 684.750 45.600 685.800 46.500 ;
        RECT 693.300 46.500 697.050 47.700 ;
        RECT 693.300 45.600 694.350 46.500 ;
        RECT 675.000 44.700 678.750 45.600 ;
        RECT 676.950 42.600 678.750 44.700 ;
        RECT 684.750 42.600 686.550 45.600 ;
        RECT 692.550 42.600 694.350 45.600 ;
        RECT 700.650 42.600 702.450 48.600 ;
        RECT 716.400 45.600 717.600 58.950 ;
        RECT 734.700 58.050 735.600 65.400 ;
        RECT 752.400 64.500 753.600 71.400 ;
        RECT 758.700 65.400 760.500 77.400 ;
        RECT 779.400 71.400 781.200 77.400 ;
        RECT 802.800 71.400 804.600 77.400 ;
        RECT 752.400 63.600 758.400 64.500 ;
        RECT 756.150 62.700 758.400 63.600 ;
        RECT 752.100 58.050 753.900 59.850 ;
        RECT 731.100 55.050 732.900 56.850 ;
        RECT 733.950 55.950 736.050 58.050 ;
        RECT 730.950 52.950 733.050 55.050 ;
        RECT 734.700 45.600 735.600 55.950 ;
        RECT 737.100 55.050 738.900 56.850 ;
        RECT 751.950 55.950 754.050 58.050 ;
        RECT 736.950 52.950 739.050 55.050 ;
        RECT 756.150 51.300 757.050 62.700 ;
        RECT 759.300 58.050 760.500 65.400 ;
        RECT 775.950 58.950 778.050 61.050 ;
        RECT 757.950 55.950 760.500 58.050 ;
        RECT 776.100 57.150 777.900 58.950 ;
        RECT 779.850 58.050 781.050 71.400 ;
        RECT 781.950 58.950 784.050 61.050 ;
        RECT 756.150 50.400 758.400 51.300 ;
        RECT 752.400 49.500 758.400 50.400 ;
        RECT 752.400 45.600 753.600 49.500 ;
        RECT 759.300 48.600 760.500 55.950 ;
        RECT 778.950 55.950 781.050 58.050 ;
        RECT 782.100 57.150 783.900 58.950 ;
        RECT 785.100 58.050 786.900 59.850 ;
        RECT 799.950 58.950 802.050 61.050 ;
        RECT 784.950 55.950 787.050 58.050 ;
        RECT 800.100 57.150 801.900 58.950 ;
        RECT 803.400 58.050 804.600 71.400 ;
        RECT 809.550 65.400 811.350 77.400 ;
        RECT 817.050 71.400 818.850 77.400 ;
        RECT 814.950 69.300 818.850 71.400 ;
        RECT 824.850 70.500 826.650 77.400 ;
        RECT 832.650 71.400 834.450 77.400 ;
        RECT 833.250 70.500 834.450 71.400 ;
        RECT 823.950 69.450 830.550 70.500 ;
        RECT 823.950 68.700 825.750 69.450 ;
        RECT 828.750 68.700 830.550 69.450 ;
        RECT 833.250 68.400 838.050 70.500 ;
        RECT 816.150 66.600 818.850 68.400 ;
        RECT 819.750 67.800 821.550 68.400 ;
        RECT 819.750 66.900 826.050 67.800 ;
        RECT 833.250 67.500 834.450 68.400 ;
        RECT 819.750 66.600 821.550 66.900 ;
        RECT 817.950 65.700 818.850 66.600 ;
        RECT 805.950 58.950 808.050 61.050 ;
        RECT 802.950 55.950 805.050 58.050 ;
        RECT 806.100 57.150 807.900 58.950 ;
        RECT 809.550 58.050 810.750 65.400 ;
        RECT 814.950 64.800 817.050 65.700 ;
        RECT 817.950 64.800 823.050 65.700 ;
        RECT 812.850 63.600 817.050 64.800 ;
        RECT 811.950 61.800 813.750 63.600 ;
        RECT 809.550 57.750 814.050 58.050 ;
        RECT 809.550 55.950 815.850 57.750 ;
        RECT 778.950 51.750 780.150 55.950 ;
        RECT 776.400 50.700 780.150 51.750 ;
        RECT 803.400 50.700 804.600 55.950 ;
        RECT 776.400 48.600 777.600 50.700 ;
        RECT 800.400 49.800 804.600 50.700 ;
        RECT 716.400 42.600 718.200 45.600 ;
        RECT 734.400 42.600 736.200 45.600 ;
        RECT 752.400 42.600 754.200 45.600 ;
        RECT 758.700 42.600 760.500 48.600 ;
        RECT 775.800 42.600 777.600 48.600 ;
        RECT 778.800 47.700 786.600 49.050 ;
        RECT 778.800 42.600 780.600 47.700 ;
        RECT 784.800 42.600 786.600 47.700 ;
        RECT 800.400 42.600 802.200 49.800 ;
        RECT 809.550 48.600 810.750 55.950 ;
        RECT 822.150 52.200 823.050 64.800 ;
        RECT 825.150 64.800 826.050 66.900 ;
        RECT 826.950 66.300 834.450 67.500 ;
        RECT 826.950 65.700 828.750 66.300 ;
        RECT 841.050 65.400 842.850 77.400 ;
        RECT 859.800 71.400 861.600 77.400 ;
        RECT 825.150 64.500 833.550 64.800 ;
        RECT 841.950 64.500 842.850 65.400 ;
        RECT 844.950 64.950 847.050 67.050 ;
        RECT 825.150 63.900 842.850 64.500 ;
        RECT 831.750 63.300 842.850 63.900 ;
        RECT 831.750 63.000 833.550 63.300 ;
        RECT 829.950 56.400 832.050 58.050 ;
        RECT 829.950 55.200 837.900 56.400 ;
        RECT 838.950 55.950 841.050 58.050 ;
        RECT 836.100 54.600 837.900 55.200 ;
        RECT 839.100 54.150 840.900 55.950 ;
        RECT 833.100 53.400 834.900 54.000 ;
        RECT 839.100 53.400 840.000 54.150 ;
        RECT 833.100 52.200 840.000 53.400 ;
        RECT 822.150 51.000 834.150 52.200 ;
        RECT 822.150 50.400 823.950 51.000 ;
        RECT 833.100 49.200 834.150 51.000 ;
        RECT 809.550 42.600 811.350 48.600 ;
        RECT 814.950 47.700 817.050 48.600 ;
        RECT 814.950 46.500 818.700 47.700 ;
        RECT 829.350 47.550 831.150 48.300 ;
        RECT 817.650 45.600 818.700 46.500 ;
        RECT 826.200 46.500 831.150 47.550 ;
        RECT 832.650 47.400 834.450 49.200 ;
        RECT 841.950 48.600 842.850 63.300 ;
        RECT 845.550 49.050 846.450 64.950 ;
        RECT 854.100 58.050 855.900 59.850 ;
        RECT 856.950 58.950 859.050 61.050 ;
        RECT 853.950 55.950 856.050 58.050 ;
        RECT 857.100 57.150 858.900 58.950 ;
        RECT 859.950 58.050 861.150 71.400 ;
        RECT 880.800 65.400 882.600 77.400 ;
        RECT 883.800 66.300 885.600 77.400 ;
        RECT 889.800 66.300 891.600 77.400 ;
        RECT 883.800 65.400 891.600 66.300 ;
        RECT 902.400 71.400 904.200 77.400 ;
        RECT 862.950 58.950 865.050 61.050 ;
        RECT 859.950 55.950 862.050 58.050 ;
        RECT 863.100 57.150 864.900 58.950 ;
        RECT 881.400 58.050 882.600 65.400 ;
        RECT 902.400 64.050 903.600 71.400 ;
        RECT 883.950 58.950 886.050 61.050 ;
        RECT 880.950 55.950 883.050 58.050 ;
        RECT 884.100 57.150 885.900 58.950 ;
        RECT 887.100 58.050 888.900 59.850 ;
        RECT 889.950 58.950 892.050 61.050 ;
        RECT 886.950 55.950 889.050 58.050 ;
        RECT 890.100 57.150 891.900 58.950 ;
        RECT 899.100 58.050 900.900 59.850 ;
        RECT 901.950 58.950 904.050 64.050 ;
        RECT 898.950 55.950 901.050 58.050 ;
        RECT 860.850 51.750 862.050 55.950 ;
        RECT 860.850 50.700 864.600 51.750 ;
        RECT 835.950 46.500 838.050 48.600 ;
        RECT 826.200 45.600 827.250 46.500 ;
        RECT 835.950 45.600 837.000 46.500 ;
        RECT 817.650 42.600 819.450 45.600 ;
        RECT 825.450 42.600 827.250 45.600 ;
        RECT 833.250 44.700 837.000 45.600 ;
        RECT 833.250 42.600 835.050 44.700 ;
        RECT 841.050 42.600 842.850 48.600 ;
        RECT 844.950 46.950 847.050 49.050 ;
        RECT 854.400 47.700 862.200 49.050 ;
        RECT 854.400 42.600 856.200 47.700 ;
        RECT 860.400 42.600 862.200 47.700 ;
        RECT 863.400 48.600 864.600 50.700 ;
        RECT 881.400 48.600 882.600 55.950 ;
        RECT 863.400 42.600 865.200 48.600 ;
        RECT 881.400 47.400 886.500 48.600 ;
        RECT 884.700 42.600 886.500 47.400 ;
        RECT 902.400 45.600 903.600 58.950 ;
        RECT 902.400 42.600 904.200 45.600 ;
        RECT 13.800 35.400 15.600 38.400 ;
        RECT 14.400 22.050 15.600 35.400 ;
        RECT 22.950 34.950 25.050 37.050 ;
        RECT 16.950 22.950 19.050 25.050 ;
        RECT 13.950 16.950 16.050 22.050 ;
        RECT 17.100 21.150 18.900 22.950 ;
        RECT 14.400 9.600 15.600 16.950 ;
        RECT 13.800 3.600 15.600 9.600 ;
        RECT 23.550 7.050 24.450 34.950 ;
        RECT 29.400 33.300 31.200 38.400 ;
        RECT 35.400 33.300 37.200 38.400 ;
        RECT 29.400 31.950 37.200 33.300 ;
        RECT 38.400 32.400 40.200 38.400 ;
        RECT 44.550 32.400 46.350 38.400 ;
        RECT 52.650 35.400 54.450 38.400 ;
        RECT 60.450 35.400 62.250 38.400 ;
        RECT 68.250 36.300 70.050 38.400 ;
        RECT 68.250 35.400 72.000 36.300 ;
        RECT 52.650 34.500 53.700 35.400 ;
        RECT 49.950 33.300 53.700 34.500 ;
        RECT 61.200 34.500 62.250 35.400 ;
        RECT 70.950 34.500 72.000 35.400 ;
        RECT 61.200 33.450 66.150 34.500 ;
        RECT 49.950 32.400 52.050 33.300 ;
        RECT 64.350 32.700 66.150 33.450 ;
        RECT 38.400 30.300 39.600 32.400 ;
        RECT 35.850 29.250 39.600 30.300 ;
        RECT 35.850 25.050 37.050 29.250 ;
        RECT 28.950 22.950 31.050 25.050 ;
        RECT 29.100 21.150 30.900 22.950 ;
        RECT 32.100 22.050 33.900 23.850 ;
        RECT 34.950 22.950 37.050 25.050 ;
        RECT 44.550 25.050 45.750 32.400 ;
        RECT 67.650 31.800 69.450 33.600 ;
        RECT 70.950 32.400 73.050 34.500 ;
        RECT 76.050 32.400 77.850 38.400 ;
        RECT 91.800 32.400 93.600 38.400 ;
        RECT 57.150 30.000 58.950 30.600 ;
        RECT 68.100 30.000 69.150 31.800 ;
        RECT 57.150 28.800 69.150 30.000 ;
        RECT 31.950 19.950 34.050 22.050 ;
        RECT 34.950 9.600 36.150 22.950 ;
        RECT 38.100 22.050 39.900 23.850 ;
        RECT 44.550 23.250 50.850 25.050 ;
        RECT 44.550 22.950 49.050 23.250 ;
        RECT 37.950 19.950 40.050 22.050 ;
        RECT 44.550 15.600 45.750 22.950 ;
        RECT 46.950 17.400 48.750 19.200 ;
        RECT 47.850 16.200 52.050 17.400 ;
        RECT 57.150 16.200 58.050 28.800 ;
        RECT 68.100 27.600 75.000 28.800 ;
        RECT 68.100 27.000 69.900 27.600 ;
        RECT 74.100 26.850 75.000 27.600 ;
        RECT 71.100 25.800 72.900 26.400 ;
        RECT 64.950 24.600 72.900 25.800 ;
        RECT 74.100 25.050 75.900 26.850 ;
        RECT 64.950 22.950 67.050 24.600 ;
        RECT 73.950 22.950 76.050 25.050 ;
        RECT 66.750 17.700 68.550 18.000 ;
        RECT 76.950 17.700 77.850 32.400 ;
        RECT 92.400 30.300 93.600 32.400 ;
        RECT 94.800 33.300 96.600 38.400 ;
        RECT 100.800 33.300 102.600 38.400 ;
        RECT 94.800 31.950 102.600 33.300 ;
        RECT 113.400 30.600 115.200 38.400 ;
        RECT 120.900 34.200 122.700 38.400 ;
        RECT 120.900 32.400 123.600 34.200 ;
        RECT 119.100 30.600 120.900 31.500 ;
        RECT 92.400 29.250 96.150 30.300 ;
        RECT 113.400 29.700 120.900 30.600 ;
        RECT 94.950 25.050 96.150 29.250 ;
        RECT 113.100 25.050 114.900 26.850 ;
        RECT 92.100 22.050 93.900 23.850 ;
        RECT 94.950 22.950 97.050 25.050 ;
        RECT 91.950 19.950 94.050 22.050 ;
        RECT 66.750 17.100 77.850 17.700 ;
        RECT 22.950 4.950 25.050 7.050 ;
        RECT 34.800 3.600 36.600 9.600 ;
        RECT 44.550 3.600 46.350 15.600 ;
        RECT 49.950 15.300 52.050 16.200 ;
        RECT 52.950 15.300 58.050 16.200 ;
        RECT 60.150 16.500 77.850 17.100 ;
        RECT 60.150 16.200 68.550 16.500 ;
        RECT 52.950 14.400 53.850 15.300 ;
        RECT 51.150 12.600 53.850 14.400 ;
        RECT 54.750 14.100 56.550 14.400 ;
        RECT 60.150 14.100 61.050 16.200 ;
        RECT 76.950 15.600 77.850 16.500 ;
        RECT 54.750 13.200 61.050 14.100 ;
        RECT 61.950 14.700 63.750 15.300 ;
        RECT 61.950 13.500 69.450 14.700 ;
        RECT 54.750 12.600 56.550 13.200 ;
        RECT 68.250 12.600 69.450 13.500 ;
        RECT 49.950 9.600 53.850 11.700 ;
        RECT 58.950 11.550 60.750 12.300 ;
        RECT 63.750 11.550 65.550 12.300 ;
        RECT 58.950 10.500 65.550 11.550 ;
        RECT 68.250 10.500 73.050 12.600 ;
        RECT 52.050 3.600 53.850 9.600 ;
        RECT 59.850 3.600 61.650 10.500 ;
        RECT 68.250 9.600 69.450 10.500 ;
        RECT 67.650 3.600 69.450 9.600 ;
        RECT 76.050 3.600 77.850 15.600 ;
        RECT 95.850 9.600 97.050 22.950 ;
        RECT 98.100 22.050 99.900 23.850 ;
        RECT 100.950 22.950 103.050 25.050 ;
        RECT 112.950 22.950 115.050 25.050 ;
        RECT 97.950 19.950 100.050 22.050 ;
        RECT 101.100 21.150 102.900 22.950 ;
        RECT 116.400 9.600 117.300 29.700 ;
        RECT 122.700 25.050 123.600 32.400 ;
        RECT 137.400 33.300 139.200 38.400 ;
        RECT 143.400 33.300 145.200 38.400 ;
        RECT 137.400 31.950 145.200 33.300 ;
        RECT 146.400 32.400 148.200 38.400 ;
        RECT 153.150 32.400 154.950 38.400 ;
        RECT 160.950 36.300 162.750 38.400 ;
        RECT 159.000 35.400 162.750 36.300 ;
        RECT 168.750 35.400 170.550 38.400 ;
        RECT 176.550 35.400 178.350 38.400 ;
        RECT 159.000 34.500 160.050 35.400 ;
        RECT 168.750 34.500 169.800 35.400 ;
        RECT 157.950 32.400 160.050 34.500 ;
        RECT 146.400 30.300 147.600 32.400 ;
        RECT 143.850 29.250 147.600 30.300 ;
        RECT 143.850 25.050 145.050 29.250 ;
        RECT 118.950 22.950 121.050 25.050 ;
        RECT 121.950 22.950 124.050 25.050 ;
        RECT 136.950 22.950 139.050 25.050 ;
        RECT 119.100 21.150 120.900 22.950 ;
        RECT 122.700 15.600 123.600 22.950 ;
        RECT 137.100 21.150 138.900 22.950 ;
        RECT 140.100 22.050 141.900 23.850 ;
        RECT 142.950 22.950 145.050 25.050 ;
        RECT 139.950 19.950 142.050 22.050 ;
        RECT 95.400 3.600 97.200 9.600 ;
        RECT 116.400 3.600 118.200 9.600 ;
        RECT 122.700 3.600 124.500 15.600 ;
        RECT 142.950 9.600 144.150 22.950 ;
        RECT 146.100 22.050 147.900 23.850 ;
        RECT 145.950 19.950 148.050 22.050 ;
        RECT 153.150 17.700 154.050 32.400 ;
        RECT 161.550 31.800 163.350 33.600 ;
        RECT 164.850 33.450 169.800 34.500 ;
        RECT 177.300 34.500 178.350 35.400 ;
        RECT 164.850 32.700 166.650 33.450 ;
        RECT 177.300 33.300 181.050 34.500 ;
        RECT 178.950 32.400 181.050 33.300 ;
        RECT 184.650 32.400 186.450 38.400 ;
        RECT 161.850 30.000 162.900 31.800 ;
        RECT 172.050 30.000 173.850 30.600 ;
        RECT 161.850 28.800 173.850 30.000 ;
        RECT 156.000 27.600 162.900 28.800 ;
        RECT 156.000 26.850 156.900 27.600 ;
        RECT 161.100 27.000 162.900 27.600 ;
        RECT 155.100 25.050 156.900 26.850 ;
        RECT 158.100 25.800 159.900 26.400 ;
        RECT 154.950 22.950 157.050 25.050 ;
        RECT 158.100 24.600 166.050 25.800 ;
        RECT 163.950 22.950 166.050 24.600 ;
        RECT 162.450 17.700 164.250 18.000 ;
        RECT 153.150 17.100 164.250 17.700 ;
        RECT 153.150 16.500 170.850 17.100 ;
        RECT 153.150 15.600 154.050 16.500 ;
        RECT 162.450 16.200 170.850 16.500 ;
        RECT 142.800 3.600 144.600 9.600 ;
        RECT 153.150 3.600 154.950 15.600 ;
        RECT 167.250 14.700 169.050 15.300 ;
        RECT 161.550 13.500 169.050 14.700 ;
        RECT 169.950 14.100 170.850 16.200 ;
        RECT 172.950 16.200 173.850 28.800 ;
        RECT 185.250 25.050 186.450 32.400 ;
        RECT 202.800 31.200 204.600 38.400 ;
        RECT 218.400 33.300 220.200 38.400 ;
        RECT 224.400 33.300 226.200 38.400 ;
        RECT 218.400 31.950 226.200 33.300 ;
        RECT 227.400 32.400 229.200 38.400 ;
        RECT 234.150 32.400 235.950 38.400 ;
        RECT 241.950 36.300 243.750 38.400 ;
        RECT 240.000 35.400 243.750 36.300 ;
        RECT 249.750 35.400 251.550 38.400 ;
        RECT 257.550 35.400 259.350 38.400 ;
        RECT 240.000 34.500 241.050 35.400 ;
        RECT 249.750 34.500 250.800 35.400 ;
        RECT 238.950 32.400 241.050 34.500 ;
        RECT 200.400 30.300 204.600 31.200 ;
        RECT 227.400 30.300 228.600 32.400 ;
        RECT 200.400 25.050 201.600 30.300 ;
        RECT 224.850 29.250 228.600 30.300 ;
        RECT 224.850 25.050 226.050 29.250 ;
        RECT 180.150 23.250 186.450 25.050 ;
        RECT 181.950 22.950 186.450 23.250 ;
        RECT 182.250 17.400 184.050 19.200 ;
        RECT 178.950 16.200 183.150 17.400 ;
        RECT 172.950 15.300 178.050 16.200 ;
        RECT 178.950 15.300 181.050 16.200 ;
        RECT 185.250 15.600 186.450 22.950 ;
        RECT 197.100 22.050 198.900 23.850 ;
        RECT 199.950 22.950 202.050 25.050 ;
        RECT 196.950 19.950 199.050 22.050 ;
        RECT 177.150 14.400 178.050 15.300 ;
        RECT 174.450 14.100 176.250 14.400 ;
        RECT 161.550 12.600 162.750 13.500 ;
        RECT 169.950 13.200 176.250 14.100 ;
        RECT 174.450 12.600 176.250 13.200 ;
        RECT 177.150 12.600 179.850 14.400 ;
        RECT 157.950 10.500 162.750 12.600 ;
        RECT 165.450 11.550 167.250 12.300 ;
        RECT 170.250 11.550 172.050 12.300 ;
        RECT 165.450 10.500 172.050 11.550 ;
        RECT 161.550 9.600 162.750 10.500 ;
        RECT 161.550 3.600 163.350 9.600 ;
        RECT 169.350 3.600 171.150 10.500 ;
        RECT 177.150 9.600 181.050 11.700 ;
        RECT 177.150 3.600 178.950 9.600 ;
        RECT 184.650 3.600 186.450 15.600 ;
        RECT 200.400 9.600 201.600 22.950 ;
        RECT 203.100 22.050 204.900 23.850 ;
        RECT 217.950 22.950 220.050 25.050 ;
        RECT 202.950 19.950 205.050 22.050 ;
        RECT 218.100 21.150 219.900 22.950 ;
        RECT 221.100 22.050 222.900 23.850 ;
        RECT 223.950 22.950 226.050 25.050 ;
        RECT 220.950 19.950 223.050 22.050 ;
        RECT 223.950 9.600 225.150 22.950 ;
        RECT 227.100 22.050 228.900 23.850 ;
        RECT 226.950 19.950 229.050 22.050 ;
        RECT 234.150 17.700 235.050 32.400 ;
        RECT 242.550 31.800 244.350 33.600 ;
        RECT 245.850 33.450 250.800 34.500 ;
        RECT 258.300 34.500 259.350 35.400 ;
        RECT 245.850 32.700 247.650 33.450 ;
        RECT 258.300 33.300 262.050 34.500 ;
        RECT 259.950 32.400 262.050 33.300 ;
        RECT 265.650 32.400 267.450 38.400 ;
        RECT 242.850 30.000 243.900 31.800 ;
        RECT 253.050 30.000 254.850 30.600 ;
        RECT 242.850 28.800 254.850 30.000 ;
        RECT 237.000 27.600 243.900 28.800 ;
        RECT 237.000 26.850 237.900 27.600 ;
        RECT 242.100 27.000 243.900 27.600 ;
        RECT 236.100 25.050 237.900 26.850 ;
        RECT 239.100 25.800 240.900 26.400 ;
        RECT 235.950 22.950 238.050 25.050 ;
        RECT 239.100 24.600 247.050 25.800 ;
        RECT 244.950 22.950 247.050 24.600 ;
        RECT 243.450 17.700 245.250 18.000 ;
        RECT 234.150 17.100 245.250 17.700 ;
        RECT 234.150 16.500 251.850 17.100 ;
        RECT 234.150 15.600 235.050 16.500 ;
        RECT 243.450 16.200 251.850 16.500 ;
        RECT 200.400 3.600 202.200 9.600 ;
        RECT 223.800 3.600 225.600 9.600 ;
        RECT 234.150 3.600 235.950 15.600 ;
        RECT 248.250 14.700 250.050 15.300 ;
        RECT 242.550 13.500 250.050 14.700 ;
        RECT 250.950 14.100 251.850 16.200 ;
        RECT 253.950 16.200 254.850 28.800 ;
        RECT 266.250 25.050 267.450 32.400 ;
        RECT 283.800 31.200 285.600 38.400 ;
        RECT 304.200 32.400 306.000 38.400 ;
        RECT 281.400 30.300 285.600 31.200 ;
        RECT 268.950 25.950 271.050 28.050 ;
        RECT 261.150 23.250 267.450 25.050 ;
        RECT 262.950 22.950 267.450 23.250 ;
        RECT 263.250 17.400 265.050 19.200 ;
        RECT 259.950 16.200 264.150 17.400 ;
        RECT 253.950 15.300 259.050 16.200 ;
        RECT 259.950 15.300 262.050 16.200 ;
        RECT 266.250 15.600 267.450 22.950 ;
        RECT 258.150 14.400 259.050 15.300 ;
        RECT 255.450 14.100 257.250 14.400 ;
        RECT 242.550 12.600 243.750 13.500 ;
        RECT 250.950 13.200 257.250 14.100 ;
        RECT 255.450 12.600 257.250 13.200 ;
        RECT 258.150 12.600 260.850 14.400 ;
        RECT 238.950 10.500 243.750 12.600 ;
        RECT 246.450 11.550 248.250 12.300 ;
        RECT 251.250 11.550 253.050 12.300 ;
        RECT 246.450 10.500 253.050 11.550 ;
        RECT 242.550 9.600 243.750 10.500 ;
        RECT 242.550 3.600 244.350 9.600 ;
        RECT 250.350 3.600 252.150 10.500 ;
        RECT 258.150 9.600 262.050 11.700 ;
        RECT 258.150 3.600 259.950 9.600 ;
        RECT 265.650 3.600 267.450 15.600 ;
        RECT 269.550 7.050 270.450 25.950 ;
        RECT 281.400 25.050 282.600 30.300 ;
        RECT 299.100 25.050 300.900 26.850 ;
        RECT 301.950 25.950 304.050 28.050 ;
        RECT 278.100 22.050 279.900 23.850 ;
        RECT 280.950 22.950 283.050 25.050 ;
        RECT 277.950 19.950 280.050 22.050 ;
        RECT 281.400 9.600 282.600 22.950 ;
        RECT 284.100 22.050 285.900 23.850 ;
        RECT 298.950 22.950 301.050 25.050 ;
        RECT 302.100 24.150 303.900 25.950 ;
        RECT 304.950 25.050 306.000 32.400 ;
        RECT 336.000 32.400 337.800 38.400 ;
        RECT 316.950 28.950 319.050 31.050 ;
        RECT 307.950 25.950 310.050 28.050 ;
        RECT 304.950 22.950 307.050 25.050 ;
        RECT 308.100 24.150 309.900 25.950 ;
        RECT 311.100 25.050 312.900 26.850 ;
        RECT 310.950 22.950 313.050 25.050 ;
        RECT 283.950 19.950 286.050 22.050 ;
        RECT 305.100 17.400 306.000 22.950 ;
        RECT 305.100 16.500 310.200 17.400 ;
        RECT 299.400 14.400 307.200 15.300 ;
        RECT 268.950 4.950 271.050 7.050 ;
        RECT 281.400 3.600 283.200 9.600 ;
        RECT 299.400 3.600 301.200 14.400 ;
        RECT 305.400 4.500 307.200 14.400 ;
        RECT 308.400 5.400 310.200 16.500 ;
        RECT 311.400 4.500 313.200 15.600 ;
        RECT 317.550 13.050 318.450 28.950 ;
        RECT 329.100 25.050 330.900 26.850 ;
        RECT 331.950 25.950 334.050 28.050 ;
        RECT 328.950 22.950 331.050 25.050 ;
        RECT 332.100 24.150 333.900 25.950 ;
        RECT 336.000 25.050 337.050 32.400 ;
        RECT 356.400 31.200 358.200 38.400 ;
        RECT 376.800 32.400 378.600 38.400 ;
        RECT 356.400 30.300 360.600 31.200 ;
        RECT 337.950 25.950 340.050 28.050 ;
        RECT 334.950 22.950 337.050 25.050 ;
        RECT 338.100 24.150 339.900 25.950 ;
        RECT 341.100 25.050 342.900 26.850 ;
        RECT 359.400 25.050 360.600 30.300 ;
        RECT 377.400 30.300 378.600 32.400 ;
        RECT 379.800 33.300 381.600 38.400 ;
        RECT 385.800 33.300 387.600 38.400 ;
        RECT 379.800 31.950 387.600 33.300 ;
        RECT 389.550 32.400 391.350 38.400 ;
        RECT 397.650 35.400 399.450 38.400 ;
        RECT 405.450 35.400 407.250 38.400 ;
        RECT 413.250 36.300 415.050 38.400 ;
        RECT 413.250 35.400 417.000 36.300 ;
        RECT 397.650 34.500 398.700 35.400 ;
        RECT 394.950 33.300 398.700 34.500 ;
        RECT 406.200 34.500 407.250 35.400 ;
        RECT 415.950 34.500 417.000 35.400 ;
        RECT 406.200 33.450 411.150 34.500 ;
        RECT 394.950 32.400 397.050 33.300 ;
        RECT 409.350 32.700 411.150 33.450 ;
        RECT 377.400 29.250 381.150 30.300 ;
        RECT 379.950 25.050 381.150 29.250 ;
        RECT 389.550 25.050 390.750 32.400 ;
        RECT 412.650 31.800 414.450 33.600 ;
        RECT 415.950 32.400 418.050 34.500 ;
        RECT 421.050 32.400 422.850 38.400 ;
        RECT 402.150 30.000 403.950 30.600 ;
        RECT 413.100 30.000 414.150 31.800 ;
        RECT 402.150 28.800 414.150 30.000 ;
        RECT 340.950 22.950 343.050 25.050 ;
        RECT 336.000 17.400 336.900 22.950 ;
        RECT 356.100 22.050 357.900 23.850 ;
        RECT 358.950 22.950 361.050 25.050 ;
        RECT 355.950 19.950 358.050 22.050 ;
        RECT 331.800 16.500 336.900 17.400 ;
        RECT 316.950 10.950 319.050 13.050 ;
        RECT 305.400 3.600 313.200 4.500 ;
        RECT 328.800 4.500 330.600 15.600 ;
        RECT 331.800 5.400 333.600 16.500 ;
        RECT 334.800 14.400 342.600 15.300 ;
        RECT 334.800 4.500 336.600 14.400 ;
        RECT 328.800 3.600 336.600 4.500 ;
        RECT 340.800 3.600 342.600 14.400 ;
        RECT 359.400 9.600 360.600 22.950 ;
        RECT 362.100 22.050 363.900 23.850 ;
        RECT 377.100 22.050 378.900 23.850 ;
        RECT 379.950 22.950 382.050 25.050 ;
        RECT 361.950 19.950 364.050 22.050 ;
        RECT 376.950 19.950 379.050 22.050 ;
        RECT 380.850 9.600 382.050 22.950 ;
        RECT 383.100 22.050 384.900 23.850 ;
        RECT 385.950 22.950 388.050 25.050 ;
        RECT 389.550 23.250 395.850 25.050 ;
        RECT 389.550 22.950 394.050 23.250 ;
        RECT 382.950 19.950 385.050 22.050 ;
        RECT 386.100 21.150 387.900 22.950 ;
        RECT 389.550 15.600 390.750 22.950 ;
        RECT 391.950 17.400 393.750 19.200 ;
        RECT 392.850 16.200 397.050 17.400 ;
        RECT 402.150 16.200 403.050 28.800 ;
        RECT 413.100 27.600 420.000 28.800 ;
        RECT 413.100 27.000 414.900 27.600 ;
        RECT 419.100 26.850 420.000 27.600 ;
        RECT 416.100 25.800 417.900 26.400 ;
        RECT 409.950 24.600 417.900 25.800 ;
        RECT 419.100 25.050 420.900 26.850 ;
        RECT 409.950 22.950 412.050 24.600 ;
        RECT 418.950 22.950 421.050 25.050 ;
        RECT 411.750 17.700 413.550 18.000 ;
        RECT 421.950 17.700 422.850 32.400 ;
        RECT 437.400 35.400 439.200 38.400 ;
        RECT 433.950 22.950 436.050 25.050 ;
        RECT 434.100 21.150 435.900 22.950 ;
        RECT 437.400 22.050 438.600 35.400 ;
        RECT 442.950 34.950 445.050 37.050 ;
        RECT 411.750 17.100 422.850 17.700 ;
        RECT 358.800 3.600 360.600 9.600 ;
        RECT 380.400 3.600 382.200 9.600 ;
        RECT 389.550 3.600 391.350 15.600 ;
        RECT 394.950 15.300 397.050 16.200 ;
        RECT 397.950 15.300 403.050 16.200 ;
        RECT 405.150 16.500 422.850 17.100 ;
        RECT 436.950 16.950 439.050 22.050 ;
        RECT 443.550 19.050 444.450 34.950 ;
        RECT 462.000 32.400 463.800 38.400 ;
        RECT 471.150 32.400 472.950 38.400 ;
        RECT 478.950 36.300 480.750 38.400 ;
        RECT 477.000 35.400 480.750 36.300 ;
        RECT 486.750 35.400 488.550 38.400 ;
        RECT 494.550 35.400 496.350 38.400 ;
        RECT 477.000 34.500 478.050 35.400 ;
        RECT 486.750 34.500 487.800 35.400 ;
        RECT 475.950 32.400 478.050 34.500 ;
        RECT 455.100 25.050 456.900 26.850 ;
        RECT 457.950 25.950 460.050 28.050 ;
        RECT 454.950 22.950 457.050 25.050 ;
        RECT 458.100 24.150 459.900 25.950 ;
        RECT 462.000 25.050 463.050 32.400 ;
        RECT 463.950 25.950 466.050 28.050 ;
        RECT 460.950 22.950 463.050 25.050 ;
        RECT 464.100 24.150 465.900 25.950 ;
        RECT 467.100 25.050 468.900 26.850 ;
        RECT 466.950 22.950 469.050 25.050 ;
        RECT 442.950 16.950 445.050 19.050 ;
        RECT 462.000 17.400 462.900 22.950 ;
        RECT 405.150 16.200 413.550 16.500 ;
        RECT 397.950 14.400 398.850 15.300 ;
        RECT 396.150 12.600 398.850 14.400 ;
        RECT 399.750 14.100 401.550 14.400 ;
        RECT 405.150 14.100 406.050 16.200 ;
        RECT 421.950 15.600 422.850 16.500 ;
        RECT 399.750 13.200 406.050 14.100 ;
        RECT 406.950 14.700 408.750 15.300 ;
        RECT 406.950 13.500 414.450 14.700 ;
        RECT 399.750 12.600 401.550 13.200 ;
        RECT 413.250 12.600 414.450 13.500 ;
        RECT 394.950 9.600 398.850 11.700 ;
        RECT 403.950 11.550 405.750 12.300 ;
        RECT 408.750 11.550 410.550 12.300 ;
        RECT 403.950 10.500 410.550 11.550 ;
        RECT 413.250 10.500 418.050 12.600 ;
        RECT 397.050 3.600 398.850 9.600 ;
        RECT 404.850 3.600 406.650 10.500 ;
        RECT 413.250 9.600 414.450 10.500 ;
        RECT 412.650 3.600 414.450 9.600 ;
        RECT 421.050 3.600 422.850 15.600 ;
        RECT 437.400 9.600 438.600 16.950 ;
        RECT 457.800 16.500 462.900 17.400 ;
        RECT 471.150 17.700 472.050 32.400 ;
        RECT 479.550 31.800 481.350 33.600 ;
        RECT 482.850 33.450 487.800 34.500 ;
        RECT 495.300 34.500 496.350 35.400 ;
        RECT 482.850 32.700 484.650 33.450 ;
        RECT 495.300 33.300 499.050 34.500 ;
        RECT 496.950 32.400 499.050 33.300 ;
        RECT 502.650 32.400 504.450 38.400 ;
        RECT 479.850 30.000 480.900 31.800 ;
        RECT 490.050 30.000 491.850 30.600 ;
        RECT 479.850 28.800 491.850 30.000 ;
        RECT 474.000 27.600 480.900 28.800 ;
        RECT 474.000 26.850 474.900 27.600 ;
        RECT 479.100 27.000 480.900 27.600 ;
        RECT 473.100 25.050 474.900 26.850 ;
        RECT 476.100 25.800 477.900 26.400 ;
        RECT 472.950 22.950 475.050 25.050 ;
        RECT 476.100 24.600 484.050 25.800 ;
        RECT 481.950 22.950 484.050 24.600 ;
        RECT 480.450 17.700 482.250 18.000 ;
        RECT 471.150 17.100 482.250 17.700 ;
        RECT 471.150 16.500 488.850 17.100 ;
        RECT 437.400 3.600 439.200 9.600 ;
        RECT 454.800 4.500 456.600 15.600 ;
        RECT 457.800 5.400 459.600 16.500 ;
        RECT 471.150 15.600 472.050 16.500 ;
        RECT 480.450 16.200 488.850 16.500 ;
        RECT 460.800 14.400 468.600 15.300 ;
        RECT 460.800 4.500 462.600 14.400 ;
        RECT 454.800 3.600 462.600 4.500 ;
        RECT 466.800 3.600 468.600 14.400 ;
        RECT 471.150 3.600 472.950 15.600 ;
        RECT 485.250 14.700 487.050 15.300 ;
        RECT 479.550 13.500 487.050 14.700 ;
        RECT 487.950 14.100 488.850 16.200 ;
        RECT 490.950 16.200 491.850 28.800 ;
        RECT 503.250 25.050 504.450 32.400 ;
        RECT 518.400 35.400 520.200 38.400 ;
        RECT 498.150 23.250 504.450 25.050 ;
        RECT 499.950 22.950 504.450 23.250 ;
        RECT 514.950 22.950 517.050 25.050 ;
        RECT 500.250 17.400 502.050 19.200 ;
        RECT 496.950 16.200 501.150 17.400 ;
        RECT 490.950 15.300 496.050 16.200 ;
        RECT 496.950 15.300 499.050 16.200 ;
        RECT 503.250 15.600 504.450 22.950 ;
        RECT 515.100 21.150 516.900 22.950 ;
        RECT 518.400 22.050 519.600 35.400 ;
        RECT 536.400 31.200 538.200 38.400 ;
        RECT 556.800 32.400 558.600 38.400 ;
        RECT 536.400 30.300 540.600 31.200 ;
        RECT 539.400 25.050 540.600 30.300 ;
        RECT 557.400 30.300 558.600 32.400 ;
        RECT 559.800 33.300 561.600 38.400 ;
        RECT 565.800 33.300 567.600 38.400 ;
        RECT 559.800 31.950 567.600 33.300 ;
        RECT 580.800 32.400 582.600 38.400 ;
        RECT 581.400 30.300 582.600 32.400 ;
        RECT 583.800 33.300 585.600 38.400 ;
        RECT 589.800 33.300 591.600 38.400 ;
        RECT 583.800 31.950 591.600 33.300 ;
        RECT 605.400 35.400 607.200 38.400 ;
        RECT 557.400 29.250 561.150 30.300 ;
        RECT 581.400 29.250 585.150 30.300 ;
        RECT 559.950 25.050 561.150 29.250 ;
        RECT 583.950 25.050 585.150 29.250 ;
        RECT 536.100 22.050 537.900 23.850 ;
        RECT 538.950 22.950 541.050 25.050 ;
        RECT 517.950 16.950 520.050 22.050 ;
        RECT 535.950 19.950 538.050 22.050 ;
        RECT 495.150 14.400 496.050 15.300 ;
        RECT 492.450 14.100 494.250 14.400 ;
        RECT 479.550 12.600 480.750 13.500 ;
        RECT 487.950 13.200 494.250 14.100 ;
        RECT 492.450 12.600 494.250 13.200 ;
        RECT 495.150 12.600 497.850 14.400 ;
        RECT 475.950 10.500 480.750 12.600 ;
        RECT 483.450 11.550 485.250 12.300 ;
        RECT 488.250 11.550 490.050 12.300 ;
        RECT 483.450 10.500 490.050 11.550 ;
        RECT 479.550 9.600 480.750 10.500 ;
        RECT 479.550 3.600 481.350 9.600 ;
        RECT 487.350 3.600 489.150 10.500 ;
        RECT 495.150 9.600 499.050 11.700 ;
        RECT 495.150 3.600 496.950 9.600 ;
        RECT 502.650 3.600 504.450 15.600 ;
        RECT 518.400 9.600 519.600 16.950 ;
        RECT 539.400 9.600 540.600 22.950 ;
        RECT 542.100 22.050 543.900 23.850 ;
        RECT 557.100 22.050 558.900 23.850 ;
        RECT 559.950 22.950 562.050 25.050 ;
        RECT 541.950 19.950 544.050 22.050 ;
        RECT 556.950 19.950 559.050 22.050 ;
        RECT 560.850 9.600 562.050 22.950 ;
        RECT 563.100 22.050 564.900 23.850 ;
        RECT 565.950 22.950 568.050 25.050 ;
        RECT 562.950 19.950 565.050 22.050 ;
        RECT 566.100 21.150 567.900 22.950 ;
        RECT 581.100 22.050 582.900 23.850 ;
        RECT 583.950 22.950 586.050 25.050 ;
        RECT 580.950 19.950 583.050 22.050 ;
        RECT 584.850 9.600 586.050 22.950 ;
        RECT 587.100 22.050 588.900 23.850 ;
        RECT 589.950 22.950 592.050 25.050 ;
        RECT 601.950 22.950 604.050 25.050 ;
        RECT 586.950 19.950 589.050 22.050 ;
        RECT 590.100 21.150 591.900 22.950 ;
        RECT 602.100 21.150 603.900 22.950 ;
        RECT 605.400 22.050 606.600 35.400 ;
        RECT 622.800 32.400 624.600 38.400 ;
        RECT 623.400 30.300 624.600 32.400 ;
        RECT 625.800 33.300 627.600 38.400 ;
        RECT 631.800 33.300 633.600 38.400 ;
        RECT 625.800 31.950 633.600 33.300 ;
        RECT 644.400 35.400 646.200 38.400 ;
        RECT 644.400 31.500 645.600 35.400 ;
        RECT 650.700 32.400 652.500 38.400 ;
        RECT 644.400 30.600 650.400 31.500 ;
        RECT 623.400 29.250 627.150 30.300 ;
        RECT 625.950 25.050 627.150 29.250 ;
        RECT 648.150 29.700 650.400 30.600 ;
        RECT 623.100 22.050 624.900 23.850 ;
        RECT 625.950 22.950 628.050 25.050 ;
        RECT 604.950 16.950 607.050 22.050 ;
        RECT 622.950 19.950 625.050 22.050 ;
        RECT 605.400 9.600 606.600 16.950 ;
        RECT 626.850 9.600 628.050 22.950 ;
        RECT 629.100 22.050 630.900 23.850 ;
        RECT 631.950 22.950 634.050 25.050 ;
        RECT 643.950 22.950 646.050 25.050 ;
        RECT 628.950 19.950 631.050 22.050 ;
        RECT 632.100 21.150 633.900 22.950 ;
        RECT 644.100 21.150 645.900 22.950 ;
        RECT 648.150 18.300 649.050 29.700 ;
        RECT 651.300 25.050 652.500 32.400 ;
        RECT 665.400 35.400 667.200 38.400 ;
        RECT 665.400 31.500 666.600 35.400 ;
        RECT 671.700 32.400 673.500 38.400 ;
        RECT 665.400 30.600 671.400 31.500 ;
        RECT 669.150 29.700 671.400 30.600 ;
        RECT 649.950 22.950 652.500 25.050 ;
        RECT 664.950 22.950 667.050 25.050 ;
        RECT 648.150 17.400 650.400 18.300 ;
        RECT 644.400 16.500 650.400 17.400 ;
        RECT 644.400 9.600 645.600 16.500 ;
        RECT 651.300 15.600 652.500 22.950 ;
        RECT 665.100 21.150 666.900 22.950 ;
        RECT 669.150 18.300 670.050 29.700 ;
        RECT 672.300 25.050 673.500 32.400 ;
        RECT 686.400 35.400 688.200 38.400 ;
        RECT 686.400 31.500 687.600 35.400 ;
        RECT 692.700 32.400 694.500 38.400 ;
        RECT 686.400 30.600 692.400 31.500 ;
        RECT 690.150 29.700 692.400 30.600 ;
        RECT 670.950 22.950 673.500 25.050 ;
        RECT 685.950 22.950 688.050 25.050 ;
        RECT 669.150 17.400 671.400 18.300 ;
        RECT 518.400 3.600 520.200 9.600 ;
        RECT 538.800 3.600 540.600 9.600 ;
        RECT 560.400 3.600 562.200 9.600 ;
        RECT 584.400 3.600 586.200 9.600 ;
        RECT 605.400 3.600 607.200 9.600 ;
        RECT 626.400 3.600 628.200 9.600 ;
        RECT 644.400 3.600 646.200 9.600 ;
        RECT 650.700 3.600 652.500 15.600 ;
        RECT 665.400 16.500 671.400 17.400 ;
        RECT 665.400 9.600 666.600 16.500 ;
        RECT 672.300 15.600 673.500 22.950 ;
        RECT 686.100 21.150 687.900 22.950 ;
        RECT 690.150 18.300 691.050 29.700 ;
        RECT 693.300 25.050 694.500 32.400 ;
        RECT 707.400 35.400 709.200 38.400 ;
        RECT 707.400 31.500 708.600 35.400 ;
        RECT 713.700 32.400 715.500 38.400 ;
        RECT 707.400 30.600 713.400 31.500 ;
        RECT 711.150 29.700 713.400 30.600 ;
        RECT 691.950 22.950 694.500 25.050 ;
        RECT 706.950 22.950 709.050 25.050 ;
        RECT 690.150 17.400 692.400 18.300 ;
        RECT 665.400 3.600 667.200 9.600 ;
        RECT 671.700 3.600 673.500 15.600 ;
        RECT 686.400 16.500 692.400 17.400 ;
        RECT 686.400 9.600 687.600 16.500 ;
        RECT 693.300 15.600 694.500 22.950 ;
        RECT 707.100 21.150 708.900 22.950 ;
        RECT 711.150 18.300 712.050 29.700 ;
        RECT 714.300 25.050 715.500 32.400 ;
        RECT 731.400 31.200 733.200 38.400 ;
        RECT 751.800 32.400 753.600 38.400 ;
        RECT 731.400 30.300 735.600 31.200 ;
        RECT 734.400 25.050 735.600 30.300 ;
        RECT 752.400 30.300 753.600 32.400 ;
        RECT 754.800 33.300 756.600 38.400 ;
        RECT 760.800 33.300 762.600 38.400 ;
        RECT 766.800 34.950 768.900 37.050 ;
        RECT 754.800 31.950 762.600 33.300 ;
        RECT 752.400 29.250 756.150 30.300 ;
        RECT 754.950 25.050 756.150 29.250 ;
        RECT 712.950 22.950 715.500 25.050 ;
        RECT 711.150 17.400 713.400 18.300 ;
        RECT 686.400 3.600 688.200 9.600 ;
        RECT 692.700 3.600 694.500 15.600 ;
        RECT 707.400 16.500 713.400 17.400 ;
        RECT 707.400 9.600 708.600 16.500 ;
        RECT 714.300 15.600 715.500 22.950 ;
        RECT 731.100 22.050 732.900 23.850 ;
        RECT 733.950 22.950 736.050 25.050 ;
        RECT 730.950 19.950 733.050 22.050 ;
        RECT 707.400 3.600 709.200 9.600 ;
        RECT 713.700 3.600 715.500 15.600 ;
        RECT 734.400 9.600 735.600 22.950 ;
        RECT 737.100 22.050 738.900 23.850 ;
        RECT 752.100 22.050 753.900 23.850 ;
        RECT 754.950 22.950 757.050 25.050 ;
        RECT 736.950 19.950 739.050 22.050 ;
        RECT 751.950 19.950 754.050 22.050 ;
        RECT 755.850 9.600 757.050 22.950 ;
        RECT 758.100 22.050 759.900 23.850 ;
        RECT 760.950 22.950 763.050 25.050 ;
        RECT 757.950 19.950 760.050 22.050 ;
        RECT 761.100 21.150 762.900 22.950 ;
        RECT 733.800 3.600 735.600 9.600 ;
        RECT 755.400 3.600 757.200 9.600 ;
        RECT 767.550 7.050 768.450 34.950 ;
        RECT 778.800 31.200 780.600 38.400 ;
        RECT 776.400 30.300 780.600 31.200 ;
        RECT 785.550 32.400 787.350 38.400 ;
        RECT 793.650 35.400 795.450 38.400 ;
        RECT 801.450 35.400 803.250 38.400 ;
        RECT 809.250 36.300 811.050 38.400 ;
        RECT 809.250 35.400 813.000 36.300 ;
        RECT 793.650 34.500 794.700 35.400 ;
        RECT 790.950 33.300 794.700 34.500 ;
        RECT 802.200 34.500 803.250 35.400 ;
        RECT 811.950 34.500 813.000 35.400 ;
        RECT 802.200 33.450 807.150 34.500 ;
        RECT 790.950 32.400 793.050 33.300 ;
        RECT 805.350 32.700 807.150 33.450 ;
        RECT 776.400 25.050 777.600 30.300 ;
        RECT 785.550 25.050 786.750 32.400 ;
        RECT 808.650 31.800 810.450 33.600 ;
        RECT 811.950 32.400 814.050 34.500 ;
        RECT 817.050 32.400 818.850 38.400 ;
        RECT 798.150 30.000 799.950 30.600 ;
        RECT 809.100 30.000 810.150 31.800 ;
        RECT 798.150 28.800 810.150 30.000 ;
        RECT 773.100 22.050 774.900 23.850 ;
        RECT 775.950 22.950 778.050 25.050 ;
        RECT 772.950 19.950 775.050 22.050 ;
        RECT 776.400 9.600 777.600 22.950 ;
        RECT 779.100 22.050 780.900 23.850 ;
        RECT 785.550 23.250 791.850 25.050 ;
        RECT 785.550 22.950 790.050 23.250 ;
        RECT 778.950 19.950 781.050 22.050 ;
        RECT 785.550 15.600 786.750 22.950 ;
        RECT 787.950 17.400 789.750 19.200 ;
        RECT 788.850 16.200 793.050 17.400 ;
        RECT 798.150 16.200 799.050 28.800 ;
        RECT 809.100 27.600 816.000 28.800 ;
        RECT 809.100 27.000 810.900 27.600 ;
        RECT 815.100 26.850 816.000 27.600 ;
        RECT 812.100 25.800 813.900 26.400 ;
        RECT 805.950 24.600 813.900 25.800 ;
        RECT 815.100 25.050 816.900 26.850 ;
        RECT 805.950 22.950 808.050 24.600 ;
        RECT 814.950 22.950 817.050 25.050 ;
        RECT 807.750 17.700 809.550 18.000 ;
        RECT 817.950 17.700 818.850 32.400 ;
        RECT 807.750 17.100 818.850 17.700 ;
        RECT 766.950 4.950 769.050 7.050 ;
        RECT 776.400 3.600 778.200 9.600 ;
        RECT 785.550 3.600 787.350 15.600 ;
        RECT 790.950 15.300 793.050 16.200 ;
        RECT 793.950 15.300 799.050 16.200 ;
        RECT 801.150 16.500 818.850 17.100 ;
        RECT 801.150 16.200 809.550 16.500 ;
        RECT 793.950 14.400 794.850 15.300 ;
        RECT 792.150 12.600 794.850 14.400 ;
        RECT 795.750 14.100 797.550 14.400 ;
        RECT 801.150 14.100 802.050 16.200 ;
        RECT 817.950 15.600 818.850 16.500 ;
        RECT 795.750 13.200 802.050 14.100 ;
        RECT 802.950 14.700 804.750 15.300 ;
        RECT 802.950 13.500 810.450 14.700 ;
        RECT 795.750 12.600 797.550 13.200 ;
        RECT 809.250 12.600 810.450 13.500 ;
        RECT 790.950 9.600 794.850 11.700 ;
        RECT 799.950 11.550 801.750 12.300 ;
        RECT 804.750 11.550 806.550 12.300 ;
        RECT 799.950 10.500 806.550 11.550 ;
        RECT 809.250 10.500 814.050 12.600 ;
        RECT 793.050 3.600 794.850 9.600 ;
        RECT 800.850 3.600 802.650 10.500 ;
        RECT 809.250 9.600 810.450 10.500 ;
        RECT 808.650 3.600 810.450 9.600 ;
        RECT 817.050 3.600 818.850 15.600 ;
        RECT 821.550 32.400 823.350 38.400 ;
        RECT 829.650 35.400 831.450 38.400 ;
        RECT 837.450 35.400 839.250 38.400 ;
        RECT 845.250 36.300 847.050 38.400 ;
        RECT 845.250 35.400 849.000 36.300 ;
        RECT 829.650 34.500 830.700 35.400 ;
        RECT 826.950 33.300 830.700 34.500 ;
        RECT 838.200 34.500 839.250 35.400 ;
        RECT 847.950 34.500 849.000 35.400 ;
        RECT 838.200 33.450 843.150 34.500 ;
        RECT 826.950 32.400 829.050 33.300 ;
        RECT 841.350 32.700 843.150 33.450 ;
        RECT 821.550 25.050 822.750 32.400 ;
        RECT 844.650 31.800 846.450 33.600 ;
        RECT 847.950 32.400 850.050 34.500 ;
        RECT 853.050 32.400 854.850 38.400 ;
        RECT 834.150 30.000 835.950 30.600 ;
        RECT 845.100 30.000 846.150 31.800 ;
        RECT 834.150 28.800 846.150 30.000 ;
        RECT 821.550 23.250 827.850 25.050 ;
        RECT 821.550 22.950 826.050 23.250 ;
        RECT 821.550 15.600 822.750 22.950 ;
        RECT 823.950 17.400 825.750 19.200 ;
        RECT 824.850 16.200 829.050 17.400 ;
        RECT 834.150 16.200 835.050 28.800 ;
        RECT 845.100 27.600 852.000 28.800 ;
        RECT 845.100 27.000 846.900 27.600 ;
        RECT 851.100 26.850 852.000 27.600 ;
        RECT 848.100 25.800 849.900 26.400 ;
        RECT 841.950 24.600 849.900 25.800 ;
        RECT 851.100 25.050 852.900 26.850 ;
        RECT 841.950 22.950 844.050 24.600 ;
        RECT 850.950 22.950 853.050 25.050 ;
        RECT 843.750 17.700 845.550 18.000 ;
        RECT 853.950 17.700 854.850 32.400 ;
        RECT 869.400 35.400 871.200 38.400 ;
        RECT 865.950 22.950 868.050 25.050 ;
        RECT 866.100 21.150 867.900 22.950 ;
        RECT 869.400 22.050 870.600 35.400 ;
        RECT 889.200 32.400 891.000 38.400 ;
        RECT 884.100 25.050 885.900 26.850 ;
        RECT 886.950 25.950 889.050 28.050 ;
        RECT 883.950 22.950 886.050 25.050 ;
        RECT 887.100 24.150 888.900 25.950 ;
        RECT 889.950 25.050 891.000 32.400 ;
        RECT 892.950 25.950 895.050 28.050 ;
        RECT 889.950 22.950 892.050 25.050 ;
        RECT 893.100 24.150 894.900 25.950 ;
        RECT 896.100 25.050 897.900 26.850 ;
        RECT 895.950 22.950 898.050 25.050 ;
        RECT 843.750 17.100 854.850 17.700 ;
        RECT 821.550 3.600 823.350 15.600 ;
        RECT 826.950 15.300 829.050 16.200 ;
        RECT 829.950 15.300 835.050 16.200 ;
        RECT 837.150 16.500 854.850 17.100 ;
        RECT 868.950 16.950 871.050 22.050 ;
        RECT 890.100 17.400 891.000 22.950 ;
        RECT 837.150 16.200 845.550 16.500 ;
        RECT 829.950 14.400 830.850 15.300 ;
        RECT 828.150 12.600 830.850 14.400 ;
        RECT 831.750 14.100 833.550 14.400 ;
        RECT 837.150 14.100 838.050 16.200 ;
        RECT 853.950 15.600 854.850 16.500 ;
        RECT 831.750 13.200 838.050 14.100 ;
        RECT 838.950 14.700 840.750 15.300 ;
        RECT 838.950 13.500 846.450 14.700 ;
        RECT 831.750 12.600 833.550 13.200 ;
        RECT 845.250 12.600 846.450 13.500 ;
        RECT 826.950 9.600 830.850 11.700 ;
        RECT 835.950 11.550 837.750 12.300 ;
        RECT 840.750 11.550 842.550 12.300 ;
        RECT 835.950 10.500 842.550 11.550 ;
        RECT 845.250 10.500 850.050 12.600 ;
        RECT 829.050 3.600 830.850 9.600 ;
        RECT 836.850 3.600 838.650 10.500 ;
        RECT 845.250 9.600 846.450 10.500 ;
        RECT 844.650 3.600 846.450 9.600 ;
        RECT 853.050 3.600 854.850 15.600 ;
        RECT 869.400 9.600 870.600 16.950 ;
        RECT 890.100 16.500 895.200 17.400 ;
        RECT 884.400 14.400 892.200 15.300 ;
        RECT 869.400 3.600 871.200 9.600 ;
        RECT 884.400 3.600 886.200 14.400 ;
        RECT 890.400 4.500 892.200 14.400 ;
        RECT 893.400 5.400 895.200 16.500 ;
        RECT 896.400 4.500 898.200 15.600 ;
        RECT 890.400 3.600 898.200 4.500 ;
      LAYER metal2 ;
        RECT 550.950 900.450 553.050 901.050 ;
        RECT 619.950 900.450 622.050 901.050 ;
        RECT 691.950 900.450 694.050 901.050 ;
        RECT 775.950 900.450 778.050 901.050 ;
        RECT 550.950 899.400 690.450 900.450 ;
        RECT 550.950 898.950 553.050 899.400 ;
        RECT 619.950 898.950 622.050 899.400 ;
        RECT 19.950 897.450 22.050 898.050 ;
        RECT 31.950 897.450 34.050 898.050 ;
        RECT 124.950 897.450 127.050 898.050 ;
        RECT 19.950 896.400 127.050 897.450 ;
        RECT 19.950 895.950 22.050 896.400 ;
        RECT 31.950 895.950 34.050 896.400 ;
        RECT 124.950 895.950 127.050 896.400 ;
        RECT 133.950 897.450 136.050 898.050 ;
        RECT 169.950 897.450 172.050 898.050 ;
        RECT 193.950 897.450 196.050 898.050 ;
        RECT 133.950 896.400 196.050 897.450 ;
        RECT 133.950 895.950 136.050 896.400 ;
        RECT 169.950 895.950 172.050 896.400 ;
        RECT 193.950 895.950 196.050 896.400 ;
        RECT 343.950 897.450 346.050 898.050 ;
        RECT 397.950 897.450 400.050 898.050 ;
        RECT 343.950 896.400 400.050 897.450 ;
        RECT 343.950 895.950 346.050 896.400 ;
        RECT 397.950 895.950 400.050 896.400 ;
        RECT 412.950 897.450 415.050 898.050 ;
        RECT 433.950 897.450 436.050 898.050 ;
        RECT 412.950 896.400 436.050 897.450 ;
        RECT 412.950 895.950 415.050 896.400 ;
        RECT 433.950 895.950 436.050 896.400 ;
        RECT 439.950 897.450 442.050 898.050 ;
        RECT 460.950 897.450 463.050 898.050 ;
        RECT 481.950 897.450 484.050 898.050 ;
        RECT 439.950 896.400 484.050 897.450 ;
        RECT 439.950 895.950 442.050 896.400 ;
        RECT 460.950 895.950 463.050 896.400 ;
        RECT 481.950 895.950 484.050 896.400 ;
        RECT 496.950 897.450 499.050 898.050 ;
        RECT 523.950 897.450 526.050 898.050 ;
        RECT 496.950 896.400 526.050 897.450 ;
        RECT 496.950 895.950 499.050 896.400 ;
        RECT 523.950 895.950 526.050 896.400 ;
        RECT 562.950 897.450 565.050 898.050 ;
        RECT 574.950 897.450 577.050 898.050 ;
        RECT 643.950 897.450 646.050 898.050 ;
        RECT 658.950 897.450 661.050 898.050 ;
        RECT 562.950 896.400 661.050 897.450 ;
        RECT 689.400 897.450 690.450 899.400 ;
        RECT 691.950 899.400 778.050 900.450 ;
        RECT 691.950 898.950 694.050 899.400 ;
        RECT 775.950 898.950 778.050 899.400 ;
        RECT 787.950 900.450 790.050 901.050 ;
        RECT 826.950 900.450 829.050 901.050 ;
        RECT 787.950 899.400 829.050 900.450 ;
        RECT 787.950 898.950 790.050 899.400 ;
        RECT 826.950 898.950 829.050 899.400 ;
        RECT 736.950 897.450 739.050 898.050 ;
        RECT 689.400 896.400 739.050 897.450 ;
        RECT 562.950 895.950 565.050 896.400 ;
        RECT 574.950 895.950 577.050 896.400 ;
        RECT 643.950 895.950 646.050 896.400 ;
        RECT 658.950 895.950 661.050 896.400 ;
        RECT 736.950 895.950 739.050 896.400 ;
        RECT 64.950 894.450 67.050 895.050 ;
        RECT 76.950 894.450 79.050 895.050 ;
        RECT 250.950 894.450 253.050 895.050 ;
        RECT 64.950 893.400 253.050 894.450 ;
        RECT 64.950 892.950 67.050 893.400 ;
        RECT 76.950 892.950 79.050 893.400 ;
        RECT 250.950 892.950 253.050 893.400 ;
        RECT 724.950 894.450 727.050 895.050 ;
        RECT 766.950 894.450 769.050 895.050 ;
        RECT 787.800 894.450 789.900 895.050 ;
        RECT 724.950 893.400 789.900 894.450 ;
        RECT 724.950 892.950 727.050 893.400 ;
        RECT 766.950 892.950 769.050 893.400 ;
        RECT 787.800 892.950 789.900 893.400 ;
        RECT 67.950 891.450 70.050 892.050 ;
        RECT 91.950 891.450 94.050 892.050 ;
        RECT 184.950 891.450 187.050 892.050 ;
        RECT 67.950 890.400 187.050 891.450 ;
        RECT 67.950 889.950 70.050 890.400 ;
        RECT 91.950 889.950 94.050 890.400 ;
        RECT 184.950 889.950 187.050 890.400 ;
        RECT 241.950 891.450 244.050 892.050 ;
        RECT 280.950 891.450 283.050 892.050 ;
        RECT 241.950 890.400 283.050 891.450 ;
        RECT 241.950 889.950 244.050 890.400 ;
        RECT 280.950 889.950 283.050 890.400 ;
        RECT 328.950 891.450 331.050 892.050 ;
        RECT 337.950 891.450 340.050 892.050 ;
        RECT 328.950 890.400 340.050 891.450 ;
        RECT 328.950 889.950 331.050 890.400 ;
        RECT 337.950 889.950 340.050 890.400 ;
        RECT 382.950 891.450 385.050 892.050 ;
        RECT 391.950 891.450 394.050 892.050 ;
        RECT 382.950 890.400 394.050 891.450 ;
        RECT 382.950 889.950 385.050 890.400 ;
        RECT 391.950 889.950 394.050 890.400 ;
        RECT 334.950 888.450 337.050 889.050 ;
        RECT 343.950 888.450 346.050 889.050 ;
        RECT 334.950 887.400 346.050 888.450 ;
        RECT 334.950 886.950 337.050 887.400 ;
        RECT 343.950 886.950 346.050 887.400 ;
        RECT 400.950 888.450 403.050 889.050 ;
        RECT 412.950 888.450 415.050 892.050 ;
        RECT 424.950 891.450 427.050 892.050 ;
        RECT 475.950 891.450 478.050 892.050 ;
        RECT 514.950 891.450 517.050 892.050 ;
        RECT 424.950 890.400 517.050 891.450 ;
        RECT 424.950 889.950 427.050 890.400 ;
        RECT 475.950 889.950 478.050 890.400 ;
        RECT 514.950 889.950 517.050 890.400 ;
        RECT 538.950 891.450 541.050 892.050 ;
        RECT 550.950 891.450 553.050 892.050 ;
        RECT 538.950 890.400 553.050 891.450 ;
        RECT 538.950 889.950 541.050 890.400 ;
        RECT 550.950 889.950 553.050 890.400 ;
        RECT 709.950 891.450 712.050 892.050 ;
        RECT 718.950 891.450 721.050 892.050 ;
        RECT 709.950 890.400 721.050 891.450 ;
        RECT 709.950 889.950 712.050 890.400 ;
        RECT 718.950 889.950 721.050 890.400 ;
        RECT 808.950 891.450 811.050 892.050 ;
        RECT 832.950 891.450 835.050 892.050 ;
        RECT 865.950 891.450 868.050 892.050 ;
        RECT 808.950 890.400 868.050 891.450 ;
        RECT 808.950 889.950 811.050 890.400 ;
        RECT 832.950 889.950 835.050 890.400 ;
        RECT 865.950 889.950 868.050 890.400 ;
        RECT 400.950 887.400 415.050 888.450 ;
        RECT 400.950 886.950 403.050 887.400 ;
        RECT 412.950 886.950 415.050 887.400 ;
        RECT 418.950 886.950 421.050 889.050 ;
        RECT 13.950 883.950 16.050 886.050 ;
        RECT 19.950 883.950 22.050 886.050 ;
        RECT 25.950 885.450 28.050 886.050 ;
        RECT 37.950 885.450 40.050 886.050 ;
        RECT 25.950 884.400 40.050 885.450 ;
        RECT 25.950 883.950 28.050 884.400 ;
        RECT 37.950 883.950 40.050 884.400 ;
        RECT 43.950 883.950 46.050 886.050 ;
        RECT 46.800 883.950 48.900 886.050 ;
        RECT 50.100 885.450 52.200 886.050 ;
        RECT 61.950 885.450 64.050 886.050 ;
        RECT 50.100 884.400 64.050 885.450 ;
        RECT 50.100 883.950 52.200 884.400 ;
        RECT 61.950 883.950 64.050 884.400 ;
        RECT 67.950 883.950 70.050 886.050 ;
        RECT 82.950 883.950 85.050 886.050 ;
        RECT 85.950 883.950 88.050 886.050 ;
        RECT 91.950 883.950 94.050 886.050 ;
        RECT 103.950 885.450 106.050 886.050 ;
        RECT 112.950 885.450 115.050 886.050 ;
        RECT 103.950 884.400 115.050 885.450 ;
        RECT 103.950 883.950 106.050 884.400 ;
        RECT 112.950 883.950 115.050 884.400 ;
        RECT 118.950 883.950 121.050 886.050 ;
        RECT 124.950 885.450 127.050 886.050 ;
        RECT 136.950 885.450 139.050 886.050 ;
        RECT 124.950 884.400 139.050 885.450 ;
        RECT 124.950 883.950 127.050 884.400 ;
        RECT 136.950 883.950 139.050 884.400 ;
        RECT 142.950 883.950 145.050 886.050 ;
        RECT 154.950 883.950 157.050 886.050 ;
        RECT 172.950 883.950 175.050 886.050 ;
        RECT 193.950 883.950 196.050 886.050 ;
        RECT 199.950 883.950 205.050 886.050 ;
        RECT 220.950 885.450 223.050 886.050 ;
        RECT 229.950 885.450 232.050 886.050 ;
        RECT 220.950 884.400 232.050 885.450 ;
        RECT 220.950 883.950 223.050 884.400 ;
        RECT 229.950 883.950 232.050 884.400 ;
        RECT 235.950 883.950 238.050 886.050 ;
        RECT 241.950 883.950 244.050 886.050 ;
        RECT 250.950 885.450 253.050 886.050 ;
        RECT 262.950 885.450 265.050 886.050 ;
        RECT 250.950 884.400 265.050 885.450 ;
        RECT 250.950 883.950 253.050 884.400 ;
        RECT 262.950 883.950 265.050 884.400 ;
        RECT 328.950 883.950 331.050 886.050 ;
        RECT 349.950 883.950 352.050 886.050 ;
        RECT 373.950 885.450 376.050 886.050 ;
        RECT 382.950 885.450 385.050 886.050 ;
        RECT 373.950 884.400 385.050 885.450 ;
        RECT 373.950 883.950 376.050 884.400 ;
        RECT 382.950 883.950 385.050 884.400 ;
        RECT 391.950 883.950 394.050 886.050 ;
        RECT 397.950 885.450 400.050 886.050 ;
        RECT 406.950 885.450 409.050 886.050 ;
        RECT 397.950 884.400 409.050 885.450 ;
        RECT 397.950 883.950 400.050 884.400 ;
        RECT 406.950 883.950 409.050 884.400 ;
        RECT 412.950 883.950 415.050 885.750 ;
        RECT 418.950 883.950 421.050 885.750 ;
        RECT 433.950 883.950 436.050 886.050 ;
        RECT 478.950 883.950 481.050 886.050 ;
        RECT 487.950 885.450 490.050 886.050 ;
        RECT 499.950 885.450 502.050 886.050 ;
        RECT 487.950 884.400 502.050 885.450 ;
        RECT 487.950 883.950 490.050 884.400 ;
        RECT 499.950 883.950 502.050 884.400 ;
        RECT 505.950 883.950 508.050 886.050 ;
        RECT 511.950 885.450 514.050 886.050 ;
        RECT 517.950 885.450 520.050 886.050 ;
        RECT 511.950 884.400 520.050 885.450 ;
        RECT 511.950 883.950 514.050 884.400 ;
        RECT 517.950 883.950 520.050 884.400 ;
        RECT 523.950 883.950 526.050 889.050 ;
        RECT 532.950 888.450 535.050 889.050 ;
        RECT 541.950 888.450 544.050 889.050 ;
        RECT 532.950 887.400 544.050 888.450 ;
        RECT 532.950 886.950 535.050 887.400 ;
        RECT 541.950 886.950 544.050 887.400 ;
        RECT 637.950 886.950 640.050 889.050 ;
        RECT 643.950 886.950 646.050 889.050 ;
        RECT 766.950 886.950 772.050 889.050 ;
        RECT 787.950 888.450 790.050 889.050 ;
        RECT 799.950 888.450 802.050 889.050 ;
        RECT 787.950 887.400 802.050 888.450 ;
        RECT 787.950 886.950 790.050 887.400 ;
        RECT 799.950 886.950 802.050 887.400 ;
        RECT 529.950 883.950 532.050 886.050 ;
        RECT 535.950 885.450 538.050 886.050 ;
        RECT 547.950 885.450 550.050 886.050 ;
        RECT 535.950 884.400 550.050 885.450 ;
        RECT 535.950 883.950 538.050 884.400 ;
        RECT 547.950 883.950 550.050 884.400 ;
        RECT 553.950 885.450 556.050 886.050 ;
        RECT 568.950 885.450 571.050 886.050 ;
        RECT 553.950 884.400 571.050 885.450 ;
        RECT 553.950 883.950 556.050 884.400 ;
        RECT 568.950 883.950 571.050 884.400 ;
        RECT 574.950 883.950 577.050 886.050 ;
        RECT 580.950 885.450 583.050 886.050 ;
        RECT 595.950 885.450 598.050 886.050 ;
        RECT 580.950 884.400 598.050 885.450 ;
        RECT 580.950 883.950 583.050 884.400 ;
        RECT 595.950 883.950 598.050 884.400 ;
        RECT 637.950 883.950 640.050 885.750 ;
        RECT 643.950 883.950 646.050 885.750 ;
        RECT 685.950 883.950 688.050 886.050 ;
        RECT 724.950 883.950 727.050 886.050 ;
        RECT 745.950 883.950 748.050 885.750 ;
        RECT 751.950 883.950 754.050 885.750 ;
        RECT 775.950 883.950 778.050 886.050 ;
        RECT 799.950 883.950 802.050 885.750 ;
        RECT 805.950 883.950 808.050 885.750 ;
        RECT 823.950 885.450 826.050 886.050 ;
        RECT 835.950 885.450 838.050 886.050 ;
        RECT 823.950 884.400 838.050 885.450 ;
        RECT 823.950 883.950 826.050 884.400 ;
        RECT 835.950 883.950 838.050 884.400 ;
        RECT 841.950 883.950 844.050 886.050 ;
        RECT 847.950 885.450 850.050 886.050 ;
        RECT 859.950 885.450 862.050 886.050 ;
        RECT 847.950 884.400 862.050 885.450 ;
        RECT 847.950 883.950 850.050 884.400 ;
        RECT 859.950 883.950 862.050 884.400 ;
        RECT 865.950 883.950 868.050 886.050 ;
        RECT 886.950 883.950 889.050 886.050 ;
        RECT 13.950 880.950 16.050 882.750 ;
        RECT 19.950 880.950 22.050 882.750 ;
        RECT 37.950 880.950 40.050 882.750 ;
        RECT 43.950 880.950 46.050 882.750 ;
        RECT 61.950 880.950 64.050 882.750 ;
        RECT 67.950 880.950 70.050 882.750 ;
        RECT 85.950 880.950 88.050 882.750 ;
        RECT 91.950 880.950 94.050 882.750 ;
        RECT 100.950 882.450 103.050 883.050 ;
        RECT 106.950 882.450 109.050 883.050 ;
        RECT 100.950 881.400 109.050 882.450 ;
        RECT 100.950 880.950 103.050 881.400 ;
        RECT 106.950 880.950 109.050 881.400 ;
        RECT 112.950 880.950 115.050 882.750 ;
        RECT 118.950 880.950 121.050 882.750 ;
        RECT 127.950 880.950 133.050 883.050 ;
        RECT 136.950 880.950 139.050 882.750 ;
        RECT 142.950 880.950 145.050 882.750 ;
        RECT 154.950 880.950 157.050 882.750 ;
        RECT 172.950 880.950 175.050 882.750 ;
        RECT 193.950 880.950 196.050 882.750 ;
        RECT 199.950 880.950 202.050 882.750 ;
        RECT 220.950 880.950 223.050 882.750 ;
        RECT 235.950 880.950 238.050 882.750 ;
        RECT 241.950 880.950 244.050 882.750 ;
        RECT 262.950 880.950 265.050 882.750 ;
        RECT 283.950 881.250 286.050 883.050 ;
        RECT 289.950 880.950 292.050 882.750 ;
        RECT 301.950 880.950 304.050 882.750 ;
        RECT 307.950 881.250 310.050 883.050 ;
        RECT 328.950 880.950 331.050 882.750 ;
        RECT 343.950 881.250 346.050 883.050 ;
        RECT 353.250 882.750 355.050 883.050 ;
        RECT 349.950 881.250 352.050 882.750 ;
        RECT 352.950 881.250 355.050 882.750 ;
        RECT 349.950 880.950 351.750 881.250 ;
        RECT 373.950 880.950 376.050 882.750 ;
        RECT 379.950 882.450 382.050 883.050 ;
        RECT 385.950 882.450 388.050 883.050 ;
        RECT 379.950 881.400 388.050 882.450 ;
        RECT 379.950 880.950 382.050 881.400 ;
        RECT 385.950 880.950 388.050 881.400 ;
        RECT 391.950 880.950 394.050 882.750 ;
        RECT 415.950 881.250 418.050 883.050 ;
        RECT 433.950 880.950 436.050 882.750 ;
        RECT 451.950 880.950 454.050 882.750 ;
        RECT 457.950 881.250 460.050 883.050 ;
        RECT 475.950 882.750 477.750 883.050 ;
        RECT 475.950 881.250 478.050 882.750 ;
        RECT 478.950 881.250 481.050 882.750 ;
        RECT 484.950 881.250 487.050 883.050 ;
        RECT 479.250 880.950 481.050 881.250 ;
        RECT 499.950 880.950 502.050 882.750 ;
        RECT 505.950 880.950 508.050 882.750 ;
        RECT 523.950 880.950 526.050 882.750 ;
        RECT 529.950 880.950 532.050 882.750 ;
        RECT 547.950 880.950 550.050 882.750 ;
        RECT 568.950 880.950 571.050 882.750 ;
        RECT 574.950 880.950 577.050 882.750 ;
        RECT 595.950 880.950 598.050 882.750 ;
        RECT 610.950 880.950 613.050 882.750 ;
        RECT 616.950 881.250 619.050 883.050 ;
        RECT 634.950 881.250 637.050 883.050 ;
        RECT 640.950 881.250 643.050 883.050 ;
        RECT 646.950 881.250 649.050 883.050 ;
        RECT 661.950 881.250 664.050 883.050 ;
        RECT 667.950 880.950 670.050 882.750 ;
        RECT 685.950 880.950 688.050 882.750 ;
        RECT 697.950 880.950 700.050 882.750 ;
        RECT 703.950 881.250 706.050 883.050 ;
        RECT 721.950 882.750 723.750 883.050 ;
        RECT 721.950 881.250 724.050 882.750 ;
        RECT 724.950 881.250 727.050 882.750 ;
        RECT 730.950 881.250 733.050 883.050 ;
        RECT 742.950 881.250 745.050 883.050 ;
        RECT 748.950 881.250 751.050 883.050 ;
        RECT 754.950 881.250 757.050 883.050 ;
        RECT 769.950 881.250 772.050 883.050 ;
        RECT 779.250 882.750 781.050 883.050 ;
        RECT 775.950 881.250 778.050 882.750 ;
        RECT 778.950 881.250 781.050 882.750 ;
        RECT 796.950 881.250 799.050 883.050 ;
        RECT 802.950 881.250 805.050 883.050 ;
        RECT 808.950 881.250 811.050 883.050 ;
        RECT 725.250 880.950 727.050 881.250 ;
        RECT 775.950 880.950 777.750 881.250 ;
        RECT 823.950 880.950 826.050 882.750 ;
        RECT 841.950 880.950 844.050 882.750 ;
        RECT 847.950 880.950 850.050 882.750 ;
        RECT 865.950 880.950 868.050 882.750 ;
        RECT 886.950 880.950 889.050 882.750 ;
        RECT 892.950 881.250 895.050 883.050 ;
        RECT 16.950 878.250 19.050 880.050 ;
        RECT 22.950 878.250 25.050 880.050 ;
        RECT 34.950 878.250 37.050 880.050 ;
        RECT 40.950 878.250 43.050 880.050 ;
        RECT 64.950 878.250 67.050 880.050 ;
        RECT 70.950 878.250 73.050 880.050 ;
        RECT 88.950 878.250 91.050 880.050 ;
        RECT 94.950 878.250 97.050 880.050 ;
        RECT 109.950 878.250 112.050 880.050 ;
        RECT 115.950 878.250 118.050 880.050 ;
        RECT 133.950 878.250 136.050 880.050 ;
        RECT 139.950 878.250 142.050 880.050 ;
        RECT 157.950 878.250 160.050 880.050 ;
        RECT 175.950 878.250 178.050 880.050 ;
        RECT 190.950 878.250 193.050 880.050 ;
        RECT 196.950 878.250 199.050 880.050 ;
        RECT 217.950 878.250 220.050 880.050 ;
        RECT 223.950 878.250 226.050 880.050 ;
        RECT 238.950 878.250 241.050 880.050 ;
        RECT 244.950 878.250 247.050 880.050 ;
        RECT 259.950 878.250 262.050 880.050 ;
        RECT 265.950 878.250 268.050 880.050 ;
        RECT 274.950 879.450 277.050 880.050 ;
        RECT 283.950 879.450 286.050 880.050 ;
        RECT 274.950 878.400 286.050 879.450 ;
        RECT 274.950 877.950 277.050 878.400 ;
        RECT 283.950 877.950 286.050 878.400 ;
        RECT 307.950 879.450 310.050 880.050 ;
        RECT 316.950 879.450 319.050 880.050 ;
        RECT 307.950 878.400 319.050 879.450 ;
        RECT 307.950 877.950 310.050 878.400 ;
        RECT 316.950 877.950 319.050 878.400 ;
        RECT 325.950 878.250 328.050 880.050 ;
        RECT 331.950 878.250 334.050 880.050 ;
        RECT 343.950 877.950 346.050 880.050 ;
        RECT 352.950 879.450 355.050 880.050 ;
        RECT 364.950 879.450 367.050 880.050 ;
        RECT 352.950 878.400 367.050 879.450 ;
        RECT 352.950 877.950 355.050 878.400 ;
        RECT 364.950 877.950 367.050 878.400 ;
        RECT 370.950 878.250 373.050 880.050 ;
        RECT 376.950 878.250 379.050 880.050 ;
        RECT 388.950 878.250 391.050 880.050 ;
        RECT 394.950 878.250 397.050 880.050 ;
        RECT 400.950 879.450 403.050 880.050 ;
        RECT 415.950 879.450 418.050 880.050 ;
        RECT 400.950 878.400 418.050 879.450 ;
        RECT 400.950 877.950 403.050 878.400 ;
        RECT 415.950 877.950 418.050 878.400 ;
        RECT 430.950 878.250 433.050 880.050 ;
        RECT 436.950 878.250 439.050 880.050 ;
        RECT 457.950 877.950 463.050 880.050 ;
        RECT 475.950 877.950 478.050 880.050 ;
        RECT 484.950 877.950 487.050 880.050 ;
        RECT 502.950 878.250 505.050 880.050 ;
        RECT 508.950 878.250 511.050 880.050 ;
        RECT 526.950 878.250 529.050 880.050 ;
        RECT 532.950 878.250 535.050 880.050 ;
        RECT 544.950 878.250 547.050 880.050 ;
        RECT 550.950 878.250 553.050 880.050 ;
        RECT 571.950 878.250 574.050 880.050 ;
        RECT 577.950 878.250 580.050 880.050 ;
        RECT 592.950 878.250 595.050 880.050 ;
        RECT 598.950 878.250 601.050 880.050 ;
        RECT 613.950 879.450 619.050 880.050 ;
        RECT 628.950 879.450 631.050 880.050 ;
        RECT 613.950 878.400 631.050 879.450 ;
        RECT 613.950 877.950 619.050 878.400 ;
        RECT 628.950 877.950 631.050 878.400 ;
        RECT 634.950 877.950 637.050 880.050 ;
        RECT 16.950 874.950 19.050 877.050 ;
        RECT 22.950 874.950 25.050 877.050 ;
        RECT 34.950 874.950 37.050 877.050 ;
        RECT 40.950 874.950 43.050 877.050 ;
        RECT 64.950 874.950 67.050 877.050 ;
        RECT 70.950 874.950 73.050 877.050 ;
        RECT 76.950 876.450 79.050 877.050 ;
        RECT 82.950 876.450 85.050 877.050 ;
        RECT 76.950 875.400 85.050 876.450 ;
        RECT 76.950 874.950 79.050 875.400 ;
        RECT 82.950 874.950 85.050 875.400 ;
        RECT 88.950 874.950 91.050 877.050 ;
        RECT 94.950 874.950 97.050 877.050 ;
        RECT 100.950 876.450 103.050 877.050 ;
        RECT 109.950 876.450 112.050 877.050 ;
        RECT 100.950 875.400 112.050 876.450 ;
        RECT 100.950 874.950 103.050 875.400 ;
        RECT 109.950 874.950 112.050 875.400 ;
        RECT 115.950 874.950 118.050 877.050 ;
        RECT 121.950 876.450 124.050 877.050 ;
        RECT 133.950 876.450 136.050 877.050 ;
        RECT 121.950 875.400 136.050 876.450 ;
        RECT 121.950 874.950 124.050 875.400 ;
        RECT 133.950 874.950 136.050 875.400 ;
        RECT 139.950 876.450 142.050 877.050 ;
        RECT 144.000 876.450 148.050 877.050 ;
        RECT 139.950 875.400 148.050 876.450 ;
        RECT 139.950 874.950 142.050 875.400 ;
        RECT 144.000 874.950 148.050 875.400 ;
        RECT 157.950 876.450 160.050 877.050 ;
        RECT 169.950 876.450 172.050 877.050 ;
        RECT 157.950 875.400 172.050 876.450 ;
        RECT 157.950 874.950 160.050 875.400 ;
        RECT 169.950 874.950 172.050 875.400 ;
        RECT 175.950 876.450 178.050 877.050 ;
        RECT 184.950 876.450 187.050 877.050 ;
        RECT 175.950 875.400 187.050 876.450 ;
        RECT 175.950 874.950 178.050 875.400 ;
        RECT 184.950 874.950 187.050 875.400 ;
        RECT 190.950 874.950 193.050 877.050 ;
        RECT 196.950 874.950 199.050 877.050 ;
        RECT 223.950 874.950 226.050 877.050 ;
        RECT 238.950 874.950 241.050 877.050 ;
        RECT 244.950 874.950 247.050 877.050 ;
        RECT 259.950 874.950 262.050 877.050 ;
        RECT 265.950 874.950 268.050 877.050 ;
        RECT 325.950 874.950 328.050 877.050 ;
        RECT 331.950 874.950 334.050 877.050 ;
        RECT 370.950 874.950 373.050 877.050 ;
        RECT 376.950 874.950 379.050 877.050 ;
        RECT 127.950 873.450 130.050 874.050 ;
        RECT 119.400 872.400 130.050 873.450 ;
        RECT 76.950 870.450 79.050 871.050 ;
        RECT 88.950 870.450 91.050 871.050 ;
        RECT 76.950 869.400 91.050 870.450 ;
        RECT 76.950 868.950 79.050 869.400 ;
        RECT 88.950 868.950 91.050 869.400 ;
        RECT 94.950 870.450 97.050 871.050 ;
        RECT 100.950 870.450 103.050 871.050 ;
        RECT 94.950 869.400 103.050 870.450 ;
        RECT 94.950 868.950 97.050 869.400 ;
        RECT 100.950 868.950 103.050 869.400 ;
        RECT 109.950 870.450 112.050 871.050 ;
        RECT 119.400 870.450 120.450 872.400 ;
        RECT 127.950 871.950 130.050 872.400 ;
        RECT 382.950 871.950 385.050 877.050 ;
        RECT 388.950 874.950 391.050 877.050 ;
        RECT 394.950 874.950 397.050 877.050 ;
        RECT 430.950 874.950 433.050 877.050 ;
        RECT 436.950 874.950 439.050 877.050 ;
        RECT 502.950 874.950 505.050 877.050 ;
        RECT 508.950 874.950 511.050 877.050 ;
        RECT 406.950 873.450 409.050 874.050 ;
        RECT 418.950 873.450 421.050 874.050 ;
        RECT 406.950 872.400 421.050 873.450 ;
        RECT 406.950 871.950 409.050 872.400 ;
        RECT 418.950 871.950 421.050 872.400 ;
        RECT 442.950 873.450 445.050 874.050 ;
        RECT 454.950 873.450 457.050 874.050 ;
        RECT 442.950 872.400 457.050 873.450 ;
        RECT 442.950 871.950 445.050 872.400 ;
        RECT 454.950 871.950 457.050 872.400 ;
        RECT 463.950 873.450 466.050 874.050 ;
        RECT 484.950 873.450 487.050 874.050 ;
        RECT 490.950 873.450 493.050 874.050 ;
        RECT 463.950 872.400 493.050 873.450 ;
        RECT 463.950 871.950 466.050 872.400 ;
        RECT 484.950 871.950 487.050 872.400 ;
        RECT 490.950 871.950 493.050 872.400 ;
        RECT 514.950 871.950 517.050 877.050 ;
        RECT 526.950 874.950 529.050 877.050 ;
        RECT 532.950 874.950 535.050 877.050 ;
        RECT 538.950 876.450 543.000 877.050 ;
        RECT 544.950 876.450 547.050 877.050 ;
        RECT 538.950 875.400 547.050 876.450 ;
        RECT 538.950 874.950 543.000 875.400 ;
        RECT 544.950 874.950 547.050 875.400 ;
        RECT 571.950 874.950 574.050 877.050 ;
        RECT 577.950 874.950 580.050 877.050 ;
        RECT 580.950 874.950 583.050 877.050 ;
        RECT 592.950 874.950 595.050 877.050 ;
        RECT 598.950 874.950 601.050 877.050 ;
        RECT 640.950 874.950 643.050 880.050 ;
        RECT 646.950 877.950 649.050 880.050 ;
        RECT 658.950 877.950 664.050 880.050 ;
        RECT 682.950 878.250 685.050 880.050 ;
        RECT 703.950 879.450 706.050 880.050 ;
        RECT 715.800 879.450 717.900 880.050 ;
        RECT 703.950 878.400 717.900 879.450 ;
        RECT 703.950 877.950 706.050 878.400 ;
        RECT 715.800 877.950 717.900 878.400 ;
        RECT 719.100 877.950 724.050 880.050 ;
        RECT 730.950 877.950 733.050 880.050 ;
        RECT 742.950 877.950 745.050 880.050 ;
        RECT 748.950 877.950 751.050 880.050 ;
        RECT 754.950 877.950 757.050 880.050 ;
        RECT 769.950 877.950 772.050 880.050 ;
        RECT 778.950 879.450 781.050 880.050 ;
        RECT 783.000 879.450 787.050 880.050 ;
        RECT 778.950 878.400 787.050 879.450 ;
        RECT 778.950 877.950 781.050 878.400 ;
        RECT 783.000 877.950 787.050 878.400 ;
        RECT 796.950 877.950 799.050 880.050 ;
        RECT 802.950 877.950 805.050 880.050 ;
        RECT 808.950 877.950 811.050 880.050 ;
        RECT 820.950 878.250 823.050 880.050 ;
        RECT 826.950 878.250 829.050 880.050 ;
        RECT 844.950 878.250 847.050 880.050 ;
        RECT 850.950 878.250 853.050 880.050 ;
        RECT 868.950 878.250 871.050 880.050 ;
        RECT 883.950 878.250 886.050 880.050 ;
        RECT 892.950 879.450 895.050 880.050 ;
        RECT 910.950 879.450 913.050 880.050 ;
        RECT 892.950 878.400 913.050 879.450 ;
        RECT 892.950 877.950 895.050 878.400 ;
        RECT 910.950 877.950 913.050 878.400 ;
        RECT 682.950 874.950 688.050 877.050 ;
        RECT 634.950 873.450 637.050 874.050 ;
        RECT 670.950 873.450 673.050 874.050 ;
        RECT 634.950 872.400 673.050 873.450 ;
        RECT 634.950 871.950 637.050 872.400 ;
        RECT 670.950 871.950 673.050 872.400 ;
        RECT 709.950 873.450 712.050 874.050 ;
        RECT 749.400 873.450 750.450 877.950 ;
        RECT 820.950 874.950 823.050 877.050 ;
        RECT 826.950 874.950 829.050 877.050 ;
        RECT 844.950 874.950 847.050 877.050 ;
        RECT 850.950 876.450 853.050 877.050 ;
        RECT 868.950 876.450 871.050 877.050 ;
        RECT 850.950 875.400 871.050 876.450 ;
        RECT 850.950 874.950 853.050 875.400 ;
        RECT 868.950 874.950 871.050 875.400 ;
        RECT 883.950 874.950 886.050 877.050 ;
        RECT 808.950 873.450 813.900 874.050 ;
        RECT 709.950 872.400 750.450 873.450 ;
        RECT 767.400 872.400 813.900 873.450 ;
        RECT 709.950 871.950 712.050 872.400 ;
        RECT 767.400 871.050 768.450 872.400 ;
        RECT 808.950 871.950 813.900 872.400 ;
        RECT 109.950 869.400 120.450 870.450 ;
        RECT 127.950 870.450 130.050 871.050 ;
        RECT 133.950 870.450 136.050 871.050 ;
        RECT 127.950 869.400 136.050 870.450 ;
        RECT 109.950 868.950 112.050 869.400 ;
        RECT 127.950 868.950 130.050 869.400 ;
        RECT 133.950 868.950 136.050 869.400 ;
        RECT 139.950 870.450 142.050 871.050 ;
        RECT 154.950 870.450 157.050 871.050 ;
        RECT 229.950 870.450 232.050 871.050 ;
        RECT 238.950 870.450 241.050 871.050 ;
        RECT 139.950 869.400 241.050 870.450 ;
        RECT 139.950 868.950 142.050 869.400 ;
        RECT 154.950 868.950 157.050 869.400 ;
        RECT 229.950 868.950 232.050 869.400 ;
        RECT 238.950 868.950 241.050 869.400 ;
        RECT 619.950 870.450 622.050 871.050 ;
        RECT 628.950 870.450 631.050 871.050 ;
        RECT 619.950 869.400 631.050 870.450 ;
        RECT 619.950 868.950 622.050 869.400 ;
        RECT 628.950 868.950 631.050 869.400 ;
        RECT 643.950 870.450 646.050 871.050 ;
        RECT 736.950 870.450 739.050 871.050 ;
        RECT 766.950 870.450 769.050 871.050 ;
        RECT 643.950 869.400 769.050 870.450 ;
        RECT 643.950 868.950 646.050 869.400 ;
        RECT 736.950 868.950 739.050 869.400 ;
        RECT 766.950 868.950 769.050 869.400 ;
        RECT 826.950 870.450 829.050 871.050 ;
        RECT 844.950 870.450 847.050 871.050 ;
        RECT 826.950 869.400 847.050 870.450 ;
        RECT 826.950 868.950 829.050 869.400 ;
        RECT 844.950 868.950 847.050 869.400 ;
        RECT 883.950 870.450 886.050 871.050 ;
        RECT 895.950 870.450 898.050 871.050 ;
        RECT 883.950 869.400 898.050 870.450 ;
        RECT 883.950 868.950 886.050 869.400 ;
        RECT 895.950 868.950 898.050 869.400 ;
        RECT 115.950 867.450 118.050 868.050 ;
        RECT 145.950 867.450 148.050 868.050 ;
        RECT 196.950 867.450 199.050 868.050 ;
        RECT 115.950 866.400 199.050 867.450 ;
        RECT 115.950 865.950 118.050 866.400 ;
        RECT 145.950 865.950 148.050 866.400 ;
        RECT 196.950 865.950 199.050 866.400 ;
        RECT 211.950 867.450 214.050 868.050 ;
        RECT 266.100 867.450 268.200 868.050 ;
        RECT 316.950 867.450 319.050 868.050 ;
        RECT 325.950 867.450 328.050 868.050 ;
        RECT 349.950 867.450 352.050 868.050 ;
        RECT 418.800 867.450 420.900 868.050 ;
        RECT 211.950 866.400 264.450 867.450 ;
        RECT 211.950 865.950 214.050 866.400 ;
        RECT 263.400 865.050 264.450 866.400 ;
        RECT 266.100 866.400 273.450 867.450 ;
        RECT 266.100 865.950 268.200 866.400 ;
        RECT 13.950 864.450 16.050 865.050 ;
        RECT 34.950 864.450 37.050 865.050 ;
        RECT 13.950 863.400 37.050 864.450 ;
        RECT 13.950 862.950 16.050 863.400 ;
        RECT 34.950 862.950 37.050 863.400 ;
        RECT 43.950 864.450 46.050 865.050 ;
        RECT 49.950 864.450 52.050 865.050 ;
        RECT 43.950 863.400 52.050 864.450 ;
        RECT 43.950 862.950 46.050 863.400 ;
        RECT 49.950 862.950 52.050 863.400 ;
        RECT 76.950 862.950 81.900 865.050 ;
        RECT 83.100 864.450 85.200 865.050 ;
        RECT 103.950 864.450 106.050 865.050 ;
        RECT 83.100 863.400 106.050 864.450 ;
        RECT 83.100 862.950 85.200 863.400 ;
        RECT 103.950 862.950 106.050 863.400 ;
        RECT 118.950 864.450 121.050 865.050 ;
        RECT 142.950 864.450 145.050 865.050 ;
        RECT 172.950 864.450 175.050 865.050 ;
        RECT 235.950 864.450 238.050 865.050 ;
        RECT 262.950 864.450 265.050 865.050 ;
        RECT 268.950 864.450 271.050 865.050 ;
        RECT 118.950 863.400 261.450 864.450 ;
        RECT 118.950 862.950 121.050 863.400 ;
        RECT 142.950 862.950 145.050 863.400 ;
        RECT 172.950 862.950 175.050 863.400 ;
        RECT 235.950 862.950 238.050 863.400 ;
        RECT 16.950 861.450 19.050 862.050 ;
        RECT 40.950 861.450 43.050 862.050 ;
        RECT 103.950 861.450 106.050 862.050 ;
        RECT 16.950 860.400 106.050 861.450 ;
        RECT 260.400 861.450 261.450 863.400 ;
        RECT 262.950 863.400 271.050 864.450 ;
        RECT 272.400 864.450 273.450 866.400 ;
        RECT 316.950 866.400 420.900 867.450 ;
        RECT 316.950 865.950 319.050 866.400 ;
        RECT 325.950 865.950 328.050 866.400 ;
        RECT 349.950 865.950 352.050 866.400 ;
        RECT 418.800 865.950 420.900 866.400 ;
        RECT 422.100 867.450 424.200 868.050 ;
        RECT 448.950 867.450 451.050 868.050 ;
        RECT 422.100 866.400 451.050 867.450 ;
        RECT 422.100 865.950 424.200 866.400 ;
        RECT 448.950 865.950 451.050 866.400 ;
        RECT 454.950 867.450 457.050 868.050 ;
        RECT 508.950 867.450 511.050 868.050 ;
        RECT 526.950 867.450 529.050 868.050 ;
        RECT 610.950 867.450 613.050 867.900 ;
        RECT 454.950 866.400 507.450 867.450 ;
        RECT 454.950 865.950 457.050 866.400 ;
        RECT 364.950 864.450 367.050 865.050 ;
        RECT 272.400 863.400 367.050 864.450 ;
        RECT 262.950 862.950 265.050 863.400 ;
        RECT 268.950 862.950 271.050 863.400 ;
        RECT 364.950 862.950 367.050 863.400 ;
        RECT 376.950 864.450 379.050 865.050 ;
        RECT 400.950 864.450 403.050 865.050 ;
        RECT 376.950 863.400 403.050 864.450 ;
        RECT 376.950 862.950 379.050 863.400 ;
        RECT 400.950 862.950 403.050 863.400 ;
        RECT 406.950 864.450 409.050 865.050 ;
        RECT 436.950 864.450 439.050 865.050 ;
        RECT 496.950 864.450 499.050 865.050 ;
        RECT 406.950 863.400 429.450 864.450 ;
        RECT 406.950 862.950 409.050 863.400 ;
        RECT 319.950 861.450 322.050 862.050 ;
        RECT 260.400 860.400 322.050 861.450 ;
        RECT 16.950 859.950 19.050 860.400 ;
        RECT 40.950 859.950 43.050 860.400 ;
        RECT 103.950 859.950 106.050 860.400 ;
        RECT 319.950 859.950 322.050 860.400 ;
        RECT 394.950 861.450 397.050 862.050 ;
        RECT 412.950 861.450 415.050 862.050 ;
        RECT 424.950 861.450 427.050 862.050 ;
        RECT 394.950 860.400 427.050 861.450 ;
        RECT 428.400 861.450 429.450 863.400 ;
        RECT 436.950 863.400 499.050 864.450 ;
        RECT 506.400 864.450 507.450 866.400 ;
        RECT 508.950 866.400 613.050 867.450 ;
        RECT 508.950 865.950 511.050 866.400 ;
        RECT 526.950 865.950 529.050 866.400 ;
        RECT 610.950 865.800 613.050 866.400 ;
        RECT 625.950 867.450 628.050 868.050 ;
        RECT 634.950 867.450 637.050 868.200 ;
        RECT 625.950 866.400 637.050 867.450 ;
        RECT 625.950 865.950 628.050 866.400 ;
        RECT 634.950 866.100 637.050 866.400 ;
        RECT 640.950 867.450 643.050 868.050 ;
        RECT 679.950 867.450 682.050 868.050 ;
        RECT 688.950 867.450 691.050 868.050 ;
        RECT 640.950 866.400 691.050 867.450 ;
        RECT 640.950 865.950 643.050 866.400 ;
        RECT 679.950 865.950 682.050 866.400 ;
        RECT 688.950 865.950 691.050 866.400 ;
        RECT 697.950 867.450 700.050 868.050 ;
        RECT 709.800 867.450 711.900 868.050 ;
        RECT 697.950 866.400 711.900 867.450 ;
        RECT 697.950 865.950 700.050 866.400 ;
        RECT 709.800 865.950 711.900 866.400 ;
        RECT 811.950 867.450 814.050 868.050 ;
        RECT 820.950 867.450 823.050 868.050 ;
        RECT 811.950 866.400 823.050 867.450 ;
        RECT 811.950 865.950 814.050 866.400 ;
        RECT 820.950 865.950 823.050 866.400 ;
        RECT 535.800 864.450 537.900 865.050 ;
        RECT 506.400 863.400 537.900 864.450 ;
        RECT 436.950 862.950 439.050 863.400 ;
        RECT 496.950 862.950 499.050 863.400 ;
        RECT 535.800 862.950 537.900 863.400 ;
        RECT 539.100 864.450 541.200 865.050 ;
        RECT 580.950 864.450 583.050 865.050 ;
        RECT 592.950 864.450 595.050 865.050 ;
        RECT 613.950 864.450 616.050 865.050 ;
        RECT 634.950 864.450 637.050 864.900 ;
        RECT 703.950 864.450 706.050 865.050 ;
        RECT 754.950 864.450 757.050 865.050 ;
        RECT 539.100 863.400 591.450 864.450 ;
        RECT 539.100 862.950 541.200 863.400 ;
        RECT 580.950 862.950 583.050 863.400 ;
        RECT 442.950 861.450 445.050 862.050 ;
        RECT 428.400 860.400 445.050 861.450 ;
        RECT 394.950 859.950 397.050 860.400 ;
        RECT 412.950 859.950 415.050 860.400 ;
        RECT 424.950 859.950 427.050 860.400 ;
        RECT 442.950 859.950 445.050 860.400 ;
        RECT 448.950 861.450 451.050 862.050 ;
        RECT 490.950 861.450 493.050 862.200 ;
        RECT 539.400 861.450 540.450 862.950 ;
        RECT 448.950 860.400 468.450 861.450 ;
        RECT 448.950 859.950 451.050 860.400 ;
        RECT 223.950 858.450 226.050 859.050 ;
        RECT 259.950 858.450 262.050 859.050 ;
        RECT 223.950 857.400 262.050 858.450 ;
        RECT 223.950 856.950 226.050 857.400 ;
        RECT 259.950 856.950 262.050 857.400 ;
        RECT 298.950 858.450 301.050 859.050 ;
        RECT 310.950 858.450 313.050 859.050 ;
        RECT 421.950 858.450 424.050 859.050 ;
        RECT 298.950 857.400 424.050 858.450 ;
        RECT 298.950 856.950 301.050 857.400 ;
        RECT 310.950 856.950 313.050 857.400 ;
        RECT 421.950 856.950 424.050 857.400 ;
        RECT 430.950 858.450 433.050 859.050 ;
        RECT 463.950 858.450 466.050 859.050 ;
        RECT 430.950 857.400 466.050 858.450 ;
        RECT 467.400 858.450 468.450 860.400 ;
        RECT 490.950 860.400 540.450 861.450 ;
        RECT 544.950 861.450 547.050 862.050 ;
        RECT 590.400 861.450 591.450 863.400 ;
        RECT 592.950 863.400 637.050 864.450 ;
        RECT 592.950 862.950 595.050 863.400 ;
        RECT 613.950 862.950 616.050 863.400 ;
        RECT 634.950 862.800 637.050 863.400 ;
        RECT 674.400 863.400 757.050 864.450 ;
        RECT 674.400 861.450 675.450 863.400 ;
        RECT 703.950 862.950 706.050 863.400 ;
        RECT 754.950 862.950 757.050 863.400 ;
        RECT 544.950 860.400 573.450 861.450 ;
        RECT 590.400 860.400 675.450 861.450 ;
        RECT 691.950 861.450 694.050 862.050 ;
        RECT 724.950 861.450 727.050 862.050 ;
        RECT 691.950 860.400 727.050 861.450 ;
        RECT 490.950 860.100 493.050 860.400 ;
        RECT 544.950 859.950 547.050 860.400 ;
        RECT 490.950 858.450 493.050 858.900 ;
        RECT 467.400 857.400 493.050 858.450 ;
        RECT 430.950 856.950 433.050 857.400 ;
        RECT 463.950 856.950 466.050 857.400 ;
        RECT 490.950 856.800 493.050 857.400 ;
        RECT 496.950 858.450 499.050 859.050 ;
        RECT 568.950 858.450 571.050 859.050 ;
        RECT 496.950 857.400 571.050 858.450 ;
        RECT 572.400 858.450 573.450 860.400 ;
        RECT 691.950 859.950 694.050 860.400 ;
        RECT 724.950 859.950 727.050 860.400 ;
        RECT 580.950 858.450 583.050 859.050 ;
        RECT 572.400 857.400 583.050 858.450 ;
        RECT 496.950 856.950 499.050 857.400 ;
        RECT 568.950 856.950 571.050 857.400 ;
        RECT 580.950 856.950 583.050 857.400 ;
        RECT 598.950 858.450 601.050 859.050 ;
        RECT 643.950 858.450 646.050 859.050 ;
        RECT 598.950 857.400 646.050 858.450 ;
        RECT 598.950 856.950 601.050 857.400 ;
        RECT 643.950 856.950 646.050 857.400 ;
        RECT 670.950 858.450 673.050 859.050 ;
        RECT 697.950 858.450 700.050 859.050 ;
        RECT 727.800 858.450 729.900 859.050 ;
        RECT 670.950 857.400 700.050 858.450 ;
        RECT 670.950 856.950 673.050 857.400 ;
        RECT 697.950 856.950 700.050 857.400 ;
        RECT 707.400 857.400 729.900 858.450 ;
        RECT 136.950 855.450 139.050 856.050 ;
        RECT 151.950 855.450 154.050 856.050 ;
        RECT 184.950 855.450 187.050 856.050 ;
        RECT 250.950 855.450 253.050 856.050 ;
        RECT 136.950 854.400 253.050 855.450 ;
        RECT 136.950 853.950 139.050 854.400 ;
        RECT 151.950 853.950 154.050 854.400 ;
        RECT 184.950 853.950 187.050 854.400 ;
        RECT 250.950 853.950 253.050 854.400 ;
        RECT 262.950 855.450 265.050 856.050 ;
        RECT 274.950 855.450 277.050 856.050 ;
        RECT 262.950 854.400 277.050 855.450 ;
        RECT 262.950 853.950 265.050 854.400 ;
        RECT 274.950 853.950 277.050 854.400 ;
        RECT 364.950 855.450 367.050 856.050 ;
        RECT 397.950 855.450 400.050 856.050 ;
        RECT 364.950 854.400 400.050 855.450 ;
        RECT 364.950 853.950 367.050 854.400 ;
        RECT 397.950 853.950 400.050 854.400 ;
        RECT 424.950 855.450 427.050 856.050 ;
        RECT 442.950 855.450 445.050 856.050 ;
        RECT 469.950 855.450 472.050 856.050 ;
        RECT 424.950 854.400 472.050 855.450 ;
        RECT 424.950 853.950 427.050 854.400 ;
        RECT 442.950 853.950 445.050 854.400 ;
        RECT 469.950 853.950 472.050 854.400 ;
        RECT 487.950 855.450 490.050 856.050 ;
        RECT 493.950 855.450 496.050 856.050 ;
        RECT 487.950 854.400 496.050 855.450 ;
        RECT 487.950 853.950 490.050 854.400 ;
        RECT 493.950 853.950 496.050 854.400 ;
        RECT 557.100 855.450 559.200 856.050 ;
        RECT 562.950 855.450 565.050 856.050 ;
        RECT 557.100 854.400 565.050 855.450 ;
        RECT 557.100 853.950 559.200 854.400 ;
        RECT 562.950 853.950 565.050 854.400 ;
        RECT 649.950 855.450 652.050 856.050 ;
        RECT 685.950 855.450 688.050 856.050 ;
        RECT 707.400 855.450 708.450 857.400 ;
        RECT 727.800 856.950 729.900 857.400 ;
        RECT 731.100 858.450 733.200 859.050 ;
        RECT 799.950 858.450 802.050 859.050 ;
        RECT 731.100 858.000 852.450 858.450 ;
        RECT 731.100 857.400 853.050 858.000 ;
        RECT 731.100 856.950 733.200 857.400 ;
        RECT 799.950 856.950 802.050 857.400 ;
        RECT 649.950 854.400 708.450 855.450 ;
        RECT 709.950 855.450 712.050 856.050 ;
        RECT 718.800 855.450 720.900 856.050 ;
        RECT 709.950 854.400 720.900 855.450 ;
        RECT 649.950 853.950 652.050 854.400 ;
        RECT 685.950 853.950 688.050 854.400 ;
        RECT 709.950 853.950 712.050 854.400 ;
        RECT 718.800 853.950 720.900 854.400 ;
        RECT 722.100 855.450 724.200 856.050 ;
        RECT 757.950 855.450 760.050 856.050 ;
        RECT 722.100 854.400 760.050 855.450 ;
        RECT 722.100 853.950 724.200 854.400 ;
        RECT 757.950 853.950 760.050 854.400 ;
        RECT 763.950 855.450 766.050 856.050 ;
        RECT 805.950 855.450 808.050 856.050 ;
        RECT 763.950 854.400 808.050 855.450 ;
        RECT 763.950 853.950 766.050 854.400 ;
        RECT 805.950 853.950 808.050 854.400 ;
        RECT 817.950 855.450 820.050 856.050 ;
        RECT 832.950 855.450 835.050 856.050 ;
        RECT 817.950 854.400 835.050 855.450 ;
        RECT 817.950 853.950 820.050 854.400 ;
        RECT 832.950 853.950 835.050 854.400 ;
        RECT 850.950 853.950 853.050 857.400 ;
        RECT 196.950 852.450 199.050 853.050 ;
        RECT 205.950 852.450 208.050 853.050 ;
        RECT 196.950 851.400 208.050 852.450 ;
        RECT 196.950 850.950 199.050 851.400 ;
        RECT 205.950 850.950 208.050 851.400 ;
        RECT 223.950 852.450 226.050 853.050 ;
        RECT 337.950 852.450 340.050 853.050 ;
        RECT 406.950 852.450 409.050 853.050 ;
        RECT 430.950 852.450 433.050 853.050 ;
        RECT 223.950 851.400 433.050 852.450 ;
        RECT 223.950 850.950 226.050 851.400 ;
        RECT 337.950 850.950 340.050 851.400 ;
        RECT 406.950 850.950 409.050 851.400 ;
        RECT 430.950 850.950 433.050 851.400 ;
        RECT 445.950 852.450 448.050 853.050 ;
        RECT 508.950 852.450 511.050 853.050 ;
        RECT 514.950 852.450 517.050 853.050 ;
        RECT 550.950 852.450 553.050 852.900 ;
        RECT 445.950 851.400 498.450 852.450 ;
        RECT 445.950 850.950 448.050 851.400 ;
        RECT 16.950 849.450 19.050 850.050 ;
        RECT 34.950 849.450 37.050 850.050 ;
        RECT 16.950 848.400 37.050 849.450 ;
        RECT 16.950 847.950 19.050 848.400 ;
        RECT 34.950 847.950 37.050 848.400 ;
        RECT 64.950 849.450 67.050 850.050 ;
        RECT 82.950 849.450 85.050 850.050 ;
        RECT 64.950 848.400 85.050 849.450 ;
        RECT 64.950 847.950 67.050 848.400 ;
        RECT 82.950 847.950 85.050 848.400 ;
        RECT 112.950 849.450 115.050 850.050 ;
        RECT 181.950 849.450 184.050 850.050 ;
        RECT 187.950 849.450 190.050 850.050 ;
        RECT 112.950 848.400 190.050 849.450 ;
        RECT 112.950 847.950 115.050 848.400 ;
        RECT 181.950 847.950 184.050 848.400 ;
        RECT 187.950 847.950 190.050 848.400 ;
        RECT 226.950 849.450 229.050 850.050 ;
        RECT 304.950 849.450 307.050 850.050 ;
        RECT 226.950 848.400 307.050 849.450 ;
        RECT 226.950 847.950 229.050 848.400 ;
        RECT 304.950 847.950 307.050 848.400 ;
        RECT 361.950 849.450 364.050 850.050 ;
        RECT 382.950 849.450 385.050 850.050 ;
        RECT 361.950 848.400 385.050 849.450 ;
        RECT 361.950 847.950 364.050 848.400 ;
        RECT 382.950 847.950 385.050 848.400 ;
        RECT 397.950 849.450 400.050 850.050 ;
        RECT 469.950 849.450 472.050 850.050 ;
        RECT 397.950 848.400 472.050 849.450 ;
        RECT 497.400 849.450 498.450 851.400 ;
        RECT 508.950 851.400 553.050 852.450 ;
        RECT 508.950 850.950 511.050 851.400 ;
        RECT 514.950 850.950 517.050 851.400 ;
        RECT 550.950 850.800 553.050 851.400 ;
        RECT 571.950 852.450 574.050 853.050 ;
        RECT 592.950 852.450 595.050 853.050 ;
        RECT 571.950 851.400 595.050 852.450 ;
        RECT 571.950 850.950 574.050 851.400 ;
        RECT 592.950 850.950 595.050 851.400 ;
        RECT 619.950 852.450 622.050 853.050 ;
        RECT 715.950 852.450 718.050 853.050 ;
        RECT 619.950 851.400 718.050 852.450 ;
        RECT 619.950 850.950 622.050 851.400 ;
        RECT 715.950 850.950 718.050 851.400 ;
        RECT 749.100 852.450 751.200 853.050 ;
        RECT 775.950 852.450 778.050 853.050 ;
        RECT 749.100 851.400 778.050 852.450 ;
        RECT 749.100 850.950 751.200 851.400 ;
        RECT 775.950 850.950 778.050 851.400 ;
        RECT 835.950 852.450 838.050 853.050 ;
        RECT 865.950 852.450 868.050 853.050 ;
        RECT 835.950 851.400 868.050 852.450 ;
        RECT 835.950 850.950 838.050 851.400 ;
        RECT 865.950 850.950 868.050 851.400 ;
        RECT 544.950 849.450 547.050 850.050 ;
        RECT 497.400 848.400 547.050 849.450 ;
        RECT 397.950 847.950 400.050 848.400 ;
        RECT 469.950 847.950 472.050 848.400 ;
        RECT 544.950 847.950 547.050 848.400 ;
        RECT 565.950 849.450 568.050 850.050 ;
        RECT 577.800 849.450 579.900 850.050 ;
        RECT 565.950 848.400 579.900 849.450 ;
        RECT 565.950 847.950 568.050 848.400 ;
        RECT 577.800 847.950 579.900 848.400 ;
        RECT 581.100 849.450 583.200 850.050 ;
        RECT 631.950 849.450 634.050 850.050 ;
        RECT 655.950 849.450 658.050 850.050 ;
        RECT 581.100 848.400 658.050 849.450 ;
        RECT 581.100 847.950 583.200 848.400 ;
        RECT 193.950 846.450 196.050 847.050 ;
        RECT 202.950 846.450 205.050 847.050 ;
        RECT 193.950 845.400 205.050 846.450 ;
        RECT 193.950 844.950 196.050 845.400 ;
        RECT 202.950 844.950 205.050 845.400 ;
        RECT 250.950 846.450 253.050 847.050 ;
        RECT 268.950 846.450 271.050 847.050 ;
        RECT 448.950 846.450 451.050 847.050 ;
        RECT 250.950 845.400 267.450 846.450 ;
        RECT 250.950 844.950 253.050 845.400 ;
        RECT 16.950 841.950 19.050 844.050 ;
        RECT 22.950 841.950 25.050 844.050 ;
        RECT 34.950 841.950 37.050 844.050 ;
        RECT 40.950 841.950 43.050 844.050 ;
        RECT 64.950 841.950 67.050 844.050 ;
        RECT 70.950 841.950 73.050 844.050 ;
        RECT 82.950 841.950 85.050 844.050 ;
        RECT 88.950 841.950 91.050 844.050 ;
        RECT 94.950 841.950 100.050 844.050 ;
        RECT 112.950 841.950 115.050 844.050 ;
        RECT 118.950 841.950 121.050 844.050 ;
        RECT 124.950 843.450 127.050 844.050 ;
        RECT 133.950 843.450 136.050 844.050 ;
        RECT 124.950 842.400 136.050 843.450 ;
        RECT 124.950 841.950 127.050 842.400 ;
        RECT 133.950 841.950 136.050 842.400 ;
        RECT 151.950 841.950 154.050 844.050 ;
        RECT 157.950 841.950 160.050 844.050 ;
        RECT 175.950 841.950 178.050 844.050 ;
        RECT 181.950 841.950 184.050 844.050 ;
        RECT 238.950 841.950 241.050 844.050 ;
        RECT 244.950 841.950 247.050 844.050 ;
        RECT 266.400 841.050 267.450 845.400 ;
        RECT 268.950 845.400 291.450 846.450 ;
        RECT 268.950 844.950 271.050 845.400 ;
        RECT 290.400 841.050 291.450 845.400 ;
        RECT 448.950 845.400 459.450 846.450 ;
        RECT 448.950 844.950 451.050 845.400 ;
        RECT 16.950 838.950 19.050 840.750 ;
        RECT 22.950 838.950 25.050 840.750 ;
        RECT 34.950 838.950 37.050 840.750 ;
        RECT 40.950 838.950 43.050 840.750 ;
        RECT 64.950 838.950 67.050 840.750 ;
        RECT 70.950 838.950 73.050 840.750 ;
        RECT 82.950 838.950 85.050 840.750 ;
        RECT 88.950 838.950 91.050 840.750 ;
        RECT 112.950 838.950 115.050 840.750 ;
        RECT 118.950 838.950 121.050 840.750 ;
        RECT 133.950 838.950 136.050 840.750 ;
        RECT 151.950 838.950 154.050 840.750 ;
        RECT 157.950 838.950 160.050 840.750 ;
        RECT 175.950 838.950 178.050 840.750 ;
        RECT 181.950 838.950 184.050 840.750 ;
        RECT 187.950 840.450 190.050 841.050 ;
        RECT 199.950 840.450 202.050 841.050 ;
        RECT 187.950 839.400 202.050 840.450 ;
        RECT 187.950 838.950 190.050 839.400 ;
        RECT 199.950 838.950 202.050 839.400 ;
        RECT 205.950 840.450 208.050 841.050 ;
        RECT 220.950 840.450 223.050 841.050 ;
        RECT 205.950 839.400 223.050 840.450 ;
        RECT 205.950 838.950 208.050 839.400 ;
        RECT 220.950 838.950 223.050 839.400 ;
        RECT 238.950 838.950 241.050 840.750 ;
        RECT 244.950 838.950 247.050 840.750 ;
        RECT 259.950 838.950 262.050 841.050 ;
        RECT 265.950 838.950 268.050 841.050 ;
        RECT 271.950 838.950 274.050 841.050 ;
        RECT 289.950 838.950 292.050 841.050 ;
        RECT 298.950 838.950 301.050 841.050 ;
        RECT 313.950 838.950 316.050 841.050 ;
        RECT 319.950 838.950 322.050 844.050 ;
        RECT 364.950 841.950 367.050 844.050 ;
        RECT 370.950 841.950 373.050 844.050 ;
        RECT 388.950 841.950 391.050 844.050 ;
        RECT 394.950 841.950 397.050 844.050 ;
        RECT 397.950 841.950 400.050 844.050 ;
        RECT 406.950 841.950 409.050 844.050 ;
        RECT 412.950 841.950 415.050 844.050 ;
        RECT 430.950 841.950 433.050 844.050 ;
        RECT 436.950 843.450 439.050 844.050 ;
        RECT 441.000 843.450 445.050 844.050 ;
        RECT 436.950 842.400 445.050 843.450 ;
        RECT 436.950 841.950 439.050 842.400 ;
        RECT 441.000 841.950 445.050 842.400 ;
        RECT 458.400 841.050 459.450 845.400 ;
        RECT 608.400 844.050 609.450 848.400 ;
        RECT 631.950 847.950 634.050 848.400 ;
        RECT 655.950 847.950 658.050 848.400 ;
        RECT 661.950 849.450 664.050 850.050 ;
        RECT 688.950 849.450 691.050 850.050 ;
        RECT 661.950 848.400 691.050 849.450 ;
        RECT 661.950 847.950 664.050 848.400 ;
        RECT 688.950 847.950 691.050 848.400 ;
        RECT 805.950 849.450 808.050 850.050 ;
        RECT 859.950 849.450 862.050 850.050 ;
        RECT 871.950 849.450 874.050 850.050 ;
        RECT 898.950 849.450 901.050 850.050 ;
        RECT 805.950 848.400 901.050 849.450 ;
        RECT 805.950 847.950 808.050 848.400 ;
        RECT 859.950 847.950 862.050 848.400 ;
        RECT 871.950 847.950 874.050 848.400 ;
        RECT 898.950 847.950 901.050 848.400 ;
        RECT 718.950 846.450 721.050 847.050 ;
        RECT 736.950 846.450 739.050 847.050 ;
        RECT 710.400 845.400 721.050 846.450 ;
        RECT 469.950 843.450 472.050 844.050 ;
        RECT 481.950 843.450 484.050 844.050 ;
        RECT 469.950 842.400 484.050 843.450 ;
        RECT 469.950 841.950 472.050 842.400 ;
        RECT 481.950 841.950 484.050 842.400 ;
        RECT 496.950 841.950 499.050 844.050 ;
        RECT 523.950 841.950 526.050 844.050 ;
        RECT 529.950 841.950 532.050 844.050 ;
        RECT 535.950 843.450 538.050 844.050 ;
        RECT 544.950 843.450 547.050 844.050 ;
        RECT 535.950 842.400 547.050 843.450 ;
        RECT 535.950 841.950 538.050 842.400 ;
        RECT 544.950 841.950 547.050 842.400 ;
        RECT 550.950 843.450 553.050 844.050 ;
        RECT 559.950 843.450 562.050 844.050 ;
        RECT 550.950 842.400 562.050 843.450 ;
        RECT 550.950 841.950 553.050 842.400 ;
        RECT 559.950 841.950 562.050 842.400 ;
        RECT 565.950 841.950 568.050 844.050 ;
        RECT 583.950 841.950 586.050 844.050 ;
        RECT 589.950 841.950 592.050 844.050 ;
        RECT 601.950 843.450 606.000 844.050 ;
        RECT 607.950 843.450 610.050 844.050 ;
        RECT 601.950 842.400 610.050 843.450 ;
        RECT 601.950 841.950 606.000 842.400 ;
        RECT 607.950 841.950 610.050 842.400 ;
        RECT 613.950 841.950 616.050 844.050 ;
        RECT 658.950 841.950 661.050 844.050 ;
        RECT 673.950 841.950 676.050 844.050 ;
        RECT 679.950 841.950 682.050 844.050 ;
        RECT 703.950 841.950 706.050 844.050 ;
        RECT 325.950 838.950 328.050 841.050 ;
        RECT 331.950 840.450 334.050 841.050 ;
        RECT 340.950 840.450 343.050 841.050 ;
        RECT 331.950 839.400 343.050 840.450 ;
        RECT 331.950 838.950 334.050 839.400 ;
        RECT 340.950 838.950 343.050 839.400 ;
        RECT 364.950 838.950 367.050 840.750 ;
        RECT 370.950 838.950 373.050 840.750 ;
        RECT 388.950 838.950 391.050 840.750 ;
        RECT 394.950 838.950 397.050 840.750 ;
        RECT 406.950 838.950 409.050 840.750 ;
        RECT 412.950 838.950 415.050 840.750 ;
        RECT 430.950 838.950 433.050 840.750 ;
        RECT 436.950 838.950 439.050 840.750 ;
        RECT 451.950 838.950 454.050 841.050 ;
        RECT 457.950 838.950 460.050 841.050 ;
        RECT 463.950 838.950 466.050 841.050 ;
        RECT 481.950 838.950 484.050 840.750 ;
        RECT 496.950 838.950 499.050 840.750 ;
        RECT 502.950 838.950 505.050 840.750 ;
        RECT 523.950 838.950 526.050 840.750 ;
        RECT 529.950 838.950 532.050 840.750 ;
        RECT 544.950 838.950 547.050 840.750 ;
        RECT 559.950 838.950 562.050 840.750 ;
        RECT 565.950 838.950 568.050 840.750 ;
        RECT 583.950 838.950 586.050 840.750 ;
        RECT 589.950 838.950 592.050 840.750 ;
        RECT 607.950 838.950 610.050 840.750 ;
        RECT 613.950 838.950 616.050 840.750 ;
        RECT 619.950 840.450 622.050 841.050 ;
        RECT 631.950 840.450 634.050 841.050 ;
        RECT 619.950 839.400 634.050 840.450 ;
        RECT 619.950 838.950 622.050 839.400 ;
        RECT 631.950 838.950 634.050 839.400 ;
        RECT 637.950 838.950 646.050 841.050 ;
        RECT 658.950 838.950 661.050 840.750 ;
        RECT 673.950 838.950 676.050 840.750 ;
        RECT 679.950 838.950 682.050 840.750 ;
        RECT 697.950 838.950 700.050 840.750 ;
        RECT 703.950 838.950 706.050 840.750 ;
        RECT 710.400 838.050 711.450 845.400 ;
        RECT 718.950 844.950 721.050 845.400 ;
        RECT 722.400 845.400 739.050 846.450 ;
        RECT 722.400 841.050 723.450 845.400 ;
        RECT 736.950 844.950 739.050 845.400 ;
        RECT 742.950 841.950 745.050 844.050 ;
        RECT 748.950 841.950 751.050 844.050 ;
        RECT 715.950 838.950 718.050 841.050 ;
        RECT 721.950 838.950 724.050 841.050 ;
        RECT 727.950 838.950 730.050 841.050 ;
        RECT 742.950 838.950 745.050 840.750 ;
        RECT 748.950 838.950 751.050 840.750 ;
        RECT 766.950 838.950 769.050 841.050 ;
        RECT 775.950 840.450 778.050 844.050 ;
        RECT 799.950 841.950 802.050 844.050 ;
        RECT 811.950 841.950 814.050 844.050 ;
        RECT 817.950 841.950 820.050 844.050 ;
        RECT 859.950 841.950 862.050 844.050 ;
        RECT 865.950 843.450 868.050 844.050 ;
        RECT 870.000 843.450 874.050 844.050 ;
        RECT 865.950 842.400 874.050 843.450 ;
        RECT 865.950 841.950 868.050 842.400 ;
        RECT 870.000 841.950 874.050 842.400 ;
        RECT 877.950 841.950 880.050 844.050 ;
        RECT 883.950 841.950 886.050 844.050 ;
        RECT 898.950 841.950 901.050 844.050 ;
        RECT 904.950 841.950 907.050 844.050 ;
        RECT 787.950 840.450 790.050 841.050 ;
        RECT 775.950 839.400 790.050 840.450 ;
        RECT 775.950 838.950 778.050 839.400 ;
        RECT 787.950 838.950 790.050 839.400 ;
        RECT 793.950 838.950 796.050 840.750 ;
        RECT 799.950 838.950 802.050 840.750 ;
        RECT 811.950 838.950 814.050 840.750 ;
        RECT 817.950 838.950 820.050 840.750 ;
        RECT 823.950 840.450 826.050 841.050 ;
        RECT 838.950 840.450 841.050 841.050 ;
        RECT 843.000 840.450 847.050 841.050 ;
        RECT 823.950 839.400 847.050 840.450 ;
        RECT 823.950 838.950 826.050 839.400 ;
        RECT 838.950 838.950 841.050 839.400 ;
        RECT 843.000 838.950 847.050 839.400 ;
        RECT 859.950 838.950 862.050 840.750 ;
        RECT 865.950 838.950 868.050 840.750 ;
        RECT 877.950 838.950 880.050 840.750 ;
        RECT 883.950 838.950 886.050 840.750 ;
        RECT 898.950 838.950 901.050 840.750 ;
        RECT 904.950 838.950 907.050 840.750 ;
        RECT 874.950 838.050 877.050 838.200 ;
        RECT 13.950 836.250 16.050 838.050 ;
        RECT 19.950 836.250 22.050 838.050 ;
        RECT 37.950 836.250 40.050 838.050 ;
        RECT 43.950 836.250 46.050 838.050 ;
        RECT 61.950 836.250 64.050 838.050 ;
        RECT 67.950 836.250 70.050 838.050 ;
        RECT 85.950 836.250 88.050 838.050 ;
        RECT 91.950 836.250 94.050 838.050 ;
        RECT 109.950 836.250 112.050 838.050 ;
        RECT 115.950 836.250 118.050 838.050 ;
        RECT 136.950 836.250 139.050 838.050 ;
        RECT 148.950 836.250 151.050 838.050 ;
        RECT 154.950 836.250 157.050 838.050 ;
        RECT 178.950 836.250 181.050 838.050 ;
        RECT 184.950 836.250 187.050 838.050 ;
        RECT 199.950 835.950 202.050 837.750 ;
        RECT 220.950 835.950 223.050 837.750 ;
        RECT 241.950 836.250 244.050 838.050 ;
        RECT 293.250 837.750 295.050 838.050 ;
        RECT 259.950 835.950 262.050 837.750 ;
        RECT 265.950 835.950 268.050 837.750 ;
        RECT 271.950 835.950 274.050 837.750 ;
        RECT 289.950 836.250 292.050 837.750 ;
        RECT 292.950 836.250 295.050 837.750 ;
        RECT 289.950 835.950 291.750 836.250 ;
        RECT 298.950 835.950 301.050 837.750 ;
        RECT 313.950 835.950 316.050 837.750 ;
        RECT 319.950 835.950 322.050 837.750 ;
        RECT 325.950 835.950 328.050 837.750 ;
        RECT 340.950 835.950 343.050 837.750 ;
        RECT 346.950 836.250 349.050 838.050 ;
        RECT 361.950 836.250 364.050 838.050 ;
        RECT 367.950 836.250 370.050 838.050 ;
        RECT 385.950 836.250 388.050 838.050 ;
        RECT 391.950 836.250 394.050 838.050 ;
        RECT 409.950 836.250 412.050 838.050 ;
        RECT 433.950 836.250 436.050 838.050 ;
        RECT 439.950 836.250 442.050 838.050 ;
        RECT 451.950 835.950 454.050 837.750 ;
        RECT 457.950 835.950 460.050 837.750 ;
        RECT 463.950 835.950 466.050 837.750 ;
        RECT 478.950 836.250 481.050 838.050 ;
        RECT 499.950 836.250 502.050 838.050 ;
        RECT 520.950 836.250 523.050 838.050 ;
        RECT 526.950 836.250 529.050 838.050 ;
        RECT 547.950 836.250 550.050 838.050 ;
        RECT 562.950 836.250 565.050 838.050 ;
        RECT 580.950 836.250 583.050 838.050 ;
        RECT 586.950 836.250 589.050 838.050 ;
        RECT 604.950 836.250 607.050 838.050 ;
        RECT 610.950 836.250 613.050 838.050 ;
        RECT 635.250 837.750 637.050 838.050 ;
        RECT 631.950 836.250 634.050 837.750 ;
        RECT 634.950 836.250 637.050 837.750 ;
        RECT 631.950 835.950 633.750 836.250 ;
        RECT 640.950 835.950 643.050 837.750 ;
        RECT 655.950 836.250 658.050 838.050 ;
        RECT 676.950 836.250 679.050 838.050 ;
        RECT 682.950 836.250 685.050 838.050 ;
        RECT 700.950 836.250 703.050 838.050 ;
        RECT 706.950 836.400 711.450 838.050 ;
        RECT 706.950 835.950 711.000 836.400 ;
        RECT 715.950 835.950 718.050 837.750 ;
        RECT 721.950 835.950 724.050 837.750 ;
        RECT 727.950 835.950 730.050 837.750 ;
        RECT 745.950 836.250 748.050 838.050 ;
        RECT 751.950 836.250 754.050 838.050 ;
        RECT 772.950 837.750 774.750 838.050 ;
        RECT 766.950 835.950 769.050 837.750 ;
        RECT 772.950 836.250 775.050 837.750 ;
        RECT 775.950 836.250 778.050 837.750 ;
        RECT 796.950 836.250 799.050 838.050 ;
        RECT 814.950 836.250 817.050 838.050 ;
        RECT 820.950 836.250 823.050 838.050 ;
        RECT 776.250 835.950 778.050 836.250 ;
        RECT 838.950 835.950 841.050 837.750 ;
        RECT 862.950 836.250 865.050 838.050 ;
        RECT 871.950 836.100 877.050 838.050 ;
        RECT 880.950 836.250 883.050 838.050 ;
        RECT 901.950 836.250 904.050 838.050 ;
        RECT 871.950 835.950 876.000 836.100 ;
        RECT 13.950 829.950 16.050 835.050 ;
        RECT 19.950 832.950 22.050 835.050 ;
        RECT 37.950 832.950 40.050 835.050 ;
        RECT 43.950 832.950 49.050 835.050 ;
        RECT 61.950 829.950 64.050 835.050 ;
        RECT 67.950 832.950 70.050 835.050 ;
        RECT 85.950 832.950 88.050 835.050 ;
        RECT 91.950 834.450 94.050 835.050 ;
        RECT 96.000 834.450 100.050 835.050 ;
        RECT 91.950 833.400 100.050 834.450 ;
        RECT 91.950 832.950 94.050 833.400 ;
        RECT 96.000 832.950 100.050 833.400 ;
        RECT 103.950 834.450 108.000 835.050 ;
        RECT 109.950 834.450 112.050 835.050 ;
        RECT 103.950 833.400 112.050 834.450 ;
        RECT 103.950 832.950 108.000 833.400 ;
        RECT 109.950 832.950 112.050 833.400 ;
        RECT 115.950 832.950 118.050 835.050 ;
        RECT 136.950 832.950 139.050 835.050 ;
        RECT 148.950 832.950 151.050 835.050 ;
        RECT 154.950 832.950 157.050 835.050 ;
        RECT 172.950 834.450 177.000 835.050 ;
        RECT 178.950 834.450 181.050 835.050 ;
        RECT 172.950 833.400 181.050 834.450 ;
        RECT 172.950 832.950 177.000 833.400 ;
        RECT 178.950 832.950 181.050 833.400 ;
        RECT 184.950 832.950 187.050 835.050 ;
        RECT 196.950 833.250 199.050 835.050 ;
        RECT 202.950 833.250 205.050 835.050 ;
        RECT 217.950 833.250 220.050 835.050 ;
        RECT 223.950 833.250 226.050 835.050 ;
        RECT 229.950 834.450 232.050 835.050 ;
        RECT 241.950 834.450 244.050 835.050 ;
        RECT 229.950 833.400 244.050 834.450 ;
        RECT 229.950 832.950 232.050 833.400 ;
        RECT 241.950 832.950 244.050 833.400 ;
        RECT 262.950 833.250 265.050 835.050 ;
        RECT 268.950 833.250 271.050 835.050 ;
        RECT 292.950 832.950 295.050 835.050 ;
        RECT 316.950 833.250 319.050 835.050 ;
        RECT 322.950 833.250 325.050 835.050 ;
        RECT 352.950 834.450 355.050 835.050 ;
        RECT 361.950 834.450 364.050 835.050 ;
        RECT 352.950 833.400 364.050 834.450 ;
        RECT 352.950 832.950 355.050 833.400 ;
        RECT 361.950 832.950 364.050 833.400 ;
        RECT 367.950 832.950 370.050 835.050 ;
        RECT 385.950 832.950 388.050 835.050 ;
        RECT 391.950 832.950 394.050 835.050 ;
        RECT 409.950 832.950 412.050 835.050 ;
        RECT 418.950 834.450 421.050 835.050 ;
        RECT 424.950 834.450 427.050 835.050 ;
        RECT 418.950 833.400 427.050 834.450 ;
        RECT 418.950 832.950 421.050 833.400 ;
        RECT 424.950 832.950 427.050 833.400 ;
        RECT 433.950 832.950 436.050 835.050 ;
        RECT 439.950 832.950 442.050 835.050 ;
        RECT 454.950 833.250 457.050 835.050 ;
        RECT 460.950 833.250 463.050 835.050 ;
        RECT 478.950 832.950 481.050 835.050 ;
        RECT 499.950 832.950 502.050 835.050 ;
        RECT 505.950 834.450 508.050 835.050 ;
        RECT 520.950 834.450 523.050 835.050 ;
        RECT 505.950 833.400 523.050 834.450 ;
        RECT 505.950 832.950 508.050 833.400 ;
        RECT 520.950 832.950 523.050 833.400 ;
        RECT 526.950 834.450 529.050 835.050 ;
        RECT 541.950 834.450 544.050 835.050 ;
        RECT 526.950 833.400 544.050 834.450 ;
        RECT 526.950 832.950 529.050 833.400 ;
        RECT 541.950 832.950 544.050 833.400 ;
        RECT 547.950 832.950 550.050 835.050 ;
        RECT 553.950 834.450 556.050 835.050 ;
        RECT 562.950 834.450 565.050 835.050 ;
        RECT 553.950 833.400 565.050 834.450 ;
        RECT 553.950 832.950 556.050 833.400 ;
        RECT 562.950 832.950 565.050 833.400 ;
        RECT 568.950 834.450 571.050 835.050 ;
        RECT 580.950 834.450 583.050 835.050 ;
        RECT 568.950 833.400 583.050 834.450 ;
        RECT 568.950 832.950 571.050 833.400 ;
        RECT 580.950 832.950 583.050 833.400 ;
        RECT 70.950 831.450 73.050 832.050 ;
        RECT 76.950 831.450 79.050 832.050 ;
        RECT 70.950 830.400 79.050 831.450 ;
        RECT 70.950 829.950 73.050 830.400 ;
        RECT 76.950 829.950 79.050 830.400 ;
        RECT 25.950 828.450 28.050 829.050 ;
        RECT 37.950 828.450 40.050 829.050 ;
        RECT 25.950 827.400 40.050 828.450 ;
        RECT 25.950 826.950 28.050 827.400 ;
        RECT 37.950 826.950 40.050 827.400 ;
        RECT 91.950 828.450 94.050 829.050 ;
        RECT 115.950 828.450 118.050 829.050 ;
        RECT 124.950 828.450 127.050 829.050 ;
        RECT 155.400 828.450 156.450 832.950 ;
        RECT 196.950 829.950 199.050 832.050 ;
        RECT 202.950 829.950 205.050 832.050 ;
        RECT 217.950 829.950 220.050 832.050 ;
        RECT 223.950 829.950 226.050 832.050 ;
        RECT 262.950 828.450 265.050 832.050 ;
        RECT 268.950 829.950 271.050 832.050 ;
        RECT 316.950 829.950 319.050 832.050 ;
        RECT 322.950 829.950 325.050 832.050 ;
        RECT 91.950 827.400 127.050 828.450 ;
        RECT 91.950 826.950 94.050 827.400 ;
        RECT 115.950 826.950 118.050 827.400 ;
        RECT 124.950 826.950 127.050 827.400 ;
        RECT 128.400 827.400 156.450 828.450 ;
        RECT 233.400 827.400 265.050 828.450 ;
        RECT 325.950 828.450 328.050 829.050 ;
        RECT 331.950 828.450 334.050 829.050 ;
        RECT 325.950 827.400 334.050 828.450 ;
        RECT 73.950 825.450 76.050 826.050 ;
        RECT 97.950 825.450 100.050 826.050 ;
        RECT 128.400 825.450 129.450 827.400 ;
        RECT 73.950 824.400 129.450 825.450 ;
        RECT 148.950 825.450 151.050 826.050 ;
        RECT 175.950 825.450 178.050 826.050 ;
        RECT 148.950 824.400 178.050 825.450 ;
        RECT 73.950 823.950 76.050 824.400 ;
        RECT 97.950 823.950 100.050 824.400 ;
        RECT 148.950 823.950 151.050 824.400 ;
        RECT 175.950 823.950 178.050 824.400 ;
        RECT 202.950 825.450 205.050 826.050 ;
        RECT 217.950 825.450 220.050 826.050 ;
        RECT 229.950 825.450 232.050 826.050 ;
        RECT 202.950 824.400 232.050 825.450 ;
        RECT 202.950 823.950 205.050 824.400 ;
        RECT 217.950 823.950 220.050 824.400 ;
        RECT 229.950 823.950 232.050 824.400 ;
        RECT 4.950 822.450 7.050 823.050 ;
        RECT 46.950 822.450 49.050 823.050 ;
        RECT 4.950 821.400 49.050 822.450 ;
        RECT 4.950 820.950 7.050 821.400 ;
        RECT 46.950 820.950 49.050 821.400 ;
        RECT 127.950 822.450 130.050 823.050 ;
        RECT 181.950 822.450 184.050 823.050 ;
        RECT 205.950 822.450 208.050 823.050 ;
        RECT 127.950 821.400 208.050 822.450 ;
        RECT 127.950 820.950 130.050 821.400 ;
        RECT 181.950 820.950 184.050 821.400 ;
        RECT 205.950 820.950 208.050 821.400 ;
        RECT 220.950 822.450 223.050 823.050 ;
        RECT 233.400 822.450 234.450 827.400 ;
        RECT 325.950 826.950 328.050 827.400 ;
        RECT 331.950 826.950 334.050 827.400 ;
        RECT 373.950 828.450 376.050 829.050 ;
        RECT 391.950 828.450 394.050 829.050 ;
        RECT 410.400 828.450 411.450 832.950 ;
        RECT 415.950 831.450 418.050 832.050 ;
        RECT 427.950 831.450 430.050 832.050 ;
        RECT 415.950 830.400 430.050 831.450 ;
        RECT 415.950 829.950 418.050 830.400 ;
        RECT 427.950 829.950 430.050 830.400 ;
        RECT 454.950 829.950 457.050 832.050 ;
        RECT 460.950 831.450 463.050 832.050 ;
        RECT 472.950 831.450 475.050 832.050 ;
        RECT 460.950 830.400 475.050 831.450 ;
        RECT 460.950 829.950 463.050 830.400 ;
        RECT 472.950 829.950 475.050 830.400 ;
        RECT 586.950 829.950 589.050 835.050 ;
        RECT 604.950 832.950 607.050 835.050 ;
        RECT 610.950 832.950 613.050 835.050 ;
        RECT 634.950 832.950 637.050 835.050 ;
        RECT 655.950 832.950 658.050 835.050 ;
        RECT 373.950 827.400 411.450 828.450 ;
        RECT 469.950 828.450 472.050 829.050 ;
        RECT 499.950 828.450 502.050 829.050 ;
        RECT 469.950 827.400 502.050 828.450 ;
        RECT 373.950 826.950 376.050 827.400 ;
        RECT 391.950 826.950 394.050 827.400 ;
        RECT 469.950 826.950 472.050 827.400 ;
        RECT 499.950 826.950 502.050 827.400 ;
        RECT 523.950 828.450 526.050 829.050 ;
        RECT 532.800 828.450 534.900 829.050 ;
        RECT 523.950 827.400 534.900 828.450 ;
        RECT 523.950 826.950 526.050 827.400 ;
        RECT 532.800 826.950 534.900 827.400 ;
        RECT 536.100 828.450 538.200 829.050 ;
        RECT 547.950 828.450 550.050 829.050 ;
        RECT 536.100 827.400 550.050 828.450 ;
        RECT 536.100 826.950 538.200 827.400 ;
        RECT 547.950 826.950 550.050 827.400 ;
        RECT 580.950 828.450 583.050 829.050 ;
        RECT 605.400 828.450 606.450 832.950 ;
        RECT 631.950 828.450 634.050 829.050 ;
        RECT 649.950 828.450 652.050 832.050 ;
        RECT 676.950 829.950 679.050 835.050 ;
        RECT 682.950 832.950 685.050 835.050 ;
        RECT 688.950 834.450 691.050 835.050 ;
        RECT 700.950 834.450 703.050 835.050 ;
        RECT 688.950 833.400 703.050 834.450 ;
        RECT 688.950 832.950 691.050 833.400 ;
        RECT 700.950 832.950 703.050 833.400 ;
        RECT 718.950 833.250 721.050 835.050 ;
        RECT 724.950 833.250 727.050 835.050 ;
        RECT 751.950 834.450 754.050 835.050 ;
        RECT 756.000 834.450 760.050 835.050 ;
        RECT 751.950 833.400 760.050 834.450 ;
        RECT 751.950 832.950 754.050 833.400 ;
        RECT 756.000 832.950 760.050 833.400 ;
        RECT 796.950 832.950 802.050 835.050 ;
        RECT 814.950 832.950 817.050 835.050 ;
        RECT 820.950 834.450 823.050 835.050 ;
        RECT 829.950 834.450 832.050 835.050 ;
        RECT 820.950 833.400 832.050 834.450 ;
        RECT 820.950 832.950 823.050 833.400 ;
        RECT 829.950 832.950 832.050 833.400 ;
        RECT 835.950 833.250 838.050 835.050 ;
        RECT 841.950 833.250 844.050 835.050 ;
        RECT 847.950 834.450 850.050 835.050 ;
        RECT 862.950 834.450 865.050 835.050 ;
        RECT 876.000 834.900 879.000 835.050 ;
        RECT 847.950 833.400 865.050 834.450 ;
        RECT 847.950 832.950 850.050 833.400 ;
        RECT 862.950 832.950 865.050 833.400 ;
        RECT 874.950 834.450 879.000 834.900 ;
        RECT 880.950 834.450 883.050 835.050 ;
        RECT 874.950 833.400 883.050 834.450 ;
        RECT 874.950 832.950 879.000 833.400 ;
        RECT 880.950 832.950 883.050 833.400 ;
        RECT 892.950 834.450 895.050 835.050 ;
        RECT 901.950 834.450 904.050 835.050 ;
        RECT 892.950 833.400 904.050 834.450 ;
        RECT 892.950 832.950 895.050 833.400 ;
        RECT 901.950 832.950 904.050 833.400 ;
        RECT 874.950 832.800 877.050 832.950 ;
        RECT 709.950 831.450 712.050 832.050 ;
        RECT 718.950 831.450 721.050 832.050 ;
        RECT 709.950 830.400 721.050 831.450 ;
        RECT 709.950 829.950 712.050 830.400 ;
        RECT 718.950 829.950 721.050 830.400 ;
        RECT 724.950 829.950 727.050 832.050 ;
        RECT 790.950 831.450 793.050 832.050 ;
        RECT 782.400 830.400 793.050 831.450 ;
        RECT 580.950 827.400 630.450 828.450 ;
        RECT 580.950 826.950 583.050 827.400 ;
        RECT 244.950 825.450 247.050 826.050 ;
        RECT 268.950 825.450 271.050 826.050 ;
        RECT 292.950 825.450 295.050 826.050 ;
        RECT 322.950 825.450 325.050 826.050 ;
        RECT 244.950 824.400 325.050 825.450 ;
        RECT 244.950 823.950 247.050 824.400 ;
        RECT 268.950 823.950 271.050 824.400 ;
        RECT 292.950 823.950 295.050 824.400 ;
        RECT 322.950 823.950 325.050 824.400 ;
        RECT 328.950 825.450 331.050 826.050 ;
        RECT 385.950 825.450 388.050 826.050 ;
        RECT 328.950 824.400 388.050 825.450 ;
        RECT 328.950 823.950 331.050 824.400 ;
        RECT 385.950 823.950 388.050 824.400 ;
        RECT 397.950 825.450 400.050 826.050 ;
        RECT 412.950 825.450 415.050 826.050 ;
        RECT 397.950 824.400 415.050 825.450 ;
        RECT 397.950 823.950 400.050 824.400 ;
        RECT 412.950 823.950 415.050 824.400 ;
        RECT 424.950 825.450 427.050 826.050 ;
        RECT 454.950 825.450 457.050 826.050 ;
        RECT 424.950 824.400 457.050 825.450 ;
        RECT 424.950 823.950 427.050 824.400 ;
        RECT 454.950 823.950 457.050 824.400 ;
        RECT 469.950 825.450 472.050 826.050 ;
        RECT 487.950 825.450 490.050 826.050 ;
        RECT 469.950 824.400 490.050 825.450 ;
        RECT 469.950 823.950 472.050 824.400 ;
        RECT 487.950 823.950 490.050 824.400 ;
        RECT 505.950 825.450 508.050 826.050 ;
        RECT 577.950 825.450 580.050 826.050 ;
        RECT 505.950 824.400 580.050 825.450 ;
        RECT 629.400 825.450 630.450 827.400 ;
        RECT 631.950 827.400 652.050 828.450 ;
        RECT 631.950 826.950 634.050 827.400 ;
        RECT 649.950 826.950 652.050 827.400 ;
        RECT 667.950 828.450 670.050 829.050 ;
        RECT 715.950 828.450 718.050 829.050 ;
        RECT 667.950 827.400 718.050 828.450 ;
        RECT 667.950 826.950 670.050 827.400 ;
        RECT 715.950 826.950 718.050 827.400 ;
        RECT 736.950 828.450 739.050 829.050 ;
        RECT 763.800 828.450 765.900 829.050 ;
        RECT 782.400 828.450 783.450 830.400 ;
        RECT 790.950 829.950 793.050 830.400 ;
        RECT 835.950 829.950 838.050 832.050 ;
        RECT 841.950 831.450 844.050 832.050 ;
        RECT 856.950 831.450 859.050 832.050 ;
        RECT 841.950 830.400 859.050 831.450 ;
        RECT 841.950 829.950 844.050 830.400 ;
        RECT 856.950 829.950 859.050 830.400 ;
        RECT 907.950 829.950 913.050 832.050 ;
        RECT 736.950 827.400 765.900 828.450 ;
        RECT 736.950 826.950 739.050 827.400 ;
        RECT 763.800 826.950 765.900 827.400 ;
        RECT 767.400 827.400 783.450 828.450 ;
        RECT 784.950 828.450 787.050 829.050 ;
        RECT 814.950 828.450 817.050 829.050 ;
        RECT 784.950 827.400 817.050 828.450 ;
        RECT 658.950 825.450 661.050 826.050 ;
        RECT 629.400 824.400 661.050 825.450 ;
        RECT 505.950 823.950 508.050 824.400 ;
        RECT 577.950 823.950 580.050 824.400 ;
        RECT 658.950 823.950 661.050 824.400 ;
        RECT 700.950 825.450 703.050 826.050 ;
        RECT 706.950 825.450 709.050 826.050 ;
        RECT 700.950 824.400 709.050 825.450 ;
        RECT 700.950 823.950 703.050 824.400 ;
        RECT 706.950 823.950 709.050 824.400 ;
        RECT 737.100 825.450 739.200 826.200 ;
        RECT 767.400 826.050 768.450 827.400 ;
        RECT 784.950 826.950 787.050 827.400 ;
        RECT 814.950 826.950 817.050 827.400 ;
        RECT 865.950 828.450 868.050 829.050 ;
        RECT 883.950 828.450 886.050 829.050 ;
        RECT 901.950 828.450 904.050 829.050 ;
        RECT 865.950 827.400 904.050 828.450 ;
        RECT 865.950 826.950 868.050 827.400 ;
        RECT 883.950 826.950 886.050 827.400 ;
        RECT 901.950 826.950 904.050 827.400 ;
        RECT 745.950 825.450 748.050 826.050 ;
        RECT 737.100 824.400 748.050 825.450 ;
        RECT 737.100 824.100 739.200 824.400 ;
        RECT 745.950 823.950 748.050 824.400 ;
        RECT 754.950 825.450 757.050 826.050 ;
        RECT 766.950 825.450 769.050 826.050 ;
        RECT 805.950 825.450 808.050 826.050 ;
        RECT 754.950 824.400 769.050 825.450 ;
        RECT 754.950 823.950 757.050 824.400 ;
        RECT 766.950 823.950 769.050 824.400 ;
        RECT 788.400 824.400 808.050 825.450 ;
        RECT 220.950 821.400 234.450 822.450 ;
        RECT 238.950 822.450 241.050 823.050 ;
        RECT 271.950 822.450 274.050 823.050 ;
        RECT 298.950 822.450 301.050 823.050 ;
        RECT 238.950 821.400 301.050 822.450 ;
        RECT 220.950 820.950 223.050 821.400 ;
        RECT 238.950 820.950 241.050 821.400 ;
        RECT 271.950 820.950 274.050 821.400 ;
        RECT 298.950 820.950 301.050 821.400 ;
        RECT 304.950 822.450 307.050 823.050 ;
        RECT 445.950 822.450 448.050 823.050 ;
        RECT 304.950 821.400 448.050 822.450 ;
        RECT 304.950 820.950 307.050 821.400 ;
        RECT 445.950 820.950 448.050 821.400 ;
        RECT 472.950 822.450 475.050 823.050 ;
        RECT 481.950 822.450 484.050 823.050 ;
        RECT 472.950 821.400 484.050 822.450 ;
        RECT 472.950 820.950 475.050 821.400 ;
        RECT 481.950 820.950 484.050 821.400 ;
        RECT 493.950 822.450 496.050 823.050 ;
        RECT 529.950 822.450 532.050 823.050 ;
        RECT 553.950 822.450 556.050 823.050 ;
        RECT 493.950 821.400 556.050 822.450 ;
        RECT 493.950 820.950 496.050 821.400 ;
        RECT 529.950 820.950 532.050 821.400 ;
        RECT 553.950 820.950 556.050 821.400 ;
        RECT 703.950 822.450 706.050 823.050 ;
        RECT 736.950 822.450 739.050 822.900 ;
        RECT 703.950 821.400 739.050 822.450 ;
        RECT 703.950 820.950 706.050 821.400 ;
        RECT 736.950 820.800 739.050 821.400 ;
        RECT 193.950 819.450 196.050 820.050 ;
        RECT 262.950 819.450 265.050 820.050 ;
        RECT 310.950 819.450 313.050 820.050 ;
        RECT 193.950 818.400 313.050 819.450 ;
        RECT 193.950 817.950 196.050 818.400 ;
        RECT 262.950 817.950 265.050 818.400 ;
        RECT 310.950 817.950 313.050 818.400 ;
        RECT 340.950 819.450 343.050 820.050 ;
        RECT 370.950 819.450 373.050 820.050 ;
        RECT 433.800 819.450 435.900 820.050 ;
        RECT 340.950 818.400 373.050 819.450 ;
        RECT 340.950 817.950 343.050 818.400 ;
        RECT 370.950 817.950 373.050 818.400 ;
        RECT 416.400 818.400 435.900 819.450 ;
        RECT 13.950 816.450 16.050 817.050 ;
        RECT 28.950 816.450 31.050 817.050 ;
        RECT 13.950 815.400 31.050 816.450 ;
        RECT 13.950 814.950 16.050 815.400 ;
        RECT 28.950 814.950 31.050 815.400 ;
        RECT 46.950 816.450 49.050 817.050 ;
        RECT 97.950 816.450 100.050 817.050 ;
        RECT 46.950 815.400 100.050 816.450 ;
        RECT 46.950 814.950 49.050 815.400 ;
        RECT 97.950 814.950 100.050 815.400 ;
        RECT 112.950 816.450 115.050 817.050 ;
        RECT 118.950 816.450 121.050 817.200 ;
        RECT 124.950 816.450 127.050 817.050 ;
        RECT 112.950 815.400 127.050 816.450 ;
        RECT 112.950 814.950 115.050 815.400 ;
        RECT 118.950 815.100 121.050 815.400 ;
        RECT 124.950 814.950 127.050 815.400 ;
        RECT 163.950 816.450 166.050 817.050 ;
        RECT 211.950 816.450 214.050 817.050 ;
        RECT 163.950 815.400 214.050 816.450 ;
        RECT 163.950 814.950 166.050 815.400 ;
        RECT 211.950 814.950 214.050 815.400 ;
        RECT 256.950 814.950 262.050 817.050 ;
        RECT 280.950 816.450 283.050 817.050 ;
        RECT 286.950 816.450 289.050 817.050 ;
        RECT 280.950 815.400 289.050 816.450 ;
        RECT 280.950 814.950 283.050 815.400 ;
        RECT 286.950 814.950 289.050 815.400 ;
        RECT 295.950 816.450 298.050 817.050 ;
        RECT 319.950 816.450 322.050 817.050 ;
        RECT 352.950 816.450 355.050 817.200 ;
        RECT 416.400 816.450 417.450 818.400 ;
        RECT 433.800 817.950 435.900 818.400 ;
        RECT 437.100 819.450 439.200 820.050 ;
        RECT 448.950 819.450 451.050 820.050 ;
        RECT 437.100 818.400 451.050 819.450 ;
        RECT 437.100 817.950 439.200 818.400 ;
        RECT 448.950 817.950 451.050 818.400 ;
        RECT 454.950 819.450 457.050 820.050 ;
        RECT 478.950 819.450 481.050 820.050 ;
        RECT 499.950 819.450 502.050 820.050 ;
        RECT 523.950 819.450 526.050 820.050 ;
        RECT 454.950 819.000 468.600 819.450 ;
        RECT 454.950 818.400 469.050 819.000 ;
        RECT 454.950 817.950 457.050 818.400 ;
        RECT 466.950 817.050 469.050 818.400 ;
        RECT 478.950 818.400 526.050 819.450 ;
        RECT 478.950 817.950 481.050 818.400 ;
        RECT 499.950 817.950 502.050 818.400 ;
        RECT 523.950 817.950 526.050 818.400 ;
        RECT 538.950 819.450 541.050 820.050 ;
        RECT 559.950 819.450 562.050 820.050 ;
        RECT 538.950 818.400 562.050 819.450 ;
        RECT 538.950 817.950 541.050 818.400 ;
        RECT 559.950 817.950 562.050 818.400 ;
        RECT 577.950 819.450 580.050 820.200 ;
        RECT 788.400 820.050 789.450 824.400 ;
        RECT 805.950 823.950 808.050 824.400 ;
        RECT 817.950 825.450 820.050 826.050 ;
        RECT 823.950 825.450 826.050 826.050 ;
        RECT 817.950 824.400 826.050 825.450 ;
        RECT 817.950 823.950 820.050 824.400 ;
        RECT 823.950 823.950 826.050 824.400 ;
        RECT 835.950 825.450 838.050 826.050 ;
        RECT 841.950 825.450 844.050 826.050 ;
        RECT 835.950 824.400 844.050 825.450 ;
        RECT 835.950 823.950 838.050 824.400 ;
        RECT 841.950 823.950 844.050 824.400 ;
        RECT 847.950 823.950 853.050 826.050 ;
        RECT 907.950 823.950 913.050 826.050 ;
        RECT 814.950 822.450 817.050 823.050 ;
        RECT 853.950 822.450 856.050 823.050 ;
        RECT 814.950 821.400 856.050 822.450 ;
        RECT 814.950 820.950 817.050 821.400 ;
        RECT 853.950 820.950 856.050 821.400 ;
        RECT 607.950 819.450 610.050 820.050 ;
        RECT 661.950 819.450 664.050 820.050 ;
        RECT 577.950 818.400 664.050 819.450 ;
        RECT 577.950 818.100 580.050 818.400 ;
        RECT 607.950 817.950 610.050 818.400 ;
        RECT 661.950 817.950 664.050 818.400 ;
        RECT 676.950 819.450 679.050 820.050 ;
        RECT 778.950 819.450 781.050 820.050 ;
        RECT 676.950 818.400 781.050 819.450 ;
        RECT 676.950 817.950 679.050 818.400 ;
        RECT 778.950 817.950 781.050 818.400 ;
        RECT 784.950 818.400 789.450 820.050 ;
        RECT 799.950 819.450 804.000 820.050 ;
        RECT 805.950 819.450 808.050 820.050 ;
        RECT 865.950 819.450 868.050 820.050 ;
        RECT 799.950 819.000 804.450 819.450 ;
        RECT 784.950 817.950 789.000 818.400 ;
        RECT 799.950 817.950 805.050 819.000 ;
        RECT 805.950 818.400 868.050 819.450 ;
        RECT 805.950 817.950 808.050 818.400 ;
        RECT 865.950 817.950 868.050 818.400 ;
        RECT 892.950 819.450 895.050 820.050 ;
        RECT 898.950 819.450 901.050 820.050 ;
        RECT 892.950 818.400 901.050 819.450 ;
        RECT 892.950 817.950 895.050 818.400 ;
        RECT 898.950 817.950 901.050 818.400 ;
        RECT 295.950 815.400 355.050 816.450 ;
        RECT 295.950 814.950 298.050 815.400 ;
        RECT 319.950 814.950 322.050 815.400 ;
        RECT 352.950 815.100 355.050 815.400 ;
        RECT 410.400 815.400 417.450 816.450 ;
        RECT 418.950 816.450 421.050 817.050 ;
        RECT 463.800 816.450 465.900 817.050 ;
        RECT 418.950 815.400 465.900 816.450 ;
        RECT 466.950 816.000 469.200 817.050 ;
        RECT 19.950 813.450 22.050 814.050 ;
        RECT 61.950 813.450 64.050 814.050 ;
        RECT 19.950 812.400 64.050 813.450 ;
        RECT 19.950 811.950 22.050 812.400 ;
        RECT 61.950 811.950 64.050 812.400 ;
        RECT 70.950 813.450 73.050 814.050 ;
        RECT 82.950 813.450 85.050 814.050 ;
        RECT 100.950 813.450 103.050 814.050 ;
        RECT 70.950 812.400 85.050 813.450 ;
        RECT 70.950 811.950 73.050 812.400 ;
        RECT 82.950 811.950 85.050 812.400 ;
        RECT 86.400 812.400 103.050 813.450 ;
        RECT 86.400 808.050 87.450 812.400 ;
        RECT 100.950 811.950 103.050 812.400 ;
        RECT 118.950 813.450 121.050 813.900 ;
        RECT 157.950 813.450 160.050 814.050 ;
        RECT 118.950 812.400 160.050 813.450 ;
        RECT 118.950 811.800 121.050 812.400 ;
        RECT 157.950 811.950 160.050 812.400 ;
        RECT 178.950 813.450 181.050 814.050 ;
        RECT 226.950 813.450 229.050 814.050 ;
        RECT 178.950 812.400 229.050 813.450 ;
        RECT 178.950 811.950 181.050 812.400 ;
        RECT 226.950 811.950 229.050 812.400 ;
        RECT 352.950 813.450 355.050 813.900 ;
        RECT 358.950 813.450 361.050 814.050 ;
        RECT 352.950 812.400 361.050 813.450 ;
        RECT 352.950 811.800 355.050 812.400 ;
        RECT 358.950 811.950 361.050 812.400 ;
        RECT 370.950 813.450 373.050 814.050 ;
        RECT 410.400 813.450 411.450 815.400 ;
        RECT 418.950 814.950 421.050 815.400 ;
        RECT 463.800 814.950 465.900 815.400 ;
        RECT 467.100 814.950 469.200 816.000 ;
        RECT 472.950 816.450 475.050 817.050 ;
        RECT 511.950 816.450 514.050 817.050 ;
        RECT 472.950 815.400 514.050 816.450 ;
        RECT 472.950 814.950 475.050 815.400 ;
        RECT 511.950 814.950 514.050 815.400 ;
        RECT 517.950 816.450 520.050 817.050 ;
        RECT 532.950 816.450 535.050 817.050 ;
        RECT 517.950 815.400 535.050 816.450 ;
        RECT 517.950 814.950 520.050 815.400 ;
        RECT 532.950 814.950 535.050 815.400 ;
        RECT 550.950 816.450 553.050 817.050 ;
        RECT 571.950 816.450 574.050 817.050 ;
        RECT 577.950 816.450 580.050 816.900 ;
        RECT 550.950 815.400 580.050 816.450 ;
        RECT 550.950 814.950 553.050 815.400 ;
        RECT 571.950 814.950 574.050 815.400 ;
        RECT 577.950 814.800 580.050 815.400 ;
        RECT 610.950 816.450 613.050 817.050 ;
        RECT 622.950 816.450 625.050 817.050 ;
        RECT 655.950 816.450 658.050 817.050 ;
        RECT 670.950 816.450 673.050 817.050 ;
        RECT 610.950 815.400 673.050 816.450 ;
        RECT 610.950 814.950 613.050 815.400 ;
        RECT 622.950 814.950 625.050 815.400 ;
        RECT 655.950 814.950 658.050 815.400 ;
        RECT 670.950 814.950 673.050 815.400 ;
        RECT 703.950 816.450 706.050 817.050 ;
        RECT 709.950 816.450 712.050 817.050 ;
        RECT 703.950 815.400 712.050 816.450 ;
        RECT 703.950 814.950 706.050 815.400 ;
        RECT 709.950 814.950 712.050 815.400 ;
        RECT 718.950 816.450 721.050 817.050 ;
        RECT 742.950 816.450 745.050 817.050 ;
        RECT 718.950 815.400 745.050 816.450 ;
        RECT 779.400 816.450 780.450 817.950 ;
        RECT 796.950 816.450 799.050 817.050 ;
        RECT 779.400 815.400 799.050 816.450 ;
        RECT 718.950 814.950 721.050 815.400 ;
        RECT 742.950 814.950 745.050 815.400 ;
        RECT 796.950 814.950 799.050 815.400 ;
        RECT 802.950 816.450 805.050 817.950 ;
        RECT 826.950 816.450 829.050 817.050 ;
        RECT 856.800 816.450 858.900 817.050 ;
        RECT 802.950 815.400 858.900 816.450 ;
        RECT 802.950 814.950 805.050 815.400 ;
        RECT 826.950 814.950 829.050 815.400 ;
        RECT 856.800 814.950 858.900 815.400 ;
        RECT 860.100 816.450 862.200 817.050 ;
        RECT 874.950 816.450 877.050 817.050 ;
        RECT 860.100 815.400 877.050 816.450 ;
        RECT 860.100 814.950 862.200 815.400 ;
        RECT 874.950 814.950 877.050 815.400 ;
        RECT 889.950 816.450 892.050 817.050 ;
        RECT 901.950 816.450 904.050 817.050 ;
        RECT 889.950 815.400 904.050 816.450 ;
        RECT 889.950 814.950 892.050 815.400 ;
        RECT 901.950 814.950 904.050 815.400 ;
        RECT 370.950 812.400 411.450 813.450 ;
        RECT 412.950 813.450 415.050 814.050 ;
        RECT 439.950 813.450 442.050 814.050 ;
        RECT 475.950 813.450 478.050 814.050 ;
        RECT 493.950 813.450 496.050 814.200 ;
        RECT 541.950 813.450 544.050 814.050 ;
        RECT 412.950 812.400 435.450 813.450 ;
        RECT 370.950 811.950 373.050 812.400 ;
        RECT 205.950 810.450 208.050 811.050 ;
        RECT 211.950 810.450 214.050 811.050 ;
        RECT 205.950 809.400 214.050 810.450 ;
        RECT 205.950 808.950 208.050 809.400 ;
        RECT 211.950 808.950 214.050 809.400 ;
        RECT 367.950 810.450 370.050 811.050 ;
        RECT 373.950 810.450 376.050 811.050 ;
        RECT 367.950 809.400 376.050 810.450 ;
        RECT 367.950 808.950 370.050 809.400 ;
        RECT 373.950 808.950 376.050 809.400 ;
        RECT 401.400 808.050 402.450 812.400 ;
        RECT 412.950 811.950 415.050 812.400 ;
        RECT 434.400 808.050 435.450 812.400 ;
        RECT 439.950 812.400 474.450 813.450 ;
        RECT 439.950 811.950 442.050 812.400 ;
        RECT 13.950 805.950 16.050 808.050 ;
        RECT 19.950 805.950 22.050 808.050 ;
        RECT 34.950 807.450 39.000 808.050 ;
        RECT 40.950 807.450 43.050 808.050 ;
        RECT 34.950 806.400 43.050 807.450 ;
        RECT 34.950 805.950 39.000 806.400 ;
        RECT 40.950 805.950 43.050 806.400 ;
        RECT 46.950 807.450 49.050 808.050 ;
        RECT 55.950 807.450 58.050 808.050 ;
        RECT 46.950 806.400 58.050 807.450 ;
        RECT 46.950 805.950 49.050 806.400 ;
        RECT 55.950 805.950 58.050 806.400 ;
        RECT 64.950 805.950 67.050 808.050 ;
        RECT 70.950 805.950 73.050 808.050 ;
        RECT 85.950 805.950 88.050 808.050 ;
        RECT 91.950 805.950 94.050 808.050 ;
        RECT 106.950 805.950 112.050 808.050 ;
        RECT 115.950 805.950 118.050 808.050 ;
        RECT 136.950 807.450 139.050 808.050 ;
        RECT 148.950 807.450 151.050 808.050 ;
        RECT 136.950 806.400 151.050 807.450 ;
        RECT 136.950 805.950 139.050 806.400 ;
        RECT 148.950 805.950 151.050 806.400 ;
        RECT 154.950 805.950 160.050 808.050 ;
        RECT 166.950 807.450 169.050 808.050 ;
        RECT 175.950 807.450 178.050 808.050 ;
        RECT 166.950 806.400 178.050 807.450 ;
        RECT 166.950 805.950 169.050 806.400 ;
        RECT 175.950 805.950 178.050 806.400 ;
        RECT 181.950 805.950 184.050 808.050 ;
        RECT 196.950 807.450 202.050 808.050 ;
        RECT 191.400 807.000 202.050 807.450 ;
        RECT 190.950 806.400 202.050 807.000 ;
        RECT 13.950 802.950 16.050 804.750 ;
        RECT 19.950 802.950 22.050 804.750 ;
        RECT 40.950 802.950 43.050 804.750 ;
        RECT 46.950 802.950 49.050 804.750 ;
        RECT 64.950 802.950 67.050 804.750 ;
        RECT 70.950 802.950 73.050 804.750 ;
        RECT 85.950 802.950 88.050 804.750 ;
        RECT 91.950 802.950 94.050 804.750 ;
        RECT 109.950 802.950 112.050 804.750 ;
        RECT 115.950 802.950 118.050 804.750 ;
        RECT 136.950 802.950 139.050 804.750 ;
        RECT 154.950 802.950 157.050 804.750 ;
        RECT 175.950 802.950 178.050 804.750 ;
        RECT 181.950 802.950 184.050 804.750 ;
        RECT 190.950 802.950 193.050 806.400 ;
        RECT 196.950 805.950 202.050 806.400 ;
        RECT 220.950 805.950 223.050 808.050 ;
        RECT 259.950 805.950 265.050 808.050 ;
        RECT 268.950 805.950 271.050 808.050 ;
        RECT 277.950 807.450 280.050 808.050 ;
        RECT 289.950 807.450 292.050 808.050 ;
        RECT 277.950 806.400 292.050 807.450 ;
        RECT 277.950 805.950 280.050 806.400 ;
        RECT 289.950 805.950 292.050 806.400 ;
        RECT 295.950 805.950 298.050 808.050 ;
        RECT 313.950 805.950 316.050 808.050 ;
        RECT 319.950 805.950 322.050 808.050 ;
        RECT 325.950 807.450 328.050 808.050 ;
        RECT 334.950 807.450 337.050 808.050 ;
        RECT 325.950 806.400 337.050 807.450 ;
        RECT 325.950 805.950 328.050 806.400 ;
        RECT 334.950 805.950 337.050 806.400 ;
        RECT 340.950 805.950 343.050 808.050 ;
        RECT 358.950 805.950 361.050 808.050 ;
        RECT 364.950 805.950 367.050 808.050 ;
        RECT 385.950 805.950 388.050 808.050 ;
        RECT 400.950 805.950 403.050 808.050 ;
        RECT 406.950 807.450 409.050 808.050 ;
        RECT 411.000 807.450 415.050 808.050 ;
        RECT 406.950 806.400 415.050 807.450 ;
        RECT 406.950 805.950 409.050 806.400 ;
        RECT 411.000 805.950 415.050 806.400 ;
        RECT 427.950 805.950 430.050 808.050 ;
        RECT 433.950 805.950 436.050 808.050 ;
        RECT 451.950 805.950 454.050 811.050 ;
        RECT 473.400 808.050 474.450 812.400 ;
        RECT 475.950 812.400 496.050 813.450 ;
        RECT 475.950 811.950 478.050 812.400 ;
        RECT 493.950 812.100 496.050 812.400 ;
        RECT 527.400 812.400 544.050 813.450 ;
        RECT 481.950 810.450 484.050 811.050 ;
        RECT 493.950 810.450 496.050 810.900 ;
        RECT 481.950 809.400 496.050 810.450 ;
        RECT 481.950 808.950 484.050 809.400 ;
        RECT 493.950 808.800 496.050 809.400 ;
        RECT 499.950 808.950 502.050 811.050 ;
        RECT 505.950 810.450 508.050 811.050 ;
        RECT 514.950 810.450 517.050 811.050 ;
        RECT 505.950 809.400 517.050 810.450 ;
        RECT 505.950 808.950 508.050 809.400 ;
        RECT 514.950 808.950 517.050 809.400 ;
        RECT 527.400 808.050 528.450 812.400 ;
        RECT 541.950 811.950 544.050 812.400 ;
        RECT 565.950 813.450 568.050 814.050 ;
        RECT 586.950 813.450 589.050 814.050 ;
        RECT 565.950 812.400 589.050 813.450 ;
        RECT 565.950 811.950 568.050 812.400 ;
        RECT 586.950 811.950 589.050 812.400 ;
        RECT 601.950 813.450 604.050 814.050 ;
        RECT 610.800 813.450 612.900 814.050 ;
        RECT 601.950 812.400 612.900 813.450 ;
        RECT 601.950 811.950 604.050 812.400 ;
        RECT 610.800 811.950 612.900 812.400 ;
        RECT 614.100 813.450 616.200 814.050 ;
        RECT 625.950 813.450 628.050 814.050 ;
        RECT 614.100 812.400 628.050 813.450 ;
        RECT 614.100 811.950 616.200 812.400 ;
        RECT 625.950 811.950 628.050 812.400 ;
        RECT 646.950 813.450 649.050 814.050 ;
        RECT 658.950 813.450 661.050 814.050 ;
        RECT 691.950 813.450 694.050 814.050 ;
        RECT 646.950 812.400 694.050 813.450 ;
        RECT 646.950 811.950 649.050 812.400 ;
        RECT 658.950 811.950 661.050 812.400 ;
        RECT 691.950 811.950 694.050 812.400 ;
        RECT 697.950 813.450 700.050 814.050 ;
        RECT 724.950 813.450 727.050 814.050 ;
        RECT 697.950 812.400 727.050 813.450 ;
        RECT 697.950 811.950 700.050 812.400 ;
        RECT 724.950 811.950 727.050 812.400 ;
        RECT 748.950 813.450 751.050 814.050 ;
        RECT 757.950 813.450 760.050 814.050 ;
        RECT 823.950 813.450 826.050 814.050 ;
        RECT 838.950 813.450 841.050 814.050 ;
        RECT 748.950 812.400 841.050 813.450 ;
        RECT 748.950 811.950 751.050 812.400 ;
        RECT 757.950 811.950 760.050 812.400 ;
        RECT 823.950 811.950 826.050 812.400 ;
        RECT 838.950 811.950 841.050 812.400 ;
        RECT 886.950 813.450 889.050 814.050 ;
        RECT 898.950 813.450 901.050 814.050 ;
        RECT 886.950 812.400 901.050 813.450 ;
        RECT 886.950 811.950 889.050 812.400 ;
        RECT 898.950 811.950 901.050 812.400 ;
        RECT 550.950 808.950 553.050 811.050 ;
        RECT 556.950 808.950 559.050 811.050 ;
        RECT 628.950 810.450 631.050 811.050 ;
        RECT 634.950 810.450 637.050 811.050 ;
        RECT 628.950 809.400 637.050 810.450 ;
        RECT 628.950 808.950 631.050 809.400 ;
        RECT 634.950 808.950 637.050 809.400 ;
        RECT 676.950 810.450 679.050 811.050 ;
        RECT 682.950 810.450 685.050 811.050 ;
        RECT 676.950 809.400 685.050 810.450 ;
        RECT 676.950 808.950 679.050 809.400 ;
        RECT 682.950 808.950 685.050 809.400 ;
        RECT 700.950 808.950 706.050 811.050 ;
        RECT 865.950 808.950 868.050 811.050 ;
        RECT 871.950 808.950 874.050 811.050 ;
        RECT 457.950 805.950 460.050 808.050 ;
        RECT 472.950 805.950 475.050 808.050 ;
        RECT 478.950 805.950 481.050 808.050 ;
        RECT 499.950 805.950 502.050 807.750 ;
        RECT 505.950 805.950 508.050 807.750 ;
        RECT 526.950 805.950 529.050 808.050 ;
        RECT 532.950 805.950 535.050 808.050 ;
        RECT 550.950 805.950 553.050 807.750 ;
        RECT 556.950 805.950 559.050 807.750 ;
        RECT 577.950 805.950 580.050 808.050 ;
        RECT 601.950 807.450 604.050 808.050 ;
        RECT 610.950 807.450 613.050 808.050 ;
        RECT 601.950 806.400 613.050 807.450 ;
        RECT 601.950 805.950 604.050 806.400 ;
        RECT 610.950 805.950 613.050 806.400 ;
        RECT 616.950 805.950 622.050 808.050 ;
        RECT 625.950 805.950 628.050 808.050 ;
        RECT 640.950 805.950 646.050 808.050 ;
        RECT 649.950 805.950 652.050 808.050 ;
        RECT 670.950 805.950 673.050 808.050 ;
        RECT 688.950 805.950 691.050 808.050 ;
        RECT 694.950 807.450 697.050 808.050 ;
        RECT 709.950 807.450 712.050 808.050 ;
        RECT 694.950 806.400 712.050 807.450 ;
        RECT 694.950 805.950 697.050 806.400 ;
        RECT 709.950 805.950 712.050 806.400 ;
        RECT 715.950 805.950 718.050 808.050 ;
        RECT 733.950 807.450 736.050 808.050 ;
        RECT 748.950 807.450 751.050 808.050 ;
        RECT 733.950 806.400 751.050 807.450 ;
        RECT 733.950 805.950 736.050 806.400 ;
        RECT 748.950 805.950 751.050 806.400 ;
        RECT 754.950 805.950 757.050 808.050 ;
        RECT 760.950 805.950 763.050 808.050 ;
        RECT 766.950 807.450 769.050 808.050 ;
        RECT 775.950 807.450 778.050 808.050 ;
        RECT 781.950 807.450 784.050 808.050 ;
        RECT 766.950 806.400 784.050 807.450 ;
        RECT 766.950 805.950 769.050 806.400 ;
        RECT 775.950 805.950 778.050 806.400 ;
        RECT 781.950 805.950 784.050 806.400 ;
        RECT 802.950 805.950 805.050 808.050 ;
        RECT 814.950 805.950 817.050 808.050 ;
        RECT 820.950 805.950 823.050 808.050 ;
        RECT 838.950 805.950 841.050 808.050 ;
        RECT 844.950 807.450 847.050 808.050 ;
        RECT 859.950 807.450 862.050 808.050 ;
        RECT 844.950 806.400 862.050 807.450 ;
        RECT 844.950 805.950 847.050 806.400 ;
        RECT 859.950 805.950 862.050 806.400 ;
        RECT 865.950 805.950 868.050 807.750 ;
        RECT 871.950 805.950 874.050 807.750 ;
        RECT 886.950 805.950 889.050 808.050 ;
        RECT 892.950 807.450 895.050 808.050 ;
        RECT 897.000 807.450 901.050 808.050 ;
        RECT 892.950 806.400 901.050 807.450 ;
        RECT 892.950 805.950 895.050 806.400 ;
        RECT 897.000 805.950 901.050 806.400 ;
        RECT 217.950 804.750 219.750 805.050 ;
        RECT 199.950 802.950 202.050 804.750 ;
        RECT 217.950 803.250 220.050 804.750 ;
        RECT 220.950 803.250 223.050 804.750 ;
        RECT 226.950 803.250 229.050 805.050 ;
        RECT 241.950 803.250 244.050 805.050 ;
        RECT 221.250 802.950 223.050 803.250 ;
        RECT 247.950 802.950 250.050 804.750 ;
        RECT 262.950 802.950 265.050 804.750 ;
        RECT 268.950 802.950 271.050 804.750 ;
        RECT 289.950 802.950 292.050 804.750 ;
        RECT 295.950 802.950 298.050 804.750 ;
        RECT 313.950 802.950 316.050 804.750 ;
        RECT 319.950 802.950 322.050 804.750 ;
        RECT 334.950 802.950 337.050 804.750 ;
        RECT 340.950 802.950 343.050 804.750 ;
        RECT 358.950 802.950 361.050 804.750 ;
        RECT 364.950 802.950 367.050 804.750 ;
        RECT 385.950 802.950 388.050 804.750 ;
        RECT 400.950 802.950 403.050 804.750 ;
        RECT 406.950 802.950 409.050 804.750 ;
        RECT 427.950 802.950 430.050 804.750 ;
        RECT 433.950 802.950 436.050 804.750 ;
        RECT 451.950 802.950 454.050 804.750 ;
        RECT 457.950 802.950 460.050 804.750 ;
        RECT 472.950 802.950 475.050 804.750 ;
        RECT 478.950 802.950 481.050 804.750 ;
        RECT 496.950 803.250 499.050 805.050 ;
        RECT 502.950 803.250 505.050 805.050 ;
        RECT 508.950 803.250 511.050 805.050 ;
        RECT 526.950 802.950 529.050 804.750 ;
        RECT 532.950 802.950 535.050 804.750 ;
        RECT 547.950 803.250 550.050 805.050 ;
        RECT 553.950 803.250 556.050 805.050 ;
        RECT 559.950 803.250 562.050 805.050 ;
        RECT 571.950 803.250 574.050 805.050 ;
        RECT 581.250 804.750 583.050 805.050 ;
        RECT 577.950 803.250 580.050 804.750 ;
        RECT 580.950 803.250 583.050 804.750 ;
        RECT 577.950 802.950 579.750 803.250 ;
        RECT 601.950 802.950 604.050 804.750 ;
        RECT 619.950 802.950 622.050 804.750 ;
        RECT 625.950 802.950 628.050 804.750 ;
        RECT 643.950 802.950 646.050 804.750 ;
        RECT 649.950 802.950 652.050 804.750 ;
        RECT 670.950 802.950 673.050 804.750 ;
        RECT 682.950 803.250 685.050 805.050 ;
        RECT 692.250 804.750 694.050 805.050 ;
        RECT 688.950 803.250 691.050 804.750 ;
        RECT 691.950 803.250 694.050 804.750 ;
        RECT 688.950 802.950 690.750 803.250 ;
        RECT 709.950 802.950 712.050 804.750 ;
        RECT 715.950 802.950 718.050 804.750 ;
        RECT 733.950 802.950 736.050 804.750 ;
        RECT 754.950 802.950 757.050 804.750 ;
        RECT 760.950 802.950 763.050 804.750 ;
        RECT 781.950 802.950 784.050 804.750 ;
        RECT 802.950 802.950 805.050 804.750 ;
        RECT 814.950 802.950 817.050 804.750 ;
        RECT 820.950 802.950 823.050 804.750 ;
        RECT 838.950 802.950 841.050 804.750 ;
        RECT 844.950 802.950 847.050 804.750 ;
        RECT 868.950 803.250 871.050 805.050 ;
        RECT 886.950 802.950 889.050 804.750 ;
        RECT 892.950 802.950 895.050 804.750 ;
        RECT 634.950 802.050 637.050 802.200 ;
        RECT 16.950 800.250 19.050 802.050 ;
        RECT 22.950 800.250 25.050 802.050 ;
        RECT 37.950 800.250 40.050 802.050 ;
        RECT 43.950 800.250 46.050 802.050 ;
        RECT 61.950 800.250 64.050 802.050 ;
        RECT 67.950 800.250 70.050 802.050 ;
        RECT 88.950 800.250 91.050 802.050 ;
        RECT 94.950 800.250 97.050 802.050 ;
        RECT 112.950 800.250 115.050 802.050 ;
        RECT 118.950 800.250 121.050 802.050 ;
        RECT 133.950 800.250 136.050 802.050 ;
        RECT 151.950 800.250 154.050 802.050 ;
        RECT 157.950 800.250 160.050 802.050 ;
        RECT 172.950 800.250 175.050 802.050 ;
        RECT 178.950 800.250 181.050 802.050 ;
        RECT 196.950 800.250 199.050 802.050 ;
        RECT 202.950 800.250 205.050 802.050 ;
        RECT 16.950 796.950 19.050 799.050 ;
        RECT 22.950 796.950 25.050 799.050 ;
        RECT 37.950 796.950 40.050 799.050 ;
        RECT 43.950 796.950 46.050 799.050 ;
        RECT 61.950 796.950 64.050 799.050 ;
        RECT 67.950 796.950 70.050 799.050 ;
        RECT 88.950 796.950 91.050 799.050 ;
        RECT 94.950 796.950 97.050 799.050 ;
        RECT 100.950 798.450 103.050 799.050 ;
        RECT 112.950 798.450 115.050 799.050 ;
        RECT 100.950 797.400 115.050 798.450 ;
        RECT 100.950 796.950 103.050 797.400 ;
        RECT 112.950 796.950 115.050 797.400 ;
        RECT 118.950 796.950 121.050 799.050 ;
        RECT 124.950 798.450 127.050 799.050 ;
        RECT 133.950 798.450 136.050 799.050 ;
        RECT 124.950 797.400 136.050 798.450 ;
        RECT 124.950 796.950 127.050 797.400 ;
        RECT 133.950 796.950 136.050 797.400 ;
        RECT 151.950 796.950 154.050 799.050 ;
        RECT 157.950 796.950 160.050 799.050 ;
        RECT 163.950 798.450 166.050 799.050 ;
        RECT 172.950 798.450 175.050 799.050 ;
        RECT 163.950 797.400 175.050 798.450 ;
        RECT 163.950 796.950 166.050 797.400 ;
        RECT 172.950 796.950 175.050 797.400 ;
        RECT 178.950 796.950 181.050 799.050 ;
        RECT 196.950 796.950 199.050 799.050 ;
        RECT 202.950 796.950 205.050 799.050 ;
        RECT 217.950 796.950 220.050 802.050 ;
        RECT 226.950 799.950 229.050 802.050 ;
        RECT 241.950 799.950 244.050 802.050 ;
        RECT 265.950 800.250 268.050 802.050 ;
        RECT 271.950 800.250 274.050 802.050 ;
        RECT 286.950 800.250 289.050 802.050 ;
        RECT 292.950 800.250 295.050 802.050 ;
        RECT 310.950 800.250 313.050 802.050 ;
        RECT 316.950 800.250 319.050 802.050 ;
        RECT 337.950 800.250 340.050 802.050 ;
        RECT 343.950 800.250 346.050 802.050 ;
        RECT 361.950 800.250 364.050 802.050 ;
        RECT 367.950 800.250 370.050 802.050 ;
        RECT 382.950 800.250 385.050 802.050 ;
        RECT 397.950 800.250 400.050 802.050 ;
        RECT 403.950 800.250 406.050 802.050 ;
        RECT 424.950 800.250 427.050 802.050 ;
        RECT 430.950 800.250 433.050 802.050 ;
        RECT 448.950 800.250 451.050 802.050 ;
        RECT 454.950 800.250 457.050 802.050 ;
        RECT 475.950 800.250 478.050 802.050 ;
        RECT 481.950 800.250 484.050 802.050 ;
        RECT 493.950 799.950 499.050 802.050 ;
        RECT 208.950 795.450 211.050 796.050 ;
        RECT 242.400 795.450 243.450 799.950 ;
        RECT 262.950 796.950 268.050 799.050 ;
        RECT 271.950 796.950 274.050 799.050 ;
        RECT 286.950 796.950 289.050 799.050 ;
        RECT 292.950 796.950 295.050 799.050 ;
        RECT 310.950 796.950 313.050 799.050 ;
        RECT 316.950 796.950 319.050 799.050 ;
        RECT 337.950 796.950 340.050 799.050 ;
        RECT 343.950 796.950 346.050 799.050 ;
        RECT 361.950 796.950 364.050 799.050 ;
        RECT 367.950 796.950 370.050 799.050 ;
        RECT 373.950 798.450 376.050 799.050 ;
        RECT 382.950 798.450 385.050 799.050 ;
        RECT 373.950 797.400 385.050 798.450 ;
        RECT 373.950 796.950 376.050 797.400 ;
        RECT 382.950 796.950 385.050 797.400 ;
        RECT 388.950 798.450 391.050 799.050 ;
        RECT 397.950 798.450 400.050 799.050 ;
        RECT 388.950 797.400 400.050 798.450 ;
        RECT 388.950 796.950 391.050 797.400 ;
        RECT 397.950 796.950 400.050 797.400 ;
        RECT 403.950 796.950 406.050 799.050 ;
        RECT 409.950 798.450 412.050 799.050 ;
        RECT 424.950 798.450 427.050 799.050 ;
        RECT 409.950 797.400 427.050 798.450 ;
        RECT 409.950 796.950 412.050 797.400 ;
        RECT 424.950 796.950 427.050 797.400 ;
        RECT 430.950 796.950 433.050 799.050 ;
        RECT 436.950 798.450 439.050 799.050 ;
        RECT 442.950 798.450 445.050 799.050 ;
        RECT 436.950 797.400 445.050 798.450 ;
        RECT 436.950 796.950 439.050 797.400 ;
        RECT 442.950 796.950 445.050 797.400 ;
        RECT 448.950 796.950 451.050 799.050 ;
        RECT 454.950 796.950 457.050 799.050 ;
        RECT 208.950 794.400 243.450 795.450 ;
        RECT 208.950 793.950 211.050 794.400 ;
        RECT 415.950 793.950 421.050 796.050 ;
        RECT 466.950 793.950 469.050 799.050 ;
        RECT 475.950 796.950 478.050 799.050 ;
        RECT 481.950 796.950 484.050 799.050 ;
        RECT 502.950 796.950 505.050 802.050 ;
        RECT 508.950 799.950 511.050 802.050 ;
        RECT 523.950 800.250 526.050 802.050 ;
        RECT 529.950 800.250 532.050 802.050 ;
        RECT 535.950 801.450 538.050 802.050 ;
        RECT 547.950 801.450 550.050 802.050 ;
        RECT 535.950 800.400 550.050 801.450 ;
        RECT 535.950 799.950 538.050 800.400 ;
        RECT 547.950 799.950 550.050 800.400 ;
        RECT 553.950 799.950 556.050 802.050 ;
        RECT 559.950 799.950 562.050 802.050 ;
        RECT 523.950 796.950 526.050 799.050 ;
        RECT 529.950 796.950 532.050 799.050 ;
        RECT 496.950 795.450 499.050 796.200 ;
        RECT 517.950 795.450 520.050 796.050 ;
        RECT 496.950 794.400 520.050 795.450 ;
        RECT 496.950 794.100 499.050 794.400 ;
        RECT 517.950 793.950 520.050 794.400 ;
        RECT 532.950 795.450 535.050 796.050 ;
        RECT 554.400 795.450 555.450 799.950 ;
        RECT 571.950 796.950 574.050 802.050 ;
        RECT 580.950 801.450 583.050 802.050 ;
        RECT 592.950 801.450 595.050 802.050 ;
        RECT 580.950 800.400 595.050 801.450 ;
        RECT 580.950 799.950 583.050 800.400 ;
        RECT 592.950 799.950 595.050 800.400 ;
        RECT 598.950 800.250 601.050 802.050 ;
        RECT 604.950 800.250 607.050 802.050 ;
        RECT 622.950 800.250 625.050 802.050 ;
        RECT 628.950 800.250 631.050 802.050 ;
        RECT 634.950 800.100 640.050 802.050 ;
        RECT 646.950 800.250 649.050 802.050 ;
        RECT 652.950 800.250 655.050 802.050 ;
        RECT 667.950 800.250 670.050 802.050 ;
        RECT 636.000 799.950 640.050 800.100 ;
        RECT 682.950 799.950 685.050 802.050 ;
        RECT 691.950 801.450 694.050 802.050 ;
        RECT 696.000 801.450 700.050 802.050 ;
        RECT 691.950 800.400 700.050 801.450 ;
        RECT 691.950 799.950 694.050 800.400 ;
        RECT 696.000 799.950 700.050 800.400 ;
        RECT 712.950 800.250 715.050 802.050 ;
        RECT 718.950 800.250 721.050 802.050 ;
        RECT 730.950 800.250 733.050 802.050 ;
        RECT 736.950 800.250 739.050 802.050 ;
        RECT 757.950 800.250 760.050 802.050 ;
        RECT 763.950 800.250 766.050 802.050 ;
        RECT 778.950 800.250 781.050 802.050 ;
        RECT 784.950 800.250 787.050 802.050 ;
        RECT 793.800 801.000 795.900 802.050 ;
        RECT 793.800 799.950 796.050 801.000 ;
        RECT 799.950 800.250 802.050 802.050 ;
        RECT 817.950 800.250 820.050 802.050 ;
        RECT 823.950 800.250 826.050 802.050 ;
        RECT 841.950 800.250 844.050 802.050 ;
        RECT 847.950 800.250 850.050 802.050 ;
        RECT 598.950 796.950 601.050 799.050 ;
        RECT 604.950 796.950 607.050 799.050 ;
        RECT 622.950 796.950 625.050 799.050 ;
        RECT 628.950 796.950 631.050 799.050 ;
        RECT 634.950 798.450 637.050 798.900 ;
        RECT 646.950 798.450 649.050 799.050 ;
        RECT 634.950 797.400 649.050 798.450 ;
        RECT 634.950 796.800 637.050 797.400 ;
        RECT 646.950 796.950 649.050 797.400 ;
        RECT 652.950 796.950 655.050 799.050 ;
        RECT 658.950 798.450 661.050 799.050 ;
        RECT 667.950 798.450 670.050 799.050 ;
        RECT 658.950 797.400 670.050 798.450 ;
        RECT 658.950 796.950 661.050 797.400 ;
        RECT 667.950 796.950 670.050 797.400 ;
        RECT 700.950 798.450 703.050 799.050 ;
        RECT 706.950 798.450 709.050 799.200 ;
        RECT 793.950 799.050 796.050 799.950 ;
        RECT 700.950 797.400 709.050 798.450 ;
        RECT 700.950 796.950 703.050 797.400 ;
        RECT 706.950 797.100 709.050 797.400 ;
        RECT 712.950 796.950 715.050 799.050 ;
        RECT 718.950 796.950 721.050 799.050 ;
        RECT 730.950 796.950 733.050 799.050 ;
        RECT 736.950 796.950 739.050 799.050 ;
        RECT 757.950 796.950 760.050 799.050 ;
        RECT 763.950 796.950 766.050 799.050 ;
        RECT 778.950 796.950 781.050 799.050 ;
        RECT 784.950 796.950 787.050 799.050 ;
        RECT 793.800 798.000 796.050 799.050 ;
        RECT 797.100 798.450 802.050 799.050 ;
        RECT 808.950 798.450 811.050 799.050 ;
        RECT 793.800 796.950 795.900 798.000 ;
        RECT 797.100 797.400 811.050 798.450 ;
        RECT 797.100 796.950 802.050 797.400 ;
        RECT 808.950 796.950 811.050 797.400 ;
        RECT 817.950 796.950 820.050 799.050 ;
        RECT 823.950 796.950 826.050 799.050 ;
        RECT 841.950 796.950 844.050 799.050 ;
        RECT 847.950 796.950 850.050 799.050 ;
        RECT 868.950 796.950 871.050 802.050 ;
        RECT 883.950 800.250 886.050 802.050 ;
        RECT 889.950 800.250 892.050 802.050 ;
        RECT 895.950 801.450 898.050 802.050 ;
        RECT 904.950 801.450 907.050 802.050 ;
        RECT 895.950 800.400 907.050 801.450 ;
        RECT 895.950 799.950 898.050 800.400 ;
        RECT 904.950 799.950 907.050 800.400 ;
        RECT 883.950 796.950 886.050 799.050 ;
        RECT 889.950 796.950 892.050 799.050 ;
        RECT 532.950 794.400 555.450 795.450 ;
        RECT 637.950 795.450 642.000 796.050 ;
        RECT 694.950 795.450 697.050 796.050 ;
        RECT 706.950 795.450 709.050 795.900 ;
        RECT 532.950 793.950 535.050 794.400 ;
        RECT 637.950 793.950 642.450 795.450 ;
        RECT 694.950 794.400 709.050 795.450 ;
        RECT 694.950 793.950 697.050 794.400 ;
        RECT 16.950 792.450 19.050 793.050 ;
        RECT 22.950 792.450 25.050 793.050 ;
        RECT 16.950 791.400 25.050 792.450 ;
        RECT 16.950 790.950 19.050 791.400 ;
        RECT 22.950 790.950 25.050 791.400 ;
        RECT 55.950 792.450 58.050 793.050 ;
        RECT 67.950 792.450 70.050 793.050 ;
        RECT 55.950 791.400 70.050 792.450 ;
        RECT 55.950 790.950 58.050 791.400 ;
        RECT 67.950 790.950 70.050 791.400 ;
        RECT 88.950 792.450 91.050 793.050 ;
        RECT 118.950 792.450 121.050 793.050 ;
        RECT 88.950 791.400 121.050 792.450 ;
        RECT 88.950 790.950 91.050 791.400 ;
        RECT 118.950 790.950 121.050 791.400 ;
        RECT 151.950 792.450 154.050 793.050 ;
        RECT 163.950 792.450 166.050 793.050 ;
        RECT 151.950 791.400 166.050 792.450 ;
        RECT 151.950 790.950 154.050 791.400 ;
        RECT 163.950 790.950 166.050 791.400 ;
        RECT 196.950 792.450 199.050 793.050 ;
        RECT 214.950 792.450 217.050 793.050 ;
        RECT 196.950 791.400 217.050 792.450 ;
        RECT 196.950 790.950 199.050 791.400 ;
        RECT 214.950 790.950 217.050 791.400 ;
        RECT 226.950 792.450 229.050 793.050 ;
        RECT 247.950 792.450 250.050 793.050 ;
        RECT 256.950 792.450 259.050 793.050 ;
        RECT 226.950 791.400 259.050 792.450 ;
        RECT 226.950 790.950 229.050 791.400 ;
        RECT 247.950 790.950 250.050 791.400 ;
        RECT 256.950 790.950 259.050 791.400 ;
        RECT 271.950 792.450 274.050 793.050 ;
        RECT 280.950 792.450 283.050 793.050 ;
        RECT 271.950 791.400 283.050 792.450 ;
        RECT 271.950 790.950 274.050 791.400 ;
        RECT 280.950 790.950 283.050 791.400 ;
        RECT 292.950 792.450 295.050 793.050 ;
        RECT 316.950 792.450 319.050 793.050 ;
        RECT 325.950 792.450 328.050 793.050 ;
        RECT 292.950 791.400 328.050 792.450 ;
        RECT 292.950 790.950 295.050 791.400 ;
        RECT 316.950 790.950 319.050 791.400 ;
        RECT 325.950 790.950 328.050 791.400 ;
        RECT 337.950 792.450 340.050 793.050 ;
        RECT 346.950 792.450 349.050 793.050 ;
        RECT 424.950 792.450 427.050 793.050 ;
        RECT 337.950 791.400 349.050 792.450 ;
        RECT 337.950 790.950 340.050 791.400 ;
        RECT 346.950 790.950 349.050 791.400 ;
        RECT 350.400 791.400 427.050 792.450 ;
        RECT 28.950 784.950 31.050 790.050 ;
        RECT 145.950 789.450 148.050 790.050 ;
        RECT 208.800 789.450 210.900 790.050 ;
        RECT 145.950 788.400 210.900 789.450 ;
        RECT 145.950 787.950 148.050 788.400 ;
        RECT 208.800 787.950 210.900 788.400 ;
        RECT 212.100 789.450 214.200 790.050 ;
        RECT 217.950 789.450 220.050 790.050 ;
        RECT 212.100 788.400 220.050 789.450 ;
        RECT 212.100 787.950 214.200 788.400 ;
        RECT 217.950 787.950 220.050 788.400 ;
        RECT 235.950 789.450 238.050 790.050 ;
        RECT 350.400 789.450 351.450 791.400 ;
        RECT 424.950 790.950 427.050 791.400 ;
        RECT 430.950 792.450 433.050 793.050 ;
        RECT 436.950 792.450 439.050 793.050 ;
        RECT 430.950 791.400 439.050 792.450 ;
        RECT 430.950 790.950 433.050 791.400 ;
        RECT 436.950 790.950 439.050 791.400 ;
        RECT 445.950 792.450 448.050 793.050 ;
        RECT 454.950 792.450 457.050 793.050 ;
        RECT 487.950 792.450 490.050 793.050 ;
        RECT 445.950 791.400 490.050 792.450 ;
        RECT 445.950 790.950 448.050 791.400 ;
        RECT 454.950 790.950 457.050 791.400 ;
        RECT 487.950 790.950 490.050 791.400 ;
        RECT 496.950 792.450 499.050 792.900 ;
        RECT 514.950 792.450 517.050 793.050 ;
        RECT 496.950 791.400 517.050 792.450 ;
        RECT 496.950 790.800 499.050 791.400 ;
        RECT 514.950 790.950 517.050 791.400 ;
        RECT 550.950 792.450 553.050 793.050 ;
        RECT 637.950 792.450 640.050 793.050 ;
        RECT 550.950 791.400 640.050 792.450 ;
        RECT 641.400 792.450 642.450 793.950 ;
        RECT 706.950 793.800 709.050 794.400 ;
        RECT 790.950 795.450 795.000 796.050 ;
        RECT 805.950 795.450 808.050 796.050 ;
        RECT 790.950 793.950 795.450 795.450 ;
        RECT 805.950 794.400 816.450 795.450 ;
        RECT 805.950 793.950 808.050 794.400 ;
        RECT 736.950 792.450 739.050 793.050 ;
        RECT 641.400 791.400 739.050 792.450 ;
        RECT 550.950 790.950 553.050 791.400 ;
        RECT 637.950 790.950 640.050 791.400 ;
        RECT 736.950 790.950 739.050 791.400 ;
        RECT 742.950 792.450 745.050 793.050 ;
        RECT 778.950 792.450 781.050 793.050 ;
        RECT 742.950 791.400 781.050 792.450 ;
        RECT 794.400 792.450 795.450 793.950 ;
        RECT 802.950 792.450 805.050 793.050 ;
        RECT 794.400 791.400 805.050 792.450 ;
        RECT 815.400 792.450 816.450 794.400 ;
        RECT 835.950 792.450 838.050 793.050 ;
        RECT 868.950 792.450 871.050 793.050 ;
        RECT 889.800 792.450 891.900 793.050 ;
        RECT 815.400 791.400 838.050 792.450 ;
        RECT 742.950 790.950 745.050 791.400 ;
        RECT 778.950 790.950 781.050 791.400 ;
        RECT 802.950 790.950 805.050 791.400 ;
        RECT 835.950 790.950 838.050 791.400 ;
        RECT 839.400 791.400 891.900 792.450 ;
        RECT 235.950 788.400 351.450 789.450 ;
        RECT 358.950 789.450 361.050 790.050 ;
        RECT 379.950 789.450 382.050 790.050 ;
        RECT 406.800 789.450 408.900 790.050 ;
        RECT 358.950 788.400 408.900 789.450 ;
        RECT 235.950 787.950 238.050 788.400 ;
        RECT 358.950 787.950 361.050 788.400 ;
        RECT 379.950 787.950 382.050 788.400 ;
        RECT 406.800 787.950 408.900 788.400 ;
        RECT 410.100 787.950 414.900 790.050 ;
        RECT 416.100 787.950 421.050 790.050 ;
        RECT 427.950 789.450 430.050 790.050 ;
        RECT 436.800 789.450 438.900 790.050 ;
        RECT 427.950 788.400 438.900 789.450 ;
        RECT 427.950 787.950 430.050 788.400 ;
        RECT 436.800 787.950 438.900 788.400 ;
        RECT 440.100 789.450 442.200 790.050 ;
        RECT 469.950 789.450 472.050 790.050 ;
        RECT 440.100 788.400 472.050 789.450 ;
        RECT 440.100 787.950 442.200 788.400 ;
        RECT 469.950 787.950 472.050 788.400 ;
        RECT 517.950 789.450 520.050 790.050 ;
        RECT 541.950 789.450 544.050 790.050 ;
        RECT 565.950 789.450 568.050 790.050 ;
        RECT 517.950 788.400 568.050 789.450 ;
        RECT 517.950 787.950 520.050 788.400 ;
        RECT 541.950 787.950 544.050 788.400 ;
        RECT 565.950 787.950 568.050 788.400 ;
        RECT 571.950 789.450 574.050 790.200 ;
        RECT 613.950 789.450 616.050 790.050 ;
        RECT 571.950 788.400 616.050 789.450 ;
        RECT 571.950 788.100 574.050 788.400 ;
        RECT 613.950 787.950 616.050 788.400 ;
        RECT 634.950 789.450 637.050 790.050 ;
        RECT 649.950 789.450 652.050 790.050 ;
        RECT 634.950 788.400 652.050 789.450 ;
        RECT 634.950 787.950 637.050 788.400 ;
        RECT 649.950 787.950 652.050 788.400 ;
        RECT 682.950 789.450 685.050 790.050 ;
        RECT 694.950 789.450 697.050 790.050 ;
        RECT 700.950 789.450 703.050 790.050 ;
        RECT 682.950 788.400 703.050 789.450 ;
        RECT 682.950 787.950 685.050 788.400 ;
        RECT 694.950 787.950 697.050 788.400 ;
        RECT 700.950 787.950 703.050 788.400 ;
        RECT 763.950 789.450 766.050 790.050 ;
        RECT 772.950 789.450 775.050 790.050 ;
        RECT 817.950 789.450 820.050 790.050 ;
        RECT 839.400 789.450 840.450 791.400 ;
        RECT 868.950 790.950 871.050 791.400 ;
        RECT 889.800 790.950 891.900 791.400 ;
        RECT 893.100 792.450 895.200 793.050 ;
        RECT 901.950 792.450 904.050 793.050 ;
        RECT 893.100 791.400 904.050 792.450 ;
        RECT 893.100 790.950 895.200 791.400 ;
        RECT 901.950 790.950 904.050 791.400 ;
        RECT 763.950 788.400 798.450 789.450 ;
        RECT 763.950 787.950 766.050 788.400 ;
        RECT 772.950 787.950 775.050 788.400 ;
        RECT 91.950 786.450 94.050 787.050 ;
        RECT 100.950 786.450 103.050 787.050 ;
        RECT 91.950 785.400 103.050 786.450 ;
        RECT 91.950 784.950 94.050 785.400 ;
        RECT 100.950 784.950 103.050 785.400 ;
        RECT 166.950 784.950 172.050 787.050 ;
        RECT 181.950 786.450 184.050 787.050 ;
        RECT 199.800 786.450 201.900 787.050 ;
        RECT 181.950 785.400 201.900 786.450 ;
        RECT 181.950 784.950 184.050 785.400 ;
        RECT 199.800 784.950 201.900 785.400 ;
        RECT 203.100 786.450 205.200 787.050 ;
        RECT 247.950 786.450 250.050 787.050 ;
        RECT 203.100 785.400 250.050 786.450 ;
        RECT 203.100 784.950 205.200 785.400 ;
        RECT 247.950 784.950 250.050 785.400 ;
        RECT 268.950 786.450 271.050 787.050 ;
        RECT 274.800 786.450 276.900 787.050 ;
        RECT 268.950 785.400 276.900 786.450 ;
        RECT 268.950 784.950 271.050 785.400 ;
        RECT 274.800 784.950 276.900 785.400 ;
        RECT 278.100 786.450 280.200 787.050 ;
        RECT 286.950 786.450 289.050 787.050 ;
        RECT 278.100 785.400 289.050 786.450 ;
        RECT 278.100 784.950 280.200 785.400 ;
        RECT 286.950 784.950 289.050 785.400 ;
        RECT 298.950 786.450 301.050 787.050 ;
        RECT 340.950 786.450 343.050 787.050 ;
        RECT 298.950 785.400 343.050 786.450 ;
        RECT 298.950 784.950 301.050 785.400 ;
        RECT 340.950 784.950 343.050 785.400 ;
        RECT 346.950 786.450 349.050 787.050 ;
        RECT 373.950 786.450 376.050 787.050 ;
        RECT 382.950 786.450 385.050 787.050 ;
        RECT 346.950 785.400 376.050 786.450 ;
        RECT 346.950 784.950 349.050 785.400 ;
        RECT 373.950 784.950 376.050 785.400 ;
        RECT 377.400 785.400 385.050 786.450 ;
        RECT 100.950 783.450 103.050 784.050 ;
        RECT 127.950 783.450 130.050 784.050 ;
        RECT 100.950 782.400 130.050 783.450 ;
        RECT 100.950 781.950 103.050 782.400 ;
        RECT 127.950 781.950 130.050 782.400 ;
        RECT 136.950 783.450 139.050 784.050 ;
        RECT 166.950 783.450 169.050 784.050 ;
        RECT 136.950 782.400 169.050 783.450 ;
        RECT 136.950 781.950 139.050 782.400 ;
        RECT 166.950 781.950 169.050 782.400 ;
        RECT 178.950 783.450 181.050 784.050 ;
        RECT 208.950 783.450 211.050 784.050 ;
        RECT 178.950 782.400 211.050 783.450 ;
        RECT 178.950 781.950 181.050 782.400 ;
        RECT 208.950 781.950 211.050 782.400 ;
        RECT 226.950 783.450 229.050 784.050 ;
        RECT 235.950 783.450 238.050 784.050 ;
        RECT 226.950 782.400 238.050 783.450 ;
        RECT 287.400 783.450 288.450 784.950 ;
        RECT 307.950 783.450 310.050 784.050 ;
        RECT 287.400 782.400 310.050 783.450 ;
        RECT 226.950 781.950 229.050 782.400 ;
        RECT 235.950 781.950 238.050 782.400 ;
        RECT 307.950 781.950 310.050 782.400 ;
        RECT 343.950 783.450 346.050 784.050 ;
        RECT 358.950 783.450 361.050 784.050 ;
        RECT 343.950 782.400 361.050 783.450 ;
        RECT 343.950 781.950 346.050 782.400 ;
        RECT 358.950 781.950 361.050 782.400 ;
        RECT 364.950 783.450 367.050 784.050 ;
        RECT 377.400 783.450 378.450 785.400 ;
        RECT 382.950 784.950 385.050 785.400 ;
        RECT 403.950 786.450 406.050 787.050 ;
        RECT 415.950 786.450 418.050 787.050 ;
        RECT 403.950 785.400 418.050 786.450 ;
        RECT 403.950 784.950 406.050 785.400 ;
        RECT 415.950 784.950 418.050 785.400 ;
        RECT 424.950 786.450 427.050 787.050 ;
        RECT 439.950 786.450 442.050 787.050 ;
        RECT 424.950 785.400 442.050 786.450 ;
        RECT 424.950 784.950 427.050 785.400 ;
        RECT 439.950 784.950 442.050 785.400 ;
        RECT 448.950 786.450 451.050 787.050 ;
        RECT 478.950 786.450 481.050 787.050 ;
        RECT 448.950 785.400 481.050 786.450 ;
        RECT 448.950 784.950 451.050 785.400 ;
        RECT 478.950 784.950 481.050 785.400 ;
        RECT 484.950 786.450 487.050 787.050 ;
        RECT 490.950 786.450 493.050 787.050 ;
        RECT 505.950 786.450 508.050 787.050 ;
        RECT 484.950 785.400 508.050 786.450 ;
        RECT 484.950 784.950 487.050 785.400 ;
        RECT 490.950 784.950 493.050 785.400 ;
        RECT 505.950 784.950 508.050 785.400 ;
        RECT 529.950 786.450 532.050 787.050 ;
        RECT 535.950 786.450 538.050 787.050 ;
        RECT 529.950 785.400 538.050 786.450 ;
        RECT 529.950 784.950 532.050 785.400 ;
        RECT 535.950 784.950 538.050 785.400 ;
        RECT 541.950 786.450 544.050 787.050 ;
        RECT 550.950 786.450 553.050 787.050 ;
        RECT 541.950 785.400 553.050 786.450 ;
        RECT 541.950 784.950 544.050 785.400 ;
        RECT 550.950 784.950 553.050 785.400 ;
        RECT 556.950 786.450 559.050 787.050 ;
        RECT 571.950 786.450 574.050 786.900 ;
        RECT 670.950 786.450 673.050 787.200 ;
        RECT 556.950 785.400 673.050 786.450 ;
        RECT 556.950 784.950 559.050 785.400 ;
        RECT 571.950 784.800 574.050 785.400 ;
        RECT 670.950 785.100 673.050 785.400 ;
        RECT 703.950 786.450 706.050 787.050 ;
        RECT 712.950 786.450 715.050 787.050 ;
        RECT 703.950 785.400 715.050 786.450 ;
        RECT 703.950 784.950 706.050 785.400 ;
        RECT 712.950 784.950 715.050 785.400 ;
        RECT 724.950 786.450 727.050 787.050 ;
        RECT 733.950 786.450 736.050 787.050 ;
        RECT 724.950 785.400 789.450 786.450 ;
        RECT 724.950 784.950 727.050 785.400 ;
        RECT 733.950 784.950 736.050 785.400 ;
        RECT 397.950 783.450 400.050 784.050 ;
        RECT 442.950 783.450 445.050 784.050 ;
        RECT 364.950 782.400 378.450 783.450 ;
        RECT 380.400 782.400 445.050 783.450 ;
        RECT 364.950 781.950 367.050 782.400 ;
        RECT 106.950 780.450 109.050 781.050 ;
        RECT 118.950 780.450 121.050 781.050 ;
        RECT 106.950 779.400 121.050 780.450 ;
        RECT 106.950 778.950 109.050 779.400 ;
        RECT 118.950 778.950 121.050 779.400 ;
        RECT 169.950 780.450 172.050 781.050 ;
        RECT 193.950 780.450 196.050 781.050 ;
        RECT 169.950 779.400 196.050 780.450 ;
        RECT 169.950 778.950 172.050 779.400 ;
        RECT 193.950 778.950 196.050 779.400 ;
        RECT 199.950 780.450 202.050 781.050 ;
        RECT 211.950 780.450 214.050 781.050 ;
        RECT 199.950 779.400 214.050 780.450 ;
        RECT 199.950 778.950 202.050 779.400 ;
        RECT 211.950 778.950 214.050 779.400 ;
        RECT 232.950 780.450 235.050 781.050 ;
        RECT 380.400 780.450 381.450 782.400 ;
        RECT 397.950 781.950 400.050 782.400 ;
        RECT 442.950 781.950 445.050 782.400 ;
        RECT 457.950 783.450 460.050 784.050 ;
        RECT 499.800 783.450 501.900 784.050 ;
        RECT 457.950 782.400 501.900 783.450 ;
        RECT 457.950 781.950 460.050 782.400 ;
        RECT 499.800 781.950 501.900 782.400 ;
        RECT 503.100 783.450 505.200 784.050 ;
        RECT 589.950 783.450 592.050 784.050 ;
        RECT 503.100 782.400 592.050 783.450 ;
        RECT 503.100 781.950 505.200 782.400 ;
        RECT 589.950 781.950 592.050 782.400 ;
        RECT 598.950 783.450 601.050 784.050 ;
        RECT 610.950 783.450 613.050 784.050 ;
        RECT 598.950 782.400 613.050 783.450 ;
        RECT 598.950 781.950 601.050 782.400 ;
        RECT 610.950 781.950 613.050 782.400 ;
        RECT 616.950 783.450 619.050 784.050 ;
        RECT 628.950 783.450 631.050 784.050 ;
        RECT 661.950 783.450 664.050 784.050 ;
        RECT 616.950 782.400 631.050 783.450 ;
        RECT 616.950 781.950 619.050 782.400 ;
        RECT 628.950 781.950 631.050 782.400 ;
        RECT 644.400 782.400 664.050 783.450 ;
        RECT 232.950 779.400 381.450 780.450 ;
        RECT 382.950 780.450 385.050 781.050 ;
        RECT 415.800 780.450 417.900 781.050 ;
        RECT 382.950 779.400 417.900 780.450 ;
        RECT 232.950 778.950 235.050 779.400 ;
        RECT 382.950 778.950 385.050 779.400 ;
        RECT 415.800 778.950 417.900 779.400 ;
        RECT 419.100 780.450 421.200 781.050 ;
        RECT 448.950 780.450 451.050 781.050 ;
        RECT 458.400 780.450 459.450 781.950 ;
        RECT 644.400 780.450 645.450 782.400 ;
        RECT 661.950 781.950 664.050 782.400 ;
        RECT 670.950 783.450 673.050 783.900 ;
        RECT 703.950 783.450 706.050 784.050 ;
        RECT 670.950 782.400 706.050 783.450 ;
        RECT 670.950 781.800 673.050 782.400 ;
        RECT 703.950 781.950 706.050 782.400 ;
        RECT 709.950 783.450 712.050 784.050 ;
        RECT 727.950 783.450 730.050 784.050 ;
        RECT 709.950 782.400 730.050 783.450 ;
        RECT 709.950 781.950 712.050 782.400 ;
        RECT 727.950 781.950 730.050 782.400 ;
        RECT 736.950 783.450 739.050 784.050 ;
        RECT 754.950 783.450 757.050 784.050 ;
        RECT 736.950 782.400 757.050 783.450 ;
        RECT 788.400 783.450 789.450 785.400 ;
        RECT 790.950 784.950 796.050 787.050 ;
        RECT 797.400 786.450 798.450 788.400 ;
        RECT 817.950 788.400 840.450 789.450 ;
        RECT 817.950 787.950 820.050 788.400 ;
        RECT 859.950 786.450 862.050 787.050 ;
        RECT 797.400 785.400 862.050 786.450 ;
        RECT 859.950 784.950 862.050 785.400 ;
        RECT 889.950 786.450 892.050 787.050 ;
        RECT 898.950 786.450 901.050 787.050 ;
        RECT 889.950 785.400 901.050 786.450 ;
        RECT 889.950 784.950 892.050 785.400 ;
        RECT 898.950 784.950 901.050 785.400 ;
        RECT 883.950 783.450 886.050 784.050 ;
        RECT 788.400 782.400 886.050 783.450 ;
        RECT 736.950 781.950 739.050 782.400 ;
        RECT 754.950 781.950 757.050 782.400 ;
        RECT 883.950 781.950 886.050 782.400 ;
        RECT 706.950 780.450 709.050 781.050 ;
        RECT 790.950 780.450 793.050 781.050 ;
        RECT 419.100 779.400 435.450 780.450 ;
        RECT 419.100 778.950 421.200 779.400 ;
        RECT 434.400 778.050 435.450 779.400 ;
        RECT 448.950 779.400 459.450 780.450 ;
        RECT 536.400 779.400 645.450 780.450 ;
        RECT 653.400 779.400 709.050 780.450 ;
        RECT 448.950 778.950 451.050 779.400 ;
        RECT 16.950 777.450 19.050 778.050 ;
        RECT 37.950 777.450 40.050 778.050 ;
        RECT 82.950 777.450 85.050 778.050 ;
        RECT 253.950 777.450 256.050 778.050 ;
        RECT 16.950 776.400 256.050 777.450 ;
        RECT 16.950 775.950 19.050 776.400 ;
        RECT 37.950 775.950 40.050 776.400 ;
        RECT 82.950 775.950 85.050 776.400 ;
        RECT 253.950 775.950 256.050 776.400 ;
        RECT 280.950 777.450 283.050 778.050 ;
        RECT 313.950 777.450 316.050 778.050 ;
        RECT 280.950 776.400 316.050 777.450 ;
        RECT 280.950 775.950 283.050 776.400 ;
        RECT 313.950 775.950 316.050 776.400 ;
        RECT 319.950 777.450 322.050 778.050 ;
        RECT 406.950 777.450 409.050 778.050 ;
        RECT 319.950 776.400 409.050 777.450 ;
        RECT 319.950 775.950 322.050 776.400 ;
        RECT 406.950 775.950 409.050 776.400 ;
        RECT 433.950 777.450 436.050 778.050 ;
        RECT 439.800 777.450 441.900 778.050 ;
        RECT 433.950 776.400 441.900 777.450 ;
        RECT 433.950 775.950 436.050 776.400 ;
        RECT 439.800 775.950 441.900 776.400 ;
        RECT 443.100 777.450 445.200 778.050 ;
        RECT 469.950 777.450 472.050 778.050 ;
        RECT 493.950 777.450 496.050 778.050 ;
        RECT 536.400 777.450 537.450 779.400 ;
        RECT 443.100 776.400 537.450 777.450 ;
        RECT 538.950 777.450 541.050 778.050 ;
        RECT 653.400 777.450 654.450 779.400 ;
        RECT 706.950 778.950 709.050 779.400 ;
        RECT 776.400 779.400 793.050 780.450 ;
        RECT 538.950 776.400 654.450 777.450 ;
        RECT 676.950 777.450 679.050 778.050 ;
        RECT 739.950 777.450 742.050 778.050 ;
        RECT 676.950 776.400 742.050 777.450 ;
        RECT 443.100 775.950 445.200 776.400 ;
        RECT 469.950 775.950 472.050 776.400 ;
        RECT 493.950 775.950 496.050 776.400 ;
        RECT 538.950 775.950 541.050 776.400 ;
        RECT 676.950 775.950 679.050 776.400 ;
        RECT 739.950 775.950 742.050 776.400 ;
        RECT 754.950 777.450 757.050 778.050 ;
        RECT 776.400 777.450 777.450 779.400 ;
        RECT 790.950 778.950 793.050 779.400 ;
        RECT 754.950 776.400 777.450 777.450 ;
        RECT 778.950 777.450 781.050 778.050 ;
        RECT 826.950 777.450 829.050 778.050 ;
        RECT 778.950 776.400 829.050 777.450 ;
        RECT 754.950 775.950 757.050 776.400 ;
        RECT 778.950 775.950 781.050 776.400 ;
        RECT 826.950 775.950 829.050 776.400 ;
        RECT 85.950 774.450 88.050 775.050 ;
        RECT 85.950 773.400 108.450 774.450 ;
        RECT 85.950 772.950 88.050 773.400 ;
        RECT 107.400 772.050 108.450 773.400 ;
        RECT 208.950 772.950 214.050 775.050 ;
        RECT 217.950 774.450 220.050 775.050 ;
        RECT 235.950 774.450 238.050 775.050 ;
        RECT 217.950 773.400 238.050 774.450 ;
        RECT 217.950 772.950 220.050 773.400 ;
        RECT 235.950 772.950 238.050 773.400 ;
        RECT 265.950 774.450 268.050 775.050 ;
        RECT 286.950 774.450 289.050 775.050 ;
        RECT 310.950 774.450 313.050 775.050 ;
        RECT 352.950 774.450 355.050 775.050 ;
        RECT 364.800 774.450 366.900 775.050 ;
        RECT 265.950 773.400 355.050 774.450 ;
        RECT 265.950 772.950 268.050 773.400 ;
        RECT 286.950 772.950 289.050 773.400 ;
        RECT 310.950 772.950 313.050 773.400 ;
        RECT 352.950 772.950 355.050 773.400 ;
        RECT 356.400 773.400 366.900 774.450 ;
        RECT 97.950 769.950 103.050 772.050 ;
        RECT 106.950 771.450 109.050 772.050 ;
        RECT 124.950 771.450 127.050 772.050 ;
        RECT 172.950 771.450 175.050 772.050 ;
        RECT 106.950 770.400 175.050 771.450 ;
        RECT 106.950 769.950 109.050 770.400 ;
        RECT 124.950 769.950 127.050 770.400 ;
        RECT 172.950 769.950 175.050 770.400 ;
        RECT 178.950 771.450 181.050 772.050 ;
        RECT 184.800 771.450 186.900 772.050 ;
        RECT 178.950 770.400 186.900 771.450 ;
        RECT 178.950 769.950 181.050 770.400 ;
        RECT 184.800 769.950 186.900 770.400 ;
        RECT 188.100 771.450 190.200 772.050 ;
        RECT 193.950 771.450 196.050 772.050 ;
        RECT 188.100 770.400 196.050 771.450 ;
        RECT 188.100 769.950 190.200 770.400 ;
        RECT 193.950 769.950 196.050 770.400 ;
        RECT 277.950 771.450 280.050 772.050 ;
        RECT 292.950 771.450 295.050 772.050 ;
        RECT 356.400 771.450 357.450 773.400 ;
        RECT 364.800 772.950 366.900 773.400 ;
        RECT 368.100 774.450 370.200 775.050 ;
        RECT 376.950 774.450 379.050 775.050 ;
        RECT 385.950 774.450 388.050 775.050 ;
        RECT 368.100 773.400 388.050 774.450 ;
        RECT 368.100 772.950 370.200 773.400 ;
        RECT 376.950 772.950 379.050 773.400 ;
        RECT 385.950 772.950 388.050 773.400 ;
        RECT 400.950 774.450 403.050 775.050 ;
        RECT 490.950 774.450 493.050 775.050 ;
        RECT 400.950 773.400 493.050 774.450 ;
        RECT 400.950 772.950 403.050 773.400 ;
        RECT 490.950 772.950 493.050 773.400 ;
        RECT 496.950 774.450 499.050 775.050 ;
        RECT 547.950 774.450 550.050 775.050 ;
        RECT 496.950 773.400 550.050 774.450 ;
        RECT 496.950 772.950 499.050 773.400 ;
        RECT 547.950 772.950 550.050 773.400 ;
        RECT 610.950 774.450 613.050 775.050 ;
        RECT 640.950 774.450 643.050 775.200 ;
        RECT 730.950 774.450 733.050 775.050 ;
        RECT 610.950 773.400 643.050 774.450 ;
        RECT 610.950 772.950 613.050 773.400 ;
        RECT 640.950 773.100 643.050 773.400 ;
        RECT 701.400 773.400 733.050 774.450 ;
        RECT 277.950 770.400 291.450 771.450 ;
        RECT 277.950 769.950 280.050 770.400 ;
        RECT 290.400 766.050 291.450 770.400 ;
        RECT 292.950 770.400 357.450 771.450 ;
        RECT 361.950 771.450 364.050 772.050 ;
        RECT 394.950 771.450 397.050 772.050 ;
        RECT 361.950 770.400 397.050 771.450 ;
        RECT 292.950 769.950 295.050 770.400 ;
        RECT 361.950 769.950 364.050 770.400 ;
        RECT 394.950 769.950 397.050 770.400 ;
        RECT 409.950 771.450 412.050 772.050 ;
        RECT 460.950 771.450 463.050 772.050 ;
        RECT 409.950 770.400 463.050 771.450 ;
        RECT 409.950 769.950 412.050 770.400 ;
        RECT 460.950 769.950 463.050 770.400 ;
        RECT 466.950 771.450 469.050 772.050 ;
        RECT 484.950 771.450 487.050 772.050 ;
        RECT 466.950 770.400 487.050 771.450 ;
        RECT 466.950 769.950 469.050 770.400 ;
        RECT 484.950 769.950 487.050 770.400 ;
        RECT 496.950 771.450 499.050 772.050 ;
        RECT 502.800 771.450 504.900 772.050 ;
        RECT 496.950 770.400 504.900 771.450 ;
        RECT 496.950 769.950 499.050 770.400 ;
        RECT 502.800 769.950 504.900 770.400 ;
        RECT 506.100 771.450 508.200 772.050 ;
        RECT 532.950 771.450 535.050 772.050 ;
        RECT 506.100 770.400 535.050 771.450 ;
        RECT 506.100 769.950 508.200 770.400 ;
        RECT 532.950 769.950 535.050 770.400 ;
        RECT 550.950 771.450 553.050 772.050 ;
        RECT 559.950 771.450 562.050 772.050 ;
        RECT 550.950 770.400 562.050 771.450 ;
        RECT 550.950 769.950 553.050 770.400 ;
        RECT 559.950 769.950 562.050 770.400 ;
        RECT 613.950 771.450 616.050 772.050 ;
        RECT 640.950 771.450 643.050 771.900 ;
        RECT 613.950 770.400 643.050 771.450 ;
        RECT 613.950 769.950 616.050 770.400 ;
        RECT 640.950 769.800 643.050 770.400 ;
        RECT 652.950 771.450 655.050 772.050 ;
        RECT 667.950 771.450 670.050 772.050 ;
        RECT 652.950 770.400 670.050 771.450 ;
        RECT 652.950 769.950 655.050 770.400 ;
        RECT 667.950 769.950 670.050 770.400 ;
        RECT 688.950 771.450 691.050 772.050 ;
        RECT 701.400 771.450 702.450 773.400 ;
        RECT 730.950 772.950 733.050 773.400 ;
        RECT 688.950 770.400 702.450 771.450 ;
        RECT 703.950 771.450 706.050 772.050 ;
        RECT 724.950 771.450 727.050 772.050 ;
        RECT 703.950 770.400 727.050 771.450 ;
        RECT 688.950 769.950 691.050 770.400 ;
        RECT 445.950 768.450 448.050 769.050 ;
        RECT 451.950 768.450 454.050 769.050 ;
        RECT 514.950 768.450 517.050 769.050 ;
        RECT 445.950 767.400 454.050 768.450 ;
        RECT 445.950 766.950 448.050 767.400 ;
        RECT 451.950 766.950 454.050 767.400 ;
        RECT 508.950 767.400 517.050 768.450 ;
        RECT 13.950 765.450 16.050 766.050 ;
        RECT 22.950 765.450 25.050 766.050 ;
        RECT 13.950 764.400 25.050 765.450 ;
        RECT 13.950 763.950 16.050 764.400 ;
        RECT 22.950 763.950 25.050 764.400 ;
        RECT 28.950 763.950 31.050 766.050 ;
        RECT 34.950 763.950 37.050 766.050 ;
        RECT 55.950 763.950 58.050 766.050 ;
        RECT 61.950 763.950 64.050 766.050 ;
        RECT 82.950 763.950 85.050 766.050 ;
        RECT 88.950 765.450 91.050 766.050 ;
        RECT 100.950 765.450 103.050 766.050 ;
        RECT 88.950 764.400 103.050 765.450 ;
        RECT 88.950 763.950 91.050 764.400 ;
        RECT 100.950 763.950 103.050 764.400 ;
        RECT 106.950 763.950 109.050 766.050 ;
        RECT 112.950 763.950 115.050 766.050 ;
        RECT 124.950 763.950 127.050 766.050 ;
        RECT 130.950 763.950 133.050 766.050 ;
        RECT 154.950 763.950 157.050 766.050 ;
        RECT 160.950 763.950 163.050 766.050 ;
        RECT 166.950 765.450 169.050 766.050 ;
        RECT 178.950 765.450 181.050 766.050 ;
        RECT 166.950 764.400 181.050 765.450 ;
        RECT 166.950 763.950 169.050 764.400 ;
        RECT 178.950 763.950 181.050 764.400 ;
        RECT 184.950 763.950 190.050 766.050 ;
        RECT 196.950 763.950 199.050 766.050 ;
        RECT 220.950 763.950 223.050 766.050 ;
        RECT 226.950 763.950 229.050 766.050 ;
        RECT 247.950 763.950 250.050 766.050 ;
        RECT 265.950 763.950 268.050 766.050 ;
        RECT 271.950 763.950 274.050 766.050 ;
        RECT 280.950 763.950 286.050 766.050 ;
        RECT 289.950 763.950 292.050 766.050 ;
        RECT 307.950 763.950 310.050 766.050 ;
        RECT 313.950 765.450 316.050 766.050 ;
        RECT 328.950 765.450 331.050 766.050 ;
        RECT 313.950 764.400 331.050 765.450 ;
        RECT 313.950 763.950 316.050 764.400 ;
        RECT 328.950 763.950 331.050 764.400 ;
        RECT 334.950 763.950 337.050 766.050 ;
        RECT 340.950 763.950 343.050 766.050 ;
        RECT 361.950 763.950 364.050 766.050 ;
        RECT 367.950 763.950 370.050 766.050 ;
        RECT 385.950 763.950 388.050 766.050 ;
        RECT 391.950 763.950 394.050 766.050 ;
        RECT 409.950 763.950 412.050 766.050 ;
        RECT 415.950 763.950 418.050 766.050 ;
        RECT 427.950 763.950 430.050 766.050 ;
        RECT 433.950 763.950 436.050 766.050 ;
        RECT 454.950 763.950 457.050 766.050 ;
        RECT 460.950 763.950 463.050 766.050 ;
        RECT 475.950 763.950 478.050 766.050 ;
        RECT 481.950 763.950 484.050 766.050 ;
        RECT 502.950 763.950 505.050 766.050 ;
        RECT 508.950 763.950 511.050 767.400 ;
        RECT 514.950 766.950 517.050 767.400 ;
        RECT 661.950 768.450 664.050 769.050 ;
        RECT 673.950 768.450 676.050 769.050 ;
        RECT 661.950 767.400 676.050 768.450 ;
        RECT 695.400 768.450 696.450 770.400 ;
        RECT 703.950 769.950 706.050 770.400 ;
        RECT 724.950 769.950 727.050 770.400 ;
        RECT 739.950 771.450 742.050 771.900 ;
        RECT 751.950 771.450 754.050 772.050 ;
        RECT 739.950 770.400 754.050 771.450 ;
        RECT 739.950 769.800 742.050 770.400 ;
        RECT 751.950 769.950 754.050 770.400 ;
        RECT 766.950 771.450 769.050 772.050 ;
        RECT 775.950 771.450 778.050 772.050 ;
        RECT 766.950 770.400 778.050 771.450 ;
        RECT 766.950 769.950 769.050 770.400 ;
        RECT 775.950 769.950 778.050 770.400 ;
        RECT 784.950 771.450 787.050 772.050 ;
        RECT 793.950 771.450 796.050 772.050 ;
        RECT 784.950 770.400 796.050 771.450 ;
        RECT 784.950 769.950 787.050 770.400 ;
        RECT 793.950 769.950 796.050 770.400 ;
        RECT 808.950 771.450 811.050 772.050 ;
        RECT 820.950 771.450 823.050 772.050 ;
        RECT 808.950 770.400 823.050 771.450 ;
        RECT 808.950 769.950 811.050 770.400 ;
        RECT 820.950 769.950 823.050 770.400 ;
        RECT 895.950 771.450 898.050 772.050 ;
        RECT 904.950 771.450 907.050 772.050 ;
        RECT 895.950 770.400 907.050 771.450 ;
        RECT 895.950 769.950 898.050 770.400 ;
        RECT 904.950 769.950 907.050 770.400 ;
        RECT 700.950 768.450 703.050 769.050 ;
        RECT 695.400 767.400 703.050 768.450 ;
        RECT 661.950 766.950 664.050 767.400 ;
        RECT 673.950 766.950 676.050 767.400 ;
        RECT 700.950 766.950 703.050 767.400 ;
        RECT 826.950 768.450 829.050 769.050 ;
        RECT 853.950 768.450 856.050 769.050 ;
        RECT 826.950 767.400 856.050 768.450 ;
        RECT 826.950 766.950 829.050 767.400 ;
        RECT 853.950 766.950 856.050 767.400 ;
        RECT 886.950 768.450 889.050 769.050 ;
        RECT 910.950 768.450 913.050 769.050 ;
        RECT 886.950 767.400 913.050 768.450 ;
        RECT 886.950 766.950 889.050 767.400 ;
        RECT 910.950 766.950 913.050 767.400 ;
        RECT 529.950 765.450 532.050 766.050 ;
        RECT 534.000 765.450 538.050 766.050 ;
        RECT 529.950 764.400 538.050 765.450 ;
        RECT 529.950 763.950 532.050 764.400 ;
        RECT 534.000 763.950 538.050 764.400 ;
        RECT 544.950 763.950 550.050 766.050 ;
        RECT 553.950 763.950 556.050 766.050 ;
        RECT 559.950 765.450 564.000 766.050 ;
        RECT 565.950 765.450 568.050 766.050 ;
        RECT 559.950 764.400 568.050 765.450 ;
        RECT 559.950 763.950 564.000 764.400 ;
        RECT 565.950 763.950 568.050 764.400 ;
        RECT 571.950 763.950 574.050 766.050 ;
        RECT 592.950 763.950 595.050 766.050 ;
        RECT 598.950 763.950 601.050 766.050 ;
        RECT 616.950 763.950 619.050 766.050 ;
        RECT 622.950 763.950 625.050 766.050 ;
        RECT 637.950 763.950 640.050 766.050 ;
        RECT 643.950 765.450 646.050 766.050 ;
        RECT 652.950 765.450 655.050 766.050 ;
        RECT 643.950 764.400 655.050 765.450 ;
        RECT 643.950 763.950 646.050 764.400 ;
        RECT 652.950 763.950 655.050 764.400 ;
        RECT 682.950 763.950 685.050 766.050 ;
        RECT 688.950 763.950 691.050 766.050 ;
        RECT 709.950 765.450 712.050 766.050 ;
        RECT 718.950 765.450 721.050 766.050 ;
        RECT 709.950 764.400 721.050 765.450 ;
        RECT 709.950 763.950 712.050 764.400 ;
        RECT 718.950 763.950 721.050 764.400 ;
        RECT 724.950 763.950 727.050 766.050 ;
        RECT 730.950 763.950 733.050 766.050 ;
        RECT 766.950 763.950 769.050 766.050 ;
        RECT 772.950 763.950 775.050 766.050 ;
        RECT 790.950 763.950 793.050 766.050 ;
        RECT 796.950 765.450 799.050 766.050 ;
        RECT 808.950 765.450 811.050 766.050 ;
        RECT 796.950 764.400 811.050 765.450 ;
        RECT 796.950 763.950 799.050 764.400 ;
        RECT 808.950 763.950 811.050 764.400 ;
        RECT 814.950 763.950 817.050 766.050 ;
        RECT 820.950 763.950 823.050 766.050 ;
        RECT 856.950 763.950 859.050 766.050 ;
        RECT 862.950 763.950 865.050 766.050 ;
        RECT 13.950 760.950 16.050 762.750 ;
        RECT 28.950 760.950 31.050 762.750 ;
        RECT 34.950 760.950 37.050 762.750 ;
        RECT 55.950 760.950 58.050 762.750 ;
        RECT 61.950 760.950 64.050 762.750 ;
        RECT 82.950 760.950 85.050 762.750 ;
        RECT 88.950 760.950 91.050 762.750 ;
        RECT 106.950 760.950 109.050 762.750 ;
        RECT 112.950 760.950 115.050 762.750 ;
        RECT 16.950 758.250 19.050 760.050 ;
        RECT 31.950 758.250 34.050 760.050 ;
        RECT 37.950 758.250 40.050 760.050 ;
        RECT 58.950 758.250 61.050 760.050 ;
        RECT 64.950 758.250 67.050 760.050 ;
        RECT 79.950 758.250 82.050 760.050 ;
        RECT 85.950 758.250 88.050 760.050 ;
        RECT 103.950 758.250 106.050 760.050 ;
        RECT 109.950 758.250 112.050 760.050 ;
        RECT 118.950 757.950 121.050 763.050 ;
        RECT 124.950 760.950 127.050 762.750 ;
        RECT 130.950 760.950 133.050 762.750 ;
        RECT 127.950 758.250 130.050 760.050 ;
        RECT 133.950 758.250 136.050 760.050 ;
        RECT 145.950 757.950 148.050 763.050 ;
        RECT 154.950 760.950 157.050 762.750 ;
        RECT 160.950 760.950 163.050 762.750 ;
        RECT 178.950 760.950 181.050 762.750 ;
        RECT 184.950 760.950 187.050 762.750 ;
        RECT 196.950 760.950 199.050 762.750 ;
        RECT 202.950 760.950 205.050 762.750 ;
        RECT 220.950 760.950 223.050 762.750 ;
        RECT 226.950 760.950 229.050 762.750 ;
        RECT 247.950 760.950 250.050 762.750 ;
        RECT 265.950 760.950 268.050 762.750 ;
        RECT 271.950 760.950 274.050 762.750 ;
        RECT 283.950 760.950 286.050 762.750 ;
        RECT 289.950 760.950 292.050 762.750 ;
        RECT 307.950 760.950 310.050 762.750 ;
        RECT 313.950 760.950 316.050 762.750 ;
        RECT 334.950 760.950 337.050 762.750 ;
        RECT 340.950 760.950 343.050 762.750 ;
        RECT 361.950 760.950 364.050 762.750 ;
        RECT 367.950 760.950 370.050 762.750 ;
        RECT 373.950 762.450 376.050 763.050 ;
        RECT 379.950 762.450 382.050 763.050 ;
        RECT 373.950 761.400 382.050 762.450 ;
        RECT 373.950 760.950 376.050 761.400 ;
        RECT 379.950 760.950 382.050 761.400 ;
        RECT 385.950 760.950 388.050 762.750 ;
        RECT 391.950 760.950 394.050 762.750 ;
        RECT 409.950 760.950 412.050 762.750 ;
        RECT 415.950 760.950 418.050 762.750 ;
        RECT 427.950 760.950 430.050 762.750 ;
        RECT 433.950 760.950 436.050 762.750 ;
        RECT 454.950 760.950 457.050 762.750 ;
        RECT 460.950 760.950 463.050 762.750 ;
        RECT 475.950 760.950 478.050 762.750 ;
        RECT 481.950 760.950 484.050 762.750 ;
        RECT 502.950 760.950 505.050 762.750 ;
        RECT 508.950 760.950 511.050 762.750 ;
        RECT 529.950 760.950 532.050 762.750 ;
        RECT 547.950 760.950 550.050 762.750 ;
        RECT 553.950 760.950 556.050 762.750 ;
        RECT 565.950 760.950 568.050 762.750 ;
        RECT 571.950 760.950 574.050 762.750 ;
        RECT 592.950 760.950 595.050 762.750 ;
        RECT 598.950 760.950 601.050 762.750 ;
        RECT 616.950 760.950 619.050 762.750 ;
        RECT 622.950 760.950 625.050 762.750 ;
        RECT 637.950 760.950 640.050 762.750 ;
        RECT 643.950 760.950 646.050 762.750 ;
        RECT 661.950 762.450 664.050 763.050 ;
        RECT 670.950 762.450 673.050 763.050 ;
        RECT 661.950 761.400 673.050 762.450 ;
        RECT 661.950 760.950 664.050 761.400 ;
        RECT 670.950 760.950 673.050 761.400 ;
        RECT 682.950 760.950 685.050 762.750 ;
        RECT 688.950 760.950 691.050 762.750 ;
        RECT 709.950 760.950 712.050 762.750 ;
        RECT 724.950 760.950 727.050 762.750 ;
        RECT 730.950 760.950 733.050 762.750 ;
        RECT 754.950 760.950 757.050 762.750 ;
        RECT 766.950 760.950 769.050 762.750 ;
        RECT 772.950 760.950 775.050 762.750 ;
        RECT 790.950 760.950 793.050 762.750 ;
        RECT 796.950 760.950 799.050 762.750 ;
        RECT 814.950 760.950 817.050 762.750 ;
        RECT 820.950 760.950 823.050 762.750 ;
        RECT 856.950 760.950 859.050 762.750 ;
        RECT 862.950 760.950 865.050 762.750 ;
        RECT 901.950 762.450 904.050 763.050 ;
        RECT 910.950 762.450 913.050 763.050 ;
        RECT 901.950 761.400 913.050 762.450 ;
        RECT 901.950 760.950 904.050 761.400 ;
        RECT 910.950 760.950 913.050 761.400 ;
        RECT 394.950 760.050 397.050 760.200 ;
        RECT 151.950 758.250 154.050 760.050 ;
        RECT 157.950 758.250 160.050 760.050 ;
        RECT 163.950 759.450 166.050 760.050 ;
        RECT 169.950 759.450 172.050 760.050 ;
        RECT 163.950 758.400 172.050 759.450 ;
        RECT 163.950 757.950 166.050 758.400 ;
        RECT 169.950 757.950 172.050 758.400 ;
        RECT 175.950 758.250 178.050 760.050 ;
        RECT 181.950 758.250 184.050 760.050 ;
        RECT 199.950 758.250 202.050 760.050 ;
        RECT 223.950 758.250 226.050 760.050 ;
        RECT 229.950 758.250 232.050 760.050 ;
        RECT 244.950 758.250 247.050 760.050 ;
        RECT 262.950 758.250 265.050 760.050 ;
        RECT 268.950 758.250 271.050 760.050 ;
        RECT 286.950 758.250 289.050 760.050 ;
        RECT 292.950 758.250 295.050 760.050 ;
        RECT 310.950 758.250 313.050 760.050 ;
        RECT 316.950 758.250 319.050 760.050 ;
        RECT 337.950 758.250 340.050 760.050 ;
        RECT 343.950 758.250 346.050 760.050 ;
        RECT 358.950 758.250 361.050 760.050 ;
        RECT 364.950 758.250 367.050 760.050 ;
        RECT 382.950 758.250 385.050 760.050 ;
        RECT 388.950 758.250 391.050 760.050 ;
        RECT 394.950 758.100 400.050 760.050 ;
        RECT 406.950 758.250 409.050 760.050 ;
        RECT 412.950 758.250 415.050 760.050 ;
        RECT 430.950 758.250 433.050 760.050 ;
        RECT 436.950 758.250 439.050 760.050 ;
        RECT 451.950 758.250 454.050 760.050 ;
        RECT 457.950 758.250 460.050 760.050 ;
        RECT 396.000 757.950 400.050 758.100 ;
        RECT 463.950 757.950 469.050 760.050 ;
        RECT 478.950 758.250 481.050 760.050 ;
        RECT 484.950 758.250 487.050 760.050 ;
        RECT 505.950 758.250 508.050 760.050 ;
        RECT 511.950 758.250 514.050 760.050 ;
        RECT 526.950 758.250 529.050 760.050 ;
        RECT 544.950 758.250 547.050 760.050 ;
        RECT 550.950 758.250 553.050 760.050 ;
        RECT 568.950 758.250 571.050 760.050 ;
        RECT 574.950 758.250 577.050 760.050 ;
        RECT 595.950 758.250 598.050 760.050 ;
        RECT 601.950 758.250 604.050 760.050 ;
        RECT 619.950 758.250 622.050 760.050 ;
        RECT 640.950 758.250 643.050 760.050 ;
        RECT 646.950 758.250 649.050 760.050 ;
        RECT 661.950 757.950 664.050 759.750 ;
        RECT 679.950 758.250 682.050 760.050 ;
        RECT 685.950 758.250 688.050 760.050 ;
        RECT 691.950 758.250 694.050 760.050 ;
        RECT 712.950 758.250 715.050 760.050 ;
        RECT 727.950 758.250 730.050 760.050 ;
        RECT 733.950 758.250 736.050 760.050 ;
        RECT 751.950 758.250 754.050 760.050 ;
        RECT 769.950 758.250 772.050 760.050 ;
        RECT 787.950 758.250 790.050 760.050 ;
        RECT 793.950 758.250 796.050 760.050 ;
        RECT 817.950 758.250 820.050 760.050 ;
        RECT 832.950 758.250 835.050 760.050 ;
        RECT 838.950 757.950 841.050 759.750 ;
        RECT 853.950 758.250 856.050 760.050 ;
        RECT 859.950 758.250 862.050 760.050 ;
        RECT 877.950 758.250 880.050 760.050 ;
        RECT 892.950 759.900 897.000 760.050 ;
        RECT 883.950 757.950 886.050 759.750 ;
        RECT 892.950 757.950 898.050 759.900 ;
        RECT 901.950 757.950 904.050 759.750 ;
        RECT 895.950 757.800 898.050 757.950 ;
        RECT 16.950 754.950 19.050 757.050 ;
        RECT 31.950 754.950 34.050 757.050 ;
        RECT 37.950 754.950 40.050 757.050 ;
        RECT 43.950 756.450 46.050 757.050 ;
        RECT 58.950 756.450 61.050 757.050 ;
        RECT 43.950 755.400 61.050 756.450 ;
        RECT 43.950 754.950 46.050 755.400 ;
        RECT 58.950 754.950 61.050 755.400 ;
        RECT 64.950 754.950 67.050 757.050 ;
        RECT 73.950 756.450 78.000 757.050 ;
        RECT 79.950 756.450 82.050 757.050 ;
        RECT 73.950 755.400 82.050 756.450 ;
        RECT 73.950 754.950 78.000 755.400 ;
        RECT 79.950 754.950 82.050 755.400 ;
        RECT 85.950 754.950 88.050 757.050 ;
        RECT 91.950 756.450 94.050 757.050 ;
        RECT 103.950 756.450 106.050 757.050 ;
        RECT 91.950 755.400 106.050 756.450 ;
        RECT 91.950 754.950 94.050 755.400 ;
        RECT 103.950 754.950 106.050 755.400 ;
        RECT 109.950 756.450 112.050 757.050 ;
        RECT 121.950 756.450 124.050 757.050 ;
        RECT 109.950 755.400 124.050 756.450 ;
        RECT 109.950 754.950 112.050 755.400 ;
        RECT 121.950 754.950 124.050 755.400 ;
        RECT 127.950 754.950 130.050 757.050 ;
        RECT 133.950 751.950 136.050 757.050 ;
        RECT 139.950 756.450 142.050 757.050 ;
        RECT 151.950 756.450 154.050 757.050 ;
        RECT 139.950 755.400 154.050 756.450 ;
        RECT 139.950 754.950 142.050 755.400 ;
        RECT 151.950 751.950 154.050 755.400 ;
        RECT 157.950 754.950 160.050 757.050 ;
        RECT 166.950 756.450 169.050 757.050 ;
        RECT 175.950 756.450 178.050 757.050 ;
        RECT 166.950 755.400 178.050 756.450 ;
        RECT 166.950 754.950 169.050 755.400 ;
        RECT 175.950 754.950 178.050 755.400 ;
        RECT 181.950 754.950 184.050 757.050 ;
        RECT 187.950 756.450 190.050 757.050 ;
        RECT 199.950 756.450 202.050 757.050 ;
        RECT 187.950 755.400 202.050 756.450 ;
        RECT 187.950 754.950 190.050 755.400 ;
        RECT 199.950 754.950 202.050 755.400 ;
        RECT 211.950 756.450 214.050 757.050 ;
        RECT 223.950 756.450 226.050 757.050 ;
        RECT 211.950 755.400 226.050 756.450 ;
        RECT 211.950 754.950 214.050 755.400 ;
        RECT 223.950 754.950 226.050 755.400 ;
        RECT 229.950 754.950 232.050 757.050 ;
        RECT 235.950 756.450 238.050 757.050 ;
        RECT 244.950 756.450 247.050 757.050 ;
        RECT 235.950 755.400 247.050 756.450 ;
        RECT 235.950 754.950 238.050 755.400 ;
        RECT 244.950 754.950 247.050 755.400 ;
        RECT 262.950 754.950 265.050 757.050 ;
        RECT 268.950 754.950 271.050 757.050 ;
        RECT 286.950 754.950 289.050 757.050 ;
        RECT 292.950 756.450 295.050 757.050 ;
        RECT 297.000 756.450 301.050 757.050 ;
        RECT 292.950 755.400 301.050 756.450 ;
        RECT 292.950 754.950 295.050 755.400 ;
        RECT 297.000 754.950 301.050 755.400 ;
        RECT 310.950 754.950 313.050 757.050 ;
        RECT 316.950 754.950 319.050 757.050 ;
        RECT 328.950 756.450 331.050 757.050 ;
        RECT 337.950 756.450 340.050 757.050 ;
        RECT 328.950 755.400 340.050 756.450 ;
        RECT 328.950 754.950 331.050 755.400 ;
        RECT 337.950 754.950 340.050 755.400 ;
        RECT 343.950 751.950 346.050 757.050 ;
        RECT 358.950 751.950 361.050 757.050 ;
        RECT 364.950 754.950 367.050 757.050 ;
        RECT 370.950 756.450 373.050 757.050 ;
        RECT 382.950 756.450 385.050 757.050 ;
        RECT 370.950 755.400 385.050 756.450 ;
        RECT 370.950 754.950 373.050 755.400 ;
        RECT 382.950 754.950 385.050 755.400 ;
        RECT 388.950 754.950 391.050 757.050 ;
        RECT 394.950 756.450 397.050 756.900 ;
        RECT 406.950 756.450 409.050 757.050 ;
        RECT 394.950 755.400 409.050 756.450 ;
        RECT 394.950 754.800 397.050 755.400 ;
        RECT 406.950 754.950 409.050 755.400 ;
        RECT 412.950 754.950 415.050 757.050 ;
        RECT 391.950 751.950 397.050 754.050 ;
        RECT 415.950 753.450 418.050 754.050 ;
        RECT 430.950 753.450 433.050 757.050 ;
        RECT 436.950 754.950 442.050 757.050 ;
        RECT 451.950 754.950 454.050 757.050 ;
        RECT 457.950 754.950 462.900 757.050 ;
        RECT 464.100 756.450 466.200 757.050 ;
        RECT 472.950 756.450 475.050 757.050 ;
        RECT 464.100 755.400 475.050 756.450 ;
        RECT 464.100 754.950 466.200 755.400 ;
        RECT 472.950 754.950 475.050 755.400 ;
        RECT 478.950 754.950 481.050 757.050 ;
        RECT 484.950 756.450 487.050 757.050 ;
        RECT 489.000 756.450 493.050 757.050 ;
        RECT 484.950 755.400 493.050 756.450 ;
        RECT 484.950 754.950 487.050 755.400 ;
        RECT 489.000 754.950 493.050 755.400 ;
        RECT 496.950 756.450 499.050 757.050 ;
        RECT 505.950 756.450 508.050 757.050 ;
        RECT 496.950 755.400 508.050 756.450 ;
        RECT 496.950 754.950 499.050 755.400 ;
        RECT 505.950 754.950 508.050 755.400 ;
        RECT 415.950 752.400 433.050 753.450 ;
        RECT 463.800 753.000 465.900 754.050 ;
        RECT 415.950 751.950 418.050 752.400 ;
        RECT 463.800 751.950 466.050 753.000 ;
        RECT 467.100 751.950 472.050 754.050 ;
        RECT 493.950 751.950 499.050 754.050 ;
        RECT 511.950 751.950 514.050 757.050 ;
        RECT 526.950 754.950 529.050 757.050 ;
        RECT 538.950 756.450 543.000 757.050 ;
        RECT 544.950 756.450 547.050 757.050 ;
        RECT 538.950 755.400 547.050 756.450 ;
        RECT 538.950 754.950 543.000 755.400 ;
        RECT 544.950 754.950 547.050 755.400 ;
        RECT 550.950 754.950 553.050 757.050 ;
        RECT 568.950 754.950 571.050 757.050 ;
        RECT 574.950 754.950 579.900 757.050 ;
        RECT 581.100 756.450 583.200 757.050 ;
        RECT 595.950 756.450 598.050 757.050 ;
        RECT 581.100 755.400 598.050 756.450 ;
        RECT 581.100 754.950 583.200 755.400 ;
        RECT 595.950 754.950 598.050 755.400 ;
        RECT 601.950 756.450 604.050 757.050 ;
        RECT 613.950 756.450 616.050 757.050 ;
        RECT 601.950 755.400 616.050 756.450 ;
        RECT 553.950 753.450 556.050 754.050 ;
        RECT 559.950 753.450 562.050 754.050 ;
        RECT 553.950 752.400 562.050 753.450 ;
        RECT 553.950 751.950 556.050 752.400 ;
        RECT 559.950 751.950 562.050 752.400 ;
        RECT 601.950 751.950 604.050 755.400 ;
        RECT 613.950 754.950 616.050 755.400 ;
        RECT 619.950 756.450 622.050 757.050 ;
        RECT 634.950 756.450 637.050 757.050 ;
        RECT 619.950 755.400 637.050 756.450 ;
        RECT 619.950 754.950 622.050 755.400 ;
        RECT 634.950 754.950 637.050 755.400 ;
        RECT 640.950 754.950 643.050 757.050 ;
        RECT 646.950 754.950 649.050 757.050 ;
        RECT 658.950 755.250 661.050 757.050 ;
        RECT 664.950 755.250 667.050 757.050 ;
        RECT 679.950 754.950 682.050 757.050 ;
        RECT 685.950 754.950 688.050 757.050 ;
        RECT 691.950 754.950 694.050 757.050 ;
        RECT 697.950 756.450 700.050 757.050 ;
        RECT 712.950 756.450 715.050 757.050 ;
        RECT 697.950 755.400 715.050 756.450 ;
        RECT 697.950 754.950 700.050 755.400 ;
        RECT 712.950 754.950 715.050 755.400 ;
        RECT 727.950 754.950 730.050 757.050 ;
        RECT 733.950 754.950 736.050 757.050 ;
        RECT 748.950 754.950 754.050 757.050 ;
        RECT 757.950 756.450 760.050 757.050 ;
        RECT 769.950 756.450 772.050 757.050 ;
        RECT 757.950 755.400 772.050 756.450 ;
        RECT 757.950 754.950 760.050 755.400 ;
        RECT 769.950 754.950 772.050 755.400 ;
        RECT 787.950 754.950 790.050 757.050 ;
        RECT 793.950 756.450 796.050 757.050 ;
        RECT 811.950 756.450 814.050 757.050 ;
        RECT 793.950 755.400 814.050 756.450 ;
        RECT 793.950 754.950 796.050 755.400 ;
        RECT 811.950 754.950 814.050 755.400 ;
        RECT 817.950 756.450 820.050 757.050 ;
        RECT 822.000 756.450 825.900 757.050 ;
        RECT 817.950 755.400 825.900 756.450 ;
        RECT 817.950 754.950 820.050 755.400 ;
        RECT 822.000 754.950 825.900 755.400 ;
        RECT 827.100 756.450 831.000 757.050 ;
        RECT 832.950 756.450 835.050 757.050 ;
        RECT 827.100 755.400 835.050 756.450 ;
        RECT 827.100 754.950 831.000 755.400 ;
        RECT 832.950 754.950 835.050 755.400 ;
        RECT 853.950 754.950 856.050 757.050 ;
        RECT 859.950 756.450 862.050 757.050 ;
        RECT 864.000 756.450 868.050 757.050 ;
        RECT 859.950 755.400 868.050 756.450 ;
        RECT 859.950 754.950 862.050 755.400 ;
        RECT 864.000 754.950 868.050 755.400 ;
        RECT 877.950 754.950 880.050 757.050 ;
        RECT 898.950 755.250 901.050 757.050 ;
        RECT 904.950 755.250 907.050 757.050 ;
        RECT 658.950 753.450 661.050 754.050 ;
        RECT 653.400 752.400 661.050 753.450 ;
        RECT 31.950 750.450 34.050 751.050 ;
        RECT 43.950 750.450 46.050 751.050 ;
        RECT 31.950 749.400 46.050 750.450 ;
        RECT 31.950 748.950 34.050 749.400 ;
        RECT 43.950 748.950 46.050 749.400 ;
        RECT 58.950 750.450 61.050 751.050 ;
        RECT 97.950 750.450 100.050 751.050 ;
        RECT 58.950 749.400 100.050 750.450 ;
        RECT 58.950 748.950 61.050 749.400 ;
        RECT 97.950 748.950 100.050 749.400 ;
        RECT 112.950 750.450 115.050 751.050 ;
        RECT 130.950 750.450 133.050 751.050 ;
        RECT 112.950 749.400 133.050 750.450 ;
        RECT 112.950 748.950 115.050 749.400 ;
        RECT 130.950 748.950 133.050 749.400 ;
        RECT 154.950 750.450 157.050 751.050 ;
        RECT 220.950 750.450 223.050 751.050 ;
        RECT 154.950 749.400 223.050 750.450 ;
        RECT 154.950 748.950 157.050 749.400 ;
        RECT 220.950 748.950 223.050 749.400 ;
        RECT 247.950 750.450 250.050 751.050 ;
        RECT 256.950 750.450 259.050 751.050 ;
        RECT 355.950 750.450 358.050 751.050 ;
        RECT 370.950 750.450 373.050 751.050 ;
        RECT 247.950 749.400 259.050 750.450 ;
        RECT 247.950 748.950 250.050 749.400 ;
        RECT 256.950 748.950 259.050 749.400 ;
        RECT 260.400 749.400 321.450 750.450 ;
        RECT 85.950 747.450 88.050 748.050 ;
        RECT 97.950 747.450 100.050 748.050 ;
        RECT 85.950 746.400 100.050 747.450 ;
        RECT 85.950 745.950 88.050 746.400 ;
        RECT 97.950 745.950 100.050 746.400 ;
        RECT 106.950 747.450 109.050 748.050 ;
        RECT 118.950 747.450 124.050 748.050 ;
        RECT 106.950 746.400 124.050 747.450 ;
        RECT 106.950 745.950 109.050 746.400 ;
        RECT 118.950 745.950 124.050 746.400 ;
        RECT 145.950 747.450 148.050 748.050 ;
        RECT 157.950 747.450 160.050 748.050 ;
        RECT 163.950 747.450 166.050 748.050 ;
        RECT 145.950 746.400 166.050 747.450 ;
        RECT 145.950 745.950 148.050 746.400 ;
        RECT 157.950 745.950 160.050 746.400 ;
        RECT 163.950 745.950 166.050 746.400 ;
        RECT 169.950 747.450 172.050 748.050 ;
        RECT 178.950 747.450 181.050 748.050 ;
        RECT 169.950 746.400 198.450 747.450 ;
        RECT 169.950 745.950 172.050 746.400 ;
        RECT 178.950 745.950 181.050 746.400 ;
        RECT 197.400 745.050 198.450 746.400 ;
        RECT 205.950 745.950 211.050 748.050 ;
        RECT 260.400 747.450 261.450 749.400 ;
        RECT 320.400 748.050 321.450 749.400 ;
        RECT 355.950 749.400 373.050 750.450 ;
        RECT 355.950 748.950 358.050 749.400 ;
        RECT 370.950 748.950 373.050 749.400 ;
        RECT 376.950 750.450 379.050 751.050 ;
        RECT 463.950 750.450 466.050 751.950 ;
        RECT 376.950 750.000 466.050 750.450 ;
        RECT 478.950 750.450 481.050 751.050 ;
        RECT 484.950 750.450 487.050 751.050 ;
        RECT 376.950 749.400 465.450 750.000 ;
        RECT 478.950 749.400 487.050 750.450 ;
        RECT 376.950 748.950 379.050 749.400 ;
        RECT 478.950 748.950 481.050 749.400 ;
        RECT 484.950 748.950 487.050 749.400 ;
        RECT 490.950 750.450 493.050 751.050 ;
        RECT 538.950 750.450 541.050 751.050 ;
        RECT 490.950 749.400 541.050 750.450 ;
        RECT 490.950 748.950 493.050 749.400 ;
        RECT 538.950 748.950 541.050 749.400 ;
        RECT 544.950 750.450 547.050 751.050 ;
        RECT 568.950 750.450 571.050 751.050 ;
        RECT 544.950 749.400 571.050 750.450 ;
        RECT 544.950 748.950 547.050 749.400 ;
        RECT 568.950 748.950 571.050 749.400 ;
        RECT 587.100 750.450 589.200 751.050 ;
        RECT 616.950 750.450 619.050 751.050 ;
        RECT 587.100 749.400 619.050 750.450 ;
        RECT 587.100 748.950 589.200 749.400 ;
        RECT 616.950 748.950 619.050 749.400 ;
        RECT 622.950 750.450 625.050 751.050 ;
        RECT 643.800 750.450 645.900 751.050 ;
        RECT 622.950 749.400 645.900 750.450 ;
        RECT 622.950 748.950 625.050 749.400 ;
        RECT 643.800 748.950 645.900 749.400 ;
        RECT 647.100 750.450 649.200 751.050 ;
        RECT 653.400 750.450 654.450 752.400 ;
        RECT 658.950 751.950 661.050 752.400 ;
        RECT 664.950 751.950 667.050 754.050 ;
        RECT 647.100 749.400 654.450 750.450 ;
        RECT 673.950 750.450 676.050 751.050 ;
        RECT 679.950 750.450 682.050 751.200 ;
        RECT 673.950 749.400 682.050 750.450 ;
        RECT 686.400 751.050 687.450 754.950 ;
        RECT 734.400 753.000 735.450 754.950 ;
        RECT 686.400 749.400 691.050 751.050 ;
        RECT 727.950 750.450 730.050 751.050 ;
        RECT 647.100 748.950 649.200 749.400 ;
        RECT 673.950 748.950 676.050 749.400 ;
        RECT 679.950 749.100 682.050 749.400 ;
        RECT 687.000 748.950 691.050 749.400 ;
        RECT 692.400 749.400 730.050 750.450 ;
        RECT 242.400 746.400 261.450 747.450 ;
        RECT 265.950 747.450 268.050 748.050 ;
        RECT 301.950 747.450 304.050 748.050 ;
        RECT 265.950 746.400 304.050 747.450 ;
        RECT 16.950 744.450 19.050 745.050 ;
        RECT 25.950 744.450 28.050 745.050 ;
        RECT 16.950 743.400 28.050 744.450 ;
        RECT 16.950 742.950 19.050 743.400 ;
        RECT 25.950 742.950 28.050 743.400 ;
        RECT 55.950 744.450 58.050 745.050 ;
        RECT 82.950 744.450 85.050 745.050 ;
        RECT 91.950 744.450 94.050 745.050 ;
        RECT 55.950 743.400 94.050 744.450 ;
        RECT 55.950 742.950 58.050 743.400 ;
        RECT 82.950 742.950 85.050 743.400 ;
        RECT 91.950 742.950 94.050 743.400 ;
        RECT 97.950 744.450 100.050 745.050 ;
        RECT 133.950 744.450 136.050 745.050 ;
        RECT 97.950 743.400 136.050 744.450 ;
        RECT 97.950 742.950 100.050 743.400 ;
        RECT 133.950 742.950 136.050 743.400 ;
        RECT 196.950 744.450 199.050 745.050 ;
        RECT 223.950 744.450 226.050 745.050 ;
        RECT 242.400 744.450 243.450 746.400 ;
        RECT 265.950 745.950 268.050 746.400 ;
        RECT 301.950 745.950 304.050 746.400 ;
        RECT 319.950 747.450 322.050 748.050 ;
        RECT 346.950 747.450 349.050 748.050 ;
        RECT 400.950 747.450 403.050 748.050 ;
        RECT 319.950 746.400 403.050 747.450 ;
        RECT 319.950 745.950 322.050 746.400 ;
        RECT 346.950 745.950 349.050 746.400 ;
        RECT 400.950 745.950 403.050 746.400 ;
        RECT 406.950 747.450 409.050 748.050 ;
        RECT 412.950 747.450 415.050 748.050 ;
        RECT 406.950 746.400 415.050 747.450 ;
        RECT 406.950 745.950 409.050 746.400 ;
        RECT 412.950 745.950 415.050 746.400 ;
        RECT 451.950 747.450 454.050 748.050 ;
        RECT 466.950 747.450 469.050 748.050 ;
        RECT 451.950 746.400 469.050 747.450 ;
        RECT 451.950 745.950 454.050 746.400 ;
        RECT 466.950 745.950 469.050 746.400 ;
        RECT 481.950 747.450 484.050 748.050 ;
        RECT 502.800 747.450 504.900 748.050 ;
        RECT 481.950 746.400 504.900 747.450 ;
        RECT 481.950 745.950 484.050 746.400 ;
        RECT 502.800 745.950 504.900 746.400 ;
        RECT 577.950 747.450 580.050 748.050 ;
        RECT 595.950 747.450 598.050 748.050 ;
        RECT 577.950 746.400 598.050 747.450 ;
        RECT 577.950 745.950 580.050 746.400 ;
        RECT 595.950 745.950 598.050 746.400 ;
        RECT 640.950 747.450 643.050 748.050 ;
        RECT 652.950 747.450 655.050 748.050 ;
        RECT 640.950 746.400 655.050 747.450 ;
        RECT 640.950 745.950 643.050 746.400 ;
        RECT 652.950 745.950 655.050 746.400 ;
        RECT 664.950 747.450 667.050 748.050 ;
        RECT 679.950 747.450 682.050 747.900 ;
        RECT 685.950 747.450 688.050 748.050 ;
        RECT 692.400 747.450 693.450 749.400 ;
        RECT 727.950 748.950 730.050 749.400 ;
        RECT 733.950 748.950 736.050 753.000 ;
        RECT 739.950 750.450 742.050 751.050 ;
        RECT 878.400 750.450 879.450 754.950 ;
        RECT 898.950 751.950 901.050 754.050 ;
        RECT 904.950 751.950 907.050 754.050 ;
        RECT 739.950 749.400 879.450 750.450 ;
        RECT 739.950 748.950 742.050 749.400 ;
        RECT 664.950 746.400 693.450 747.450 ;
        RECT 808.950 747.450 811.050 748.050 ;
        RECT 814.950 747.450 817.050 748.050 ;
        RECT 808.950 746.400 817.050 747.450 ;
        RECT 664.950 745.950 667.050 746.400 ;
        RECT 679.950 745.800 682.050 746.400 ;
        RECT 685.950 745.950 688.050 746.400 ;
        RECT 808.950 745.950 811.050 746.400 ;
        RECT 814.950 745.950 817.050 746.400 ;
        RECT 820.950 747.450 823.050 748.050 ;
        RECT 850.950 747.450 853.050 748.050 ;
        RECT 820.950 746.400 853.050 747.450 ;
        RECT 820.950 745.950 823.050 746.400 ;
        RECT 850.950 745.950 853.050 746.400 ;
        RECT 880.950 747.450 883.050 748.050 ;
        RECT 898.950 747.450 901.050 748.050 ;
        RECT 880.950 746.400 901.050 747.450 ;
        RECT 880.950 745.950 883.050 746.400 ;
        RECT 898.950 745.950 901.050 746.400 ;
        RECT 196.950 743.400 243.450 744.450 ;
        RECT 244.950 744.450 247.050 745.050 ;
        RECT 307.950 744.450 310.050 745.050 ;
        RECT 376.950 744.450 379.050 745.050 ;
        RECT 244.950 743.400 310.050 744.450 ;
        RECT 196.950 742.950 199.050 743.400 ;
        RECT 223.950 742.950 226.050 743.400 ;
        RECT 244.950 742.950 247.050 743.400 ;
        RECT 307.950 742.950 310.050 743.400 ;
        RECT 317.400 743.400 379.050 744.450 ;
        RECT 13.950 741.450 16.050 742.050 ;
        RECT 28.950 741.450 31.050 742.050 ;
        RECT 13.950 740.400 31.050 741.450 ;
        RECT 13.950 739.950 16.050 740.400 ;
        RECT 28.950 739.950 31.050 740.400 ;
        RECT 70.950 741.450 73.050 742.050 ;
        RECT 88.950 741.450 91.050 742.050 ;
        RECT 70.950 740.400 91.050 741.450 ;
        RECT 70.950 739.950 73.050 740.400 ;
        RECT 88.950 739.950 91.050 740.400 ;
        RECT 124.950 741.450 127.050 742.050 ;
        RECT 166.950 741.450 169.050 742.050 ;
        RECT 124.950 740.400 169.050 741.450 ;
        RECT 124.950 739.950 127.050 740.400 ;
        RECT 166.950 739.950 169.050 740.400 ;
        RECT 250.950 741.450 253.050 742.050 ;
        RECT 280.950 741.450 283.050 742.050 ;
        RECT 250.950 740.400 283.050 741.450 ;
        RECT 250.950 739.950 253.050 740.400 ;
        RECT 280.950 739.950 283.050 740.400 ;
        RECT 289.950 741.450 292.050 742.050 ;
        RECT 317.400 741.450 318.450 743.400 ;
        RECT 376.950 742.950 379.050 743.400 ;
        RECT 394.950 744.450 397.050 745.050 ;
        RECT 436.950 744.450 439.050 745.050 ;
        RECT 649.800 744.450 651.900 745.050 ;
        RECT 394.950 743.400 439.050 744.450 ;
        RECT 394.950 742.950 397.050 743.400 ;
        RECT 436.950 742.950 439.050 743.400 ;
        RECT 572.400 743.400 651.900 744.450 ;
        RECT 289.950 740.400 318.450 741.450 ;
        RECT 334.950 741.450 337.050 742.050 ;
        RECT 358.950 741.450 361.050 742.050 ;
        RECT 334.950 740.400 361.050 741.450 ;
        RECT 289.950 739.950 292.050 740.400 ;
        RECT 334.950 739.950 337.050 740.400 ;
        RECT 358.950 739.950 361.050 740.400 ;
        RECT 385.950 741.450 388.050 742.050 ;
        RECT 430.800 741.450 432.900 742.050 ;
        RECT 385.950 740.400 432.900 741.450 ;
        RECT 385.950 739.950 388.050 740.400 ;
        RECT 430.800 739.950 432.900 740.400 ;
        RECT 511.950 741.450 514.050 742.050 ;
        RECT 572.400 741.450 573.450 743.400 ;
        RECT 649.800 742.950 651.900 743.400 ;
        RECT 653.100 744.450 655.200 745.050 ;
        RECT 736.950 744.450 739.050 745.050 ;
        RECT 757.950 744.450 760.050 745.050 ;
        RECT 653.100 743.400 735.450 744.450 ;
        RECT 653.100 742.950 655.200 743.400 ;
        RECT 511.950 740.400 573.450 741.450 ;
        RECT 589.950 741.450 592.050 742.050 ;
        RECT 619.950 741.450 622.050 742.050 ;
        RECT 589.950 740.400 622.050 741.450 ;
        RECT 511.950 739.950 514.050 740.400 ;
        RECT 589.950 739.950 592.050 740.400 ;
        RECT 619.950 739.950 622.050 740.400 ;
        RECT 722.100 741.450 724.200 742.050 ;
        RECT 730.950 741.450 733.050 742.050 ;
        RECT 722.100 740.400 733.050 741.450 ;
        RECT 734.400 741.450 735.450 743.400 ;
        RECT 736.950 743.400 760.050 744.450 ;
        RECT 736.950 742.950 739.050 743.400 ;
        RECT 757.950 742.950 760.050 743.400 ;
        RECT 847.950 744.450 850.050 745.050 ;
        RECT 904.950 744.450 907.050 748.050 ;
        RECT 847.950 744.000 907.050 744.450 ;
        RECT 847.950 743.400 906.450 744.000 ;
        RECT 847.950 742.950 850.050 743.400 ;
        RECT 742.950 741.450 745.050 742.050 ;
        RECT 772.950 741.450 775.050 742.050 ;
        RECT 787.950 741.450 790.050 742.050 ;
        RECT 808.950 741.450 811.050 742.050 ;
        RECT 734.400 740.400 790.050 741.450 ;
        RECT 722.100 739.950 724.200 740.400 ;
        RECT 730.950 739.950 733.050 740.400 ;
        RECT 742.950 739.950 745.050 740.400 ;
        RECT 772.950 739.950 775.050 740.400 ;
        RECT 787.950 739.950 790.050 740.400 ;
        RECT 800.400 740.400 811.050 741.450 ;
        RECT 1.950 738.450 4.050 739.050 ;
        RECT 37.950 738.450 40.050 739.050 ;
        RECT 61.950 738.450 64.050 739.050 ;
        RECT 1.950 737.400 40.050 738.450 ;
        RECT 41.400 738.000 64.050 738.450 ;
        RECT 1.950 736.950 4.050 737.400 ;
        RECT 37.950 736.950 40.050 737.400 ;
        RECT 40.950 737.400 64.050 738.000 ;
        RECT 7.950 735.450 10.050 736.050 ;
        RECT 7.950 734.400 36.450 735.450 ;
        RECT 7.950 733.950 10.050 734.400 ;
        RECT 35.400 730.050 36.450 734.400 ;
        RECT 40.950 733.950 43.050 737.400 ;
        RECT 61.950 736.950 64.050 737.400 ;
        RECT 79.950 738.450 82.050 739.050 ;
        RECT 97.950 738.450 100.050 739.050 ;
        RECT 175.950 738.450 178.050 739.050 ;
        RECT 79.950 737.400 178.050 738.450 ;
        RECT 79.950 736.950 82.050 737.400 ;
        RECT 97.950 736.950 100.050 737.400 ;
        RECT 175.950 736.950 178.050 737.400 ;
        RECT 190.950 738.450 193.050 739.050 ;
        RECT 196.800 738.450 198.900 739.050 ;
        RECT 190.950 737.400 198.900 738.450 ;
        RECT 190.950 736.950 193.050 737.400 ;
        RECT 196.800 736.950 198.900 737.400 ;
        RECT 200.100 738.450 202.200 739.050 ;
        RECT 214.950 738.450 217.050 739.050 ;
        RECT 200.100 737.400 217.050 738.450 ;
        RECT 200.100 736.950 202.200 737.400 ;
        RECT 214.950 736.950 217.050 737.400 ;
        RECT 247.950 738.450 250.050 739.050 ;
        RECT 256.950 738.450 259.050 739.050 ;
        RECT 247.950 737.400 259.050 738.450 ;
        RECT 247.950 736.950 250.050 737.400 ;
        RECT 256.950 736.950 259.050 737.400 ;
        RECT 271.950 738.450 274.050 739.050 ;
        RECT 343.800 738.450 345.900 739.050 ;
        RECT 271.950 737.400 345.900 738.450 ;
        RECT 271.950 736.950 274.050 737.400 ;
        RECT 343.800 736.950 345.900 737.400 ;
        RECT 347.100 738.450 349.200 739.050 ;
        RECT 376.950 738.450 379.050 739.050 ;
        RECT 347.100 737.400 379.050 738.450 ;
        RECT 347.100 736.950 349.200 737.400 ;
        RECT 376.950 736.950 379.050 737.400 ;
        RECT 397.950 738.450 400.050 739.050 ;
        RECT 406.950 738.450 409.050 739.050 ;
        RECT 397.950 737.400 409.050 738.450 ;
        RECT 397.950 736.950 400.050 737.400 ;
        RECT 406.950 736.950 409.050 737.400 ;
        RECT 427.950 738.450 430.050 739.050 ;
        RECT 472.950 738.450 475.050 739.050 ;
        RECT 517.950 738.450 520.050 739.050 ;
        RECT 628.950 738.450 631.050 739.050 ;
        RECT 427.950 737.400 471.450 738.450 ;
        RECT 427.950 736.950 430.050 737.400 ;
        RECT 46.950 735.450 49.050 736.050 ;
        RECT 55.950 735.450 58.050 736.050 ;
        RECT 46.950 734.400 58.050 735.450 ;
        RECT 46.950 733.950 49.050 734.400 ;
        RECT 55.950 733.950 58.050 734.400 ;
        RECT 112.950 735.450 115.050 736.050 ;
        RECT 127.950 735.450 130.050 736.050 ;
        RECT 157.950 735.450 160.050 736.050 ;
        RECT 178.950 735.450 181.050 736.050 ;
        RECT 112.950 734.400 126.450 735.450 ;
        RECT 112.950 733.950 115.050 734.400 ;
        RECT 16.950 727.950 19.050 730.050 ;
        RECT 28.950 727.950 31.050 730.050 ;
        RECT 34.950 727.950 37.050 730.050 ;
        RECT 55.950 727.950 58.050 730.050 ;
        RECT 61.950 727.950 64.050 733.050 ;
        RECT 67.950 732.450 70.050 733.050 ;
        RECT 73.950 732.450 76.050 733.050 ;
        RECT 67.950 731.400 76.050 732.450 ;
        RECT 67.950 730.950 70.050 731.400 ;
        RECT 73.950 730.950 76.050 731.400 ;
        RECT 125.400 730.050 126.450 734.400 ;
        RECT 127.950 734.400 150.450 735.450 ;
        RECT 127.950 733.950 130.050 734.400 ;
        RECT 149.400 730.050 150.450 734.400 ;
        RECT 157.950 734.400 181.050 735.450 ;
        RECT 157.950 733.950 160.050 734.400 ;
        RECT 178.950 733.950 181.050 734.400 ;
        RECT 208.950 735.450 211.050 736.050 ;
        RECT 259.800 735.450 261.900 736.050 ;
        RECT 208.950 734.400 261.900 735.450 ;
        RECT 208.950 733.950 211.050 734.400 ;
        RECT 259.800 733.950 261.900 734.400 ;
        RECT 263.100 735.450 265.200 736.050 ;
        RECT 280.950 735.450 283.050 736.050 ;
        RECT 298.950 735.450 301.050 736.050 ;
        RECT 313.800 735.450 315.900 736.050 ;
        RECT 263.100 734.400 279.450 735.450 ;
        RECT 263.100 733.950 265.200 734.400 ;
        RECT 70.950 729.450 73.050 730.050 ;
        RECT 82.950 729.450 85.050 730.050 ;
        RECT 70.950 728.400 85.050 729.450 ;
        RECT 70.950 727.950 73.050 728.400 ;
        RECT 82.950 727.950 85.050 728.400 ;
        RECT 88.950 729.450 91.050 730.050 ;
        RECT 100.950 729.450 103.050 730.050 ;
        RECT 88.950 728.400 103.050 729.450 ;
        RECT 88.950 727.950 91.050 728.400 ;
        RECT 100.950 727.950 103.050 728.400 ;
        RECT 106.950 727.950 109.050 730.050 ;
        RECT 118.950 727.950 121.050 730.050 ;
        RECT 124.950 727.950 127.050 730.050 ;
        RECT 142.950 727.950 145.050 730.050 ;
        RECT 148.950 727.950 151.050 730.050 ;
        RECT 169.950 727.950 172.050 730.050 ;
        RECT 175.950 727.950 178.050 733.050 ;
        RECT 190.950 730.950 193.050 733.050 ;
        RECT 196.950 730.950 199.050 733.050 ;
        RECT 278.400 730.050 279.450 734.400 ;
        RECT 280.950 734.400 315.900 735.450 ;
        RECT 280.950 733.950 283.050 734.400 ;
        RECT 298.950 733.950 301.050 734.400 ;
        RECT 313.800 733.950 315.900 734.400 ;
        RECT 317.100 735.450 319.200 736.050 ;
        RECT 331.950 735.450 334.050 736.050 ;
        RECT 454.950 735.450 457.050 736.050 ;
        RECT 466.950 735.450 469.050 736.050 ;
        RECT 317.100 734.400 375.450 735.450 ;
        RECT 317.100 733.950 319.200 734.400 ;
        RECT 331.950 733.950 334.050 734.400 ;
        RECT 374.400 732.450 375.450 734.400 ;
        RECT 454.950 734.400 469.050 735.450 ;
        RECT 470.400 735.450 471.450 737.400 ;
        RECT 472.950 737.400 631.050 738.450 ;
        RECT 472.950 736.950 475.050 737.400 ;
        RECT 517.950 736.950 520.050 737.400 ;
        RECT 628.950 736.950 631.050 737.400 ;
        RECT 634.950 738.450 637.050 739.050 ;
        RECT 646.950 738.450 649.050 739.050 ;
        RECT 634.950 737.400 649.050 738.450 ;
        RECT 634.950 736.950 637.050 737.400 ;
        RECT 646.950 736.950 649.050 737.400 ;
        RECT 655.950 738.450 658.050 739.050 ;
        RECT 694.950 738.450 697.050 739.050 ;
        RECT 655.950 737.400 697.050 738.450 ;
        RECT 655.950 736.950 658.050 737.400 ;
        RECT 694.950 736.950 697.050 737.400 ;
        RECT 700.950 738.450 703.050 739.050 ;
        RECT 715.800 738.450 717.900 739.050 ;
        RECT 700.950 737.400 717.900 738.450 ;
        RECT 700.950 736.950 703.050 737.400 ;
        RECT 715.800 736.950 717.900 737.400 ;
        RECT 719.100 738.450 721.200 738.900 ;
        RECT 724.800 738.450 726.900 739.050 ;
        RECT 719.100 737.400 726.900 738.450 ;
        RECT 719.100 736.800 721.200 737.400 ;
        RECT 724.800 736.950 726.900 737.400 ;
        RECT 728.100 738.450 730.200 739.050 ;
        RECT 748.950 738.450 751.050 739.050 ;
        RECT 728.100 737.400 751.050 738.450 ;
        RECT 728.100 736.950 730.200 737.400 ;
        RECT 748.950 736.950 751.050 737.400 ;
        RECT 781.950 738.450 784.050 739.050 ;
        RECT 800.400 738.450 801.450 740.400 ;
        RECT 808.950 739.950 811.050 740.400 ;
        RECT 889.950 741.450 892.050 742.050 ;
        RECT 904.950 741.450 907.050 742.050 ;
        RECT 889.950 740.400 907.050 741.450 ;
        RECT 889.950 739.950 892.050 740.400 ;
        RECT 904.950 739.950 907.050 740.400 ;
        RECT 781.950 737.400 801.450 738.450 ;
        RECT 802.950 738.450 805.050 739.050 ;
        RECT 814.950 738.450 817.050 739.050 ;
        RECT 802.950 737.400 817.050 738.450 ;
        RECT 781.950 736.950 784.050 737.400 ;
        RECT 802.950 736.950 805.050 737.400 ;
        RECT 814.950 736.950 817.050 737.400 ;
        RECT 886.950 738.450 889.050 739.050 ;
        RECT 892.950 738.450 895.050 739.050 ;
        RECT 886.950 737.400 895.050 738.450 ;
        RECT 886.950 736.950 889.050 737.400 ;
        RECT 892.950 736.950 895.050 737.400 ;
        RECT 898.950 738.450 901.050 739.050 ;
        RECT 904.950 738.450 907.050 739.050 ;
        RECT 898.950 737.400 907.050 738.450 ;
        RECT 898.950 736.950 901.050 737.400 ;
        RECT 904.950 736.950 907.050 737.400 ;
        RECT 484.950 735.450 487.050 736.050 ;
        RECT 470.400 734.400 487.050 735.450 ;
        RECT 454.950 733.950 457.050 734.400 ;
        RECT 466.950 733.950 469.050 734.400 ;
        RECT 484.950 733.950 487.050 734.400 ;
        RECT 493.950 735.450 496.050 736.050 ;
        RECT 526.950 735.450 529.050 736.050 ;
        RECT 532.950 735.450 535.050 736.050 ;
        RECT 601.800 735.450 603.900 736.050 ;
        RECT 493.950 734.400 516.450 735.450 ;
        RECT 493.950 733.950 496.050 734.400 ;
        RECT 385.950 732.450 388.050 733.050 ;
        RECT 374.400 731.400 388.050 732.450 ;
        RECT 385.950 730.950 388.050 731.400 ;
        RECT 190.950 727.950 193.050 729.750 ;
        RECT 196.950 727.950 199.050 729.750 ;
        RECT 211.950 727.950 214.050 730.050 ;
        RECT 217.950 729.450 220.050 730.050 ;
        RECT 232.950 729.450 235.050 730.050 ;
        RECT 217.950 728.400 235.050 729.450 ;
        RECT 217.950 727.950 220.050 728.400 ;
        RECT 232.950 727.950 235.050 728.400 ;
        RECT 253.950 727.950 259.050 730.050 ;
        RECT 262.950 727.950 265.050 730.050 ;
        RECT 277.950 727.950 280.050 730.050 ;
        RECT 292.950 729.450 295.050 730.050 ;
        RECT 301.950 729.450 304.050 730.050 ;
        RECT 292.950 728.400 304.050 729.450 ;
        RECT 292.950 727.950 295.050 728.400 ;
        RECT 301.950 727.950 304.050 728.400 ;
        RECT 307.950 727.950 310.050 730.050 ;
        RECT 313.950 729.450 316.050 730.050 ;
        RECT 322.950 729.450 325.050 730.050 ;
        RECT 313.950 728.400 325.050 729.450 ;
        RECT 313.950 727.950 316.050 728.400 ;
        RECT 322.950 727.950 325.050 728.400 ;
        RECT 343.950 727.950 346.050 730.050 ;
        RECT 367.950 727.950 370.050 730.050 ;
        RECT 373.950 729.450 376.050 730.050 ;
        RECT 388.950 729.450 391.050 730.050 ;
        RECT 373.950 728.400 391.050 729.450 ;
        RECT 373.950 727.950 376.050 728.400 ;
        RECT 388.950 727.950 391.050 728.400 ;
        RECT 394.950 727.950 397.050 730.050 ;
        RECT 400.950 729.450 403.050 730.050 ;
        RECT 412.950 729.450 415.050 733.050 ;
        RECT 515.400 730.050 516.450 734.400 ;
        RECT 526.950 734.400 603.900 735.450 ;
        RECT 526.950 733.950 529.050 734.400 ;
        RECT 532.950 733.950 535.050 734.400 ;
        RECT 601.800 733.950 603.900 734.400 ;
        RECT 634.950 735.450 637.050 736.050 ;
        RECT 649.950 735.450 652.050 736.050 ;
        RECT 634.950 734.400 652.050 735.450 ;
        RECT 634.950 733.950 637.050 734.400 ;
        RECT 649.950 733.950 652.050 734.400 ;
        RECT 661.950 735.450 664.050 736.050 ;
        RECT 673.950 735.450 676.050 736.050 ;
        RECT 661.950 734.400 676.050 735.450 ;
        RECT 661.950 733.950 664.050 734.400 ;
        RECT 673.950 733.950 676.050 734.400 ;
        RECT 682.950 735.450 685.050 736.050 ;
        RECT 706.950 735.450 709.050 736.050 ;
        RECT 682.950 734.400 709.050 735.450 ;
        RECT 682.950 733.950 685.050 734.400 ;
        RECT 706.950 733.950 709.050 734.400 ;
        RECT 745.950 735.450 748.050 736.050 ;
        RECT 763.950 735.450 766.050 736.050 ;
        RECT 745.950 734.400 766.050 735.450 ;
        RECT 745.950 733.950 748.050 734.400 ;
        RECT 763.950 733.950 766.050 734.400 ;
        RECT 769.950 735.450 772.050 736.050 ;
        RECT 802.950 735.450 805.050 736.050 ;
        RECT 769.950 734.400 805.050 735.450 ;
        RECT 769.950 733.950 772.050 734.400 ;
        RECT 802.950 733.950 805.050 734.400 ;
        RECT 811.950 735.450 814.050 736.050 ;
        RECT 826.950 735.450 829.050 736.050 ;
        RECT 811.950 734.400 829.050 735.450 ;
        RECT 811.950 733.950 814.050 734.400 ;
        RECT 826.950 733.950 829.050 734.400 ;
        RECT 850.950 735.450 853.050 736.050 ;
        RECT 859.950 735.450 862.050 736.050 ;
        RECT 850.950 734.400 862.050 735.450 ;
        RECT 850.950 733.950 853.050 734.400 ;
        RECT 859.950 733.950 862.050 734.400 ;
        RECT 886.950 735.450 889.050 736.050 ;
        RECT 907.950 735.450 910.050 736.050 ;
        RECT 886.950 734.400 910.050 735.450 ;
        RECT 886.950 733.950 889.050 734.400 ;
        RECT 907.950 733.950 910.050 734.400 ;
        RECT 649.950 732.450 652.050 733.050 ;
        RECT 655.950 732.450 658.050 733.050 ;
        RECT 649.950 731.400 658.050 732.450 ;
        RECT 649.950 730.950 652.050 731.400 ;
        RECT 655.950 730.950 658.050 731.400 ;
        RECT 724.950 730.950 727.050 733.050 ;
        RECT 730.950 730.950 733.050 733.050 ;
        RECT 883.950 732.450 886.050 733.050 ;
        RECT 889.950 732.450 892.050 733.050 ;
        RECT 883.950 731.400 892.050 732.450 ;
        RECT 883.950 730.950 886.050 731.400 ;
        RECT 889.950 730.950 892.050 731.400 ;
        RECT 400.950 728.400 415.050 729.450 ;
        RECT 400.950 727.950 403.050 728.400 ;
        RECT 412.950 727.950 415.050 728.400 ;
        RECT 418.950 729.450 421.050 730.050 ;
        RECT 423.000 729.450 427.050 730.050 ;
        RECT 418.950 728.400 427.050 729.450 ;
        RECT 418.950 727.950 421.050 728.400 ;
        RECT 423.000 727.950 427.050 728.400 ;
        RECT 430.950 727.950 436.050 730.050 ;
        RECT 454.950 727.950 457.050 730.050 ;
        RECT 469.950 727.950 472.050 730.050 ;
        RECT 475.950 727.950 478.050 730.050 ;
        RECT 487.950 729.450 490.050 730.050 ;
        RECT 496.950 729.450 499.050 730.050 ;
        RECT 487.950 728.400 499.050 729.450 ;
        RECT 487.950 727.950 490.050 728.400 ;
        RECT 496.950 727.950 499.050 728.400 ;
        RECT 514.950 727.950 517.050 730.050 ;
        RECT 520.950 729.450 523.050 730.050 ;
        RECT 529.950 729.450 532.050 730.050 ;
        RECT 520.950 728.400 532.050 729.450 ;
        RECT 520.950 727.950 523.050 728.400 ;
        RECT 529.950 727.950 532.050 728.400 ;
        RECT 583.950 729.450 586.050 730.050 ;
        RECT 592.950 729.450 595.050 730.050 ;
        RECT 583.950 728.400 595.050 729.450 ;
        RECT 583.950 727.950 586.050 728.400 ;
        RECT 592.950 727.950 595.050 728.400 ;
        RECT 598.950 727.950 601.050 730.050 ;
        RECT 604.950 729.450 609.000 730.050 ;
        RECT 610.950 729.450 613.050 730.050 ;
        RECT 604.950 728.400 613.050 729.450 ;
        RECT 604.950 727.950 609.000 728.400 ;
        RECT 610.950 727.950 613.050 728.400 ;
        RECT 616.950 729.450 619.050 730.050 ;
        RECT 634.950 729.450 637.050 730.050 ;
        RECT 616.950 728.400 637.050 729.450 ;
        RECT 616.950 727.950 619.050 728.400 ;
        RECT 634.950 727.950 637.050 728.400 ;
        RECT 640.950 729.450 643.050 730.050 ;
        RECT 652.950 729.450 655.050 730.050 ;
        RECT 640.950 728.400 655.050 729.450 ;
        RECT 640.950 727.950 643.050 728.400 ;
        RECT 652.950 727.950 655.050 728.400 ;
        RECT 661.950 727.950 664.050 730.050 ;
        RECT 667.950 727.950 670.050 730.050 ;
        RECT 685.950 729.450 688.050 730.050 ;
        RECT 694.950 729.450 697.050 730.050 ;
        RECT 685.950 728.400 697.050 729.450 ;
        RECT 685.950 727.950 688.050 728.400 ;
        RECT 694.950 727.950 697.050 728.400 ;
        RECT 700.950 727.950 703.050 730.050 ;
        RECT 706.950 727.950 709.050 730.050 ;
        RECT 724.950 727.950 727.050 729.750 ;
        RECT 730.950 727.950 733.050 729.750 ;
        RECT 745.950 727.950 748.050 730.050 ;
        RECT 751.950 729.450 754.050 730.050 ;
        RECT 763.950 729.450 766.050 730.050 ;
        RECT 772.950 729.450 775.050 730.050 ;
        RECT 751.950 728.400 766.050 729.450 ;
        RECT 751.950 727.950 754.050 728.400 ;
        RECT 763.950 727.950 766.050 728.400 ;
        RECT 767.400 728.400 775.050 729.450 ;
        RECT 16.950 724.950 19.050 726.750 ;
        RECT 28.950 724.950 31.050 726.750 ;
        RECT 34.950 724.950 37.050 726.750 ;
        RECT 55.950 724.950 58.050 726.750 ;
        RECT 61.950 724.950 64.050 726.750 ;
        RECT 82.950 724.950 85.050 726.750 ;
        RECT 100.950 724.950 103.050 726.750 ;
        RECT 106.950 724.950 109.050 726.750 ;
        RECT 118.950 724.950 121.050 726.750 ;
        RECT 124.950 724.950 127.050 726.750 ;
        RECT 142.950 724.950 145.050 726.750 ;
        RECT 148.950 724.950 151.050 726.750 ;
        RECT 169.950 724.950 172.050 726.750 ;
        RECT 175.950 724.950 178.050 726.750 ;
        RECT 193.950 725.250 196.050 727.050 ;
        RECT 211.950 724.950 214.050 726.750 ;
        RECT 232.950 724.950 235.050 726.750 ;
        RECT 256.950 724.950 259.050 726.750 ;
        RECT 262.950 724.950 265.050 726.750 ;
        RECT 277.950 724.950 280.050 726.750 ;
        RECT 301.950 724.950 304.050 726.750 ;
        RECT 307.950 724.950 310.050 726.750 ;
        RECT 322.950 724.950 325.050 726.750 ;
        RECT 328.950 724.950 334.050 727.050 ;
        RECT 343.950 724.950 346.050 726.750 ;
        RECT 361.950 725.250 364.050 727.050 ;
        RECT 371.250 726.750 373.050 727.050 ;
        RECT 367.950 725.250 370.050 726.750 ;
        RECT 370.950 725.250 373.050 726.750 ;
        RECT 367.950 724.950 369.750 725.250 ;
        RECT 376.950 724.950 382.050 727.050 ;
        RECT 541.950 726.750 543.750 727.050 ;
        RECT 388.950 724.950 391.050 726.750 ;
        RECT 394.950 724.950 397.050 726.750 ;
        RECT 412.950 724.950 415.050 726.750 ;
        RECT 418.950 724.950 421.050 726.750 ;
        RECT 433.950 724.950 436.050 726.750 ;
        RECT 454.950 724.950 457.050 726.750 ;
        RECT 469.950 724.950 472.050 726.750 ;
        RECT 475.950 724.950 478.050 726.750 ;
        RECT 496.950 724.950 499.050 726.750 ;
        RECT 514.950 724.950 517.050 726.750 ;
        RECT 520.950 724.950 523.050 726.750 ;
        RECT 541.950 725.250 544.050 726.750 ;
        RECT 544.950 725.250 547.050 726.750 ;
        RECT 550.950 725.250 553.050 727.050 ;
        RECT 565.950 726.750 567.750 727.050 ;
        RECT 565.950 725.250 568.050 726.750 ;
        RECT 568.950 725.250 571.050 726.750 ;
        RECT 574.950 725.250 577.050 727.050 ;
        RECT 545.250 724.950 547.050 725.250 ;
        RECT 569.250 724.950 571.050 725.250 ;
        RECT 592.950 724.950 595.050 726.750 ;
        RECT 598.950 724.950 601.050 726.750 ;
        RECT 610.950 724.950 613.050 726.750 ;
        RECT 616.950 724.950 619.050 726.750 ;
        RECT 640.950 724.950 643.050 726.750 ;
        RECT 661.950 724.950 664.050 726.750 ;
        RECT 667.950 724.950 670.050 726.750 ;
        RECT 685.950 724.950 688.050 726.750 ;
        RECT 700.950 724.950 703.050 726.750 ;
        RECT 706.950 724.950 709.050 726.750 ;
        RECT 727.950 725.250 730.050 727.050 ;
        RECT 745.950 724.950 748.050 726.750 ;
        RECT 751.950 724.950 754.050 726.750 ;
        RECT 757.950 726.450 760.050 727.050 ;
        RECT 767.400 726.450 768.450 728.400 ;
        RECT 772.950 727.950 775.050 728.400 ;
        RECT 793.950 727.950 796.050 730.050 ;
        RECT 814.950 727.950 817.050 730.050 ;
        RECT 829.950 727.950 832.050 730.050 ;
        RECT 835.950 729.450 838.050 730.050 ;
        RECT 847.950 729.450 850.050 730.050 ;
        RECT 835.950 728.400 850.050 729.450 ;
        RECT 835.950 727.950 838.050 728.400 ;
        RECT 847.950 727.950 850.050 728.400 ;
        RECT 868.950 727.950 874.050 730.050 ;
        RECT 757.950 725.400 768.450 726.450 ;
        RECT 757.950 724.950 760.050 725.400 ;
        RECT 772.950 724.950 775.050 726.750 ;
        RECT 793.950 724.950 796.050 726.750 ;
        RECT 814.950 724.950 817.050 726.750 ;
        RECT 829.950 724.950 832.050 726.750 ;
        RECT 847.950 724.950 850.050 726.750 ;
        RECT 853.950 725.250 856.050 727.050 ;
        RECT 871.950 724.950 874.050 726.750 ;
        RECT 886.950 724.950 889.050 730.050 ;
        RECT 892.950 727.950 895.050 730.050 ;
        RECT 898.950 727.950 901.050 730.050 ;
        RECT 892.950 724.950 895.050 726.750 ;
        RECT 898.950 724.950 901.050 726.750 ;
        RECT 13.950 722.250 16.050 724.050 ;
        RECT 31.950 722.250 34.050 724.050 ;
        RECT 37.950 722.250 40.050 724.050 ;
        RECT 52.950 722.250 55.050 724.050 ;
        RECT 58.950 722.250 61.050 724.050 ;
        RECT 79.950 722.250 82.050 724.050 ;
        RECT 97.950 722.250 100.050 724.050 ;
        RECT 103.950 722.250 106.050 724.050 ;
        RECT 121.950 722.250 124.050 724.050 ;
        RECT 127.950 722.250 130.050 724.050 ;
        RECT 145.950 722.250 148.050 724.050 ;
        RECT 151.950 722.250 154.050 724.050 ;
        RECT 166.950 722.250 169.050 724.050 ;
        RECT 172.950 722.250 175.050 724.050 ;
        RECT 181.950 723.450 184.050 724.050 ;
        RECT 193.950 723.450 196.050 724.050 ;
        RECT 181.950 722.400 196.050 723.450 ;
        RECT 181.950 721.950 184.050 722.400 ;
        RECT 193.950 721.950 196.050 722.400 ;
        RECT 214.950 722.250 217.050 724.050 ;
        RECT 229.950 722.250 232.050 724.050 ;
        RECT 235.950 722.250 238.050 724.050 ;
        RECT 253.950 722.250 256.050 724.050 ;
        RECT 259.950 722.250 262.050 724.050 ;
        RECT 274.950 722.250 277.050 724.050 ;
        RECT 280.950 722.250 283.050 724.050 ;
        RECT 298.950 722.250 301.050 724.050 ;
        RECT 304.950 722.250 307.050 724.050 ;
        RECT 319.950 722.250 322.050 724.050 ;
        RECT 325.950 722.250 328.050 724.050 ;
        RECT 340.950 722.250 343.050 724.050 ;
        RECT 346.950 722.250 349.050 724.050 ;
        RECT 361.950 721.950 364.050 724.050 ;
        RECT 370.950 721.950 373.050 724.050 ;
        RECT 385.950 722.250 388.050 724.050 ;
        RECT 391.950 722.250 394.050 724.050 ;
        RECT 409.950 722.250 412.050 724.050 ;
        RECT 415.950 722.250 418.050 724.050 ;
        RECT 436.950 722.250 439.050 724.050 ;
        RECT 451.950 722.250 454.050 724.050 ;
        RECT 472.950 722.250 475.050 724.050 ;
        RECT 478.950 722.250 481.050 724.050 ;
        RECT 493.950 722.250 496.050 724.050 ;
        RECT 499.950 722.250 502.050 724.050 ;
        RECT 517.950 722.250 520.050 724.050 ;
        RECT 523.950 722.250 526.050 724.050 ;
        RECT 529.950 723.450 532.050 724.050 ;
        RECT 541.950 723.450 544.050 724.050 ;
        RECT 529.950 722.400 544.050 723.450 ;
        RECT 529.950 721.950 532.050 722.400 ;
        RECT 541.950 721.950 544.050 722.400 ;
        RECT 550.950 721.950 556.050 724.050 ;
        RECT 565.950 721.950 568.050 724.050 ;
        RECT 574.950 723.450 577.050 724.050 ;
        RECT 583.950 723.450 586.050 724.050 ;
        RECT 574.950 722.400 586.050 723.450 ;
        RECT 574.950 721.950 577.050 722.400 ;
        RECT 583.950 721.950 586.050 722.400 ;
        RECT 589.950 722.250 592.050 724.050 ;
        RECT 595.950 722.250 598.050 724.050 ;
        RECT 613.950 722.250 616.050 724.050 ;
        RECT 619.950 722.250 622.050 724.050 ;
        RECT 637.950 722.250 640.050 724.050 ;
        RECT 643.950 722.250 646.050 724.050 ;
        RECT 658.950 722.250 661.050 724.050 ;
        RECT 664.950 722.250 667.050 724.050 ;
        RECT 682.950 722.250 685.050 724.050 ;
        RECT 688.950 722.250 691.050 724.050 ;
        RECT 703.950 722.250 706.050 724.050 ;
        RECT 709.950 722.250 712.050 724.050 ;
        RECT 715.950 723.450 718.050 724.050 ;
        RECT 727.950 723.450 730.050 724.050 ;
        RECT 715.950 722.400 730.050 723.450 ;
        RECT 715.950 721.950 718.050 722.400 ;
        RECT 727.950 721.950 730.050 722.400 ;
        RECT 748.950 722.250 751.050 724.050 ;
        RECT 754.950 722.250 757.050 724.050 ;
        RECT 769.950 722.250 772.050 724.050 ;
        RECT 775.950 722.250 778.050 724.050 ;
        RECT 790.950 722.250 793.050 724.050 ;
        RECT 796.950 722.250 799.050 724.050 ;
        RECT 817.950 722.250 820.050 724.050 ;
        RECT 832.950 722.250 835.050 724.050 ;
        RECT 868.950 722.250 871.050 724.050 ;
        RECT 874.950 722.250 877.050 724.050 ;
        RECT 889.950 722.250 892.050 724.050 ;
        RECT 895.950 722.250 898.050 724.050 ;
        RECT 901.950 721.950 906.900 724.050 ;
        RECT 13.950 718.950 16.050 721.050 ;
        RECT 31.950 718.950 34.050 721.050 ;
        RECT 37.950 718.950 40.050 721.050 ;
        RECT 52.950 718.950 55.050 721.050 ;
        RECT 58.950 718.950 61.050 721.050 ;
        RECT 64.950 720.450 67.050 721.050 ;
        RECT 79.950 720.450 82.050 721.050 ;
        RECT 64.950 719.400 82.050 720.450 ;
        RECT 64.950 718.950 67.050 719.400 ;
        RECT 79.950 718.950 82.050 719.400 ;
        RECT 97.950 718.950 100.050 721.050 ;
        RECT 103.950 718.950 106.050 721.050 ;
        RECT 14.400 714.450 15.450 718.950 ;
        RECT 106.950 717.450 109.050 718.050 ;
        RECT 121.950 717.450 124.050 721.050 ;
        RECT 127.950 718.950 130.050 721.050 ;
        RECT 145.950 718.950 148.050 721.050 ;
        RECT 151.950 718.950 154.050 721.050 ;
        RECT 166.950 718.950 169.050 721.050 ;
        RECT 172.950 718.950 175.050 721.050 ;
        RECT 214.950 720.450 217.050 721.050 ;
        RECT 200.400 719.400 217.050 720.450 ;
        RECT 106.950 716.400 124.050 717.450 ;
        RECT 187.950 717.450 190.050 718.050 ;
        RECT 200.400 717.450 201.450 719.400 ;
        RECT 214.950 718.950 217.050 719.400 ;
        RECT 229.950 718.950 232.050 721.050 ;
        RECT 253.950 718.950 256.050 721.050 ;
        RECT 259.950 718.950 262.050 721.050 ;
        RECT 274.950 718.950 277.050 721.050 ;
        RECT 298.950 718.950 301.050 721.050 ;
        RECT 304.950 718.950 307.050 721.050 ;
        RECT 319.950 718.950 322.050 721.050 ;
        RECT 340.950 718.950 343.050 721.050 ;
        RECT 346.950 720.450 349.050 721.050 ;
        RECT 355.950 720.450 358.050 721.050 ;
        RECT 346.950 719.400 358.050 720.450 ;
        RECT 346.950 718.950 349.050 719.400 ;
        RECT 355.950 718.950 358.050 719.400 ;
        RECT 385.950 718.950 388.050 721.050 ;
        RECT 391.950 718.950 394.050 721.050 ;
        RECT 397.950 720.450 400.050 721.050 ;
        RECT 409.950 720.450 412.050 721.050 ;
        RECT 397.950 719.400 412.050 720.450 ;
        RECT 397.950 718.950 400.050 719.400 ;
        RECT 409.950 718.950 412.050 719.400 ;
        RECT 415.950 718.950 418.050 721.050 ;
        RECT 421.950 720.450 424.050 721.050 ;
        RECT 436.950 720.450 439.050 721.050 ;
        RECT 421.950 719.400 439.050 720.450 ;
        RECT 421.950 718.950 424.050 719.400 ;
        RECT 436.950 718.950 439.050 719.400 ;
        RECT 451.950 718.950 454.050 721.050 ;
        RECT 472.950 718.950 475.050 721.050 ;
        RECT 478.950 718.950 481.050 721.050 ;
        RECT 493.950 718.950 496.050 721.050 ;
        RECT 499.950 718.950 502.050 721.050 ;
        RECT 517.950 718.950 520.050 721.050 ;
        RECT 523.950 718.950 526.050 721.050 ;
        RECT 187.950 716.400 201.450 717.450 ;
        RECT 106.950 715.950 109.050 716.400 ;
        RECT 187.950 715.950 190.050 716.400 ;
        RECT 244.950 715.950 250.050 718.050 ;
        RECT 352.950 717.450 355.050 718.050 ;
        RECT 361.950 717.450 364.050 718.050 ;
        RECT 352.950 716.400 364.050 717.450 ;
        RECT 352.950 715.950 355.050 716.400 ;
        RECT 361.950 715.950 364.050 716.400 ;
        RECT 367.950 717.450 370.050 718.050 ;
        RECT 373.950 717.450 376.050 718.050 ;
        RECT 566.400 717.450 567.450 721.950 ;
        RECT 589.950 718.950 592.050 721.050 ;
        RECT 595.950 720.450 598.050 721.050 ;
        RECT 607.950 720.450 610.050 721.050 ;
        RECT 595.950 719.400 610.050 720.450 ;
        RECT 595.950 718.950 598.050 719.400 ;
        RECT 607.950 718.950 610.050 719.400 ;
        RECT 613.950 718.950 616.050 721.050 ;
        RECT 619.950 718.950 622.050 721.050 ;
        RECT 637.950 718.950 640.050 721.050 ;
        RECT 643.950 718.950 646.050 721.050 ;
        RECT 652.950 720.450 657.000 721.050 ;
        RECT 658.950 720.450 661.050 721.050 ;
        RECT 652.950 719.400 661.050 720.450 ;
        RECT 652.950 718.950 657.000 719.400 ;
        RECT 658.950 718.950 661.050 719.400 ;
        RECT 664.950 718.950 667.050 721.050 ;
        RECT 682.950 718.950 685.050 721.050 ;
        RECT 688.950 720.450 691.050 721.050 ;
        RECT 697.950 720.450 700.050 721.050 ;
        RECT 688.950 719.400 700.050 720.450 ;
        RECT 688.950 718.950 691.050 719.400 ;
        RECT 697.950 718.950 700.050 719.400 ;
        RECT 703.950 718.950 706.050 721.050 ;
        RECT 709.950 718.950 712.050 721.050 ;
        RECT 748.950 718.950 751.050 721.050 ;
        RECT 754.950 718.950 757.050 721.050 ;
        RECT 760.950 720.450 763.050 721.050 ;
        RECT 769.950 720.450 772.050 721.050 ;
        RECT 760.950 719.400 772.050 720.450 ;
        RECT 760.950 718.950 763.050 719.400 ;
        RECT 769.950 718.950 772.050 719.400 ;
        RECT 790.950 718.950 793.050 721.050 ;
        RECT 796.950 718.950 799.050 721.050 ;
        RECT 817.950 718.950 820.050 721.050 ;
        RECT 829.950 720.450 835.050 721.050 ;
        RECT 844.950 720.450 847.050 721.050 ;
        RECT 829.950 719.400 847.050 720.450 ;
        RECT 829.950 718.950 835.050 719.400 ;
        RECT 844.950 718.950 847.050 719.400 ;
        RECT 868.950 718.950 871.050 721.050 ;
        RECT 874.950 718.950 877.050 721.050 ;
        RECT 889.950 718.950 892.050 721.050 ;
        RECT 895.950 718.950 898.050 721.050 ;
        RECT 367.950 716.400 376.050 717.450 ;
        RECT 367.950 715.950 370.050 716.400 ;
        RECT 373.950 715.950 376.050 716.400 ;
        RECT 530.400 716.400 567.450 717.450 ;
        RECT 715.950 717.450 718.050 718.050 ;
        RECT 739.950 717.450 742.050 718.050 ;
        RECT 715.950 716.400 742.050 717.450 ;
        RECT 31.950 714.450 34.050 715.050 ;
        RECT 14.400 713.400 34.050 714.450 ;
        RECT 31.950 712.950 34.050 713.400 ;
        RECT 40.950 714.450 43.050 715.050 ;
        RECT 52.950 714.450 55.050 715.050 ;
        RECT 40.950 713.400 55.050 714.450 ;
        RECT 40.950 712.950 43.050 713.400 ;
        RECT 52.950 712.950 55.050 713.400 ;
        RECT 64.950 714.450 67.050 715.050 ;
        RECT 229.950 714.450 232.050 715.050 ;
        RECT 271.800 714.450 273.900 715.050 ;
        RECT 64.950 713.400 213.450 714.450 ;
        RECT 64.950 712.950 67.050 713.400 ;
        RECT 34.950 711.450 37.050 712.050 ;
        RECT 46.950 711.450 49.050 712.050 ;
        RECT 88.950 711.450 91.050 712.050 ;
        RECT 34.950 710.400 91.050 711.450 ;
        RECT 34.950 709.950 37.050 710.400 ;
        RECT 46.950 709.950 49.050 710.400 ;
        RECT 88.950 709.950 91.050 710.400 ;
        RECT 121.950 711.450 124.050 712.050 ;
        RECT 172.950 711.450 175.050 712.050 ;
        RECT 181.800 711.450 183.900 712.050 ;
        RECT 121.950 710.400 183.900 711.450 ;
        RECT 121.950 709.950 124.050 710.400 ;
        RECT 172.950 709.950 175.050 710.400 ;
        RECT 181.800 709.950 183.900 710.400 ;
        RECT 185.100 711.450 187.200 712.050 ;
        RECT 208.950 711.450 211.050 712.050 ;
        RECT 185.100 710.400 211.050 711.450 ;
        RECT 212.400 711.450 213.450 713.400 ;
        RECT 229.950 713.400 273.900 714.450 ;
        RECT 229.950 712.950 232.050 713.400 ;
        RECT 271.800 712.950 273.900 713.400 ;
        RECT 391.950 714.450 394.050 715.050 ;
        RECT 400.950 714.450 403.050 715.050 ;
        RECT 391.950 713.400 403.050 714.450 ;
        RECT 391.950 712.950 394.050 713.400 ;
        RECT 400.950 712.950 403.050 713.400 ;
        RECT 415.950 714.450 418.050 715.050 ;
        RECT 421.950 714.450 424.050 715.050 ;
        RECT 415.950 713.400 424.050 714.450 ;
        RECT 415.950 712.950 418.050 713.400 ;
        RECT 421.950 712.950 424.050 713.400 ;
        RECT 436.950 714.450 439.050 715.050 ;
        RECT 466.950 714.450 469.050 715.050 ;
        RECT 436.950 713.400 469.050 714.450 ;
        RECT 436.950 712.950 439.050 713.400 ;
        RECT 466.950 712.950 469.050 713.400 ;
        RECT 496.950 714.450 499.050 715.050 ;
        RECT 523.950 714.450 526.050 715.200 ;
        RECT 530.400 714.450 531.450 716.400 ;
        RECT 715.950 715.950 718.050 716.400 ;
        RECT 739.950 715.950 742.050 716.400 ;
        RECT 496.950 713.400 531.450 714.450 ;
        RECT 550.950 714.450 553.050 715.050 ;
        RECT 568.950 714.450 571.050 715.050 ;
        RECT 607.950 714.450 610.050 715.050 ;
        RECT 550.950 713.400 610.050 714.450 ;
        RECT 496.950 712.950 499.050 713.400 ;
        RECT 523.950 713.100 526.050 713.400 ;
        RECT 550.950 712.950 553.050 713.400 ;
        RECT 568.950 712.950 571.050 713.400 ;
        RECT 607.950 712.950 610.050 713.400 ;
        RECT 613.950 714.450 616.050 715.050 ;
        RECT 628.950 714.450 631.050 715.050 ;
        RECT 661.950 714.450 664.050 715.050 ;
        RECT 613.950 713.400 664.050 714.450 ;
        RECT 613.950 712.950 616.050 713.400 ;
        RECT 628.950 712.950 631.050 713.400 ;
        RECT 661.950 712.950 664.050 713.400 ;
        RECT 682.950 714.450 685.050 715.050 ;
        RECT 694.950 714.450 697.050 715.050 ;
        RECT 703.950 714.450 706.050 715.050 ;
        RECT 724.950 714.450 727.050 715.050 ;
        RECT 682.950 713.400 727.050 714.450 ;
        RECT 682.950 712.950 685.050 713.400 ;
        RECT 694.950 712.950 697.050 713.400 ;
        RECT 703.950 712.950 706.050 713.400 ;
        RECT 724.950 712.950 727.050 713.400 ;
        RECT 730.950 714.450 733.050 715.200 ;
        RECT 754.950 714.450 757.050 715.050 ;
        RECT 781.800 714.450 783.900 715.050 ;
        RECT 730.950 713.400 757.050 714.450 ;
        RECT 730.950 713.100 733.050 713.400 ;
        RECT 754.950 712.950 757.050 713.400 ;
        RECT 764.400 713.400 783.900 714.450 ;
        RECT 259.950 711.450 262.050 712.050 ;
        RECT 212.400 710.400 262.050 711.450 ;
        RECT 272.400 711.450 273.450 712.950 ;
        RECT 289.950 711.450 292.050 712.050 ;
        RECT 272.400 710.400 292.050 711.450 ;
        RECT 185.100 709.950 187.200 710.400 ;
        RECT 208.950 709.950 211.050 710.400 ;
        RECT 259.950 709.950 262.050 710.400 ;
        RECT 289.950 709.950 292.050 710.400 ;
        RECT 304.950 711.450 307.050 712.050 ;
        RECT 349.950 711.450 352.050 712.050 ;
        RECT 424.950 711.450 427.050 712.050 ;
        RECT 304.950 710.400 352.050 711.450 ;
        RECT 304.950 709.950 307.050 710.400 ;
        RECT 349.950 709.950 352.050 710.400 ;
        RECT 353.400 710.400 427.050 711.450 ;
        RECT 55.950 708.450 58.050 709.050 ;
        RECT 67.950 708.450 70.050 709.050 ;
        RECT 55.950 707.400 70.050 708.450 ;
        RECT 55.950 706.950 58.050 707.400 ;
        RECT 67.950 706.950 70.050 707.400 ;
        RECT 106.950 708.450 109.050 709.050 ;
        RECT 166.950 708.450 169.050 709.050 ;
        RECT 265.950 708.450 268.050 709.050 ;
        RECT 106.950 707.400 169.050 708.450 ;
        RECT 212.400 708.000 268.050 708.450 ;
        RECT 106.950 706.950 109.050 707.400 ;
        RECT 166.950 706.950 169.050 707.400 ;
        RECT 211.950 707.400 268.050 708.000 ;
        RECT 100.950 705.450 103.050 706.050 ;
        RECT 139.950 705.450 142.050 706.050 ;
        RECT 100.950 704.400 142.050 705.450 ;
        RECT 100.950 703.950 103.050 704.400 ;
        RECT 139.950 703.950 142.050 704.400 ;
        RECT 151.950 705.450 154.050 706.050 ;
        RECT 151.950 704.400 195.450 705.450 ;
        RECT 151.950 703.950 154.050 704.400 ;
        RECT 136.950 702.450 139.050 703.050 ;
        RECT 157.950 702.450 160.050 703.050 ;
        RECT 136.950 701.400 160.050 702.450 ;
        RECT 136.950 700.950 139.050 701.400 ;
        RECT 157.950 700.950 160.050 701.400 ;
        RECT 166.950 702.450 169.050 703.050 ;
        RECT 187.950 702.450 190.050 703.050 ;
        RECT 166.950 701.400 190.050 702.450 ;
        RECT 194.400 702.450 195.450 704.400 ;
        RECT 211.950 703.950 214.050 707.400 ;
        RECT 265.950 706.950 268.050 707.400 ;
        RECT 292.950 708.450 295.050 709.050 ;
        RECT 301.950 708.450 304.050 709.050 ;
        RECT 292.950 707.400 304.050 708.450 ;
        RECT 292.950 706.950 295.050 707.400 ;
        RECT 301.950 706.950 304.050 707.400 ;
        RECT 319.950 708.450 322.050 709.050 ;
        RECT 331.950 708.450 334.050 709.050 ;
        RECT 319.950 707.400 334.050 708.450 ;
        RECT 319.950 706.950 322.050 707.400 ;
        RECT 331.950 706.950 334.050 707.400 ;
        RECT 337.950 708.450 340.050 709.050 ;
        RECT 353.400 708.450 354.450 710.400 ;
        RECT 424.950 709.950 427.050 710.400 ;
        RECT 472.950 711.450 475.050 712.200 ;
        RECT 490.950 711.450 493.050 712.050 ;
        RECT 472.950 710.400 493.050 711.450 ;
        RECT 472.950 710.100 475.050 710.400 ;
        RECT 490.950 709.950 493.050 710.400 ;
        RECT 499.950 711.450 502.050 712.050 ;
        RECT 505.950 711.450 508.050 712.050 ;
        RECT 499.950 710.400 508.050 711.450 ;
        RECT 499.950 709.950 502.050 710.400 ;
        RECT 505.950 709.950 508.050 710.400 ;
        RECT 523.950 711.450 526.050 711.900 ;
        RECT 532.950 711.450 535.050 712.050 ;
        RECT 523.950 710.400 535.050 711.450 ;
        RECT 523.950 709.800 526.050 710.400 ;
        RECT 532.950 709.950 535.050 710.400 ;
        RECT 559.950 711.450 562.050 712.050 ;
        RECT 577.950 711.450 580.050 712.050 ;
        RECT 589.950 711.450 592.050 712.050 ;
        RECT 559.950 710.400 592.050 711.450 ;
        RECT 559.950 709.950 562.050 710.400 ;
        RECT 577.950 709.950 580.050 710.400 ;
        RECT 589.950 709.950 592.050 710.400 ;
        RECT 625.950 711.450 628.050 712.050 ;
        RECT 637.950 711.450 640.050 712.050 ;
        RECT 625.950 710.400 640.050 711.450 ;
        RECT 625.950 709.950 628.050 710.400 ;
        RECT 637.950 709.950 640.050 710.400 ;
        RECT 649.950 709.950 655.050 712.050 ;
        RECT 670.950 711.450 673.050 712.050 ;
        RECT 688.950 711.450 691.050 712.050 ;
        RECT 670.950 710.400 691.050 711.450 ;
        RECT 670.950 709.950 673.050 710.400 ;
        RECT 688.950 709.950 691.050 710.400 ;
        RECT 694.950 711.450 697.050 712.050 ;
        RECT 709.950 711.450 712.050 712.050 ;
        RECT 694.950 710.400 712.050 711.450 ;
        RECT 694.950 709.950 697.050 710.400 ;
        RECT 709.950 709.950 712.050 710.400 ;
        RECT 730.950 711.450 733.050 711.900 ;
        RECT 748.950 711.450 751.050 712.050 ;
        RECT 730.950 710.400 751.050 711.450 ;
        RECT 337.950 707.400 354.450 708.450 ;
        RECT 355.950 708.450 358.050 709.050 ;
        RECT 391.950 708.450 394.050 709.050 ;
        RECT 424.950 708.450 427.050 709.050 ;
        RECT 355.950 707.400 427.050 708.450 ;
        RECT 337.950 706.950 340.050 707.400 ;
        RECT 355.950 706.950 358.050 707.400 ;
        RECT 391.950 706.950 394.050 707.400 ;
        RECT 424.950 706.950 427.050 707.400 ;
        RECT 439.950 708.450 442.050 709.050 ;
        RECT 472.950 708.450 475.050 708.900 ;
        RECT 478.950 708.450 481.050 709.050 ;
        RECT 439.950 707.400 481.050 708.450 ;
        RECT 439.950 706.950 442.050 707.400 ;
        RECT 472.950 706.800 475.050 707.400 ;
        RECT 478.950 706.950 481.050 707.400 ;
        RECT 520.950 708.450 523.050 709.050 ;
        RECT 529.950 708.450 532.050 709.050 ;
        RECT 520.950 707.400 532.050 708.450 ;
        RECT 520.950 706.950 523.050 707.400 ;
        RECT 529.950 706.950 532.050 707.400 ;
        RECT 544.950 708.450 547.050 709.050 ;
        RECT 560.400 708.450 561.450 709.950 ;
        RECT 544.950 707.400 561.450 708.450 ;
        RECT 583.950 708.450 586.050 709.050 ;
        RECT 592.800 708.450 594.900 709.050 ;
        RECT 583.950 707.400 594.900 708.450 ;
        RECT 544.950 706.950 547.050 707.400 ;
        RECT 583.950 706.950 586.050 707.400 ;
        RECT 592.800 706.950 594.900 707.400 ;
        RECT 596.100 708.450 598.200 709.050 ;
        RECT 619.800 708.450 621.900 709.050 ;
        RECT 596.100 707.400 621.900 708.450 ;
        RECT 596.100 706.950 598.200 707.400 ;
        RECT 619.800 706.950 621.900 707.400 ;
        RECT 623.100 708.450 625.200 709.050 ;
        RECT 631.950 708.450 634.050 709.050 ;
        RECT 623.100 707.400 634.050 708.450 ;
        RECT 623.100 706.950 625.200 707.400 ;
        RECT 631.950 706.950 634.050 707.400 ;
        RECT 643.950 708.450 646.050 709.050 ;
        RECT 671.400 708.450 672.450 709.950 ;
        RECT 730.950 709.800 733.050 710.400 ;
        RECT 748.950 709.950 751.050 710.400 ;
        RECT 757.950 711.450 760.050 712.050 ;
        RECT 764.400 711.450 765.450 713.400 ;
        RECT 781.800 712.950 783.900 713.400 ;
        RECT 826.950 714.450 829.050 715.050 ;
        RECT 868.950 714.450 871.050 715.050 ;
        RECT 889.950 714.450 892.050 715.050 ;
        RECT 826.950 713.400 892.050 714.450 ;
        RECT 826.950 712.950 829.050 713.400 ;
        RECT 868.950 712.950 871.050 713.400 ;
        RECT 889.950 712.950 892.050 713.400 ;
        RECT 757.950 710.400 765.450 711.450 ;
        RECT 766.950 711.450 769.050 712.050 ;
        RECT 835.950 711.450 838.050 712.050 ;
        RECT 766.950 710.400 838.050 711.450 ;
        RECT 757.950 709.950 760.050 710.400 ;
        RECT 766.950 709.950 769.050 710.400 ;
        RECT 835.950 709.950 838.050 710.400 ;
        RECT 844.950 711.450 847.050 712.050 ;
        RECT 883.950 711.450 886.050 712.050 ;
        RECT 844.950 710.400 886.050 711.450 ;
        RECT 908.100 711.000 910.200 712.050 ;
        RECT 844.950 709.950 847.050 710.400 ;
        RECT 883.950 709.950 886.050 710.400 ;
        RECT 907.950 709.950 910.200 711.000 ;
        RECT 907.950 709.050 910.050 709.950 ;
        RECT 643.950 707.400 672.450 708.450 ;
        RECT 727.950 708.450 730.050 709.050 ;
        RECT 742.950 708.450 745.050 709.050 ;
        RECT 727.950 707.400 745.050 708.450 ;
        RECT 643.950 706.950 646.050 707.400 ;
        RECT 727.950 706.950 730.050 707.400 ;
        RECT 742.950 706.950 745.050 707.400 ;
        RECT 754.950 708.450 757.050 709.050 ;
        RECT 760.800 708.450 762.900 709.050 ;
        RECT 754.950 707.400 762.900 708.450 ;
        RECT 754.950 706.950 757.050 707.400 ;
        RECT 760.800 706.950 762.900 707.400 ;
        RECT 764.100 708.450 766.200 709.050 ;
        RECT 787.950 708.450 790.050 709.050 ;
        RECT 764.100 707.400 790.050 708.450 ;
        RECT 764.100 706.950 766.200 707.400 ;
        RECT 787.950 706.950 790.050 707.400 ;
        RECT 796.950 708.450 799.050 709.050 ;
        RECT 802.950 708.450 805.050 709.050 ;
        RECT 796.950 707.400 805.050 708.450 ;
        RECT 907.950 708.000 910.200 709.050 ;
        RECT 796.950 706.950 799.050 707.400 ;
        RECT 802.950 706.950 805.050 707.400 ;
        RECT 908.100 706.950 910.200 708.000 ;
        RECT 235.950 705.450 238.050 706.050 ;
        RECT 253.950 705.450 256.050 706.050 ;
        RECT 235.950 704.400 256.050 705.450 ;
        RECT 235.950 703.950 238.050 704.400 ;
        RECT 253.950 703.950 256.050 704.400 ;
        RECT 292.950 705.450 295.050 706.050 ;
        RECT 304.950 705.450 307.050 706.050 ;
        RECT 397.950 705.450 400.050 706.050 ;
        RECT 292.950 704.400 307.050 705.450 ;
        RECT 292.950 703.950 295.050 704.400 ;
        RECT 304.950 703.950 307.050 704.400 ;
        RECT 308.400 704.400 400.050 705.450 ;
        RECT 238.950 702.450 241.050 703.050 ;
        RECT 308.400 702.450 309.450 704.400 ;
        RECT 397.950 703.950 400.050 704.400 ;
        RECT 403.950 705.450 406.050 706.050 ;
        RECT 409.800 705.450 411.900 706.050 ;
        RECT 403.950 704.400 411.900 705.450 ;
        RECT 403.950 703.950 406.050 704.400 ;
        RECT 409.800 703.950 411.900 704.400 ;
        RECT 413.100 705.450 415.200 706.050 ;
        RECT 460.950 705.450 463.050 706.050 ;
        RECT 413.100 704.400 463.050 705.450 ;
        RECT 413.100 703.950 415.200 704.400 ;
        RECT 460.950 703.950 463.050 704.400 ;
        RECT 481.950 705.450 484.050 706.050 ;
        RECT 493.950 705.450 496.050 706.050 ;
        RECT 481.950 704.400 496.050 705.450 ;
        RECT 481.950 703.950 484.050 704.400 ;
        RECT 493.950 703.950 496.050 704.400 ;
        RECT 541.950 705.450 544.050 706.050 ;
        RECT 568.950 705.450 571.050 706.050 ;
        RECT 541.950 704.400 571.050 705.450 ;
        RECT 541.950 703.950 544.050 704.400 ;
        RECT 568.950 703.950 571.050 704.400 ;
        RECT 685.950 705.450 688.050 706.050 ;
        RECT 736.800 705.450 738.900 706.200 ;
        RECT 685.950 704.400 738.900 705.450 ;
        RECT 685.950 703.950 688.050 704.400 ;
        RECT 736.800 704.100 738.900 704.400 ;
        RECT 740.100 705.450 742.200 706.050 ;
        RECT 766.950 705.450 769.050 706.050 ;
        RECT 740.100 704.400 769.050 705.450 ;
        RECT 740.100 703.950 742.200 704.400 ;
        RECT 766.950 703.950 769.050 704.400 ;
        RECT 799.950 705.450 802.050 706.050 ;
        RECT 814.950 705.450 817.050 706.050 ;
        RECT 799.950 704.400 817.050 705.450 ;
        RECT 799.950 703.950 802.050 704.400 ;
        RECT 814.950 703.950 817.050 704.400 ;
        RECT 820.950 705.450 823.050 706.050 ;
        RECT 841.950 705.450 844.050 706.050 ;
        RECT 820.950 704.400 844.050 705.450 ;
        RECT 820.950 703.950 823.050 704.400 ;
        RECT 841.950 703.950 844.050 704.400 ;
        RECT 194.400 701.400 241.050 702.450 ;
        RECT 166.950 700.950 169.050 701.400 ;
        RECT 187.950 700.950 190.050 701.400 ;
        RECT 238.950 700.950 241.050 701.400 ;
        RECT 293.400 701.400 309.450 702.450 ;
        RECT 310.950 702.450 313.050 703.050 ;
        RECT 358.800 702.450 360.900 703.050 ;
        RECT 310.950 701.400 360.900 702.450 ;
        RECT 58.950 699.450 61.050 700.050 ;
        RECT 112.950 699.450 115.050 700.050 ;
        RECT 58.950 698.400 115.050 699.450 ;
        RECT 58.950 697.950 61.050 698.400 ;
        RECT 112.950 697.950 115.050 698.400 ;
        RECT 127.950 699.450 130.050 700.050 ;
        RECT 142.950 699.450 145.050 700.050 ;
        RECT 214.950 699.450 217.050 700.050 ;
        RECT 127.950 698.400 217.050 699.450 ;
        RECT 127.950 697.950 130.050 698.400 ;
        RECT 142.950 697.950 145.050 698.400 ;
        RECT 214.950 697.950 217.050 698.400 ;
        RECT 268.950 699.450 271.050 700.050 ;
        RECT 293.400 699.450 294.450 701.400 ;
        RECT 310.950 700.950 313.050 701.400 ;
        RECT 358.800 700.950 360.900 701.400 ;
        RECT 362.100 702.450 364.200 703.200 ;
        RECT 388.950 702.450 391.050 703.050 ;
        RECT 362.100 701.400 391.050 702.450 ;
        RECT 362.100 701.100 364.200 701.400 ;
        RECT 388.950 700.950 391.050 701.400 ;
        RECT 400.950 702.450 403.050 703.050 ;
        RECT 505.950 702.450 508.050 703.050 ;
        RECT 529.950 702.450 532.050 703.050 ;
        RECT 400.950 701.400 532.050 702.450 ;
        RECT 400.950 700.950 403.050 701.400 ;
        RECT 505.950 700.950 508.050 701.400 ;
        RECT 529.950 700.950 532.050 701.400 ;
        RECT 586.950 702.450 589.050 703.050 ;
        RECT 682.950 702.450 685.050 703.050 ;
        RECT 586.950 701.400 685.050 702.450 ;
        RECT 586.950 700.950 589.050 701.400 ;
        RECT 682.950 700.950 685.050 701.400 ;
        RECT 772.950 702.450 775.050 703.050 ;
        RECT 811.950 702.450 814.050 703.050 ;
        RECT 772.950 701.400 814.050 702.450 ;
        RECT 772.950 700.950 775.050 701.400 ;
        RECT 811.950 700.950 814.050 701.400 ;
        RECT 823.950 702.450 826.050 703.050 ;
        RECT 877.950 702.450 880.050 703.050 ;
        RECT 895.950 702.450 898.050 703.050 ;
        RECT 823.950 701.400 898.050 702.450 ;
        RECT 823.950 700.950 826.050 701.400 ;
        RECT 877.950 700.950 880.050 701.400 ;
        RECT 895.950 700.950 898.050 701.400 ;
        RECT 907.950 702.450 910.050 703.050 ;
        RECT 907.950 701.400 915.450 702.450 ;
        RECT 907.950 700.950 910.050 701.400 ;
        RECT 659.100 700.050 661.200 700.200 ;
        RECT 268.950 698.400 294.450 699.450 ;
        RECT 295.950 699.450 298.050 700.050 ;
        RECT 307.950 699.450 310.050 700.050 ;
        RECT 295.950 698.400 310.050 699.450 ;
        RECT 268.950 697.950 271.050 698.400 ;
        RECT 295.950 697.950 298.050 698.400 ;
        RECT 307.950 697.950 310.050 698.400 ;
        RECT 328.950 699.450 331.050 700.050 ;
        RECT 343.800 699.450 345.900 700.050 ;
        RECT 328.950 698.400 345.900 699.450 ;
        RECT 328.950 697.950 331.050 698.400 ;
        RECT 343.800 697.950 345.900 698.400 ;
        RECT 370.950 699.450 373.050 700.050 ;
        RECT 376.950 699.450 379.050 700.050 ;
        RECT 496.950 699.450 499.050 700.050 ;
        RECT 520.800 699.450 522.900 700.050 ;
        RECT 370.950 698.400 379.050 699.450 ;
        RECT 370.950 697.950 373.050 698.400 ;
        RECT 376.950 697.950 379.050 698.400 ;
        RECT 458.400 698.400 499.050 699.450 ;
        RECT 16.950 696.450 19.050 697.050 ;
        RECT 64.950 696.450 67.050 697.050 ;
        RECT 16.950 695.400 67.050 696.450 ;
        RECT 16.950 694.950 19.050 695.400 ;
        RECT 64.950 694.950 67.050 695.400 ;
        RECT 88.950 694.950 93.900 697.050 ;
        RECT 95.100 696.450 97.200 697.050 ;
        RECT 175.800 696.450 177.900 697.050 ;
        RECT 95.100 695.400 177.900 696.450 ;
        RECT 95.100 694.950 97.200 695.400 ;
        RECT 175.800 694.950 177.900 695.400 ;
        RECT 179.100 696.450 181.200 697.050 ;
        RECT 184.950 696.450 187.050 697.050 ;
        RECT 179.100 695.400 187.050 696.450 ;
        RECT 179.100 694.950 181.200 695.400 ;
        RECT 184.950 694.950 187.050 695.400 ;
        RECT 190.950 696.450 193.050 697.050 ;
        RECT 205.950 696.450 208.050 697.050 ;
        RECT 190.950 695.400 208.050 696.450 ;
        RECT 190.950 694.950 193.050 695.400 ;
        RECT 205.950 694.950 208.050 695.400 ;
        RECT 238.950 696.450 241.050 697.050 ;
        RECT 250.950 696.450 253.050 697.050 ;
        RECT 238.950 695.400 253.050 696.450 ;
        RECT 238.950 694.950 241.050 695.400 ;
        RECT 250.950 694.950 253.050 695.400 ;
        RECT 265.950 696.450 268.050 697.050 ;
        RECT 277.950 696.450 280.050 697.050 ;
        RECT 310.950 696.450 313.050 697.050 ;
        RECT 265.950 695.400 313.050 696.450 ;
        RECT 265.950 694.950 268.050 695.400 ;
        RECT 277.950 694.950 280.050 695.400 ;
        RECT 310.950 694.950 313.050 695.400 ;
        RECT 316.950 696.450 319.050 697.050 ;
        RECT 337.800 696.450 339.900 697.050 ;
        RECT 316.950 695.400 339.900 696.450 ;
        RECT 316.950 694.950 319.050 695.400 ;
        RECT 337.800 694.950 339.900 695.400 ;
        RECT 341.100 696.450 343.200 697.050 ;
        RECT 373.950 696.450 376.050 697.050 ;
        RECT 341.100 695.400 376.050 696.450 ;
        RECT 341.100 694.950 343.200 695.400 ;
        RECT 373.950 694.950 376.050 695.400 ;
        RECT 379.950 696.450 382.050 697.050 ;
        RECT 403.800 696.450 405.900 697.050 ;
        RECT 379.950 695.400 405.900 696.450 ;
        RECT 379.950 694.950 382.050 695.400 ;
        RECT 403.800 694.950 405.900 695.400 ;
        RECT 407.100 696.450 412.050 697.050 ;
        RECT 430.950 696.450 433.050 697.050 ;
        RECT 458.400 696.450 459.450 698.400 ;
        RECT 496.950 697.950 499.050 698.400 ;
        RECT 500.400 698.400 522.900 699.450 ;
        RECT 407.100 695.400 429.450 696.450 ;
        RECT 407.100 694.950 412.050 695.400 ;
        RECT 28.950 693.450 31.050 694.050 ;
        RECT 37.950 693.450 40.050 694.050 ;
        RECT 14.400 692.400 40.050 693.450 ;
        RECT 14.400 688.050 15.450 692.400 ;
        RECT 28.950 691.950 31.050 692.400 ;
        RECT 37.950 691.950 40.050 692.400 ;
        RECT 85.950 693.450 88.050 694.050 ;
        RECT 118.950 693.450 121.050 694.050 ;
        RECT 148.950 693.450 151.050 694.050 ;
        RECT 85.950 692.400 151.050 693.450 ;
        RECT 85.950 691.950 88.050 692.400 ;
        RECT 118.950 691.950 121.050 692.400 ;
        RECT 148.950 691.950 151.050 692.400 ;
        RECT 172.950 693.450 175.050 694.050 ;
        RECT 199.950 693.450 202.050 694.050 ;
        RECT 172.950 692.400 202.050 693.450 ;
        RECT 172.950 691.950 175.050 692.400 ;
        RECT 199.950 691.950 202.050 692.400 ;
        RECT 223.950 693.450 226.050 694.050 ;
        RECT 232.950 693.450 235.050 694.050 ;
        RECT 223.950 692.400 235.050 693.450 ;
        RECT 223.950 691.950 226.050 692.400 ;
        RECT 232.950 691.950 235.050 692.400 ;
        RECT 250.950 693.450 253.050 694.050 ;
        RECT 355.950 693.450 358.050 694.050 ;
        RECT 250.950 692.400 358.050 693.450 ;
        RECT 250.950 691.950 253.050 692.400 ;
        RECT 355.950 691.950 358.050 692.400 ;
        RECT 361.950 693.450 364.050 694.050 ;
        RECT 406.800 693.450 408.900 694.050 ;
        RECT 361.950 692.400 408.900 693.450 ;
        RECT 361.950 691.950 364.050 692.400 ;
        RECT 406.800 691.950 408.900 692.400 ;
        RECT 410.100 693.450 412.200 694.050 ;
        RECT 428.400 693.450 429.450 695.400 ;
        RECT 430.950 695.400 459.450 696.450 ;
        RECT 460.950 696.450 463.050 697.050 ;
        RECT 500.400 696.450 501.450 698.400 ;
        RECT 520.800 697.950 522.900 698.400 ;
        RECT 524.100 697.950 529.050 700.050 ;
        RECT 532.950 699.450 535.050 700.050 ;
        RECT 550.950 699.450 556.050 700.050 ;
        RECT 532.950 698.400 556.050 699.450 ;
        RECT 532.950 697.950 535.050 698.400 ;
        RECT 550.950 697.950 556.050 698.400 ;
        RECT 559.950 699.450 562.050 700.050 ;
        RECT 574.950 699.450 577.050 700.050 ;
        RECT 622.950 699.450 625.050 700.050 ;
        RECT 559.950 698.400 625.050 699.450 ;
        RECT 559.950 697.950 562.050 698.400 ;
        RECT 574.950 697.950 577.050 698.400 ;
        RECT 622.950 697.950 625.050 698.400 ;
        RECT 637.950 699.450 640.050 700.050 ;
        RECT 643.950 699.450 646.050 700.050 ;
        RECT 637.950 698.400 646.050 699.450 ;
        RECT 637.950 697.950 640.050 698.400 ;
        RECT 643.950 697.950 646.050 698.400 ;
        RECT 649.950 699.450 652.050 700.050 ;
        RECT 655.800 699.450 657.900 700.050 ;
        RECT 649.950 698.400 657.900 699.450 ;
        RECT 649.950 697.950 652.050 698.400 ;
        RECT 655.800 697.950 657.900 698.400 ;
        RECT 659.100 698.100 664.050 700.050 ;
        RECT 660.000 697.950 664.050 698.100 ;
        RECT 721.950 697.950 727.050 700.050 ;
        RECT 751.950 699.450 754.050 700.050 ;
        RECT 757.950 699.450 760.050 700.050 ;
        RECT 751.950 698.400 760.050 699.450 ;
        RECT 751.950 697.950 754.050 698.400 ;
        RECT 757.950 697.950 760.050 698.400 ;
        RECT 763.950 699.450 766.050 700.050 ;
        RECT 772.950 699.450 775.050 700.050 ;
        RECT 763.950 698.400 775.050 699.450 ;
        RECT 763.950 697.950 766.050 698.400 ;
        RECT 772.950 697.950 775.050 698.400 ;
        RECT 841.950 699.450 844.050 700.050 ;
        RECT 862.950 699.450 865.050 700.050 ;
        RECT 871.950 699.450 874.050 700.050 ;
        RECT 841.950 698.400 874.050 699.450 ;
        RECT 841.950 697.950 844.050 698.400 ;
        RECT 862.950 697.950 865.050 698.400 ;
        RECT 871.950 697.950 874.050 698.400 ;
        RECT 586.950 696.450 589.050 697.050 ;
        RECT 460.950 695.400 501.450 696.450 ;
        RECT 503.400 695.400 589.050 696.450 ;
        RECT 430.950 694.950 433.050 695.400 ;
        RECT 460.950 694.950 463.050 695.400 ;
        RECT 448.950 693.450 451.050 694.050 ;
        RECT 410.100 692.400 426.450 693.450 ;
        RECT 428.400 692.400 451.050 693.450 ;
        RECT 410.100 691.950 412.200 692.400 ;
        RECT 425.400 691.050 426.450 692.400 ;
        RECT 448.950 691.950 451.050 692.400 ;
        RECT 481.950 693.450 484.050 694.050 ;
        RECT 503.400 693.450 504.450 695.400 ;
        RECT 586.950 694.950 589.050 695.400 ;
        RECT 601.950 696.450 604.050 697.050 ;
        RECT 625.950 696.450 628.050 697.050 ;
        RECT 715.950 696.450 718.050 697.050 ;
        RECT 601.950 695.400 628.050 696.450 ;
        RECT 601.950 694.950 604.050 695.400 ;
        RECT 625.950 694.950 628.050 695.400 ;
        RECT 659.400 695.400 718.050 696.450 ;
        RECT 659.400 694.050 660.450 695.400 ;
        RECT 715.950 694.950 718.050 695.400 ;
        RECT 721.950 696.450 724.050 697.050 ;
        RECT 730.950 696.450 733.050 697.050 ;
        RECT 721.950 695.400 733.050 696.450 ;
        RECT 721.950 694.950 724.050 695.400 ;
        RECT 730.950 694.950 733.050 695.400 ;
        RECT 742.950 696.450 745.050 697.050 ;
        RECT 754.950 696.450 757.050 697.050 ;
        RECT 742.950 695.400 757.050 696.450 ;
        RECT 742.950 694.950 745.050 695.400 ;
        RECT 754.950 694.950 757.050 695.400 ;
        RECT 865.950 696.450 868.050 697.050 ;
        RECT 880.950 696.450 883.050 697.050 ;
        RECT 865.950 695.400 883.050 696.450 ;
        RECT 865.950 694.950 868.050 695.400 ;
        RECT 880.950 694.950 883.050 695.400 ;
        RECT 886.950 694.950 889.050 700.050 ;
        RECT 904.950 699.450 907.050 700.050 ;
        RECT 910.950 699.450 913.050 700.050 ;
        RECT 904.950 698.400 913.050 699.450 ;
        RECT 904.950 697.950 907.050 698.400 ;
        RECT 910.950 697.950 913.050 698.400 ;
        RECT 914.400 696.450 915.450 701.400 ;
        RECT 911.400 696.000 915.450 696.450 ;
        RECT 910.950 695.400 915.450 696.000 ;
        RECT 481.950 692.400 504.450 693.450 ;
        RECT 511.950 693.450 514.050 694.050 ;
        RECT 520.950 693.450 523.050 694.050 ;
        RECT 511.950 692.400 523.050 693.450 ;
        RECT 481.950 691.950 484.050 692.400 ;
        RECT 511.950 691.950 514.050 692.400 ;
        RECT 520.950 691.950 523.050 692.400 ;
        RECT 529.950 693.450 532.050 694.050 ;
        RECT 550.950 693.450 553.050 694.050 ;
        RECT 529.950 692.400 553.050 693.450 ;
        RECT 614.100 693.000 616.200 694.050 ;
        RECT 529.950 691.950 532.050 692.400 ;
        RECT 550.950 691.950 553.050 692.400 ;
        RECT 613.950 691.950 616.200 693.000 ;
        RECT 652.950 693.450 655.050 694.050 ;
        RECT 658.800 693.450 660.900 694.050 ;
        RECT 652.950 692.400 660.900 693.450 ;
        RECT 652.950 691.950 655.050 692.400 ;
        RECT 658.800 691.950 660.900 692.400 ;
        RECT 662.100 693.450 664.200 694.050 ;
        RECT 730.950 693.450 733.050 694.050 ;
        RECT 748.950 693.450 751.050 694.050 ;
        RECT 662.100 692.400 751.050 693.450 ;
        RECT 662.100 691.950 664.200 692.400 ;
        RECT 730.950 691.950 733.050 692.400 ;
        RECT 748.950 691.950 751.050 692.400 ;
        RECT 757.950 693.450 760.050 694.050 ;
        RECT 784.950 693.450 787.050 694.050 ;
        RECT 793.950 693.450 796.050 694.050 ;
        RECT 757.950 692.400 780.450 693.450 ;
        RECT 757.950 691.950 760.050 692.400 ;
        RECT 313.950 690.450 316.050 691.050 ;
        RECT 322.950 690.450 325.050 691.050 ;
        RECT 313.950 689.400 325.050 690.450 ;
        RECT 313.950 688.950 316.050 689.400 ;
        RECT 322.950 688.950 325.050 689.400 ;
        RECT 340.950 688.950 346.050 691.050 ;
        RECT 391.950 690.450 396.000 691.050 ;
        RECT 391.950 688.950 397.050 690.450 ;
        RECT 425.400 689.400 430.050 691.050 ;
        RECT 426.000 688.950 430.050 689.400 ;
        RECT 613.950 688.950 616.050 691.950 ;
        RECT 679.950 690.450 682.050 691.050 ;
        RECT 691.950 690.450 694.050 691.050 ;
        RECT 709.950 690.450 712.050 691.050 ;
        RECT 679.950 689.400 712.050 690.450 ;
        RECT 679.950 688.950 682.050 689.400 ;
        RECT 691.950 688.950 694.050 689.400 ;
        RECT 709.950 688.950 712.050 689.400 ;
        RECT 13.950 685.950 16.050 688.050 ;
        RECT 34.950 685.950 37.050 688.050 ;
        RECT 40.950 685.950 43.050 688.050 ;
        RECT 58.950 685.950 61.050 688.050 ;
        RECT 64.950 685.950 67.050 688.050 ;
        RECT 79.950 687.450 82.050 688.050 ;
        RECT 94.950 687.450 97.050 688.050 ;
        RECT 79.950 686.400 97.050 687.450 ;
        RECT 79.950 685.950 82.050 686.400 ;
        RECT 94.950 685.950 97.050 686.400 ;
        RECT 100.950 685.950 103.050 688.050 ;
        RECT 106.950 685.950 109.050 688.050 ;
        RECT 121.950 685.950 124.050 688.050 ;
        RECT 127.950 685.950 130.050 688.050 ;
        RECT 13.950 682.950 16.050 684.750 ;
        RECT 34.950 682.950 37.050 684.750 ;
        RECT 40.950 682.950 43.050 684.750 ;
        RECT 58.950 682.950 61.050 684.750 ;
        RECT 64.950 682.950 67.050 684.750 ;
        RECT 79.950 682.950 82.050 684.750 ;
        RECT 100.950 682.950 103.050 684.750 ;
        RECT 106.950 682.950 109.050 684.750 ;
        RECT 121.950 682.950 124.050 684.750 ;
        RECT 127.950 682.950 130.050 684.750 ;
        RECT 142.950 682.950 145.050 685.050 ;
        RECT 148.950 682.950 151.050 688.050 ;
        RECT 160.950 687.450 163.050 688.050 ;
        RECT 172.950 687.450 175.050 688.050 ;
        RECT 160.950 686.400 175.050 687.450 ;
        RECT 160.950 685.950 163.050 686.400 ;
        RECT 172.950 685.950 175.050 686.400 ;
        RECT 178.950 685.950 181.050 688.050 ;
        RECT 193.950 685.950 196.050 688.050 ;
        RECT 199.950 685.950 202.050 688.050 ;
        RECT 217.950 685.950 220.050 688.050 ;
        RECT 223.950 685.950 226.050 688.050 ;
        RECT 232.950 687.450 237.000 688.050 ;
        RECT 238.950 687.450 241.050 688.050 ;
        RECT 232.950 686.400 241.050 687.450 ;
        RECT 232.950 685.950 237.000 686.400 ;
        RECT 238.950 685.950 241.050 686.400 ;
        RECT 262.950 687.450 265.050 688.050 ;
        RECT 271.950 687.450 274.050 688.050 ;
        RECT 262.950 686.400 274.050 687.450 ;
        RECT 262.950 685.950 265.050 686.400 ;
        RECT 271.950 685.950 274.050 686.400 ;
        RECT 277.950 685.950 280.050 688.050 ;
        RECT 283.950 685.950 286.050 688.050 ;
        RECT 301.950 685.950 304.050 688.050 ;
        RECT 307.950 685.950 310.050 688.050 ;
        RECT 328.950 685.950 331.050 688.050 ;
        RECT 334.950 687.450 337.050 688.050 ;
        RECT 339.000 687.450 343.050 688.050 ;
        RECT 334.950 686.400 343.050 687.450 ;
        RECT 334.950 685.950 337.050 686.400 ;
        RECT 339.000 685.950 343.050 686.400 ;
        RECT 349.950 685.950 352.050 688.050 ;
        RECT 370.950 685.950 373.050 688.050 ;
        RECT 394.950 685.950 397.050 688.950 ;
        RECT 779.400 688.050 780.450 692.400 ;
        RECT 784.950 692.400 796.050 693.450 ;
        RECT 784.950 691.950 787.050 692.400 ;
        RECT 793.950 691.950 796.050 692.400 ;
        RECT 883.950 693.450 886.050 694.050 ;
        RECT 904.950 693.450 907.050 694.050 ;
        RECT 883.950 692.400 907.050 693.450 ;
        RECT 883.950 691.950 886.050 692.400 ;
        RECT 904.950 691.950 907.050 692.400 ;
        RECT 910.950 691.950 913.050 695.400 ;
        RECT 859.950 690.450 862.050 691.050 ;
        RECT 859.950 689.400 877.050 690.450 ;
        RECT 859.950 688.950 862.050 689.400 ;
        RECT 400.950 685.950 403.050 688.050 ;
        RECT 409.950 687.450 412.050 688.050 ;
        RECT 418.950 687.450 421.050 688.050 ;
        RECT 409.950 686.400 421.050 687.450 ;
        RECT 409.950 685.950 412.050 686.400 ;
        RECT 418.950 685.950 421.050 686.400 ;
        RECT 430.950 685.950 433.050 688.050 ;
        RECT 433.950 685.950 436.050 688.050 ;
        RECT 454.950 685.950 457.050 688.050 ;
        RECT 460.950 685.950 463.050 688.050 ;
        RECT 484.950 685.950 487.050 688.050 ;
        RECT 520.950 685.950 523.050 688.050 ;
        RECT 538.950 685.950 541.050 688.050 ;
        RECT 544.950 685.950 547.050 688.050 ;
        RECT 550.950 687.450 555.000 688.050 ;
        RECT 556.950 687.450 559.050 688.050 ;
        RECT 550.950 686.400 559.050 687.450 ;
        RECT 550.950 685.950 555.000 686.400 ;
        RECT 556.950 685.950 559.050 686.400 ;
        RECT 562.950 687.450 565.050 688.050 ;
        RECT 574.950 687.450 577.050 688.050 ;
        RECT 562.950 686.400 577.050 687.450 ;
        RECT 562.950 685.950 565.050 686.400 ;
        RECT 574.950 685.950 577.050 686.400 ;
        RECT 580.950 685.950 583.050 688.050 ;
        RECT 586.950 685.950 589.050 688.050 ;
        RECT 622.950 685.950 625.050 688.050 ;
        RECT 646.950 685.950 649.050 688.050 ;
        RECT 652.950 685.950 655.050 688.050 ;
        RECT 667.950 685.950 670.050 688.050 ;
        RECT 712.950 685.950 715.050 688.050 ;
        RECT 718.950 685.950 721.050 688.050 ;
        RECT 742.950 685.950 745.050 688.050 ;
        RECT 757.950 685.950 760.050 688.050 ;
        RECT 763.950 685.950 766.050 688.050 ;
        RECT 778.950 685.950 781.050 688.050 ;
        RECT 784.950 685.950 787.050 688.050 ;
        RECT 802.950 685.950 805.050 688.050 ;
        RECT 823.950 685.950 826.050 688.050 ;
        RECT 829.950 685.950 832.050 688.050 ;
        RECT 850.950 685.950 853.050 688.050 ;
        RECT 856.950 685.950 859.050 688.050 ;
        RECT 874.950 685.950 877.050 689.400 ;
        RECT 880.950 685.950 883.050 688.050 ;
        RECT 890.100 687.450 892.200 688.050 ;
        RECT 898.950 687.450 901.050 688.050 ;
        RECT 890.100 686.400 901.050 687.450 ;
        RECT 890.100 685.950 892.200 686.400 ;
        RECT 898.950 685.950 901.050 686.400 ;
        RECT 154.950 684.450 157.050 685.050 ;
        RECT 163.950 684.450 166.050 685.050 ;
        RECT 154.950 683.400 166.050 684.450 ;
        RECT 154.950 682.950 157.050 683.400 ;
        RECT 163.950 682.950 166.050 683.400 ;
        RECT 172.950 682.950 175.050 684.750 ;
        RECT 178.950 682.950 181.050 684.750 ;
        RECT 193.950 682.950 196.050 684.750 ;
        RECT 199.950 682.950 202.050 684.750 ;
        RECT 217.950 682.950 220.050 684.750 ;
        RECT 223.950 682.950 226.050 684.750 ;
        RECT 238.950 682.950 241.050 684.750 ;
        RECT 244.950 682.950 247.050 684.750 ;
        RECT 262.950 682.950 265.050 684.750 ;
        RECT 277.950 682.950 280.050 684.750 ;
        RECT 283.950 682.950 286.050 684.750 ;
        RECT 301.950 682.950 304.050 684.750 ;
        RECT 307.950 682.950 310.050 684.750 ;
        RECT 328.950 682.950 331.050 684.750 ;
        RECT 334.950 682.950 337.050 684.750 ;
        RECT 349.950 682.950 352.050 684.750 ;
        RECT 355.950 682.950 358.050 684.750 ;
        RECT 370.950 682.950 373.050 684.750 ;
        RECT 376.950 682.950 379.050 684.750 ;
        RECT 394.950 682.950 397.050 684.750 ;
        RECT 400.950 682.950 403.050 684.750 ;
        RECT 418.950 682.950 421.050 684.750 ;
        RECT 424.950 682.950 430.050 685.050 ;
        RECT 433.950 682.950 436.050 684.750 ;
        RECT 439.950 682.950 442.050 684.750 ;
        RECT 454.950 682.950 457.050 684.750 ;
        RECT 460.950 682.950 463.050 684.750 ;
        RECT 484.950 682.950 487.050 684.750 ;
        RECT 502.950 682.950 505.050 684.750 ;
        RECT 520.950 682.950 523.050 684.750 ;
        RECT 538.950 682.950 541.050 684.750 ;
        RECT 544.950 682.950 547.050 684.750 ;
        RECT 556.950 682.950 559.050 684.750 ;
        RECT 562.950 682.950 565.050 684.750 ;
        RECT 580.950 682.950 583.050 684.750 ;
        RECT 586.950 682.950 589.050 684.750 ;
        RECT 604.950 682.950 607.050 684.750 ;
        RECT 622.950 682.950 625.050 684.750 ;
        RECT 628.950 682.950 631.050 684.750 ;
        RECT 646.950 682.950 649.050 684.750 ;
        RECT 652.950 682.950 655.050 684.750 ;
        RECT 667.950 682.950 670.050 684.750 ;
        RECT 673.950 682.950 676.050 684.750 ;
        RECT 694.950 684.450 697.050 685.050 ;
        RECT 703.950 684.450 706.050 685.050 ;
        RECT 694.950 683.400 706.050 684.450 ;
        RECT 694.950 682.950 697.050 683.400 ;
        RECT 703.950 682.950 706.050 683.400 ;
        RECT 712.950 682.950 715.050 684.750 ;
        RECT 718.950 682.950 721.050 684.750 ;
        RECT 727.950 682.950 733.050 685.050 ;
        RECT 736.950 682.950 739.050 684.750 ;
        RECT 742.950 682.950 745.050 684.750 ;
        RECT 757.950 682.950 760.050 684.750 ;
        RECT 763.950 682.950 766.050 684.750 ;
        RECT 778.950 682.950 781.050 684.750 ;
        RECT 784.950 682.950 787.050 684.750 ;
        RECT 802.950 682.950 805.050 684.750 ;
        RECT 808.950 682.950 811.050 684.750 ;
        RECT 823.950 682.950 826.050 684.750 ;
        RECT 829.950 682.950 832.050 684.750 ;
        RECT 850.950 682.950 853.050 684.750 ;
        RECT 856.950 682.950 859.050 684.750 ;
        RECT 874.950 682.950 877.050 684.750 ;
        RECT 880.950 682.950 883.050 684.750 ;
        RECT 898.950 682.950 901.050 684.750 ;
        RECT 16.950 680.250 19.050 682.050 ;
        RECT 31.950 680.250 34.050 682.050 ;
        RECT 37.950 680.250 40.050 682.050 ;
        RECT 55.950 680.250 58.050 682.050 ;
        RECT 61.950 680.250 64.050 682.050 ;
        RECT 82.950 680.250 85.050 682.050 ;
        RECT 97.950 680.250 100.050 682.050 ;
        RECT 103.950 680.250 106.050 682.050 ;
        RECT 118.950 680.250 121.050 682.050 ;
        RECT 124.950 680.250 127.050 682.050 ;
        RECT 142.950 679.950 145.050 681.750 ;
        RECT 148.950 679.950 151.050 681.750 ;
        RECT 154.950 679.950 157.050 681.750 ;
        RECT 175.950 680.250 178.050 682.050 ;
        RECT 196.950 680.250 199.050 682.050 ;
        RECT 202.950 680.250 205.050 682.050 ;
        RECT 214.950 680.250 217.050 682.050 ;
        RECT 220.950 680.250 223.050 682.050 ;
        RECT 241.950 680.250 244.050 682.050 ;
        RECT 250.950 681.450 253.050 682.050 ;
        RECT 259.950 681.450 262.050 682.050 ;
        RECT 250.950 680.400 262.050 681.450 ;
        RECT 250.950 679.950 253.050 680.400 ;
        RECT 259.950 679.950 262.050 680.400 ;
        RECT 265.950 680.250 268.050 682.050 ;
        RECT 280.950 680.250 283.050 682.050 ;
        RECT 286.950 680.250 289.050 682.050 ;
        RECT 304.950 680.250 307.050 682.050 ;
        RECT 310.950 680.250 313.050 682.050 ;
        RECT 325.950 680.250 328.050 682.050 ;
        RECT 331.950 680.250 334.050 682.050 ;
        RECT 337.950 681.450 340.050 682.050 ;
        RECT 346.950 681.450 349.050 682.050 ;
        RECT 337.950 680.400 349.050 681.450 ;
        RECT 337.950 679.950 340.050 680.400 ;
        RECT 346.950 679.950 349.050 680.400 ;
        RECT 352.950 680.250 355.050 682.050 ;
        RECT 373.950 680.250 376.050 682.050 ;
        RECT 391.950 680.250 394.050 682.050 ;
        RECT 397.950 680.250 400.050 682.050 ;
        RECT 421.950 680.250 424.050 682.050 ;
        RECT 436.950 680.250 439.050 682.050 ;
        RECT 457.950 680.250 460.050 682.050 ;
        RECT 463.950 680.250 466.050 682.050 ;
        RECT 481.950 680.250 484.050 682.050 ;
        RECT 499.950 680.250 502.050 682.050 ;
        RECT 517.950 680.250 520.050 682.050 ;
        RECT 523.950 681.450 526.050 682.050 ;
        RECT 529.950 681.450 532.050 682.050 ;
        RECT 523.950 680.400 532.050 681.450 ;
        RECT 523.950 679.950 526.050 680.400 ;
        RECT 529.950 679.950 532.050 680.400 ;
        RECT 535.950 680.250 538.050 682.050 ;
        RECT 541.950 680.250 544.050 682.050 ;
        RECT 559.950 680.250 562.050 682.050 ;
        RECT 565.950 680.250 568.050 682.050 ;
        RECT 583.950 680.250 586.050 682.050 ;
        RECT 589.950 680.250 592.050 682.050 ;
        RECT 607.950 680.250 610.050 682.050 ;
        RECT 625.950 680.250 628.050 682.050 ;
        RECT 643.950 680.250 646.050 682.050 ;
        RECT 649.950 680.250 652.050 682.050 ;
        RECT 670.950 680.250 673.050 682.050 ;
        RECT 694.950 679.950 697.050 681.750 ;
        RECT 709.950 680.250 712.050 682.050 ;
        RECT 715.950 680.250 718.050 682.050 ;
        RECT 739.950 680.250 742.050 682.050 ;
        RECT 745.950 681.450 748.050 682.050 ;
        RECT 751.950 681.450 754.050 682.050 ;
        RECT 745.950 680.400 754.050 681.450 ;
        RECT 745.950 679.950 748.050 680.400 ;
        RECT 751.950 679.950 754.050 680.400 ;
        RECT 760.950 680.250 763.050 682.050 ;
        RECT 766.950 680.250 769.050 682.050 ;
        RECT 781.950 680.250 784.050 682.050 ;
        RECT 787.950 680.250 790.050 682.050 ;
        RECT 805.950 680.250 808.050 682.050 ;
        RECT 826.950 680.250 829.050 682.050 ;
        RECT 832.950 680.250 835.050 682.050 ;
        RECT 853.950 680.250 856.050 682.050 ;
        RECT 859.950 680.250 862.050 682.050 ;
        RECT 871.950 680.250 874.050 682.050 ;
        RECT 877.950 680.250 880.050 682.050 ;
        RECT 883.950 681.450 886.050 682.050 ;
        RECT 889.950 681.450 892.050 682.050 ;
        RECT 883.950 680.400 892.050 681.450 ;
        RECT 883.950 679.950 886.050 680.400 ;
        RECT 889.950 679.950 892.050 680.400 ;
        RECT 895.950 680.250 898.050 682.050 ;
        RECT 901.950 681.450 904.050 682.050 ;
        RECT 907.950 681.450 910.050 682.050 ;
        RECT 901.950 680.400 910.050 681.450 ;
        RECT 901.950 679.950 904.050 680.400 ;
        RECT 907.950 679.950 910.050 680.400 ;
        RECT 16.950 676.950 19.050 679.050 ;
        RECT 31.950 673.950 34.050 679.050 ;
        RECT 37.950 676.950 40.050 679.050 ;
        RECT 43.950 678.450 46.050 679.050 ;
        RECT 55.950 678.450 58.050 679.050 ;
        RECT 43.950 677.400 58.050 678.450 ;
        RECT 43.950 676.950 46.050 677.400 ;
        RECT 55.950 676.950 58.050 677.400 ;
        RECT 61.950 676.950 64.050 679.050 ;
        RECT 82.950 676.950 85.050 679.050 ;
        RECT 97.950 676.950 100.050 679.050 ;
        RECT 103.950 676.950 106.050 679.050 ;
        RECT 118.950 676.950 121.050 679.050 ;
        RECT 124.950 676.950 127.050 679.050 ;
        RECT 145.950 677.250 148.050 679.050 ;
        RECT 151.950 677.250 154.050 679.050 ;
        RECT 157.950 676.950 163.050 679.050 ;
        RECT 169.950 678.450 174.000 679.050 ;
        RECT 175.950 678.450 178.050 679.050 ;
        RECT 169.950 677.400 178.050 678.450 ;
        RECT 169.950 676.950 174.000 677.400 ;
        RECT 175.950 676.950 178.050 677.400 ;
        RECT 190.950 678.450 195.000 679.050 ;
        RECT 196.950 678.450 199.050 679.050 ;
        RECT 190.950 677.400 199.050 678.450 ;
        RECT 190.950 676.950 195.000 677.400 ;
        RECT 196.950 676.950 199.050 677.400 ;
        RECT 202.950 676.950 205.050 679.050 ;
        RECT 214.950 676.950 217.050 679.050 ;
        RECT 220.950 678.450 223.050 679.050 ;
        RECT 235.950 678.450 238.050 679.050 ;
        RECT 220.950 677.400 238.050 678.450 ;
        RECT 220.950 676.950 223.050 677.400 ;
        RECT 235.950 676.950 238.050 677.400 ;
        RECT 241.950 676.950 244.050 679.050 ;
        RECT 265.950 676.950 268.050 679.050 ;
        RECT 280.950 676.950 283.050 679.050 ;
        RECT 286.950 678.450 289.050 679.050 ;
        RECT 298.950 678.450 301.050 679.050 ;
        RECT 286.950 677.400 301.050 678.450 ;
        RECT 286.950 676.950 289.050 677.400 ;
        RECT 298.950 676.950 301.050 677.400 ;
        RECT 304.950 676.950 307.050 679.050 ;
        RECT 310.950 676.950 313.050 679.050 ;
        RECT 37.950 672.450 40.050 673.050 ;
        RECT 70.950 672.450 73.050 673.050 ;
        RECT 37.950 671.400 73.050 672.450 ;
        RECT 37.950 670.950 40.050 671.400 ;
        RECT 70.950 670.950 73.050 671.400 ;
        RECT 88.950 667.950 91.050 673.050 ;
        RECT 98.400 672.450 99.450 676.950 ;
        RECT 106.950 672.450 109.050 673.050 ;
        RECT 98.400 671.400 109.050 672.450 ;
        RECT 106.950 670.950 109.050 671.400 ;
        RECT 112.950 672.450 115.050 673.050 ;
        RECT 125.400 672.450 126.450 676.950 ;
        RECT 145.950 673.950 148.050 676.050 ;
        RECT 151.950 673.950 154.050 676.050 ;
        RECT 325.950 673.950 328.050 679.050 ;
        RECT 331.950 676.950 334.050 679.050 ;
        RECT 343.950 678.450 346.050 679.050 ;
        RECT 352.950 678.450 355.050 679.050 ;
        RECT 343.950 677.400 355.050 678.450 ;
        RECT 343.950 676.950 346.050 677.400 ;
        RECT 352.950 676.950 355.050 677.400 ;
        RECT 358.950 678.450 361.050 679.050 ;
        RECT 373.950 678.450 376.050 679.050 ;
        RECT 358.950 677.400 376.050 678.450 ;
        RECT 358.950 676.950 361.050 677.400 ;
        RECT 373.950 676.950 376.050 677.400 ;
        RECT 112.950 671.400 126.450 672.450 ;
        RECT 172.950 672.450 175.050 673.050 ;
        RECT 184.950 672.450 187.050 673.050 ;
        RECT 172.950 671.400 187.050 672.450 ;
        RECT 112.950 670.950 115.050 671.400 ;
        RECT 172.950 670.950 175.050 671.400 ;
        RECT 184.950 670.950 187.050 671.400 ;
        RECT 193.950 672.450 196.050 673.050 ;
        RECT 202.950 672.450 205.050 673.050 ;
        RECT 214.950 672.450 217.050 673.050 ;
        RECT 193.950 671.400 217.050 672.450 ;
        RECT 193.950 670.950 196.050 671.400 ;
        RECT 202.950 670.950 205.050 671.400 ;
        RECT 214.950 670.950 217.050 671.400 ;
        RECT 232.950 670.950 238.050 673.050 ;
        RECT 271.950 672.450 274.050 673.050 ;
        RECT 301.950 672.450 304.050 673.050 ;
        RECT 271.950 671.400 304.050 672.450 ;
        RECT 271.950 670.950 274.050 671.400 ;
        RECT 301.950 670.950 304.050 671.400 ;
        RECT 307.950 672.450 310.050 673.050 ;
        RECT 332.400 672.450 333.450 676.950 ;
        RECT 379.950 675.450 382.050 676.050 ;
        RECT 385.950 675.450 388.050 676.050 ;
        RECT 379.950 674.400 388.050 675.450 ;
        RECT 379.950 673.950 382.050 674.400 ;
        RECT 385.950 673.950 388.050 674.400 ;
        RECT 391.950 673.950 394.050 679.050 ;
        RECT 397.950 678.450 400.050 679.050 ;
        RECT 412.950 678.450 415.050 679.050 ;
        RECT 397.950 677.400 415.050 678.450 ;
        RECT 397.950 676.950 400.050 677.400 ;
        RECT 412.950 676.950 415.050 677.400 ;
        RECT 421.950 676.950 424.050 679.050 ;
        RECT 427.950 678.450 430.050 679.200 ;
        RECT 436.950 678.450 439.050 679.050 ;
        RECT 451.950 678.450 454.050 679.200 ;
        RECT 427.950 677.400 454.050 678.450 ;
        RECT 427.950 677.100 430.050 677.400 ;
        RECT 436.950 676.950 439.050 677.400 ;
        RECT 451.950 677.100 454.050 677.400 ;
        RECT 457.950 676.950 460.050 679.050 ;
        RECT 429.000 675.900 433.050 676.050 ;
        RECT 427.950 673.950 433.050 675.900 ;
        RECT 442.950 675.450 445.050 676.050 ;
        RECT 451.950 675.450 454.050 675.900 ;
        RECT 442.950 674.400 454.050 675.450 ;
        RECT 442.950 673.950 445.050 674.400 ;
        RECT 427.950 673.800 430.050 673.950 ;
        RECT 451.950 673.800 454.050 674.400 ;
        RECT 463.950 673.950 466.050 679.050 ;
        RECT 469.950 678.450 472.050 679.050 ;
        RECT 481.950 678.450 484.050 679.050 ;
        RECT 469.950 677.400 484.050 678.450 ;
        RECT 469.950 676.950 472.050 677.400 ;
        RECT 481.950 676.950 484.050 677.400 ;
        RECT 499.950 676.950 502.050 679.050 ;
        RECT 517.950 676.950 520.050 679.050 ;
        RECT 527.100 675.000 529.200 676.050 ;
        RECT 526.950 673.950 529.200 675.000 ;
        RECT 535.950 673.950 538.050 679.050 ;
        RECT 541.950 676.950 544.050 679.050 ;
        RECT 559.950 676.950 562.050 679.050 ;
        RECT 565.950 673.950 568.050 679.050 ;
        RECT 574.950 676.950 580.050 679.050 ;
        RECT 583.950 676.950 586.050 679.050 ;
        RECT 589.950 673.950 592.050 679.050 ;
        RECT 607.950 676.950 610.050 679.050 ;
        RECT 625.950 673.950 628.050 679.050 ;
        RECT 643.950 676.950 646.050 679.050 ;
        RECT 649.950 673.950 652.050 679.050 ;
        RECT 658.950 678.450 661.050 679.200 ;
        RECT 670.950 678.450 673.050 679.050 ;
        RECT 658.950 677.400 673.050 678.450 ;
        RECT 658.950 677.100 661.050 677.400 ;
        RECT 670.950 676.950 673.050 677.400 ;
        RECT 691.950 677.250 694.050 679.050 ;
        RECT 697.950 677.250 700.050 679.050 ;
        RECT 709.950 676.950 712.050 679.050 ;
        RECT 715.950 678.450 718.050 679.050 ;
        RECT 733.950 678.450 736.050 679.050 ;
        RECT 715.950 677.400 736.050 678.450 ;
        RECT 715.950 676.950 718.050 677.400 ;
        RECT 733.950 676.950 736.050 677.400 ;
        RECT 739.950 678.450 742.050 679.050 ;
        RECT 754.950 678.450 757.050 679.050 ;
        RECT 739.950 677.400 757.050 678.450 ;
        RECT 739.950 676.950 742.050 677.400 ;
        RECT 754.950 676.950 757.050 677.400 ;
        RECT 655.950 675.900 660.000 676.050 ;
        RECT 655.950 673.950 661.050 675.900 ;
        RECT 691.950 673.950 694.050 676.050 ;
        RECT 697.950 673.950 700.050 676.050 ;
        RECT 760.950 673.950 763.050 679.050 ;
        RECT 766.950 676.950 769.050 679.050 ;
        RECT 781.950 676.950 784.050 679.050 ;
        RECT 787.950 676.950 790.050 679.050 ;
        RECT 805.950 678.450 808.050 679.050 ;
        RECT 820.950 678.450 823.050 679.050 ;
        RECT 805.950 677.400 823.050 678.450 ;
        RECT 805.950 676.950 808.050 677.400 ;
        RECT 820.950 676.950 823.050 677.400 ;
        RECT 826.950 676.950 829.050 679.050 ;
        RECT 832.950 678.450 835.050 679.050 ;
        RECT 841.950 678.450 844.050 679.050 ;
        RECT 832.950 677.400 844.050 678.450 ;
        RECT 832.950 676.950 835.050 677.400 ;
        RECT 841.950 676.950 844.050 677.400 ;
        RECT 526.950 673.050 529.050 673.950 ;
        RECT 658.950 673.800 661.050 673.950 ;
        RECT 788.400 673.050 789.450 676.950 ;
        RECT 853.950 673.950 856.050 679.050 ;
        RECT 859.950 676.950 862.050 679.050 ;
        RECT 871.950 676.950 874.050 679.050 ;
        RECT 877.950 673.950 880.050 679.050 ;
        RECT 895.950 676.950 898.050 679.050 ;
        RECT 307.950 671.400 333.450 672.450 ;
        RECT 340.950 672.450 343.050 673.050 ;
        RECT 352.950 672.450 355.050 673.050 ;
        RECT 424.950 672.450 427.050 673.050 ;
        RECT 487.950 672.450 490.050 673.050 ;
        RECT 340.950 671.400 355.050 672.450 ;
        RECT 307.950 670.950 310.050 671.400 ;
        RECT 340.950 670.950 343.050 671.400 ;
        RECT 352.950 670.950 355.050 671.400 ;
        RECT 386.400 671.400 420.450 672.450 ;
        RECT 151.950 669.450 154.050 670.050 ;
        RECT 166.950 669.450 169.050 670.050 ;
        RECT 151.950 668.400 183.450 669.450 ;
        RECT 151.950 667.950 154.050 668.400 ;
        RECT 166.950 667.950 169.050 668.400 ;
        RECT 136.950 666.450 139.050 667.050 ;
        RECT 175.950 666.450 178.050 667.050 ;
        RECT 136.950 665.400 178.050 666.450 ;
        RECT 182.400 666.450 183.450 668.400 ;
        RECT 184.950 667.950 190.050 670.050 ;
        RECT 217.950 669.450 220.050 670.050 ;
        RECT 250.950 669.450 253.050 670.050 ;
        RECT 256.950 669.450 259.050 670.050 ;
        RECT 217.950 668.400 259.050 669.450 ;
        RECT 217.950 667.950 220.050 668.400 ;
        RECT 250.950 667.950 253.050 668.400 ;
        RECT 256.950 667.950 259.050 668.400 ;
        RECT 298.950 669.450 301.050 670.050 ;
        RECT 313.800 669.450 315.900 670.050 ;
        RECT 298.950 668.400 315.900 669.450 ;
        RECT 298.950 667.950 301.050 668.400 ;
        RECT 313.800 667.950 315.900 668.400 ;
        RECT 317.100 669.450 319.200 670.050 ;
        RECT 334.950 669.450 337.050 670.050 ;
        RECT 317.100 668.400 337.050 669.450 ;
        RECT 317.100 667.950 319.200 668.400 ;
        RECT 334.950 667.950 337.050 668.400 ;
        RECT 343.950 667.950 349.050 670.050 ;
        RECT 361.950 669.450 364.050 670.050 ;
        RECT 350.400 668.400 364.050 669.450 ;
        RECT 208.950 666.450 211.050 667.050 ;
        RECT 182.400 665.400 211.050 666.450 ;
        RECT 136.950 664.950 139.050 665.400 ;
        RECT 175.950 664.950 178.050 665.400 ;
        RECT 208.950 664.950 211.050 665.400 ;
        RECT 223.950 666.450 226.050 667.050 ;
        RECT 310.950 666.450 313.050 667.050 ;
        RECT 331.950 666.450 334.050 667.050 ;
        RECT 350.400 666.450 351.450 668.400 ;
        RECT 361.950 667.950 364.050 668.400 ;
        RECT 370.950 669.450 373.050 670.050 ;
        RECT 386.400 669.450 387.450 671.400 ;
        RECT 370.950 668.400 387.450 669.450 ;
        RECT 370.950 667.950 373.050 668.400 ;
        RECT 403.950 667.950 409.050 670.050 ;
        RECT 412.950 669.450 417.000 670.050 ;
        RECT 419.400 669.450 420.450 671.400 ;
        RECT 424.950 671.400 490.050 672.450 ;
        RECT 424.950 670.950 427.050 671.400 ;
        RECT 487.950 670.950 490.050 671.400 ;
        RECT 496.950 672.450 499.050 673.050 ;
        RECT 523.800 672.450 525.900 673.050 ;
        RECT 496.950 671.400 525.900 672.450 ;
        RECT 526.950 672.000 529.200 673.050 ;
        RECT 496.950 670.950 499.050 671.400 ;
        RECT 523.800 670.950 525.900 671.400 ;
        RECT 527.100 670.950 529.200 672.000 ;
        RECT 532.950 672.450 535.050 673.050 ;
        RECT 544.950 672.450 547.050 673.050 ;
        RECT 532.950 671.400 547.050 672.450 ;
        RECT 532.950 670.950 535.050 671.400 ;
        RECT 544.950 670.950 547.050 671.400 ;
        RECT 550.950 672.450 553.050 673.050 ;
        RECT 568.950 672.450 571.050 673.050 ;
        RECT 601.950 672.450 604.050 673.050 ;
        RECT 550.950 671.400 604.050 672.450 ;
        RECT 550.950 670.950 553.050 671.400 ;
        RECT 568.950 670.950 571.050 671.400 ;
        RECT 601.950 670.950 604.050 671.400 ;
        RECT 607.950 672.450 610.050 673.050 ;
        RECT 613.950 672.450 616.050 673.050 ;
        RECT 607.950 671.400 616.050 672.450 ;
        RECT 607.950 670.950 610.050 671.400 ;
        RECT 613.950 670.950 616.050 671.400 ;
        RECT 634.950 672.450 637.050 673.050 ;
        RECT 643.800 672.450 645.900 673.050 ;
        RECT 634.950 671.400 645.900 672.450 ;
        RECT 634.950 670.950 637.050 671.400 ;
        RECT 643.800 670.950 645.900 671.400 ;
        RECT 647.100 672.450 649.200 673.050 ;
        RECT 661.950 672.450 664.050 673.050 ;
        RECT 647.100 671.400 664.050 672.450 ;
        RECT 647.100 670.950 649.200 671.400 ;
        RECT 661.950 670.950 664.050 671.400 ;
        RECT 703.950 672.450 706.050 673.050 ;
        RECT 781.950 672.450 784.050 673.050 ;
        RECT 703.950 671.400 784.050 672.450 ;
        RECT 703.950 670.950 706.050 671.400 ;
        RECT 781.950 670.950 784.050 671.400 ;
        RECT 787.950 672.450 790.050 673.050 ;
        RECT 826.950 672.450 829.050 673.050 ;
        RECT 787.950 671.400 829.050 672.450 ;
        RECT 787.950 670.950 790.050 671.400 ;
        RECT 826.950 670.950 829.050 671.400 ;
        RECT 850.950 672.450 853.050 673.050 ;
        RECT 859.800 672.450 861.900 673.050 ;
        RECT 850.950 671.400 861.900 672.450 ;
        RECT 850.950 670.950 853.050 671.400 ;
        RECT 859.800 670.950 861.900 671.400 ;
        RECT 863.100 670.950 868.050 673.050 ;
        RECT 886.950 672.450 889.050 673.050 ;
        RECT 898.950 672.450 901.050 673.050 ;
        RECT 886.950 671.400 901.050 672.450 ;
        RECT 886.950 670.950 889.050 671.400 ;
        RECT 898.950 670.950 901.050 671.400 ;
        RECT 442.950 669.450 445.050 670.050 ;
        RECT 412.950 667.950 417.450 669.450 ;
        RECT 419.400 668.400 445.050 669.450 ;
        RECT 442.950 667.950 445.050 668.400 ;
        RECT 448.950 669.450 451.050 670.050 ;
        RECT 484.950 669.450 487.050 670.050 ;
        RECT 448.950 668.400 487.050 669.450 ;
        RECT 448.950 667.950 451.050 668.400 ;
        RECT 484.950 667.950 487.050 668.400 ;
        RECT 490.950 669.450 493.050 670.050 ;
        RECT 517.950 669.450 520.050 670.050 ;
        RECT 541.950 669.450 544.050 670.050 ;
        RECT 550.950 669.450 553.050 670.050 ;
        RECT 490.950 668.400 534.450 669.450 ;
        RECT 490.950 667.950 493.050 668.400 ;
        RECT 517.950 667.950 520.050 668.400 ;
        RECT 223.950 665.400 243.450 666.450 ;
        RECT 223.950 664.950 226.050 665.400 ;
        RECT 242.400 664.050 243.450 665.400 ;
        RECT 310.950 665.400 351.450 666.450 ;
        RECT 364.950 666.450 367.050 667.050 ;
        RECT 385.800 666.450 387.900 667.050 ;
        RECT 364.950 665.400 387.900 666.450 ;
        RECT 310.950 664.950 313.050 665.400 ;
        RECT 331.950 664.950 334.050 665.400 ;
        RECT 364.950 664.950 367.050 665.400 ;
        RECT 385.800 664.950 387.900 665.400 ;
        RECT 389.100 666.450 391.200 667.050 ;
        RECT 406.950 666.450 409.050 667.050 ;
        RECT 389.100 665.400 409.050 666.450 ;
        RECT 416.400 666.450 417.450 667.950 ;
        RECT 457.950 666.450 460.050 667.050 ;
        RECT 416.400 665.400 460.050 666.450 ;
        RECT 389.100 664.950 391.200 665.400 ;
        RECT 406.950 664.950 409.050 665.400 ;
        RECT 457.950 664.950 460.050 665.400 ;
        RECT 478.950 666.450 481.050 667.050 ;
        RECT 499.950 666.450 502.050 667.050 ;
        RECT 478.950 665.400 502.050 666.450 ;
        RECT 478.950 664.950 481.050 665.400 ;
        RECT 499.950 664.950 502.050 665.400 ;
        RECT 511.950 666.450 514.050 667.050 ;
        RECT 529.950 666.450 532.050 667.050 ;
        RECT 511.950 665.400 532.050 666.450 ;
        RECT 533.400 666.450 534.450 668.400 ;
        RECT 541.950 668.400 553.050 669.450 ;
        RECT 541.950 667.950 544.050 668.400 ;
        RECT 550.950 667.950 553.050 668.400 ;
        RECT 559.950 669.450 562.050 670.050 ;
        RECT 595.800 669.450 597.900 670.050 ;
        RECT 559.950 668.400 597.900 669.450 ;
        RECT 559.950 667.950 562.050 668.400 ;
        RECT 595.800 667.950 597.900 668.400 ;
        RECT 604.950 669.450 607.050 670.050 ;
        RECT 622.950 669.450 625.050 670.050 ;
        RECT 604.950 668.400 625.050 669.450 ;
        RECT 604.950 667.950 607.050 668.400 ;
        RECT 622.950 667.950 625.050 668.400 ;
        RECT 631.950 669.450 634.050 670.050 ;
        RECT 637.950 669.450 640.050 670.050 ;
        RECT 631.950 668.400 640.050 669.450 ;
        RECT 631.950 667.950 634.050 668.400 ;
        RECT 637.950 667.950 640.050 668.400 ;
        RECT 655.950 669.450 658.050 670.050 ;
        RECT 667.950 669.450 670.050 670.050 ;
        RECT 679.950 669.450 682.050 670.050 ;
        RECT 655.950 668.400 682.050 669.450 ;
        RECT 655.950 667.950 658.050 668.400 ;
        RECT 667.950 667.950 670.050 668.400 ;
        RECT 679.950 667.950 682.050 668.400 ;
        RECT 697.950 669.450 700.050 670.050 ;
        RECT 709.950 669.450 712.050 670.050 ;
        RECT 697.950 668.400 712.050 669.450 ;
        RECT 697.950 667.950 700.050 668.400 ;
        RECT 709.950 667.950 712.050 668.400 ;
        RECT 718.950 669.450 721.050 670.050 ;
        RECT 724.950 669.450 727.050 670.050 ;
        RECT 718.950 668.400 727.050 669.450 ;
        RECT 718.950 667.950 721.050 668.400 ;
        RECT 724.950 667.950 727.050 668.400 ;
        RECT 733.950 669.450 736.050 670.050 ;
        RECT 754.950 669.450 757.050 670.050 ;
        RECT 766.800 669.450 768.900 670.050 ;
        RECT 733.950 668.400 753.450 669.450 ;
        RECT 733.950 667.950 736.050 668.400 ;
        RECT 553.950 666.450 556.050 667.050 ;
        RECT 652.950 666.450 655.050 667.050 ;
        RECT 533.400 665.400 556.050 666.450 ;
        RECT 511.950 664.950 514.050 665.400 ;
        RECT 529.950 664.950 532.050 665.400 ;
        RECT 553.950 664.950 556.050 665.400 ;
        RECT 614.400 665.400 655.050 666.450 ;
        RECT 7.950 661.950 10.050 664.050 ;
        RECT 13.950 663.450 16.050 664.050 ;
        RECT 55.950 663.450 58.050 664.050 ;
        RECT 13.950 662.400 58.050 663.450 ;
        RECT 13.950 661.950 16.050 662.400 ;
        RECT 55.950 661.950 58.050 662.400 ;
        RECT 85.950 663.450 88.050 664.050 ;
        RECT 97.950 663.450 100.050 664.050 ;
        RECT 85.950 662.400 100.050 663.450 ;
        RECT 85.950 661.950 88.050 662.400 ;
        RECT 97.950 661.950 100.050 662.400 ;
        RECT 205.950 663.450 208.050 664.050 ;
        RECT 217.950 663.450 220.050 664.050 ;
        RECT 205.950 662.400 220.050 663.450 ;
        RECT 205.950 661.950 208.050 662.400 ;
        RECT 217.950 661.950 220.050 662.400 ;
        RECT 8.400 658.050 9.450 661.950 ;
        RECT 10.950 660.450 13.050 661.050 ;
        RECT 31.950 660.450 34.050 661.050 ;
        RECT 37.950 660.450 40.050 661.050 ;
        RECT 10.950 659.400 40.050 660.450 ;
        RECT 10.950 658.950 13.050 659.400 ;
        RECT 31.950 658.950 34.050 659.400 ;
        RECT 37.950 658.950 40.050 659.400 ;
        RECT 64.950 660.450 67.050 661.050 ;
        RECT 130.950 660.450 133.050 661.050 ;
        RECT 64.950 659.400 133.050 660.450 ;
        RECT 64.950 658.950 67.050 659.400 ;
        RECT 130.950 658.950 133.050 659.400 ;
        RECT 169.950 660.450 172.050 661.050 ;
        RECT 181.950 660.450 184.050 661.050 ;
        RECT 169.950 659.400 184.050 660.450 ;
        RECT 169.950 658.950 172.050 659.400 ;
        RECT 181.950 658.950 184.050 659.400 ;
        RECT 187.950 660.450 190.050 661.050 ;
        RECT 223.950 660.450 226.050 661.050 ;
        RECT 229.950 660.450 232.050 661.050 ;
        RECT 187.950 659.400 232.050 660.450 ;
        RECT 187.950 658.950 190.050 659.400 ;
        RECT 223.950 658.950 226.050 659.400 ;
        RECT 229.950 658.950 232.050 659.400 ;
        RECT 235.950 658.950 238.050 664.050 ;
        RECT 241.950 663.450 244.050 664.050 ;
        RECT 283.950 663.450 286.050 664.050 ;
        RECT 301.800 663.450 303.900 664.050 ;
        RECT 241.950 662.400 279.450 663.450 ;
        RECT 241.950 661.950 244.050 662.400 ;
        RECT 247.950 660.450 250.050 661.050 ;
        RECT 256.800 660.450 258.900 661.050 ;
        RECT 247.950 659.400 258.900 660.450 ;
        RECT 278.400 660.450 279.450 662.400 ;
        RECT 283.950 662.400 303.900 663.450 ;
        RECT 283.950 661.950 286.050 662.400 ;
        RECT 301.800 661.950 303.900 662.400 ;
        RECT 305.100 663.450 307.200 664.050 ;
        RECT 442.800 663.450 444.900 664.050 ;
        RECT 305.100 662.400 444.900 663.450 ;
        RECT 305.100 661.950 307.200 662.400 ;
        RECT 442.800 661.950 444.900 662.400 ;
        RECT 446.100 663.450 448.200 664.050 ;
        RECT 472.950 663.450 475.050 664.050 ;
        RECT 496.800 663.450 498.900 664.050 ;
        RECT 446.100 662.400 498.900 663.450 ;
        RECT 500.400 663.450 501.450 664.950 ;
        RECT 614.400 663.450 615.450 665.400 ;
        RECT 652.950 664.950 655.050 665.400 ;
        RECT 715.950 666.450 718.050 667.050 ;
        RECT 727.950 666.450 730.050 667.050 ;
        RECT 715.950 665.400 730.050 666.450 ;
        RECT 752.400 666.450 753.450 668.400 ;
        RECT 754.950 668.400 768.900 669.450 ;
        RECT 754.950 667.950 757.050 668.400 ;
        RECT 766.800 667.950 768.900 668.400 ;
        RECT 770.100 667.950 774.900 670.050 ;
        RECT 820.950 669.450 823.050 670.050 ;
        RECT 832.950 669.450 835.050 670.050 ;
        RECT 877.950 669.450 880.050 670.050 ;
        RECT 820.950 668.400 831.450 669.450 ;
        RECT 820.950 667.950 823.050 668.400 ;
        RECT 823.950 666.450 826.050 667.050 ;
        RECT 752.400 665.400 826.050 666.450 ;
        RECT 830.400 666.450 831.450 668.400 ;
        RECT 832.950 668.400 880.050 669.450 ;
        RECT 832.950 667.950 835.050 668.400 ;
        RECT 877.950 667.950 880.050 668.400 ;
        RECT 904.950 667.950 910.050 670.050 ;
        RECT 838.800 666.450 840.900 667.050 ;
        RECT 830.400 665.400 840.900 666.450 ;
        RECT 715.950 664.950 718.050 665.400 ;
        RECT 727.950 664.950 730.050 665.400 ;
        RECT 823.950 664.950 826.050 665.400 ;
        RECT 838.800 664.950 840.900 665.400 ;
        RECT 842.100 666.450 844.200 667.050 ;
        RECT 856.950 666.450 859.050 667.050 ;
        RECT 842.100 665.400 859.050 666.450 ;
        RECT 842.100 664.950 844.200 665.400 ;
        RECT 856.950 664.950 859.050 665.400 ;
        RECT 500.400 662.400 615.450 663.450 ;
        RECT 685.950 663.450 688.050 664.200 ;
        RECT 709.950 663.450 712.050 664.050 ;
        RECT 685.950 662.400 712.050 663.450 ;
        RECT 446.100 661.950 448.200 662.400 ;
        RECT 472.950 661.950 475.050 662.400 ;
        RECT 496.800 661.950 498.900 662.400 ;
        RECT 685.950 662.100 688.050 662.400 ;
        RECT 709.950 661.950 712.050 662.400 ;
        RECT 724.950 663.450 727.050 664.050 ;
        RECT 760.950 663.450 763.050 664.050 ;
        RECT 724.950 662.400 763.050 663.450 ;
        RECT 724.950 661.950 727.050 662.400 ;
        RECT 760.950 661.950 763.050 662.400 ;
        RECT 790.950 663.450 793.050 664.050 ;
        RECT 796.950 663.450 799.050 664.050 ;
        RECT 790.950 662.400 799.050 663.450 ;
        RECT 790.950 661.950 793.050 662.400 ;
        RECT 796.950 661.950 799.050 662.400 ;
        RECT 349.950 660.450 352.050 661.050 ;
        RECT 373.950 660.450 376.050 661.050 ;
        RECT 278.400 659.400 285.450 660.450 ;
        RECT 247.950 658.950 250.050 659.400 ;
        RECT 256.800 658.950 258.900 659.400 ;
        RECT 7.950 655.950 10.050 658.050 ;
        RECT 19.950 657.450 22.050 658.050 ;
        RECT 43.950 657.450 46.050 658.050 ;
        RECT 49.950 657.450 52.050 658.050 ;
        RECT 19.950 656.400 52.050 657.450 ;
        RECT 19.950 655.950 22.050 656.400 ;
        RECT 43.950 655.950 46.050 656.400 ;
        RECT 49.950 655.950 52.050 656.400 ;
        RECT 94.950 657.450 97.050 658.050 ;
        RECT 136.950 657.450 139.050 658.050 ;
        RECT 94.950 656.400 139.050 657.450 ;
        RECT 142.950 656.400 145.050 658.500 ;
        RECT 163.950 656.400 166.050 658.500 ;
        RECT 208.950 657.450 211.050 658.050 ;
        RECT 238.950 657.450 241.050 658.050 ;
        RECT 208.950 656.400 241.050 657.450 ;
        RECT 94.950 655.950 97.050 656.400 ;
        RECT 136.950 655.950 139.050 656.400 ;
        RECT 13.950 649.950 16.050 655.050 ;
        RECT 79.950 652.950 82.050 655.050 ;
        RECT 85.950 652.950 88.050 655.050 ;
        RECT 19.950 649.950 22.050 652.050 ;
        RECT 37.950 649.950 40.050 652.050 ;
        RECT 43.950 651.450 46.050 652.050 ;
        RECT 48.000 651.450 52.050 652.050 ;
        RECT 43.950 650.400 52.050 651.450 ;
        RECT 43.950 649.950 46.050 650.400 ;
        RECT 48.000 649.950 52.050 650.400 ;
        RECT 64.950 649.950 67.050 652.050 ;
        RECT 79.950 649.950 82.050 651.750 ;
        RECT 85.950 649.950 88.050 651.750 ;
        RECT 97.950 649.950 103.050 652.050 ;
        RECT 106.950 651.450 109.050 652.050 ;
        RECT 118.950 651.450 121.050 652.050 ;
        RECT 106.950 650.400 121.050 651.450 ;
        RECT 106.950 649.950 109.050 650.400 ;
        RECT 118.950 649.950 121.050 650.400 ;
        RECT 124.950 649.950 127.050 652.050 ;
        RECT 130.950 649.950 133.050 655.050 ;
        RECT 13.950 646.950 16.050 648.750 ;
        RECT 19.950 646.950 22.050 648.750 ;
        RECT 16.950 644.250 19.050 646.050 ;
        RECT 22.950 644.250 25.050 646.050 ;
        RECT 28.950 643.950 31.050 649.050 ;
        RECT 37.950 646.950 40.050 648.750 ;
        RECT 43.950 646.950 46.050 648.750 ;
        RECT 64.950 646.950 67.050 648.750 ;
        RECT 82.950 647.250 85.050 649.050 ;
        RECT 100.950 646.950 103.050 648.750 ;
        RECT 106.950 646.950 109.050 648.750 ;
        RECT 124.950 646.950 127.050 648.750 ;
        RECT 130.950 646.950 133.050 648.750 ;
        RECT 139.950 647.250 142.050 649.050 ;
        RECT 34.950 644.250 37.050 646.050 ;
        RECT 40.950 644.250 43.050 646.050 ;
        RECT 61.950 644.250 64.050 646.050 ;
        RECT 70.950 645.450 73.050 646.050 ;
        RECT 82.950 645.450 85.050 646.050 ;
        RECT 70.950 644.400 85.050 645.450 ;
        RECT 70.950 643.950 73.050 644.400 ;
        RECT 82.950 643.950 85.050 644.400 ;
        RECT 103.950 644.250 106.050 646.050 ;
        RECT 109.950 644.250 112.050 646.050 ;
        RECT 121.950 644.250 124.050 646.050 ;
        RECT 127.950 644.250 130.050 646.050 ;
        RECT 139.950 643.950 142.050 646.050 ;
        RECT 16.950 640.950 19.050 643.050 ;
        RECT 22.950 640.950 25.050 643.050 ;
        RECT 34.950 640.950 37.050 643.050 ;
        RECT 40.950 640.950 43.050 643.050 ;
        RECT 46.950 642.450 49.050 643.050 ;
        RECT 61.950 642.450 64.050 643.050 ;
        RECT 76.950 642.450 79.050 643.050 ;
        RECT 46.950 641.400 79.050 642.450 ;
        RECT 46.950 640.950 49.050 641.400 ;
        RECT 61.950 640.950 64.050 641.400 ;
        RECT 76.950 640.950 79.050 641.400 ;
        RECT 103.950 640.950 106.050 643.050 ;
        RECT 109.950 640.950 112.050 643.050 ;
        RECT 121.950 640.950 124.050 643.050 ;
        RECT 127.950 640.950 130.050 643.050 ;
        RECT 82.950 639.450 85.050 640.050 ;
        RECT 91.950 639.450 94.050 640.050 ;
        RECT 82.950 638.400 94.050 639.450 ;
        RECT 82.950 637.950 85.050 638.400 ;
        RECT 91.950 637.950 94.050 638.400 ;
        RECT 34.950 636.450 37.050 637.050 ;
        RECT 49.950 636.450 52.050 637.050 ;
        RECT 34.950 635.400 52.050 636.450 ;
        RECT 34.950 634.950 37.050 635.400 ;
        RECT 49.950 634.950 52.050 635.400 ;
        RECT 112.950 636.450 115.050 637.050 ;
        RECT 127.950 636.450 130.050 637.050 ;
        RECT 143.700 636.600 144.900 656.400 ;
        RECT 148.950 647.250 151.050 649.050 ;
        RECT 148.950 643.950 151.050 646.050 ;
        RECT 163.950 641.400 165.150 656.400 ;
        RECT 208.950 655.950 211.050 656.400 ;
        RECT 238.950 655.950 241.050 656.400 ;
        RECT 244.950 657.450 247.050 658.050 ;
        RECT 280.950 657.450 283.050 658.050 ;
        RECT 244.950 656.400 283.050 657.450 ;
        RECT 284.400 657.450 285.450 659.400 ;
        RECT 349.950 659.400 376.050 660.450 ;
        RECT 349.950 658.950 352.050 659.400 ;
        RECT 373.950 658.950 376.050 659.400 ;
        RECT 406.950 660.450 409.050 661.050 ;
        RECT 430.950 660.450 433.050 661.050 ;
        RECT 406.950 659.400 433.050 660.450 ;
        RECT 406.950 658.950 409.050 659.400 ;
        RECT 430.950 658.950 433.050 659.400 ;
        RECT 442.950 660.450 445.050 661.050 ;
        RECT 448.800 660.450 450.900 661.050 ;
        RECT 442.950 659.400 450.900 660.450 ;
        RECT 442.950 658.950 445.050 659.400 ;
        RECT 448.800 658.950 450.900 659.400 ;
        RECT 452.100 660.450 454.200 661.050 ;
        RECT 469.950 660.450 472.050 661.050 ;
        RECT 452.100 659.400 472.050 660.450 ;
        RECT 452.100 658.950 454.200 659.400 ;
        RECT 469.950 658.950 472.050 659.400 ;
        RECT 493.950 660.450 496.050 661.050 ;
        RECT 517.950 660.450 520.050 661.050 ;
        RECT 493.950 659.400 520.050 660.450 ;
        RECT 493.950 658.950 496.050 659.400 ;
        RECT 517.950 658.950 520.050 659.400 ;
        RECT 553.950 660.450 556.050 661.050 ;
        RECT 577.800 660.450 579.900 661.050 ;
        RECT 553.950 659.400 579.900 660.450 ;
        RECT 553.950 658.950 556.050 659.400 ;
        RECT 577.800 658.950 579.900 659.400 ;
        RECT 581.100 660.450 583.200 661.050 ;
        RECT 592.950 660.450 595.050 661.050 ;
        RECT 604.950 660.450 607.050 661.050 ;
        RECT 581.100 659.400 595.050 660.450 ;
        RECT 581.100 658.950 583.200 659.400 ;
        RECT 592.950 658.950 595.050 659.400 ;
        RECT 596.400 659.400 607.050 660.450 ;
        RECT 325.800 657.450 327.900 658.050 ;
        RECT 284.400 656.400 327.900 657.450 ;
        RECT 379.950 656.400 382.050 658.500 ;
        RECT 400.950 656.400 403.050 658.500 ;
        RECT 409.950 657.450 412.050 658.050 ;
        RECT 421.950 657.450 424.050 658.050 ;
        RECT 409.950 656.400 424.050 657.450 ;
        RECT 244.950 655.950 247.050 656.400 ;
        RECT 280.950 655.950 283.050 656.400 ;
        RECT 325.800 655.950 327.900 656.400 ;
        RECT 181.950 652.950 184.050 655.050 ;
        RECT 187.950 652.950 190.050 655.050 ;
        RECT 166.950 649.950 169.050 652.050 ;
        RECT 181.950 649.950 184.050 651.750 ;
        RECT 187.950 649.950 190.050 651.750 ;
        RECT 199.950 651.450 202.050 652.050 ;
        RECT 205.950 651.450 208.050 652.050 ;
        RECT 194.400 650.400 208.050 651.450 ;
        RECT 194.400 649.050 195.450 650.400 ;
        RECT 199.950 649.950 202.050 650.400 ;
        RECT 205.950 649.950 208.050 650.400 ;
        RECT 229.950 649.950 232.050 652.050 ;
        RECT 235.950 651.450 238.050 652.050 ;
        RECT 247.950 651.450 250.050 652.050 ;
        RECT 235.950 650.400 250.050 651.450 ;
        RECT 235.950 649.950 238.050 650.400 ;
        RECT 247.950 649.950 250.050 650.400 ;
        RECT 253.950 649.950 256.050 652.050 ;
        RECT 295.950 649.950 298.050 655.050 ;
        RECT 301.950 651.450 304.050 652.050 ;
        RECT 316.950 651.450 319.050 652.050 ;
        RECT 301.950 650.400 319.050 651.450 ;
        RECT 301.950 649.950 304.050 650.400 ;
        RECT 316.950 649.950 319.050 650.400 ;
        RECT 322.950 649.950 325.050 652.050 ;
        RECT 334.950 649.950 337.050 652.050 ;
        RECT 340.950 651.450 343.050 652.050 ;
        RECT 355.950 651.450 358.050 652.050 ;
        RECT 340.950 650.400 358.050 651.450 ;
        RECT 340.950 649.950 343.050 650.400 ;
        RECT 355.950 649.950 358.050 650.400 ;
        RECT 364.950 649.950 367.050 652.050 ;
        RECT 370.950 649.950 373.050 652.050 ;
        RECT 166.950 646.950 169.050 648.750 ;
        RECT 184.950 647.250 187.050 649.050 ;
        RECT 190.950 647.400 195.450 649.050 ;
        RECT 190.950 646.950 195.000 647.400 ;
        RECT 205.950 646.950 208.050 648.750 ;
        RECT 229.950 646.950 232.050 648.750 ;
        RECT 247.950 646.950 250.050 648.750 ;
        RECT 253.950 646.950 256.050 648.750 ;
        RECT 265.950 647.250 268.050 649.050 ;
        RECT 275.250 648.750 277.050 649.050 ;
        RECT 271.950 647.250 274.050 648.750 ;
        RECT 274.950 647.250 277.050 648.750 ;
        RECT 271.950 646.950 273.750 647.250 ;
        RECT 295.950 646.950 298.050 648.750 ;
        RECT 316.950 646.950 319.050 648.750 ;
        RECT 322.950 646.950 325.050 648.750 ;
        RECT 334.950 646.950 337.050 648.750 ;
        RECT 340.950 646.950 343.050 648.750 ;
        RECT 364.950 646.950 367.050 648.750 ;
        RECT 370.950 646.950 373.050 648.750 ;
        RECT 376.950 647.250 379.050 649.050 ;
        RECT 184.950 643.950 190.050 646.050 ;
        RECT 202.950 644.250 205.050 646.050 ;
        RECT 208.950 644.250 211.050 646.050 ;
        RECT 226.950 644.250 229.050 646.050 ;
        RECT 232.950 643.950 238.050 646.050 ;
        RECT 244.950 644.250 247.050 646.050 ;
        RECT 250.950 644.250 253.050 646.050 ;
        RECT 262.950 643.950 268.050 646.050 ;
        RECT 274.950 645.450 277.050 646.050 ;
        RECT 280.950 645.450 283.050 646.050 ;
        RECT 286.950 645.450 289.050 646.050 ;
        RECT 274.950 644.400 289.050 645.450 ;
        RECT 274.950 643.950 277.050 644.400 ;
        RECT 280.950 643.950 283.050 644.400 ;
        RECT 286.950 643.950 289.050 644.400 ;
        RECT 292.950 644.250 295.050 646.050 ;
        RECT 298.950 644.250 301.050 646.050 ;
        RECT 313.950 644.250 316.050 646.050 ;
        RECT 319.950 644.250 322.050 646.050 ;
        RECT 325.950 643.950 331.050 646.050 ;
        RECT 337.950 644.250 340.050 646.050 ;
        RECT 343.950 644.250 346.050 646.050 ;
        RECT 361.950 644.250 364.050 646.050 ;
        RECT 367.950 644.250 370.050 646.050 ;
        RECT 376.950 643.950 379.050 646.050 ;
        RECT 169.950 642.450 172.050 643.200 ;
        RECT 178.950 642.450 181.050 643.050 ;
        RECT 169.950 641.400 181.050 642.450 ;
        RECT 151.950 639.450 154.050 640.050 ;
        RECT 157.950 639.450 160.050 640.050 ;
        RECT 151.950 638.400 160.050 639.450 ;
        RECT 151.950 637.950 154.050 638.400 ;
        RECT 157.950 637.950 160.050 638.400 ;
        RECT 163.950 639.300 166.050 641.400 ;
        RECT 169.950 641.100 172.050 641.400 ;
        RECT 178.950 640.950 181.050 641.400 ;
        RECT 202.950 640.950 205.050 643.050 ;
        RECT 208.950 640.950 211.050 643.050 ;
        RECT 226.950 640.950 229.050 643.050 ;
        RECT 244.950 640.950 247.050 643.050 ;
        RECT 250.950 640.950 253.050 643.050 ;
        RECT 292.950 640.950 295.050 643.050 ;
        RECT 298.950 640.950 301.050 643.050 ;
        RECT 313.950 640.950 316.050 643.050 ;
        RECT 319.950 640.950 322.050 643.050 ;
        RECT 169.950 639.450 172.050 639.900 ;
        RECT 196.950 639.450 199.050 640.050 ;
        RECT 112.950 635.400 130.050 636.450 ;
        RECT 112.950 634.950 115.050 635.400 ;
        RECT 127.950 634.950 130.050 635.400 ;
        RECT 142.950 634.500 145.050 636.600 ;
        RECT 163.950 635.700 165.150 639.300 ;
        RECT 169.950 638.400 199.050 639.450 ;
        RECT 169.950 637.800 172.050 638.400 ;
        RECT 196.950 637.950 199.050 638.400 ;
        RECT 265.950 639.450 268.050 640.200 ;
        RECT 286.950 639.450 289.050 640.050 ;
        RECT 265.950 638.400 289.050 639.450 ;
        RECT 265.950 638.100 268.050 638.400 ;
        RECT 286.950 637.950 289.050 638.400 ;
        RECT 322.950 639.450 325.050 640.050 ;
        RECT 337.950 639.450 340.050 643.050 ;
        RECT 343.950 640.950 346.050 643.050 ;
        RECT 361.950 640.950 364.050 643.050 ;
        RECT 367.950 640.950 370.050 643.050 ;
        RECT 322.950 638.400 340.050 639.450 ;
        RECT 322.950 637.950 325.050 638.400 ;
        RECT 178.950 636.450 181.050 637.050 ;
        RECT 184.950 636.450 187.050 637.050 ;
        RECT 202.950 636.450 205.050 637.050 ;
        RECT 91.950 633.450 94.050 634.050 ;
        RECT 133.950 633.450 136.050 634.050 ;
        RECT 163.950 633.600 166.050 635.700 ;
        RECT 178.950 635.400 187.050 636.450 ;
        RECT 178.950 634.950 181.050 635.400 ;
        RECT 184.950 634.950 187.050 635.400 ;
        RECT 194.400 635.400 205.050 636.450 ;
        RECT 91.950 632.400 136.050 633.450 ;
        RECT 91.950 631.950 94.050 632.400 ;
        RECT 133.950 631.950 136.050 632.400 ;
        RECT 175.950 633.450 178.050 634.050 ;
        RECT 194.400 633.450 195.450 635.400 ;
        RECT 202.950 634.950 205.050 635.400 ;
        RECT 226.950 636.450 229.050 637.050 ;
        RECT 256.950 636.450 259.050 637.050 ;
        RECT 226.950 635.400 259.050 636.450 ;
        RECT 226.950 634.950 229.050 635.400 ;
        RECT 256.950 634.950 259.050 635.400 ;
        RECT 265.950 636.450 268.050 636.900 ;
        RECT 277.950 636.450 280.050 637.050 ;
        RECT 313.950 636.450 316.050 637.050 ;
        RECT 380.700 636.600 381.900 656.400 ;
        RECT 385.950 647.250 388.050 649.050 ;
        RECT 385.950 643.950 388.050 646.050 ;
        RECT 400.950 641.400 402.150 656.400 ;
        RECT 409.950 655.950 412.050 656.400 ;
        RECT 421.950 655.950 424.050 656.400 ;
        RECT 427.950 657.450 430.050 658.050 ;
        RECT 478.800 657.450 480.900 658.050 ;
        RECT 427.950 656.400 480.900 657.450 ;
        RECT 427.950 655.950 430.050 656.400 ;
        RECT 478.800 655.950 480.900 656.400 ;
        RECT 482.100 657.450 484.200 658.050 ;
        RECT 508.950 657.450 511.050 658.050 ;
        RECT 482.100 656.400 511.050 657.450 ;
        RECT 526.950 656.400 529.050 658.500 ;
        RECT 547.950 656.400 550.050 658.500 ;
        RECT 589.950 657.450 592.050 658.050 ;
        RECT 596.400 657.450 597.450 659.400 ;
        RECT 604.950 658.950 607.050 659.400 ;
        RECT 625.950 660.450 628.050 661.050 ;
        RECT 637.950 660.450 640.050 661.050 ;
        RECT 625.950 659.400 640.050 660.450 ;
        RECT 625.950 658.950 628.050 659.400 ;
        RECT 637.950 658.950 640.050 659.400 ;
        RECT 643.950 660.450 646.050 661.050 ;
        RECT 655.950 660.450 658.050 661.050 ;
        RECT 643.950 659.400 658.050 660.450 ;
        RECT 643.950 658.950 646.050 659.400 ;
        RECT 655.950 658.950 658.050 659.400 ;
        RECT 703.950 660.450 706.050 661.050 ;
        RECT 730.800 660.450 732.900 661.050 ;
        RECT 703.950 659.400 732.900 660.450 ;
        RECT 703.950 658.950 706.050 659.400 ;
        RECT 730.800 658.950 732.900 659.400 ;
        RECT 734.100 660.450 736.200 661.200 ;
        RECT 739.950 660.450 742.050 661.050 ;
        RECT 835.950 660.450 838.050 661.050 ;
        RECT 734.100 659.400 742.050 660.450 ;
        RECT 734.100 659.100 736.200 659.400 ;
        RECT 739.950 658.950 742.050 659.400 ;
        RECT 764.400 659.400 838.050 660.450 ;
        RECT 764.400 658.050 765.450 659.400 ;
        RECT 835.950 658.950 838.050 659.400 ;
        RECT 856.950 660.450 859.050 661.050 ;
        RECT 862.800 660.450 864.900 661.050 ;
        RECT 856.950 659.400 864.900 660.450 ;
        RECT 856.950 658.950 859.050 659.400 ;
        RECT 862.800 658.950 864.900 659.400 ;
        RECT 866.100 660.450 868.200 661.050 ;
        RECT 880.950 660.450 883.050 661.050 ;
        RECT 866.100 659.400 883.050 660.450 ;
        RECT 866.100 658.950 868.200 659.400 ;
        RECT 880.950 658.950 883.050 659.400 ;
        RECT 589.950 656.400 597.450 657.450 ;
        RECT 598.950 657.450 601.050 658.050 ;
        RECT 613.950 657.450 616.050 658.050 ;
        RECT 598.950 656.400 616.050 657.450 ;
        RECT 482.100 655.950 484.200 656.400 ;
        RECT 508.950 655.950 511.050 656.400 ;
        RECT 454.950 654.450 457.050 655.050 ;
        RECT 463.950 654.450 466.050 655.050 ;
        RECT 454.950 653.400 466.050 654.450 ;
        RECT 454.950 652.950 457.050 653.400 ;
        RECT 463.950 652.950 466.050 653.400 ;
        RECT 403.950 649.950 406.050 652.050 ;
        RECT 421.950 649.950 424.050 652.050 ;
        RECT 427.950 651.450 430.050 652.050 ;
        RECT 442.950 651.450 445.050 652.050 ;
        RECT 427.950 650.400 445.050 651.450 ;
        RECT 427.950 649.950 430.050 650.400 ;
        RECT 442.950 649.950 445.050 650.400 ;
        RECT 448.950 649.950 451.050 652.050 ;
        RECT 466.950 649.950 472.050 652.050 ;
        RECT 493.950 649.950 496.050 652.050 ;
        RECT 511.950 649.950 514.050 652.050 ;
        RECT 517.950 649.950 520.050 652.050 ;
        RECT 445.950 648.750 447.750 649.050 ;
        RECT 403.950 646.950 406.050 648.750 ;
        RECT 421.950 646.950 424.050 648.750 ;
        RECT 427.950 646.950 430.050 648.750 ;
        RECT 445.950 647.250 448.050 648.750 ;
        RECT 448.950 647.250 451.050 648.750 ;
        RECT 454.950 647.250 457.050 649.050 ;
        RECT 449.250 646.950 451.050 647.250 ;
        RECT 469.950 646.950 472.050 648.750 ;
        RECT 475.950 648.450 478.050 649.050 ;
        RECT 481.950 648.450 484.050 649.050 ;
        RECT 475.950 647.400 484.050 648.450 ;
        RECT 475.950 646.950 478.050 647.400 ;
        RECT 481.950 646.950 484.050 647.400 ;
        RECT 493.950 646.950 496.050 648.750 ;
        RECT 511.950 646.950 514.050 648.750 ;
        RECT 517.950 646.950 520.050 648.750 ;
        RECT 523.950 647.250 526.050 649.050 ;
        RECT 418.950 644.250 421.050 646.050 ;
        RECT 424.950 644.250 427.050 646.050 ;
        RECT 445.950 643.950 448.050 646.050 ;
        RECT 454.950 643.950 457.050 646.050 ;
        RECT 466.950 644.250 469.050 646.050 ;
        RECT 472.950 644.250 475.050 646.050 ;
        RECT 490.950 644.250 493.050 646.050 ;
        RECT 508.950 644.250 511.050 646.050 ;
        RECT 514.950 644.250 517.050 646.050 ;
        RECT 523.950 643.950 526.050 646.050 ;
        RECT 400.950 639.300 403.050 641.400 ;
        RECT 418.950 640.950 421.050 643.050 ;
        RECT 424.950 640.950 430.050 643.050 ;
        RECT 436.950 639.450 439.050 640.050 ;
        RECT 446.400 639.450 447.450 643.950 ;
        RECT 466.950 640.950 469.050 643.050 ;
        RECT 472.950 640.950 475.050 643.050 ;
        RECT 478.950 642.450 481.050 643.050 ;
        RECT 490.950 642.450 493.050 643.050 ;
        RECT 478.950 641.400 493.050 642.450 ;
        RECT 478.950 640.950 481.050 641.400 ;
        RECT 490.950 640.950 493.050 641.400 ;
        RECT 508.950 640.950 511.050 643.050 ;
        RECT 514.950 640.950 517.050 643.050 ;
        RECT 454.950 639.450 457.050 640.050 ;
        RECT 265.950 635.400 280.050 636.450 ;
        RECT 265.950 634.800 268.050 635.400 ;
        RECT 277.950 634.950 280.050 635.400 ;
        RECT 296.400 635.400 316.050 636.450 ;
        RECT 296.400 634.050 297.450 635.400 ;
        RECT 313.950 634.950 316.050 635.400 ;
        RECT 379.950 634.500 382.050 636.600 ;
        RECT 400.950 635.700 402.150 639.300 ;
        RECT 436.950 638.400 457.050 639.450 ;
        RECT 436.950 637.950 439.050 638.400 ;
        RECT 454.950 637.950 457.050 638.400 ;
        RECT 175.950 632.400 195.450 633.450 ;
        RECT 196.950 633.450 199.050 634.050 ;
        RECT 295.950 633.450 298.050 634.050 ;
        RECT 196.950 632.400 298.050 633.450 ;
        RECT 175.950 631.950 178.050 632.400 ;
        RECT 196.950 631.950 199.050 632.400 ;
        RECT 295.950 631.950 298.050 632.400 ;
        RECT 322.950 633.450 325.050 634.050 ;
        RECT 349.950 633.450 352.050 634.050 ;
        RECT 322.950 632.400 352.050 633.450 ;
        RECT 322.950 631.950 325.050 632.400 ;
        RECT 349.950 631.950 352.050 632.400 ;
        RECT 355.950 633.450 358.050 634.050 ;
        RECT 373.950 633.450 376.050 634.050 ;
        RECT 400.950 633.600 403.050 635.700 ;
        RECT 412.950 634.950 418.050 637.050 ;
        RECT 451.950 636.450 454.050 637.050 ;
        RECT 481.950 636.450 484.050 637.050 ;
        RECT 451.950 635.400 484.050 636.450 ;
        RECT 451.950 634.950 454.050 635.400 ;
        RECT 481.950 634.950 484.050 635.400 ;
        RECT 502.950 636.450 505.050 637.050 ;
        RECT 508.950 636.450 511.050 637.050 ;
        RECT 527.700 636.600 528.900 656.400 ;
        RECT 532.950 647.250 535.050 649.050 ;
        RECT 532.950 643.950 535.050 646.050 ;
        RECT 547.950 641.400 549.150 656.400 ;
        RECT 589.950 655.950 592.050 656.400 ;
        RECT 598.950 655.950 601.050 656.400 ;
        RECT 613.950 655.950 616.050 656.400 ;
        RECT 622.950 657.450 625.050 658.050 ;
        RECT 733.950 657.450 736.050 657.900 ;
        RECT 763.950 657.450 766.050 658.050 ;
        RECT 622.950 656.400 663.450 657.450 ;
        RECT 622.950 655.950 625.050 656.400 ;
        RECT 559.950 654.450 562.050 655.050 ;
        RECT 565.950 654.450 568.050 655.050 ;
        RECT 559.950 653.400 568.050 654.450 ;
        RECT 559.950 652.950 562.050 653.400 ;
        RECT 565.950 652.950 568.050 653.400 ;
        RECT 662.400 652.050 663.450 656.400 ;
        RECT 733.950 656.400 766.050 657.450 ;
        RECT 733.950 655.800 736.050 656.400 ;
        RECT 763.950 655.950 766.050 656.400 ;
        RECT 772.950 657.450 775.050 658.200 ;
        RECT 796.950 657.450 799.050 658.050 ;
        RECT 772.950 656.400 799.050 657.450 ;
        RECT 772.950 656.100 775.050 656.400 ;
        RECT 796.950 655.950 799.050 656.400 ;
        RECT 817.950 657.450 820.050 658.050 ;
        RECT 823.950 657.450 826.050 658.050 ;
        RECT 817.950 656.400 826.050 657.450 ;
        RECT 817.950 655.950 820.050 656.400 ;
        RECT 823.950 655.950 826.050 656.400 ;
        RECT 886.950 657.450 889.050 658.050 ;
        RECT 895.950 657.450 898.050 658.050 ;
        RECT 886.950 656.400 898.050 657.450 ;
        RECT 886.950 655.950 889.050 656.400 ;
        RECT 895.950 655.950 898.050 656.400 ;
        RECT 703.950 652.950 706.050 655.050 ;
        RECT 709.950 654.450 712.050 655.050 ;
        RECT 718.950 654.450 721.050 655.050 ;
        RECT 709.950 653.400 721.050 654.450 ;
        RECT 709.950 652.950 712.050 653.400 ;
        RECT 718.950 652.950 721.050 653.400 ;
        RECT 874.950 654.450 877.050 655.050 ;
        RECT 874.950 653.400 892.050 654.450 ;
        RECT 874.950 652.950 877.050 653.400 ;
        RECT 550.950 649.950 553.050 652.050 ;
        RECT 586.950 651.450 589.050 652.050 ;
        RECT 595.950 651.450 598.050 652.050 ;
        RECT 586.950 650.400 598.050 651.450 ;
        RECT 586.950 649.950 589.050 650.400 ;
        RECT 595.950 649.950 598.050 650.400 ;
        RECT 601.950 651.450 604.050 652.050 ;
        RECT 610.950 651.450 613.050 652.050 ;
        RECT 601.950 650.400 613.050 651.450 ;
        RECT 601.950 649.950 604.050 650.400 ;
        RECT 610.950 649.950 613.050 650.400 ;
        RECT 616.950 649.950 619.050 652.050 ;
        RECT 622.950 649.950 625.050 652.050 ;
        RECT 637.950 649.950 640.050 652.050 ;
        RECT 655.950 649.950 658.050 652.050 ;
        RECT 661.950 649.950 664.050 652.050 ;
        RECT 703.950 649.950 706.050 651.750 ;
        RECT 709.950 649.950 712.050 651.750 ;
        RECT 724.950 649.950 727.050 652.050 ;
        RECT 730.950 651.450 733.050 652.050 ;
        RECT 742.950 651.450 745.050 652.050 ;
        RECT 730.950 650.400 745.050 651.450 ;
        RECT 730.950 649.950 733.050 650.400 ;
        RECT 742.950 649.950 745.050 650.400 ;
        RECT 748.950 649.950 751.050 652.050 ;
        RECT 754.950 651.450 757.050 652.050 ;
        RECT 763.950 651.450 766.050 652.050 ;
        RECT 778.950 651.450 781.050 652.050 ;
        RECT 754.950 650.400 762.450 651.450 ;
        RECT 754.950 649.950 757.050 650.400 ;
        RECT 550.950 646.950 553.050 648.750 ;
        RECT 565.950 647.250 568.050 649.050 ;
        RECT 575.250 648.750 577.050 649.050 ;
        RECT 571.950 647.250 574.050 648.750 ;
        RECT 574.950 647.250 577.050 648.750 ;
        RECT 571.950 646.950 573.750 647.250 ;
        RECT 595.950 646.950 598.050 648.750 ;
        RECT 601.950 646.950 604.050 648.750 ;
        RECT 616.950 646.950 619.050 648.750 ;
        RECT 622.950 646.950 625.050 648.750 ;
        RECT 637.950 646.950 640.050 648.750 ;
        RECT 655.950 646.950 658.050 648.750 ;
        RECT 661.950 646.950 664.050 648.750 ;
        RECT 679.950 647.250 682.050 649.050 ;
        RECT 689.250 648.750 691.050 649.050 ;
        RECT 685.950 647.250 688.050 648.750 ;
        RECT 688.950 647.250 691.050 648.750 ;
        RECT 706.950 647.250 709.050 649.050 ;
        RECT 685.950 646.950 687.750 647.250 ;
        RECT 724.950 646.950 727.050 648.750 ;
        RECT 730.950 646.950 733.050 648.750 ;
        RECT 748.950 646.950 751.050 648.750 ;
        RECT 754.950 646.950 757.050 648.750 ;
        RECT 761.400 648.450 762.450 650.400 ;
        RECT 763.950 650.400 781.050 651.450 ;
        RECT 763.950 649.950 766.050 650.400 ;
        RECT 778.950 649.950 781.050 650.400 ;
        RECT 784.950 649.950 787.050 652.050 ;
        RECT 790.950 651.450 793.050 652.050 ;
        RECT 799.950 651.450 802.050 652.050 ;
        RECT 790.950 650.400 802.050 651.450 ;
        RECT 790.950 649.950 793.050 650.400 ;
        RECT 799.950 649.950 802.050 650.400 ;
        RECT 817.950 651.450 822.000 652.050 ;
        RECT 823.950 651.450 826.050 652.050 ;
        RECT 817.950 650.400 826.050 651.450 ;
        RECT 817.950 649.950 822.000 650.400 ;
        RECT 823.950 649.950 826.050 650.400 ;
        RECT 841.950 649.950 844.050 652.050 ;
        RECT 859.950 651.450 864.000 652.050 ;
        RECT 865.950 651.450 868.050 652.050 ;
        RECT 859.950 650.400 868.050 651.450 ;
        RECT 859.950 649.950 864.000 650.400 ;
        RECT 865.950 649.950 868.050 650.400 ;
        RECT 871.950 649.950 874.050 652.050 ;
        RECT 889.950 649.950 892.050 653.400 ;
        RECT 895.950 651.450 898.050 652.050 ;
        RECT 900.000 651.450 904.050 652.050 ;
        RECT 895.950 650.400 904.050 651.450 ;
        RECT 895.950 649.950 898.050 650.400 ;
        RECT 900.000 649.950 904.050 650.400 ;
        RECT 772.950 648.450 775.050 649.050 ;
        RECT 761.400 647.400 775.050 648.450 ;
        RECT 772.950 646.950 775.050 647.400 ;
        RECT 778.950 646.950 781.050 648.750 ;
        RECT 784.950 646.950 787.050 648.750 ;
        RECT 799.950 646.950 802.050 648.750 ;
        RECT 823.950 646.950 826.050 648.750 ;
        RECT 841.950 646.950 844.050 648.750 ;
        RECT 847.950 647.250 850.050 649.050 ;
        RECT 865.950 646.950 868.050 648.750 ;
        RECT 871.950 646.950 874.050 648.750 ;
        RECT 889.950 646.950 892.050 648.750 ;
        RECT 895.950 646.950 898.050 648.750 ;
        RECT 565.950 643.950 568.050 646.050 ;
        RECT 574.950 645.450 577.050 646.050 ;
        RECT 586.950 645.450 589.050 646.050 ;
        RECT 574.950 644.400 589.050 645.450 ;
        RECT 574.950 643.950 577.050 644.400 ;
        RECT 586.950 643.950 589.050 644.400 ;
        RECT 592.950 644.250 595.050 646.050 ;
        RECT 598.950 644.250 601.050 646.050 ;
        RECT 619.950 644.250 622.050 646.050 ;
        RECT 625.950 644.250 628.050 646.050 ;
        RECT 640.950 644.250 643.050 646.050 ;
        RECT 658.950 644.250 661.050 646.050 ;
        RECT 664.950 644.250 667.050 646.050 ;
        RECT 679.950 643.950 682.050 646.050 ;
        RECT 688.950 643.950 691.050 646.050 ;
        RECT 706.950 643.950 712.050 646.050 ;
        RECT 727.950 644.250 730.050 646.050 ;
        RECT 733.950 644.250 736.050 646.050 ;
        RECT 742.950 643.950 748.050 646.050 ;
        RECT 751.950 644.250 754.050 646.050 ;
        RECT 757.950 644.250 760.050 646.050 ;
        RECT 775.950 644.250 778.050 646.050 ;
        RECT 781.950 644.250 784.050 646.050 ;
        RECT 796.950 644.250 799.050 646.050 ;
        RECT 802.950 644.250 805.050 646.050 ;
        RECT 820.950 644.250 823.050 646.050 ;
        RECT 826.950 644.250 829.050 646.050 ;
        RECT 838.950 644.250 841.050 646.050 ;
        RECT 547.950 639.300 550.050 641.400 ;
        RECT 592.950 640.950 595.050 643.050 ;
        RECT 598.950 640.950 601.050 643.050 ;
        RECT 619.950 640.950 622.050 643.050 ;
        RECT 625.950 640.950 628.050 643.050 ;
        RECT 640.950 640.950 646.050 643.050 ;
        RECT 658.950 640.950 661.050 643.050 ;
        RECT 664.950 640.950 667.050 643.050 ;
        RECT 689.400 639.450 690.450 643.950 ;
        RECT 727.950 640.950 730.050 643.050 ;
        RECT 733.950 640.950 736.050 643.050 ;
        RECT 751.950 640.950 754.050 643.050 ;
        RECT 757.950 640.950 760.050 643.050 ;
        RECT 775.950 640.950 778.050 643.050 ;
        RECT 781.950 640.950 784.050 643.050 ;
        RECT 793.950 640.950 799.050 643.050 ;
        RECT 826.950 640.950 829.050 643.050 ;
        RECT 838.950 640.950 841.050 643.050 ;
        RECT 847.950 640.950 850.050 646.050 ;
        RECT 868.950 644.250 871.050 646.050 ;
        RECT 874.950 644.250 877.050 646.050 ;
        RECT 886.950 644.250 889.050 646.050 ;
        RECT 892.950 644.250 895.050 646.050 ;
        RECT 868.950 640.950 871.050 643.050 ;
        RECT 874.950 640.950 877.050 643.050 ;
        RECT 886.950 640.950 889.050 643.050 ;
        RECT 892.950 640.950 895.050 643.050 ;
        RECT 502.950 635.400 511.050 636.450 ;
        RECT 502.950 634.950 505.050 635.400 ;
        RECT 508.950 634.950 511.050 635.400 ;
        RECT 526.950 634.500 529.050 636.600 ;
        RECT 547.950 635.700 549.150 639.300 ;
        RECT 671.400 638.400 690.450 639.450 ;
        RECT 691.950 639.450 694.050 640.050 ;
        RECT 724.950 639.450 727.050 640.050 ;
        RECT 691.950 638.400 727.050 639.450 ;
        RECT 671.400 637.050 672.450 638.400 ;
        RECT 691.950 637.950 694.050 638.400 ;
        RECT 724.950 637.950 727.050 638.400 ;
        RECT 739.950 639.450 742.050 640.050 ;
        RECT 745.950 639.450 748.050 640.050 ;
        RECT 739.950 638.400 748.050 639.450 ;
        RECT 739.950 637.950 742.050 638.400 ;
        RECT 745.950 637.950 748.050 638.400 ;
        RECT 784.950 639.450 787.050 640.050 ;
        RECT 790.950 639.450 793.050 640.050 ;
        RECT 784.950 638.400 793.050 639.450 ;
        RECT 784.950 637.950 787.050 638.400 ;
        RECT 790.950 637.950 793.050 638.400 ;
        RECT 562.950 636.450 565.050 637.050 ;
        RECT 580.950 636.450 583.050 637.050 ;
        RECT 355.950 632.400 376.050 633.450 ;
        RECT 355.950 631.950 358.050 632.400 ;
        RECT 373.950 631.950 376.050 632.400 ;
        RECT 409.950 633.450 412.050 634.050 ;
        RECT 445.800 633.450 447.900 634.050 ;
        RECT 409.950 632.400 447.900 633.450 ;
        RECT 409.950 631.950 412.050 632.400 ;
        RECT 445.800 631.950 447.900 632.400 ;
        RECT 449.100 633.450 451.200 634.050 ;
        RECT 457.950 633.450 460.050 634.050 ;
        RECT 466.950 633.450 469.050 634.050 ;
        RECT 449.100 632.400 469.050 633.450 ;
        RECT 449.100 631.950 451.200 632.400 ;
        RECT 457.950 631.950 460.050 632.400 ;
        RECT 466.950 631.950 469.050 632.400 ;
        RECT 484.950 633.450 487.050 634.050 ;
        RECT 547.950 633.600 550.050 635.700 ;
        RECT 562.950 635.400 583.050 636.450 ;
        RECT 562.950 634.950 565.050 635.400 ;
        RECT 580.950 634.950 583.050 635.400 ;
        RECT 586.950 636.450 589.050 637.050 ;
        RECT 619.950 636.450 622.050 637.050 ;
        RECT 586.950 635.400 622.050 636.450 ;
        RECT 586.950 634.950 589.050 635.400 ;
        RECT 619.950 634.950 622.050 635.400 ;
        RECT 631.950 636.450 634.050 637.050 ;
        RECT 637.950 636.450 640.050 637.050 ;
        RECT 631.950 635.400 640.050 636.450 ;
        RECT 631.950 634.950 634.050 635.400 ;
        RECT 637.950 634.950 640.050 635.400 ;
        RECT 652.950 636.450 655.050 637.050 ;
        RECT 658.950 636.450 661.050 637.050 ;
        RECT 652.950 635.400 661.050 636.450 ;
        RECT 652.950 634.950 655.050 635.400 ;
        RECT 658.950 634.950 661.050 635.400 ;
        RECT 664.950 636.450 667.050 637.050 ;
        RECT 671.400 636.450 676.050 637.050 ;
        RECT 664.950 635.400 676.050 636.450 ;
        RECT 664.950 634.950 667.050 635.400 ;
        RECT 672.000 634.950 676.050 635.400 ;
        RECT 700.950 636.450 703.050 637.050 ;
        RECT 745.950 636.450 751.050 637.050 ;
        RECT 700.950 635.400 751.050 636.450 ;
        RECT 700.950 634.950 703.050 635.400 ;
        RECT 745.950 634.950 751.050 635.400 ;
        RECT 769.950 636.450 772.050 637.050 ;
        RECT 791.400 636.450 792.450 637.950 ;
        RECT 808.950 636.450 811.050 636.900 ;
        RECT 769.950 635.400 783.450 636.450 ;
        RECT 791.400 635.400 811.050 636.450 ;
        RECT 769.950 634.950 772.050 635.400 ;
        RECT 742.950 633.450 745.050 634.050 ;
        RECT 782.400 633.450 783.450 635.400 ;
        RECT 808.950 634.800 811.050 635.400 ;
        RECT 838.950 636.450 841.050 637.050 ;
        RECT 859.950 636.450 862.050 637.050 ;
        RECT 838.950 635.400 862.050 636.450 ;
        RECT 838.950 634.950 841.050 635.400 ;
        RECT 859.950 634.950 862.050 635.400 ;
        RECT 868.950 636.450 871.050 637.050 ;
        RECT 880.950 636.450 883.050 637.050 ;
        RECT 886.950 636.450 889.050 637.050 ;
        RECT 868.950 635.400 889.050 636.450 ;
        RECT 868.950 634.950 871.050 635.400 ;
        RECT 880.950 634.950 883.050 635.400 ;
        RECT 886.950 634.950 889.050 635.400 ;
        RECT 823.950 633.450 826.050 634.050 ;
        RECT 484.950 632.400 495.450 633.450 ;
        RECT 484.950 631.950 487.050 632.400 ;
        RECT 16.950 630.450 19.050 631.050 ;
        RECT 28.800 630.450 30.900 631.050 ;
        RECT 16.950 629.400 30.900 630.450 ;
        RECT 16.950 628.950 19.050 629.400 ;
        RECT 28.800 628.950 30.900 629.400 ;
        RECT 325.950 630.450 328.050 631.050 ;
        RECT 391.950 630.450 394.050 631.050 ;
        RECT 325.950 629.400 394.050 630.450 ;
        RECT 325.950 628.950 328.050 629.400 ;
        RECT 391.950 628.950 394.050 629.400 ;
        RECT 413.100 628.950 418.050 631.050 ;
        RECT 439.950 630.450 442.050 631.050 ;
        RECT 490.950 630.450 493.050 631.050 ;
        RECT 439.950 629.400 493.050 630.450 ;
        RECT 494.400 630.450 495.450 632.400 ;
        RECT 742.950 632.400 780.450 633.450 ;
        RECT 782.400 632.400 826.050 633.450 ;
        RECT 742.950 631.950 745.050 632.400 ;
        RECT 526.950 630.450 529.050 631.050 ;
        RECT 494.400 629.400 529.050 630.450 ;
        RECT 439.950 628.950 442.050 629.400 ;
        RECT 490.950 628.950 493.050 629.400 ;
        RECT 526.950 628.950 529.050 629.400 ;
        RECT 568.950 630.450 571.050 631.050 ;
        RECT 646.950 630.450 649.050 631.050 ;
        RECT 700.950 630.450 703.050 631.050 ;
        RECT 568.950 629.400 703.050 630.450 ;
        RECT 568.950 628.950 571.050 629.400 ;
        RECT 646.950 628.950 649.050 629.400 ;
        RECT 700.950 628.950 703.050 629.400 ;
        RECT 718.950 630.450 721.050 631.050 ;
        RECT 739.950 630.450 742.050 631.050 ;
        RECT 718.950 629.400 742.050 630.450 ;
        RECT 779.400 630.450 780.450 632.400 ;
        RECT 823.950 631.950 826.050 632.400 ;
        RECT 844.950 630.450 847.050 631.050 ;
        RECT 855.000 630.450 859.050 631.050 ;
        RECT 779.400 629.400 847.050 630.450 ;
        RECT 718.950 628.950 721.050 629.400 ;
        RECT 739.950 628.950 742.050 629.400 ;
        RECT 844.950 628.950 847.050 629.400 ;
        RECT 854.400 628.950 859.050 630.450 ;
        RECT 1.950 627.450 4.050 628.050 ;
        RECT 10.950 627.450 13.050 628.050 ;
        RECT 1.950 626.400 13.050 627.450 ;
        RECT 1.950 625.950 4.050 626.400 ;
        RECT 10.950 625.950 13.050 626.400 ;
        RECT 19.950 627.450 22.050 628.050 ;
        RECT 154.950 627.450 157.050 628.050 ;
        RECT 19.950 626.400 157.050 627.450 ;
        RECT 19.950 625.950 22.050 626.400 ;
        RECT 154.950 625.950 157.050 626.400 ;
        RECT 160.950 627.450 163.050 628.050 ;
        RECT 268.950 627.450 271.050 628.050 ;
        RECT 160.950 626.400 271.050 627.450 ;
        RECT 160.950 625.950 163.050 626.400 ;
        RECT 268.950 625.950 271.050 626.400 ;
        RECT 286.950 627.450 289.050 628.050 ;
        RECT 322.950 627.450 325.050 628.050 ;
        RECT 286.950 626.400 325.050 627.450 ;
        RECT 286.950 625.950 289.050 626.400 ;
        RECT 322.950 625.950 325.050 626.400 ;
        RECT 334.950 627.450 337.050 628.050 ;
        RECT 346.950 627.450 349.050 628.050 ;
        RECT 334.950 626.400 349.050 627.450 ;
        RECT 334.950 625.950 337.050 626.400 ;
        RECT 346.950 625.950 349.050 626.400 ;
        RECT 367.950 627.450 370.050 628.050 ;
        RECT 442.950 627.450 445.050 628.050 ;
        RECT 502.800 627.450 504.900 628.050 ;
        RECT 367.950 626.400 438.450 627.450 ;
        RECT 367.950 625.950 370.050 626.400 ;
        RECT 25.950 624.450 28.050 625.050 ;
        RECT 49.950 624.450 52.050 625.050 ;
        RECT 25.950 623.400 52.050 624.450 ;
        RECT 25.950 622.950 28.050 623.400 ;
        RECT 49.950 622.950 52.050 623.400 ;
        RECT 103.950 624.450 106.050 625.050 ;
        RECT 121.950 624.450 124.050 625.050 ;
        RECT 187.950 624.450 190.050 625.050 ;
        RECT 226.950 624.450 229.050 625.050 ;
        RECT 103.950 623.400 190.050 624.450 ;
        RECT 103.950 622.950 106.050 623.400 ;
        RECT 121.950 622.950 124.050 623.400 ;
        RECT 187.950 622.950 190.050 623.400 ;
        RECT 200.400 623.400 229.050 624.450 ;
        RECT 4.950 621.450 7.050 622.050 ;
        RECT 37.950 621.450 40.050 622.050 ;
        RECT 4.950 620.400 40.050 621.450 ;
        RECT 4.950 619.950 7.050 620.400 ;
        RECT 37.950 619.950 40.050 620.400 ;
        RECT 43.950 621.450 46.050 622.050 ;
        RECT 100.950 621.450 103.050 622.050 ;
        RECT 172.950 621.450 175.050 622.050 ;
        RECT 43.950 620.400 175.050 621.450 ;
        RECT 43.950 619.950 46.050 620.400 ;
        RECT 100.950 619.950 103.050 620.400 ;
        RECT 172.950 619.950 175.050 620.400 ;
        RECT 184.950 621.450 187.050 622.050 ;
        RECT 200.400 621.450 201.450 623.400 ;
        RECT 226.950 622.950 229.050 623.400 ;
        RECT 253.950 624.450 256.050 625.050 ;
        RECT 361.800 624.450 363.900 625.050 ;
        RECT 253.950 623.400 363.900 624.450 ;
        RECT 253.950 622.950 256.050 623.400 ;
        RECT 361.800 622.950 363.900 623.400 ;
        RECT 373.950 624.450 376.050 625.050 ;
        RECT 418.950 624.450 421.050 625.050 ;
        RECT 373.950 623.400 421.050 624.450 ;
        RECT 437.400 624.450 438.450 626.400 ;
        RECT 442.950 626.400 504.900 627.450 ;
        RECT 442.950 625.950 445.050 626.400 ;
        RECT 502.800 625.950 504.900 626.400 ;
        RECT 506.100 627.450 508.200 628.050 ;
        RECT 523.950 627.450 526.050 628.050 ;
        RECT 506.100 626.400 526.050 627.450 ;
        RECT 506.100 625.950 508.200 626.400 ;
        RECT 523.950 625.950 526.050 626.400 ;
        RECT 529.950 627.450 532.050 628.050 ;
        RECT 535.950 627.450 538.050 628.050 ;
        RECT 529.950 626.400 538.050 627.450 ;
        RECT 529.950 625.950 532.050 626.400 ;
        RECT 535.950 625.950 538.050 626.400 ;
        RECT 550.950 627.450 553.050 628.050 ;
        RECT 577.950 627.450 580.050 628.050 ;
        RECT 610.950 627.450 613.050 628.050 ;
        RECT 667.950 627.450 670.050 628.050 ;
        RECT 697.950 627.450 700.050 628.050 ;
        RECT 550.950 626.400 573.450 627.450 ;
        RECT 550.950 625.950 553.050 626.400 ;
        RECT 514.800 624.450 516.900 625.050 ;
        RECT 437.400 623.400 516.900 624.450 ;
        RECT 373.950 622.950 376.050 623.400 ;
        RECT 418.950 622.950 421.050 623.400 ;
        RECT 184.950 620.400 201.450 621.450 ;
        RECT 202.950 621.450 205.050 622.050 ;
        RECT 232.800 621.450 234.900 622.050 ;
        RECT 202.950 620.400 234.900 621.450 ;
        RECT 184.950 619.950 187.050 620.400 ;
        RECT 202.950 619.950 205.050 620.400 ;
        RECT 232.800 619.950 234.900 620.400 ;
        RECT 236.100 621.450 238.200 622.050 ;
        RECT 265.950 621.450 268.050 622.050 ;
        RECT 236.100 620.400 268.050 621.450 ;
        RECT 236.100 619.950 238.200 620.400 ;
        RECT 265.950 619.950 268.050 620.400 ;
        RECT 280.950 621.450 283.050 622.050 ;
        RECT 346.950 621.450 349.050 622.050 ;
        RECT 373.950 621.450 376.050 622.050 ;
        RECT 280.950 620.400 349.050 621.450 ;
        RECT 280.950 619.950 283.050 620.400 ;
        RECT 346.950 619.950 349.050 620.400 ;
        RECT 350.400 620.400 376.050 621.450 ;
        RECT 73.950 618.450 76.050 619.050 ;
        RECT 91.950 618.450 94.050 619.050 ;
        RECT 73.950 617.400 94.050 618.450 ;
        RECT 127.950 618.450 130.050 619.050 ;
        RECT 139.950 618.450 142.050 619.050 ;
        RECT 127.950 617.400 142.050 618.450 ;
        RECT 205.950 618.450 208.050 619.050 ;
        RECT 229.950 618.450 232.050 619.050 ;
        RECT 205.950 617.400 232.050 618.450 ;
        RECT 73.950 616.950 76.050 617.400 ;
        RECT 91.950 616.950 94.050 617.400 ;
        RECT 97.950 615.300 100.050 617.400 ;
        RECT 127.950 616.950 130.050 617.400 ;
        RECT 139.950 616.950 142.050 617.400 ;
        RECT 98.850 611.700 100.050 615.300 ;
        RECT 118.950 614.400 121.050 616.500 ;
        RECT 133.950 615.450 136.050 616.050 ;
        RECT 148.950 615.450 151.050 616.050 ;
        RECT 133.950 614.400 151.050 615.450 ;
        RECT 157.950 614.400 160.050 616.500 ;
        RECT 178.950 615.300 181.050 617.400 ;
        RECT 205.950 616.950 208.050 617.400 ;
        RECT 229.950 616.950 232.050 617.400 ;
        RECT 271.950 618.450 274.050 619.050 ;
        RECT 310.800 618.450 312.900 619.050 ;
        RECT 271.950 617.400 312.900 618.450 ;
        RECT 271.950 616.950 274.050 617.400 ;
        RECT 310.800 616.950 312.900 617.400 ;
        RECT 314.100 618.450 316.200 619.050 ;
        RECT 334.950 618.450 337.050 619.050 ;
        RECT 314.100 617.400 337.050 618.450 ;
        RECT 314.100 616.950 316.200 617.400 ;
        RECT 334.950 616.950 337.050 617.400 ;
        RECT 343.950 618.450 346.050 619.050 ;
        RECT 350.400 618.450 351.450 620.400 ;
        RECT 373.950 619.950 376.050 620.400 ;
        RECT 385.950 621.450 388.050 622.050 ;
        RECT 415.950 621.450 418.050 622.050 ;
        RECT 457.950 621.450 460.050 622.050 ;
        RECT 385.950 620.400 460.050 621.450 ;
        RECT 385.950 619.950 388.050 620.400 ;
        RECT 415.950 619.950 418.050 620.400 ;
        RECT 457.950 619.950 460.050 620.400 ;
        RECT 496.950 619.950 499.050 623.400 ;
        RECT 514.800 622.950 516.900 623.400 ;
        RECT 518.100 624.450 520.200 625.050 ;
        RECT 568.950 624.450 571.050 625.050 ;
        RECT 518.100 623.400 571.050 624.450 ;
        RECT 572.400 624.450 573.450 626.400 ;
        RECT 577.950 626.400 700.050 627.450 ;
        RECT 577.950 625.950 580.050 626.400 ;
        RECT 610.950 625.950 613.050 626.400 ;
        RECT 667.950 625.950 670.050 626.400 ;
        RECT 697.950 625.950 700.050 626.400 ;
        RECT 703.950 627.450 706.050 628.050 ;
        RECT 733.950 627.450 736.050 628.050 ;
        RECT 703.950 626.400 736.050 627.450 ;
        RECT 703.950 625.950 706.050 626.400 ;
        RECT 733.950 625.950 736.050 626.400 ;
        RECT 781.950 627.450 784.050 628.050 ;
        RECT 841.950 627.450 844.050 628.050 ;
        RECT 854.400 627.450 855.450 628.950 ;
        RECT 781.950 626.400 819.450 627.450 ;
        RECT 781.950 625.950 784.050 626.400 ;
        RECT 818.400 625.050 819.450 626.400 ;
        RECT 841.950 626.400 855.450 627.450 ;
        RECT 856.950 627.450 859.050 628.050 ;
        RECT 880.950 627.450 883.050 628.050 ;
        RECT 856.950 626.400 883.050 627.450 ;
        RECT 841.950 625.950 844.050 626.400 ;
        RECT 856.950 625.950 859.050 626.400 ;
        RECT 880.950 625.950 883.050 626.400 ;
        RECT 910.950 625.050 913.050 625.200 ;
        RECT 724.950 624.450 727.050 625.050 ;
        RECT 817.950 624.450 820.050 625.050 ;
        RECT 826.950 624.450 829.050 625.050 ;
        RECT 572.400 623.400 600.450 624.450 ;
        RECT 518.100 622.950 520.200 623.400 ;
        RECT 568.950 622.950 571.050 623.400 ;
        RECT 505.950 621.450 508.050 622.050 ;
        RECT 520.950 621.450 523.050 622.050 ;
        RECT 505.950 620.400 523.050 621.450 ;
        RECT 505.950 619.950 508.050 620.400 ;
        RECT 520.950 619.950 523.050 620.400 ;
        RECT 532.950 621.450 535.050 622.050 ;
        RECT 544.950 621.450 547.050 622.050 ;
        RECT 532.950 620.400 547.050 621.450 ;
        RECT 599.400 621.450 600.450 623.400 ;
        RECT 724.950 623.400 783.450 624.450 ;
        RECT 724.950 622.950 727.050 623.400 ;
        RECT 769.950 621.450 772.050 622.050 ;
        RECT 599.400 620.400 772.050 621.450 ;
        RECT 782.400 621.450 783.450 623.400 ;
        RECT 817.950 623.400 829.050 624.450 ;
        RECT 817.950 622.950 820.050 623.400 ;
        RECT 826.950 622.950 829.050 623.400 ;
        RECT 835.950 624.450 838.050 625.050 ;
        RECT 847.800 624.450 849.900 625.050 ;
        RECT 835.950 623.400 849.900 624.450 ;
        RECT 835.950 622.950 838.050 623.400 ;
        RECT 847.800 622.950 849.900 623.400 ;
        RECT 851.100 624.450 853.200 625.050 ;
        RECT 859.950 624.450 862.050 625.050 ;
        RECT 851.100 623.400 862.050 624.450 ;
        RECT 851.100 622.950 853.200 623.400 ;
        RECT 859.950 622.950 862.050 623.400 ;
        RECT 895.950 624.450 898.050 625.050 ;
        RECT 901.950 624.450 904.050 625.050 ;
        RECT 895.950 623.400 904.050 624.450 ;
        RECT 895.950 622.950 898.050 623.400 ;
        RECT 901.950 622.950 904.050 623.400 ;
        RECT 910.950 624.450 915.000 625.050 ;
        RECT 910.950 623.100 915.450 624.450 ;
        RECT 912.000 622.950 915.450 623.100 ;
        RECT 790.800 621.450 792.900 622.050 ;
        RECT 782.400 620.400 792.900 621.450 ;
        RECT 532.950 619.950 535.050 620.400 ;
        RECT 544.950 619.950 547.050 620.400 ;
        RECT 769.950 619.950 772.050 620.400 ;
        RECT 790.800 619.950 792.900 620.400 ;
        RECT 794.100 621.450 796.200 622.050 ;
        RECT 811.950 621.450 814.050 622.050 ;
        RECT 794.100 620.400 814.050 621.450 ;
        RECT 794.100 619.950 796.200 620.400 ;
        RECT 811.950 619.950 814.050 620.400 ;
        RECT 358.950 618.450 361.050 619.050 ;
        RECT 343.950 617.400 351.450 618.450 ;
        RECT 353.400 617.400 361.050 618.450 ;
        RECT 484.950 618.450 487.050 619.050 ;
        RECT 499.950 618.450 502.050 619.050 ;
        RECT 484.950 617.400 502.050 618.450 ;
        RECT 562.950 618.450 565.050 619.050 ;
        RECT 577.950 618.450 580.050 619.050 ;
        RECT 562.950 617.400 580.050 618.450 ;
        RECT 343.950 616.950 346.050 617.400 ;
        RECT 184.950 615.450 187.050 616.050 ;
        RECT 211.950 615.450 214.050 616.050 ;
        RECT 13.950 607.950 16.050 610.050 ;
        RECT 19.950 607.950 22.050 610.050 ;
        RECT 37.950 607.950 40.050 610.050 ;
        RECT 43.950 607.950 46.050 610.050 ;
        RECT 64.950 607.950 67.050 610.050 ;
        RECT 79.950 607.950 82.050 610.050 ;
        RECT 85.950 607.950 88.050 610.050 ;
        RECT 97.950 609.600 100.050 611.700 ;
        RECT 13.950 604.950 16.050 606.750 ;
        RECT 19.950 604.950 22.050 606.750 ;
        RECT 37.950 604.950 40.050 606.750 ;
        RECT 43.950 604.950 46.050 606.750 ;
        RECT 58.950 604.950 61.050 606.750 ;
        RECT 64.950 604.950 67.050 606.750 ;
        RECT 16.950 602.250 19.050 604.050 ;
        RECT 34.950 602.250 37.050 604.050 ;
        RECT 40.950 602.250 43.050 604.050 ;
        RECT 61.950 602.250 64.050 604.050 ;
        RECT 70.950 601.950 73.050 607.050 ;
        RECT 79.950 604.950 82.050 606.750 ;
        RECT 85.950 604.950 88.050 606.750 ;
        RECT 82.950 602.250 85.050 604.050 ;
        RECT 88.950 602.250 91.050 604.050 ;
        RECT 94.950 602.250 97.050 604.050 ;
        RECT 16.950 598.950 19.050 601.050 ;
        RECT 34.950 595.950 37.050 601.050 ;
        RECT 40.950 598.950 43.050 601.050 ;
        RECT 61.950 600.450 64.050 601.050 ;
        RECT 73.800 600.450 75.900 601.050 ;
        RECT 61.950 599.400 75.900 600.450 ;
        RECT 61.950 598.950 64.050 599.400 ;
        RECT 73.800 598.950 75.900 599.400 ;
        RECT 77.100 600.450 81.000 601.050 ;
        RECT 82.950 600.450 85.050 601.050 ;
        RECT 77.100 599.400 85.050 600.450 ;
        RECT 77.100 598.950 81.000 599.400 ;
        RECT 82.950 598.950 85.050 599.400 ;
        RECT 88.950 598.950 91.050 601.050 ;
        RECT 94.950 598.950 97.050 601.050 ;
        RECT 16.950 594.450 19.050 595.050 ;
        RECT 46.950 594.450 49.050 595.050 ;
        RECT 16.950 593.400 49.050 594.450 ;
        RECT 16.950 592.950 19.050 593.400 ;
        RECT 46.950 592.950 49.050 593.400 ;
        RECT 49.950 591.450 52.050 592.050 ;
        RECT 55.950 591.450 58.050 592.050 ;
        RECT 49.950 590.400 58.050 591.450 ;
        RECT 49.950 589.950 52.050 590.400 ;
        RECT 55.950 589.950 58.050 590.400 ;
        RECT 70.950 589.950 73.050 595.050 ;
        RECT 98.850 594.600 100.050 609.600 ;
        RECT 112.950 604.950 115.050 607.050 ;
        RECT 112.950 601.950 115.050 603.750 ;
        RECT 119.100 594.600 120.300 614.400 ;
        RECT 133.950 613.950 136.050 614.400 ;
        RECT 148.950 613.950 151.050 614.400 ;
        RECT 121.950 612.450 124.050 613.050 ;
        RECT 127.950 612.450 130.050 613.050 ;
        RECT 151.950 612.450 154.050 613.050 ;
        RECT 121.950 611.400 130.050 612.450 ;
        RECT 121.950 610.950 124.050 611.400 ;
        RECT 127.950 610.950 130.050 611.400 ;
        RECT 145.950 611.400 154.050 612.450 ;
        RECT 139.950 607.950 142.050 610.050 ;
        RECT 145.950 607.950 148.050 611.400 ;
        RECT 151.950 610.950 154.050 611.400 ;
        RECT 121.950 606.450 124.050 607.050 ;
        RECT 126.000 606.450 130.050 607.050 ;
        RECT 121.950 605.400 130.050 606.450 ;
        RECT 121.950 604.950 124.050 605.400 ;
        RECT 126.000 604.950 130.050 605.400 ;
        RECT 139.950 604.950 142.050 606.750 ;
        RECT 145.950 604.950 148.050 606.750 ;
        RECT 154.950 604.950 157.050 607.050 ;
        RECT 121.950 601.950 124.050 603.750 ;
        RECT 142.950 602.250 145.050 604.050 ;
        RECT 148.950 602.250 151.050 604.050 ;
        RECT 154.950 601.950 157.050 603.750 ;
        RECT 127.950 600.450 130.050 601.050 ;
        RECT 142.950 600.450 145.050 601.050 ;
        RECT 127.950 599.400 145.050 600.450 ;
        RECT 127.950 598.950 130.050 599.400 ;
        RECT 142.950 598.950 145.050 599.400 ;
        RECT 148.950 598.950 151.050 601.050 ;
        RECT 97.950 592.500 100.050 594.600 ;
        RECT 118.950 592.500 121.050 594.600 ;
        RECT 139.950 594.450 142.050 595.050 ;
        RECT 145.950 594.450 148.050 595.050 ;
        RECT 158.700 594.600 159.900 614.400 ;
        RECT 178.950 611.700 180.150 615.300 ;
        RECT 184.950 614.400 214.050 615.450 ;
        RECT 184.950 613.950 187.050 614.400 ;
        RECT 211.950 613.950 214.050 614.400 ;
        RECT 256.950 615.450 259.050 616.050 ;
        RECT 304.950 615.450 307.050 616.050 ;
        RECT 256.950 614.400 307.050 615.450 ;
        RECT 256.950 613.950 259.050 614.400 ;
        RECT 304.950 613.950 307.050 614.400 ;
        RECT 319.950 615.450 322.050 616.050 ;
        RECT 325.800 615.450 327.900 616.050 ;
        RECT 319.950 614.400 327.900 615.450 ;
        RECT 319.950 613.950 322.050 614.400 ;
        RECT 325.800 613.950 327.900 614.400 ;
        RECT 329.100 615.450 331.200 616.050 ;
        RECT 340.950 615.450 343.050 616.050 ;
        RECT 353.400 615.450 354.450 617.400 ;
        RECT 358.950 616.950 361.050 617.400 ;
        RECT 373.950 615.450 376.050 616.050 ;
        RECT 329.100 614.400 354.450 615.450 ;
        RECT 356.400 614.400 376.050 615.450 ;
        RECT 329.100 613.950 331.200 614.400 ;
        RECT 340.950 613.950 343.050 614.400 ;
        RECT 346.950 612.450 349.050 613.050 ;
        RECT 356.400 612.450 357.450 614.400 ;
        RECT 373.950 613.950 376.050 614.400 ;
        RECT 391.950 615.450 394.050 616.050 ;
        RECT 409.950 615.450 412.050 616.050 ;
        RECT 391.950 614.400 412.050 615.450 ;
        RECT 424.950 614.400 427.050 616.500 ;
        RECT 445.950 615.300 448.050 617.400 ;
        RECT 484.950 616.950 487.050 617.400 ;
        RECT 499.950 616.950 502.050 617.400 ;
        RECT 454.950 615.450 457.050 616.050 ;
        RECT 463.950 615.450 466.050 616.050 ;
        RECT 391.950 613.950 394.050 614.400 ;
        RECT 409.950 613.950 412.050 614.400 ;
        RECT 178.950 609.600 181.050 611.700 ;
        RECT 346.950 611.400 357.450 612.450 ;
        RECT 346.950 610.950 349.050 611.400 ;
        RECT 163.950 604.950 166.050 607.050 ;
        RECT 163.950 601.950 166.050 603.750 ;
        RECT 178.950 594.600 180.150 609.600 ;
        RECT 199.950 607.950 202.050 610.050 ;
        RECT 205.950 607.950 208.050 610.050 ;
        RECT 220.950 607.950 223.050 610.050 ;
        RECT 247.950 607.950 250.050 610.050 ;
        RECT 268.950 607.950 271.050 610.050 ;
        RECT 313.950 607.950 316.050 610.050 ;
        RECT 319.950 607.950 322.050 610.050 ;
        RECT 334.950 607.950 337.050 610.050 ;
        RECT 340.950 607.950 343.050 610.050 ;
        RECT 358.950 607.950 361.050 610.050 ;
        RECT 364.950 607.950 367.050 610.050 ;
        RECT 385.950 607.950 388.050 610.050 ;
        RECT 391.950 607.950 394.050 610.050 ;
        RECT 406.950 607.950 412.050 610.050 ;
        RECT 415.950 607.950 418.050 610.050 ;
        RECT 199.950 604.950 202.050 606.750 ;
        RECT 205.950 604.950 208.050 606.750 ;
        RECT 220.950 604.950 223.050 606.750 ;
        RECT 226.950 604.950 229.050 606.750 ;
        RECT 241.950 604.950 244.050 606.750 ;
        RECT 247.950 604.950 250.050 606.750 ;
        RECT 262.950 604.950 265.050 606.750 ;
        RECT 268.950 604.950 271.050 606.750 ;
        RECT 283.950 604.950 286.050 607.050 ;
        RECT 292.950 604.950 298.050 607.050 ;
        RECT 313.950 604.950 316.050 606.750 ;
        RECT 319.950 604.950 322.050 606.750 ;
        RECT 334.950 604.950 337.050 606.750 ;
        RECT 340.950 604.950 343.050 606.750 ;
        RECT 358.950 604.950 361.050 606.750 ;
        RECT 364.950 604.950 367.050 606.750 ;
        RECT 385.950 604.950 388.050 606.750 ;
        RECT 391.950 604.950 394.050 606.750 ;
        RECT 409.950 604.950 412.050 606.750 ;
        RECT 415.950 604.950 418.050 606.750 ;
        RECT 421.950 604.950 424.050 607.050 ;
        RECT 181.950 602.250 184.050 604.050 ;
        RECT 202.950 602.250 205.050 604.050 ;
        RECT 208.950 602.250 211.050 604.050 ;
        RECT 223.950 602.250 226.050 604.050 ;
        RECT 244.950 602.250 247.050 604.050 ;
        RECT 265.950 602.250 268.050 604.050 ;
        RECT 289.950 603.750 291.750 604.050 ;
        RECT 283.950 601.950 286.050 603.750 ;
        RECT 289.950 602.250 292.050 603.750 ;
        RECT 292.950 602.250 295.050 603.750 ;
        RECT 310.950 602.250 313.050 604.050 ;
        RECT 316.950 602.250 319.050 604.050 ;
        RECT 337.950 602.250 340.050 604.050 ;
        RECT 343.950 602.250 346.050 604.050 ;
        RECT 355.950 602.250 358.050 604.050 ;
        RECT 361.950 602.250 364.050 604.050 ;
        RECT 382.950 602.250 385.050 604.050 ;
        RECT 388.950 602.250 391.050 604.050 ;
        RECT 406.950 602.250 409.050 604.050 ;
        RECT 412.950 602.250 415.050 604.050 ;
        RECT 293.250 601.950 295.050 602.250 ;
        RECT 421.950 601.950 424.050 603.750 ;
        RECT 181.950 598.950 184.050 601.050 ;
        RECT 202.950 595.950 205.050 601.050 ;
        RECT 208.950 598.950 211.050 601.050 ;
        RECT 223.950 598.950 226.050 601.050 ;
        RECT 244.950 600.450 247.050 601.050 ;
        RECT 256.950 600.450 259.050 601.050 ;
        RECT 244.950 599.400 259.050 600.450 ;
        RECT 244.950 598.950 247.050 599.400 ;
        RECT 256.950 598.950 259.050 599.400 ;
        RECT 265.950 600.450 268.050 601.050 ;
        RECT 280.950 600.450 283.050 601.050 ;
        RECT 265.950 599.400 283.050 600.450 ;
        RECT 265.950 598.950 268.050 599.400 ;
        RECT 280.950 598.950 283.050 599.400 ;
        RECT 301.950 600.450 304.050 601.050 ;
        RECT 310.950 600.450 313.050 601.050 ;
        RECT 301.950 599.400 313.050 600.450 ;
        RECT 301.950 598.950 304.050 599.400 ;
        RECT 310.950 598.950 313.050 599.400 ;
        RECT 316.950 598.950 319.050 601.050 ;
        RECT 139.950 593.400 148.050 594.450 ;
        RECT 139.950 592.950 142.050 593.400 ;
        RECT 145.950 592.950 148.050 593.400 ;
        RECT 157.950 592.500 160.050 594.600 ;
        RECT 178.950 592.500 181.050 594.600 ;
        RECT 199.950 594.450 202.050 595.050 ;
        RECT 224.400 594.450 225.450 598.950 ;
        RECT 337.950 595.950 340.050 601.050 ;
        RECT 343.950 600.450 346.050 601.050 ;
        RECT 348.000 600.450 352.050 601.050 ;
        RECT 343.950 599.400 352.050 600.450 ;
        RECT 343.950 598.950 346.050 599.400 ;
        RECT 348.000 598.950 352.050 599.400 ;
        RECT 355.950 598.950 358.050 601.050 ;
        RECT 361.950 598.950 364.050 601.050 ;
        RECT 370.950 600.450 373.050 601.050 ;
        RECT 382.950 600.450 385.050 601.050 ;
        RECT 370.950 599.400 385.050 600.450 ;
        RECT 370.950 598.950 373.050 599.400 ;
        RECT 382.950 598.950 385.050 599.400 ;
        RECT 388.950 598.950 391.050 601.050 ;
        RECT 406.950 598.950 409.050 601.050 ;
        RECT 412.950 598.950 415.050 601.050 ;
        RECT 199.950 593.400 225.450 594.450 ;
        RECT 247.950 594.450 250.050 595.050 ;
        RECT 268.950 594.450 271.050 595.050 ;
        RECT 247.950 593.400 271.050 594.450 ;
        RECT 199.950 592.950 202.050 593.400 ;
        RECT 247.950 592.950 250.050 593.400 ;
        RECT 268.950 592.950 271.050 593.400 ;
        RECT 304.950 594.450 307.050 595.050 ;
        RECT 362.400 594.450 363.450 598.950 ;
        RECT 304.950 593.400 363.450 594.450 ;
        RECT 373.950 594.450 376.050 595.050 ;
        RECT 407.400 594.450 408.450 598.950 ;
        RECT 425.700 594.600 426.900 614.400 ;
        RECT 445.950 611.700 447.150 615.300 ;
        RECT 454.950 614.400 466.050 615.450 ;
        RECT 454.950 613.950 457.050 614.400 ;
        RECT 463.950 613.950 466.050 614.400 ;
        RECT 469.950 615.450 472.050 616.050 ;
        RECT 478.950 615.450 481.050 616.050 ;
        RECT 469.950 614.400 481.050 615.450 ;
        RECT 508.950 614.400 511.050 616.500 ;
        RECT 529.950 615.300 532.050 617.400 ;
        RECT 562.950 616.950 565.050 617.400 ;
        RECT 577.950 616.950 580.050 617.400 ;
        RECT 592.950 618.450 595.050 619.050 ;
        RECT 664.950 618.450 667.050 619.050 ;
        RECT 592.950 617.400 667.050 618.450 ;
        RECT 592.950 616.950 595.050 617.400 ;
        RECT 664.950 616.950 667.050 617.400 ;
        RECT 706.950 618.450 709.050 619.050 ;
        RECT 715.950 618.450 718.050 619.050 ;
        RECT 706.950 617.400 718.050 618.450 ;
        RECT 706.950 616.950 709.050 617.400 ;
        RECT 715.950 616.950 718.050 617.400 ;
        RECT 766.950 618.450 769.050 619.050 ;
        RECT 772.950 618.450 775.050 619.050 ;
        RECT 814.950 618.450 817.050 619.050 ;
        RECT 766.950 617.400 775.050 618.450 ;
        RECT 766.950 616.950 769.050 617.400 ;
        RECT 772.950 616.950 775.050 617.400 ;
        RECT 806.400 617.400 817.050 618.450 ;
        RECT 559.950 615.450 562.050 616.050 ;
        RECT 568.950 615.450 571.050 616.050 ;
        RECT 469.950 613.950 472.050 614.400 ;
        RECT 478.950 613.950 481.050 614.400 ;
        RECT 445.950 609.600 448.050 611.700 ;
        RECT 430.950 604.950 436.050 607.050 ;
        RECT 430.950 601.950 433.050 603.750 ;
        RECT 445.950 594.600 447.150 609.600 ;
        RECT 463.950 607.950 466.050 610.050 ;
        RECT 469.950 607.950 472.050 610.050 ;
        RECT 490.950 607.950 493.050 610.050 ;
        RECT 496.950 607.950 499.050 610.050 ;
        RECT 463.950 604.950 466.050 606.750 ;
        RECT 469.950 604.950 472.050 606.750 ;
        RECT 490.950 604.950 493.050 606.750 ;
        RECT 496.950 604.950 499.050 606.750 ;
        RECT 505.950 604.950 508.050 607.050 ;
        RECT 448.950 602.250 451.050 604.050 ;
        RECT 466.950 602.250 469.050 604.050 ;
        RECT 472.950 602.250 475.050 604.050 ;
        RECT 493.950 602.250 496.050 604.050 ;
        RECT 499.950 602.250 502.050 604.050 ;
        RECT 505.950 601.950 508.050 603.750 ;
        RECT 448.950 598.950 451.050 601.050 ;
        RECT 466.950 598.950 469.050 601.050 ;
        RECT 472.950 598.950 478.050 601.050 ;
        RECT 493.950 598.950 496.050 601.050 ;
        RECT 499.950 598.950 502.050 601.050 ;
        RECT 373.950 593.400 408.450 594.450 ;
        RECT 304.950 592.950 307.050 593.400 ;
        RECT 373.950 592.950 376.050 593.400 ;
        RECT 424.950 592.500 427.050 594.600 ;
        RECT 445.950 592.500 448.050 594.600 ;
        RECT 457.950 594.450 460.050 595.050 ;
        RECT 466.950 594.450 469.050 595.050 ;
        RECT 457.950 593.400 469.050 594.450 ;
        RECT 457.950 592.950 460.050 593.400 ;
        RECT 466.950 592.950 469.050 593.400 ;
        RECT 493.950 594.450 496.050 595.050 ;
        RECT 502.950 594.450 505.050 595.050 ;
        RECT 509.700 594.600 510.900 614.400 ;
        RECT 529.950 611.700 531.150 615.300 ;
        RECT 559.950 614.400 571.050 615.450 ;
        RECT 559.950 613.950 562.050 614.400 ;
        RECT 568.950 613.950 571.050 614.400 ;
        RECT 616.950 615.450 619.050 616.050 ;
        RECT 622.950 615.450 625.050 616.050 ;
        RECT 616.950 614.400 625.050 615.450 ;
        RECT 616.950 613.950 619.050 614.400 ;
        RECT 622.950 613.950 625.050 614.400 ;
        RECT 634.950 615.450 637.050 616.050 ;
        RECT 655.950 615.450 658.050 616.050 ;
        RECT 806.400 615.450 807.450 617.400 ;
        RECT 814.950 616.950 817.050 617.400 ;
        RECT 838.950 616.950 841.050 622.050 ;
        RECT 886.950 621.450 889.050 622.050 ;
        RECT 898.950 621.450 901.050 622.050 ;
        RECT 886.950 620.400 901.050 621.450 ;
        RECT 886.950 619.950 889.050 620.400 ;
        RECT 898.950 619.950 901.050 620.400 ;
        RECT 904.950 621.450 907.050 622.200 ;
        RECT 910.950 621.450 913.050 621.900 ;
        RECT 904.950 620.400 913.050 621.450 ;
        RECT 904.950 620.100 907.050 620.400 ;
        RECT 910.950 619.800 913.050 620.400 ;
        RECT 847.950 618.450 850.050 619.050 ;
        RECT 853.950 618.450 856.050 619.050 ;
        RECT 847.950 617.400 856.050 618.450 ;
        RECT 847.950 616.950 850.050 617.400 ;
        RECT 853.950 616.950 856.050 617.400 ;
        RECT 904.950 618.450 907.050 618.900 ;
        RECT 914.400 618.450 915.450 622.950 ;
        RECT 904.950 617.400 915.450 618.450 ;
        RECT 904.950 616.800 907.050 617.400 ;
        RECT 634.950 614.400 658.050 615.450 ;
        RECT 634.950 613.950 637.050 614.400 ;
        RECT 655.950 613.950 658.050 614.400 ;
        RECT 770.400 614.400 807.450 615.450 ;
        RECT 808.950 615.450 811.050 616.050 ;
        RECT 817.950 615.450 820.050 616.050 ;
        RECT 808.950 614.400 820.050 615.450 ;
        RECT 770.400 613.050 771.450 614.400 ;
        RECT 808.950 613.950 811.050 614.400 ;
        RECT 817.950 613.950 820.050 614.400 ;
        RECT 865.950 615.450 868.050 616.050 ;
        RECT 874.950 615.450 877.050 616.050 ;
        RECT 898.950 615.450 901.050 616.050 ;
        RECT 865.950 614.400 901.050 615.450 ;
        RECT 865.950 613.950 868.050 614.400 ;
        RECT 874.950 613.950 877.050 614.400 ;
        RECT 898.950 613.950 901.050 614.400 ;
        RECT 697.950 612.450 700.050 613.050 ;
        RECT 529.950 609.600 532.050 611.700 ;
        RECT 697.950 611.400 715.050 612.450 ;
        RECT 697.950 610.950 700.050 611.400 ;
        RECT 514.950 604.950 517.050 607.050 ;
        RECT 514.950 601.950 517.050 603.750 ;
        RECT 529.950 594.600 531.150 609.600 ;
        RECT 553.950 607.950 556.050 610.050 ;
        RECT 559.950 607.950 562.050 610.050 ;
        RECT 577.950 607.950 580.050 610.050 ;
        RECT 583.950 607.950 586.050 610.050 ;
        RECT 598.950 607.950 601.050 610.050 ;
        RECT 604.950 607.950 607.050 610.050 ;
        RECT 622.950 607.950 625.050 610.050 ;
        RECT 628.950 607.950 631.050 610.050 ;
        RECT 646.950 607.950 649.050 610.050 ;
        RECT 652.950 607.950 655.050 610.050 ;
        RECT 664.950 607.950 667.050 610.050 ;
        RECT 670.950 607.950 673.050 610.050 ;
        RECT 688.950 607.950 691.050 610.050 ;
        RECT 694.950 607.950 697.050 610.050 ;
        RECT 712.950 607.950 715.050 611.400 ;
        RECT 766.950 611.400 771.450 613.050 ;
        RECT 790.950 612.450 793.050 613.050 ;
        RECT 799.950 612.450 802.050 613.050 ;
        RECT 790.950 611.400 802.050 612.450 ;
        RECT 766.950 610.950 771.000 611.400 ;
        RECT 790.950 610.950 793.050 611.400 ;
        RECT 799.950 610.950 802.050 611.400 ;
        RECT 718.950 607.950 721.050 610.050 ;
        RECT 733.950 607.950 736.050 610.050 ;
        RECT 739.950 607.950 742.050 610.050 ;
        RECT 754.950 607.950 757.050 610.050 ;
        RECT 778.950 607.950 781.050 610.050 ;
        RECT 784.950 607.950 787.050 610.050 ;
        RECT 802.950 607.950 805.050 610.050 ;
        RECT 808.950 607.950 811.050 610.050 ;
        RECT 814.950 609.450 817.050 610.050 ;
        RECT 826.950 609.450 829.050 610.050 ;
        RECT 814.950 608.400 829.050 609.450 ;
        RECT 814.950 607.950 817.050 608.400 ;
        RECT 826.950 607.950 829.050 608.400 ;
        RECT 832.950 607.950 835.050 610.050 ;
        RECT 847.950 607.950 850.050 610.050 ;
        RECT 853.950 607.950 856.050 610.050 ;
        RECT 874.950 607.950 877.050 610.050 ;
        RECT 880.950 607.950 886.050 610.050 ;
        RECT 892.950 607.950 895.050 610.050 ;
        RECT 898.950 607.950 901.050 610.050 ;
        RECT 553.950 604.950 556.050 606.750 ;
        RECT 559.950 604.950 562.050 606.750 ;
        RECT 577.950 604.950 580.050 606.750 ;
        RECT 583.950 604.950 586.050 606.750 ;
        RECT 598.950 604.950 601.050 606.750 ;
        RECT 604.950 604.950 607.050 606.750 ;
        RECT 622.950 604.950 625.050 606.750 ;
        RECT 628.950 604.950 631.050 606.750 ;
        RECT 646.950 604.950 649.050 606.750 ;
        RECT 652.950 604.950 655.050 606.750 ;
        RECT 664.950 604.950 667.050 606.750 ;
        RECT 670.950 604.950 673.050 606.750 ;
        RECT 688.950 604.950 691.050 606.750 ;
        RECT 694.950 604.950 697.050 606.750 ;
        RECT 712.950 604.950 715.050 606.750 ;
        RECT 718.950 604.950 721.050 606.750 ;
        RECT 733.950 604.950 736.050 606.750 ;
        RECT 739.950 604.950 742.050 606.750 ;
        RECT 754.950 604.950 757.050 606.750 ;
        RECT 760.950 604.950 763.050 606.750 ;
        RECT 778.950 604.950 781.050 606.750 ;
        RECT 784.950 604.950 787.050 606.750 ;
        RECT 802.950 604.950 805.050 606.750 ;
        RECT 808.950 604.950 811.050 606.750 ;
        RECT 826.950 604.950 829.050 606.750 ;
        RECT 832.950 604.950 835.050 606.750 ;
        RECT 847.950 604.950 850.050 606.750 ;
        RECT 853.950 604.950 856.050 606.750 ;
        RECT 874.950 604.950 877.050 606.750 ;
        RECT 880.950 604.950 883.050 606.750 ;
        RECT 892.950 604.950 895.050 606.750 ;
        RECT 898.950 604.950 901.050 606.750 ;
        RECT 532.950 602.250 535.050 604.050 ;
        RECT 550.950 602.250 553.050 604.050 ;
        RECT 556.950 602.250 559.050 604.050 ;
        RECT 574.950 602.250 577.050 604.050 ;
        RECT 580.950 602.250 583.050 604.050 ;
        RECT 601.950 602.250 604.050 604.050 ;
        RECT 607.950 602.250 610.050 604.050 ;
        RECT 625.950 602.250 628.050 604.050 ;
        RECT 643.950 602.250 646.050 604.050 ;
        RECT 649.950 602.250 652.050 604.050 ;
        RECT 667.950 602.250 670.050 604.050 ;
        RECT 691.950 602.250 694.050 604.050 ;
        RECT 697.950 602.250 700.050 604.050 ;
        RECT 709.950 602.250 712.050 604.050 ;
        RECT 715.950 602.250 718.050 604.050 ;
        RECT 736.950 602.250 739.050 604.050 ;
        RECT 757.950 602.250 760.050 604.050 ;
        RECT 775.950 602.250 778.050 604.050 ;
        RECT 781.950 602.250 784.050 604.050 ;
        RECT 532.950 598.950 535.050 601.050 ;
        RECT 538.950 600.450 541.050 601.050 ;
        RECT 550.950 600.450 553.050 601.050 ;
        RECT 538.950 599.400 553.050 600.450 ;
        RECT 538.950 598.950 541.050 599.400 ;
        RECT 550.950 598.950 553.050 599.400 ;
        RECT 556.950 598.950 559.050 601.050 ;
        RECT 574.950 595.950 577.050 601.050 ;
        RECT 580.950 598.950 583.050 601.050 ;
        RECT 601.950 595.950 604.050 601.050 ;
        RECT 607.950 598.950 610.050 601.050 ;
        RECT 625.950 598.950 628.050 601.050 ;
        RECT 631.950 600.450 634.050 601.050 ;
        RECT 643.950 600.450 646.050 601.050 ;
        RECT 631.950 599.400 646.050 600.450 ;
        RECT 631.950 598.950 634.050 599.400 ;
        RECT 643.950 598.950 646.050 599.400 ;
        RECT 649.950 598.950 652.050 601.050 ;
        RECT 667.950 598.950 670.050 601.050 ;
        RECT 673.950 600.450 676.050 601.050 ;
        RECT 691.950 600.450 694.050 601.050 ;
        RECT 673.950 599.400 694.050 600.450 ;
        RECT 673.950 598.950 676.050 599.400 ;
        RECT 691.950 598.950 694.050 599.400 ;
        RECT 697.950 598.950 700.050 601.050 ;
        RECT 709.950 598.950 712.050 601.050 ;
        RECT 493.950 593.400 505.050 594.450 ;
        RECT 493.950 592.950 496.050 593.400 ;
        RECT 502.950 592.950 505.050 593.400 ;
        RECT 508.950 592.500 511.050 594.600 ;
        RECT 529.950 592.500 532.050 594.600 ;
        RECT 553.950 594.450 556.050 595.050 ;
        RECT 586.950 594.450 589.050 595.050 ;
        RECT 607.950 594.450 610.050 595.050 ;
        RECT 626.400 594.450 627.450 598.950 ;
        RECT 553.950 593.400 627.450 594.450 ;
        RECT 646.950 594.450 649.050 595.050 ;
        RECT 668.400 594.450 669.450 598.950 ;
        RECT 715.950 595.950 718.050 601.050 ;
        RECT 736.950 595.950 739.050 601.050 ;
        RECT 757.950 600.450 760.050 601.050 ;
        RECT 769.950 600.450 772.050 601.050 ;
        RECT 757.950 599.400 772.050 600.450 ;
        RECT 757.950 598.950 760.050 599.400 ;
        RECT 769.950 598.950 772.050 599.400 ;
        RECT 775.950 598.950 778.050 601.050 ;
        RECT 781.950 598.950 784.050 601.050 ;
        RECT 790.950 598.950 793.050 604.050 ;
        RECT 799.950 602.250 802.050 604.050 ;
        RECT 805.950 602.250 808.050 604.050 ;
        RECT 823.950 602.250 826.050 604.050 ;
        RECT 829.950 602.250 832.050 604.050 ;
        RECT 850.950 602.250 853.050 604.050 ;
        RECT 871.950 602.250 874.050 604.050 ;
        RECT 877.950 602.250 880.050 604.050 ;
        RECT 883.950 603.450 886.050 604.050 ;
        RECT 889.950 603.450 892.050 604.050 ;
        RECT 883.950 602.400 892.050 603.450 ;
        RECT 883.950 601.950 886.050 602.400 ;
        RECT 889.950 601.950 892.050 602.400 ;
        RECT 895.950 602.250 898.050 604.050 ;
        RECT 901.950 602.250 904.050 604.050 ;
        RECT 799.950 598.950 802.050 601.050 ;
        RECT 805.950 598.950 811.050 601.050 ;
        RECT 823.950 598.950 826.050 601.050 ;
        RECT 829.950 600.450 832.050 601.050 ;
        RECT 834.000 600.450 838.050 601.050 ;
        RECT 829.950 599.400 838.050 600.450 ;
        RECT 829.950 598.950 832.050 599.400 ;
        RECT 834.000 598.950 838.050 599.400 ;
        RECT 850.950 600.450 853.050 601.050 ;
        RECT 865.800 600.450 867.900 601.050 ;
        RECT 850.950 599.400 867.900 600.450 ;
        RECT 850.950 598.950 853.050 599.400 ;
        RECT 865.800 598.950 867.900 599.400 ;
        RECT 869.100 598.950 874.050 601.050 ;
        RECT 877.950 598.950 880.050 601.050 ;
        RECT 895.950 598.950 898.050 601.050 ;
        RECT 901.950 598.950 904.050 601.050 ;
        RECT 646.950 593.400 669.450 594.450 ;
        RECT 697.950 594.450 700.050 595.050 ;
        RECT 706.950 594.450 709.050 595.050 ;
        RECT 697.950 593.400 709.050 594.450 ;
        RECT 553.950 592.950 556.050 593.400 ;
        RECT 586.950 592.950 589.050 593.400 ;
        RECT 607.950 592.950 610.050 593.400 ;
        RECT 646.950 592.950 649.050 593.400 ;
        RECT 697.950 592.950 700.050 593.400 ;
        RECT 706.950 592.950 709.050 593.400 ;
        RECT 754.950 594.450 757.050 595.050 ;
        RECT 769.950 594.450 772.050 595.050 ;
        RECT 778.950 594.450 781.050 595.050 ;
        RECT 754.950 593.400 762.450 594.450 ;
        RECT 754.950 592.950 757.050 593.400 ;
        RECT 208.950 591.450 211.050 592.050 ;
        RECT 220.950 591.450 223.050 592.050 ;
        RECT 208.950 590.400 223.050 591.450 ;
        RECT 208.950 589.950 211.050 590.400 ;
        RECT 220.950 589.950 223.050 590.400 ;
        RECT 232.950 591.450 235.050 592.050 ;
        RECT 283.950 591.450 286.050 592.050 ;
        RECT 232.950 590.400 286.050 591.450 ;
        RECT 232.950 589.950 235.050 590.400 ;
        RECT 283.950 589.950 286.050 590.400 ;
        RECT 325.950 591.450 328.050 592.050 ;
        RECT 340.950 591.450 343.050 592.050 ;
        RECT 364.950 591.450 367.050 592.050 ;
        RECT 325.950 590.400 367.050 591.450 ;
        RECT 325.950 589.950 328.050 590.400 ;
        RECT 340.950 589.950 343.050 590.400 ;
        RECT 364.950 589.950 367.050 590.400 ;
        RECT 376.950 591.450 379.050 592.050 ;
        RECT 418.950 591.450 421.050 592.050 ;
        RECT 376.950 590.400 421.050 591.450 ;
        RECT 376.950 589.950 379.050 590.400 ;
        RECT 418.950 589.950 421.050 590.400 ;
        RECT 559.950 591.450 562.050 592.050 ;
        RECT 568.950 591.450 571.050 592.050 ;
        RECT 580.950 591.450 583.050 592.050 ;
        RECT 559.950 590.400 583.050 591.450 ;
        RECT 559.950 589.950 562.050 590.400 ;
        RECT 568.950 589.950 571.050 590.400 ;
        RECT 580.950 589.950 583.050 590.400 ;
        RECT 589.950 591.450 592.050 592.050 ;
        RECT 634.950 591.450 637.050 592.050 ;
        RECT 589.950 590.400 637.050 591.450 ;
        RECT 589.950 589.950 592.050 590.400 ;
        RECT 634.950 589.950 637.050 590.400 ;
        RECT 643.950 591.450 646.050 592.050 ;
        RECT 649.950 591.450 652.050 592.050 ;
        RECT 643.950 590.400 652.050 591.450 ;
        RECT 643.950 589.950 646.050 590.400 ;
        RECT 649.950 589.950 652.050 590.400 ;
        RECT 661.950 591.450 664.050 592.050 ;
        RECT 742.950 591.450 745.050 592.050 ;
        RECT 661.950 590.400 745.050 591.450 ;
        RECT 761.400 591.450 762.450 593.400 ;
        RECT 769.950 593.400 781.050 594.450 ;
        RECT 782.400 594.450 783.450 598.950 ;
        RECT 787.950 597.450 790.050 598.050 ;
        RECT 793.950 597.450 796.050 598.050 ;
        RECT 787.950 596.400 796.050 597.450 ;
        RECT 787.950 595.950 790.050 596.400 ;
        RECT 793.950 595.950 796.050 596.400 ;
        RECT 886.950 597.450 889.050 598.050 ;
        RECT 892.950 597.450 895.050 598.050 ;
        RECT 886.950 596.400 895.050 597.450 ;
        RECT 886.950 595.950 889.050 596.400 ;
        RECT 892.950 595.950 895.050 596.400 ;
        RECT 793.950 594.450 796.050 595.050 ;
        RECT 799.950 594.450 802.050 595.050 ;
        RECT 782.400 593.400 786.450 594.450 ;
        RECT 769.950 592.950 772.050 593.400 ;
        RECT 778.950 592.950 781.050 593.400 ;
        RECT 781.950 591.450 784.050 592.050 ;
        RECT 761.400 590.400 784.050 591.450 ;
        RECT 661.950 589.950 664.050 590.400 ;
        RECT 742.950 589.950 745.050 590.400 ;
        RECT 781.950 589.950 784.050 590.400 ;
        RECT 785.400 589.050 786.450 593.400 ;
        RECT 793.950 593.400 802.050 594.450 ;
        RECT 793.950 592.950 796.050 593.400 ;
        RECT 799.950 592.950 802.050 593.400 ;
        RECT 817.950 594.450 820.050 595.050 ;
        RECT 823.950 594.450 826.050 595.050 ;
        RECT 817.950 593.400 826.050 594.450 ;
        RECT 817.950 592.950 820.050 593.400 ;
        RECT 823.950 592.950 826.050 593.400 ;
        RECT 850.950 594.450 853.050 595.050 ;
        RECT 859.950 594.450 862.050 595.050 ;
        RECT 850.950 593.400 862.050 594.450 ;
        RECT 850.950 592.950 853.050 593.400 ;
        RECT 859.950 592.950 862.050 593.400 ;
        RECT 880.950 594.450 883.050 595.050 ;
        RECT 902.400 594.450 903.450 598.950 ;
        RECT 880.950 593.400 903.450 594.450 ;
        RECT 880.950 592.950 883.050 593.400 ;
        RECT 787.950 589.950 793.050 592.050 ;
        RECT 826.950 591.450 829.050 592.050 ;
        RECT 838.950 591.450 841.050 592.050 ;
        RECT 826.950 590.400 841.050 591.450 ;
        RECT 826.950 589.950 829.050 590.400 ;
        RECT 838.950 589.950 841.050 590.400 ;
        RECT 886.950 589.950 892.050 592.050 ;
        RECT 43.950 588.450 46.050 589.050 ;
        RECT 52.950 588.450 55.050 589.050 ;
        RECT 43.950 587.400 55.050 588.450 ;
        RECT 43.950 586.950 46.050 587.400 ;
        RECT 52.950 586.950 55.050 587.400 ;
        RECT 316.950 588.450 319.050 589.050 ;
        RECT 349.950 588.450 352.050 589.050 ;
        RECT 316.950 587.400 352.050 588.450 ;
        RECT 316.950 586.950 319.050 587.400 ;
        RECT 349.950 586.950 352.050 587.400 ;
        RECT 373.950 588.450 376.050 589.050 ;
        RECT 487.950 588.450 490.050 589.050 ;
        RECT 373.950 587.400 490.050 588.450 ;
        RECT 373.950 586.950 376.050 587.400 ;
        RECT 487.950 586.950 490.050 587.400 ;
        RECT 556.950 588.450 559.050 589.050 ;
        RECT 598.950 588.450 601.050 589.050 ;
        RECT 556.950 587.400 601.050 588.450 ;
        RECT 556.950 586.950 559.050 587.400 ;
        RECT 598.950 586.950 601.050 587.400 ;
        RECT 610.950 588.450 613.050 589.050 ;
        RECT 688.950 588.450 691.050 589.050 ;
        RECT 610.950 587.400 691.050 588.450 ;
        RECT 610.950 586.950 613.050 587.400 ;
        RECT 688.950 586.950 691.050 587.400 ;
        RECT 724.950 588.450 727.050 589.050 ;
        RECT 757.950 588.450 760.050 589.050 ;
        RECT 724.950 587.400 760.050 588.450 ;
        RECT 724.950 586.950 727.050 587.400 ;
        RECT 757.950 586.950 760.050 587.400 ;
        RECT 784.950 586.950 787.050 589.050 ;
        RECT 823.950 588.450 826.050 589.050 ;
        RECT 844.950 588.450 847.050 589.050 ;
        RECT 823.950 587.400 847.050 588.450 ;
        RECT 823.950 586.950 826.050 587.400 ;
        RECT 844.950 586.950 847.050 587.400 ;
        RECT 10.950 585.450 13.050 586.050 ;
        RECT 2.400 585.000 13.050 585.450 ;
        RECT 1.950 584.400 13.050 585.000 ;
        RECT 1.950 583.050 4.050 584.400 ;
        RECT 10.950 583.950 13.050 584.400 ;
        RECT 40.950 585.450 43.050 586.050 ;
        RECT 94.950 585.450 97.050 586.050 ;
        RECT 100.950 585.450 103.050 586.050 ;
        RECT 112.950 585.450 115.050 586.050 ;
        RECT 40.950 584.400 87.450 585.450 ;
        RECT 40.950 583.950 43.050 584.400 ;
        RECT 1.800 582.000 4.050 583.050 ;
        RECT 5.100 582.450 7.200 583.050 ;
        RECT 19.950 582.450 22.050 583.050 ;
        RECT 1.800 580.950 3.900 582.000 ;
        RECT 5.100 581.400 22.050 582.450 ;
        RECT 5.100 580.950 7.200 581.400 ;
        RECT 19.950 580.950 22.050 581.400 ;
        RECT 73.950 582.450 76.050 583.050 ;
        RECT 82.950 582.450 85.050 583.050 ;
        RECT 73.950 581.400 85.050 582.450 ;
        RECT 86.400 582.450 87.450 584.400 ;
        RECT 94.950 584.400 115.050 585.450 ;
        RECT 94.950 583.950 97.050 584.400 ;
        RECT 100.950 583.950 103.050 584.400 ;
        RECT 112.950 583.950 115.050 584.400 ;
        RECT 121.950 585.450 124.050 586.050 ;
        RECT 139.950 585.450 142.050 586.050 ;
        RECT 154.950 585.450 157.050 586.050 ;
        RECT 121.950 584.400 157.050 585.450 ;
        RECT 121.950 583.950 124.050 584.400 ;
        RECT 139.950 583.950 142.050 584.400 ;
        RECT 154.950 583.950 157.050 584.400 ;
        RECT 163.950 585.450 166.050 586.050 ;
        RECT 202.950 585.450 205.050 586.050 ;
        RECT 163.950 584.400 205.050 585.450 ;
        RECT 163.950 583.950 166.050 584.400 ;
        RECT 202.950 583.950 205.050 584.400 ;
        RECT 229.950 585.450 232.050 586.050 ;
        RECT 271.950 585.450 274.050 586.050 ;
        RECT 388.950 585.450 391.050 586.050 ;
        RECT 406.950 585.450 409.050 586.050 ;
        RECT 436.950 585.450 439.050 586.050 ;
        RECT 229.950 584.400 274.050 585.450 ;
        RECT 229.950 583.950 232.050 584.400 ;
        RECT 271.950 583.950 274.050 584.400 ;
        RECT 323.400 584.400 369.450 585.450 ;
        RECT 91.950 582.450 94.050 583.050 ;
        RECT 142.950 582.450 145.050 583.050 ;
        RECT 148.950 582.450 151.050 583.050 ;
        RECT 175.950 582.450 178.050 583.050 ;
        RECT 220.950 582.450 223.050 583.050 ;
        RECT 86.400 581.400 94.050 582.450 ;
        RECT 73.950 580.950 76.050 581.400 ;
        RECT 82.950 580.950 85.050 581.400 ;
        RECT 91.950 580.950 94.050 581.400 ;
        RECT 95.400 581.400 223.050 582.450 ;
        RECT 13.950 579.450 16.050 580.050 ;
        RECT 58.950 579.450 61.050 580.050 ;
        RECT 13.950 578.400 61.050 579.450 ;
        RECT 13.950 577.950 16.050 578.400 ;
        RECT 58.950 577.950 61.050 578.400 ;
        RECT 64.950 579.450 67.050 580.050 ;
        RECT 88.950 579.450 91.050 580.050 ;
        RECT 95.400 579.450 96.450 581.400 ;
        RECT 142.950 580.950 145.050 581.400 ;
        RECT 148.950 580.950 151.050 581.400 ;
        RECT 175.950 580.950 178.050 581.400 ;
        RECT 220.950 580.950 223.050 581.400 ;
        RECT 247.950 582.450 250.050 583.050 ;
        RECT 256.950 582.450 259.050 583.050 ;
        RECT 323.400 582.450 324.450 584.400 ;
        RECT 247.950 581.400 324.450 582.450 ;
        RECT 325.950 582.450 328.050 583.200 ;
        RECT 368.400 583.050 369.450 584.400 ;
        RECT 388.950 584.400 439.050 585.450 ;
        RECT 388.950 583.950 391.050 584.400 ;
        RECT 406.950 583.950 409.050 584.400 ;
        RECT 436.950 583.950 439.050 584.400 ;
        RECT 481.950 585.450 484.050 586.050 ;
        RECT 538.950 585.450 541.050 586.050 ;
        RECT 481.950 584.400 541.050 585.450 ;
        RECT 481.950 583.950 484.050 584.400 ;
        RECT 538.950 583.950 541.050 584.400 ;
        RECT 544.950 585.450 547.050 586.050 ;
        RECT 601.950 585.450 604.050 586.050 ;
        RECT 718.950 585.450 721.050 586.050 ;
        RECT 544.950 584.400 600.450 585.450 ;
        RECT 544.950 583.950 547.050 584.400 ;
        RECT 346.950 582.450 349.050 583.050 ;
        RECT 355.950 582.450 358.050 583.050 ;
        RECT 325.950 581.400 358.050 582.450 ;
        RECT 247.950 580.950 250.050 581.400 ;
        RECT 256.950 580.950 259.050 581.400 ;
        RECT 325.950 581.100 328.050 581.400 ;
        RECT 346.950 580.950 349.050 581.400 ;
        RECT 355.950 580.950 358.050 581.400 ;
        RECT 367.950 582.450 370.050 583.050 ;
        RECT 412.950 582.450 415.050 583.050 ;
        RECT 367.950 581.400 415.050 582.450 ;
        RECT 367.950 580.950 370.050 581.400 ;
        RECT 412.950 580.950 415.050 581.400 ;
        RECT 496.950 582.450 499.050 583.050 ;
        RECT 514.950 582.450 517.050 583.050 ;
        RECT 496.950 581.400 517.050 582.450 ;
        RECT 496.950 580.950 499.050 581.400 ;
        RECT 514.950 580.950 517.050 581.400 ;
        RECT 529.950 582.450 532.050 583.050 ;
        RECT 556.950 582.450 559.050 583.050 ;
        RECT 529.950 581.400 559.050 582.450 ;
        RECT 599.400 582.450 600.450 584.400 ;
        RECT 601.950 584.400 721.050 585.450 ;
        RECT 601.950 583.950 604.050 584.400 ;
        RECT 718.950 583.950 721.050 584.400 ;
        RECT 820.950 585.450 823.050 586.050 ;
        RECT 898.950 585.450 901.050 586.050 ;
        RECT 820.950 584.400 901.050 585.450 ;
        RECT 820.950 583.950 823.050 584.400 ;
        RECT 898.950 583.950 901.050 584.400 ;
        RECT 719.400 583.050 720.450 583.950 ;
        RECT 607.950 582.450 610.050 583.050 ;
        RECT 599.400 581.400 610.050 582.450 ;
        RECT 529.950 580.950 532.050 581.400 ;
        RECT 556.950 580.950 559.050 581.400 ;
        RECT 607.950 580.950 610.050 581.400 ;
        RECT 622.950 580.950 628.050 583.050 ;
        RECT 637.950 582.450 640.050 583.050 ;
        RECT 667.950 582.450 670.050 583.050 ;
        RECT 637.950 581.400 670.050 582.450 ;
        RECT 637.950 580.950 640.050 581.400 ;
        RECT 667.950 580.950 670.050 581.400 ;
        RECT 691.950 582.450 694.050 583.050 ;
        RECT 691.950 581.400 717.450 582.450 ;
        RECT 719.400 581.400 723.900 583.050 ;
        RECT 691.950 580.950 694.050 581.400 ;
        RECT 716.400 580.050 717.450 581.400 ;
        RECT 720.000 580.950 723.900 581.400 ;
        RECT 725.100 582.450 727.200 583.050 ;
        RECT 787.950 582.450 790.050 583.050 ;
        RECT 725.100 581.400 790.050 582.450 ;
        RECT 725.100 580.950 727.200 581.400 ;
        RECT 787.950 580.950 790.050 581.400 ;
        RECT 817.950 582.450 820.050 583.050 ;
        RECT 856.950 582.450 859.050 583.050 ;
        RECT 817.950 581.400 859.050 582.450 ;
        RECT 817.950 580.950 820.050 581.400 ;
        RECT 856.950 580.950 859.050 581.400 ;
        RECT 64.950 578.400 96.450 579.450 ;
        RECT 157.950 579.450 160.050 580.050 ;
        RECT 172.950 579.450 175.050 580.050 ;
        RECT 223.950 579.450 226.050 580.050 ;
        RECT 157.950 578.400 226.050 579.450 ;
        RECT 64.950 577.950 67.050 578.400 ;
        RECT 88.950 577.950 91.050 578.400 ;
        RECT 157.950 577.950 160.050 578.400 ;
        RECT 172.950 577.950 175.050 578.400 ;
        RECT 223.950 577.950 226.050 578.400 ;
        RECT 280.950 579.450 283.050 580.050 ;
        RECT 304.800 579.450 306.900 580.050 ;
        RECT 280.950 578.400 306.900 579.450 ;
        RECT 280.950 577.950 283.050 578.400 ;
        RECT 304.800 577.950 306.900 578.400 ;
        RECT 308.100 579.450 310.200 580.050 ;
        RECT 316.950 579.450 319.050 580.050 ;
        RECT 325.950 579.450 328.050 579.900 ;
        RECT 308.100 578.400 328.050 579.450 ;
        RECT 308.100 577.950 310.200 578.400 ;
        RECT 316.950 577.950 319.050 578.400 ;
        RECT 325.950 577.800 328.050 578.400 ;
        RECT 349.950 579.450 352.050 580.050 ;
        RECT 370.950 579.450 373.050 580.050 ;
        RECT 349.950 578.400 373.050 579.450 ;
        RECT 349.950 577.950 352.050 578.400 ;
        RECT 370.950 577.950 373.050 578.400 ;
        RECT 379.950 579.450 382.050 580.050 ;
        RECT 394.950 579.450 397.050 580.050 ;
        RECT 379.950 578.400 397.050 579.450 ;
        RECT 379.950 577.950 382.050 578.400 ;
        RECT 394.950 577.950 397.050 578.400 ;
        RECT 427.950 579.450 430.050 580.050 ;
        RECT 460.950 579.450 463.050 580.050 ;
        RECT 427.950 578.400 463.050 579.450 ;
        RECT 427.950 577.950 430.050 578.400 ;
        RECT 460.950 577.950 463.050 578.400 ;
        RECT 484.950 579.450 487.050 580.050 ;
        RECT 505.950 579.450 508.050 580.050 ;
        RECT 484.950 578.400 508.050 579.450 ;
        RECT 484.950 577.950 487.050 578.400 ;
        RECT 505.950 577.950 508.050 578.400 ;
        RECT 553.950 579.450 556.050 580.050 ;
        RECT 562.950 579.450 565.050 580.050 ;
        RECT 553.950 578.400 565.050 579.450 ;
        RECT 553.950 577.950 556.050 578.400 ;
        RECT 562.950 577.950 565.050 578.400 ;
        RECT 574.950 579.450 577.050 580.050 ;
        RECT 580.950 579.450 583.050 580.050 ;
        RECT 574.950 578.400 583.050 579.450 ;
        RECT 574.950 577.950 577.050 578.400 ;
        RECT 580.950 577.950 583.050 578.400 ;
        RECT 619.950 579.450 622.050 580.050 ;
        RECT 631.950 579.450 634.050 580.050 ;
        RECT 640.950 579.450 643.050 580.050 ;
        RECT 619.950 578.400 643.050 579.450 ;
        RECT 619.950 577.950 622.050 578.400 ;
        RECT 631.950 577.950 634.050 578.400 ;
        RECT 640.950 577.950 643.050 578.400 ;
        RECT 652.950 579.450 655.050 580.050 ;
        RECT 712.800 579.450 714.900 580.050 ;
        RECT 652.950 578.400 714.900 579.450 ;
        RECT 652.950 577.950 655.050 578.400 ;
        RECT 712.800 577.950 714.900 578.400 ;
        RECT 716.100 579.450 718.200 580.050 ;
        RECT 736.950 579.450 739.050 580.050 ;
        RECT 716.100 578.400 739.050 579.450 ;
        RECT 716.100 577.950 718.200 578.400 ;
        RECT 736.950 577.950 739.050 578.400 ;
        RECT 772.950 579.450 775.050 580.050 ;
        RECT 778.800 579.450 780.900 580.050 ;
        RECT 772.950 578.400 780.900 579.450 ;
        RECT 772.950 577.950 775.050 578.400 ;
        RECT 778.800 577.950 780.900 578.400 ;
        RECT 782.100 579.450 784.200 580.050 ;
        RECT 892.950 579.450 895.050 580.050 ;
        RECT 782.100 578.400 825.450 579.450 ;
        RECT 782.100 577.950 784.200 578.400 ;
        RECT 1.950 574.950 7.050 577.050 ;
        RECT 16.950 571.950 19.050 574.050 ;
        RECT 34.950 571.950 37.050 574.050 ;
        RECT 40.950 571.950 43.050 574.050 ;
        RECT 46.950 573.450 49.050 574.050 ;
        RECT 61.950 573.450 64.050 574.050 ;
        RECT 46.950 572.400 64.050 573.450 ;
        RECT 46.950 571.950 49.050 572.400 ;
        RECT 61.950 571.950 64.050 572.400 ;
        RECT 67.950 573.450 70.050 574.050 ;
        RECT 82.950 573.450 85.050 574.050 ;
        RECT 67.950 572.400 85.050 573.450 ;
        RECT 67.950 571.950 70.050 572.400 ;
        RECT 82.950 571.950 85.050 572.400 ;
        RECT 97.950 571.950 103.050 574.050 ;
        RECT 106.950 573.450 109.050 574.050 ;
        RECT 118.800 573.450 120.900 574.050 ;
        RECT 106.950 572.400 120.900 573.450 ;
        RECT 106.950 571.950 109.050 572.400 ;
        RECT 118.800 571.950 120.900 572.400 ;
        RECT 122.100 571.950 127.050 574.050 ;
        RECT 130.950 571.950 133.050 574.050 ;
        RECT 145.950 571.950 151.050 574.050 ;
        RECT 172.950 571.950 175.050 574.050 ;
        RECT 184.950 571.950 187.050 574.050 ;
        RECT 199.950 573.450 204.000 574.050 ;
        RECT 205.950 573.450 208.050 574.050 ;
        RECT 199.950 572.400 208.050 573.450 ;
        RECT 199.950 571.950 204.000 572.400 ;
        RECT 205.950 571.950 208.050 572.400 ;
        RECT 211.950 571.950 214.050 574.050 ;
        RECT 223.950 573.450 228.000 574.050 ;
        RECT 229.950 573.450 232.050 574.050 ;
        RECT 223.950 572.400 232.050 573.450 ;
        RECT 223.950 571.950 228.000 572.400 ;
        RECT 229.950 571.950 232.050 572.400 ;
        RECT 235.950 571.950 238.050 574.050 ;
        RECT 253.950 571.950 256.050 577.050 ;
        RECT 622.950 574.950 628.050 577.050 ;
        RECT 721.950 574.950 730.050 577.050 ;
        RECT 751.950 574.950 754.050 577.050 ;
        RECT 757.950 574.950 760.050 577.050 ;
        RECT 802.950 576.450 805.050 577.050 ;
        RECT 802.950 575.400 820.050 576.450 ;
        RECT 802.950 574.950 805.050 575.400 ;
        RECT 262.950 573.450 265.050 574.050 ;
        RECT 274.950 573.450 277.050 574.050 ;
        RECT 262.950 572.400 277.050 573.450 ;
        RECT 262.950 571.950 265.050 572.400 ;
        RECT 274.950 571.950 277.050 572.400 ;
        RECT 280.950 571.950 283.050 574.050 ;
        RECT 295.950 571.950 301.050 574.050 ;
        RECT 304.950 571.950 307.050 574.050 ;
        RECT 325.950 571.950 328.050 574.050 ;
        RECT 334.950 573.450 339.000 574.050 ;
        RECT 340.950 573.450 343.050 574.050 ;
        RECT 334.950 572.400 343.050 573.450 ;
        RECT 334.950 571.950 339.000 572.400 ;
        RECT 340.950 571.950 343.050 572.400 ;
        RECT 346.950 571.950 349.050 574.050 ;
        RECT 355.950 573.450 358.050 574.050 ;
        RECT 364.950 573.450 367.050 574.050 ;
        RECT 355.950 572.400 367.050 573.450 ;
        RECT 355.950 571.950 358.050 572.400 ;
        RECT 364.950 571.950 367.050 572.400 ;
        RECT 370.950 571.950 373.050 574.050 ;
        RECT 391.950 573.450 394.050 574.050 ;
        RECT 400.950 573.450 403.050 574.050 ;
        RECT 391.950 572.400 403.050 573.450 ;
        RECT 391.950 571.950 394.050 572.400 ;
        RECT 400.950 571.950 403.050 572.400 ;
        RECT 409.950 573.450 412.050 574.050 ;
        RECT 427.950 573.450 430.050 574.050 ;
        RECT 409.950 572.400 430.050 573.450 ;
        RECT 409.950 571.950 412.050 572.400 ;
        RECT 427.950 571.950 430.050 572.400 ;
        RECT 433.950 571.950 436.050 574.050 ;
        RECT 439.950 571.950 442.050 574.050 ;
        RECT 457.950 573.450 460.050 574.050 ;
        RECT 466.800 573.450 468.900 574.050 ;
        RECT 457.950 572.400 468.900 573.450 ;
        RECT 457.950 571.950 460.050 572.400 ;
        RECT 466.800 571.950 468.900 572.400 ;
        RECT 470.100 573.450 472.200 574.050 ;
        RECT 478.950 573.450 481.050 574.050 ;
        RECT 470.100 572.400 481.050 573.450 ;
        RECT 470.100 571.950 472.200 572.400 ;
        RECT 478.950 571.950 481.050 572.400 ;
        RECT 484.950 571.950 487.050 574.050 ;
        RECT 490.950 573.450 495.000 574.050 ;
        RECT 496.950 573.450 499.050 574.050 ;
        RECT 490.950 572.400 499.050 573.450 ;
        RECT 490.950 571.950 495.000 572.400 ;
        RECT 496.950 571.950 499.050 572.400 ;
        RECT 502.950 573.450 505.050 574.050 ;
        RECT 511.800 573.450 513.900 574.050 ;
        RECT 502.950 572.400 513.900 573.450 ;
        RECT 502.950 571.950 505.050 572.400 ;
        RECT 511.800 571.950 513.900 572.400 ;
        RECT 515.100 573.450 517.200 574.050 ;
        RECT 523.950 573.450 526.050 574.050 ;
        RECT 515.100 572.400 526.050 573.450 ;
        RECT 515.100 571.950 517.200 572.400 ;
        RECT 523.950 571.950 526.050 572.400 ;
        RECT 529.950 571.950 532.050 574.050 ;
        RECT 538.950 573.450 541.050 574.050 ;
        RECT 547.950 573.450 550.050 574.050 ;
        RECT 538.950 572.400 550.050 573.450 ;
        RECT 538.950 571.950 541.050 572.400 ;
        RECT 547.950 571.950 550.050 572.400 ;
        RECT 553.950 571.950 556.050 574.050 ;
        RECT 574.950 571.950 577.050 574.050 ;
        RECT 580.950 573.450 583.050 574.050 ;
        RECT 589.950 573.450 592.050 574.050 ;
        RECT 580.950 572.400 592.050 573.450 ;
        RECT 580.950 571.950 583.050 572.400 ;
        RECT 589.950 571.950 592.050 572.400 ;
        RECT 595.950 573.450 598.050 574.050 ;
        RECT 610.950 573.450 613.050 574.050 ;
        RECT 595.950 572.400 613.050 573.450 ;
        RECT 595.950 571.950 598.050 572.400 ;
        RECT 610.950 571.950 613.050 572.400 ;
        RECT 616.950 571.950 619.050 574.050 ;
        RECT 625.950 573.450 628.050 574.050 ;
        RECT 637.950 573.450 640.050 574.050 ;
        RECT 625.950 572.400 640.050 573.450 ;
        RECT 625.950 571.950 628.050 572.400 ;
        RECT 637.950 571.950 640.050 572.400 ;
        RECT 661.950 571.950 664.050 574.050 ;
        RECT 667.950 571.950 670.050 574.050 ;
        RECT 679.950 571.950 685.050 574.050 ;
        RECT 688.950 571.950 691.050 574.050 ;
        RECT 697.950 573.450 700.050 574.050 ;
        RECT 706.950 573.450 709.050 574.050 ;
        RECT 697.950 572.400 709.050 573.450 ;
        RECT 697.950 571.950 700.050 572.400 ;
        RECT 706.950 571.950 709.050 572.400 ;
        RECT 712.950 571.950 715.050 574.050 ;
        RECT 730.950 571.950 733.050 574.050 ;
        RECT 736.950 571.950 742.050 574.050 ;
        RECT 751.950 571.950 754.050 573.750 ;
        RECT 757.950 571.950 760.050 573.750 ;
        RECT 772.950 571.950 775.050 574.050 ;
        RECT 778.950 573.450 781.050 574.050 ;
        RECT 793.950 573.450 796.050 574.050 ;
        RECT 778.950 572.400 796.050 573.450 ;
        RECT 778.950 571.950 781.050 572.400 ;
        RECT 793.950 571.950 796.050 572.400 ;
        RECT 799.950 571.950 802.050 574.050 ;
        RECT 817.950 571.950 820.050 575.400 ;
        RECT 824.400 574.050 825.450 578.400 ;
        RECT 863.400 578.400 895.050 579.450 ;
        RECT 863.400 574.050 864.450 578.400 ;
        RECT 892.950 577.950 895.050 578.400 ;
        RECT 823.950 571.950 826.050 574.050 ;
        RECT 844.950 571.950 847.050 574.050 ;
        RECT 862.950 571.950 865.050 574.050 ;
        RECT 868.950 571.950 871.050 574.050 ;
        RECT 880.950 571.950 883.050 574.050 ;
        RECT 886.950 573.450 889.050 574.050 ;
        RECT 898.950 573.450 901.050 574.050 ;
        RECT 886.950 572.400 901.050 573.450 ;
        RECT 886.950 571.950 889.050 572.400 ;
        RECT 898.950 571.950 901.050 572.400 ;
        RECT 613.950 570.750 615.750 571.050 ;
        RECT 16.950 568.950 19.050 570.750 ;
        RECT 34.950 568.950 37.050 570.750 ;
        RECT 40.950 568.950 43.050 570.750 ;
        RECT 61.950 568.950 64.050 570.750 ;
        RECT 82.950 568.950 85.050 570.750 ;
        RECT 100.950 568.950 103.050 570.750 ;
        RECT 106.950 568.950 109.050 570.750 ;
        RECT 124.950 568.950 127.050 570.750 ;
        RECT 130.950 568.950 133.050 570.750 ;
        RECT 148.950 568.950 151.050 570.750 ;
        RECT 172.950 568.950 175.050 570.750 ;
        RECT 184.950 568.950 187.050 570.750 ;
        RECT 205.950 568.950 208.050 570.750 ;
        RECT 211.950 568.950 214.050 570.750 ;
        RECT 229.950 568.950 232.050 570.750 ;
        RECT 235.950 568.950 238.050 570.750 ;
        RECT 253.950 568.950 256.050 570.750 ;
        RECT 274.950 568.950 277.050 570.750 ;
        RECT 280.950 568.950 283.050 570.750 ;
        RECT 298.950 568.950 301.050 570.750 ;
        RECT 304.950 568.950 307.050 570.750 ;
        RECT 325.950 568.950 328.050 570.750 ;
        RECT 340.950 568.950 343.050 570.750 ;
        RECT 346.950 568.950 349.050 570.750 ;
        RECT 364.950 568.950 367.050 570.750 ;
        RECT 370.950 568.950 373.050 570.750 ;
        RECT 391.950 568.950 394.050 570.750 ;
        RECT 409.950 568.950 412.050 570.750 ;
        RECT 433.950 568.950 436.050 570.750 ;
        RECT 439.950 568.950 442.050 570.750 ;
        RECT 457.950 568.950 460.050 570.750 ;
        RECT 478.950 568.950 481.050 570.750 ;
        RECT 484.950 568.950 487.050 570.750 ;
        RECT 496.950 568.950 499.050 570.750 ;
        RECT 502.950 568.950 505.050 570.750 ;
        RECT 523.950 568.950 526.050 570.750 ;
        RECT 529.950 568.950 532.050 570.750 ;
        RECT 547.950 568.950 550.050 570.750 ;
        RECT 553.950 568.950 556.050 570.750 ;
        RECT 574.950 568.950 577.050 570.750 ;
        RECT 589.950 568.950 592.050 570.750 ;
        RECT 595.950 568.950 598.050 570.750 ;
        RECT 613.950 569.250 616.050 570.750 ;
        RECT 616.950 569.250 619.050 570.750 ;
        RECT 622.950 569.250 625.050 571.050 ;
        RECT 617.250 568.950 619.050 569.250 ;
        RECT 637.950 568.950 640.050 570.750 ;
        RECT 661.950 568.950 664.050 570.750 ;
        RECT 667.950 568.950 670.050 570.750 ;
        RECT 682.950 568.950 685.050 570.750 ;
        RECT 688.950 568.950 691.050 570.750 ;
        RECT 706.950 568.950 709.050 570.750 ;
        RECT 712.950 568.950 715.050 570.750 ;
        RECT 730.950 568.950 733.050 570.750 ;
        RECT 736.950 568.950 739.050 570.750 ;
        RECT 754.950 569.250 757.050 571.050 ;
        RECT 772.950 568.950 775.050 570.750 ;
        RECT 793.950 568.950 796.050 570.750 ;
        RECT 799.950 568.950 802.050 570.750 ;
        RECT 817.950 568.950 820.050 570.750 ;
        RECT 823.950 568.950 826.050 570.750 ;
        RECT 844.950 568.950 847.050 570.750 ;
        RECT 862.950 568.950 865.050 570.750 ;
        RECT 868.950 568.950 871.050 570.750 ;
        RECT 880.950 568.950 883.050 570.750 ;
        RECT 898.950 568.950 901.050 570.750 ;
        RECT 904.950 569.250 907.050 571.050 ;
        RECT 13.950 566.250 16.050 568.050 ;
        RECT 19.950 566.250 22.050 568.050 ;
        RECT 31.950 566.250 34.050 568.050 ;
        RECT 37.950 566.250 40.050 568.050 ;
        RECT 58.950 566.250 61.050 568.050 ;
        RECT 64.950 566.250 67.050 568.050 ;
        RECT 79.950 566.250 82.050 568.050 ;
        RECT 85.950 566.250 88.050 568.050 ;
        RECT 103.950 566.250 106.050 568.050 ;
        RECT 109.950 566.250 112.050 568.050 ;
        RECT 127.950 566.250 130.050 568.050 ;
        RECT 133.950 566.250 136.050 568.050 ;
        RECT 145.950 566.250 148.050 568.050 ;
        RECT 151.950 566.250 154.050 568.050 ;
        RECT 169.950 566.250 172.050 568.050 ;
        RECT 187.950 566.250 190.050 568.050 ;
        RECT 208.950 566.250 211.050 568.050 ;
        RECT 214.950 566.250 217.050 568.050 ;
        RECT 232.950 566.250 235.050 568.050 ;
        RECT 238.950 566.250 241.050 568.050 ;
        RECT 250.950 566.250 253.050 568.050 ;
        RECT 256.950 566.250 259.050 568.050 ;
        RECT 277.950 566.250 280.050 568.050 ;
        RECT 283.950 566.250 286.050 568.050 ;
        RECT 301.950 566.250 304.050 568.050 ;
        RECT 307.950 566.250 310.050 568.050 ;
        RECT 322.950 566.250 325.050 568.050 ;
        RECT 343.950 566.250 346.050 568.050 ;
        RECT 349.950 566.250 352.050 568.050 ;
        RECT 367.950 566.250 370.050 568.050 ;
        RECT 373.950 566.250 376.050 568.050 ;
        RECT 388.950 566.250 391.050 568.050 ;
        RECT 394.950 566.250 397.050 568.050 ;
        RECT 406.950 566.250 409.050 568.050 ;
        RECT 412.950 566.250 415.050 568.050 ;
        RECT 430.950 566.250 433.050 568.050 ;
        RECT 436.950 566.250 439.050 568.050 ;
        RECT 454.950 566.250 457.050 568.050 ;
        RECT 460.950 566.250 463.050 568.050 ;
        RECT 475.950 566.250 478.050 568.050 ;
        RECT 481.950 566.250 484.050 568.050 ;
        RECT 499.950 566.250 502.050 568.050 ;
        RECT 505.950 566.250 508.050 568.050 ;
        RECT 526.950 566.250 529.050 568.050 ;
        RECT 532.950 566.250 535.050 568.050 ;
        RECT 550.950 566.250 553.050 568.050 ;
        RECT 556.950 566.250 559.050 568.050 ;
        RECT 571.950 566.250 574.050 568.050 ;
        RECT 586.950 566.250 589.050 568.050 ;
        RECT 592.950 566.250 595.050 568.050 ;
        RECT 598.950 567.450 601.050 568.050 ;
        RECT 613.950 567.450 616.050 568.050 ;
        RECT 598.950 566.400 616.050 567.450 ;
        RECT 598.950 565.950 601.050 566.400 ;
        RECT 613.950 565.950 616.050 566.400 ;
        RECT 622.950 565.950 625.050 568.050 ;
        RECT 634.950 566.250 637.050 568.050 ;
        RECT 640.950 566.250 643.050 568.050 ;
        RECT 658.950 566.250 661.050 568.050 ;
        RECT 664.950 566.250 667.050 568.050 ;
        RECT 685.950 566.250 688.050 568.050 ;
        RECT 691.950 566.250 694.050 568.050 ;
        RECT 709.950 566.250 712.050 568.050 ;
        RECT 715.950 566.250 718.050 568.050 ;
        RECT 727.950 566.250 730.050 568.050 ;
        RECT 733.950 566.250 736.050 568.050 ;
        RECT 754.950 565.950 757.050 568.050 ;
        RECT 775.950 566.250 778.050 568.050 ;
        RECT 796.950 566.250 799.050 568.050 ;
        RECT 802.950 566.250 805.050 568.050 ;
        RECT 814.950 566.250 817.050 568.050 ;
        RECT 820.950 566.250 823.050 568.050 ;
        RECT 841.950 566.250 844.050 568.050 ;
        RECT 859.950 566.250 862.050 568.050 ;
        RECT 865.950 566.250 868.050 568.050 ;
        RECT 883.950 566.250 886.050 568.050 ;
        RECT 13.950 562.950 16.050 565.050 ;
        RECT 19.950 562.950 22.050 565.050 ;
        RECT 31.950 562.950 34.050 565.050 ;
        RECT 37.950 562.950 40.050 565.050 ;
        RECT 58.950 562.950 61.050 565.050 ;
        RECT 64.950 562.950 67.050 565.050 ;
        RECT 79.950 562.950 82.050 565.050 ;
        RECT 85.950 562.950 88.050 565.050 ;
        RECT 103.950 562.950 106.050 565.050 ;
        RECT 109.950 562.950 114.900 565.050 ;
        RECT 116.100 564.450 118.200 565.050 ;
        RECT 127.950 564.450 130.050 565.050 ;
        RECT 116.100 563.400 130.050 564.450 ;
        RECT 116.100 562.950 118.200 563.400 ;
        RECT 127.950 562.950 130.050 563.400 ;
        RECT 133.950 562.950 136.050 565.050 ;
        RECT 142.950 562.950 148.050 565.050 ;
        RECT 169.950 562.950 172.050 565.050 ;
        RECT 187.950 564.450 190.050 565.050 ;
        RECT 202.950 564.450 205.050 565.050 ;
        RECT 187.950 563.400 205.050 564.450 ;
        RECT 187.950 562.950 190.050 563.400 ;
        RECT 202.950 562.950 205.050 563.400 ;
        RECT 208.950 562.950 211.050 565.050 ;
        RECT 214.950 562.950 217.050 565.050 ;
        RECT 220.950 564.450 223.050 565.050 ;
        RECT 232.950 564.450 235.050 565.050 ;
        RECT 220.950 563.400 235.050 564.450 ;
        RECT 220.950 562.950 223.050 563.400 ;
        RECT 232.950 562.950 235.050 563.400 ;
        RECT 238.950 562.950 241.050 565.050 ;
        RECT 256.950 562.950 259.050 565.050 ;
        RECT 277.950 562.950 280.050 565.050 ;
        RECT 283.950 562.950 286.050 565.050 ;
        RECT 289.950 564.450 292.050 565.050 ;
        RECT 301.950 564.450 304.050 565.050 ;
        RECT 289.950 563.400 304.050 564.450 ;
        RECT 289.950 562.950 292.050 563.400 ;
        RECT 301.950 562.950 304.050 563.400 ;
        RECT 307.950 562.950 310.050 565.050 ;
        RECT 322.950 562.950 325.050 565.050 ;
        RECT 343.950 562.950 346.050 565.050 ;
        RECT 349.950 562.950 352.050 565.050 ;
        RECT 367.950 562.950 370.050 565.050 ;
        RECT 373.950 562.950 376.050 565.050 ;
        RECT 388.950 562.950 391.050 565.050 ;
        RECT 394.950 562.950 397.050 565.050 ;
        RECT 412.950 562.950 415.050 565.050 ;
        RECT 430.950 562.950 433.050 565.050 ;
        RECT 436.950 562.950 439.050 565.050 ;
        RECT 454.950 562.950 457.050 565.050 ;
        RECT 460.950 562.950 463.050 565.050 ;
        RECT 466.950 564.450 469.050 565.050 ;
        RECT 475.950 564.450 478.050 565.050 ;
        RECT 466.950 563.400 478.050 564.450 ;
        RECT 466.950 562.950 469.050 563.400 ;
        RECT 475.950 562.950 478.050 563.400 ;
        RECT 16.950 558.450 19.050 559.050 ;
        RECT 31.950 558.450 34.050 559.050 ;
        RECT 16.950 557.400 34.050 558.450 ;
        RECT 16.950 556.950 19.050 557.400 ;
        RECT 31.950 556.950 34.050 557.400 ;
        RECT 37.950 558.450 40.050 559.050 ;
        RECT 46.950 558.450 49.050 559.050 ;
        RECT 37.950 557.400 49.050 558.450 ;
        RECT 37.950 556.950 40.050 557.400 ;
        RECT 46.950 556.950 49.050 557.400 ;
        RECT 64.950 558.450 67.050 559.050 ;
        RECT 73.950 558.450 76.050 559.050 ;
        RECT 104.400 558.450 105.450 562.950 ;
        RECT 112.950 558.450 115.050 559.050 ;
        RECT 133.950 558.450 136.050 559.050 ;
        RECT 64.950 557.400 111.450 558.450 ;
        RECT 64.950 556.950 67.050 557.400 ;
        RECT 73.950 556.950 76.050 557.400 ;
        RECT 52.950 555.450 55.050 556.050 ;
        RECT 79.950 555.450 82.050 556.050 ;
        RECT 106.950 555.450 109.050 556.050 ;
        RECT 52.950 554.400 109.050 555.450 ;
        RECT 110.400 555.450 111.450 557.400 ;
        RECT 112.950 557.400 136.050 558.450 ;
        RECT 112.950 556.950 115.050 557.400 ;
        RECT 133.950 556.950 136.050 557.400 ;
        RECT 169.950 558.450 172.050 559.050 ;
        RECT 193.950 558.450 196.050 559.050 ;
        RECT 169.950 557.400 196.050 558.450 ;
        RECT 169.950 556.950 172.050 557.400 ;
        RECT 193.950 556.950 196.050 557.400 ;
        RECT 277.950 558.450 280.050 559.050 ;
        RECT 307.950 558.450 310.050 559.050 ;
        RECT 323.400 558.450 324.450 562.950 ;
        RECT 481.950 561.450 484.050 565.050 ;
        RECT 499.950 562.950 502.050 565.050 ;
        RECT 505.950 564.450 508.050 565.050 ;
        RECT 517.950 564.450 520.050 565.050 ;
        RECT 505.950 563.400 520.050 564.450 ;
        RECT 505.950 562.950 508.050 563.400 ;
        RECT 517.950 562.950 520.050 563.400 ;
        RECT 526.950 562.950 529.050 565.050 ;
        RECT 532.950 562.950 535.050 565.050 ;
        RECT 550.950 562.950 553.050 565.050 ;
        RECT 556.950 564.450 559.050 565.050 ;
        RECT 565.950 564.450 568.050 565.050 ;
        RECT 556.950 563.400 568.050 564.450 ;
        RECT 556.950 562.950 559.050 563.400 ;
        RECT 565.950 562.950 568.050 563.400 ;
        RECT 571.950 564.450 574.050 565.050 ;
        RECT 576.000 564.450 580.050 565.050 ;
        RECT 571.950 563.400 580.050 564.450 ;
        RECT 571.950 562.950 574.050 563.400 ;
        RECT 576.000 562.950 580.050 563.400 ;
        RECT 586.950 562.950 589.050 565.050 ;
        RECT 592.950 562.950 595.050 565.050 ;
        RECT 634.950 562.950 637.050 565.050 ;
        RECT 640.950 562.950 643.050 565.050 ;
        RECT 658.950 562.950 661.050 565.050 ;
        RECT 664.950 562.950 667.050 565.050 ;
        RECT 685.950 562.950 688.050 565.050 ;
        RECT 691.950 562.950 694.050 565.050 ;
        RECT 709.950 562.950 712.050 565.050 ;
        RECT 715.950 562.950 718.050 565.050 ;
        RECT 727.950 562.950 730.050 565.050 ;
        RECT 733.950 562.950 736.050 565.050 ;
        RECT 496.950 561.450 499.050 562.050 ;
        RECT 481.950 560.400 499.050 561.450 ;
        RECT 496.950 559.950 499.050 560.400 ;
        RECT 577.950 559.950 583.050 562.050 ;
        RECT 755.400 561.450 756.450 565.950 ;
        RECT 760.950 564.450 763.050 565.050 ;
        RECT 766.950 564.450 769.050 565.050 ;
        RECT 775.950 564.450 778.050 565.050 ;
        RECT 760.950 563.400 778.050 564.450 ;
        RECT 760.950 562.950 763.050 563.400 ;
        RECT 766.950 562.950 769.050 563.400 ;
        RECT 775.950 562.950 778.050 563.400 ;
        RECT 796.950 562.950 799.050 565.050 ;
        RECT 802.950 562.950 805.050 565.050 ;
        RECT 814.950 562.950 817.050 565.050 ;
        RECT 820.950 562.950 823.050 565.050 ;
        RECT 841.950 562.950 844.050 565.050 ;
        RECT 859.950 562.950 862.050 565.050 ;
        RECT 865.950 562.950 868.050 565.050 ;
        RECT 883.950 562.950 886.050 565.050 ;
        RECT 763.950 561.450 766.050 562.050 ;
        RECT 755.400 560.400 766.050 561.450 ;
        RECT 763.950 559.950 766.050 560.400 ;
        RECT 340.950 558.450 343.050 559.050 ;
        RECT 277.950 557.400 343.050 558.450 ;
        RECT 277.950 556.950 280.050 557.400 ;
        RECT 307.950 556.950 310.050 557.400 ;
        RECT 340.950 556.950 343.050 557.400 ;
        RECT 355.950 558.450 358.050 559.050 ;
        RECT 373.950 558.450 376.050 559.050 ;
        RECT 379.950 558.450 382.050 559.050 ;
        RECT 355.950 557.400 382.050 558.450 ;
        RECT 355.950 556.950 358.050 557.400 ;
        RECT 373.950 556.950 376.050 557.400 ;
        RECT 379.950 556.950 382.050 557.400 ;
        RECT 412.950 558.450 415.050 559.050 ;
        RECT 427.950 558.450 430.050 559.050 ;
        RECT 436.950 558.450 439.050 559.050 ;
        RECT 412.950 557.400 439.050 558.450 ;
        RECT 412.950 556.950 415.050 557.400 ;
        RECT 427.950 556.950 430.050 557.400 ;
        RECT 436.950 556.950 439.050 557.400 ;
        RECT 463.950 558.450 466.050 559.050 ;
        RECT 520.950 558.450 523.050 559.050 ;
        RECT 463.950 557.400 523.050 558.450 ;
        RECT 463.950 556.950 466.050 557.400 ;
        RECT 520.950 556.950 523.050 557.400 ;
        RECT 526.950 558.450 529.050 559.050 ;
        RECT 562.950 558.450 565.050 559.050 ;
        RECT 586.950 558.450 589.050 559.050 ;
        RECT 598.950 558.450 601.050 559.050 ;
        RECT 526.950 557.400 601.050 558.450 ;
        RECT 526.950 556.950 529.050 557.400 ;
        RECT 562.950 556.950 565.050 557.400 ;
        RECT 586.950 556.950 589.050 557.400 ;
        RECT 598.950 556.950 601.050 557.400 ;
        RECT 634.950 558.450 637.050 559.050 ;
        RECT 646.950 558.450 649.050 559.050 ;
        RECT 634.950 557.400 649.050 558.450 ;
        RECT 634.950 556.950 637.050 557.400 ;
        RECT 646.950 556.950 649.050 557.400 ;
        RECT 709.950 558.450 712.050 559.050 ;
        RECT 721.950 558.450 724.050 559.050 ;
        RECT 727.950 558.450 730.050 559.050 ;
        RECT 709.950 557.400 730.050 558.450 ;
        RECT 842.400 558.450 843.450 562.950 ;
        RECT 859.950 558.450 862.050 559.050 ;
        RECT 842.400 557.400 862.050 558.450 ;
        RECT 709.950 556.950 712.050 557.400 ;
        RECT 721.950 556.950 724.050 557.400 ;
        RECT 727.950 556.950 730.050 557.400 ;
        RECT 859.950 556.950 862.050 557.400 ;
        RECT 865.950 558.450 868.050 559.050 ;
        RECT 884.400 558.450 885.450 562.950 ;
        RECT 865.950 557.400 885.450 558.450 ;
        RECT 865.950 556.950 868.050 557.400 ;
        RECT 115.800 555.450 117.900 556.050 ;
        RECT 110.400 554.400 117.900 555.450 ;
        RECT 52.950 553.950 55.050 554.400 ;
        RECT 79.950 553.950 82.050 554.400 ;
        RECT 106.950 553.950 109.050 554.400 ;
        RECT 115.800 553.950 117.900 554.400 ;
        RECT 119.100 555.450 121.200 556.050 ;
        RECT 130.950 555.450 133.050 556.050 ;
        RECT 160.950 555.450 163.050 556.050 ;
        RECT 119.100 554.400 163.050 555.450 ;
        RECT 119.100 553.950 121.200 554.400 ;
        RECT 130.950 553.950 133.050 554.400 ;
        RECT 160.950 553.950 163.050 554.400 ;
        RECT 199.950 555.450 202.050 556.050 ;
        RECT 214.950 555.450 217.050 556.050 ;
        RECT 199.950 554.400 217.050 555.450 ;
        RECT 199.950 553.950 202.050 554.400 ;
        RECT 214.950 553.950 217.050 554.400 ;
        RECT 238.950 555.450 241.050 556.050 ;
        RECT 328.950 555.450 331.050 556.050 ;
        RECT 238.950 554.400 331.050 555.450 ;
        RECT 238.950 553.950 241.050 554.400 ;
        RECT 328.950 553.950 331.050 554.400 ;
        RECT 400.950 555.450 403.050 556.050 ;
        RECT 544.950 555.450 547.050 556.050 ;
        RECT 400.950 554.400 547.050 555.450 ;
        RECT 400.950 553.950 403.050 554.400 ;
        RECT 544.950 553.950 547.050 554.400 ;
        RECT 568.950 555.450 571.050 556.050 ;
        RECT 589.950 555.450 592.050 556.050 ;
        RECT 673.950 555.450 676.050 556.050 ;
        RECT 568.950 554.400 676.050 555.450 ;
        RECT 568.950 553.950 571.050 554.400 ;
        RECT 589.950 553.950 592.050 554.400 ;
        RECT 673.950 553.950 676.050 554.400 ;
        RECT 691.950 555.450 694.050 556.050 ;
        RECT 706.950 555.450 709.050 556.050 ;
        RECT 721.950 555.450 724.050 556.050 ;
        RECT 691.950 554.400 724.050 555.450 ;
        RECT 691.950 553.950 694.050 554.400 ;
        RECT 706.950 553.950 709.050 554.400 ;
        RECT 721.950 553.950 724.050 554.400 ;
        RECT 784.950 555.450 787.050 556.050 ;
        RECT 844.950 555.450 847.050 556.050 ;
        RECT 862.950 555.450 865.050 556.050 ;
        RECT 874.950 555.450 877.050 556.050 ;
        RECT 784.950 554.400 877.050 555.450 ;
        RECT 784.950 553.950 787.050 554.400 ;
        RECT 844.950 553.950 847.050 554.400 ;
        RECT 862.950 553.950 865.050 554.400 ;
        RECT 874.950 553.950 877.050 554.400 ;
        RECT 70.950 552.450 73.050 553.050 ;
        RECT 85.950 552.450 88.050 553.050 ;
        RECT 70.950 551.400 88.050 552.450 ;
        RECT 70.950 550.950 73.050 551.400 ;
        RECT 85.950 550.950 88.050 551.400 ;
        RECT 91.950 552.450 94.050 553.050 ;
        RECT 112.950 552.450 115.050 553.050 ;
        RECT 91.950 551.400 115.050 552.450 ;
        RECT 91.950 550.950 94.050 551.400 ;
        RECT 112.950 550.950 115.050 551.400 ;
        RECT 118.950 550.950 124.050 553.050 ;
        RECT 127.950 552.450 130.050 553.050 ;
        RECT 145.950 552.450 148.050 553.050 ;
        RECT 127.950 551.400 148.050 552.450 ;
        RECT 127.950 550.950 130.050 551.400 ;
        RECT 145.950 550.950 148.050 551.400 ;
        RECT 334.950 552.450 337.050 553.050 ;
        RECT 343.950 552.450 346.050 553.050 ;
        RECT 334.950 551.400 346.050 552.450 ;
        RECT 334.950 550.950 337.050 551.400 ;
        RECT 343.950 550.950 346.050 551.400 ;
        RECT 349.950 552.450 352.050 553.050 ;
        RECT 355.950 552.450 358.050 553.050 ;
        RECT 367.950 552.450 370.050 553.050 ;
        RECT 349.950 551.400 370.050 552.450 ;
        RECT 349.950 550.950 352.050 551.400 ;
        RECT 355.950 550.950 358.050 551.400 ;
        RECT 367.950 550.950 370.050 551.400 ;
        RECT 412.950 552.450 415.050 553.050 ;
        RECT 418.950 552.450 421.050 553.050 ;
        RECT 463.800 552.450 465.900 553.050 ;
        RECT 412.950 551.400 465.900 552.450 ;
        RECT 467.100 552.000 469.200 553.050 ;
        RECT 412.950 550.950 415.050 551.400 ;
        RECT 418.950 550.950 421.050 551.400 ;
        RECT 463.800 550.950 465.900 551.400 ;
        RECT 466.950 550.950 469.200 552.000 ;
        RECT 502.950 552.450 505.050 553.050 ;
        RECT 511.950 552.450 514.050 553.050 ;
        RECT 502.950 551.400 514.050 552.450 ;
        RECT 502.950 550.950 505.050 551.400 ;
        RECT 511.950 550.950 514.050 551.400 ;
        RECT 565.950 552.450 568.050 553.050 ;
        RECT 574.800 552.450 576.900 553.050 ;
        RECT 565.950 551.400 576.900 552.450 ;
        RECT 565.950 550.950 568.050 551.400 ;
        RECT 574.800 550.950 576.900 551.400 ;
        RECT 578.100 552.450 580.200 553.050 ;
        RECT 592.950 552.450 595.050 553.050 ;
        RECT 578.100 551.400 595.050 552.450 ;
        RECT 578.100 550.950 580.200 551.400 ;
        RECT 592.950 550.950 595.050 551.400 ;
        RECT 634.950 552.450 637.050 553.050 ;
        RECT 652.950 552.450 655.050 553.050 ;
        RECT 634.950 551.400 655.050 552.450 ;
        RECT 634.950 550.950 637.050 551.400 ;
        RECT 652.950 550.950 655.050 551.400 ;
        RECT 754.950 552.450 757.050 553.050 ;
        RECT 781.950 552.450 784.050 553.050 ;
        RECT 754.950 551.400 784.050 552.450 ;
        RECT 754.950 550.950 757.050 551.400 ;
        RECT 781.950 550.950 784.050 551.400 ;
        RECT 796.950 552.450 799.050 553.050 ;
        RECT 820.950 552.450 823.050 553.050 ;
        RECT 796.950 551.400 823.050 552.450 ;
        RECT 796.950 550.950 799.050 551.400 ;
        RECT 820.950 550.950 823.050 551.400 ;
        RECT 133.950 549.450 136.050 550.050 ;
        RECT 139.950 549.450 142.050 550.050 ;
        RECT 160.950 549.450 163.050 550.050 ;
        RECT 238.950 549.450 241.050 550.050 ;
        RECT 133.950 548.400 156.450 549.450 ;
        RECT 133.950 547.950 136.050 548.400 ;
        RECT 139.950 547.950 142.050 548.400 ;
        RECT 31.950 546.450 34.050 547.050 ;
        RECT 76.950 546.450 79.050 547.050 ;
        RECT 31.950 545.400 79.050 546.450 ;
        RECT 155.400 546.450 156.450 548.400 ;
        RECT 160.950 548.400 241.050 549.450 ;
        RECT 160.950 547.950 163.050 548.400 ;
        RECT 238.950 547.950 241.050 548.400 ;
        RECT 280.950 549.450 283.050 550.050 ;
        RECT 322.950 549.450 325.050 550.050 ;
        RECT 337.950 549.450 340.050 550.050 ;
        RECT 280.950 548.400 340.050 549.450 ;
        RECT 280.950 547.950 283.050 548.400 ;
        RECT 322.950 547.950 325.050 548.400 ;
        RECT 337.950 547.950 340.050 548.400 ;
        RECT 460.950 549.450 463.050 550.050 ;
        RECT 466.950 549.450 469.050 550.950 ;
        RECT 460.950 549.000 469.050 549.450 ;
        RECT 532.950 549.450 535.050 550.050 ;
        RECT 550.950 549.450 553.050 550.050 ;
        RECT 577.950 549.450 580.050 550.050 ;
        RECT 460.950 548.400 468.450 549.000 ;
        RECT 532.950 548.400 580.050 549.450 ;
        RECT 460.950 547.950 463.050 548.400 ;
        RECT 532.950 547.950 535.050 548.400 ;
        RECT 550.950 547.950 553.050 548.400 ;
        RECT 577.950 547.950 580.050 548.400 ;
        RECT 607.950 549.450 610.050 550.050 ;
        RECT 658.950 549.450 661.050 550.050 ;
        RECT 607.950 548.400 661.050 549.450 ;
        RECT 607.950 547.950 610.050 548.400 ;
        RECT 658.950 547.950 661.050 548.400 ;
        RECT 742.950 549.450 745.050 550.050 ;
        RECT 886.950 549.450 889.050 550.050 ;
        RECT 742.950 548.400 889.050 549.450 ;
        RECT 742.950 547.950 745.050 548.400 ;
        RECT 886.950 547.950 889.050 548.400 ;
        RECT 166.950 546.450 169.050 547.050 ;
        RECT 155.400 545.400 169.050 546.450 ;
        RECT 31.950 544.950 34.050 545.400 ;
        RECT 76.950 544.950 79.050 545.400 ;
        RECT 166.950 544.950 169.050 545.400 ;
        RECT 418.950 546.450 421.050 547.050 ;
        RECT 442.950 546.450 445.050 547.050 ;
        RECT 418.950 545.400 445.050 546.450 ;
        RECT 418.950 544.950 421.050 545.400 ;
        RECT 442.950 544.950 445.050 545.400 ;
        RECT 463.950 546.450 466.050 547.050 ;
        RECT 469.950 546.450 472.050 547.200 ;
        RECT 478.950 546.450 481.050 547.050 ;
        RECT 463.950 545.400 481.050 546.450 ;
        RECT 463.950 544.950 466.050 545.400 ;
        RECT 469.950 545.100 472.050 545.400 ;
        RECT 478.950 544.950 481.050 545.400 ;
        RECT 496.950 546.450 499.050 547.050 ;
        RECT 517.950 546.450 520.050 547.050 ;
        RECT 496.950 545.400 520.050 546.450 ;
        RECT 496.950 544.950 499.050 545.400 ;
        RECT 517.950 544.950 520.050 545.400 ;
        RECT 772.950 546.450 775.050 547.050 ;
        RECT 784.950 546.450 787.050 547.050 ;
        RECT 772.950 545.400 787.050 546.450 ;
        RECT 772.950 544.950 775.050 545.400 ;
        RECT 784.950 544.950 787.050 545.400 ;
        RECT 808.950 546.450 811.050 547.050 ;
        RECT 814.950 546.450 817.050 547.050 ;
        RECT 808.950 545.400 817.050 546.450 ;
        RECT 808.950 544.950 811.050 545.400 ;
        RECT 814.950 544.950 817.050 545.400 ;
        RECT 355.950 543.450 358.050 544.050 ;
        RECT 412.950 543.450 415.050 544.050 ;
        RECT 457.950 543.450 460.050 544.050 ;
        RECT 355.950 542.400 415.050 543.450 ;
        RECT 355.950 541.950 358.050 542.400 ;
        RECT 412.950 541.950 415.050 542.400 ;
        RECT 437.400 542.400 460.050 543.450 ;
        RECT 25.950 540.450 28.050 541.050 ;
        RECT 43.950 540.450 46.050 541.050 ;
        RECT 25.950 539.400 46.050 540.450 ;
        RECT 25.950 538.950 28.050 539.400 ;
        RECT 43.950 538.950 46.050 539.400 ;
        RECT 61.950 540.450 64.050 541.050 ;
        RECT 103.950 540.450 106.050 541.050 ;
        RECT 121.950 540.450 124.050 541.050 ;
        RECT 61.950 539.400 124.050 540.450 ;
        RECT 217.950 540.450 220.050 541.050 ;
        RECT 268.950 540.450 271.050 541.050 ;
        RECT 316.950 540.450 319.050 541.050 ;
        RECT 217.950 539.400 271.050 540.450 ;
        RECT 275.250 540.000 319.050 540.450 ;
        RECT 61.950 538.950 64.050 539.400 ;
        RECT 103.950 538.950 106.050 539.400 ;
        RECT 121.950 538.950 124.050 539.400 ;
        RECT 34.950 537.450 37.050 538.050 ;
        RECT 40.950 537.450 43.050 538.050 ;
        RECT 34.950 536.400 43.050 537.450 ;
        RECT 34.950 535.950 37.050 536.400 ;
        RECT 40.950 535.950 43.050 536.400 ;
        RECT 46.950 537.450 49.050 538.050 ;
        RECT 70.950 537.450 73.050 538.050 ;
        RECT 85.950 537.450 88.050 538.050 ;
        RECT 46.950 536.400 88.050 537.450 ;
        RECT 136.950 536.400 139.050 538.500 ;
        RECT 157.950 537.300 160.050 539.400 ;
        RECT 217.950 538.950 220.050 539.400 ;
        RECT 268.950 538.950 271.050 539.400 ;
        RECT 274.950 539.400 319.050 540.000 ;
        RECT 274.950 538.050 277.050 539.400 ;
        RECT 316.950 538.950 319.050 539.400 ;
        RECT 328.950 540.450 331.050 541.050 ;
        RECT 388.950 540.450 391.050 541.050 ;
        RECT 328.950 539.400 391.050 540.450 ;
        RECT 328.950 538.950 331.050 539.400 ;
        RECT 388.950 538.950 391.050 539.400 ;
        RECT 397.950 540.450 400.050 541.050 ;
        RECT 437.400 540.450 438.450 542.400 ;
        RECT 457.950 541.950 460.050 542.400 ;
        RECT 469.950 543.450 472.050 543.900 ;
        RECT 484.950 543.450 487.050 544.050 ;
        RECT 502.950 543.450 505.050 544.050 ;
        RECT 538.950 543.450 541.050 544.050 ;
        RECT 469.950 542.400 541.050 543.450 ;
        RECT 469.950 541.800 472.050 542.400 ;
        RECT 484.950 541.950 487.050 542.400 ;
        RECT 502.950 541.950 505.050 542.400 ;
        RECT 538.950 541.950 541.050 542.400 ;
        RECT 559.950 543.450 562.050 544.050 ;
        RECT 577.950 543.450 580.050 544.050 ;
        RECT 640.950 543.450 643.050 544.050 ;
        RECT 664.950 543.450 667.050 544.050 ;
        RECT 679.950 543.450 682.050 544.050 ;
        RECT 559.950 542.400 609.450 543.450 ;
        RECT 559.950 541.950 562.050 542.400 ;
        RECT 577.950 541.950 580.050 542.400 ;
        RECT 608.400 541.050 609.450 542.400 ;
        RECT 640.950 542.400 682.050 543.450 ;
        RECT 640.950 541.950 643.050 542.400 ;
        RECT 664.950 541.950 667.050 542.400 ;
        RECT 679.950 541.950 682.050 542.400 ;
        RECT 724.950 543.450 727.050 544.050 ;
        RECT 757.950 543.450 760.050 544.050 ;
        RECT 778.950 543.450 781.050 544.050 ;
        RECT 724.950 542.400 781.050 543.450 ;
        RECT 724.950 541.950 727.050 542.400 ;
        RECT 757.950 541.950 760.050 542.400 ;
        RECT 778.950 541.950 781.050 542.400 ;
        RECT 802.950 541.950 808.050 544.050 ;
        RECT 397.950 539.400 438.450 540.450 ;
        RECT 442.950 540.450 445.050 541.050 ;
        RECT 463.950 540.450 466.050 541.050 ;
        RECT 442.950 539.400 466.050 540.450 ;
        RECT 397.950 538.950 400.050 539.400 ;
        RECT 442.950 538.950 445.050 539.400 ;
        RECT 463.950 538.950 466.050 539.400 ;
        RECT 472.950 540.450 475.050 541.050 ;
        RECT 490.950 540.450 493.050 541.050 ;
        RECT 508.950 540.450 511.050 541.050 ;
        RECT 580.950 540.450 583.050 541.050 ;
        RECT 472.950 539.400 583.050 540.450 ;
        RECT 472.950 538.950 475.050 539.400 ;
        RECT 490.950 538.950 493.050 539.400 ;
        RECT 508.950 538.950 511.050 539.400 ;
        RECT 580.950 538.950 583.050 539.400 ;
        RECT 607.950 540.450 610.050 541.050 ;
        RECT 625.950 540.450 628.050 541.050 ;
        RECT 607.950 539.400 628.050 540.450 ;
        RECT 607.950 538.950 610.050 539.400 ;
        RECT 625.950 538.950 628.050 539.400 ;
        RECT 676.950 540.450 679.050 541.050 ;
        RECT 709.950 540.450 712.050 541.050 ;
        RECT 676.950 539.400 712.050 540.450 ;
        RECT 676.950 538.950 679.050 539.400 ;
        RECT 709.950 538.950 712.050 539.400 ;
        RECT 772.950 540.450 775.050 541.050 ;
        RECT 835.950 540.450 838.050 541.050 ;
        RECT 844.950 540.450 847.050 541.050 ;
        RECT 772.950 539.400 816.450 540.450 ;
        RECT 772.950 538.950 775.050 539.400 ;
        RECT 199.950 537.450 202.050 538.050 ;
        RECT 208.950 537.450 211.050 538.050 ;
        RECT 46.950 535.950 49.050 536.400 ;
        RECT 70.950 535.950 73.050 536.400 ;
        RECT 85.950 535.950 88.050 536.400 ;
        RECT 13.950 529.950 16.050 532.050 ;
        RECT 19.950 531.450 22.050 532.050 ;
        RECT 28.950 531.450 31.050 535.050 ;
        RECT 19.950 530.400 31.050 531.450 ;
        RECT 19.950 529.950 22.050 530.400 ;
        RECT 28.950 529.950 31.050 530.400 ;
        RECT 34.950 529.950 37.050 532.050 ;
        RECT 40.950 531.450 43.050 532.050 ;
        RECT 55.950 531.450 58.050 532.050 ;
        RECT 40.950 530.400 58.050 531.450 ;
        RECT 40.950 529.950 43.050 530.400 ;
        RECT 55.950 529.950 58.050 530.400 ;
        RECT 70.950 529.950 73.050 532.050 ;
        RECT 76.950 529.950 79.050 532.050 ;
        RECT 97.950 529.950 100.050 532.050 ;
        RECT 103.950 529.950 106.050 535.050 ;
        RECT 13.950 526.950 16.050 528.750 ;
        RECT 28.950 526.950 31.050 528.750 ;
        RECT 34.950 526.950 37.050 528.750 ;
        RECT 55.950 526.950 58.050 528.750 ;
        RECT 70.950 526.950 73.050 528.750 ;
        RECT 76.950 526.950 79.050 528.750 ;
        RECT 97.950 526.950 100.050 528.750 ;
        RECT 103.950 526.950 106.050 528.750 ;
        RECT 124.950 526.950 130.050 529.050 ;
        RECT 133.950 526.950 136.050 529.050 ;
        RECT 16.950 524.250 19.050 526.050 ;
        RECT 31.950 524.250 34.050 526.050 ;
        RECT 37.950 524.250 40.050 526.050 ;
        RECT 58.950 524.250 61.050 526.050 ;
        RECT 73.950 524.250 76.050 526.050 ;
        RECT 79.950 524.250 82.050 526.050 ;
        RECT 94.950 524.250 97.050 526.050 ;
        RECT 100.950 524.250 103.050 526.050 ;
        RECT 118.950 524.250 121.050 526.050 ;
        RECT 124.950 523.950 127.050 525.750 ;
        RECT 133.950 523.950 136.050 525.750 ;
        RECT 16.950 520.950 19.050 523.050 ;
        RECT 31.950 520.950 34.050 523.050 ;
        RECT 37.950 522.450 40.050 523.050 ;
        RECT 49.950 522.450 52.050 523.050 ;
        RECT 37.950 521.400 52.050 522.450 ;
        RECT 37.950 520.950 40.050 521.400 ;
        RECT 49.950 520.950 52.050 521.400 ;
        RECT 58.950 522.450 61.050 523.050 ;
        RECT 67.950 522.450 70.050 523.050 ;
        RECT 58.950 521.400 70.050 522.450 ;
        RECT 58.950 520.950 61.050 521.400 ;
        RECT 67.950 520.950 70.050 521.400 ;
        RECT 73.950 520.950 76.050 523.050 ;
        RECT 79.950 520.950 82.050 523.050 ;
        RECT 85.950 522.450 88.050 523.050 ;
        RECT 94.950 522.450 97.050 523.050 ;
        RECT 85.950 521.400 97.050 522.450 ;
        RECT 85.950 520.950 88.050 521.400 ;
        RECT 94.950 520.950 97.050 521.400 ;
        RECT 100.950 520.950 103.050 523.050 ;
        RECT 118.950 520.950 121.050 523.050 ;
        RECT 16.950 516.450 19.050 517.050 ;
        RECT 85.950 516.450 88.050 517.050 ;
        RECT 16.950 515.400 88.050 516.450 ;
        RECT 101.400 516.450 102.450 520.950 ;
        RECT 127.950 519.450 130.050 520.050 ;
        RECT 133.950 519.450 136.050 520.050 ;
        RECT 127.950 518.400 136.050 519.450 ;
        RECT 127.950 517.950 130.050 518.400 ;
        RECT 133.950 517.950 136.050 518.400 ;
        RECT 130.950 516.450 133.050 517.050 ;
        RECT 137.700 516.600 138.900 536.400 ;
        RECT 157.950 533.700 159.150 537.300 ;
        RECT 199.950 536.400 211.050 537.450 ;
        RECT 199.950 535.950 202.050 536.400 ;
        RECT 208.950 535.950 211.050 536.400 ;
        RECT 229.950 537.450 232.050 538.050 ;
        RECT 238.950 537.450 241.050 538.050 ;
        RECT 229.950 536.400 241.050 537.450 ;
        RECT 229.950 535.950 232.050 536.400 ;
        RECT 238.950 535.950 241.050 536.400 ;
        RECT 253.950 537.450 256.050 538.050 ;
        RECT 262.950 537.450 265.050 538.050 ;
        RECT 253.950 536.400 265.050 537.450 ;
        RECT 253.950 535.950 256.050 536.400 ;
        RECT 262.950 535.950 265.050 536.400 ;
        RECT 274.800 537.000 277.050 538.050 ;
        RECT 278.100 537.450 280.200 538.050 ;
        RECT 319.950 537.450 322.050 538.050 ;
        RECT 349.950 537.450 352.050 538.050 ;
        RECT 274.800 535.950 276.900 537.000 ;
        RECT 278.100 536.400 352.050 537.450 ;
        RECT 278.100 535.950 280.200 536.400 ;
        RECT 319.950 535.950 322.050 536.400 ;
        RECT 349.950 535.950 352.050 536.400 ;
        RECT 424.950 537.450 427.050 538.050 ;
        RECT 448.950 537.450 451.050 538.050 ;
        RECT 466.950 537.450 469.050 538.050 ;
        RECT 538.950 537.450 541.050 538.050 ;
        RECT 424.950 536.400 541.050 537.450 ;
        RECT 424.950 535.950 427.050 536.400 ;
        RECT 448.950 535.950 451.050 536.400 ;
        RECT 466.950 535.950 469.050 536.400 ;
        RECT 538.950 535.950 541.050 536.400 ;
        RECT 565.950 537.450 568.050 538.050 ;
        RECT 583.950 537.450 586.050 538.050 ;
        RECT 682.950 537.450 685.050 538.050 ;
        RECT 703.950 537.450 706.050 538.050 ;
        RECT 745.950 537.450 748.050 538.200 ;
        RECT 815.400 538.050 816.450 539.400 ;
        RECT 835.950 539.400 847.050 540.450 ;
        RECT 835.950 538.950 838.050 539.400 ;
        RECT 844.950 538.950 847.050 539.400 ;
        RECT 880.950 540.450 883.050 541.200 ;
        RECT 886.950 540.450 889.050 541.050 ;
        RECT 880.950 539.400 889.050 540.450 ;
        RECT 880.950 539.100 883.050 539.400 ;
        RECT 886.950 538.950 889.050 539.400 ;
        RECT 778.950 537.450 781.050 538.050 ;
        RECT 796.950 537.450 799.050 538.050 ;
        RECT 565.950 536.400 741.450 537.450 ;
        RECT 565.950 535.950 568.050 536.400 ;
        RECT 583.950 535.950 586.050 536.400 ;
        RECT 682.950 535.950 685.050 536.400 ;
        RECT 703.950 535.950 706.050 536.400 ;
        RECT 740.400 535.050 741.450 536.400 ;
        RECT 745.950 536.400 799.050 537.450 ;
        RECT 745.950 536.100 748.050 536.400 ;
        RECT 778.950 535.950 781.050 536.400 ;
        RECT 796.950 535.950 799.050 536.400 ;
        RECT 802.950 537.450 805.050 538.050 ;
        RECT 808.950 537.450 811.050 538.050 ;
        RECT 802.950 536.400 811.050 537.450 ;
        RECT 802.950 535.950 805.050 536.400 ;
        RECT 808.950 535.950 811.050 536.400 ;
        RECT 814.950 537.450 817.050 538.050 ;
        RECT 829.950 537.450 832.050 538.050 ;
        RECT 814.950 536.400 832.050 537.450 ;
        RECT 814.950 535.950 817.050 536.400 ;
        RECT 829.950 535.950 832.050 536.400 ;
        RECT 838.950 537.450 841.050 538.050 ;
        RECT 868.950 537.450 871.050 538.050 ;
        RECT 880.950 537.450 883.050 537.900 ;
        RECT 838.950 536.400 883.050 537.450 ;
        RECT 838.950 535.950 841.050 536.400 ;
        RECT 868.950 535.950 871.050 536.400 ;
        RECT 880.950 535.800 883.050 536.400 ;
        RECT 169.950 534.450 172.050 535.050 ;
        RECT 382.950 534.450 385.050 535.050 ;
        RECT 157.950 531.600 160.050 533.700 ;
        RECT 169.950 533.400 181.050 534.450 ;
        RECT 169.950 532.950 172.050 533.400 ;
        RECT 142.950 526.950 145.050 529.050 ;
        RECT 142.950 523.950 145.050 525.750 ;
        RECT 101.400 515.400 133.050 516.450 ;
        RECT 16.950 514.950 19.050 515.400 ;
        RECT 85.950 514.950 88.050 515.400 ;
        RECT 130.950 514.950 133.050 515.400 ;
        RECT 136.950 514.500 139.050 516.600 ;
        RECT 142.950 516.450 145.050 517.050 ;
        RECT 151.950 516.450 154.050 517.050 ;
        RECT 142.950 515.400 154.050 516.450 ;
        RECT 142.950 514.950 145.050 515.400 ;
        RECT 151.950 514.950 154.050 515.400 ;
        RECT 157.950 516.600 159.150 531.600 ;
        RECT 178.950 529.950 181.050 533.400 ;
        RECT 371.400 533.400 385.050 534.450 ;
        RECT 184.950 529.950 187.050 532.050 ;
        RECT 208.950 529.950 211.050 532.050 ;
        RECT 223.950 529.950 226.050 532.050 ;
        RECT 229.950 529.950 232.050 532.050 ;
        RECT 247.950 529.950 250.050 532.050 ;
        RECT 253.950 529.950 256.050 532.050 ;
        RECT 274.950 529.950 277.050 532.050 ;
        RECT 280.950 529.950 283.050 532.050 ;
        RECT 298.950 529.950 301.050 532.050 ;
        RECT 304.950 529.950 307.050 532.050 ;
        RECT 316.950 529.950 319.050 532.050 ;
        RECT 322.950 529.950 325.050 532.050 ;
        RECT 343.950 529.950 346.050 532.050 ;
        RECT 349.950 529.950 352.050 532.050 ;
        RECT 371.400 529.050 372.450 533.400 ;
        RECT 382.950 532.950 385.050 533.400 ;
        RECT 544.950 534.450 547.050 535.050 ;
        RECT 553.950 534.450 556.050 535.050 ;
        RECT 544.950 533.400 556.050 534.450 ;
        RECT 544.950 532.950 547.050 533.400 ;
        RECT 553.950 532.950 556.050 533.400 ;
        RECT 739.950 534.450 742.050 535.050 ;
        RECT 745.950 534.450 748.050 534.900 ;
        RECT 739.950 533.400 748.050 534.450 ;
        RECT 739.950 532.950 742.050 533.400 ;
        RECT 745.950 532.800 748.050 533.400 ;
        RECT 892.950 532.950 895.050 538.050 ;
        RECT 898.950 537.450 901.050 538.050 ;
        RECT 910.950 537.450 913.050 538.050 ;
        RECT 898.950 536.400 913.050 537.450 ;
        RECT 898.950 535.950 901.050 536.400 ;
        RECT 910.950 535.950 913.050 536.400 ;
        RECT 418.950 529.950 421.050 532.050 ;
        RECT 424.950 529.950 427.050 532.050 ;
        RECT 442.950 529.950 445.050 532.050 ;
        RECT 448.950 529.950 451.050 532.050 ;
        RECT 466.950 529.950 469.050 532.050 ;
        RECT 472.950 529.950 475.050 532.050 ;
        RECT 484.950 531.450 489.000 532.050 ;
        RECT 490.950 531.450 493.050 532.050 ;
        RECT 484.950 530.400 493.050 531.450 ;
        RECT 484.950 529.950 489.000 530.400 ;
        RECT 490.950 529.950 493.050 530.400 ;
        RECT 496.950 529.950 499.050 532.050 ;
        RECT 508.950 529.950 511.050 532.050 ;
        RECT 514.950 529.950 517.050 532.050 ;
        RECT 535.950 529.950 538.050 532.050 ;
        RECT 541.950 529.950 544.050 532.050 ;
        RECT 562.950 529.950 565.050 532.050 ;
        RECT 568.950 529.950 571.050 532.050 ;
        RECT 580.950 529.950 583.050 532.050 ;
        RECT 586.950 529.950 589.050 532.050 ;
        RECT 607.950 531.450 610.050 532.050 ;
        RECT 622.950 531.450 625.050 532.050 ;
        RECT 607.950 530.400 625.050 531.450 ;
        RECT 607.950 529.950 610.050 530.400 ;
        RECT 622.950 529.950 625.050 530.400 ;
        RECT 628.950 529.950 631.050 532.050 ;
        RECT 634.950 529.950 637.050 532.050 ;
        RECT 652.950 529.950 655.050 532.050 ;
        RECT 658.950 531.450 661.050 532.050 ;
        RECT 670.950 531.450 673.050 532.050 ;
        RECT 658.950 530.400 673.050 531.450 ;
        RECT 658.950 529.950 661.050 530.400 ;
        RECT 670.950 529.950 673.050 530.400 ;
        RECT 676.950 529.950 679.050 532.050 ;
        RECT 682.950 529.950 685.050 532.050 ;
        RECT 697.950 529.950 700.050 532.050 ;
        RECT 703.950 529.950 706.050 532.050 ;
        RECT 718.950 529.950 721.050 532.050 ;
        RECT 724.950 531.450 727.050 532.050 ;
        RECT 729.000 531.450 733.050 532.050 ;
        RECT 724.950 530.400 733.050 531.450 ;
        RECT 724.950 529.950 727.050 530.400 ;
        RECT 729.000 529.950 733.050 530.400 ;
        RECT 772.950 529.950 775.050 532.050 ;
        RECT 778.950 529.950 781.050 532.050 ;
        RECT 793.950 531.450 796.050 532.050 ;
        RECT 802.950 531.450 805.050 532.050 ;
        RECT 793.950 530.400 805.050 531.450 ;
        RECT 793.950 529.950 796.050 530.400 ;
        RECT 802.950 529.950 805.050 530.400 ;
        RECT 808.950 529.950 811.050 532.050 ;
        RECT 814.950 529.950 817.050 532.050 ;
        RECT 835.950 531.450 838.050 532.050 ;
        RECT 850.950 531.450 853.050 532.050 ;
        RECT 835.950 530.400 853.050 531.450 ;
        RECT 835.950 529.950 838.050 530.400 ;
        RECT 850.950 529.950 853.050 530.400 ;
        RECT 856.950 529.950 859.050 532.050 ;
        RECT 862.950 529.950 865.050 532.050 ;
        RECT 874.950 529.950 877.050 532.050 ;
        RECT 880.950 529.950 883.050 532.050 ;
        RECT 889.950 531.450 892.050 532.050 ;
        RECT 901.950 531.450 904.050 532.050 ;
        RECT 889.950 530.400 904.050 531.450 ;
        RECT 889.950 529.950 892.050 530.400 ;
        RECT 901.950 529.950 904.050 530.400 ;
        RECT 178.950 526.950 181.050 528.750 ;
        RECT 184.950 526.950 187.050 528.750 ;
        RECT 202.950 526.950 205.050 528.750 ;
        RECT 208.950 526.950 211.050 528.750 ;
        RECT 223.950 526.950 226.050 528.750 ;
        RECT 229.950 526.950 232.050 528.750 ;
        RECT 247.950 526.950 250.050 528.750 ;
        RECT 253.950 526.950 256.050 528.750 ;
        RECT 274.950 526.950 277.050 528.750 ;
        RECT 280.950 526.950 283.050 528.750 ;
        RECT 298.950 526.950 301.050 528.750 ;
        RECT 304.950 526.950 307.050 528.750 ;
        RECT 316.950 526.950 319.050 528.750 ;
        RECT 322.950 526.950 325.050 528.750 ;
        RECT 343.950 526.950 346.050 528.750 ;
        RECT 349.950 526.950 352.050 528.750 ;
        RECT 364.950 526.950 367.050 529.050 ;
        RECT 370.950 526.950 373.050 529.050 ;
        RECT 376.950 526.950 379.050 529.050 ;
        RECT 394.950 526.950 400.050 529.050 ;
        RECT 418.950 526.950 421.050 528.750 ;
        RECT 424.950 526.950 427.050 528.750 ;
        RECT 442.950 526.950 445.050 528.750 ;
        RECT 448.950 526.950 451.050 528.750 ;
        RECT 466.950 526.950 469.050 528.750 ;
        RECT 472.950 526.950 475.050 528.750 ;
        RECT 490.950 526.950 493.050 528.750 ;
        RECT 496.950 526.950 499.050 528.750 ;
        RECT 508.950 526.950 511.050 528.750 ;
        RECT 514.950 526.950 517.050 528.750 ;
        RECT 535.950 526.950 538.050 528.750 ;
        RECT 541.950 526.950 544.050 528.750 ;
        RECT 562.950 526.950 565.050 528.750 ;
        RECT 568.950 526.950 571.050 528.750 ;
        RECT 580.950 526.950 583.050 528.750 ;
        RECT 586.950 526.950 589.050 528.750 ;
        RECT 607.950 526.950 610.050 528.750 ;
        RECT 628.950 526.950 631.050 528.750 ;
        RECT 634.950 526.950 637.050 528.750 ;
        RECT 645.000 528.450 649.050 529.050 ;
        RECT 644.400 526.950 649.050 528.450 ;
        RECT 652.950 526.950 655.050 528.750 ;
        RECT 658.950 526.950 661.050 528.750 ;
        RECT 676.950 526.950 679.050 528.750 ;
        RECT 682.950 526.950 685.050 528.750 ;
        RECT 697.950 526.950 700.050 528.750 ;
        RECT 703.950 526.950 706.050 528.750 ;
        RECT 718.950 526.950 721.050 528.750 ;
        RECT 724.950 526.950 727.050 528.750 ;
        RECT 742.950 526.950 745.050 529.050 ;
        RECT 748.950 526.950 751.050 529.050 ;
        RECT 754.950 526.950 757.050 529.050 ;
        RECT 772.950 526.950 775.050 528.750 ;
        RECT 778.950 526.950 781.050 528.750 ;
        RECT 793.950 526.950 796.050 528.750 ;
        RECT 808.950 526.950 811.050 528.750 ;
        RECT 814.950 526.950 817.050 528.750 ;
        RECT 835.950 526.950 838.050 528.750 ;
        RECT 856.950 526.950 859.050 528.750 ;
        RECT 862.950 526.950 865.050 528.750 ;
        RECT 874.950 526.950 877.050 528.750 ;
        RECT 880.950 526.950 883.050 528.750 ;
        RECT 901.950 526.950 904.050 528.750 ;
        RECT 160.950 524.250 163.050 526.050 ;
        RECT 175.950 524.250 178.050 526.050 ;
        RECT 181.950 524.250 184.050 526.050 ;
        RECT 205.950 524.250 208.050 526.050 ;
        RECT 226.950 524.250 229.050 526.050 ;
        RECT 232.950 524.250 235.050 526.050 ;
        RECT 250.950 524.250 253.050 526.050 ;
        RECT 256.950 524.250 259.050 526.050 ;
        RECT 271.950 524.250 274.050 526.050 ;
        RECT 277.950 524.250 280.050 526.050 ;
        RECT 295.950 524.250 298.050 526.050 ;
        RECT 301.950 524.250 304.050 526.050 ;
        RECT 319.950 524.250 322.050 526.050 ;
        RECT 325.950 524.250 328.050 526.050 ;
        RECT 340.950 524.250 343.050 526.050 ;
        RECT 346.950 524.250 349.050 526.050 ;
        RECT 364.950 523.950 367.050 525.750 ;
        RECT 370.950 523.950 373.050 525.750 ;
        RECT 376.950 523.950 379.050 525.750 ;
        RECT 394.950 523.950 397.050 525.750 ;
        RECT 400.950 524.250 403.050 526.050 ;
        RECT 415.950 524.250 418.050 526.050 ;
        RECT 421.950 524.250 424.050 526.050 ;
        RECT 439.950 524.250 442.050 526.050 ;
        RECT 445.950 524.250 448.050 526.050 ;
        RECT 463.950 524.250 466.050 526.050 ;
        RECT 469.950 524.250 472.050 526.050 ;
        RECT 487.950 524.250 490.050 526.050 ;
        RECT 493.950 524.250 496.050 526.050 ;
        RECT 511.950 524.250 514.050 526.050 ;
        RECT 517.950 524.250 520.050 526.050 ;
        RECT 538.950 524.250 541.050 526.050 ;
        RECT 544.950 524.250 547.050 526.050 ;
        RECT 559.950 524.250 562.050 526.050 ;
        RECT 565.950 524.250 568.050 526.050 ;
        RECT 583.950 524.250 586.050 526.050 ;
        RECT 589.950 524.250 592.050 526.050 ;
        RECT 604.950 524.250 607.050 526.050 ;
        RECT 625.950 524.250 628.050 526.050 ;
        RECT 631.950 524.250 634.050 526.050 ;
        RECT 637.950 525.450 640.050 526.050 ;
        RECT 644.400 525.450 645.450 526.950 ;
        RECT 637.950 524.400 645.450 525.450 ;
        RECT 637.950 523.950 640.050 524.400 ;
        RECT 649.950 524.250 652.050 526.050 ;
        RECT 655.950 524.250 658.050 526.050 ;
        RECT 673.950 524.250 676.050 526.050 ;
        RECT 679.950 524.250 682.050 526.050 ;
        RECT 694.950 524.250 697.050 526.050 ;
        RECT 700.950 524.250 703.050 526.050 ;
        RECT 721.950 524.250 724.050 526.050 ;
        RECT 742.950 523.950 745.050 525.750 ;
        RECT 748.950 523.950 751.050 525.750 ;
        RECT 754.950 523.950 757.050 525.750 ;
        RECT 769.950 524.250 772.050 526.050 ;
        RECT 775.950 524.250 778.050 526.050 ;
        RECT 796.950 524.250 799.050 526.050 ;
        RECT 811.950 524.250 814.050 526.050 ;
        RECT 817.950 524.250 820.050 526.050 ;
        RECT 838.950 524.250 841.050 526.050 ;
        RECT 853.950 524.250 856.050 526.050 ;
        RECT 859.950 524.250 862.050 526.050 ;
        RECT 877.950 524.250 880.050 526.050 ;
        RECT 883.950 524.250 886.050 526.050 ;
        RECT 898.950 524.250 901.050 526.050 ;
        RECT 160.950 520.950 163.050 523.050 ;
        RECT 175.950 520.950 178.050 523.050 ;
        RECT 181.950 517.950 184.050 523.050 ;
        RECT 187.950 522.450 190.050 523.050 ;
        RECT 205.950 522.450 208.050 523.050 ;
        RECT 187.950 521.400 208.050 522.450 ;
        RECT 187.950 520.950 190.050 521.400 ;
        RECT 205.950 520.950 208.050 521.400 ;
        RECT 226.950 520.950 229.050 523.050 ;
        RECT 232.950 520.950 235.050 523.050 ;
        RECT 238.950 522.450 241.050 523.050 ;
        RECT 244.950 522.450 247.050 523.050 ;
        RECT 238.950 521.400 247.050 522.450 ;
        RECT 238.950 520.950 241.050 521.400 ;
        RECT 244.950 520.950 247.050 521.400 ;
        RECT 250.950 517.950 253.050 523.050 ;
        RECT 256.950 520.950 259.050 523.050 ;
        RECT 262.950 522.450 265.050 523.050 ;
        RECT 271.950 522.450 274.050 523.050 ;
        RECT 262.950 521.400 274.050 522.450 ;
        RECT 262.950 520.950 265.050 521.400 ;
        RECT 271.950 520.950 274.050 521.400 ;
        RECT 277.950 520.950 280.050 523.050 ;
        RECT 295.950 520.950 298.050 523.050 ;
        RECT 301.950 520.950 304.050 523.050 ;
        RECT 319.950 520.950 322.050 523.050 ;
        RECT 157.950 514.500 160.050 516.600 ;
        RECT 163.950 516.450 166.050 517.050 ;
        RECT 292.950 516.450 295.050 517.050 ;
        RECT 163.950 515.400 295.050 516.450 ;
        RECT 296.400 516.450 297.450 520.950 ;
        RECT 325.950 517.950 328.050 523.050 ;
        RECT 340.950 520.950 343.050 523.050 ;
        RECT 346.950 522.450 349.050 523.050 ;
        RECT 361.950 522.450 364.050 523.050 ;
        RECT 346.950 521.400 364.050 522.450 ;
        RECT 346.950 520.950 349.050 521.400 ;
        RECT 361.950 520.950 364.050 521.400 ;
        RECT 367.950 521.250 370.050 523.050 ;
        RECT 373.950 521.250 376.050 523.050 ;
        RECT 400.950 520.950 403.050 523.050 ;
        RECT 409.950 522.450 414.000 523.050 ;
        RECT 415.950 522.450 418.050 523.050 ;
        RECT 409.950 521.400 418.050 522.450 ;
        RECT 409.950 520.950 414.000 521.400 ;
        RECT 415.950 520.950 418.050 521.400 ;
        RECT 421.950 520.950 424.050 523.050 ;
        RECT 430.950 522.450 433.050 523.050 ;
        RECT 439.950 522.450 442.050 523.050 ;
        RECT 430.950 521.400 442.050 522.450 ;
        RECT 430.950 520.950 433.050 521.400 ;
        RECT 439.950 520.950 442.050 521.400 ;
        RECT 445.950 520.950 448.050 523.050 ;
        RECT 463.950 520.950 466.050 523.050 ;
        RECT 469.950 520.950 472.050 523.050 ;
        RECT 367.950 517.950 370.050 520.050 ;
        RECT 373.950 517.950 376.050 520.050 ;
        RECT 337.950 516.450 340.050 517.050 ;
        RECT 296.400 515.400 340.050 516.450 ;
        RECT 163.950 514.950 166.050 515.400 ;
        RECT 292.950 514.950 295.050 515.400 ;
        RECT 337.950 514.950 340.050 515.400 ;
        RECT 442.950 516.450 445.050 517.050 ;
        RECT 464.400 516.450 465.450 520.950 ;
        RECT 487.950 517.950 490.050 523.050 ;
        RECT 493.950 520.950 496.050 523.050 ;
        RECT 511.950 520.950 514.050 523.050 ;
        RECT 517.950 522.450 520.050 523.050 ;
        RECT 532.950 522.450 535.050 523.050 ;
        RECT 517.950 521.400 535.050 522.450 ;
        RECT 517.950 520.950 520.050 521.400 ;
        RECT 532.950 520.950 535.050 521.400 ;
        RECT 538.950 520.950 541.050 523.050 ;
        RECT 544.950 520.950 547.050 523.050 ;
        RECT 550.950 522.450 553.050 523.050 ;
        RECT 559.950 522.450 562.050 523.050 ;
        RECT 550.950 521.400 562.050 522.450 ;
        RECT 550.950 520.950 553.050 521.400 ;
        RECT 559.950 520.950 562.050 521.400 ;
        RECT 565.950 520.950 568.050 523.050 ;
        RECT 583.950 520.950 586.050 523.050 ;
        RECT 589.950 522.450 592.050 523.050 ;
        RECT 598.950 522.450 601.050 523.050 ;
        RECT 589.950 521.400 601.050 522.450 ;
        RECT 589.950 520.950 592.050 521.400 ;
        RECT 598.950 520.950 601.050 521.400 ;
        RECT 604.950 520.950 607.050 523.050 ;
        RECT 610.950 522.450 613.050 523.050 ;
        RECT 625.950 522.450 628.050 523.050 ;
        RECT 610.950 521.400 628.050 522.450 ;
        RECT 610.950 520.950 613.050 521.400 ;
        RECT 625.950 520.950 628.050 521.400 ;
        RECT 631.950 520.950 634.050 523.050 ;
        RECT 646.950 520.950 652.050 523.050 ;
        RECT 655.950 520.950 658.050 523.050 ;
        RECT 670.950 520.950 676.050 523.050 ;
        RECT 679.950 520.950 682.050 523.050 ;
        RECT 694.950 520.950 697.050 523.050 ;
        RECT 700.950 522.450 703.050 523.050 ;
        RECT 709.950 522.450 712.050 523.050 ;
        RECT 721.950 522.450 724.050 523.050 ;
        RECT 700.950 521.400 708.450 522.450 ;
        RECT 700.950 520.950 703.050 521.400 ;
        RECT 496.950 516.450 499.050 517.050 ;
        RECT 442.950 515.400 499.050 516.450 ;
        RECT 442.950 514.950 445.050 515.400 ;
        RECT 496.950 514.950 499.050 515.400 ;
        RECT 502.950 516.450 505.050 517.050 ;
        RECT 511.950 516.450 514.050 517.050 ;
        RECT 502.950 515.400 514.050 516.450 ;
        RECT 539.400 516.450 540.450 520.950 ;
        RECT 637.950 517.950 643.050 520.050 ;
        RECT 658.950 519.450 661.050 520.050 ;
        RECT 664.950 519.450 667.050 520.050 ;
        RECT 658.950 518.400 667.050 519.450 ;
        RECT 707.400 519.450 708.450 521.400 ;
        RECT 709.950 521.400 724.050 522.450 ;
        RECT 709.950 520.950 712.050 521.400 ;
        RECT 721.950 520.950 724.050 521.400 ;
        RECT 745.950 521.250 748.050 523.050 ;
        RECT 751.950 521.250 754.050 523.050 ;
        RECT 769.950 522.450 772.050 523.050 ;
        RECT 758.400 521.400 772.050 522.450 ;
        RECT 712.950 519.450 715.050 520.050 ;
        RECT 707.400 518.400 715.050 519.450 ;
        RECT 658.950 517.950 661.050 518.400 ;
        RECT 664.950 517.950 667.050 518.400 ;
        RECT 712.950 517.950 715.050 518.400 ;
        RECT 745.950 517.950 748.050 520.050 ;
        RECT 751.950 519.450 754.050 520.050 ;
        RECT 758.400 519.450 759.450 521.400 ;
        RECT 769.950 520.950 772.050 521.400 ;
        RECT 775.950 520.950 778.050 523.050 ;
        RECT 796.950 520.950 799.050 523.050 ;
        RECT 811.950 520.950 814.050 523.050 ;
        RECT 817.950 522.450 820.050 523.050 ;
        RECT 832.950 522.450 835.050 523.050 ;
        RECT 817.950 521.400 835.050 522.450 ;
        RECT 817.950 520.950 820.050 521.400 ;
        RECT 832.950 520.950 835.050 521.400 ;
        RECT 838.950 520.950 841.050 523.050 ;
        RECT 751.950 518.400 759.450 519.450 ;
        RECT 751.950 517.950 754.050 518.400 ;
        RECT 853.950 517.950 856.050 523.050 ;
        RECT 859.950 520.950 862.050 523.050 ;
        RECT 865.950 522.450 868.050 523.050 ;
        RECT 877.950 522.450 880.050 523.050 ;
        RECT 865.950 521.400 880.050 522.450 ;
        RECT 865.950 520.950 868.050 521.400 ;
        RECT 877.950 520.950 880.050 521.400 ;
        RECT 883.950 517.950 886.050 523.050 ;
        RECT 898.950 520.950 901.050 523.050 ;
        RECT 592.950 516.450 595.050 517.050 ;
        RECT 539.400 515.400 595.050 516.450 ;
        RECT 502.950 514.950 505.050 515.400 ;
        RECT 511.950 514.950 514.050 515.400 ;
        RECT 592.950 514.950 595.050 515.400 ;
        RECT 598.950 516.450 601.050 517.050 ;
        RECT 679.950 516.450 682.050 517.050 ;
        RECT 739.950 516.450 742.050 517.050 ;
        RECT 598.950 515.400 742.050 516.450 ;
        RECT 598.950 514.950 601.050 515.400 ;
        RECT 679.950 514.950 682.050 515.400 ;
        RECT 739.950 514.950 742.050 515.400 ;
        RECT 811.950 516.450 814.050 517.050 ;
        RECT 826.950 516.450 829.050 517.050 ;
        RECT 811.950 515.400 829.050 516.450 ;
        RECT 811.950 514.950 814.050 515.400 ;
        RECT 826.950 514.950 829.050 515.400 ;
        RECT 841.950 516.450 844.050 517.050 ;
        RECT 847.950 516.450 850.050 517.050 ;
        RECT 841.950 515.400 850.050 516.450 ;
        RECT 841.950 514.950 844.050 515.400 ;
        RECT 847.950 514.950 850.050 515.400 ;
        RECT 40.950 511.950 46.050 514.050 ;
        RECT 166.950 513.450 169.050 514.050 ;
        RECT 175.950 513.450 178.050 514.050 ;
        RECT 217.950 513.450 220.050 514.050 ;
        RECT 166.950 512.400 220.050 513.450 ;
        RECT 166.950 511.950 169.050 512.400 ;
        RECT 175.950 511.950 178.050 512.400 ;
        RECT 217.950 511.950 220.050 512.400 ;
        RECT 268.950 513.450 271.050 514.050 ;
        RECT 307.950 513.450 310.050 514.050 ;
        RECT 325.950 513.450 328.050 514.050 ;
        RECT 358.800 513.450 360.900 514.050 ;
        RECT 268.950 512.400 306.450 513.450 ;
        RECT 268.950 511.950 271.050 512.400 ;
        RECT 49.950 510.450 52.050 511.050 ;
        RECT 238.950 510.450 241.050 511.050 ;
        RECT 298.950 510.450 301.050 511.050 ;
        RECT 49.950 509.400 241.050 510.450 ;
        RECT 49.950 508.950 52.050 509.400 ;
        RECT 238.950 508.950 241.050 509.400 ;
        RECT 245.400 509.400 301.050 510.450 ;
        RECT 305.400 510.450 306.450 512.400 ;
        RECT 307.950 512.400 360.900 513.450 ;
        RECT 307.950 511.950 310.050 512.400 ;
        RECT 325.950 511.950 328.050 512.400 ;
        RECT 358.800 511.950 360.900 512.400 ;
        RECT 362.100 513.450 364.200 514.050 ;
        RECT 418.950 513.450 421.050 514.050 ;
        RECT 454.800 513.450 456.900 514.050 ;
        RECT 362.100 512.400 456.900 513.450 ;
        RECT 362.100 511.950 364.200 512.400 ;
        RECT 418.950 511.950 421.050 512.400 ;
        RECT 454.800 511.950 456.900 512.400 ;
        RECT 458.100 513.450 460.200 514.050 ;
        RECT 664.950 513.450 667.050 514.050 ;
        RECT 458.100 512.400 667.050 513.450 ;
        RECT 458.100 511.950 460.200 512.400 ;
        RECT 664.950 511.950 667.050 512.400 ;
        RECT 718.950 513.450 721.050 514.050 ;
        RECT 724.950 513.450 727.050 514.050 ;
        RECT 718.950 512.400 727.050 513.450 ;
        RECT 718.950 511.950 721.050 512.400 ;
        RECT 724.950 511.950 727.050 512.400 ;
        RECT 763.950 513.450 766.050 514.050 ;
        RECT 781.950 513.450 784.050 514.050 ;
        RECT 763.950 512.400 784.050 513.450 ;
        RECT 763.950 511.950 766.050 512.400 ;
        RECT 781.950 511.950 784.050 512.400 ;
        RECT 802.950 511.950 808.050 514.050 ;
        RECT 880.950 513.450 883.050 514.050 ;
        RECT 892.950 513.450 895.050 517.050 ;
        RECT 880.950 512.400 895.050 513.450 ;
        RECT 880.950 511.950 883.050 512.400 ;
        RECT 892.950 511.950 895.050 512.400 ;
        RECT 316.950 510.450 319.050 511.050 ;
        RECT 355.950 510.450 358.050 511.050 ;
        RECT 305.400 509.400 358.050 510.450 ;
        RECT 79.950 507.450 82.050 508.050 ;
        RECT 109.950 507.450 112.050 508.050 ;
        RECT 79.950 506.400 112.050 507.450 ;
        RECT 79.950 505.950 82.050 506.400 ;
        RECT 109.950 505.950 112.050 506.400 ;
        RECT 127.950 507.450 130.050 508.050 ;
        RECT 181.950 507.450 184.050 508.050 ;
        RECT 127.950 506.400 184.050 507.450 ;
        RECT 127.950 505.950 130.050 506.400 ;
        RECT 181.950 505.950 184.050 506.400 ;
        RECT 199.950 507.450 202.050 508.050 ;
        RECT 245.400 507.450 246.450 509.400 ;
        RECT 298.950 508.950 301.050 509.400 ;
        RECT 316.950 508.950 319.050 509.400 ;
        RECT 355.950 508.950 358.050 509.400 ;
        RECT 376.950 510.450 379.050 511.050 ;
        RECT 430.950 510.450 433.050 511.050 ;
        RECT 376.950 509.400 433.050 510.450 ;
        RECT 376.950 508.950 379.050 509.400 ;
        RECT 430.950 508.950 433.050 509.400 ;
        RECT 445.950 510.450 448.050 511.050 ;
        RECT 502.950 510.450 505.050 511.050 ;
        RECT 445.950 509.400 505.050 510.450 ;
        RECT 445.950 508.950 448.050 509.400 ;
        RECT 502.950 508.950 505.050 509.400 ;
        RECT 553.950 510.450 556.050 511.050 ;
        RECT 610.950 510.450 613.050 511.050 ;
        RECT 553.950 509.400 613.050 510.450 ;
        RECT 553.950 508.950 556.050 509.400 ;
        RECT 610.950 508.950 613.050 509.400 ;
        RECT 775.950 510.450 778.050 511.050 ;
        RECT 811.950 510.450 814.050 511.050 ;
        RECT 775.950 509.400 814.050 510.450 ;
        RECT 775.950 508.950 778.050 509.400 ;
        RECT 811.950 508.950 814.050 509.400 ;
        RECT 199.950 506.400 246.450 507.450 ;
        RECT 250.950 507.450 253.050 508.050 ;
        RECT 343.950 507.450 346.050 508.050 ;
        RECT 250.950 506.400 346.050 507.450 ;
        RECT 199.950 505.950 202.050 506.400 ;
        RECT 250.950 505.950 253.050 506.400 ;
        RECT 343.950 505.950 346.050 506.400 ;
        RECT 373.950 507.450 376.050 508.050 ;
        RECT 469.950 507.450 472.050 508.050 ;
        RECT 505.950 507.450 508.050 508.050 ;
        RECT 373.950 506.400 508.050 507.450 ;
        RECT 373.950 505.950 376.050 506.400 ;
        RECT 469.950 505.950 472.050 506.400 ;
        RECT 505.950 505.950 508.050 506.400 ;
        RECT 532.950 507.450 535.050 508.050 ;
        RECT 544.950 507.450 547.050 508.050 ;
        RECT 532.950 506.400 547.050 507.450 ;
        RECT 532.950 505.950 535.050 506.400 ;
        RECT 544.950 505.950 547.050 506.400 ;
        RECT 739.950 507.450 742.050 508.050 ;
        RECT 748.950 507.450 751.050 508.050 ;
        RECT 739.950 506.400 751.050 507.450 ;
        RECT 739.950 505.950 742.050 506.400 ;
        RECT 748.950 505.950 751.050 506.400 ;
        RECT 760.950 507.450 763.050 508.050 ;
        RECT 787.950 507.450 790.050 508.050 ;
        RECT 760.950 506.400 790.050 507.450 ;
        RECT 760.950 505.950 763.050 506.400 ;
        RECT 787.950 505.950 790.050 506.400 ;
        RECT 904.950 507.450 907.050 508.200 ;
        RECT 910.950 507.450 913.050 508.050 ;
        RECT 904.950 506.400 913.050 507.450 ;
        RECT 904.950 506.100 907.050 506.400 ;
        RECT 910.950 505.950 913.050 506.400 ;
        RECT 40.950 504.450 43.050 505.050 ;
        RECT 52.950 504.450 55.050 505.050 ;
        RECT 40.950 503.400 55.050 504.450 ;
        RECT 40.950 502.950 43.050 503.400 ;
        RECT 52.950 502.950 55.050 503.400 ;
        RECT 94.950 504.450 97.050 505.050 ;
        RECT 103.950 504.450 106.050 505.050 ;
        RECT 94.950 503.400 106.050 504.450 ;
        RECT 94.950 502.950 97.050 503.400 ;
        RECT 103.950 502.950 106.050 503.400 ;
        RECT 124.950 504.450 127.050 505.050 ;
        RECT 130.950 504.450 133.050 505.050 ;
        RECT 124.950 503.400 133.050 504.450 ;
        RECT 124.950 502.950 127.050 503.400 ;
        RECT 130.950 502.950 133.050 503.400 ;
        RECT 388.950 504.450 391.050 505.050 ;
        RECT 394.950 504.450 397.050 505.050 ;
        RECT 388.950 503.400 397.050 504.450 ;
        RECT 388.950 502.950 391.050 503.400 ;
        RECT 394.950 502.950 397.050 503.400 ;
        RECT 430.950 504.450 433.050 505.050 ;
        RECT 460.950 504.450 463.050 505.050 ;
        RECT 430.950 503.400 463.050 504.450 ;
        RECT 430.950 502.950 433.050 503.400 ;
        RECT 460.950 502.950 463.050 503.400 ;
        RECT 478.950 504.450 481.050 505.050 ;
        RECT 484.950 504.450 487.050 505.050 ;
        RECT 478.950 503.400 487.050 504.450 ;
        RECT 478.950 502.950 481.050 503.400 ;
        RECT 484.950 502.950 487.050 503.400 ;
        RECT 535.950 504.450 538.050 505.050 ;
        RECT 571.950 504.450 574.050 505.050 ;
        RECT 535.950 503.400 574.050 504.450 ;
        RECT 535.950 502.950 538.050 503.400 ;
        RECT 571.950 502.950 574.050 503.400 ;
        RECT 607.950 504.450 610.050 505.050 ;
        RECT 646.950 504.450 649.050 505.050 ;
        RECT 607.950 503.400 649.050 504.450 ;
        RECT 607.950 502.950 610.050 503.400 ;
        RECT 646.950 502.950 649.050 503.400 ;
        RECT 652.950 504.450 655.050 505.050 ;
        RECT 658.950 504.450 661.050 505.050 ;
        RECT 652.950 503.400 661.050 504.450 ;
        RECT 652.950 502.950 655.050 503.400 ;
        RECT 658.950 502.950 661.050 503.400 ;
        RECT 724.950 504.450 727.050 505.050 ;
        RECT 724.950 503.400 771.450 504.450 ;
        RECT 724.950 502.950 727.050 503.400 ;
        RECT 7.950 501.450 10.050 502.050 ;
        RECT 19.950 501.450 22.050 502.050 ;
        RECT 37.950 501.450 40.050 502.050 ;
        RECT 7.950 500.400 40.050 501.450 ;
        RECT 7.950 499.950 10.050 500.400 ;
        RECT 19.950 499.950 22.050 500.400 ;
        RECT 37.950 499.950 40.050 500.400 ;
        RECT 52.950 501.450 55.050 502.050 ;
        RECT 58.950 501.450 61.050 502.050 ;
        RECT 52.950 500.400 61.050 501.450 ;
        RECT 52.950 499.950 55.050 500.400 ;
        RECT 58.950 499.950 61.050 500.400 ;
        RECT 109.950 501.450 112.050 502.050 ;
        RECT 127.950 501.450 130.050 502.050 ;
        RECT 109.950 500.400 130.050 501.450 ;
        RECT 103.950 496.950 106.050 499.050 ;
        RECT 109.950 496.950 112.050 500.400 ;
        RECT 127.950 499.950 130.050 500.400 ;
        RECT 205.950 501.450 208.050 502.050 ;
        RECT 214.950 501.450 217.050 502.050 ;
        RECT 205.950 500.400 217.050 501.450 ;
        RECT 220.950 500.400 223.050 502.500 ;
        RECT 241.950 500.400 244.050 502.500 ;
        RECT 292.950 500.400 295.050 502.500 ;
        RECT 313.950 500.400 316.050 502.500 ;
        RECT 770.400 502.050 771.450 503.400 ;
        RECT 820.950 502.950 826.050 505.050 ;
        RECT 841.950 504.450 844.050 505.050 ;
        RECT 883.950 504.450 886.050 505.050 ;
        RECT 841.950 503.400 886.050 504.450 ;
        RECT 841.950 502.950 844.050 503.400 ;
        RECT 883.950 502.950 886.050 503.400 ;
        RECT 898.950 504.450 901.050 505.050 ;
        RECT 904.950 504.450 907.050 504.900 ;
        RECT 898.950 503.400 907.050 504.450 ;
        RECT 898.950 502.950 901.050 503.400 ;
        RECT 904.950 502.800 907.050 503.400 ;
        RECT 349.950 501.450 352.050 502.050 ;
        RECT 358.950 501.450 361.050 502.050 ;
        RECT 349.950 500.400 361.050 501.450 ;
        RECT 205.950 499.950 208.050 500.400 ;
        RECT 214.950 499.950 217.050 500.400 ;
        RECT 10.950 493.950 16.050 496.050 ;
        RECT 19.950 493.950 22.050 496.050 ;
        RECT 37.950 493.950 40.050 496.050 ;
        RECT 43.950 493.950 46.050 496.050 ;
        RECT 58.950 493.950 61.050 496.050 ;
        RECT 82.950 495.450 85.050 496.050 ;
        RECT 94.950 495.450 97.050 496.050 ;
        RECT 82.950 494.400 97.050 495.450 ;
        RECT 82.950 493.950 85.050 494.400 ;
        RECT 94.950 493.950 97.050 494.400 ;
        RECT 103.950 493.950 106.050 495.750 ;
        RECT 109.950 493.950 112.050 495.750 ;
        RECT 124.950 493.950 127.050 496.050 ;
        RECT 130.950 495.450 133.050 496.050 ;
        RECT 145.950 495.450 148.050 496.050 ;
        RECT 130.950 494.400 148.050 495.450 ;
        RECT 130.950 493.950 133.050 494.400 ;
        RECT 145.950 493.950 148.050 494.400 ;
        RECT 211.950 493.950 214.050 496.050 ;
        RECT 13.950 490.950 16.050 492.750 ;
        RECT 19.950 490.950 22.050 492.750 ;
        RECT 37.950 490.950 40.050 492.750 ;
        RECT 43.950 490.950 46.050 492.750 ;
        RECT 58.950 490.950 61.050 492.750 ;
        RECT 82.950 490.950 85.050 492.750 ;
        RECT 100.950 491.250 103.050 493.050 ;
        RECT 106.950 491.250 109.050 493.050 ;
        RECT 112.950 491.250 115.050 493.050 ;
        RECT 124.950 490.950 127.050 492.750 ;
        RECT 145.950 490.950 148.050 492.750 ;
        RECT 151.950 491.250 154.050 493.050 ;
        RECT 169.950 491.250 172.050 493.050 ;
        RECT 190.950 491.250 193.050 493.050 ;
        RECT 211.950 490.950 214.050 492.750 ;
        RECT 217.950 491.250 220.050 493.050 ;
        RECT 16.950 488.250 19.050 490.050 ;
        RECT 22.950 488.250 25.050 490.050 ;
        RECT 34.950 488.250 37.050 490.050 ;
        RECT 40.950 488.250 43.050 490.050 ;
        RECT 61.950 488.250 64.050 490.050 ;
        RECT 79.950 488.250 82.050 490.050 ;
        RECT 85.950 488.250 88.050 490.050 ;
        RECT 100.950 487.950 103.050 490.050 ;
        RECT 16.950 484.950 19.050 487.050 ;
        RECT 22.950 484.950 25.050 487.050 ;
        RECT 34.950 484.950 37.050 487.050 ;
        RECT 40.950 484.950 43.050 487.050 ;
        RECT 61.950 481.950 64.050 487.050 ;
        RECT 79.950 484.950 82.050 487.050 ;
        RECT 85.950 486.450 88.050 487.050 ;
        RECT 85.950 485.400 96.450 486.450 ;
        RECT 85.950 484.950 88.050 485.400 ;
        RECT 43.950 480.450 46.050 481.050 ;
        RECT 80.400 480.450 81.450 484.950 ;
        RECT 95.400 483.450 96.450 485.400 ;
        RECT 106.950 484.950 109.050 490.050 ;
        RECT 112.950 487.950 118.050 490.050 ;
        RECT 121.950 488.250 124.050 490.050 ;
        RECT 127.950 488.250 130.050 490.050 ;
        RECT 142.950 488.250 145.050 490.050 ;
        RECT 151.950 489.450 154.050 490.050 ;
        RECT 160.950 489.450 163.050 490.050 ;
        RECT 151.950 488.400 163.050 489.450 ;
        RECT 151.950 487.950 154.050 488.400 ;
        RECT 160.950 487.950 163.050 488.400 ;
        RECT 169.950 489.450 172.050 490.050 ;
        RECT 174.000 489.450 178.050 490.050 ;
        RECT 169.950 488.400 178.050 489.450 ;
        RECT 169.950 487.950 172.050 488.400 ;
        RECT 174.000 487.950 178.050 488.400 ;
        RECT 208.950 488.250 211.050 490.050 ;
        RECT 217.950 487.950 220.050 490.050 ;
        RECT 121.950 484.950 124.050 487.050 ;
        RECT 127.950 484.950 130.050 487.050 ;
        RECT 142.950 484.950 145.050 487.050 ;
        RECT 208.950 484.950 211.050 487.050 ;
        RECT 100.950 483.450 103.050 484.050 ;
        RECT 95.400 482.400 103.050 483.450 ;
        RECT 100.950 481.950 103.050 482.400 ;
        RECT 94.950 480.450 97.050 481.050 ;
        RECT 43.950 479.400 97.050 480.450 ;
        RECT 43.950 478.950 46.050 479.400 ;
        RECT 94.950 478.950 97.050 479.400 ;
        RECT 115.950 480.450 118.050 481.050 ;
        RECT 121.950 480.450 124.050 481.050 ;
        RECT 115.950 479.400 124.050 480.450 ;
        RECT 115.950 478.950 118.050 479.400 ;
        RECT 121.950 478.950 124.050 479.400 ;
        RECT 184.950 480.450 187.050 481.050 ;
        RECT 209.400 480.450 210.450 484.950 ;
        RECT 221.700 480.600 222.900 500.400 ;
        RECT 226.950 491.250 229.050 493.050 ;
        RECT 226.950 487.950 229.050 490.050 ;
        RECT 241.950 485.400 243.150 500.400 ;
        RECT 244.950 495.450 247.050 496.050 ;
        RECT 253.950 495.450 256.050 496.050 ;
        RECT 244.950 494.400 256.050 495.450 ;
        RECT 244.950 493.950 247.050 494.400 ;
        RECT 253.950 493.950 256.050 494.400 ;
        RECT 259.950 493.950 262.050 496.050 ;
        RECT 283.950 495.450 286.050 496.050 ;
        RECT 289.950 495.450 292.050 496.050 ;
        RECT 283.950 494.400 292.050 495.450 ;
        RECT 283.950 493.950 286.050 494.400 ;
        RECT 289.950 493.950 292.050 494.400 ;
        RECT 244.950 490.950 247.050 492.750 ;
        RECT 259.950 490.950 262.050 492.750 ;
        RECT 283.950 490.950 286.050 492.750 ;
        RECT 289.950 490.950 292.050 492.750 ;
        RECT 262.950 488.250 265.050 490.050 ;
        RECT 280.950 488.250 283.050 490.050 ;
        RECT 241.950 483.300 244.050 485.400 ;
        RECT 262.950 484.950 265.050 487.050 ;
        RECT 280.950 484.950 283.050 487.050 ;
        RECT 293.850 485.400 295.050 500.400 ;
        RECT 307.950 491.250 310.050 493.050 ;
        RECT 292.950 483.300 295.050 485.400 ;
        RECT 307.950 484.950 310.050 490.050 ;
        RECT 184.950 479.400 210.450 480.450 ;
        RECT 184.950 478.950 187.050 479.400 ;
        RECT 220.950 478.500 223.050 480.600 ;
        RECT 241.950 479.700 243.150 483.300 ;
        RECT 262.950 480.450 265.050 481.050 ;
        RECT 271.950 480.450 274.050 481.050 ;
        RECT 16.950 477.450 19.050 478.050 ;
        RECT 40.950 477.450 43.050 478.050 ;
        RECT 61.950 477.450 64.050 478.050 ;
        RECT 16.950 476.400 64.050 477.450 ;
        RECT 16.950 475.950 19.050 476.400 ;
        RECT 40.950 475.950 43.050 476.400 ;
        RECT 61.950 475.950 64.050 476.400 ;
        RECT 94.950 477.450 97.050 478.050 ;
        RECT 142.950 477.450 145.050 478.050 ;
        RECT 241.950 477.600 244.050 479.700 ;
        RECT 262.950 479.400 274.050 480.450 ;
        RECT 262.950 478.950 265.050 479.400 ;
        RECT 271.950 478.950 274.050 479.400 ;
        RECT 280.950 480.450 283.050 481.050 ;
        RECT 286.950 480.450 289.050 481.050 ;
        RECT 280.950 479.400 289.050 480.450 ;
        RECT 293.850 479.700 295.050 483.300 ;
        RECT 314.100 480.600 315.300 500.400 ;
        RECT 349.950 499.950 352.050 500.400 ;
        RECT 358.950 499.950 361.050 500.400 ;
        RECT 424.950 501.450 427.050 502.050 ;
        RECT 487.950 501.450 490.050 502.050 ;
        RECT 523.950 501.450 526.050 502.050 ;
        RECT 565.950 501.450 568.050 502.050 ;
        RECT 424.950 500.400 568.050 501.450 ;
        RECT 424.950 499.950 427.050 500.400 ;
        RECT 487.950 499.950 490.050 500.400 ;
        RECT 523.950 499.950 526.050 500.400 ;
        RECT 565.950 499.950 568.050 500.400 ;
        RECT 592.950 501.450 595.050 502.050 ;
        RECT 625.950 501.450 628.050 502.050 ;
        RECT 592.950 500.400 628.050 501.450 ;
        RECT 592.950 499.950 595.050 500.400 ;
        RECT 625.950 499.950 628.050 500.400 ;
        RECT 757.950 501.450 760.050 502.050 ;
        RECT 763.950 501.450 766.050 502.050 ;
        RECT 757.950 500.400 766.050 501.450 ;
        RECT 757.950 499.950 760.050 500.400 ;
        RECT 763.950 499.950 766.050 500.400 ;
        RECT 769.950 501.450 772.050 502.050 ;
        RECT 832.950 501.450 835.050 502.050 ;
        RECT 769.950 500.400 835.050 501.450 ;
        RECT 769.950 499.950 772.050 500.400 ;
        RECT 832.950 499.950 835.050 500.400 ;
        RECT 853.950 501.450 856.050 502.050 ;
        RECT 877.950 501.450 880.050 502.050 ;
        RECT 895.950 501.450 898.050 502.050 ;
        RECT 853.950 500.400 898.050 501.450 ;
        RECT 853.950 499.950 856.050 500.400 ;
        RECT 877.950 499.950 880.050 500.400 ;
        RECT 895.950 499.950 898.050 500.400 ;
        RECT 382.950 496.950 385.050 499.050 ;
        RECT 388.950 496.950 391.050 499.050 ;
        RECT 646.950 496.950 649.050 499.050 ;
        RECT 652.950 496.950 655.050 499.050 ;
        RECT 721.950 498.450 724.050 499.050 ;
        RECT 727.950 498.450 730.050 499.050 ;
        RECT 721.950 497.400 730.050 498.450 ;
        RECT 721.950 496.950 724.050 497.400 ;
        RECT 727.950 496.950 730.050 497.400 ;
        RECT 733.950 496.950 736.050 499.050 ;
        RECT 739.950 496.950 742.050 499.050 ;
        RECT 337.950 493.950 340.050 496.050 ;
        RECT 358.950 493.950 361.050 496.050 ;
        RECT 364.950 495.450 367.050 496.050 ;
        RECT 376.950 495.450 379.050 496.050 ;
        RECT 364.950 494.400 379.050 495.450 ;
        RECT 364.950 493.950 367.050 494.400 ;
        RECT 376.950 493.950 379.050 494.400 ;
        RECT 382.950 493.950 385.050 495.750 ;
        RECT 388.950 493.950 391.050 495.750 ;
        RECT 394.950 495.450 397.050 496.050 ;
        RECT 403.950 495.450 406.050 496.050 ;
        RECT 394.950 494.400 406.050 495.450 ;
        RECT 394.950 493.950 397.050 494.400 ;
        RECT 403.950 493.950 406.050 494.400 ;
        RECT 409.950 495.450 412.050 496.050 ;
        RECT 427.950 495.450 430.050 496.050 ;
        RECT 409.950 494.400 430.050 495.450 ;
        RECT 409.950 493.950 412.050 494.400 ;
        RECT 427.950 493.950 430.050 494.400 ;
        RECT 433.950 495.450 436.050 496.050 ;
        RECT 438.000 495.450 442.050 496.050 ;
        RECT 433.950 494.400 442.050 495.450 ;
        RECT 433.950 493.950 436.050 494.400 ;
        RECT 438.000 493.950 442.050 494.400 ;
        RECT 454.950 493.950 457.050 496.050 ;
        RECT 469.950 493.950 472.050 496.050 ;
        RECT 475.950 495.450 478.050 496.050 ;
        RECT 484.800 495.450 486.900 496.050 ;
        RECT 475.950 494.400 486.900 495.450 ;
        RECT 475.950 493.950 478.050 494.400 ;
        RECT 484.800 493.950 486.900 494.400 ;
        RECT 488.100 495.450 492.000 496.050 ;
        RECT 493.950 495.450 496.050 496.050 ;
        RECT 488.100 494.400 496.050 495.450 ;
        RECT 488.100 493.950 492.000 494.400 ;
        RECT 493.950 493.950 496.050 494.400 ;
        RECT 499.950 493.950 502.050 496.050 ;
        RECT 505.950 495.450 508.050 496.050 ;
        RECT 517.950 495.450 520.050 496.050 ;
        RECT 505.950 494.400 520.050 495.450 ;
        RECT 505.950 493.950 508.050 494.400 ;
        RECT 517.950 493.950 520.050 494.400 ;
        RECT 523.950 493.950 526.050 496.050 ;
        RECT 538.950 493.950 541.050 496.050 ;
        RECT 556.950 493.950 559.050 496.050 ;
        RECT 562.950 495.450 565.050 496.050 ;
        RECT 580.950 495.450 583.050 496.050 ;
        RECT 562.950 494.400 583.050 495.450 ;
        RECT 562.950 493.950 565.050 494.400 ;
        RECT 580.950 493.950 583.050 494.400 ;
        RECT 586.950 495.450 589.050 496.050 ;
        RECT 595.950 495.450 598.050 496.050 ;
        RECT 586.950 494.400 598.050 495.450 ;
        RECT 586.950 493.950 589.050 494.400 ;
        RECT 595.950 493.950 598.050 494.400 ;
        RECT 601.950 493.950 604.050 496.050 ;
        RECT 607.950 495.450 610.050 496.050 ;
        RECT 616.950 495.450 619.050 496.050 ;
        RECT 607.950 494.400 619.050 495.450 ;
        RECT 607.950 493.950 610.050 494.400 ;
        RECT 616.950 493.950 619.050 494.400 ;
        RECT 628.950 495.450 631.050 496.050 ;
        RECT 640.950 495.450 643.050 496.050 ;
        RECT 628.950 494.400 643.050 495.450 ;
        RECT 628.950 493.950 631.050 494.400 ;
        RECT 640.950 493.950 643.050 494.400 ;
        RECT 646.950 493.950 649.050 495.750 ;
        RECT 652.950 493.950 655.050 495.750 ;
        RECT 658.950 495.450 661.050 496.050 ;
        RECT 670.950 495.450 673.050 496.050 ;
        RECT 658.950 494.400 673.050 495.450 ;
        RECT 658.950 493.950 661.050 494.400 ;
        RECT 670.950 493.950 673.050 494.400 ;
        RECT 685.950 493.950 688.050 496.050 ;
        RECT 691.950 495.450 694.050 496.050 ;
        RECT 700.800 495.450 702.900 496.050 ;
        RECT 691.950 494.400 702.900 495.450 ;
        RECT 691.950 493.950 694.050 494.400 ;
        RECT 700.800 493.950 702.900 494.400 ;
        RECT 704.100 495.450 706.200 496.050 ;
        RECT 712.950 495.450 715.050 496.050 ;
        RECT 704.100 494.400 715.050 495.450 ;
        RECT 704.100 493.950 706.200 494.400 ;
        RECT 712.950 493.950 715.050 494.400 ;
        RECT 718.950 493.950 721.050 496.050 ;
        RECT 733.950 493.950 736.050 495.750 ;
        RECT 739.950 493.950 742.050 495.750 ;
        RECT 745.950 495.450 748.050 496.050 ;
        RECT 757.950 495.450 760.050 496.050 ;
        RECT 745.950 494.400 760.050 495.450 ;
        RECT 745.950 493.950 748.050 494.400 ;
        RECT 757.950 493.950 760.050 494.400 ;
        RECT 763.950 493.950 766.050 496.050 ;
        RECT 784.950 495.450 787.050 496.050 ;
        RECT 796.950 495.450 799.050 496.050 ;
        RECT 784.950 494.400 799.050 495.450 ;
        RECT 784.950 493.950 787.050 494.400 ;
        RECT 796.950 493.950 799.050 494.400 ;
        RECT 805.950 493.950 808.050 496.050 ;
        RECT 820.950 495.450 825.000 496.050 ;
        RECT 826.950 495.450 829.050 496.050 ;
        RECT 820.950 494.400 829.050 495.450 ;
        RECT 820.950 493.950 825.000 494.400 ;
        RECT 826.950 493.950 829.050 494.400 ;
        RECT 832.950 495.450 835.050 496.050 ;
        RECT 847.950 495.450 850.050 496.050 ;
        RECT 832.950 494.400 850.050 495.450 ;
        RECT 832.950 493.950 835.050 494.400 ;
        RECT 847.950 493.950 850.050 494.400 ;
        RECT 853.950 495.450 856.050 496.050 ;
        RECT 862.800 495.450 864.900 496.050 ;
        RECT 853.950 494.400 864.900 495.450 ;
        RECT 853.950 493.950 856.050 494.400 ;
        RECT 862.800 493.950 864.900 494.400 ;
        RECT 866.100 495.450 870.000 496.050 ;
        RECT 871.950 495.450 874.050 496.050 ;
        RECT 866.100 494.400 874.050 495.450 ;
        RECT 866.100 493.950 870.000 494.400 ;
        RECT 871.950 493.950 874.050 494.400 ;
        RECT 877.950 493.950 880.050 496.050 ;
        RECT 883.950 495.450 886.050 496.050 ;
        RECT 895.950 495.450 898.050 496.050 ;
        RECT 883.950 494.400 898.050 495.450 ;
        RECT 883.950 493.950 886.050 494.400 ;
        RECT 895.950 493.950 898.050 494.400 ;
        RECT 316.950 491.250 319.050 493.050 ;
        RECT 334.950 492.750 336.750 493.050 ;
        RECT 334.950 491.250 337.050 492.750 ;
        RECT 337.950 491.250 340.050 492.750 ;
        RECT 343.950 491.250 346.050 493.050 ;
        RECT 338.250 490.950 340.050 491.250 ;
        RECT 358.950 490.950 361.050 492.750 ;
        RECT 364.950 490.950 367.050 492.750 ;
        RECT 385.950 491.250 388.050 493.050 ;
        RECT 403.950 490.950 406.050 492.750 ;
        RECT 409.950 490.950 412.050 492.750 ;
        RECT 427.950 490.950 430.050 492.750 ;
        RECT 433.950 490.950 436.050 492.750 ;
        RECT 454.950 490.950 457.050 492.750 ;
        RECT 469.950 490.950 472.050 492.750 ;
        RECT 475.950 490.950 478.050 492.750 ;
        RECT 493.950 490.950 496.050 492.750 ;
        RECT 499.950 490.950 502.050 492.750 ;
        RECT 517.950 490.950 520.050 492.750 ;
        RECT 523.950 490.950 526.050 492.750 ;
        RECT 538.950 490.950 541.050 492.750 ;
        RECT 556.950 490.950 559.050 492.750 ;
        RECT 562.950 490.950 565.050 492.750 ;
        RECT 586.950 490.950 589.050 492.750 ;
        RECT 601.950 490.950 604.050 492.750 ;
        RECT 607.950 490.950 610.050 492.750 ;
        RECT 628.950 490.950 631.050 492.750 ;
        RECT 649.950 491.250 652.050 493.050 ;
        RECT 670.950 490.950 673.050 492.750 ;
        RECT 685.950 490.950 688.050 492.750 ;
        RECT 691.950 490.950 694.050 492.750 ;
        RECT 712.950 490.950 715.050 492.750 ;
        RECT 718.950 490.950 721.050 492.750 ;
        RECT 736.950 491.250 739.050 493.050 ;
        RECT 757.950 490.950 760.050 492.750 ;
        RECT 763.950 490.950 766.050 492.750 ;
        RECT 784.950 490.950 787.050 492.750 ;
        RECT 799.950 491.250 802.050 493.050 ;
        RECT 809.250 492.750 811.050 493.050 ;
        RECT 805.950 491.250 808.050 492.750 ;
        RECT 808.950 491.250 811.050 492.750 ;
        RECT 805.950 490.950 807.750 491.250 ;
        RECT 826.950 490.950 829.050 492.750 ;
        RECT 832.950 490.950 835.050 492.750 ;
        RECT 853.950 490.950 856.050 492.750 ;
        RECT 871.950 490.950 874.050 492.750 ;
        RECT 877.950 490.950 880.050 492.750 ;
        RECT 895.950 490.950 898.050 492.750 ;
        RECT 316.950 487.950 319.050 490.050 ;
        RECT 322.950 489.450 325.050 490.050 ;
        RECT 334.950 489.450 337.050 490.050 ;
        RECT 322.950 488.400 337.050 489.450 ;
        RECT 322.950 487.950 325.050 488.400 ;
        RECT 334.950 487.950 337.050 488.400 ;
        RECT 343.950 487.950 346.050 490.050 ;
        RECT 355.950 488.250 358.050 490.050 ;
        RECT 361.950 488.250 364.050 490.050 ;
        RECT 385.950 489.450 388.050 490.050 ;
        RECT 390.000 489.450 394.050 490.050 ;
        RECT 385.950 488.400 394.050 489.450 ;
        RECT 385.950 487.950 388.050 488.400 ;
        RECT 390.000 487.950 394.050 488.400 ;
        RECT 406.950 488.250 409.050 490.050 ;
        RECT 412.950 488.250 415.050 490.050 ;
        RECT 424.950 488.250 427.050 490.050 ;
        RECT 430.950 488.250 433.050 490.050 ;
        RECT 451.950 488.250 454.050 490.050 ;
        RECT 466.950 488.250 469.050 490.050 ;
        RECT 472.950 488.250 475.050 490.050 ;
        RECT 496.950 488.250 499.050 490.050 ;
        RECT 502.950 488.250 505.050 490.050 ;
        RECT 520.950 488.250 523.050 490.050 ;
        RECT 526.950 488.250 529.050 490.050 ;
        RECT 541.950 488.250 544.050 490.050 ;
        RECT 559.950 488.250 562.050 490.050 ;
        RECT 565.950 488.250 568.050 490.050 ;
        RECT 583.950 488.250 586.050 490.050 ;
        RECT 598.950 488.250 601.050 490.050 ;
        RECT 604.950 488.250 607.050 490.050 ;
        RECT 625.950 488.250 628.050 490.050 ;
        RECT 631.950 488.250 634.050 490.050 ;
        RECT 640.950 489.450 643.050 490.050 ;
        RECT 649.950 489.450 652.050 490.050 ;
        RECT 640.950 488.400 652.050 489.450 ;
        RECT 640.950 487.950 643.050 488.400 ;
        RECT 649.950 487.950 652.050 488.400 ;
        RECT 667.950 488.250 670.050 490.050 ;
        RECT 673.950 488.250 676.050 490.050 ;
        RECT 688.950 488.250 691.050 490.050 ;
        RECT 694.950 488.250 697.050 490.050 ;
        RECT 715.950 488.250 718.050 490.050 ;
        RECT 721.950 488.250 724.050 490.050 ;
        RECT 727.950 489.450 730.050 490.050 ;
        RECT 736.950 489.450 739.050 490.050 ;
        RECT 727.950 488.400 739.050 489.450 ;
        RECT 727.950 487.950 730.050 488.400 ;
        RECT 736.950 487.950 739.050 488.400 ;
        RECT 760.950 488.250 763.050 490.050 ;
        RECT 766.950 488.250 769.050 490.050 ;
        RECT 781.950 488.250 784.050 490.050 ;
        RECT 787.950 488.250 790.050 490.050 ;
        RECT 799.950 487.950 802.050 490.050 ;
        RECT 808.950 489.450 811.050 490.050 ;
        RECT 823.950 489.450 826.050 490.050 ;
        RECT 808.950 488.400 826.050 489.450 ;
        RECT 808.950 487.950 811.050 488.400 ;
        RECT 823.950 487.950 826.050 488.400 ;
        RECT 829.950 488.250 832.050 490.050 ;
        RECT 835.950 488.250 838.050 490.050 ;
        RECT 850.950 488.250 853.050 490.050 ;
        RECT 856.950 488.250 859.050 490.050 ;
        RECT 874.950 488.250 877.050 490.050 ;
        RECT 880.950 488.250 883.050 490.050 ;
        RECT 892.950 488.250 895.050 490.050 ;
        RECT 898.950 488.250 901.050 490.050 ;
        RECT 355.950 484.950 358.050 487.050 ;
        RECT 361.950 484.950 364.050 487.050 ;
        RECT 406.950 484.950 409.050 487.050 ;
        RECT 412.950 484.950 415.050 487.050 ;
        RECT 424.950 484.950 427.050 487.050 ;
        RECT 430.950 484.950 433.050 487.050 ;
        RECT 451.950 486.450 454.050 487.050 ;
        RECT 456.000 486.450 460.050 487.050 ;
        RECT 451.950 485.400 460.050 486.450 ;
        RECT 451.950 484.950 454.050 485.400 ;
        RECT 456.000 484.950 460.050 485.400 ;
        RECT 466.950 484.950 469.050 487.050 ;
        RECT 472.950 484.950 475.050 487.050 ;
        RECT 496.950 484.950 499.050 487.050 ;
        RECT 502.950 484.950 505.050 487.050 ;
        RECT 508.950 486.450 511.050 487.050 ;
        RECT 514.950 486.450 517.050 487.050 ;
        RECT 508.950 485.400 517.050 486.450 ;
        RECT 508.950 484.950 511.050 485.400 ;
        RECT 514.950 484.950 517.050 485.400 ;
        RECT 520.950 484.950 523.050 487.050 ;
        RECT 526.950 484.950 529.050 487.050 ;
        RECT 532.950 486.450 535.050 487.050 ;
        RECT 541.950 486.450 544.050 487.050 ;
        RECT 553.950 486.450 556.050 487.050 ;
        RECT 532.950 485.400 556.050 486.450 ;
        RECT 532.950 484.950 535.050 485.400 ;
        RECT 541.950 484.950 544.050 485.400 ;
        RECT 553.950 484.950 556.050 485.400 ;
        RECT 559.950 484.950 562.050 487.050 ;
        RECT 565.950 484.950 568.050 487.050 ;
        RECT 571.950 486.450 574.050 487.050 ;
        RECT 583.950 486.450 586.050 487.050 ;
        RECT 571.950 485.400 586.050 486.450 ;
        RECT 571.950 484.950 574.050 485.400 ;
        RECT 583.950 484.950 586.050 485.400 ;
        RECT 598.950 484.950 601.050 487.050 ;
        RECT 604.950 484.950 607.050 487.050 ;
        RECT 625.950 484.950 628.050 487.050 ;
        RECT 631.950 484.950 634.050 487.050 ;
        RECT 667.950 484.950 670.050 487.050 ;
        RECT 673.950 484.950 676.050 487.050 ;
        RECT 688.950 484.950 691.050 487.050 ;
        RECT 694.950 484.950 697.050 487.050 ;
        RECT 715.950 484.950 718.050 487.050 ;
        RECT 721.950 484.950 724.050 487.050 ;
        RECT 760.950 484.950 763.050 487.050 ;
        RECT 766.950 484.950 769.050 487.050 ;
        RECT 781.950 484.950 784.050 487.050 ;
        RECT 787.950 484.950 790.050 487.050 ;
        RECT 829.950 484.950 832.050 487.050 ;
        RECT 835.950 484.950 838.050 487.050 ;
        RECT 850.950 484.950 853.050 487.050 ;
        RECT 856.950 484.950 859.050 487.050 ;
        RECT 874.950 484.950 877.050 487.050 ;
        RECT 880.950 484.950 883.050 487.050 ;
        RECT 892.950 484.950 895.050 487.050 ;
        RECT 898.950 484.950 901.050 487.050 ;
        RECT 733.950 483.450 736.050 484.050 ;
        RECT 745.950 483.450 748.050 484.050 ;
        RECT 733.950 482.400 748.050 483.450 ;
        RECT 733.950 481.950 736.050 482.400 ;
        RECT 745.950 481.950 748.050 482.400 ;
        RECT 280.950 478.950 283.050 479.400 ;
        RECT 286.950 478.950 289.050 479.400 ;
        RECT 292.950 477.600 295.050 479.700 ;
        RECT 313.950 478.500 316.050 480.600 ;
        RECT 343.950 480.450 346.050 481.050 ;
        RECT 361.950 480.450 364.050 481.050 ;
        RECT 343.950 479.400 364.050 480.450 ;
        RECT 343.950 478.950 346.050 479.400 ;
        RECT 361.950 478.950 364.050 479.400 ;
        RECT 406.950 480.450 409.050 481.050 ;
        RECT 418.950 480.450 421.050 481.050 ;
        RECT 424.950 480.450 427.050 481.050 ;
        RECT 406.950 479.400 427.050 480.450 ;
        RECT 406.950 478.950 409.050 479.400 ;
        RECT 418.950 478.950 421.050 479.400 ;
        RECT 424.950 478.950 427.050 479.400 ;
        RECT 430.950 480.450 433.050 481.050 ;
        RECT 454.950 480.450 457.050 481.050 ;
        RECT 430.950 479.400 457.050 480.450 ;
        RECT 430.950 478.950 433.050 479.400 ;
        RECT 454.950 478.950 457.050 479.400 ;
        RECT 460.950 480.450 463.050 481.050 ;
        RECT 466.950 480.450 469.050 481.050 ;
        RECT 460.950 479.400 469.050 480.450 ;
        RECT 460.950 478.950 463.050 479.400 ;
        RECT 466.950 478.950 469.050 479.400 ;
        RECT 484.950 480.450 487.050 481.050 ;
        RECT 520.950 480.450 523.050 481.050 ;
        RECT 484.950 479.400 523.050 480.450 ;
        RECT 484.950 478.950 487.050 479.400 ;
        RECT 520.950 478.950 523.050 479.400 ;
        RECT 544.950 480.450 547.050 481.050 ;
        RECT 559.950 480.450 562.050 481.050 ;
        RECT 544.950 479.400 562.050 480.450 ;
        RECT 544.950 478.950 547.050 479.400 ;
        RECT 559.950 478.950 562.050 479.400 ;
        RECT 616.950 480.450 619.050 481.050 ;
        RECT 631.950 480.450 634.050 481.050 ;
        RECT 655.950 480.450 658.050 481.050 ;
        RECT 682.950 480.450 685.050 481.050 ;
        RECT 616.950 479.400 685.050 480.450 ;
        RECT 616.950 478.950 619.050 479.400 ;
        RECT 631.950 478.950 634.050 479.400 ;
        RECT 655.950 478.950 658.050 479.400 ;
        RECT 682.950 478.950 685.050 479.400 ;
        RECT 694.950 480.450 697.050 481.050 ;
        RECT 703.950 480.450 706.050 481.050 ;
        RECT 694.950 479.400 706.050 480.450 ;
        RECT 694.950 478.950 697.050 479.400 ;
        RECT 703.950 478.950 706.050 479.400 ;
        RECT 715.950 480.450 718.050 481.050 ;
        RECT 760.950 480.450 763.050 481.050 ;
        RECT 715.950 479.400 763.050 480.450 ;
        RECT 715.950 478.950 718.050 479.400 ;
        RECT 760.950 478.950 763.050 479.400 ;
        RECT 811.950 480.450 814.050 481.050 ;
        RECT 835.950 480.450 838.050 481.050 ;
        RECT 856.950 480.450 859.050 481.050 ;
        RECT 811.950 479.400 859.050 480.450 ;
        RECT 811.950 478.950 814.050 479.400 ;
        RECT 835.950 478.950 838.050 479.400 ;
        RECT 856.950 478.950 859.050 479.400 ;
        RECT 862.950 480.450 865.050 481.050 ;
        RECT 874.950 480.450 877.050 481.050 ;
        RECT 862.950 479.400 877.050 480.450 ;
        RECT 862.950 478.950 865.050 479.400 ;
        RECT 874.950 478.950 877.050 479.400 ;
        RECT 94.950 476.400 145.050 477.450 ;
        RECT 94.950 475.950 97.050 476.400 ;
        RECT 142.950 475.950 145.050 476.400 ;
        RECT 337.950 477.450 340.050 478.050 ;
        RECT 355.950 477.450 358.050 478.050 ;
        RECT 403.950 477.450 406.050 478.050 ;
        RECT 337.950 476.400 406.050 477.450 ;
        RECT 337.950 475.950 340.050 476.400 ;
        RECT 355.950 475.950 358.050 476.400 ;
        RECT 403.950 475.950 406.050 476.400 ;
        RECT 412.950 477.450 415.050 478.050 ;
        RECT 431.400 477.450 432.450 478.950 ;
        RECT 412.950 476.400 432.450 477.450 ;
        RECT 457.950 477.450 460.050 478.050 ;
        RECT 472.800 477.450 474.900 478.050 ;
        RECT 457.950 476.400 474.900 477.450 ;
        RECT 412.950 475.950 415.050 476.400 ;
        RECT 457.950 475.950 460.050 476.400 ;
        RECT 472.800 475.950 474.900 476.400 ;
        RECT 476.100 477.450 478.200 478.050 ;
        RECT 487.950 477.450 490.050 478.050 ;
        RECT 476.100 476.400 490.050 477.450 ;
        RECT 476.100 475.950 478.200 476.400 ;
        RECT 487.950 475.950 490.050 476.400 ;
        RECT 688.950 477.450 691.050 478.050 ;
        RECT 733.950 477.450 736.050 478.050 ;
        RECT 688.950 476.400 736.050 477.450 ;
        RECT 688.950 475.950 691.050 476.400 ;
        RECT 733.950 475.950 736.050 476.400 ;
        RECT 829.950 477.450 832.050 478.050 ;
        RECT 841.950 477.450 844.050 478.050 ;
        RECT 829.950 476.400 844.050 477.450 ;
        RECT 829.950 475.950 832.050 476.400 ;
        RECT 841.950 475.950 844.050 476.400 ;
        RECT 49.950 472.950 55.050 475.050 ;
        RECT 106.950 474.450 109.050 475.050 ;
        RECT 208.950 474.450 211.050 475.050 ;
        RECT 280.950 474.450 283.050 475.050 ;
        RECT 106.950 473.400 283.050 474.450 ;
        RECT 106.950 472.950 109.050 473.400 ;
        RECT 208.950 472.950 211.050 473.400 ;
        RECT 280.950 472.950 283.050 473.400 ;
        RECT 286.950 474.450 289.050 475.050 ;
        RECT 310.950 474.450 313.050 475.050 ;
        RECT 286.950 473.400 313.050 474.450 ;
        RECT 286.950 472.950 289.050 473.400 ;
        RECT 310.950 472.950 313.050 473.400 ;
        RECT 409.950 474.450 412.050 475.050 ;
        RECT 427.950 474.450 430.050 475.050 ;
        RECT 409.950 473.400 430.050 474.450 ;
        RECT 409.950 472.950 412.050 473.400 ;
        RECT 427.950 472.950 430.050 473.400 ;
        RECT 673.950 474.450 676.050 475.050 ;
        RECT 694.950 474.450 697.050 475.050 ;
        RECT 673.950 473.400 697.050 474.450 ;
        RECT 673.950 472.950 676.050 473.400 ;
        RECT 694.950 472.950 697.050 473.400 ;
        RECT 820.950 474.450 823.050 475.050 ;
        RECT 835.950 474.450 838.050 475.050 ;
        RECT 820.950 473.400 838.050 474.450 ;
        RECT 820.950 472.950 823.050 473.400 ;
        RECT 835.950 472.950 838.050 473.400 ;
        RECT 4.950 471.450 7.050 472.050 ;
        RECT 22.950 471.450 25.050 472.050 ;
        RECT 34.950 471.450 37.050 472.050 ;
        RECT 100.950 471.450 103.050 472.050 ;
        RECT 4.950 470.400 103.050 471.450 ;
        RECT 4.950 469.950 7.050 470.400 ;
        RECT 22.950 469.950 25.050 470.400 ;
        RECT 34.950 469.950 37.050 470.400 ;
        RECT 100.950 469.950 103.050 470.400 ;
        RECT 289.950 471.450 292.050 472.050 ;
        RECT 322.950 471.450 325.050 472.050 ;
        RECT 370.950 471.450 373.050 472.050 ;
        RECT 289.950 470.400 373.050 471.450 ;
        RECT 289.950 469.950 292.050 470.400 ;
        RECT 322.950 469.950 325.050 470.400 ;
        RECT 370.950 469.950 373.050 470.400 ;
        RECT 403.950 471.450 406.050 472.050 ;
        RECT 421.950 471.450 424.050 472.050 ;
        RECT 463.950 471.450 466.050 472.050 ;
        RECT 403.950 470.400 466.050 471.450 ;
        RECT 403.950 469.950 406.050 470.400 ;
        RECT 421.950 469.950 424.050 470.400 ;
        RECT 463.950 469.950 466.050 470.400 ;
        RECT 625.950 471.450 628.050 472.050 ;
        RECT 652.950 471.450 655.050 472.050 ;
        RECT 625.950 470.400 655.050 471.450 ;
        RECT 625.950 469.950 628.050 470.400 ;
        RECT 652.950 469.950 655.050 470.400 ;
        RECT 781.950 471.450 784.050 472.050 ;
        RECT 808.950 471.450 811.050 472.050 ;
        RECT 781.950 470.400 811.050 471.450 ;
        RECT 781.950 469.950 784.050 470.400 ;
        RECT 808.950 469.950 811.050 470.400 ;
        RECT 184.950 468.450 187.050 469.050 ;
        RECT 361.950 468.450 364.050 469.050 ;
        RECT 184.950 467.400 364.050 468.450 ;
        RECT 371.400 468.450 372.450 469.950 ;
        RECT 442.950 468.450 445.050 469.050 ;
        RECT 371.400 467.400 445.050 468.450 ;
        RECT 184.950 466.950 187.050 467.400 ;
        RECT 361.950 466.950 364.050 467.400 ;
        RECT 442.950 466.950 445.050 467.400 ;
        RECT 634.950 468.450 637.050 469.050 ;
        RECT 640.950 468.450 643.050 469.200 ;
        RECT 634.950 467.400 643.050 468.450 ;
        RECT 634.950 466.950 637.050 467.400 ;
        RECT 640.950 467.100 643.050 467.400 ;
        RECT 814.950 468.450 817.050 469.050 ;
        RECT 826.950 468.450 829.050 469.050 ;
        RECT 814.950 467.400 829.050 468.450 ;
        RECT 814.950 466.950 817.050 467.400 ;
        RECT 826.950 466.950 829.050 467.400 ;
        RECT 160.950 465.450 163.050 466.050 ;
        RECT 193.950 465.450 196.050 466.050 ;
        RECT 160.950 464.400 196.050 465.450 ;
        RECT 160.950 463.950 163.050 464.400 ;
        RECT 193.950 463.950 196.050 464.400 ;
        RECT 232.950 465.450 235.050 466.050 ;
        RECT 271.950 465.450 274.050 466.050 ;
        RECT 232.950 464.400 274.050 465.450 ;
        RECT 232.950 463.950 235.050 464.400 ;
        RECT 271.950 463.950 274.050 464.400 ;
        RECT 280.950 465.450 283.050 466.050 ;
        RECT 349.950 465.450 352.050 466.050 ;
        RECT 436.950 465.450 439.050 466.050 ;
        RECT 280.950 464.400 439.050 465.450 ;
        RECT 280.950 463.950 283.050 464.400 ;
        RECT 349.950 463.950 352.050 464.400 ;
        RECT 436.950 463.950 439.050 464.400 ;
        RECT 469.950 465.450 472.050 466.050 ;
        RECT 481.950 465.450 484.050 466.050 ;
        RECT 469.950 464.400 484.050 465.450 ;
        RECT 469.950 463.950 472.050 464.400 ;
        RECT 481.950 463.950 484.050 464.400 ;
        RECT 592.950 465.450 595.050 466.050 ;
        RECT 640.950 465.450 643.050 465.900 ;
        RECT 703.950 465.450 706.050 466.050 ;
        RECT 592.950 464.400 706.050 465.450 ;
        RECT 592.950 463.950 595.050 464.400 ;
        RECT 640.950 463.800 643.050 464.400 ;
        RECT 703.950 463.950 706.050 464.400 ;
        RECT 787.950 465.450 790.050 466.050 ;
        RECT 802.950 465.450 805.050 466.050 ;
        RECT 787.950 464.400 805.050 465.450 ;
        RECT 787.950 463.950 790.050 464.400 ;
        RECT 802.950 463.950 805.050 464.400 ;
        RECT 808.950 465.450 811.050 466.050 ;
        RECT 817.950 465.450 820.050 466.050 ;
        RECT 808.950 464.400 820.050 465.450 ;
        RECT 808.950 463.950 811.050 464.400 ;
        RECT 817.950 463.950 820.050 464.400 ;
        RECT 823.950 465.450 826.050 466.050 ;
        RECT 847.950 465.450 850.050 466.050 ;
        RECT 874.950 465.450 877.050 466.050 ;
        RECT 823.950 464.400 877.050 465.450 ;
        RECT 823.950 463.950 826.050 464.400 ;
        RECT 847.950 463.950 850.050 464.400 ;
        RECT 874.950 463.950 877.050 464.400 ;
        RECT 151.950 462.450 154.050 463.050 ;
        RECT 172.950 462.450 175.050 463.050 ;
        RECT 151.950 461.400 175.050 462.450 ;
        RECT 151.950 460.950 154.050 461.400 ;
        RECT 172.950 460.950 175.050 461.400 ;
        RECT 205.950 462.450 208.050 463.050 ;
        RECT 214.950 462.450 217.050 463.050 ;
        RECT 205.950 461.400 217.050 462.450 ;
        RECT 205.950 460.950 208.050 461.400 ;
        RECT 214.950 460.950 217.050 461.400 ;
        RECT 241.950 462.450 244.050 463.050 ;
        RECT 259.950 462.450 262.050 463.050 ;
        RECT 319.950 462.450 322.050 463.050 ;
        RECT 241.950 461.400 322.050 462.450 ;
        RECT 241.950 460.950 244.050 461.400 ;
        RECT 259.950 460.950 262.050 461.400 ;
        RECT 319.950 460.950 322.050 461.400 ;
        RECT 358.950 462.450 361.050 463.050 ;
        RECT 364.950 462.450 367.050 463.050 ;
        RECT 358.950 461.400 367.050 462.450 ;
        RECT 358.950 460.950 361.050 461.400 ;
        RECT 364.950 460.950 367.050 461.400 ;
        RECT 376.950 462.450 379.050 463.050 ;
        RECT 385.950 462.450 388.050 463.050 ;
        RECT 376.950 461.400 388.050 462.450 ;
        RECT 376.950 460.950 379.050 461.400 ;
        RECT 385.950 460.950 388.050 461.400 ;
        RECT 391.950 462.450 394.050 463.050 ;
        RECT 418.950 462.450 421.050 463.050 ;
        RECT 430.950 462.450 433.050 463.050 ;
        RECT 391.950 461.400 433.050 462.450 ;
        RECT 391.950 460.950 394.050 461.400 ;
        RECT 418.950 460.950 421.050 461.400 ;
        RECT 430.950 460.950 433.050 461.400 ;
        RECT 457.950 462.450 460.050 463.050 ;
        RECT 523.950 462.450 526.050 463.050 ;
        RECT 457.950 461.400 526.050 462.450 ;
        RECT 457.950 460.950 460.050 461.400 ;
        RECT 523.950 460.950 526.050 461.400 ;
        RECT 550.950 462.450 553.050 463.050 ;
        RECT 571.950 462.450 574.050 463.050 ;
        RECT 622.950 462.450 625.050 463.050 ;
        RECT 550.950 461.400 625.050 462.450 ;
        RECT 550.950 460.950 553.050 461.400 ;
        RECT 571.950 460.950 574.050 461.400 ;
        RECT 622.950 460.950 625.050 461.400 ;
        RECT 664.950 462.450 667.050 463.050 ;
        RECT 694.950 462.450 697.050 463.050 ;
        RECT 727.950 462.450 730.050 463.050 ;
        RECT 664.950 461.400 730.050 462.450 ;
        RECT 664.950 460.950 667.050 461.400 ;
        RECT 694.950 460.950 697.050 461.400 ;
        RECT 727.950 460.950 730.050 461.400 ;
        RECT 751.950 462.450 754.050 463.050 ;
        RECT 820.950 462.450 823.050 463.050 ;
        RECT 751.950 461.400 823.050 462.450 ;
        RECT 751.950 460.950 754.050 461.400 ;
        RECT 820.950 460.950 823.050 461.400 ;
        RECT 844.950 462.450 847.050 463.050 ;
        RECT 859.950 462.450 862.050 463.050 ;
        RECT 844.950 461.400 862.050 462.450 ;
        RECT 844.950 460.950 847.050 461.400 ;
        RECT 859.950 460.950 862.050 461.400 ;
        RECT 16.950 459.450 19.050 460.050 ;
        RECT 31.950 459.450 34.050 460.050 ;
        RECT 118.950 459.450 121.050 460.050 ;
        RECT 400.950 459.450 403.050 460.050 ;
        RECT 412.950 459.450 415.050 460.050 ;
        RECT 16.950 458.400 27.450 459.450 ;
        RECT 16.950 457.950 19.050 458.400 ;
        RECT 26.400 456.450 27.450 458.400 ;
        RECT 31.950 458.400 415.050 459.450 ;
        RECT 31.950 457.950 34.050 458.400 ;
        RECT 118.950 457.950 121.050 458.400 ;
        RECT 400.950 457.950 403.050 458.400 ;
        RECT 412.950 457.950 415.050 458.400 ;
        RECT 439.950 459.450 442.050 460.050 ;
        RECT 469.950 459.450 472.050 460.050 ;
        RECT 439.950 458.400 472.050 459.450 ;
        RECT 439.950 457.950 442.050 458.400 ;
        RECT 469.950 457.950 472.050 458.400 ;
        RECT 475.950 459.450 478.050 460.050 ;
        RECT 508.950 459.450 511.050 460.050 ;
        RECT 475.950 458.400 511.050 459.450 ;
        RECT 475.950 457.950 478.050 458.400 ;
        RECT 508.950 457.950 511.050 458.400 ;
        RECT 577.950 459.450 580.050 460.050 ;
        RECT 589.950 459.450 592.050 460.050 ;
        RECT 733.950 459.450 736.050 460.050 ;
        RECT 745.950 459.450 748.050 460.050 ;
        RECT 853.950 459.450 856.050 460.050 ;
        RECT 865.950 459.450 868.050 460.050 ;
        RECT 577.950 458.400 868.050 459.450 ;
        RECT 577.950 457.950 580.050 458.400 ;
        RECT 589.950 457.950 592.050 458.400 ;
        RECT 733.950 457.950 736.050 458.400 ;
        RECT 745.950 457.950 748.050 458.400 ;
        RECT 853.950 457.950 856.050 458.400 ;
        RECT 865.950 457.950 868.050 458.400 ;
        RECT 889.950 459.450 892.050 460.050 ;
        RECT 901.950 459.450 904.050 460.050 ;
        RECT 889.950 458.400 904.050 459.450 ;
        RECT 889.950 457.950 892.050 458.400 ;
        RECT 901.950 457.950 904.050 458.400 ;
        RECT 31.950 456.450 34.050 457.050 ;
        RECT 26.400 455.400 34.050 456.450 ;
        RECT 31.950 454.950 34.050 455.400 ;
        RECT 271.950 456.450 274.050 457.050 ;
        RECT 778.950 456.450 783.000 457.050 ;
        RECT 271.950 455.400 297.450 456.450 ;
        RECT 271.950 454.950 274.050 455.400 ;
        RECT 296.400 454.050 297.450 455.400 ;
        RECT 778.950 454.950 783.450 456.450 ;
        RECT 16.950 451.950 19.050 454.050 ;
        RECT 22.950 451.950 25.050 454.050 ;
        RECT 37.950 451.950 40.050 454.050 ;
        RECT 43.950 451.950 46.050 454.050 ;
        RECT 61.950 451.950 64.050 454.050 ;
        RECT 67.950 451.950 70.050 454.050 ;
        RECT 82.950 451.950 85.050 454.050 ;
        RECT 88.950 451.950 91.050 454.050 ;
        RECT 103.950 451.950 106.050 454.050 ;
        RECT 109.950 451.950 112.050 454.050 ;
        RECT 148.950 453.450 151.050 454.050 ;
        RECT 160.950 453.450 163.050 454.050 ;
        RECT 148.950 452.400 163.050 453.450 ;
        RECT 148.950 451.950 151.050 452.400 ;
        RECT 160.950 451.950 163.050 452.400 ;
        RECT 166.950 451.950 169.050 454.050 ;
        RECT 172.950 451.950 175.050 454.050 ;
        RECT 193.950 451.950 196.050 454.050 ;
        RECT 199.950 451.950 202.050 454.050 ;
        RECT 214.950 451.950 217.050 454.050 ;
        RECT 220.950 451.950 223.050 454.050 ;
        RECT 259.950 451.950 262.050 454.050 ;
        RECT 265.950 451.950 268.050 454.050 ;
        RECT 295.950 453.450 298.050 454.050 ;
        RECT 301.950 453.450 304.050 454.050 ;
        RECT 295.950 452.400 304.050 453.450 ;
        RECT 295.950 451.950 298.050 452.400 ;
        RECT 301.950 451.950 304.050 452.400 ;
        RECT 307.950 451.950 310.050 454.050 ;
        RECT 313.950 453.450 316.050 454.050 ;
        RECT 322.950 453.450 325.050 454.050 ;
        RECT 313.950 452.400 325.050 453.450 ;
        RECT 313.950 451.950 316.050 452.400 ;
        RECT 322.950 451.950 325.050 452.400 ;
        RECT 328.950 451.950 331.050 454.050 ;
        RECT 334.950 451.950 337.050 454.050 ;
        RECT 352.950 451.950 355.050 454.050 ;
        RECT 358.950 451.950 361.050 454.050 ;
        RECT 364.950 453.450 367.050 454.050 ;
        RECT 376.950 453.450 379.050 454.050 ;
        RECT 388.950 453.450 391.050 454.050 ;
        RECT 364.950 452.400 391.050 453.450 ;
        RECT 364.950 451.950 367.050 452.400 ;
        RECT 376.950 451.950 379.050 452.400 ;
        RECT 388.950 451.950 391.050 452.400 ;
        RECT 394.950 451.950 397.050 454.050 ;
        RECT 400.950 451.950 403.050 454.050 ;
        RECT 418.950 451.950 421.050 454.050 ;
        RECT 424.950 451.950 427.050 454.050 ;
        RECT 436.950 451.950 439.050 454.050 ;
        RECT 442.950 451.950 445.050 454.050 ;
        RECT 463.950 451.950 466.050 454.050 ;
        RECT 469.950 451.950 472.050 454.050 ;
        RECT 481.950 451.950 484.050 454.050 ;
        RECT 487.950 453.450 490.050 454.050 ;
        RECT 496.950 453.450 499.050 454.050 ;
        RECT 487.950 452.400 499.050 453.450 ;
        RECT 487.950 451.950 490.050 452.400 ;
        RECT 496.950 451.950 499.050 452.400 ;
        RECT 502.950 451.950 505.050 454.050 ;
        RECT 508.950 451.950 511.050 454.050 ;
        RECT 523.950 451.950 526.050 454.050 ;
        RECT 529.950 451.950 532.050 454.050 ;
        RECT 550.950 451.950 553.050 454.050 ;
        RECT 556.950 451.950 559.050 454.050 ;
        RECT 571.950 451.950 574.050 454.050 ;
        RECT 577.950 451.950 580.050 454.050 ;
        RECT 595.950 451.950 598.050 454.050 ;
        RECT 601.950 451.950 604.050 454.050 ;
        RECT 607.950 453.450 610.050 454.050 ;
        RECT 619.950 453.450 622.050 454.050 ;
        RECT 607.950 452.400 622.050 453.450 ;
        RECT 607.950 451.950 610.050 452.400 ;
        RECT 619.950 451.950 622.050 452.400 ;
        RECT 640.950 451.950 643.050 454.050 ;
        RECT 646.950 451.950 649.050 454.050 ;
        RECT 658.950 451.950 661.050 454.050 ;
        RECT 664.950 451.950 667.050 454.050 ;
        RECT 706.950 451.950 712.050 454.050 ;
        RECT 727.950 451.950 730.050 454.050 ;
        RECT 733.950 451.950 736.050 454.050 ;
        RECT 745.950 451.950 748.050 454.050 ;
        RECT 751.950 451.950 754.050 454.050 ;
        RECT 769.950 451.950 772.050 454.050 ;
        RECT 775.950 451.950 778.050 454.050 ;
        RECT 782.400 453.450 783.450 454.950 ;
        RECT 793.950 453.450 796.050 454.050 ;
        RECT 798.000 453.450 802.050 454.050 ;
        RECT 782.400 452.400 802.050 453.450 ;
        RECT 793.950 451.950 796.050 452.400 ;
        RECT 798.000 451.950 802.050 452.400 ;
        RECT 814.950 451.950 817.050 454.050 ;
        RECT 820.950 451.950 823.050 454.050 ;
        RECT 826.950 453.450 829.050 454.050 ;
        RECT 835.950 453.450 838.050 454.050 ;
        RECT 826.950 452.400 838.050 453.450 ;
        RECT 826.950 451.950 829.050 452.400 ;
        RECT 835.950 451.950 838.050 452.400 ;
        RECT 850.950 451.950 853.050 454.050 ;
        RECT 856.950 453.450 859.050 454.050 ;
        RECT 865.950 453.450 868.050 454.050 ;
        RECT 856.950 452.400 868.050 453.450 ;
        RECT 856.950 451.950 859.050 452.400 ;
        RECT 865.950 451.950 868.050 452.400 ;
        RECT 871.950 451.950 874.050 454.050 ;
        RECT 895.950 451.950 898.050 454.050 ;
        RECT 901.950 451.950 904.050 454.050 ;
        RECT 16.950 448.950 19.050 450.750 ;
        RECT 22.950 448.950 25.050 450.750 ;
        RECT 37.950 448.950 40.050 450.750 ;
        RECT 43.950 448.950 46.050 450.750 ;
        RECT 61.950 448.950 64.050 450.750 ;
        RECT 67.950 448.950 70.050 450.750 ;
        RECT 82.950 448.950 85.050 450.750 ;
        RECT 88.950 448.950 91.050 450.750 ;
        RECT 103.950 448.950 106.050 450.750 ;
        RECT 109.950 448.950 112.050 450.750 ;
        RECT 130.950 448.950 133.050 451.050 ;
        RECT 148.950 448.950 151.050 450.750 ;
        RECT 166.950 448.950 169.050 450.750 ;
        RECT 172.950 448.950 175.050 450.750 ;
        RECT 193.950 448.950 196.050 450.750 ;
        RECT 199.950 448.950 202.050 450.750 ;
        RECT 214.950 448.950 217.050 450.750 ;
        RECT 220.950 448.950 223.050 450.750 ;
        RECT 226.950 450.450 229.050 451.050 ;
        RECT 238.950 450.450 241.050 451.050 ;
        RECT 226.950 449.400 241.050 450.450 ;
        RECT 226.950 448.950 229.050 449.400 ;
        RECT 238.950 448.950 241.050 449.400 ;
        RECT 259.950 448.950 262.050 450.750 ;
        RECT 265.950 448.950 268.050 450.750 ;
        RECT 271.950 450.450 274.050 451.050 ;
        RECT 286.950 450.450 289.050 451.050 ;
        RECT 271.950 449.400 289.050 450.450 ;
        RECT 271.950 448.950 274.050 449.400 ;
        RECT 286.950 448.950 289.050 449.400 ;
        RECT 307.950 448.950 310.050 450.750 ;
        RECT 313.950 448.950 316.050 450.750 ;
        RECT 328.950 448.950 331.050 450.750 ;
        RECT 334.950 448.950 337.050 450.750 ;
        RECT 352.950 448.950 355.050 450.750 ;
        RECT 358.950 448.950 361.050 450.750 ;
        RECT 376.950 448.950 379.050 450.750 ;
        RECT 394.950 448.950 397.050 450.750 ;
        RECT 400.950 448.950 403.050 450.750 ;
        RECT 418.950 448.950 421.050 450.750 ;
        RECT 424.950 448.950 427.050 450.750 ;
        RECT 436.950 448.950 439.050 450.750 ;
        RECT 442.950 448.950 445.050 450.750 ;
        RECT 463.950 448.950 466.050 450.750 ;
        RECT 469.950 448.950 472.050 450.750 ;
        RECT 481.950 448.950 484.050 450.750 ;
        RECT 487.950 448.950 490.050 450.750 ;
        RECT 502.950 448.950 505.050 450.750 ;
        RECT 508.950 448.950 511.050 450.750 ;
        RECT 523.950 448.950 526.050 450.750 ;
        RECT 529.950 448.950 532.050 450.750 ;
        RECT 550.950 448.950 553.050 450.750 ;
        RECT 556.950 448.950 559.050 450.750 ;
        RECT 571.950 448.950 574.050 450.750 ;
        RECT 577.950 448.950 580.050 450.750 ;
        RECT 595.950 448.950 598.050 450.750 ;
        RECT 601.950 448.950 604.050 450.750 ;
        RECT 619.950 448.950 622.050 450.750 ;
        RECT 640.950 448.950 643.050 450.750 ;
        RECT 646.950 448.950 649.050 450.750 ;
        RECT 658.950 448.950 661.050 450.750 ;
        RECT 664.950 448.950 667.050 450.750 ;
        RECT 685.950 448.950 688.050 451.050 ;
        RECT 706.950 448.950 709.050 450.750 ;
        RECT 727.950 448.950 730.050 450.750 ;
        RECT 733.950 448.950 736.050 450.750 ;
        RECT 745.950 448.950 748.050 450.750 ;
        RECT 751.950 448.950 754.050 450.750 ;
        RECT 769.950 448.950 772.050 450.750 ;
        RECT 775.950 448.950 778.050 450.750 ;
        RECT 781.950 450.450 784.050 451.050 ;
        RECT 787.950 450.450 790.050 451.050 ;
        RECT 781.950 449.400 790.050 450.450 ;
        RECT 781.950 448.950 784.050 449.400 ;
        RECT 787.950 448.950 790.050 449.400 ;
        RECT 793.950 448.950 796.050 450.750 ;
        RECT 799.950 450.450 802.050 451.050 ;
        RECT 808.950 450.450 811.050 451.050 ;
        RECT 799.950 449.400 811.050 450.450 ;
        RECT 799.950 448.950 802.050 449.400 ;
        RECT 808.950 448.950 811.050 449.400 ;
        RECT 814.950 448.950 817.050 450.750 ;
        RECT 820.950 448.950 823.050 450.750 ;
        RECT 835.950 448.950 838.050 450.750 ;
        RECT 850.950 448.950 853.050 450.750 ;
        RECT 856.950 448.950 859.050 450.750 ;
        RECT 871.950 448.950 874.050 450.750 ;
        RECT 880.950 450.450 883.050 451.050 ;
        RECT 889.950 450.450 892.050 451.050 ;
        RECT 880.950 449.400 892.050 450.450 ;
        RECT 880.950 448.950 883.050 449.400 ;
        RECT 889.950 448.950 892.050 449.400 ;
        RECT 895.950 448.950 898.050 450.750 ;
        RECT 901.950 448.950 904.050 450.750 ;
        RECT 13.950 446.250 16.050 448.050 ;
        RECT 19.950 446.250 22.050 448.050 ;
        RECT 25.950 446.250 28.050 448.050 ;
        RECT 40.950 446.250 43.050 448.050 ;
        RECT 64.950 446.250 67.050 448.050 ;
        RECT 85.950 446.250 88.050 448.050 ;
        RECT 106.950 446.250 109.050 448.050 ;
        RECT 112.950 446.250 115.050 448.050 ;
        RECT 130.950 445.950 133.050 447.750 ;
        RECT 145.950 446.250 148.050 448.050 ;
        RECT 163.950 446.250 166.050 448.050 ;
        RECT 169.950 446.250 172.050 448.050 ;
        RECT 190.950 446.250 193.050 448.050 ;
        RECT 196.950 446.250 199.050 448.050 ;
        RECT 217.950 446.250 220.050 448.050 ;
        RECT 223.950 446.250 226.050 448.050 ;
        RECT 238.950 445.950 241.050 447.750 ;
        RECT 244.950 446.250 247.050 448.050 ;
        RECT 256.950 446.250 259.050 448.050 ;
        RECT 262.950 446.250 265.050 448.050 ;
        RECT 268.950 446.250 271.050 448.050 ;
        RECT 286.950 445.950 289.050 447.750 ;
        RECT 310.950 446.250 313.050 448.050 ;
        RECT 325.950 446.250 328.050 448.050 ;
        RECT 331.950 446.250 334.050 448.050 ;
        RECT 355.950 446.250 358.050 448.050 ;
        RECT 361.950 446.250 364.050 448.050 ;
        RECT 373.950 446.250 376.050 448.050 ;
        RECT 391.950 446.250 394.050 448.050 ;
        RECT 397.950 446.250 400.050 448.050 ;
        RECT 415.950 446.250 418.050 448.050 ;
        RECT 421.950 446.250 424.050 448.050 ;
        RECT 439.950 446.250 442.050 448.050 ;
        RECT 445.950 446.250 448.050 448.050 ;
        RECT 466.950 446.250 469.050 448.050 ;
        RECT 484.950 446.250 487.050 448.050 ;
        RECT 505.950 446.250 508.050 448.050 ;
        RECT 526.950 446.250 529.050 448.050 ;
        RECT 532.950 446.250 535.050 448.050 ;
        RECT 553.950 446.250 556.050 448.050 ;
        RECT 568.950 446.250 571.050 448.050 ;
        RECT 574.950 446.250 577.050 448.050 ;
        RECT 592.950 446.250 595.050 448.050 ;
        RECT 598.950 446.250 601.050 448.050 ;
        RECT 616.950 446.250 619.050 448.050 ;
        RECT 637.950 446.250 640.050 448.050 ;
        RECT 643.950 446.250 646.050 448.050 ;
        RECT 661.950 446.250 664.050 448.050 ;
        RECT 667.950 446.250 670.050 448.050 ;
        RECT 685.950 445.950 688.050 447.750 ;
        RECT 691.950 446.250 694.050 448.050 ;
        RECT 703.950 446.250 706.050 448.050 ;
        RECT 724.950 446.250 727.050 448.050 ;
        RECT 730.950 446.250 733.050 448.050 ;
        RECT 748.950 446.250 751.050 448.050 ;
        RECT 772.950 446.250 775.050 448.050 ;
        RECT 778.950 446.250 781.050 448.050 ;
        RECT 790.950 446.250 793.050 448.050 ;
        RECT 811.950 446.250 814.050 448.050 ;
        RECT 817.950 446.250 820.050 448.050 ;
        RECT 832.950 446.250 835.050 448.050 ;
        RECT 853.950 446.250 856.050 448.050 ;
        RECT 874.950 446.250 877.050 448.050 ;
        RECT 880.950 445.950 883.050 447.750 ;
        RECT 898.950 446.250 901.050 448.050 ;
        RECT 13.950 442.950 16.050 445.050 ;
        RECT 19.950 442.950 22.050 445.050 ;
        RECT 25.950 442.950 28.050 445.050 ;
        RECT 31.950 444.450 34.050 445.050 ;
        RECT 40.950 444.450 43.050 445.050 ;
        RECT 31.950 443.400 43.050 444.450 ;
        RECT 31.950 442.950 34.050 443.400 ;
        RECT 40.950 442.950 43.050 443.400 ;
        RECT 46.950 444.450 49.050 445.050 ;
        RECT 64.950 444.450 67.050 445.050 ;
        RECT 46.950 443.400 67.050 444.450 ;
        RECT 46.950 442.950 49.050 443.400 ;
        RECT 64.950 442.950 67.050 443.400 ;
        RECT 85.950 444.450 88.050 445.050 ;
        RECT 100.950 444.450 103.050 445.050 ;
        RECT 85.950 443.400 103.050 444.450 ;
        RECT 85.950 442.950 88.050 443.400 ;
        RECT 100.950 442.950 103.050 443.400 ;
        RECT 106.950 442.950 109.050 445.050 ;
        RECT 112.950 442.950 115.050 445.050 ;
        RECT 127.950 443.250 130.050 445.050 ;
        RECT 133.950 443.250 136.050 445.050 ;
        RECT 145.950 442.950 148.050 445.050 ;
        RECT 163.950 442.950 166.050 445.050 ;
        RECT 169.950 442.950 172.050 445.050 ;
        RECT 127.950 441.450 130.050 442.050 ;
        RECT 119.400 440.400 130.050 441.450 ;
        RECT 16.950 438.450 19.050 439.050 ;
        RECT 25.950 438.450 28.050 439.050 ;
        RECT 16.950 437.400 28.050 438.450 ;
        RECT 16.950 436.950 19.050 437.400 ;
        RECT 25.950 436.950 28.050 437.400 ;
        RECT 37.950 438.450 40.050 439.050 ;
        RECT 79.950 438.450 82.050 439.050 ;
        RECT 106.950 438.450 109.050 439.050 ;
        RECT 37.950 437.400 69.450 438.450 ;
        RECT 37.950 436.950 40.050 437.400 ;
        RECT 68.400 436.050 69.450 437.400 ;
        RECT 79.950 437.400 109.050 438.450 ;
        RECT 79.950 436.950 82.050 437.400 ;
        RECT 106.950 436.950 109.050 437.400 ;
        RECT 112.950 438.450 115.050 439.050 ;
        RECT 119.400 438.450 120.450 440.400 ;
        RECT 127.950 439.950 130.050 440.400 ;
        RECT 133.950 441.450 136.050 442.050 ;
        RECT 138.000 441.450 142.050 442.050 ;
        RECT 133.950 440.400 142.050 441.450 ;
        RECT 133.950 439.950 136.050 440.400 ;
        RECT 138.000 439.950 142.050 440.400 ;
        RECT 190.950 439.950 193.050 445.050 ;
        RECT 196.950 442.950 199.050 445.050 ;
        RECT 217.950 442.950 220.050 445.050 ;
        RECT 223.950 442.950 226.050 445.050 ;
        RECT 244.950 442.950 247.050 445.050 ;
        RECT 256.950 442.950 259.050 445.050 ;
        RECT 262.950 442.950 265.050 445.050 ;
        RECT 268.950 442.950 271.050 445.050 ;
        RECT 283.950 443.250 286.050 445.050 ;
        RECT 289.950 443.250 292.050 445.050 ;
        RECT 112.950 437.400 120.450 438.450 ;
        RECT 163.950 438.450 166.050 439.050 ;
        RECT 199.950 438.450 202.050 439.050 ;
        RECT 220.950 438.450 223.050 439.050 ;
        RECT 163.950 437.400 223.050 438.450 ;
        RECT 112.950 436.950 115.050 437.400 ;
        RECT 163.950 436.950 166.050 437.400 ;
        RECT 199.950 436.950 202.050 437.400 ;
        RECT 220.950 436.950 223.050 437.400 ;
        RECT 232.950 438.450 235.050 439.050 ;
        RECT 263.400 438.450 264.450 442.950 ;
        RECT 283.950 439.950 286.050 442.050 ;
        RECT 289.950 439.950 292.050 442.050 ;
        RECT 310.950 439.950 313.050 445.050 ;
        RECT 319.950 444.450 324.000 445.050 ;
        RECT 325.950 444.450 328.050 445.050 ;
        RECT 319.950 443.400 328.050 444.450 ;
        RECT 319.950 442.950 324.000 443.400 ;
        RECT 325.950 442.950 328.050 443.400 ;
        RECT 331.950 442.950 334.050 445.050 ;
        RECT 337.950 444.450 340.050 445.050 ;
        RECT 355.950 444.450 358.050 445.050 ;
        RECT 337.950 443.400 358.050 444.450 ;
        RECT 337.950 442.950 340.050 443.400 ;
        RECT 355.950 442.950 358.050 443.400 ;
        RECT 361.950 442.950 364.050 445.050 ;
        RECT 373.950 442.950 376.050 445.050 ;
        RECT 391.950 442.950 394.050 445.050 ;
        RECT 397.950 442.950 403.050 445.050 ;
        RECT 415.950 439.950 418.050 445.050 ;
        RECT 421.950 442.950 424.050 445.050 ;
        RECT 439.950 442.950 442.050 445.050 ;
        RECT 445.950 444.450 448.050 445.050 ;
        RECT 457.950 444.450 460.050 445.050 ;
        RECT 445.950 443.400 460.050 444.450 ;
        RECT 445.950 442.950 448.050 443.400 ;
        RECT 457.950 442.950 460.050 443.400 ;
        RECT 466.950 444.450 469.050 445.050 ;
        RECT 475.800 444.450 477.900 445.050 ;
        RECT 466.950 443.400 477.900 444.450 ;
        RECT 466.950 442.950 469.050 443.400 ;
        RECT 475.800 442.950 477.900 443.400 ;
        RECT 479.100 444.450 483.000 445.050 ;
        RECT 484.950 444.450 487.050 445.050 ;
        RECT 479.100 443.400 487.050 444.450 ;
        RECT 479.100 442.950 483.000 443.400 ;
        RECT 484.950 442.950 487.050 443.400 ;
        RECT 496.950 444.450 499.050 445.050 ;
        RECT 505.950 444.450 508.050 445.050 ;
        RECT 520.950 444.450 523.050 445.050 ;
        RECT 496.950 443.400 523.050 444.450 ;
        RECT 496.950 442.950 499.050 443.400 ;
        RECT 505.950 442.950 508.050 443.400 ;
        RECT 520.950 442.950 523.050 443.400 ;
        RECT 526.950 442.950 529.050 445.050 ;
        RECT 532.950 444.450 535.050 445.050 ;
        RECT 547.950 444.450 550.050 445.050 ;
        RECT 532.950 443.400 550.050 444.450 ;
        RECT 532.950 442.950 535.050 443.400 ;
        RECT 547.950 442.950 550.050 443.400 ;
        RECT 553.950 442.950 556.050 445.050 ;
        RECT 559.950 444.450 562.050 445.050 ;
        RECT 568.950 444.450 571.050 445.050 ;
        RECT 559.950 443.400 571.050 444.450 ;
        RECT 559.950 442.950 562.050 443.400 ;
        RECT 568.950 442.950 571.050 443.400 ;
        RECT 574.950 442.950 577.050 445.050 ;
        RECT 592.950 442.950 595.050 445.050 ;
        RECT 232.950 437.400 264.450 438.450 ;
        RECT 316.950 438.450 319.050 439.050 ;
        RECT 331.950 438.450 334.050 439.050 ;
        RECT 316.950 437.400 334.050 438.450 ;
        RECT 232.950 436.950 235.050 437.400 ;
        RECT 316.950 436.950 319.050 437.400 ;
        RECT 331.950 436.950 334.050 437.400 ;
        RECT 385.950 438.450 388.050 439.050 ;
        RECT 427.800 438.450 429.900 439.050 ;
        RECT 385.950 437.400 429.900 438.450 ;
        RECT 385.950 436.950 388.050 437.400 ;
        RECT 427.800 436.950 429.900 437.400 ;
        RECT 431.100 438.450 433.200 439.050 ;
        RECT 439.950 438.450 442.050 439.050 ;
        RECT 431.100 437.400 442.050 438.450 ;
        RECT 431.100 436.950 433.200 437.400 ;
        RECT 439.950 436.950 442.050 437.400 ;
        RECT 520.950 438.450 523.050 439.050 ;
        RECT 554.400 438.450 555.450 442.950 ;
        RECT 520.950 437.400 555.450 438.450 ;
        RECT 562.950 438.450 565.050 439.050 ;
        RECT 575.400 438.450 576.450 442.950 ;
        RECT 598.950 439.950 601.050 445.050 ;
        RECT 616.950 442.950 619.050 445.050 ;
        RECT 622.950 444.450 625.050 445.050 ;
        RECT 637.950 444.450 640.050 445.050 ;
        RECT 622.950 443.400 640.050 444.450 ;
        RECT 622.950 442.950 625.050 443.400 ;
        RECT 637.950 442.950 640.050 443.400 ;
        RECT 643.950 442.950 646.050 445.050 ;
        RECT 661.950 442.950 664.050 445.050 ;
        RECT 667.950 444.450 670.050 445.050 ;
        RECT 676.950 444.450 679.050 445.050 ;
        RECT 667.950 443.400 679.050 444.450 ;
        RECT 667.950 442.950 670.050 443.400 ;
        RECT 676.950 442.950 679.050 443.400 ;
        RECT 688.950 442.950 694.050 445.050 ;
        RECT 703.950 442.950 706.050 445.050 ;
        RECT 715.950 444.450 718.050 445.050 ;
        RECT 724.950 444.450 727.050 445.050 ;
        RECT 715.950 443.400 727.050 444.450 ;
        RECT 715.950 442.950 718.050 443.400 ;
        RECT 724.950 442.950 727.050 443.400 ;
        RECT 730.950 442.950 733.050 445.050 ;
        RECT 748.950 442.950 751.050 445.050 ;
        RECT 766.950 444.450 771.000 445.050 ;
        RECT 772.950 444.450 775.050 445.050 ;
        RECT 766.950 443.400 775.050 444.450 ;
        RECT 766.950 442.950 771.000 443.400 ;
        RECT 772.950 442.950 775.050 443.400 ;
        RECT 778.950 442.950 781.050 445.050 ;
        RECT 790.950 442.950 793.050 445.050 ;
        RECT 796.950 444.450 799.050 445.050 ;
        RECT 811.950 444.450 814.050 445.050 ;
        RECT 796.950 443.400 814.050 444.450 ;
        RECT 796.950 442.950 799.050 443.400 ;
        RECT 811.950 442.950 814.050 443.400 ;
        RECT 817.950 442.950 820.050 445.050 ;
        RECT 832.950 442.950 835.050 445.050 ;
        RECT 853.950 442.950 856.050 445.050 ;
        RECT 874.950 442.950 877.050 445.050 ;
        RECT 892.950 444.450 897.000 445.050 ;
        RECT 898.950 444.450 901.050 445.050 ;
        RECT 892.950 443.400 901.050 444.450 ;
        RECT 892.950 442.950 897.000 443.400 ;
        RECT 898.950 442.950 901.050 443.400 ;
        RECT 562.950 437.400 576.450 438.450 ;
        RECT 577.950 438.450 580.050 439.050 ;
        RECT 616.950 438.450 619.050 439.050 ;
        RECT 749.400 438.450 750.450 442.950 ;
        RECT 577.950 437.400 750.450 438.450 ;
        RECT 799.800 438.000 801.900 439.050 ;
        RECT 808.950 438.450 811.050 439.050 ;
        RECT 832.950 438.450 835.050 439.050 ;
        RECT 854.400 438.450 855.450 442.950 ;
        RECT 892.950 438.450 895.050 439.050 ;
        RECT 520.950 436.950 523.050 437.400 ;
        RECT 562.950 436.950 565.050 437.400 ;
        RECT 577.950 436.950 580.050 437.400 ;
        RECT 616.950 436.950 619.050 437.400 ;
        RECT 799.800 436.950 802.050 438.000 ;
        RECT 808.950 437.400 895.050 438.450 ;
        RECT 808.950 436.950 811.050 437.400 ;
        RECT 832.950 436.950 835.050 437.400 ;
        RECT 892.950 436.950 895.050 437.400 ;
        RECT 22.950 435.450 25.050 436.050 ;
        RECT 67.950 435.450 70.050 436.050 ;
        RECT 88.950 435.450 91.050 436.050 ;
        RECT 109.950 435.450 112.050 436.050 ;
        RECT 164.400 435.450 165.450 436.950 ;
        RECT 22.950 434.400 165.450 435.450 ;
        RECT 184.950 435.450 187.050 436.050 ;
        RECT 196.950 435.450 199.050 436.200 ;
        RECT 799.950 436.050 802.050 436.950 ;
        RECT 184.950 434.400 199.050 435.450 ;
        RECT 22.950 433.950 25.050 434.400 ;
        RECT 67.950 433.950 70.050 434.400 ;
        RECT 88.950 433.950 91.050 434.400 ;
        RECT 109.950 433.950 112.050 434.400 ;
        RECT 184.950 433.950 187.050 434.400 ;
        RECT 196.950 434.100 199.050 434.400 ;
        RECT 238.950 435.450 241.050 436.050 ;
        RECT 256.950 435.450 259.050 436.050 ;
        RECT 238.950 434.400 259.050 435.450 ;
        RECT 238.950 433.950 241.050 434.400 ;
        RECT 256.950 433.950 259.050 434.400 ;
        RECT 262.950 435.450 265.050 436.050 ;
        RECT 337.950 435.450 340.050 436.050 ;
        RECT 262.950 434.400 340.050 435.450 ;
        RECT 262.950 433.950 265.050 434.400 ;
        RECT 337.950 433.950 340.050 434.400 ;
        RECT 361.950 435.450 364.050 436.050 ;
        RECT 391.950 435.450 394.050 436.050 ;
        RECT 361.950 434.400 394.050 435.450 ;
        RECT 361.950 433.950 364.050 434.400 ;
        RECT 391.950 433.950 394.050 434.400 ;
        RECT 547.950 435.450 550.050 436.050 ;
        RECT 604.950 435.450 607.050 436.050 ;
        RECT 547.950 434.400 607.050 435.450 ;
        RECT 547.950 433.950 550.050 434.400 ;
        RECT 604.950 433.950 607.050 434.400 ;
        RECT 634.950 435.450 637.050 436.050 ;
        RECT 643.950 435.450 646.050 436.050 ;
        RECT 634.950 434.400 646.050 435.450 ;
        RECT 634.950 433.950 637.050 434.400 ;
        RECT 643.950 433.950 646.050 434.400 ;
        RECT 652.950 435.450 655.050 436.050 ;
        RECT 661.950 435.450 664.050 436.050 ;
        RECT 652.950 434.400 664.050 435.450 ;
        RECT 652.950 433.950 655.050 434.400 ;
        RECT 661.950 433.950 664.050 434.400 ;
        RECT 685.950 435.450 688.050 436.050 ;
        RECT 730.950 435.450 733.050 436.050 ;
        RECT 751.950 435.450 754.050 436.050 ;
        RECT 685.950 434.400 729.450 435.450 ;
        RECT 685.950 433.950 688.050 434.400 ;
        RECT 196.950 432.450 199.050 432.900 ;
        RECT 232.950 432.450 235.050 433.050 ;
        RECT 196.950 431.400 235.050 432.450 ;
        RECT 196.950 430.800 199.050 431.400 ;
        RECT 232.950 430.950 235.050 431.400 ;
        RECT 244.950 432.450 247.050 433.050 ;
        RECT 334.950 432.450 337.050 433.050 ;
        RECT 244.950 431.400 337.050 432.450 ;
        RECT 244.950 430.950 247.050 431.400 ;
        RECT 334.950 430.950 337.050 431.400 ;
        RECT 628.950 432.450 631.050 433.050 ;
        RECT 646.950 432.450 649.050 433.050 ;
        RECT 628.950 431.400 649.050 432.450 ;
        RECT 628.950 430.950 631.050 431.400 ;
        RECT 646.950 430.950 649.050 431.400 ;
        RECT 655.950 432.450 658.050 433.050 ;
        RECT 682.950 432.450 685.050 433.050 ;
        RECT 655.950 431.400 685.050 432.450 ;
        RECT 728.400 432.450 729.450 434.400 ;
        RECT 730.950 434.400 754.050 435.450 ;
        RECT 730.950 433.950 733.050 434.400 ;
        RECT 751.950 433.950 754.050 434.400 ;
        RECT 799.800 435.000 802.050 436.050 ;
        RECT 803.100 435.000 805.200 436.050 ;
        RECT 799.800 433.950 801.900 435.000 ;
        RECT 802.950 433.950 805.200 435.000 ;
        RECT 892.950 433.950 898.050 436.050 ;
        RECT 769.950 432.450 772.050 433.050 ;
        RECT 796.950 432.450 799.050 433.050 ;
        RECT 802.950 432.450 805.050 433.950 ;
        RECT 728.400 431.400 783.450 432.450 ;
        RECT 655.950 430.950 658.050 431.400 ;
        RECT 682.950 430.950 685.050 431.400 ;
        RECT 769.950 430.950 772.050 431.400 ;
        RECT 7.950 429.450 10.050 430.050 ;
        RECT 40.950 429.450 43.050 430.050 ;
        RECT 7.950 428.400 43.050 429.450 ;
        RECT 7.950 427.950 10.050 428.400 ;
        RECT 40.950 427.950 43.050 428.400 ;
        RECT 61.950 429.450 64.050 430.050 ;
        RECT 85.950 429.450 88.050 430.050 ;
        RECT 61.950 428.400 88.050 429.450 ;
        RECT 61.950 427.950 64.050 428.400 ;
        RECT 85.950 427.950 88.050 428.400 ;
        RECT 136.950 429.450 139.050 430.050 ;
        RECT 142.950 429.450 145.050 430.050 ;
        RECT 136.950 428.400 145.050 429.450 ;
        RECT 136.950 427.950 139.050 428.400 ;
        RECT 142.950 427.950 145.050 428.400 ;
        RECT 160.950 429.450 163.050 430.050 ;
        RECT 169.950 429.450 172.050 430.050 ;
        RECT 160.950 428.400 172.050 429.450 ;
        RECT 160.950 427.950 163.050 428.400 ;
        RECT 169.950 427.950 172.050 428.400 ;
        RECT 214.950 429.450 217.050 430.050 ;
        RECT 223.950 429.450 226.050 430.050 ;
        RECT 214.950 428.400 226.050 429.450 ;
        RECT 214.950 427.950 217.050 428.400 ;
        RECT 223.950 427.950 226.050 428.400 ;
        RECT 427.950 429.450 430.050 430.050 ;
        RECT 487.950 429.450 490.050 430.050 ;
        RECT 427.950 428.400 490.050 429.450 ;
        RECT 427.950 427.950 430.050 428.400 ;
        RECT 487.950 427.950 490.050 428.400 ;
        RECT 565.950 429.450 568.050 430.050 ;
        RECT 604.950 429.450 607.050 430.050 ;
        RECT 727.950 429.450 730.050 430.050 ;
        RECT 772.950 429.450 775.050 430.050 ;
        RECT 565.950 428.400 775.050 429.450 ;
        RECT 782.400 429.450 783.450 431.400 ;
        RECT 796.950 432.000 805.050 432.450 ;
        RECT 796.950 431.400 804.450 432.000 ;
        RECT 796.950 430.950 799.050 431.400 ;
        RECT 859.950 429.450 862.050 430.050 ;
        RECT 782.400 428.400 862.050 429.450 ;
        RECT 565.950 427.950 568.050 428.400 ;
        RECT 604.950 427.950 607.050 428.400 ;
        RECT 727.950 427.950 730.050 428.400 ;
        RECT 772.950 427.950 775.050 428.400 ;
        RECT 859.950 427.950 862.050 428.400 ;
        RECT 259.950 426.450 262.050 427.050 ;
        RECT 301.950 426.450 304.050 427.050 ;
        RECT 397.950 426.450 400.050 427.050 ;
        RECT 259.950 425.400 282.450 426.450 ;
        RECT 259.950 424.950 262.050 425.400 ;
        RECT 7.950 422.400 10.050 424.500 ;
        RECT 28.950 422.400 31.050 424.500 ;
        RECT 43.950 423.450 46.050 424.050 ;
        RECT 55.950 423.450 58.050 424.050 ;
        RECT 43.950 422.400 58.050 423.450 ;
        RECT 70.950 422.400 73.050 424.500 ;
        RECT 91.950 422.400 94.050 424.500 ;
        RECT 109.950 423.450 112.050 424.050 ;
        RECT 115.950 423.450 118.050 424.050 ;
        RECT 109.950 422.400 118.050 423.450 ;
        RECT 4.950 413.250 7.050 415.050 ;
        RECT 4.950 409.950 7.050 412.050 ;
        RECT 8.700 402.600 9.900 422.400 ;
        RECT 13.950 413.250 16.050 415.050 ;
        RECT 28.950 407.400 30.150 422.400 ;
        RECT 43.950 421.950 46.050 422.400 ;
        RECT 55.950 421.950 58.050 422.400 ;
        RECT 31.950 415.950 34.050 418.050 ;
        RECT 49.950 415.950 52.050 418.050 ;
        RECT 55.950 415.950 58.050 418.050 ;
        RECT 61.950 415.950 64.050 418.050 ;
        RECT 31.950 412.950 34.050 414.750 ;
        RECT 49.950 412.950 52.050 414.750 ;
        RECT 55.950 412.950 58.050 414.750 ;
        RECT 61.950 412.950 64.050 414.750 ;
        RECT 67.950 413.250 70.050 415.050 ;
        RECT 52.950 410.250 55.050 412.050 ;
        RECT 58.950 410.250 61.050 412.050 ;
        RECT 67.950 409.950 70.050 412.050 ;
        RECT 28.950 405.300 31.050 407.400 ;
        RECT 52.950 406.950 55.050 409.050 ;
        RECT 58.950 406.950 61.050 409.050 ;
        RECT 7.950 400.500 10.050 402.600 ;
        RECT 28.950 401.700 30.150 405.300 ;
        RECT 43.950 402.450 46.050 403.050 ;
        RECT 49.950 402.450 52.050 403.050 ;
        RECT 71.700 402.600 72.900 422.400 ;
        RECT 76.950 413.250 79.050 415.050 ;
        RECT 76.950 409.950 82.050 412.050 ;
        RECT 91.950 407.400 93.150 422.400 ;
        RECT 109.950 421.950 112.050 422.400 ;
        RECT 115.950 421.950 118.050 422.400 ;
        RECT 121.950 420.450 124.050 421.050 ;
        RECT 130.950 420.450 133.050 421.050 ;
        RECT 121.950 419.400 133.050 420.450 ;
        RECT 121.950 418.950 124.050 419.400 ;
        RECT 130.950 418.950 133.050 419.400 ;
        RECT 136.950 418.950 139.050 424.050 ;
        RECT 145.950 422.400 148.050 424.500 ;
        RECT 166.950 422.400 169.050 424.500 ;
        RECT 181.950 422.400 184.050 424.500 ;
        RECT 202.950 422.400 205.050 424.500 ;
        RECT 217.950 422.400 220.050 424.500 ;
        RECT 238.950 422.400 241.050 424.500 ;
        RECT 94.950 415.950 97.050 418.050 ;
        RECT 100.950 417.450 103.050 418.050 ;
        RECT 115.950 417.450 118.050 418.050 ;
        RECT 100.950 416.400 118.050 417.450 ;
        RECT 100.950 415.950 103.050 416.400 ;
        RECT 115.950 415.950 118.050 416.400 ;
        RECT 130.950 415.950 133.050 417.750 ;
        RECT 136.950 415.950 139.050 417.750 ;
        RECT 142.950 415.950 145.050 418.050 ;
        RECT 94.950 412.950 97.050 414.750 ;
        RECT 115.950 412.950 118.050 414.750 ;
        RECT 133.950 413.250 136.050 415.050 ;
        RECT 142.950 412.950 145.050 414.750 ;
        RECT 112.950 410.250 115.050 412.050 ;
        RECT 91.950 405.300 94.050 407.400 ;
        RECT 112.950 406.950 115.050 409.050 ;
        RECT 133.950 406.950 136.050 412.050 ;
        RECT 146.850 407.400 148.050 422.400 ;
        RECT 160.950 413.250 163.050 415.050 ;
        RECT 160.950 409.950 163.050 412.050 ;
        RECT 145.950 405.300 148.050 407.400 ;
        RECT 28.950 399.600 31.050 401.700 ;
        RECT 43.950 401.400 52.050 402.450 ;
        RECT 43.950 400.950 46.050 401.400 ;
        RECT 49.950 400.950 52.050 401.400 ;
        RECT 70.950 400.500 73.050 402.600 ;
        RECT 91.950 401.700 93.150 405.300 ;
        RECT 146.850 401.700 148.050 405.300 ;
        RECT 167.100 402.600 168.300 422.400 ;
        RECT 178.950 415.950 181.050 418.050 ;
        RECT 169.950 413.250 172.050 415.050 ;
        RECT 178.950 412.950 181.050 414.750 ;
        RECT 169.950 409.950 172.050 412.050 ;
        RECT 182.850 407.400 184.050 422.400 ;
        RECT 196.950 413.250 199.050 415.050 ;
        RECT 196.950 409.950 199.050 412.050 ;
        RECT 181.950 405.300 184.050 407.400 ;
        RECT 91.950 399.600 94.050 401.700 ;
        RECT 145.950 399.600 148.050 401.700 ;
        RECT 166.950 400.500 169.050 402.600 ;
        RECT 182.850 401.700 184.050 405.300 ;
        RECT 203.100 402.600 204.300 422.400 ;
        RECT 205.950 413.250 208.050 415.050 ;
        RECT 214.950 413.250 217.050 415.050 ;
        RECT 205.950 409.950 208.050 412.050 ;
        RECT 214.950 409.950 217.050 412.050 ;
        RECT 205.950 405.450 208.050 406.050 ;
        RECT 214.950 405.450 217.050 406.050 ;
        RECT 205.950 404.400 217.050 405.450 ;
        RECT 205.950 403.950 208.050 404.400 ;
        RECT 214.950 403.950 217.050 404.400 ;
        RECT 218.700 402.600 219.900 422.400 ;
        RECT 223.950 413.250 226.050 415.050 ;
        RECT 223.950 409.950 226.050 412.050 ;
        RECT 238.950 407.400 240.150 422.400 ;
        RECT 281.400 421.050 282.450 425.400 ;
        RECT 301.950 425.400 400.050 426.450 ;
        RECT 301.950 424.950 304.050 425.400 ;
        RECT 397.950 424.950 400.050 425.400 ;
        RECT 406.950 426.450 409.050 427.050 ;
        RECT 478.950 426.450 481.050 427.050 ;
        RECT 484.950 426.450 487.050 427.050 ;
        RECT 406.950 425.400 487.050 426.450 ;
        RECT 406.950 424.950 409.050 425.400 ;
        RECT 478.950 424.950 481.050 425.400 ;
        RECT 484.950 424.950 487.050 425.400 ;
        RECT 529.950 426.450 532.050 427.050 ;
        RECT 676.950 426.450 679.050 427.050 ;
        RECT 697.950 426.450 700.050 427.050 ;
        RECT 529.950 425.400 700.050 426.450 ;
        RECT 529.950 424.950 532.050 425.400 ;
        RECT 676.950 424.950 679.050 425.400 ;
        RECT 697.950 424.950 700.050 425.400 ;
        RECT 703.950 426.450 706.050 427.050 ;
        RECT 715.950 426.450 718.050 427.050 ;
        RECT 703.950 425.400 718.050 426.450 ;
        RECT 703.950 424.950 706.050 425.400 ;
        RECT 715.950 424.950 718.050 425.400 ;
        RECT 781.950 426.450 784.050 427.050 ;
        RECT 844.950 426.450 847.050 427.050 ;
        RECT 781.950 425.400 847.050 426.450 ;
        RECT 781.950 424.950 784.050 425.400 ;
        RECT 844.950 424.950 847.050 425.400 ;
        RECT 874.950 426.450 877.050 427.050 ;
        RECT 883.950 426.450 886.050 427.050 ;
        RECT 889.950 426.450 892.050 427.050 ;
        RECT 874.950 425.400 892.050 426.450 ;
        RECT 874.950 424.950 877.050 425.400 ;
        RECT 883.950 424.950 886.050 425.400 ;
        RECT 889.950 424.950 892.050 425.400 ;
        RECT 265.950 420.450 268.050 421.050 ;
        RECT 274.950 420.450 277.050 421.050 ;
        RECT 265.950 419.400 277.050 420.450 ;
        RECT 265.950 418.950 268.050 419.400 ;
        RECT 274.950 418.950 277.050 419.400 ;
        RECT 280.950 418.950 283.050 421.050 ;
        RECT 292.950 420.450 297.000 421.050 ;
        RECT 298.950 420.450 301.050 421.050 ;
        RECT 292.950 419.400 301.050 420.450 ;
        RECT 292.950 418.950 297.000 419.400 ;
        RECT 298.950 418.950 301.050 419.400 ;
        RECT 304.950 418.950 307.050 424.050 ;
        RECT 310.950 418.950 313.050 424.050 ;
        RECT 322.950 423.450 325.050 424.050 ;
        RECT 355.950 423.450 358.050 424.050 ;
        RECT 376.950 423.450 379.050 424.050 ;
        RECT 322.950 422.400 379.050 423.450 ;
        RECT 322.950 421.950 325.050 422.400 ;
        RECT 355.950 421.950 358.050 422.400 ;
        RECT 376.950 421.950 379.050 422.400 ;
        RECT 460.950 423.450 463.050 424.050 ;
        RECT 514.950 423.450 517.050 424.050 ;
        RECT 637.950 423.450 640.050 424.050 ;
        RECT 658.950 423.450 661.050 424.050 ;
        RECT 460.950 422.400 513.450 423.450 ;
        RECT 460.950 421.950 463.050 422.400 ;
        RECT 400.950 418.950 403.050 421.050 ;
        RECT 406.950 418.950 409.050 421.050 ;
        RECT 512.400 418.050 513.450 422.400 ;
        RECT 514.950 422.400 600.450 423.450 ;
        RECT 514.950 421.950 517.050 422.400 ;
        RECT 599.400 421.050 600.450 422.400 ;
        RECT 637.950 422.400 661.050 423.450 ;
        RECT 637.950 421.950 640.050 422.400 ;
        RECT 658.950 421.950 661.050 422.400 ;
        RECT 589.950 420.450 592.050 421.050 ;
        RECT 598.950 420.450 601.050 421.050 ;
        RECT 589.950 419.400 601.050 420.450 ;
        RECT 589.950 418.950 592.050 419.400 ;
        RECT 598.950 418.950 601.050 419.400 ;
        RECT 697.950 418.950 700.050 421.050 ;
        RECT 703.950 418.950 706.050 421.050 ;
        RECT 241.950 415.950 244.050 418.050 ;
        RECT 247.950 417.450 250.050 418.050 ;
        RECT 256.950 417.450 259.050 418.050 ;
        RECT 247.950 416.400 259.050 417.450 ;
        RECT 247.950 415.950 250.050 416.400 ;
        RECT 256.950 415.950 259.050 416.400 ;
        RECT 274.950 415.950 277.050 417.750 ;
        RECT 280.950 415.950 283.050 417.750 ;
        RECT 298.950 415.950 301.050 417.750 ;
        RECT 304.950 415.950 307.050 417.750 ;
        RECT 316.950 415.950 319.050 418.050 ;
        RECT 334.950 415.950 337.050 418.050 ;
        RECT 343.950 417.450 346.050 418.050 ;
        RECT 361.950 417.450 364.050 418.050 ;
        RECT 343.950 416.400 364.050 417.450 ;
        RECT 343.950 415.950 346.050 416.400 ;
        RECT 361.950 415.950 364.050 416.400 ;
        RECT 370.950 417.450 373.050 418.050 ;
        RECT 379.950 417.450 382.050 418.050 ;
        RECT 370.950 416.400 382.050 417.450 ;
        RECT 370.950 415.950 373.050 416.400 ;
        RECT 379.950 415.950 382.050 416.400 ;
        RECT 400.950 415.950 403.050 417.750 ;
        RECT 406.950 415.950 409.050 417.750 ;
        RECT 418.950 415.950 421.050 418.050 ;
        RECT 424.950 417.450 427.050 418.050 ;
        RECT 433.950 417.450 436.050 418.050 ;
        RECT 424.950 416.400 436.050 417.450 ;
        RECT 424.950 415.950 427.050 416.400 ;
        RECT 433.950 415.950 436.050 416.400 ;
        RECT 442.950 415.950 445.050 418.050 ;
        RECT 472.950 415.950 475.050 418.050 ;
        RECT 484.950 415.950 487.050 418.050 ;
        RECT 490.950 417.450 493.050 418.050 ;
        RECT 505.950 417.450 508.050 418.050 ;
        RECT 490.950 416.400 508.050 417.450 ;
        RECT 490.950 415.950 493.050 416.400 ;
        RECT 505.950 415.950 508.050 416.400 ;
        RECT 511.950 415.950 514.050 418.050 ;
        RECT 517.950 415.950 520.050 418.050 ;
        RECT 526.950 417.450 529.050 418.050 ;
        RECT 535.950 417.450 538.050 418.050 ;
        RECT 526.950 416.400 538.050 417.450 ;
        RECT 526.950 415.950 529.050 416.400 ;
        RECT 535.950 415.950 538.050 416.400 ;
        RECT 541.950 415.950 544.050 418.050 ;
        RECT 547.950 417.450 550.050 418.050 ;
        RECT 562.950 417.450 565.050 418.050 ;
        RECT 547.950 416.400 565.050 417.450 ;
        RECT 547.950 415.950 550.050 416.400 ;
        RECT 562.950 415.950 565.050 416.400 ;
        RECT 568.950 417.450 571.050 418.050 ;
        RECT 580.950 417.450 583.050 418.050 ;
        RECT 568.950 416.400 583.050 417.450 ;
        RECT 568.950 415.950 571.050 416.400 ;
        RECT 580.950 415.950 583.050 416.400 ;
        RECT 586.950 415.950 589.050 418.050 ;
        RECT 604.950 415.950 607.050 418.050 ;
        RECT 622.950 417.450 625.050 418.050 ;
        RECT 627.000 417.450 631.050 418.050 ;
        RECT 622.950 416.400 631.050 417.450 ;
        RECT 622.950 415.950 625.050 416.400 ;
        RECT 627.000 415.950 631.050 416.400 ;
        RECT 634.950 415.950 637.050 418.050 ;
        RECT 640.950 417.450 643.050 418.050 ;
        RECT 649.950 417.450 652.050 418.050 ;
        RECT 640.950 416.400 652.050 417.450 ;
        RECT 640.950 415.950 643.050 416.400 ;
        RECT 649.950 415.950 652.050 416.400 ;
        RECT 658.950 415.950 661.050 418.050 ;
        RECT 682.950 415.950 685.050 418.050 ;
        RECT 697.950 415.950 700.050 417.750 ;
        RECT 703.950 415.950 706.050 417.750 ;
        RECT 709.950 415.950 712.050 421.050 ;
        RECT 760.950 418.950 763.050 421.050 ;
        RECT 766.950 418.950 769.050 421.050 ;
        RECT 781.950 418.950 784.050 421.050 ;
        RECT 787.950 418.950 790.050 421.050 ;
        RECT 823.950 418.950 826.050 421.050 ;
        RECT 829.950 418.950 832.050 421.050 ;
        RECT 844.950 418.950 847.050 421.050 ;
        RECT 850.950 418.950 853.050 421.050 ;
        RECT 889.950 418.950 892.050 421.050 ;
        RECT 895.950 418.950 898.050 421.050 ;
        RECT 715.950 415.950 718.050 418.050 ;
        RECT 721.950 417.450 724.050 418.050 ;
        RECT 730.950 417.450 733.050 418.050 ;
        RECT 721.950 416.400 733.050 417.450 ;
        RECT 721.950 415.950 724.050 416.400 ;
        RECT 730.950 415.950 733.050 416.400 ;
        RECT 745.950 415.950 748.050 418.050 ;
        RECT 760.950 415.950 763.050 417.750 ;
        RECT 766.950 415.950 769.050 417.750 ;
        RECT 781.950 415.950 784.050 417.750 ;
        RECT 787.950 415.950 790.050 417.750 ;
        RECT 799.950 415.950 802.050 418.050 ;
        RECT 805.950 417.450 808.050 418.050 ;
        RECT 814.950 417.450 817.050 418.050 ;
        RECT 805.950 416.400 817.050 417.450 ;
        RECT 805.950 415.950 808.050 416.400 ;
        RECT 814.950 415.950 817.050 416.400 ;
        RECT 823.950 415.950 826.050 417.750 ;
        RECT 829.950 415.950 832.050 417.750 ;
        RECT 844.950 415.950 847.050 417.750 ;
        RECT 850.950 415.950 853.050 417.750 ;
        RECT 871.950 415.950 874.050 418.050 ;
        RECT 889.950 415.950 892.050 417.750 ;
        RECT 895.950 415.950 898.050 417.750 ;
        RECT 241.950 412.950 244.050 414.750 ;
        RECT 256.950 412.950 259.050 414.750 ;
        RECT 277.950 413.250 280.050 415.050 ;
        RECT 301.950 413.250 304.050 415.050 ;
        RECT 316.950 412.950 319.050 414.750 ;
        RECT 334.950 412.950 337.050 414.750 ;
        RECT 340.950 413.250 343.050 415.050 ;
        RECT 361.950 412.950 364.050 414.750 ;
        RECT 379.950 412.950 382.050 414.750 ;
        RECT 403.950 413.250 406.050 415.050 ;
        RECT 418.950 412.950 421.050 414.750 ;
        RECT 424.950 412.950 427.050 414.750 ;
        RECT 442.950 412.950 445.050 414.750 ;
        RECT 448.950 413.250 451.050 415.050 ;
        RECT 466.950 413.250 469.050 415.050 ;
        RECT 472.950 412.950 475.050 414.750 ;
        RECT 484.950 412.950 487.050 414.750 ;
        RECT 490.950 412.950 493.050 414.750 ;
        RECT 511.950 412.950 514.050 414.750 ;
        RECT 517.950 412.950 520.050 414.750 ;
        RECT 535.950 412.950 538.050 414.750 ;
        RECT 541.950 412.950 544.050 414.750 ;
        RECT 562.950 412.950 565.050 414.750 ;
        RECT 580.950 412.950 583.050 414.750 ;
        RECT 586.950 412.950 589.050 414.750 ;
        RECT 604.950 412.950 607.050 414.750 ;
        RECT 622.950 412.950 625.050 414.750 ;
        RECT 634.950 412.950 637.050 414.750 ;
        RECT 640.950 412.950 643.050 414.750 ;
        RECT 658.950 412.950 661.050 414.750 ;
        RECT 682.950 412.950 685.050 414.750 ;
        RECT 700.950 413.250 703.050 415.050 ;
        RECT 715.950 412.950 718.050 414.750 ;
        RECT 721.950 412.950 724.050 414.750 ;
        RECT 745.950 412.950 748.050 414.750 ;
        RECT 763.950 413.250 766.050 415.050 ;
        RECT 784.950 413.250 787.050 415.050 ;
        RECT 799.950 412.950 802.050 414.750 ;
        RECT 805.950 412.950 808.050 414.750 ;
        RECT 826.950 413.250 829.050 415.050 ;
        RECT 847.950 413.250 850.050 415.050 ;
        RECT 868.950 414.750 870.750 415.050 ;
        RECT 868.950 413.250 871.050 414.750 ;
        RECT 871.950 413.250 874.050 414.750 ;
        RECT 877.950 413.250 880.050 415.050 ;
        RECT 892.950 413.250 895.050 415.050 ;
        RECT 872.250 412.950 874.050 413.250 ;
        RECT 259.950 410.250 262.050 412.050 ;
        RECT 277.950 409.950 280.050 412.050 ;
        RECT 289.950 411.450 292.050 412.050 ;
        RECT 301.950 411.450 304.050 412.050 ;
        RECT 310.950 411.450 313.050 412.050 ;
        RECT 289.950 410.400 313.050 411.450 ;
        RECT 289.950 409.950 292.050 410.400 ;
        RECT 301.950 409.950 304.050 410.400 ;
        RECT 310.950 409.950 313.050 410.400 ;
        RECT 319.950 410.250 322.050 412.050 ;
        RECT 340.950 411.450 343.050 412.050 ;
        RECT 352.950 411.450 355.050 412.050 ;
        RECT 340.950 410.400 355.050 411.450 ;
        RECT 340.950 409.950 343.050 410.400 ;
        RECT 352.950 409.950 355.050 410.400 ;
        RECT 358.950 410.250 361.050 412.050 ;
        RECT 364.950 410.250 367.050 412.050 ;
        RECT 376.950 410.250 379.050 412.050 ;
        RECT 382.950 410.250 385.050 412.050 ;
        RECT 403.950 411.450 406.050 412.050 ;
        RECT 415.950 411.450 418.050 412.050 ;
        RECT 403.950 410.400 418.050 411.450 ;
        RECT 403.950 409.950 406.050 410.400 ;
        RECT 415.950 409.950 418.050 410.400 ;
        RECT 421.950 410.250 424.050 412.050 ;
        RECT 427.950 410.250 430.050 412.050 ;
        RECT 448.950 411.450 451.050 412.050 ;
        RECT 453.000 411.450 457.050 412.050 ;
        RECT 448.950 410.400 457.050 411.450 ;
        RECT 448.950 409.950 451.050 410.400 ;
        RECT 453.000 409.950 457.050 410.400 ;
        RECT 466.950 409.950 469.050 412.050 ;
        RECT 487.950 410.250 490.050 412.050 ;
        RECT 493.950 410.250 496.050 412.050 ;
        RECT 514.950 410.250 517.050 412.050 ;
        RECT 520.950 410.250 523.050 412.050 ;
        RECT 538.950 410.250 541.050 412.050 ;
        RECT 544.950 410.250 547.050 412.050 ;
        RECT 559.950 410.250 562.050 412.050 ;
        RECT 565.950 410.250 568.050 412.050 ;
        RECT 583.950 410.250 586.050 412.050 ;
        RECT 589.950 410.250 592.050 412.050 ;
        RECT 601.950 410.250 604.050 412.050 ;
        RECT 619.950 410.250 622.050 412.050 ;
        RECT 637.950 410.250 640.050 412.050 ;
        RECT 643.950 410.250 646.050 412.050 ;
        RECT 661.950 410.250 664.050 412.050 ;
        RECT 679.950 410.250 682.050 412.050 ;
        RECT 700.950 411.450 703.050 412.050 ;
        RECT 709.950 411.450 712.050 412.050 ;
        RECT 700.950 410.400 712.050 411.450 ;
        RECT 700.950 409.950 703.050 410.400 ;
        RECT 709.950 409.950 712.050 410.400 ;
        RECT 718.950 410.250 721.050 412.050 ;
        RECT 724.950 410.250 727.050 412.050 ;
        RECT 742.950 410.250 745.050 412.050 ;
        RECT 763.950 411.450 766.050 412.050 ;
        RECT 768.000 411.450 771.900 412.050 ;
        RECT 763.950 410.400 771.900 411.450 ;
        RECT 763.950 409.950 766.050 410.400 ;
        RECT 768.000 409.950 771.900 410.400 ;
        RECT 773.100 411.450 775.200 412.050 ;
        RECT 784.950 411.450 787.050 412.050 ;
        RECT 773.100 410.400 787.050 411.450 ;
        RECT 773.100 409.950 775.200 410.400 ;
        RECT 784.950 409.950 787.050 410.400 ;
        RECT 802.950 410.250 805.050 412.050 ;
        RECT 808.950 410.250 811.050 412.050 ;
        RECT 814.950 411.450 817.050 412.050 ;
        RECT 826.950 411.450 829.050 412.050 ;
        RECT 814.950 410.400 829.050 411.450 ;
        RECT 814.950 409.950 817.050 410.400 ;
        RECT 826.950 409.950 829.050 410.400 ;
        RECT 832.950 411.450 835.050 412.050 ;
        RECT 847.950 411.450 850.050 412.050 ;
        RECT 832.950 410.400 850.050 411.450 ;
        RECT 832.950 409.950 835.050 410.400 ;
        RECT 847.950 409.950 850.050 410.400 ;
        RECT 868.950 409.950 871.050 412.050 ;
        RECT 877.950 409.950 880.050 412.050 ;
        RECT 883.950 411.450 886.050 412.050 ;
        RECT 892.950 411.450 895.050 412.050 ;
        RECT 883.950 410.400 895.050 411.450 ;
        RECT 883.950 409.950 886.050 410.400 ;
        RECT 892.950 409.950 895.050 410.400 ;
        RECT 238.950 405.300 241.050 407.400 ;
        RECT 259.950 406.950 262.050 409.050 ;
        RECT 278.400 405.450 279.450 409.950 ;
        RECT 313.950 408.450 318.000 409.050 ;
        RECT 319.950 408.450 322.050 409.050 ;
        RECT 313.950 407.400 322.050 408.450 ;
        RECT 313.950 406.950 318.000 407.400 ;
        RECT 319.950 406.950 322.050 407.400 ;
        RECT 358.950 406.950 361.050 409.050 ;
        RECT 364.950 406.950 367.050 409.050 ;
        RECT 376.950 406.950 379.050 409.050 ;
        RECT 382.950 406.950 385.050 409.050 ;
        RECT 421.950 406.950 424.050 409.050 ;
        RECT 427.950 406.950 430.050 409.050 ;
        RECT 298.950 405.450 301.050 406.050 ;
        RECT 181.950 399.600 184.050 401.700 ;
        RECT 202.950 400.500 205.050 402.600 ;
        RECT 217.950 400.500 220.050 402.600 ;
        RECT 238.950 401.700 240.150 405.300 ;
        RECT 278.400 404.400 301.050 405.450 ;
        RECT 298.950 403.950 301.050 404.400 ;
        RECT 448.950 405.450 451.050 406.050 ;
        RECT 467.400 405.450 468.450 409.950 ;
        RECT 487.950 406.950 490.050 409.050 ;
        RECT 493.950 406.950 496.050 409.050 ;
        RECT 514.950 406.950 517.050 409.050 ;
        RECT 520.950 406.950 523.050 409.050 ;
        RECT 538.950 406.950 541.050 409.050 ;
        RECT 544.950 406.950 547.050 409.050 ;
        RECT 559.950 406.950 562.050 409.050 ;
        RECT 565.950 406.950 568.050 409.050 ;
        RECT 583.950 406.950 586.050 409.050 ;
        RECT 589.950 406.950 592.050 409.050 ;
        RECT 595.950 408.450 600.000 409.050 ;
        RECT 601.950 408.450 604.050 409.050 ;
        RECT 595.950 407.400 604.050 408.450 ;
        RECT 595.950 406.950 600.000 407.400 ;
        RECT 601.950 406.950 604.050 407.400 ;
        RECT 619.950 408.450 622.050 409.050 ;
        RECT 631.950 408.450 634.050 409.050 ;
        RECT 619.950 407.400 634.050 408.450 ;
        RECT 619.950 406.950 622.050 407.400 ;
        RECT 631.950 406.950 634.050 407.400 ;
        RECT 637.950 406.950 640.050 409.050 ;
        RECT 643.950 406.950 646.050 409.050 ;
        RECT 661.950 408.450 664.050 409.050 ;
        RECT 673.950 408.450 676.050 409.050 ;
        RECT 661.950 407.400 676.050 408.450 ;
        RECT 661.950 406.950 664.050 407.400 ;
        RECT 673.950 406.950 676.050 407.400 ;
        RECT 679.950 406.950 682.050 409.050 ;
        RECT 718.950 406.950 721.050 409.050 ;
        RECT 724.950 406.950 727.050 409.050 ;
        RECT 742.950 408.450 745.050 409.050 ;
        RECT 757.950 408.450 760.050 409.050 ;
        RECT 742.950 407.400 760.050 408.450 ;
        RECT 742.950 406.950 745.050 407.400 ;
        RECT 757.950 406.950 760.050 407.400 ;
        RECT 802.950 406.950 805.050 409.050 ;
        RECT 808.950 406.950 811.050 409.050 ;
        RECT 448.950 404.400 468.450 405.450 ;
        RECT 448.950 403.950 451.050 404.400 ;
        RECT 247.950 402.450 250.050 403.050 ;
        RECT 370.950 402.450 373.050 403.050 ;
        RECT 238.950 399.600 241.050 401.700 ;
        RECT 247.950 401.400 373.050 402.450 ;
        RECT 247.950 400.950 250.050 401.400 ;
        RECT 370.950 400.950 373.050 401.400 ;
        RECT 427.950 402.450 430.050 403.050 ;
        RECT 449.400 402.450 450.450 403.950 ;
        RECT 508.950 402.450 511.050 403.050 ;
        RECT 520.950 402.450 523.050 403.050 ;
        RECT 544.950 402.450 547.050 403.050 ;
        RECT 559.950 402.450 562.050 403.050 ;
        RECT 583.950 402.450 586.050 403.050 ;
        RECT 427.950 401.400 586.050 402.450 ;
        RECT 680.400 402.450 681.450 406.950 ;
        RECT 709.950 405.450 712.050 406.050 ;
        RECT 715.950 405.450 718.050 406.050 ;
        RECT 709.950 404.400 718.050 405.450 ;
        RECT 709.950 403.950 712.050 404.400 ;
        RECT 715.950 403.950 718.050 404.400 ;
        RECT 844.950 405.450 847.050 406.050 ;
        RECT 869.400 405.450 870.450 409.950 ;
        RECT 844.950 404.400 870.450 405.450 ;
        RECT 877.950 405.450 880.050 406.050 ;
        RECT 895.950 405.450 898.050 406.050 ;
        RECT 877.950 404.400 898.050 405.450 ;
        RECT 844.950 403.950 847.050 404.400 ;
        RECT 877.950 403.950 880.050 404.400 ;
        RECT 895.950 403.950 898.050 404.400 ;
        RECT 703.950 402.450 706.050 403.050 ;
        RECT 680.400 401.400 706.050 402.450 ;
        RECT 427.950 400.950 430.050 401.400 ;
        RECT 508.950 400.950 511.050 401.400 ;
        RECT 520.950 400.950 523.050 401.400 ;
        RECT 544.950 400.950 547.050 401.400 ;
        RECT 559.950 400.950 562.050 401.400 ;
        RECT 583.950 400.950 586.050 401.400 ;
        RECT 703.950 400.950 706.050 401.400 ;
        RECT 727.950 402.450 730.050 403.050 ;
        RECT 733.950 402.450 736.050 403.050 ;
        RECT 727.950 401.400 736.050 402.450 ;
        RECT 727.950 400.950 730.050 401.400 ;
        RECT 733.950 400.950 736.050 401.400 ;
        RECT 787.950 402.450 790.050 403.050 ;
        RECT 826.950 402.450 829.050 403.050 ;
        RECT 883.950 402.450 886.050 403.050 ;
        RECT 787.950 401.400 886.050 402.450 ;
        RECT 787.950 400.950 790.050 401.400 ;
        RECT 826.950 400.950 829.050 401.400 ;
        RECT 883.950 400.950 886.050 401.400 ;
        RECT 244.950 399.450 247.050 400.050 ;
        RECT 265.950 399.450 268.050 400.050 ;
        RECT 244.950 398.400 268.050 399.450 ;
        RECT 244.950 397.950 247.050 398.400 ;
        RECT 265.950 397.950 268.050 398.400 ;
        RECT 334.950 399.450 337.050 400.050 ;
        RECT 472.950 399.450 475.050 400.050 ;
        RECT 334.950 398.400 475.050 399.450 ;
        RECT 334.950 397.950 337.050 398.400 ;
        RECT 472.950 397.950 475.050 398.400 ;
        RECT 505.950 399.450 508.050 400.050 ;
        RECT 622.950 399.450 625.050 400.050 ;
        RECT 697.950 399.450 700.050 400.050 ;
        RECT 724.950 399.450 727.050 400.050 ;
        RECT 505.950 398.400 727.050 399.450 ;
        RECT 505.950 397.950 508.050 398.400 ;
        RECT 622.950 397.950 625.050 398.400 ;
        RECT 697.950 397.950 700.050 398.400 ;
        RECT 724.950 397.950 727.050 398.400 ;
        RECT 745.950 399.450 748.050 400.050 ;
        RECT 793.950 399.450 796.050 400.050 ;
        RECT 745.950 398.400 796.050 399.450 ;
        RECT 745.950 397.950 748.050 398.400 ;
        RECT 793.950 397.950 796.050 398.400 ;
        RECT 58.950 396.450 61.050 397.050 ;
        RECT 88.950 396.450 91.050 397.050 ;
        RECT 58.950 395.400 91.050 396.450 ;
        RECT 58.950 394.950 61.050 395.400 ;
        RECT 88.950 394.950 91.050 395.400 ;
        RECT 151.950 396.450 154.050 397.050 ;
        RECT 247.950 396.450 250.050 397.050 ;
        RECT 151.950 395.400 250.050 396.450 ;
        RECT 151.950 394.950 154.050 395.400 ;
        RECT 247.950 394.950 250.050 395.400 ;
        RECT 310.950 396.450 313.050 397.050 ;
        RECT 322.950 396.450 325.050 397.050 ;
        RECT 310.950 395.400 325.050 396.450 ;
        RECT 310.950 394.950 313.050 395.400 ;
        RECT 322.950 394.950 325.050 395.400 ;
        RECT 331.950 396.450 334.050 397.050 ;
        RECT 412.950 396.450 415.050 397.050 ;
        RECT 442.950 396.450 445.050 397.050 ;
        RECT 331.950 395.400 445.050 396.450 ;
        RECT 331.950 394.950 334.050 395.400 ;
        RECT 412.950 394.950 415.050 395.400 ;
        RECT 442.950 394.950 445.050 395.400 ;
        RECT 538.950 396.450 541.050 397.050 ;
        RECT 568.950 396.450 571.050 397.050 ;
        RECT 538.950 395.400 571.050 396.450 ;
        RECT 538.950 394.950 541.050 395.400 ;
        RECT 568.950 394.950 571.050 395.400 ;
        RECT 577.950 396.450 580.050 397.050 ;
        RECT 595.950 396.450 598.050 397.050 ;
        RECT 688.950 396.450 691.050 397.050 ;
        RECT 577.950 395.400 598.050 396.450 ;
        RECT 577.950 394.950 580.050 395.400 ;
        RECT 595.950 394.950 598.050 395.400 ;
        RECT 599.400 395.400 691.050 396.450 ;
        RECT 160.950 393.450 163.050 394.050 ;
        RECT 196.950 393.450 199.050 394.050 ;
        RECT 160.950 392.400 199.050 393.450 ;
        RECT 160.950 391.950 163.050 392.400 ;
        RECT 196.950 391.950 199.050 392.400 ;
        RECT 247.950 393.450 250.050 394.050 ;
        RECT 259.950 393.450 262.050 394.050 ;
        RECT 247.950 392.400 262.050 393.450 ;
        RECT 247.950 391.950 250.050 392.400 ;
        RECT 259.950 391.950 262.050 392.400 ;
        RECT 382.950 393.450 385.050 394.050 ;
        RECT 403.950 393.450 406.050 394.050 ;
        RECT 382.950 392.400 406.050 393.450 ;
        RECT 382.950 391.950 385.050 392.400 ;
        RECT 403.950 391.950 406.050 392.400 ;
        RECT 466.950 393.450 469.050 394.050 ;
        RECT 472.950 393.450 475.050 394.050 ;
        RECT 599.400 393.450 600.450 395.400 ;
        RECT 688.950 394.950 691.050 395.400 ;
        RECT 727.950 394.950 733.050 397.050 ;
        RECT 808.950 396.450 811.050 397.050 ;
        RECT 814.950 396.450 817.050 397.050 ;
        RECT 808.950 395.400 817.050 396.450 ;
        RECT 808.950 394.950 811.050 395.400 ;
        RECT 814.950 394.950 817.050 395.400 ;
        RECT 466.950 392.400 600.450 393.450 ;
        RECT 733.950 393.450 736.050 394.050 ;
        RECT 814.950 393.450 817.050 394.050 ;
        RECT 733.950 392.400 817.050 393.450 ;
        RECT 466.950 391.950 469.050 392.400 ;
        RECT 472.950 391.950 475.050 392.400 ;
        RECT 733.950 391.950 736.050 392.400 ;
        RECT 814.950 391.950 817.050 392.400 ;
        RECT 214.950 390.450 217.050 391.050 ;
        RECT 170.400 389.400 217.050 390.450 ;
        RECT 170.400 388.050 171.450 389.400 ;
        RECT 214.950 388.950 217.050 389.400 ;
        RECT 397.950 390.450 400.050 391.050 ;
        RECT 412.950 390.450 415.050 391.050 ;
        RECT 454.950 390.450 457.050 391.050 ;
        RECT 397.950 389.400 457.050 390.450 ;
        RECT 397.950 388.950 400.050 389.400 ;
        RECT 412.950 388.950 415.050 389.400 ;
        RECT 454.950 388.950 457.050 389.400 ;
        RECT 802.950 390.450 805.050 391.050 ;
        RECT 835.950 390.450 838.050 391.050 ;
        RECT 802.950 389.400 838.050 390.450 ;
        RECT 802.950 388.950 805.050 389.400 ;
        RECT 835.950 388.950 838.050 389.400 ;
        RECT 40.950 387.450 43.050 388.050 ;
        RECT 67.950 387.450 70.050 388.050 ;
        RECT 169.950 387.450 172.050 388.050 ;
        RECT 40.950 386.400 172.050 387.450 ;
        RECT 40.950 385.950 43.050 386.400 ;
        RECT 67.950 385.950 70.050 386.400 ;
        RECT 169.950 385.950 172.050 386.400 ;
        RECT 178.950 387.450 181.050 388.050 ;
        RECT 184.950 387.450 187.050 388.050 ;
        RECT 178.950 386.400 187.050 387.450 ;
        RECT 178.950 385.950 181.050 386.400 ;
        RECT 184.950 385.950 187.050 386.400 ;
        RECT 229.950 387.450 232.050 388.050 ;
        RECT 433.950 387.450 436.050 388.050 ;
        RECT 229.950 386.400 436.050 387.450 ;
        RECT 229.950 385.950 232.050 386.400 ;
        RECT 433.950 385.950 436.050 386.400 ;
        RECT 475.950 387.450 478.050 388.050 ;
        RECT 520.950 387.450 523.050 388.050 ;
        RECT 475.950 386.400 523.050 387.450 ;
        RECT 475.950 385.950 478.050 386.400 ;
        RECT 520.950 385.950 523.050 386.400 ;
        RECT 826.950 387.450 829.050 388.050 ;
        RECT 844.950 387.450 847.050 388.050 ;
        RECT 826.950 386.400 847.050 387.450 ;
        RECT 826.950 385.950 829.050 386.400 ;
        RECT 844.950 385.950 847.050 386.400 ;
        RECT 643.950 384.450 646.050 385.050 ;
        RECT 652.950 384.450 655.050 385.050 ;
        RECT 685.950 384.450 688.050 385.050 ;
        RECT 643.950 383.400 688.050 384.450 ;
        RECT 7.950 381.300 10.050 383.400 ;
        RECT 8.850 377.700 10.050 381.300 ;
        RECT 28.950 380.400 31.050 382.500 ;
        RECT 43.950 380.400 46.050 382.500 ;
        RECT 64.950 381.300 67.050 383.400 ;
        RECT 106.950 381.450 109.050 382.050 ;
        RECT 130.950 381.450 133.050 382.050 ;
        RECT 7.950 375.600 10.050 377.700 ;
        RECT 4.950 368.250 7.050 370.050 ;
        RECT 4.950 364.950 7.050 367.050 ;
        RECT 8.850 360.600 10.050 375.600 ;
        RECT 19.950 370.950 25.050 373.050 ;
        RECT 22.950 367.950 25.050 369.750 ;
        RECT 29.100 360.600 30.300 380.400 ;
        RECT 31.950 370.950 34.050 373.050 ;
        RECT 40.950 370.950 43.050 373.050 ;
        RECT 31.950 367.950 34.050 369.750 ;
        RECT 40.950 367.950 43.050 369.750 ;
        RECT 44.700 360.600 45.900 380.400 ;
        RECT 64.950 377.700 66.150 381.300 ;
        RECT 106.950 380.400 133.050 381.450 ;
        RECT 106.950 379.950 109.050 380.400 ;
        RECT 130.950 379.950 133.050 380.400 ;
        RECT 190.950 381.450 193.050 382.050 ;
        RECT 202.950 381.450 205.050 382.050 ;
        RECT 190.950 380.400 205.050 381.450 ;
        RECT 190.950 379.950 193.050 380.400 ;
        RECT 202.950 379.950 205.050 380.400 ;
        RECT 274.950 381.450 277.050 382.050 ;
        RECT 280.950 381.450 283.050 382.050 ;
        RECT 274.950 380.400 283.050 381.450 ;
        RECT 274.950 379.950 277.050 380.400 ;
        RECT 280.950 379.950 283.050 380.400 ;
        RECT 316.950 381.450 319.050 382.050 ;
        RECT 352.950 381.450 355.050 382.050 ;
        RECT 316.950 380.400 355.050 381.450 ;
        RECT 406.950 381.300 409.050 383.400 ;
        RECT 316.950 379.950 319.050 380.400 ;
        RECT 352.950 379.950 355.050 380.400 ;
        RECT 223.950 378.450 226.050 379.050 ;
        RECT 229.950 378.450 232.050 379.050 ;
        RECT 247.950 378.450 250.050 379.050 ;
        RECT 49.950 370.950 52.050 376.050 ;
        RECT 64.950 375.600 67.050 377.700 ;
        RECT 223.950 377.400 250.050 378.450 ;
        RECT 407.850 377.700 409.050 381.300 ;
        RECT 427.950 380.400 430.050 382.500 ;
        RECT 454.950 381.450 457.050 382.050 ;
        RECT 460.950 381.450 463.050 382.050 ;
        RECT 454.950 380.400 463.050 381.450 ;
        RECT 490.950 380.400 493.050 382.500 ;
        RECT 511.950 381.300 514.050 383.400 ;
        RECT 610.950 381.300 613.050 383.400 ;
        RECT 643.950 382.950 646.050 383.400 ;
        RECT 652.950 382.950 655.050 383.400 ;
        RECT 685.950 382.950 688.050 383.400 ;
        RECT 223.950 376.950 226.050 377.400 ;
        RECT 229.950 376.950 232.050 377.400 ;
        RECT 247.950 376.950 250.050 377.400 ;
        RECT 49.950 367.950 52.050 369.750 ;
        RECT 64.950 360.600 66.150 375.600 ;
        RECT 85.950 373.950 88.050 376.050 ;
        RECT 106.950 373.950 109.050 376.050 ;
        RECT 112.950 373.950 115.050 376.050 ;
        RECT 145.950 373.950 148.050 376.050 ;
        RECT 169.950 373.950 172.050 376.050 ;
        RECT 175.950 373.950 178.050 376.050 ;
        RECT 181.950 373.950 187.050 376.050 ;
        RECT 190.950 373.950 193.050 376.050 ;
        RECT 196.950 373.950 199.050 376.050 ;
        RECT 214.950 373.950 217.050 376.050 ;
        RECT 220.950 373.950 223.050 376.050 ;
        RECT 280.950 373.950 283.050 376.050 ;
        RECT 286.950 373.950 289.050 376.050 ;
        RECT 292.950 375.450 295.050 376.050 ;
        RECT 301.950 375.450 304.050 376.050 ;
        RECT 292.950 374.400 304.050 375.450 ;
        RECT 292.950 373.950 295.050 374.400 ;
        RECT 301.950 373.950 304.050 374.400 ;
        RECT 307.950 375.450 310.050 376.050 ;
        RECT 316.950 375.450 319.050 376.050 ;
        RECT 307.950 374.400 319.050 375.450 ;
        RECT 307.950 373.950 310.050 374.400 ;
        RECT 316.950 373.950 319.050 374.400 ;
        RECT 322.950 373.950 325.050 376.050 ;
        RECT 328.950 373.950 331.050 376.050 ;
        RECT 346.950 373.950 349.050 376.050 ;
        RECT 352.950 373.950 355.050 376.050 ;
        RECT 391.950 373.950 394.050 376.050 ;
        RECT 397.950 373.950 400.050 376.050 ;
        RECT 406.950 375.600 409.050 377.700 ;
        RECT 85.950 370.950 88.050 372.750 ;
        RECT 106.950 370.950 109.050 372.750 ;
        RECT 112.950 370.950 115.050 372.750 ;
        RECT 118.950 372.450 121.050 373.050 ;
        RECT 130.950 372.450 133.050 373.050 ;
        RECT 139.950 372.450 142.050 373.050 ;
        RECT 118.950 371.400 142.050 372.450 ;
        RECT 118.950 370.950 121.050 371.400 ;
        RECT 130.950 370.950 133.050 371.400 ;
        RECT 139.950 370.950 142.050 371.400 ;
        RECT 145.950 370.950 148.050 372.750 ;
        RECT 154.950 372.450 157.050 373.050 ;
        RECT 159.000 372.450 163.050 373.050 ;
        RECT 154.950 371.400 163.050 372.450 ;
        RECT 154.950 370.950 157.050 371.400 ;
        RECT 159.000 370.950 163.050 371.400 ;
        RECT 169.950 370.950 172.050 372.750 ;
        RECT 175.950 370.950 178.050 372.750 ;
        RECT 190.950 370.950 193.050 372.750 ;
        RECT 196.950 370.950 199.050 372.750 ;
        RECT 214.950 370.950 217.050 372.750 ;
        RECT 220.950 370.950 223.050 372.750 ;
        RECT 238.950 372.450 241.050 373.050 ;
        RECT 256.950 372.450 259.050 373.050 ;
        RECT 238.950 371.400 259.050 372.450 ;
        RECT 238.950 370.950 241.050 371.400 ;
        RECT 256.950 370.950 259.050 371.400 ;
        RECT 262.950 372.450 265.050 373.050 ;
        RECT 274.950 372.450 277.050 373.050 ;
        RECT 262.950 371.400 277.050 372.450 ;
        RECT 262.950 370.950 265.050 371.400 ;
        RECT 274.950 370.950 277.050 371.400 ;
        RECT 280.950 370.950 283.050 372.750 ;
        RECT 286.950 370.950 289.050 372.750 ;
        RECT 301.950 370.950 304.050 372.750 ;
        RECT 307.950 370.950 310.050 372.750 ;
        RECT 322.950 370.950 325.050 372.750 ;
        RECT 328.950 370.950 331.050 372.750 ;
        RECT 346.950 370.950 349.050 372.750 ;
        RECT 352.950 370.950 355.050 372.750 ;
        RECT 370.950 372.450 373.050 373.050 ;
        RECT 385.950 372.450 388.050 373.050 ;
        RECT 370.950 371.400 388.050 372.450 ;
        RECT 370.950 370.950 373.050 371.400 ;
        RECT 385.950 370.950 388.050 371.400 ;
        RECT 391.950 370.950 394.050 372.750 ;
        RECT 397.950 370.950 400.050 372.750 ;
        RECT 67.950 368.250 70.050 370.050 ;
        RECT 88.950 368.250 91.050 370.050 ;
        RECT 103.950 368.250 106.050 370.050 ;
        RECT 109.950 368.250 112.050 370.050 ;
        RECT 130.950 367.950 133.050 369.750 ;
        RECT 148.950 368.250 151.050 370.050 ;
        RECT 154.950 367.950 157.050 369.750 ;
        RECT 172.950 368.250 175.050 370.050 ;
        RECT 184.950 367.050 187.050 370.050 ;
        RECT 193.950 368.250 196.050 370.050 ;
        RECT 217.950 368.250 220.050 370.050 ;
        RECT 223.950 368.250 226.050 370.050 ;
        RECT 238.950 367.950 241.050 369.750 ;
        RECT 262.950 367.950 265.050 369.750 ;
        RECT 268.950 369.450 271.050 370.050 ;
        RECT 277.950 369.450 280.050 370.050 ;
        RECT 268.950 368.400 280.050 369.450 ;
        RECT 268.950 367.950 271.050 368.400 ;
        RECT 277.950 367.950 280.050 368.400 ;
        RECT 283.950 368.250 286.050 370.050 ;
        RECT 298.950 368.250 301.050 370.050 ;
        RECT 304.950 368.250 307.050 370.050 ;
        RECT 325.950 368.250 328.050 370.050 ;
        RECT 349.950 368.250 352.050 370.050 ;
        RECT 370.950 367.950 373.050 369.750 ;
        RECT 388.950 368.250 391.050 370.050 ;
        RECT 394.950 368.250 397.050 370.050 ;
        RECT 403.950 368.250 406.050 370.050 ;
        RECT 67.950 364.950 70.050 367.050 ;
        RECT 88.950 364.950 91.050 367.050 ;
        RECT 103.950 361.950 106.050 367.050 ;
        RECT 109.950 364.950 112.050 367.050 ;
        RECT 127.950 365.250 130.050 367.050 ;
        RECT 133.950 365.250 136.050 367.050 ;
        RECT 148.950 364.950 151.050 367.050 ;
        RECT 172.950 366.450 175.050 367.050 ;
        RECT 181.800 366.450 183.900 367.050 ;
        RECT 172.950 365.400 183.900 366.450 ;
        RECT 184.950 366.000 187.200 367.050 ;
        RECT 172.950 364.950 175.050 365.400 ;
        RECT 181.800 364.950 183.900 365.400 ;
        RECT 185.100 364.950 187.200 366.000 ;
        RECT 193.950 366.450 196.050 367.050 ;
        RECT 198.000 366.450 202.050 367.050 ;
        RECT 193.950 365.400 202.050 366.450 ;
        RECT 193.950 364.950 196.050 365.400 ;
        RECT 198.000 364.950 202.050 365.400 ;
        RECT 205.950 366.450 208.050 367.050 ;
        RECT 217.950 366.450 220.050 367.050 ;
        RECT 205.950 365.400 220.050 366.450 ;
        RECT 205.950 364.950 208.050 365.400 ;
        RECT 217.950 364.950 220.050 365.400 ;
        RECT 223.950 364.950 226.050 367.050 ;
        RECT 235.950 365.250 238.050 367.050 ;
        RECT 241.950 365.250 244.050 367.050 ;
        RECT 259.950 365.250 262.050 367.050 ;
        RECT 265.950 365.250 268.050 367.050 ;
        RECT 283.950 364.950 286.050 367.050 ;
        RECT 298.950 364.950 301.050 367.050 ;
        RECT 304.950 366.450 307.050 367.050 ;
        RECT 316.950 366.450 319.050 367.050 ;
        RECT 304.950 365.400 319.050 366.450 ;
        RECT 304.950 364.950 307.050 365.400 ;
        RECT 316.950 364.950 319.050 365.400 ;
        RECT 127.950 361.950 130.050 364.050 ;
        RECT 133.950 361.950 136.050 364.050 ;
        RECT 235.950 363.450 238.050 364.050 ;
        RECT 230.400 362.400 238.050 363.450 ;
        RECT 7.950 358.500 10.050 360.600 ;
        RECT 28.950 358.500 31.050 360.600 ;
        RECT 43.950 358.500 46.050 360.600 ;
        RECT 64.950 358.500 67.050 360.600 ;
        RECT 109.950 360.450 112.050 361.050 ;
        RECT 118.950 360.450 121.050 361.050 ;
        RECT 109.950 359.400 121.050 360.450 ;
        RECT 109.950 358.950 112.050 359.400 ;
        RECT 118.950 358.950 121.050 359.400 ;
        RECT 139.950 360.450 142.050 361.050 ;
        RECT 148.950 360.450 151.050 361.050 ;
        RECT 166.950 360.450 169.050 361.050 ;
        RECT 139.950 359.400 169.050 360.450 ;
        RECT 139.950 358.950 142.050 359.400 ;
        RECT 148.950 358.950 151.050 359.400 ;
        RECT 166.950 358.950 169.050 359.400 ;
        RECT 223.950 360.450 226.050 361.050 ;
        RECT 230.400 360.450 231.450 362.400 ;
        RECT 235.950 361.950 238.050 362.400 ;
        RECT 241.950 363.450 244.050 364.050 ;
        RECT 246.000 363.450 250.050 364.050 ;
        RECT 241.950 362.400 250.050 363.450 ;
        RECT 241.950 361.950 244.050 362.400 ;
        RECT 246.000 361.950 250.050 362.400 ;
        RECT 259.950 361.950 262.050 364.050 ;
        RECT 265.950 361.950 268.050 364.050 ;
        RECT 223.950 359.400 231.450 360.450 ;
        RECT 271.950 360.450 274.050 361.050 ;
        RECT 284.400 360.450 285.450 364.950 ;
        RECT 325.950 361.950 328.050 367.050 ;
        RECT 349.950 361.950 352.050 367.050 ;
        RECT 367.950 365.250 370.050 367.050 ;
        RECT 373.950 365.250 376.050 367.050 ;
        RECT 379.950 366.450 382.050 367.050 ;
        RECT 388.950 366.450 391.050 367.050 ;
        RECT 379.950 365.400 391.050 366.450 ;
        RECT 379.950 364.950 382.050 365.400 ;
        RECT 388.950 364.950 391.050 365.400 ;
        RECT 394.950 364.950 397.050 367.050 ;
        RECT 403.950 364.950 406.050 367.050 ;
        RECT 364.950 361.950 370.050 364.050 ;
        RECT 373.950 361.950 376.050 364.050 ;
        RECT 346.950 360.450 349.050 361.050 ;
        RECT 407.850 360.600 409.050 375.600 ;
        RECT 421.950 370.950 424.050 373.050 ;
        RECT 421.950 367.950 424.050 369.750 ;
        RECT 428.100 360.600 429.300 380.400 ;
        RECT 454.950 379.950 457.050 380.400 ;
        RECT 460.950 379.950 463.050 380.400 ;
        RECT 448.950 373.950 451.050 376.050 ;
        RECT 454.950 373.950 457.050 376.050 ;
        RECT 469.950 373.950 472.050 376.050 ;
        RECT 475.950 373.950 478.050 376.050 ;
        RECT 430.950 370.950 433.050 373.050 ;
        RECT 448.950 370.950 451.050 372.750 ;
        RECT 454.950 370.950 457.050 372.750 ;
        RECT 469.950 370.950 472.050 372.750 ;
        RECT 475.950 370.950 478.050 372.750 ;
        RECT 487.950 370.950 490.050 373.050 ;
        RECT 430.950 367.950 433.050 369.750 ;
        RECT 445.950 368.250 448.050 370.050 ;
        RECT 451.950 368.250 454.050 370.050 ;
        RECT 472.950 368.250 475.050 370.050 ;
        RECT 478.950 368.250 481.050 370.050 ;
        RECT 487.950 367.950 490.050 369.750 ;
        RECT 445.950 364.950 448.050 367.050 ;
        RECT 451.950 361.950 454.050 367.050 ;
        RECT 472.950 364.950 475.050 367.050 ;
        RECT 478.950 364.950 484.050 367.050 ;
        RECT 271.950 359.400 349.050 360.450 ;
        RECT 223.950 358.950 226.050 359.400 ;
        RECT 271.950 358.950 274.050 359.400 ;
        RECT 346.950 358.950 349.050 359.400 ;
        RECT 406.950 358.500 409.050 360.600 ;
        RECT 427.950 358.500 430.050 360.600 ;
        RECT 475.950 360.450 478.050 361.050 ;
        RECT 484.950 360.450 487.050 361.050 ;
        RECT 491.700 360.600 492.900 380.400 ;
        RECT 511.950 377.700 513.150 381.300 ;
        RECT 517.950 378.450 520.050 379.050 ;
        RECT 547.950 378.450 550.050 379.050 ;
        RECT 511.950 375.600 514.050 377.700 ;
        RECT 517.950 377.400 550.050 378.450 ;
        RECT 611.850 377.700 613.050 381.300 ;
        RECT 631.950 380.400 634.050 382.500 ;
        RECT 649.950 381.450 652.050 382.050 ;
        RECT 658.950 381.450 661.050 382.050 ;
        RECT 649.950 380.400 661.050 381.450 ;
        RECT 517.950 376.950 520.050 377.400 ;
        RECT 547.950 376.950 550.050 377.400 ;
        RECT 496.950 370.950 499.050 373.050 ;
        RECT 496.950 367.950 499.050 369.750 ;
        RECT 511.950 360.600 513.150 375.600 ;
        RECT 553.950 373.950 556.050 376.050 ;
        RECT 559.950 373.950 562.050 376.050 ;
        RECT 574.950 373.950 577.050 376.050 ;
        RECT 580.950 373.950 583.050 376.050 ;
        RECT 598.950 373.950 601.050 376.050 ;
        RECT 610.950 375.600 613.050 377.700 ;
        RECT 520.950 372.450 523.050 373.050 ;
        RECT 532.950 372.450 535.050 373.050 ;
        RECT 520.950 371.400 535.050 372.450 ;
        RECT 520.950 370.950 523.050 371.400 ;
        RECT 532.950 370.950 535.050 371.400 ;
        RECT 553.950 370.950 556.050 372.750 ;
        RECT 559.950 370.950 562.050 372.750 ;
        RECT 574.950 370.950 577.050 372.750 ;
        RECT 580.950 370.950 583.050 372.750 ;
        RECT 598.950 370.950 601.050 372.750 ;
        RECT 514.950 368.250 517.050 370.050 ;
        RECT 532.950 367.950 535.050 369.750 ;
        RECT 556.950 368.250 559.050 370.050 ;
        RECT 577.950 368.250 580.050 370.050 ;
        RECT 583.950 368.250 586.050 370.050 ;
        RECT 595.950 368.250 598.050 370.050 ;
        RECT 607.950 368.250 610.050 370.050 ;
        RECT 514.950 364.950 517.050 367.050 ;
        RECT 529.950 365.250 532.050 367.050 ;
        RECT 535.950 365.250 538.050 367.050 ;
        RECT 556.950 366.450 559.050 367.050 ;
        RECT 571.950 366.450 574.050 367.050 ;
        RECT 556.950 365.400 574.050 366.450 ;
        RECT 556.950 364.950 559.050 365.400 ;
        RECT 571.950 364.950 574.050 365.400 ;
        RECT 577.950 364.950 580.050 367.050 ;
        RECT 583.950 364.950 586.050 367.050 ;
        RECT 595.950 364.950 598.050 367.050 ;
        RECT 607.950 364.950 610.050 367.050 ;
        RECT 520.950 363.450 523.050 364.050 ;
        RECT 529.950 363.450 532.050 364.050 ;
        RECT 520.950 362.400 532.050 363.450 ;
        RECT 520.950 361.950 523.050 362.400 ;
        RECT 529.950 361.950 532.050 362.400 ;
        RECT 535.950 361.950 538.050 364.050 ;
        RECT 475.950 359.400 487.050 360.450 ;
        RECT 475.950 358.950 478.050 359.400 ;
        RECT 484.950 358.950 487.050 359.400 ;
        RECT 490.950 358.500 493.050 360.600 ;
        RECT 511.950 358.500 514.050 360.600 ;
        RECT 571.950 360.450 574.050 361.050 ;
        RECT 577.950 360.450 580.050 361.050 ;
        RECT 611.850 360.600 613.050 375.600 ;
        RECT 625.950 370.950 628.050 373.050 ;
        RECT 625.950 367.950 628.050 369.750 ;
        RECT 632.100 360.600 633.300 380.400 ;
        RECT 649.950 379.950 652.050 380.400 ;
        RECT 658.950 379.950 661.050 380.400 ;
        RECT 709.950 381.450 712.050 382.050 ;
        RECT 721.950 381.450 724.050 382.050 ;
        RECT 709.950 380.400 724.050 381.450 ;
        RECT 742.950 380.400 745.050 382.500 ;
        RECT 763.950 381.300 766.050 383.400 ;
        RECT 769.950 381.450 772.050 382.200 ;
        RECT 787.950 381.450 790.050 382.050 ;
        RECT 709.950 379.950 712.050 380.400 ;
        RECT 721.950 379.950 724.050 380.400 ;
        RECT 634.950 378.450 637.050 379.050 ;
        RECT 640.950 378.450 643.050 379.050 ;
        RECT 634.950 377.400 643.050 378.450 ;
        RECT 634.950 376.950 637.050 377.400 ;
        RECT 640.950 376.950 643.050 377.400 ;
        RECT 673.950 378.450 676.050 379.050 ;
        RECT 691.950 378.450 694.050 379.050 ;
        RECT 673.950 377.400 694.050 378.450 ;
        RECT 673.950 376.950 676.050 377.400 ;
        RECT 691.950 376.950 694.050 377.400 ;
        RECT 652.950 373.950 655.050 376.050 ;
        RECT 658.950 373.950 661.050 376.050 ;
        RECT 685.950 375.450 688.050 376.050 ;
        RECT 697.950 375.450 700.050 376.050 ;
        RECT 685.950 374.400 700.050 375.450 ;
        RECT 685.950 373.950 688.050 374.400 ;
        RECT 697.950 373.950 700.050 374.400 ;
        RECT 703.950 373.950 706.050 376.050 ;
        RECT 721.950 373.950 724.050 376.050 ;
        RECT 727.950 373.950 730.050 376.050 ;
        RECT 634.950 370.950 637.050 373.050 ;
        RECT 652.950 370.950 655.050 372.750 ;
        RECT 658.950 370.950 661.050 372.750 ;
        RECT 664.950 372.450 667.050 373.050 ;
        RECT 679.950 372.450 682.050 373.050 ;
        RECT 664.950 371.400 682.050 372.450 ;
        RECT 664.950 370.950 667.050 371.400 ;
        RECT 679.950 370.950 682.050 371.400 ;
        RECT 697.950 370.950 700.050 372.750 ;
        RECT 703.950 370.950 706.050 372.750 ;
        RECT 721.950 370.950 724.050 372.750 ;
        RECT 727.950 370.950 730.050 372.750 ;
        RECT 739.950 370.950 742.050 373.050 ;
        RECT 634.950 367.950 637.050 369.750 ;
        RECT 649.950 368.250 652.050 370.050 ;
        RECT 655.950 368.250 658.050 370.050 ;
        RECT 661.950 368.250 664.050 370.050 ;
        RECT 679.950 367.950 682.050 369.750 ;
        RECT 700.950 368.250 703.050 370.050 ;
        RECT 706.950 368.250 709.050 370.050 ;
        RECT 724.950 368.250 727.050 370.050 ;
        RECT 730.950 368.250 733.050 370.050 ;
        RECT 739.950 367.950 742.050 369.750 ;
        RECT 649.950 364.950 652.050 367.050 ;
        RECT 655.950 364.950 658.050 367.050 ;
        RECT 661.950 364.950 664.050 367.050 ;
        RECT 676.950 365.250 679.050 367.050 ;
        RECT 682.950 365.250 685.050 367.050 ;
        RECT 700.950 364.950 703.050 367.050 ;
        RECT 706.950 364.950 712.050 367.050 ;
        RECT 724.950 364.950 727.050 367.050 ;
        RECT 730.950 366.450 733.050 367.050 ;
        RECT 735.000 366.450 739.050 367.050 ;
        RECT 730.950 365.400 739.050 366.450 ;
        RECT 730.950 364.950 733.050 365.400 ;
        RECT 735.000 364.950 739.050 365.400 ;
        RECT 571.950 359.400 580.050 360.450 ;
        RECT 571.950 358.950 574.050 359.400 ;
        RECT 577.950 358.950 580.050 359.400 ;
        RECT 610.950 358.500 613.050 360.600 ;
        RECT 631.950 358.500 634.050 360.600 ;
        RECT 640.950 360.450 643.050 361.050 ;
        RECT 656.400 360.450 657.450 364.950 ;
        RECT 676.950 361.950 679.050 364.050 ;
        RECT 682.950 361.950 685.050 364.050 ;
        RECT 640.950 359.400 657.450 360.450 ;
        RECT 691.950 360.450 694.050 361.050 ;
        RECT 700.950 360.450 703.050 361.050 ;
        RECT 743.700 360.600 744.900 380.400 ;
        RECT 748.950 378.450 751.050 379.050 ;
        RECT 757.950 378.450 760.050 379.050 ;
        RECT 748.950 377.400 760.050 378.450 ;
        RECT 748.950 376.950 751.050 377.400 ;
        RECT 757.950 376.950 760.050 377.400 ;
        RECT 763.950 377.700 765.150 381.300 ;
        RECT 769.950 380.400 790.050 381.450 ;
        RECT 769.950 380.100 772.050 380.400 ;
        RECT 787.950 379.950 790.050 380.400 ;
        RECT 793.950 381.450 796.050 382.050 ;
        RECT 814.950 381.450 817.050 382.050 ;
        RECT 793.950 380.400 817.050 381.450 ;
        RECT 874.950 380.400 877.050 382.500 ;
        RECT 895.950 381.300 898.050 383.400 ;
        RECT 793.950 379.950 796.050 380.400 ;
        RECT 814.950 379.950 817.050 380.400 ;
        RECT 769.950 378.450 772.050 378.900 ;
        RECT 763.950 375.600 766.050 377.700 ;
        RECT 769.950 377.400 789.450 378.450 ;
        RECT 769.950 376.800 772.050 377.400 ;
        RECT 748.950 370.950 751.050 373.050 ;
        RECT 748.950 367.950 751.050 369.750 ;
        RECT 763.950 360.600 765.150 375.600 ;
        RECT 788.400 373.050 789.450 377.400 ;
        RECT 808.950 373.950 811.050 376.050 ;
        RECT 814.950 373.950 817.050 376.050 ;
        RECT 841.950 373.950 844.050 376.050 ;
        RECT 856.950 373.950 859.050 376.050 ;
        RECT 862.950 373.950 865.050 376.050 ;
        RECT 781.950 370.950 784.050 373.050 ;
        RECT 787.950 370.950 790.050 373.050 ;
        RECT 793.950 370.950 796.050 373.050 ;
        RECT 808.950 370.950 811.050 372.750 ;
        RECT 814.950 370.950 817.050 372.750 ;
        RECT 820.950 372.450 823.050 373.050 ;
        RECT 832.950 372.450 835.050 373.050 ;
        RECT 820.950 371.400 835.050 372.450 ;
        RECT 820.950 370.950 823.050 371.400 ;
        RECT 832.950 370.950 835.050 371.400 ;
        RECT 841.950 370.950 844.050 372.750 ;
        RECT 856.950 370.950 859.050 372.750 ;
        RECT 862.950 370.950 865.050 372.750 ;
        RECT 871.950 370.950 874.050 373.050 ;
        RECT 766.950 368.250 769.050 370.050 ;
        RECT 781.950 367.950 784.050 369.750 ;
        RECT 787.950 367.950 790.050 369.750 ;
        RECT 793.950 367.950 796.050 369.750 ;
        RECT 811.950 368.250 814.050 370.050 ;
        RECT 832.950 367.950 835.050 369.750 ;
        RECT 838.950 368.250 841.050 370.050 ;
        RECT 853.950 368.250 856.050 370.050 ;
        RECT 859.950 368.250 862.050 370.050 ;
        RECT 871.950 367.950 874.050 369.750 ;
        RECT 766.950 364.950 769.050 367.050 ;
        RECT 784.950 365.250 787.050 367.050 ;
        RECT 790.950 365.250 793.050 367.050 ;
        RECT 811.950 366.450 814.050 367.050 ;
        RECT 829.950 366.450 832.050 367.050 ;
        RECT 811.950 365.400 832.050 366.450 ;
        RECT 811.950 364.950 814.050 365.400 ;
        RECT 829.950 364.950 832.050 365.400 ;
        RECT 838.950 366.450 841.050 367.050 ;
        RECT 847.950 366.450 850.050 367.050 ;
        RECT 838.950 365.400 850.050 366.450 ;
        RECT 838.950 364.950 841.050 365.400 ;
        RECT 847.950 364.950 850.050 365.400 ;
        RECT 853.950 364.950 856.050 367.050 ;
        RECT 859.950 364.950 865.050 367.050 ;
        RECT 784.950 361.950 787.050 364.050 ;
        RECT 790.950 361.950 793.050 364.050 ;
        RECT 691.950 359.400 703.050 360.450 ;
        RECT 640.950 358.950 643.050 359.400 ;
        RECT 691.950 358.950 694.050 359.400 ;
        RECT 700.950 358.950 703.050 359.400 ;
        RECT 742.950 358.500 745.050 360.600 ;
        RECT 763.950 358.500 766.050 360.600 ;
        RECT 796.950 360.450 799.050 361.050 ;
        RECT 820.950 360.450 823.050 361.050 ;
        RECT 796.950 359.400 823.050 360.450 ;
        RECT 796.950 358.950 799.050 359.400 ;
        RECT 820.950 358.950 823.050 359.400 ;
        RECT 829.950 360.450 832.050 361.050 ;
        RECT 838.800 360.450 840.900 361.050 ;
        RECT 829.950 359.400 840.900 360.450 ;
        RECT 829.950 358.950 832.050 359.400 ;
        RECT 838.800 358.950 840.900 359.400 ;
        RECT 842.100 360.450 844.200 361.050 ;
        RECT 856.950 360.450 859.050 361.050 ;
        RECT 875.700 360.600 876.900 380.400 ;
        RECT 895.950 377.700 897.150 381.300 ;
        RECT 895.950 375.600 898.050 377.700 ;
        RECT 880.950 370.950 883.050 373.050 ;
        RECT 880.950 367.950 883.050 369.750 ;
        RECT 895.950 360.600 897.150 375.600 ;
        RECT 898.950 368.250 901.050 370.050 ;
        RECT 898.950 364.950 901.050 367.050 ;
        RECT 842.100 359.400 859.050 360.450 ;
        RECT 842.100 358.950 844.200 359.400 ;
        RECT 856.950 358.950 859.050 359.400 ;
        RECT 874.950 358.500 877.050 360.600 ;
        RECT 895.950 358.500 898.050 360.600 ;
        RECT 112.950 357.450 115.050 358.050 ;
        RECT 145.950 357.450 148.050 358.050 ;
        RECT 193.950 357.450 196.050 358.050 ;
        RECT 202.950 357.450 205.050 358.050 ;
        RECT 112.950 356.400 177.450 357.450 ;
        RECT 112.950 355.950 115.050 356.400 ;
        RECT 145.950 355.950 148.050 356.400 ;
        RECT 176.400 355.050 177.450 356.400 ;
        RECT 193.950 356.400 205.050 357.450 ;
        RECT 193.950 355.950 196.050 356.400 ;
        RECT 202.950 355.950 205.050 356.400 ;
        RECT 229.950 355.950 235.050 358.050 ;
        RECT 265.950 357.450 268.050 358.050 ;
        RECT 292.950 357.450 295.050 358.050 ;
        RECT 265.950 356.400 295.050 357.450 ;
        RECT 265.950 355.950 268.050 356.400 ;
        RECT 292.950 355.950 295.050 356.400 ;
        RECT 664.950 357.450 667.050 358.050 ;
        RECT 694.950 357.450 697.050 358.050 ;
        RECT 715.950 357.450 718.050 358.050 ;
        RECT 664.950 356.400 718.050 357.450 ;
        RECT 664.950 355.950 667.050 356.400 ;
        RECT 694.950 355.950 697.050 356.400 ;
        RECT 715.950 355.950 718.050 356.400 ;
        RECT 823.950 355.950 829.050 358.050 ;
        RECT 25.950 354.450 28.050 355.050 ;
        RECT 31.950 354.450 34.050 355.050 ;
        RECT 40.950 354.450 43.050 355.050 ;
        RECT 25.950 353.400 43.050 354.450 ;
        RECT 25.950 352.950 28.050 353.400 ;
        RECT 31.950 352.950 34.050 353.400 ;
        RECT 40.950 352.950 43.050 353.400 ;
        RECT 67.950 354.450 70.050 355.050 ;
        RECT 88.950 354.450 91.050 355.050 ;
        RECT 67.950 353.400 91.050 354.450 ;
        RECT 67.950 352.950 70.050 353.400 ;
        RECT 88.950 352.950 91.050 353.400 ;
        RECT 175.950 354.450 178.050 355.050 ;
        RECT 205.950 354.450 208.050 355.050 ;
        RECT 175.950 353.400 208.050 354.450 ;
        RECT 175.950 352.950 178.050 353.400 ;
        RECT 205.950 352.950 208.050 353.400 ;
        RECT 220.950 354.450 223.050 355.050 ;
        RECT 244.950 354.450 247.050 355.050 ;
        RECT 220.950 353.400 247.050 354.450 ;
        RECT 220.950 352.950 223.050 353.400 ;
        RECT 244.950 352.950 247.050 353.400 ;
        RECT 295.950 354.450 298.050 355.050 ;
        RECT 334.950 354.450 337.050 355.050 ;
        RECT 295.950 353.400 337.050 354.450 ;
        RECT 295.950 352.950 298.050 353.400 ;
        RECT 334.950 352.950 337.050 353.400 ;
        RECT 355.950 354.450 358.050 355.050 ;
        RECT 373.950 354.450 376.050 355.050 ;
        RECT 412.950 354.450 415.050 355.050 ;
        RECT 355.950 353.400 415.050 354.450 ;
        RECT 355.950 352.950 358.050 353.400 ;
        RECT 373.950 352.950 376.050 353.400 ;
        RECT 412.950 352.950 415.050 353.400 ;
        RECT 424.950 354.450 427.050 355.050 ;
        RECT 475.950 354.450 478.050 355.050 ;
        RECT 424.950 353.400 478.050 354.450 ;
        RECT 424.950 352.950 427.050 353.400 ;
        RECT 475.950 352.950 478.050 353.400 ;
        RECT 481.950 354.450 484.050 355.050 ;
        RECT 496.950 354.450 499.050 355.050 ;
        RECT 481.950 353.400 499.050 354.450 ;
        RECT 481.950 352.950 484.050 353.400 ;
        RECT 496.950 352.950 499.050 353.400 ;
        RECT 505.950 354.450 508.050 355.050 ;
        RECT 526.950 354.450 529.050 355.050 ;
        RECT 505.950 353.400 529.050 354.450 ;
        RECT 505.950 352.950 508.050 353.400 ;
        RECT 526.950 352.950 529.050 353.400 ;
        RECT 574.950 354.450 577.050 355.050 ;
        RECT 601.950 354.450 604.050 355.050 ;
        RECT 637.950 354.450 640.050 355.050 ;
        RECT 574.950 353.400 640.050 354.450 ;
        RECT 574.950 352.950 577.050 353.400 ;
        RECT 601.950 352.950 604.050 353.400 ;
        RECT 637.950 352.950 640.050 353.400 ;
        RECT 736.950 354.450 739.050 355.050 ;
        RECT 856.950 354.450 859.050 355.050 ;
        RECT 736.950 353.400 859.050 354.450 ;
        RECT 736.950 352.950 739.050 353.400 ;
        RECT 196.950 351.450 199.050 352.050 ;
        RECT 208.950 351.450 211.050 352.050 ;
        RECT 196.950 350.400 211.050 351.450 ;
        RECT 196.950 349.950 199.050 350.400 ;
        RECT 208.950 349.950 211.050 350.400 ;
        RECT 214.950 351.450 217.050 352.050 ;
        RECT 271.950 351.450 274.050 352.050 ;
        RECT 214.950 350.400 274.050 351.450 ;
        RECT 214.950 349.950 217.050 350.400 ;
        RECT 271.950 349.950 274.050 350.400 ;
        RECT 388.950 351.450 391.050 352.050 ;
        RECT 430.950 351.450 433.050 352.050 ;
        RECT 442.950 351.450 445.050 352.050 ;
        RECT 388.950 350.400 445.050 351.450 ;
        RECT 388.950 349.950 391.050 350.400 ;
        RECT 430.950 349.950 433.050 350.400 ;
        RECT 442.950 349.950 445.050 350.400 ;
        RECT 460.950 351.450 463.050 352.050 ;
        RECT 469.950 351.450 472.050 352.050 ;
        RECT 460.950 350.400 472.050 351.450 ;
        RECT 460.950 349.950 463.050 350.400 ;
        RECT 469.950 349.950 472.050 350.400 ;
        RECT 487.950 351.450 490.050 352.200 ;
        RECT 502.950 351.450 505.050 352.050 ;
        RECT 535.950 351.450 538.050 352.050 ;
        RECT 487.950 350.400 505.050 351.450 ;
        RECT 487.950 350.100 490.050 350.400 ;
        RECT 502.950 349.950 505.050 350.400 ;
        RECT 512.400 350.400 538.050 351.450 ;
        RECT 512.400 349.050 513.450 350.400 ;
        RECT 535.950 349.950 538.050 350.400 ;
        RECT 586.950 351.450 589.050 352.050 ;
        RECT 595.950 351.450 598.050 352.050 ;
        RECT 586.950 350.400 598.050 351.450 ;
        RECT 586.950 349.950 589.050 350.400 ;
        RECT 595.950 349.950 598.050 350.400 ;
        RECT 685.950 351.450 688.050 352.050 ;
        RECT 784.950 351.450 787.050 352.050 ;
        RECT 685.950 350.400 787.050 351.450 ;
        RECT 685.950 349.950 688.050 350.400 ;
        RECT 784.950 349.950 787.050 350.400 ;
        RECT 832.950 349.950 835.050 353.400 ;
        RECT 856.950 352.950 859.050 353.400 ;
        RECT 865.950 354.450 868.050 355.050 ;
        RECT 871.950 354.450 874.050 355.050 ;
        RECT 865.950 353.400 874.050 354.450 ;
        RECT 865.950 352.950 868.050 353.400 ;
        RECT 871.950 352.950 874.050 353.400 ;
        RECT 85.950 348.450 88.050 349.050 ;
        RECT 68.400 347.400 88.050 348.450 ;
        RECT 68.400 343.050 69.450 347.400 ;
        RECT 85.950 346.950 88.050 347.400 ;
        RECT 217.950 348.450 220.050 349.050 ;
        RECT 238.950 348.450 241.050 349.050 ;
        RECT 217.950 347.400 241.050 348.450 ;
        RECT 217.950 346.950 220.050 347.400 ;
        RECT 238.950 346.950 241.050 347.400 ;
        RECT 412.950 348.450 415.050 349.050 ;
        RECT 436.950 348.450 439.050 349.050 ;
        RECT 412.950 347.400 439.050 348.450 ;
        RECT 412.950 346.950 415.050 347.400 ;
        RECT 436.950 346.950 439.050 347.400 ;
        RECT 487.950 348.450 490.050 348.900 ;
        RECT 511.950 348.450 514.050 349.050 ;
        RECT 487.950 347.400 514.050 348.450 ;
        RECT 487.950 346.800 490.050 347.400 ;
        RECT 511.950 346.950 514.050 347.400 ;
        RECT 607.950 348.450 610.050 349.050 ;
        RECT 613.950 348.450 616.050 349.050 ;
        RECT 607.950 347.400 616.050 348.450 ;
        RECT 607.950 346.950 610.050 347.400 ;
        RECT 613.950 346.950 616.050 347.400 ;
        RECT 631.950 348.450 634.050 349.050 ;
        RECT 646.950 348.450 649.050 349.050 ;
        RECT 631.950 347.400 649.050 348.450 ;
        RECT 631.950 346.950 634.050 347.400 ;
        RECT 646.950 346.950 649.050 347.400 ;
        RECT 862.950 348.450 865.050 349.050 ;
        RECT 871.950 348.450 874.050 349.050 ;
        RECT 862.950 347.400 874.050 348.450 ;
        RECT 862.950 346.950 865.050 347.400 ;
        RECT 871.950 346.950 874.050 347.400 ;
        RECT 67.950 340.950 70.050 343.050 ;
        RECT 73.950 342.450 76.050 343.050 ;
        RECT 82.950 342.450 85.050 343.050 ;
        RECT 73.950 341.400 85.050 342.450 ;
        RECT 73.950 340.950 76.050 341.400 ;
        RECT 82.950 340.950 85.050 341.400 ;
        RECT 88.950 340.950 91.050 346.050 ;
        RECT 112.950 345.450 115.050 346.050 ;
        RECT 107.400 344.400 115.050 345.450 ;
        RECT 121.950 344.400 124.050 346.500 ;
        RECT 142.950 344.400 145.050 346.500 ;
        RECT 181.950 344.400 184.050 346.500 ;
        RECT 202.950 344.400 205.050 346.500 ;
        RECT 208.950 345.450 211.050 346.050 ;
        RECT 244.950 345.450 247.050 346.050 ;
        RECT 208.950 344.400 247.050 345.450 ;
        RECT 94.950 342.450 97.050 343.050 ;
        RECT 107.400 342.450 108.450 344.400 ;
        RECT 112.950 343.950 115.050 344.400 ;
        RECT 94.950 341.400 108.450 342.450 ;
        RECT 94.950 340.950 97.050 341.400 ;
        RECT 4.950 339.450 9.000 340.050 ;
        RECT 10.950 339.450 13.050 340.050 ;
        RECT 4.950 338.400 13.050 339.450 ;
        RECT 4.950 337.950 9.000 338.400 ;
        RECT 10.950 337.950 13.050 338.400 ;
        RECT 34.950 337.950 37.050 340.050 ;
        RECT 52.950 337.950 55.050 340.050 ;
        RECT 67.950 337.950 70.050 339.750 ;
        RECT 73.950 337.950 76.050 339.750 ;
        RECT 88.950 337.950 91.050 339.750 ;
        RECT 94.950 337.950 97.050 339.750 ;
        RECT 112.950 337.950 115.050 340.050 ;
        RECT 118.950 337.950 121.050 340.050 ;
        RECT 10.950 334.950 13.050 336.750 ;
        RECT 34.950 334.950 37.050 336.750 ;
        RECT 52.950 334.950 55.050 336.750 ;
        RECT 70.950 335.250 73.050 337.050 ;
        RECT 91.950 335.250 94.050 337.050 ;
        RECT 112.950 334.950 115.050 336.750 ;
        RECT 118.950 334.950 121.050 336.750 ;
        RECT 13.950 332.250 16.050 334.050 ;
        RECT 31.950 332.250 34.050 334.050 ;
        RECT 49.950 332.250 52.050 334.050 ;
        RECT 55.950 333.450 58.050 334.050 ;
        RECT 70.950 333.450 73.050 334.050 ;
        RECT 75.000 333.450 79.050 334.050 ;
        RECT 55.950 332.400 79.050 333.450 ;
        RECT 55.950 331.950 58.050 332.400 ;
        RECT 70.950 331.950 73.050 332.400 ;
        RECT 75.000 331.950 79.050 332.400 ;
        RECT 85.950 333.450 90.000 334.050 ;
        RECT 91.950 333.450 94.050 334.050 ;
        RECT 85.950 332.400 94.050 333.450 ;
        RECT 85.950 331.950 90.000 332.400 ;
        RECT 91.950 331.950 94.050 332.400 ;
        RECT 109.950 332.250 112.050 334.050 ;
        RECT 13.950 328.950 19.050 331.050 ;
        RECT 31.950 325.950 34.050 331.050 ;
        RECT 49.950 328.950 55.050 331.050 ;
        RECT 109.950 328.950 112.050 331.050 ;
        RECT 122.850 329.400 124.050 344.400 ;
        RECT 136.950 335.250 139.050 337.050 ;
        RECT 136.950 331.950 139.050 334.050 ;
        RECT 121.950 327.300 124.050 329.400 ;
        RECT 82.950 324.450 85.050 325.050 ;
        RECT 109.950 324.450 112.050 325.050 ;
        RECT 82.950 323.400 112.050 324.450 ;
        RECT 122.850 323.700 124.050 327.300 ;
        RECT 143.100 324.600 144.300 344.400 ;
        RECT 145.950 342.450 148.050 343.050 ;
        RECT 160.950 342.450 163.050 343.050 ;
        RECT 145.950 341.400 163.050 342.450 ;
        RECT 145.950 340.950 148.050 341.400 ;
        RECT 160.950 340.950 163.050 341.400 ;
        RECT 166.950 337.950 169.050 340.050 ;
        RECT 172.950 337.950 175.050 340.050 ;
        RECT 145.950 335.250 148.050 337.050 ;
        RECT 166.950 334.950 169.050 336.750 ;
        RECT 172.950 334.950 175.050 336.750 ;
        RECT 178.950 335.250 181.050 337.050 ;
        RECT 145.950 331.950 148.050 334.050 ;
        RECT 163.950 332.250 166.050 334.050 ;
        RECT 169.950 332.250 172.050 334.050 ;
        RECT 178.950 331.950 181.050 334.050 ;
        RECT 163.950 328.950 166.050 331.050 ;
        RECT 169.950 328.950 172.050 331.050 ;
        RECT 182.700 324.600 183.900 344.400 ;
        RECT 187.950 335.250 190.050 337.050 ;
        RECT 187.950 333.450 190.050 334.050 ;
        RECT 196.950 333.450 199.050 334.050 ;
        RECT 187.950 332.400 199.050 333.450 ;
        RECT 187.950 331.950 190.050 332.400 ;
        RECT 196.950 331.950 199.050 332.400 ;
        RECT 202.950 329.400 204.150 344.400 ;
        RECT 208.950 343.950 211.050 344.400 ;
        RECT 244.950 343.950 247.050 344.400 ;
        RECT 262.950 345.450 265.050 346.050 ;
        RECT 295.950 345.450 298.050 346.050 ;
        RECT 262.950 344.400 298.050 345.450 ;
        RECT 262.950 343.950 265.050 344.400 ;
        RECT 295.950 343.950 298.050 344.400 ;
        RECT 316.950 345.450 319.050 346.050 ;
        RECT 328.950 345.450 331.050 346.050 ;
        RECT 316.950 344.400 336.450 345.450 ;
        RECT 364.950 344.400 367.050 346.500 ;
        RECT 385.950 344.400 388.050 346.500 ;
        RECT 424.950 345.450 427.050 346.050 ;
        RECT 433.950 345.450 436.050 346.050 ;
        RECT 424.950 344.400 436.050 345.450 ;
        RECT 445.950 344.400 448.050 346.500 ;
        RECT 466.950 344.400 469.050 346.500 ;
        RECT 526.950 344.400 529.050 346.500 ;
        RECT 547.950 344.400 550.050 346.500 ;
        RECT 562.950 344.400 565.050 346.500 ;
        RECT 583.950 344.400 586.050 346.500 ;
        RECT 676.950 345.450 679.050 346.050 ;
        RECT 685.950 345.450 688.050 346.050 ;
        RECT 676.950 344.400 688.050 345.450 ;
        RECT 733.950 344.400 736.050 346.500 ;
        RECT 754.950 344.400 757.050 346.500 ;
        RECT 760.950 345.450 763.050 346.050 ;
        RECT 778.950 345.450 781.050 346.050 ;
        RECT 811.950 345.450 814.050 346.050 ;
        RECT 760.950 344.400 781.050 345.450 ;
        RECT 316.950 343.950 319.050 344.400 ;
        RECT 328.950 343.950 331.050 344.400 ;
        RECT 335.400 340.050 336.450 344.400 ;
        RECT 340.950 342.450 343.050 343.050 ;
        RECT 349.950 342.450 352.050 343.050 ;
        RECT 340.950 341.400 352.050 342.450 ;
        RECT 340.950 340.950 343.050 341.400 ;
        RECT 349.950 340.950 352.050 341.400 ;
        RECT 355.950 340.950 358.050 343.050 ;
        RECT 205.950 337.950 208.050 340.050 ;
        RECT 211.950 339.450 214.050 340.050 ;
        RECT 220.950 339.450 223.050 340.050 ;
        RECT 211.950 338.400 223.050 339.450 ;
        RECT 211.950 337.950 214.050 338.400 ;
        RECT 220.950 337.950 223.050 338.400 ;
        RECT 238.950 337.950 241.050 340.050 ;
        RECT 244.950 337.950 247.050 340.050 ;
        RECT 262.950 337.950 265.050 340.050 ;
        RECT 271.950 339.450 274.050 340.050 ;
        RECT 286.950 339.450 289.050 340.050 ;
        RECT 271.950 338.400 289.050 339.450 ;
        RECT 271.950 337.950 274.050 338.400 ;
        RECT 286.950 337.950 289.050 338.400 ;
        RECT 313.950 337.950 316.050 340.050 ;
        RECT 334.950 337.950 337.050 340.050 ;
        RECT 349.950 337.950 352.050 339.750 ;
        RECT 355.950 337.950 358.050 339.750 ;
        RECT 361.950 337.950 364.050 340.050 ;
        RECT 205.950 334.950 208.050 336.750 ;
        RECT 220.950 334.950 223.050 336.750 ;
        RECT 238.950 334.950 241.050 336.750 ;
        RECT 244.950 334.950 247.050 336.750 ;
        RECT 262.950 334.950 265.050 336.750 ;
        RECT 268.950 335.250 271.050 337.050 ;
        RECT 286.950 334.950 289.050 336.750 ;
        RECT 307.950 335.250 310.050 337.050 ;
        RECT 313.950 334.950 316.050 336.750 ;
        RECT 328.950 335.250 331.050 337.050 ;
        RECT 334.950 334.950 337.050 336.750 ;
        RECT 352.950 335.250 355.050 337.050 ;
        RECT 361.950 334.950 364.050 336.750 ;
        RECT 223.950 332.250 226.050 334.050 ;
        RECT 241.950 332.250 244.050 334.050 ;
        RECT 247.950 332.250 250.050 334.050 ;
        RECT 268.950 331.950 274.050 334.050 ;
        RECT 283.950 332.250 286.050 334.050 ;
        RECT 289.950 332.250 292.050 334.050 ;
        RECT 307.950 331.950 313.050 334.050 ;
        RECT 316.950 333.450 319.050 334.050 ;
        RECT 328.950 333.450 331.050 334.050 ;
        RECT 316.950 332.400 331.050 333.450 ;
        RECT 316.950 331.950 319.050 332.400 ;
        RECT 328.950 331.950 331.050 332.400 ;
        RECT 352.950 331.950 358.050 334.050 ;
        RECT 223.950 330.450 226.050 331.050 ;
        RECT 223.950 329.400 237.450 330.450 ;
        RECT 202.950 327.300 205.050 329.400 ;
        RECT 223.950 328.950 226.050 329.400 ;
        RECT 236.400 328.050 237.450 329.400 ;
        RECT 241.950 328.950 244.050 331.050 ;
        RECT 247.950 328.950 250.050 331.050 ;
        RECT 253.950 330.450 256.050 331.050 ;
        RECT 262.950 330.450 265.050 331.050 ;
        RECT 253.950 329.400 265.050 330.450 ;
        RECT 253.950 328.950 256.050 329.400 ;
        RECT 262.950 328.950 265.050 329.400 ;
        RECT 283.950 328.950 286.050 331.050 ;
        RECT 289.950 328.950 292.050 331.050 ;
        RECT 365.850 329.400 367.050 344.400 ;
        RECT 379.950 335.250 382.050 337.050 ;
        RECT 379.950 331.950 382.050 334.050 ;
        RECT 82.950 322.950 85.050 323.400 ;
        RECT 109.950 322.950 112.050 323.400 ;
        RECT 121.950 321.600 124.050 323.700 ;
        RECT 142.950 322.500 145.050 324.600 ;
        RECT 181.950 322.500 184.050 324.600 ;
        RECT 202.950 323.700 204.150 327.300 ;
        RECT 236.400 326.400 241.050 328.050 ;
        RECT 364.950 327.300 367.050 329.400 ;
        RECT 237.000 325.950 241.050 326.400 ;
        RECT 220.950 324.450 223.050 325.050 ;
        RECT 235.950 324.450 238.050 325.050 ;
        RECT 271.950 324.450 274.050 325.050 ;
        RECT 283.950 324.450 286.050 325.050 ;
        RECT 202.950 321.600 205.050 323.700 ;
        RECT 220.950 323.400 286.050 324.450 ;
        RECT 220.950 322.950 223.050 323.400 ;
        RECT 235.950 322.950 238.050 323.400 ;
        RECT 271.950 322.950 274.050 323.400 ;
        RECT 283.950 322.950 286.050 323.400 ;
        RECT 289.950 324.450 292.050 325.050 ;
        RECT 340.950 324.450 343.050 325.050 ;
        RECT 289.950 323.400 343.050 324.450 ;
        RECT 365.850 323.700 367.050 327.300 ;
        RECT 386.100 324.600 387.300 344.400 ;
        RECT 424.950 343.950 427.050 344.400 ;
        RECT 433.950 343.950 436.050 344.400 ;
        RECT 403.950 340.950 409.050 343.050 ;
        RECT 412.950 340.950 415.050 343.050 ;
        RECT 406.950 337.950 409.050 339.750 ;
        RECT 412.950 337.950 415.050 339.750 ;
        RECT 421.950 339.450 426.000 340.050 ;
        RECT 427.950 339.450 430.050 340.050 ;
        RECT 421.950 338.400 430.050 339.450 ;
        RECT 421.950 337.950 426.000 338.400 ;
        RECT 427.950 337.950 430.050 338.400 ;
        RECT 433.950 337.950 436.050 340.050 ;
        RECT 388.950 335.250 391.050 337.050 ;
        RECT 409.950 335.250 412.050 337.050 ;
        RECT 427.950 334.950 430.050 336.750 ;
        RECT 433.950 334.950 436.050 336.750 ;
        RECT 442.950 335.250 445.050 337.050 ;
        RECT 388.950 331.950 391.050 334.050 ;
        RECT 409.950 333.450 412.050 334.050 ;
        RECT 421.950 333.450 424.050 334.050 ;
        RECT 409.950 332.400 424.050 333.450 ;
        RECT 409.950 331.950 412.050 332.400 ;
        RECT 421.950 331.950 424.050 332.400 ;
        RECT 430.950 332.250 433.050 334.050 ;
        RECT 436.950 332.250 439.050 334.050 ;
        RECT 442.950 331.950 445.050 334.050 ;
        RECT 430.950 328.950 433.050 331.050 ;
        RECT 436.950 328.950 439.050 331.050 ;
        RECT 446.700 324.600 447.900 344.400 ;
        RECT 451.950 335.250 454.050 337.050 ;
        RECT 451.950 331.950 454.050 334.050 ;
        RECT 466.950 329.400 468.150 344.400 ;
        RECT 511.950 340.950 514.050 343.050 ;
        RECT 517.950 340.950 520.050 343.050 ;
        RECT 469.950 337.950 472.050 340.050 ;
        RECT 487.950 337.950 490.050 340.050 ;
        RECT 493.950 339.450 496.050 340.050 ;
        RECT 505.950 339.450 508.050 340.050 ;
        RECT 493.950 338.400 508.050 339.450 ;
        RECT 493.950 337.950 496.050 338.400 ;
        RECT 505.950 337.950 508.050 338.400 ;
        RECT 511.950 337.950 514.050 339.750 ;
        RECT 517.950 337.950 520.050 339.750 ;
        RECT 523.950 337.950 526.050 340.050 ;
        RECT 469.950 334.950 472.050 336.750 ;
        RECT 487.950 334.950 490.050 336.750 ;
        RECT 493.950 334.950 496.050 336.750 ;
        RECT 514.950 335.250 517.050 337.050 ;
        RECT 523.950 334.950 526.050 336.750 ;
        RECT 484.950 332.250 487.050 334.050 ;
        RECT 490.950 332.250 493.050 334.050 ;
        RECT 496.950 333.450 499.050 334.050 ;
        RECT 514.950 333.450 517.050 334.050 ;
        RECT 496.950 332.400 517.050 333.450 ;
        RECT 496.950 331.950 499.050 332.400 ;
        RECT 514.950 331.950 517.050 332.400 ;
        RECT 475.950 330.450 478.050 331.050 ;
        RECT 484.950 330.450 487.050 331.050 ;
        RECT 475.950 329.400 487.050 330.450 ;
        RECT 466.950 327.300 469.050 329.400 ;
        RECT 475.950 328.950 478.050 329.400 ;
        RECT 484.950 328.950 487.050 329.400 ;
        RECT 490.950 328.950 493.050 331.050 ;
        RECT 527.850 329.400 529.050 344.400 ;
        RECT 541.950 335.250 544.050 337.050 ;
        RECT 541.950 331.950 544.050 334.050 ;
        RECT 505.950 327.450 508.050 328.050 ;
        RECT 520.950 327.450 523.050 328.050 ;
        RECT 289.950 322.950 292.050 323.400 ;
        RECT 340.950 322.950 343.050 323.400 ;
        RECT 364.950 321.600 367.050 323.700 ;
        RECT 385.950 322.500 388.050 324.600 ;
        RECT 445.950 322.500 448.050 324.600 ;
        RECT 466.950 323.700 468.150 327.300 ;
        RECT 505.950 326.400 523.050 327.450 ;
        RECT 526.950 327.300 529.050 329.400 ;
        RECT 505.950 325.950 508.050 326.400 ;
        RECT 520.950 325.950 523.050 326.400 ;
        RECT 481.950 324.450 484.050 325.050 ;
        RECT 487.950 324.450 490.050 325.050 ;
        RECT 466.950 321.600 469.050 323.700 ;
        RECT 481.950 323.400 490.050 324.450 ;
        RECT 527.850 323.700 529.050 327.300 ;
        RECT 532.950 327.450 535.050 328.050 ;
        RECT 541.950 327.450 544.050 328.050 ;
        RECT 532.950 326.400 544.050 327.450 ;
        RECT 532.950 325.950 535.050 326.400 ;
        RECT 541.950 325.950 544.050 326.400 ;
        RECT 548.100 324.600 549.300 344.400 ;
        RECT 550.950 335.250 553.050 337.050 ;
        RECT 559.950 335.250 562.050 337.050 ;
        RECT 550.950 331.950 553.050 334.050 ;
        RECT 559.950 331.950 562.050 334.050 ;
        RECT 563.700 324.600 564.900 344.400 ;
        RECT 568.950 335.250 571.050 337.050 ;
        RECT 568.950 331.950 574.050 334.050 ;
        RECT 583.950 329.400 585.150 344.400 ;
        RECT 676.950 343.950 679.050 344.400 ;
        RECT 685.950 343.950 688.050 344.400 ;
        RECT 595.950 342.450 600.000 343.050 ;
        RECT 601.950 342.450 604.050 343.050 ;
        RECT 595.950 341.400 604.050 342.450 ;
        RECT 595.950 340.950 600.000 341.400 ;
        RECT 601.950 340.950 604.050 341.400 ;
        RECT 607.950 340.950 610.050 343.050 ;
        RECT 637.950 340.950 643.050 343.050 ;
        RECT 646.950 340.950 649.050 343.050 ;
        RECT 688.950 340.950 691.050 343.050 ;
        RECT 694.950 340.950 697.050 343.050 ;
        RECT 586.950 337.950 589.050 340.050 ;
        RECT 601.950 337.950 604.050 339.750 ;
        RECT 607.950 337.950 610.050 339.750 ;
        RECT 613.950 339.450 616.050 340.050 ;
        RECT 622.950 339.450 625.050 340.050 ;
        RECT 613.950 338.400 625.050 339.450 ;
        RECT 613.950 337.950 616.050 338.400 ;
        RECT 622.950 337.950 625.050 338.400 ;
        RECT 640.950 337.950 643.050 339.750 ;
        RECT 646.950 337.950 649.050 339.750 ;
        RECT 664.950 337.950 667.050 340.050 ;
        RECT 670.950 339.450 673.050 340.050 ;
        RECT 682.950 339.450 685.050 340.050 ;
        RECT 670.950 338.400 685.050 339.450 ;
        RECT 670.950 337.950 673.050 338.400 ;
        RECT 682.950 337.950 685.050 338.400 ;
        RECT 688.950 337.950 691.050 339.750 ;
        RECT 694.950 337.950 697.050 339.750 ;
        RECT 715.950 337.950 718.050 340.050 ;
        RECT 586.950 334.950 589.050 336.750 ;
        RECT 604.950 335.250 607.050 337.050 ;
        RECT 622.950 334.950 625.050 336.750 ;
        RECT 643.950 335.250 646.050 337.050 ;
        RECT 664.950 334.950 667.050 336.750 ;
        RECT 670.950 334.950 673.050 336.750 ;
        RECT 685.950 335.250 688.050 337.050 ;
        RECT 691.950 335.250 694.050 337.050 ;
        RECT 697.950 335.250 700.050 337.050 ;
        RECT 715.950 334.950 718.050 336.750 ;
        RECT 721.950 335.250 724.050 337.050 ;
        RECT 730.950 335.250 733.050 337.050 ;
        RECT 583.950 327.300 586.050 329.400 ;
        RECT 604.950 328.950 607.050 334.050 ;
        RECT 625.950 332.250 628.050 334.050 ;
        RECT 640.950 331.950 646.050 334.050 ;
        RECT 661.950 332.250 664.050 334.050 ;
        RECT 667.950 332.250 670.050 334.050 ;
        RECT 685.950 331.950 688.050 334.050 ;
        RECT 625.950 330.450 628.050 331.050 ;
        RECT 630.000 330.450 634.050 331.050 ;
        RECT 625.950 329.400 634.050 330.450 ;
        RECT 625.950 328.950 628.050 329.400 ;
        RECT 630.000 328.950 634.050 329.400 ;
        RECT 661.950 328.950 664.050 331.050 ;
        RECT 667.950 330.450 670.050 331.050 ;
        RECT 676.950 330.450 679.050 331.050 ;
        RECT 667.950 329.400 679.050 330.450 ;
        RECT 667.950 328.950 670.050 329.400 ;
        RECT 676.950 328.950 679.050 329.400 ;
        RECT 691.950 328.950 694.050 334.050 ;
        RECT 697.950 331.950 700.050 334.050 ;
        RECT 712.950 332.250 715.050 334.050 ;
        RECT 718.950 331.950 724.050 334.050 ;
        RECT 730.950 331.950 733.050 334.050 ;
        RECT 712.950 328.950 715.050 331.050 ;
        RECT 481.950 322.950 484.050 323.400 ;
        RECT 487.950 322.950 490.050 323.400 ;
        RECT 526.950 321.600 529.050 323.700 ;
        RECT 547.950 322.500 550.050 324.600 ;
        RECT 562.950 322.500 565.050 324.600 ;
        RECT 583.950 323.700 585.150 327.300 ;
        RECT 661.950 324.450 664.050 325.050 ;
        RECT 712.950 324.450 715.050 325.050 ;
        RECT 734.700 324.600 735.900 344.400 ;
        RECT 739.950 335.250 742.050 337.050 ;
        RECT 739.950 333.450 742.050 334.050 ;
        RECT 748.950 333.450 751.050 334.050 ;
        RECT 739.950 332.400 751.050 333.450 ;
        RECT 739.950 331.950 742.050 332.400 ;
        RECT 748.950 331.950 751.050 332.400 ;
        RECT 754.950 329.400 756.150 344.400 ;
        RECT 760.950 343.950 763.050 344.400 ;
        RECT 778.950 343.950 781.050 344.400 ;
        RECT 806.400 344.400 814.050 345.450 ;
        RECT 793.950 340.950 796.050 343.050 ;
        RECT 799.950 342.450 802.050 343.050 ;
        RECT 806.400 342.450 807.450 344.400 ;
        RECT 811.950 343.950 814.050 344.400 ;
        RECT 859.950 345.450 862.050 346.050 ;
        RECT 880.950 345.450 883.050 346.050 ;
        RECT 859.950 344.400 883.050 345.450 ;
        RECT 859.950 343.950 862.050 344.400 ;
        RECT 880.950 343.950 883.050 344.400 ;
        RECT 886.950 345.450 889.050 346.050 ;
        RECT 892.950 345.450 895.050 346.050 ;
        RECT 886.950 344.400 895.050 345.450 ;
        RECT 886.950 343.950 889.050 344.400 ;
        RECT 892.950 343.950 895.050 344.400 ;
        RECT 799.950 341.400 807.450 342.450 ;
        RECT 799.950 340.950 802.050 341.400 ;
        RECT 757.950 337.950 760.050 340.050 ;
        RECT 766.950 339.450 771.000 340.050 ;
        RECT 772.950 339.450 775.050 340.050 ;
        RECT 787.950 339.450 790.050 340.050 ;
        RECT 766.950 338.400 790.050 339.450 ;
        RECT 766.950 337.950 771.000 338.400 ;
        RECT 772.950 337.950 775.050 338.400 ;
        RECT 787.950 337.950 790.050 338.400 ;
        RECT 793.950 337.950 796.050 339.750 ;
        RECT 799.950 337.950 802.050 339.750 ;
        RECT 811.950 337.950 814.050 340.050 ;
        RECT 835.950 339.450 838.050 340.050 ;
        RECT 844.950 339.450 847.050 340.050 ;
        RECT 835.950 338.400 847.050 339.450 ;
        RECT 835.950 337.950 838.050 338.400 ;
        RECT 844.950 337.950 847.050 338.400 ;
        RECT 850.950 337.950 853.050 340.050 ;
        RECT 871.950 337.950 874.050 340.050 ;
        RECT 877.950 337.950 880.050 343.050 ;
        RECT 883.950 337.950 886.050 340.050 ;
        RECT 889.950 339.450 892.050 340.050 ;
        RECT 898.950 339.450 904.050 340.050 ;
        RECT 889.950 338.400 904.050 339.450 ;
        RECT 889.950 337.950 892.050 338.400 ;
        RECT 898.950 337.950 904.050 338.400 ;
        RECT 757.950 334.950 760.050 336.750 ;
        RECT 772.950 334.950 775.050 336.750 ;
        RECT 778.950 336.450 781.050 337.050 ;
        RECT 790.950 336.450 793.050 337.050 ;
        RECT 778.950 335.400 793.050 336.450 ;
        RECT 778.950 334.950 781.050 335.400 ;
        RECT 790.950 334.950 793.050 335.400 ;
        RECT 796.950 335.250 799.050 337.050 ;
        RECT 811.950 334.950 814.050 336.750 ;
        RECT 835.950 334.950 838.050 336.750 ;
        RECT 850.950 334.950 853.050 336.750 ;
        RECT 871.950 334.950 874.050 336.750 ;
        RECT 877.950 334.950 880.050 336.750 ;
        RECT 883.950 334.950 886.050 336.750 ;
        RECT 901.950 334.950 904.050 336.750 ;
        RECT 775.950 332.250 778.050 334.050 ;
        RECT 796.950 333.450 799.050 334.050 ;
        RECT 801.000 333.450 805.050 334.050 ;
        RECT 796.950 332.400 805.050 333.450 ;
        RECT 796.950 331.950 799.050 332.400 ;
        RECT 801.000 331.950 805.050 332.400 ;
        RECT 814.950 332.250 817.050 334.050 ;
        RECT 832.950 332.250 835.050 334.050 ;
        RECT 838.950 332.250 841.050 334.050 ;
        RECT 853.950 332.250 856.050 334.050 ;
        RECT 874.950 332.250 877.050 334.050 ;
        RECT 880.950 332.250 883.050 334.050 ;
        RECT 898.950 332.250 901.050 334.050 ;
        RECT 754.950 327.300 757.050 329.400 ;
        RECT 775.950 328.950 781.050 331.050 ;
        RECT 814.950 328.950 817.050 331.050 ;
        RECT 832.950 328.950 835.050 331.050 ;
        RECT 838.950 328.950 841.050 331.050 ;
        RECT 853.950 330.450 856.050 331.050 ;
        RECT 868.950 330.450 871.050 331.050 ;
        RECT 853.950 329.400 871.050 330.450 ;
        RECT 853.950 328.950 856.050 329.400 ;
        RECT 868.950 328.950 871.050 329.400 ;
        RECT 874.950 328.950 877.050 331.050 ;
        RECT 880.950 328.950 883.050 331.050 ;
        RECT 886.950 330.450 889.050 331.050 ;
        RECT 898.950 330.450 901.050 331.050 ;
        RECT 886.950 329.400 901.050 330.450 ;
        RECT 886.950 328.950 889.050 329.400 ;
        RECT 898.950 328.950 901.050 329.400 ;
        RECT 583.950 321.600 586.050 323.700 ;
        RECT 661.950 323.400 715.050 324.450 ;
        RECT 661.950 322.950 664.050 323.400 ;
        RECT 712.950 322.950 715.050 323.400 ;
        RECT 733.950 322.500 736.050 324.600 ;
        RECT 754.950 323.700 756.150 327.300 ;
        RECT 776.400 324.450 777.450 328.950 ;
        RECT 802.950 324.450 805.050 325.050 ;
        RECT 697.950 321.450 700.050 322.050 ;
        RECT 718.950 321.450 721.050 322.050 ;
        RECT 754.950 321.600 757.050 323.700 ;
        RECT 776.400 323.400 805.050 324.450 ;
        RECT 802.950 322.950 805.050 323.400 ;
        RECT 808.950 324.450 811.050 325.050 ;
        RECT 814.950 324.450 817.050 325.050 ;
        RECT 808.950 323.400 817.050 324.450 ;
        RECT 808.950 322.950 811.050 323.400 ;
        RECT 814.950 322.950 817.050 323.400 ;
        RECT 880.950 324.450 883.050 325.050 ;
        RECT 895.950 324.450 898.050 325.050 ;
        RECT 880.950 323.400 898.050 324.450 ;
        RECT 880.950 322.950 883.050 323.400 ;
        RECT 895.950 322.950 898.050 323.400 ;
        RECT 697.950 320.400 721.050 321.450 ;
        RECT 697.950 319.950 700.050 320.400 ;
        RECT 718.950 319.950 721.050 320.400 ;
        RECT 109.950 318.450 112.050 319.050 ;
        RECT 169.950 318.450 172.050 319.050 ;
        RECT 109.950 317.400 172.050 318.450 ;
        RECT 109.950 316.950 112.050 317.400 ;
        RECT 169.950 316.950 172.050 317.400 ;
        RECT 178.950 318.450 181.050 319.050 ;
        RECT 184.950 318.450 187.050 319.050 ;
        RECT 178.950 317.400 187.050 318.450 ;
        RECT 178.950 316.950 181.050 317.400 ;
        RECT 184.950 316.950 187.050 317.400 ;
        RECT 310.950 318.450 313.050 319.050 ;
        RECT 319.950 318.450 322.050 319.050 ;
        RECT 487.950 318.450 490.050 319.050 ;
        RECT 310.950 317.400 490.050 318.450 ;
        RECT 310.950 316.950 313.050 317.400 ;
        RECT 319.950 316.950 322.050 317.400 ;
        RECT 487.950 316.950 490.050 317.400 ;
        RECT 508.950 318.450 511.050 319.050 ;
        RECT 724.950 318.450 727.050 319.050 ;
        RECT 508.950 317.400 727.050 318.450 ;
        RECT 508.950 316.950 511.050 317.400 ;
        RECT 724.950 316.950 727.050 317.400 ;
        RECT 748.950 318.450 751.050 319.050 ;
        RECT 778.950 318.450 781.050 319.050 ;
        RECT 748.950 317.400 781.050 318.450 ;
        RECT 748.950 316.950 751.050 317.400 ;
        RECT 778.950 316.950 781.050 317.400 ;
        RECT 880.950 318.450 883.050 319.050 ;
        RECT 889.950 318.450 892.050 319.050 ;
        RECT 880.950 317.400 892.050 318.450 ;
        RECT 880.950 316.950 883.050 317.400 ;
        RECT 889.950 316.950 892.050 317.400 ;
        RECT 145.950 315.450 148.050 316.050 ;
        RECT 181.950 315.450 184.050 316.050 ;
        RECT 145.950 314.400 184.050 315.450 ;
        RECT 145.950 313.950 148.050 314.400 ;
        RECT 181.950 313.950 184.050 314.400 ;
        RECT 211.950 315.450 214.050 316.050 ;
        RECT 229.950 315.450 232.050 316.050 ;
        RECT 211.950 314.400 232.050 315.450 ;
        RECT 211.950 313.950 214.050 314.400 ;
        RECT 229.950 313.950 232.050 314.400 ;
        RECT 466.950 315.450 469.050 316.050 ;
        RECT 523.950 315.450 526.050 316.050 ;
        RECT 466.950 314.400 526.050 315.450 ;
        RECT 466.950 313.950 469.050 314.400 ;
        RECT 523.950 313.950 526.050 314.400 ;
        RECT 559.950 315.450 562.050 316.050 ;
        RECT 625.950 315.450 628.050 316.050 ;
        RECT 634.950 315.450 637.050 316.050 ;
        RECT 709.950 315.450 712.050 316.050 ;
        RECT 730.950 315.450 733.050 316.050 ;
        RECT 739.950 315.450 742.050 316.050 ;
        RECT 820.950 315.450 823.050 316.050 ;
        RECT 865.950 315.450 868.050 316.050 ;
        RECT 871.950 315.450 874.050 316.050 ;
        RECT 559.950 314.400 874.050 315.450 ;
        RECT 559.950 313.950 562.050 314.400 ;
        RECT 625.950 313.950 628.050 314.400 ;
        RECT 634.950 313.950 637.050 314.400 ;
        RECT 709.950 313.950 712.050 314.400 ;
        RECT 730.950 313.950 733.050 314.400 ;
        RECT 739.950 313.950 742.050 314.400 ;
        RECT 820.950 313.950 823.050 314.400 ;
        RECT 865.950 313.950 868.050 314.400 ;
        RECT 871.950 313.950 874.050 314.400 ;
        RECT 76.950 312.450 79.050 313.050 ;
        RECT 100.950 312.450 103.050 313.050 ;
        RECT 76.950 311.400 103.050 312.450 ;
        RECT 76.950 310.950 79.050 311.400 ;
        RECT 100.950 310.950 103.050 311.400 ;
        RECT 163.950 312.450 166.050 313.050 ;
        RECT 232.950 312.450 235.050 313.050 ;
        RECT 163.950 311.400 235.050 312.450 ;
        RECT 163.950 310.950 166.050 311.400 ;
        RECT 232.950 310.950 235.050 311.400 ;
        RECT 241.950 312.450 244.050 313.050 ;
        RECT 316.950 312.450 319.050 313.050 ;
        RECT 241.950 311.400 319.050 312.450 ;
        RECT 241.950 310.950 244.050 311.400 ;
        RECT 316.950 310.950 319.050 311.400 ;
        RECT 394.950 312.450 397.050 313.050 ;
        RECT 472.950 312.450 475.050 313.050 ;
        RECT 577.950 312.450 580.050 313.050 ;
        RECT 394.950 311.400 580.050 312.450 ;
        RECT 394.950 310.950 397.050 311.400 ;
        RECT 472.950 310.950 475.050 311.400 ;
        RECT 577.950 310.950 580.050 311.400 ;
        RECT 34.950 309.450 37.050 310.050 ;
        RECT 64.950 309.450 67.050 310.050 ;
        RECT 103.950 309.450 106.050 310.050 ;
        RECT 34.950 308.400 106.050 309.450 ;
        RECT 34.950 307.950 37.050 308.400 ;
        RECT 64.950 307.950 67.050 308.400 ;
        RECT 103.950 307.950 106.050 308.400 ;
        RECT 172.950 309.450 175.050 310.050 ;
        RECT 199.950 309.450 202.050 310.050 ;
        RECT 220.950 309.450 223.050 310.050 ;
        RECT 172.950 308.400 223.050 309.450 ;
        RECT 172.950 307.950 175.050 308.400 ;
        RECT 199.950 307.950 202.050 308.400 ;
        RECT 220.950 307.950 223.050 308.400 ;
        RECT 340.950 309.450 343.050 310.050 ;
        RECT 406.950 309.450 409.050 310.050 ;
        RECT 340.950 308.400 409.050 309.450 ;
        RECT 340.950 307.950 343.050 308.400 ;
        RECT 406.950 307.950 409.050 308.400 ;
        RECT 442.950 309.450 445.050 310.050 ;
        RECT 496.950 309.450 499.050 310.050 ;
        RECT 502.950 309.450 505.050 310.050 ;
        RECT 535.950 309.450 538.050 310.050 ;
        RECT 553.950 309.450 556.050 310.050 ;
        RECT 442.950 308.400 556.050 309.450 ;
        RECT 442.950 307.950 445.050 308.400 ;
        RECT 496.950 307.950 499.050 308.400 ;
        RECT 502.950 307.950 505.050 308.400 ;
        RECT 535.950 307.950 538.050 308.400 ;
        RECT 553.950 307.950 556.050 308.400 ;
        RECT 721.950 309.450 724.050 310.050 ;
        RECT 784.950 309.450 787.050 310.050 ;
        RECT 721.950 308.400 787.050 309.450 ;
        RECT 721.950 307.950 724.050 308.400 ;
        RECT 784.950 307.950 787.050 308.400 ;
        RECT 814.950 309.450 817.050 310.050 ;
        RECT 826.950 309.450 829.050 310.050 ;
        RECT 892.950 309.450 895.050 310.050 ;
        RECT 814.950 308.400 895.050 309.450 ;
        RECT 814.950 307.950 817.050 308.400 ;
        RECT 826.950 307.950 829.050 308.400 ;
        RECT 892.950 307.950 895.050 308.400 ;
        RECT 28.950 306.450 31.050 307.050 ;
        RECT 127.950 306.450 130.050 307.050 ;
        RECT 28.950 305.400 130.050 306.450 ;
        RECT 196.950 306.450 199.050 307.050 ;
        RECT 211.950 306.450 214.050 307.050 ;
        RECT 196.950 305.400 214.050 306.450 ;
        RECT 349.950 306.450 352.050 307.050 ;
        RECT 373.950 306.450 376.050 307.050 ;
        RECT 349.950 305.400 376.050 306.450 ;
        RECT 28.950 304.950 31.050 305.400 ;
        RECT 127.950 304.950 130.050 305.400 ;
        RECT 43.950 303.450 46.050 304.050 ;
        RECT 43.950 302.400 84.450 303.450 ;
        RECT 157.950 303.300 160.050 305.400 ;
        RECT 196.950 304.950 199.050 305.400 ;
        RECT 211.950 304.950 214.050 305.400 ;
        RECT 43.950 301.950 46.050 302.400 ;
        RECT 83.400 298.050 84.450 302.400 ;
        RECT 158.850 299.700 160.050 303.300 ;
        RECT 178.950 302.400 181.050 304.500 ;
        RECT 193.950 303.450 196.050 304.050 ;
        RECT 205.950 303.450 208.050 304.050 ;
        RECT 193.950 302.400 208.050 303.450 ;
        RECT 259.950 303.300 262.050 305.400 ;
        RECT 349.950 304.950 352.050 305.400 ;
        RECT 373.950 304.950 376.050 305.400 ;
        RECT 37.950 295.950 40.050 298.050 ;
        RECT 43.950 295.950 46.050 298.050 ;
        RECT 58.950 295.950 61.050 298.050 ;
        RECT 64.950 295.950 67.050 298.050 ;
        RECT 82.950 295.950 85.050 298.050 ;
        RECT 100.950 295.950 103.050 298.050 ;
        RECT 106.950 295.950 109.050 298.050 ;
        RECT 121.950 295.950 124.050 298.050 ;
        RECT 127.950 295.950 130.050 298.050 ;
        RECT 145.950 295.950 148.050 298.050 ;
        RECT 157.950 297.600 160.050 299.700 ;
        RECT 16.950 292.950 19.050 295.050 ;
        RECT 37.950 292.950 40.050 294.750 ;
        RECT 43.950 292.950 46.050 294.750 ;
        RECT 58.950 292.950 61.050 294.750 ;
        RECT 64.950 292.950 67.050 294.750 ;
        RECT 82.950 292.950 85.050 294.750 ;
        RECT 100.950 292.950 103.050 294.750 ;
        RECT 106.950 292.950 109.050 294.750 ;
        RECT 121.950 292.950 124.050 294.750 ;
        RECT 127.950 292.950 130.050 294.750 ;
        RECT 145.950 292.950 148.050 294.750 ;
        RECT 16.950 289.950 19.050 291.750 ;
        RECT 34.950 290.250 37.050 292.050 ;
        RECT 40.950 290.250 43.050 292.050 ;
        RECT 61.950 290.250 64.050 292.050 ;
        RECT 67.950 290.250 70.050 292.050 ;
        RECT 85.950 290.250 88.050 292.050 ;
        RECT 97.950 290.250 100.050 292.050 ;
        RECT 103.950 290.250 106.050 292.050 ;
        RECT 124.950 290.250 127.050 292.050 ;
        RECT 142.950 290.250 145.050 292.050 ;
        RECT 154.950 290.250 157.050 292.050 ;
        RECT 13.950 287.250 16.050 289.050 ;
        RECT 19.950 287.250 22.050 289.050 ;
        RECT 28.950 288.450 33.000 289.050 ;
        RECT 34.950 288.450 37.050 289.050 ;
        RECT 28.950 287.400 37.050 288.450 ;
        RECT 28.950 286.950 33.000 287.400 ;
        RECT 34.950 286.950 37.050 287.400 ;
        RECT 40.950 286.950 43.050 289.050 ;
        RECT 46.950 288.450 49.050 289.050 ;
        RECT 61.950 288.450 64.050 289.050 ;
        RECT 46.950 287.400 64.050 288.450 ;
        RECT 46.950 286.950 49.050 287.400 ;
        RECT 61.950 286.950 64.050 287.400 ;
        RECT 67.950 286.950 70.050 289.050 ;
        RECT 73.950 288.450 76.050 289.050 ;
        RECT 85.950 288.450 88.050 289.050 ;
        RECT 90.000 288.450 94.050 289.050 ;
        RECT 73.950 287.400 94.050 288.450 ;
        RECT 73.950 286.950 76.050 287.400 ;
        RECT 85.950 286.950 88.050 287.400 ;
        RECT 90.000 286.950 94.050 287.400 ;
        RECT 97.950 286.950 100.050 289.050 ;
        RECT 103.950 288.450 106.050 289.050 ;
        RECT 118.950 288.450 121.050 289.050 ;
        RECT 103.950 287.400 121.050 288.450 ;
        RECT 103.950 286.950 106.050 287.400 ;
        RECT 118.950 286.950 121.050 287.400 ;
        RECT 124.950 288.450 127.050 289.050 ;
        RECT 136.950 288.450 139.050 289.050 ;
        RECT 124.950 287.400 139.050 288.450 ;
        RECT 124.950 286.950 127.050 287.400 ;
        RECT 136.950 286.950 139.050 287.400 ;
        RECT 142.950 286.950 145.050 289.050 ;
        RECT 154.950 286.950 157.050 289.050 ;
        RECT 13.950 283.950 16.050 286.050 ;
        RECT 19.950 283.950 25.050 286.050 ;
        RECT 43.950 285.450 46.050 286.050 ;
        RECT 52.950 285.450 55.050 286.050 ;
        RECT 43.950 284.400 55.050 285.450 ;
        RECT 43.950 283.950 46.050 284.400 ;
        RECT 52.950 283.950 55.050 284.400 ;
        RECT 112.950 282.450 115.050 283.050 ;
        RECT 142.950 282.450 145.050 283.050 ;
        RECT 151.950 282.450 154.050 283.050 ;
        RECT 158.850 282.600 160.050 297.600 ;
        RECT 172.950 292.950 175.050 295.050 ;
        RECT 172.950 289.950 175.050 291.750 ;
        RECT 179.100 282.600 180.300 302.400 ;
        RECT 193.950 301.950 196.050 302.400 ;
        RECT 205.950 301.950 208.050 302.400 ;
        RECT 181.950 300.450 184.050 301.050 ;
        RECT 196.950 300.450 199.050 301.050 ;
        RECT 181.950 299.400 199.050 300.450 ;
        RECT 260.850 299.700 262.050 303.300 ;
        RECT 280.950 302.400 283.050 304.500 ;
        RECT 355.950 303.450 358.050 304.050 ;
        RECT 367.950 303.450 370.050 304.050 ;
        RECT 355.950 302.400 370.050 303.450 ;
        RECT 382.950 302.400 385.050 304.500 ;
        RECT 403.950 303.300 406.050 305.400 ;
        RECT 418.950 303.300 421.050 305.400 ;
        RECT 181.950 298.950 184.050 299.400 ;
        RECT 196.950 298.950 199.050 299.400 ;
        RECT 187.950 297.450 190.050 298.050 ;
        RECT 199.950 297.450 202.050 298.050 ;
        RECT 187.950 296.400 202.050 297.450 ;
        RECT 187.950 295.950 190.050 296.400 ;
        RECT 199.950 295.950 202.050 296.400 ;
        RECT 205.950 295.950 208.050 298.050 ;
        RECT 220.950 295.950 223.050 298.050 ;
        RECT 226.950 295.950 229.050 298.050 ;
        RECT 259.950 297.600 262.050 299.700 ;
        RECT 265.950 300.450 268.050 301.050 ;
        RECT 274.950 300.450 277.050 301.050 ;
        RECT 265.950 299.400 277.050 300.450 ;
        RECT 265.950 298.950 268.050 299.400 ;
        RECT 274.950 298.950 277.050 299.400 ;
        RECT 181.950 292.950 184.050 295.050 ;
        RECT 199.950 292.950 202.050 294.750 ;
        RECT 205.950 292.950 208.050 294.750 ;
        RECT 220.950 292.950 223.050 294.750 ;
        RECT 226.950 292.950 229.050 294.750 ;
        RECT 247.950 294.450 250.050 295.050 ;
        RECT 252.000 294.450 256.050 295.050 ;
        RECT 247.950 293.400 256.050 294.450 ;
        RECT 247.950 292.950 250.050 293.400 ;
        RECT 252.000 292.950 256.050 293.400 ;
        RECT 181.950 289.950 184.050 291.750 ;
        RECT 196.950 290.250 199.050 292.050 ;
        RECT 202.950 290.250 205.050 292.050 ;
        RECT 223.950 290.250 226.050 292.050 ;
        RECT 247.950 289.950 250.050 291.750 ;
        RECT 256.950 290.250 259.050 292.050 ;
        RECT 184.950 288.450 187.050 289.050 ;
        RECT 196.950 288.450 199.050 289.050 ;
        RECT 184.950 287.400 199.050 288.450 ;
        RECT 184.950 286.950 187.050 287.400 ;
        RECT 196.950 286.950 199.050 287.400 ;
        RECT 202.950 283.950 205.050 289.050 ;
        RECT 223.950 288.450 226.050 289.050 ;
        RECT 232.950 288.450 235.050 289.050 ;
        RECT 223.950 287.400 235.050 288.450 ;
        RECT 223.950 286.950 226.050 287.400 ;
        RECT 232.950 286.950 235.050 287.400 ;
        RECT 244.950 287.250 247.050 289.050 ;
        RECT 250.950 287.250 253.050 289.050 ;
        RECT 256.950 286.950 259.050 289.050 ;
        RECT 229.950 285.450 232.050 286.050 ;
        RECT 244.950 285.450 247.050 286.050 ;
        RECT 229.950 284.400 247.050 285.450 ;
        RECT 229.950 283.950 232.050 284.400 ;
        RECT 244.950 283.950 247.050 284.400 ;
        RECT 250.950 283.950 253.050 286.050 ;
        RECT 260.850 282.600 262.050 297.600 ;
        RECT 274.950 292.950 277.050 295.050 ;
        RECT 274.950 289.950 277.050 291.750 ;
        RECT 281.100 282.600 282.300 302.400 ;
        RECT 355.950 301.950 358.050 302.400 ;
        RECT 367.950 301.950 370.050 302.400 ;
        RECT 283.950 300.450 286.050 301.050 ;
        RECT 298.950 300.450 301.050 301.050 ;
        RECT 283.950 299.400 301.050 300.450 ;
        RECT 283.950 298.950 286.050 299.400 ;
        RECT 298.950 298.950 301.050 299.400 ;
        RECT 304.950 295.950 307.050 298.050 ;
        RECT 310.950 295.950 313.050 298.050 ;
        RECT 361.950 295.950 364.050 298.050 ;
        RECT 367.950 295.950 370.050 298.050 ;
        RECT 283.950 292.950 286.050 295.050 ;
        RECT 304.950 292.950 307.050 294.750 ;
        RECT 310.950 292.950 313.050 294.750 ;
        RECT 316.950 294.450 319.050 295.050 ;
        RECT 325.950 294.450 328.050 295.050 ;
        RECT 316.950 293.400 328.050 294.450 ;
        RECT 316.950 292.950 319.050 293.400 ;
        RECT 325.950 292.950 328.050 293.400 ;
        RECT 361.950 292.950 364.050 294.750 ;
        RECT 367.950 292.950 370.050 294.750 ;
        RECT 379.950 292.950 382.050 295.050 ;
        RECT 283.950 289.950 286.050 291.750 ;
        RECT 301.950 290.250 304.050 292.050 ;
        RECT 307.950 290.250 310.050 292.050 ;
        RECT 325.950 289.950 328.050 291.750 ;
        RECT 346.950 289.950 349.050 291.750 ;
        RECT 364.950 290.250 367.050 292.050 ;
        RECT 370.950 290.250 373.050 292.050 ;
        RECT 379.950 289.950 382.050 291.750 ;
        RECT 295.950 288.450 300.000 289.050 ;
        RECT 301.950 288.450 304.050 289.050 ;
        RECT 295.950 287.400 304.050 288.450 ;
        RECT 295.950 286.950 300.000 287.400 ;
        RECT 301.950 286.950 304.050 287.400 ;
        RECT 307.950 286.950 310.050 289.050 ;
        RECT 364.950 286.950 367.050 289.050 ;
        RECT 283.950 285.450 288.000 286.050 ;
        RECT 313.950 285.450 316.050 286.050 ;
        RECT 352.950 285.450 355.050 286.050 ;
        RECT 358.950 285.450 361.050 286.050 ;
        RECT 283.950 283.950 288.450 285.450 ;
        RECT 313.950 284.400 361.050 285.450 ;
        RECT 313.950 283.950 316.050 284.400 ;
        RECT 352.950 283.950 355.050 284.400 ;
        RECT 358.950 283.950 361.050 284.400 ;
        RECT 370.950 283.950 373.050 289.050 ;
        RECT 112.950 281.400 154.050 282.450 ;
        RECT 112.950 280.950 115.050 281.400 ;
        RECT 142.950 280.950 145.050 281.400 ;
        RECT 151.950 280.950 154.050 281.400 ;
        RECT 157.950 280.500 160.050 282.600 ;
        RECT 178.950 280.500 181.050 282.600 ;
        RECT 259.950 280.500 262.050 282.600 ;
        RECT 280.950 280.500 283.050 282.600 ;
        RECT 287.400 282.450 288.450 283.950 ;
        RECT 355.950 282.450 358.050 283.050 ;
        RECT 383.700 282.600 384.900 302.400 ;
        RECT 403.950 299.700 405.150 303.300 ;
        RECT 419.850 299.700 421.050 303.300 ;
        RECT 439.950 302.400 442.050 304.500 ;
        RECT 472.950 303.300 475.050 305.400 ;
        RECT 403.950 297.600 406.050 299.700 ;
        RECT 418.950 297.600 421.050 299.700 ;
        RECT 388.950 292.950 391.050 295.050 ;
        RECT 388.950 289.950 391.050 291.750 ;
        RECT 403.950 282.600 405.150 297.600 ;
        RECT 406.950 290.250 409.050 292.050 ;
        RECT 415.950 290.250 418.050 292.050 ;
        RECT 406.950 286.950 409.050 289.050 ;
        RECT 415.950 286.950 418.050 289.050 ;
        RECT 419.850 282.600 421.050 297.600 ;
        RECT 433.950 292.950 436.050 295.050 ;
        RECT 433.950 289.950 436.050 291.750 ;
        RECT 440.100 282.600 441.300 302.400 ;
        RECT 473.850 299.700 475.050 303.300 ;
        RECT 493.950 302.400 496.050 304.500 ;
        RECT 529.950 303.300 532.050 305.400 ;
        RECT 448.950 297.450 451.050 298.050 ;
        RECT 460.950 297.450 463.050 298.050 ;
        RECT 472.950 297.600 475.050 299.700 ;
        RECT 448.950 296.400 463.050 297.450 ;
        RECT 448.950 295.950 451.050 296.400 ;
        RECT 460.950 295.950 463.050 296.400 ;
        RECT 442.950 292.950 445.050 295.050 ;
        RECT 460.950 292.950 463.050 294.750 ;
        RECT 442.950 289.950 445.050 291.750 ;
        RECT 463.950 290.250 466.050 292.050 ;
        RECT 469.950 290.250 472.050 292.050 ;
        RECT 460.950 286.950 466.050 289.050 ;
        RECT 469.950 283.950 472.050 289.050 ;
        RECT 287.400 281.400 358.050 282.450 ;
        RECT 355.950 280.950 358.050 281.400 ;
        RECT 382.950 280.500 385.050 282.600 ;
        RECT 403.950 280.500 406.050 282.600 ;
        RECT 418.950 280.500 421.050 282.600 ;
        RECT 439.950 280.500 442.050 282.600 ;
        RECT 451.950 282.450 454.050 283.050 ;
        RECT 466.950 282.450 469.050 283.050 ;
        RECT 473.850 282.600 475.050 297.600 ;
        RECT 487.950 292.950 490.050 295.050 ;
        RECT 487.950 289.950 490.050 291.750 ;
        RECT 494.100 282.600 495.300 302.400 ;
        RECT 530.850 299.700 532.050 303.300 ;
        RECT 550.950 302.400 553.050 304.500 ;
        RECT 628.950 302.400 631.050 304.500 ;
        RECT 649.950 303.300 652.050 305.400 ;
        RECT 685.950 303.300 688.050 305.400 ;
        RECT 511.950 295.950 514.050 298.050 ;
        RECT 517.950 295.950 520.050 298.050 ;
        RECT 529.950 297.600 532.050 299.700 ;
        RECT 496.950 292.950 499.050 295.050 ;
        RECT 511.950 292.950 514.050 294.750 ;
        RECT 517.950 292.950 520.050 294.750 ;
        RECT 496.950 289.950 499.050 291.750 ;
        RECT 514.950 290.250 517.050 292.050 ;
        RECT 526.950 290.250 529.050 292.050 ;
        RECT 514.950 283.950 517.050 289.050 ;
        RECT 526.950 286.950 529.050 289.050 ;
        RECT 530.850 282.600 532.050 297.600 ;
        RECT 538.950 294.450 543.000 295.050 ;
        RECT 544.950 294.450 547.050 295.050 ;
        RECT 538.950 293.400 547.050 294.450 ;
        RECT 538.950 292.950 543.000 293.400 ;
        RECT 544.950 292.950 547.050 293.400 ;
        RECT 544.950 289.950 547.050 291.750 ;
        RECT 551.100 282.600 552.300 302.400 ;
        RECT 553.950 300.450 556.050 301.050 ;
        RECT 553.950 299.400 573.450 300.450 ;
        RECT 553.950 298.950 556.050 299.400 ;
        RECT 572.400 295.050 573.450 299.400 ;
        RECT 610.950 295.950 613.050 298.050 ;
        RECT 616.950 295.950 619.050 298.050 ;
        RECT 553.950 292.950 556.050 295.050 ;
        RECT 571.950 292.950 574.050 295.050 ;
        RECT 610.950 292.950 613.050 294.750 ;
        RECT 616.950 292.950 619.050 294.750 ;
        RECT 625.950 292.950 628.050 295.050 ;
        RECT 553.950 289.950 556.050 291.750 ;
        RECT 571.950 289.950 574.050 291.750 ;
        RECT 592.950 289.950 595.050 291.750 ;
        RECT 607.950 290.250 610.050 292.050 ;
        RECT 613.950 290.250 616.050 292.050 ;
        RECT 625.950 289.950 628.050 291.750 ;
        RECT 607.950 286.950 610.050 289.050 ;
        RECT 613.950 288.450 616.050 289.050 ;
        RECT 622.950 288.450 625.050 289.050 ;
        RECT 613.950 287.400 625.050 288.450 ;
        RECT 613.950 286.950 616.050 287.400 ;
        RECT 622.950 286.950 625.050 287.400 ;
        RECT 629.700 282.600 630.900 302.400 ;
        RECT 649.950 299.700 651.150 303.300 ;
        RECT 686.850 299.700 688.050 303.300 ;
        RECT 706.950 302.400 709.050 304.500 ;
        RECT 742.950 302.400 745.050 304.500 ;
        RECT 763.950 303.300 766.050 305.400 ;
        RECT 790.950 303.450 793.050 304.050 ;
        RECT 808.950 303.450 811.050 304.050 ;
        RECT 649.950 297.600 652.050 299.700 ;
        RECT 634.950 292.950 637.050 295.050 ;
        RECT 634.950 289.950 637.050 291.750 ;
        RECT 649.950 282.600 651.150 297.600 ;
        RECT 655.950 297.450 658.050 298.050 ;
        RECT 667.950 297.450 670.050 298.050 ;
        RECT 655.950 296.400 670.050 297.450 ;
        RECT 655.950 295.950 658.050 296.400 ;
        RECT 667.950 295.950 670.050 296.400 ;
        RECT 673.950 295.950 676.050 298.050 ;
        RECT 685.950 297.600 688.050 299.700 ;
        RECT 691.950 300.450 694.050 301.050 ;
        RECT 700.950 300.450 703.050 301.050 ;
        RECT 691.950 299.400 703.050 300.450 ;
        RECT 691.950 298.950 694.050 299.400 ;
        RECT 700.950 298.950 703.050 299.400 ;
        RECT 667.950 292.950 670.050 294.750 ;
        RECT 673.950 292.950 676.050 294.750 ;
        RECT 652.950 290.250 655.050 292.050 ;
        RECT 670.950 290.250 673.050 292.050 ;
        RECT 682.950 290.250 685.050 292.050 ;
        RECT 652.950 286.950 655.050 289.050 ;
        RECT 664.950 288.450 669.000 289.050 ;
        RECT 670.950 288.450 673.050 289.050 ;
        RECT 664.950 287.400 673.050 288.450 ;
        RECT 664.950 286.950 669.000 287.400 ;
        RECT 670.950 286.950 673.050 287.400 ;
        RECT 682.950 286.950 685.050 289.050 ;
        RECT 686.850 282.600 688.050 297.600 ;
        RECT 700.950 292.950 703.050 295.050 ;
        RECT 700.950 289.950 703.050 291.750 ;
        RECT 707.100 282.600 708.300 302.400 ;
        RECT 724.950 295.950 727.050 298.050 ;
        RECT 730.950 295.950 733.050 298.050 ;
        RECT 709.950 292.950 712.050 295.050 ;
        RECT 724.950 292.950 727.050 294.750 ;
        RECT 730.950 292.950 733.050 294.750 ;
        RECT 739.950 292.950 742.050 295.050 ;
        RECT 709.950 289.950 712.050 291.750 ;
        RECT 727.950 290.250 730.050 292.050 ;
        RECT 739.950 289.950 742.050 291.750 ;
        RECT 721.950 288.450 726.000 289.050 ;
        RECT 727.950 288.450 730.050 289.050 ;
        RECT 721.950 287.400 730.050 288.450 ;
        RECT 721.950 286.950 726.000 287.400 ;
        RECT 727.950 286.950 730.050 287.400 ;
        RECT 743.700 282.600 744.900 302.400 ;
        RECT 763.950 299.700 765.150 303.300 ;
        RECT 790.950 302.400 811.050 303.450 ;
        RECT 823.950 302.400 826.050 304.500 ;
        RECT 844.950 303.300 847.050 305.400 ;
        RECT 790.950 301.950 793.050 302.400 ;
        RECT 808.950 301.950 811.050 302.400 ;
        RECT 763.950 297.600 766.050 299.700 ;
        RECT 748.950 292.950 751.050 295.050 ;
        RECT 748.950 289.950 751.050 291.750 ;
        RECT 763.950 282.600 765.150 297.600 ;
        RECT 784.950 295.950 787.050 298.050 ;
        RECT 790.950 295.950 793.050 298.050 ;
        RECT 784.950 292.950 787.050 294.750 ;
        RECT 790.950 292.950 793.050 294.750 ;
        RECT 811.950 292.950 817.050 295.050 ;
        RECT 820.950 292.950 823.050 295.050 ;
        RECT 766.950 290.250 769.050 292.050 ;
        RECT 787.950 290.250 790.050 292.050 ;
        RECT 793.950 290.250 796.050 292.050 ;
        RECT 811.950 289.950 814.050 291.750 ;
        RECT 820.950 289.950 823.050 291.750 ;
        RECT 766.950 286.950 769.050 289.050 ;
        RECT 787.950 286.950 790.050 289.050 ;
        RECT 793.950 286.950 796.050 289.050 ;
        RECT 808.950 287.250 811.050 289.050 ;
        RECT 814.950 287.250 817.050 289.050 ;
        RECT 808.950 283.950 811.050 286.050 ;
        RECT 814.950 283.950 817.050 286.050 ;
        RECT 451.950 281.400 469.050 282.450 ;
        RECT 451.950 280.950 454.050 281.400 ;
        RECT 466.950 280.950 469.050 281.400 ;
        RECT 472.950 280.500 475.050 282.600 ;
        RECT 493.950 280.500 496.050 282.600 ;
        RECT 529.950 280.500 532.050 282.600 ;
        RECT 550.950 280.500 553.050 282.600 ;
        RECT 628.950 280.500 631.050 282.600 ;
        RECT 649.950 280.500 652.050 282.600 ;
        RECT 685.950 280.500 688.050 282.600 ;
        RECT 706.950 280.500 709.050 282.600 ;
        RECT 742.950 280.500 745.050 282.600 ;
        RECT 763.950 280.500 766.050 282.600 ;
        RECT 778.950 282.450 781.050 283.050 ;
        RECT 787.950 282.450 790.050 283.050 ;
        RECT 824.700 282.600 825.900 302.400 ;
        RECT 844.950 299.700 846.150 303.300 ;
        RECT 844.950 297.600 847.050 299.700 ;
        RECT 829.950 292.950 832.050 295.050 ;
        RECT 829.950 289.950 832.050 291.750 ;
        RECT 844.950 282.600 846.150 297.600 ;
        RECT 871.950 294.450 874.050 295.050 ;
        RECT 886.950 294.450 889.050 295.050 ;
        RECT 871.950 293.400 889.050 294.450 ;
        RECT 871.950 292.950 874.050 293.400 ;
        RECT 886.950 292.950 889.050 293.400 ;
        RECT 847.950 290.250 850.050 292.050 ;
        RECT 865.950 289.950 868.050 291.750 ;
        RECT 886.950 289.950 889.050 291.750 ;
        RECT 847.950 286.950 850.050 289.050 ;
        RECT 778.950 281.400 790.050 282.450 ;
        RECT 778.950 280.950 781.050 281.400 ;
        RECT 787.950 280.950 790.050 281.400 ;
        RECT 823.950 280.500 826.050 282.600 ;
        RECT 844.950 280.500 847.050 282.600 ;
        RECT 208.950 277.950 214.050 280.050 ;
        RECT 241.950 279.450 244.050 280.050 ;
        RECT 250.950 279.450 253.050 280.050 ;
        RECT 241.950 278.400 253.050 279.450 ;
        RECT 241.950 277.950 244.050 278.400 ;
        RECT 250.950 277.950 253.050 278.400 ;
        RECT 286.950 279.450 289.050 280.050 ;
        RECT 316.950 279.450 319.050 280.050 ;
        RECT 376.950 279.450 379.050 280.050 ;
        RECT 286.950 278.400 379.050 279.450 ;
        RECT 286.950 277.950 289.050 278.400 ;
        RECT 316.950 277.950 319.050 278.400 ;
        RECT 376.950 277.950 379.050 278.400 ;
        RECT 517.950 279.450 520.050 280.050 ;
        RECT 523.950 279.450 526.050 280.050 ;
        RECT 517.950 278.400 526.050 279.450 ;
        RECT 517.950 277.950 520.050 278.400 ;
        RECT 523.950 277.950 526.050 278.400 ;
        RECT 802.950 279.450 805.050 280.050 ;
        RECT 808.950 279.450 811.050 280.050 ;
        RECT 802.950 278.400 811.050 279.450 ;
        RECT 802.950 277.950 805.050 278.400 ;
        RECT 808.950 277.950 811.050 278.400 ;
        RECT 55.950 276.450 58.050 277.050 ;
        RECT 145.950 276.450 148.050 277.050 ;
        RECT 184.950 276.450 187.050 277.050 ;
        RECT 202.950 276.450 205.050 277.050 ;
        RECT 55.950 275.400 187.050 276.450 ;
        RECT 55.950 274.950 58.050 275.400 ;
        RECT 145.950 274.950 148.050 275.400 ;
        RECT 184.950 274.950 187.050 275.400 ;
        RECT 188.400 275.400 205.050 276.450 ;
        RECT 79.950 273.450 82.050 274.050 ;
        RECT 23.400 272.400 82.050 273.450 ;
        RECT 23.400 271.050 24.450 272.400 ;
        RECT 79.950 271.950 82.050 272.400 ;
        RECT 136.950 273.450 139.050 274.050 ;
        RECT 148.950 273.450 151.050 274.050 ;
        RECT 136.950 272.400 151.050 273.450 ;
        RECT 136.950 271.950 139.050 272.400 ;
        RECT 148.950 271.950 151.050 272.400 ;
        RECT 172.950 273.450 175.050 274.050 ;
        RECT 188.400 273.450 189.450 275.400 ;
        RECT 202.950 274.950 205.050 275.400 ;
        RECT 265.950 276.450 268.050 277.050 ;
        RECT 292.950 276.450 295.050 277.050 ;
        RECT 265.950 275.400 295.050 276.450 ;
        RECT 265.950 274.950 268.050 275.400 ;
        RECT 292.950 274.950 295.050 275.400 ;
        RECT 340.950 276.450 343.050 277.050 ;
        RECT 364.950 276.450 367.050 277.050 ;
        RECT 391.950 276.450 394.050 277.050 ;
        RECT 415.950 276.450 418.050 277.050 ;
        RECT 340.950 275.400 390.450 276.450 ;
        RECT 340.950 274.950 343.050 275.400 ;
        RECT 364.950 274.950 367.050 275.400 ;
        RECT 172.950 272.400 189.450 273.450 ;
        RECT 199.950 273.450 202.050 274.050 ;
        RECT 286.950 273.450 289.050 274.050 ;
        RECT 199.950 272.400 289.050 273.450 ;
        RECT 172.950 271.950 175.050 272.400 ;
        RECT 199.950 271.950 202.050 272.400 ;
        RECT 286.950 271.950 289.050 272.400 ;
        RECT 307.950 273.450 310.050 274.050 ;
        RECT 319.950 273.450 322.050 274.050 ;
        RECT 307.950 272.400 322.050 273.450 ;
        RECT 307.950 271.950 310.050 272.400 ;
        RECT 319.950 271.950 322.050 272.400 ;
        RECT 370.950 273.450 373.050 274.050 ;
        RECT 385.950 273.450 388.050 274.050 ;
        RECT 370.950 272.400 388.050 273.450 ;
        RECT 389.400 273.450 390.450 275.400 ;
        RECT 391.950 275.400 418.050 276.450 ;
        RECT 391.950 274.950 394.050 275.400 ;
        RECT 415.950 274.950 418.050 275.400 ;
        RECT 481.950 276.450 484.050 277.050 ;
        RECT 490.950 276.450 493.050 277.050 ;
        RECT 481.950 275.400 493.050 276.450 ;
        RECT 481.950 274.950 484.050 275.400 ;
        RECT 490.950 274.950 493.050 275.400 ;
        RECT 502.950 276.450 505.050 277.050 ;
        RECT 520.950 276.450 523.050 277.050 ;
        RECT 607.950 276.450 610.050 277.050 ;
        RECT 502.950 275.400 523.050 276.450 ;
        RECT 502.950 274.950 505.050 275.400 ;
        RECT 520.950 274.950 523.050 275.400 ;
        RECT 530.400 275.400 610.050 276.450 ;
        RECT 433.950 273.450 436.050 274.050 ;
        RECT 530.400 273.450 531.450 275.400 ;
        RECT 607.950 274.950 610.050 275.400 ;
        RECT 655.950 276.450 658.050 277.050 ;
        RECT 730.950 276.450 733.050 277.050 ;
        RECT 655.950 275.400 733.050 276.450 ;
        RECT 655.950 274.950 658.050 275.400 ;
        RECT 730.950 274.950 733.050 275.400 ;
        RECT 742.950 276.450 745.050 277.050 ;
        RECT 766.950 276.450 769.050 277.050 ;
        RECT 742.950 275.400 769.050 276.450 ;
        RECT 742.950 274.950 745.050 275.400 ;
        RECT 766.950 274.950 769.050 275.400 ;
        RECT 841.950 276.450 844.050 277.050 ;
        RECT 847.950 276.450 850.050 277.050 ;
        RECT 868.950 276.450 871.050 277.050 ;
        RECT 841.950 275.400 871.050 276.450 ;
        RECT 841.950 274.950 844.050 275.400 ;
        RECT 847.950 274.950 850.050 275.400 ;
        RECT 868.950 274.950 871.050 275.400 ;
        RECT 538.950 273.450 541.050 274.050 ;
        RECT 389.400 272.400 531.450 273.450 ;
        RECT 533.400 272.400 541.050 273.450 ;
        RECT 370.950 271.950 373.050 272.400 ;
        RECT 385.950 271.950 388.050 272.400 ;
        RECT 433.950 271.950 436.050 272.400 ;
        RECT 22.950 270.450 25.050 271.050 ;
        RECT 28.950 270.450 31.050 271.050 ;
        RECT 22.950 269.400 31.050 270.450 ;
        RECT 22.950 268.950 25.050 269.400 ;
        RECT 28.950 268.950 31.050 269.400 ;
        RECT 85.950 270.450 88.050 271.050 ;
        RECT 97.950 270.450 100.050 271.050 ;
        RECT 85.950 269.400 100.050 270.450 ;
        RECT 85.950 268.950 88.050 269.400 ;
        RECT 97.950 268.950 100.050 269.400 ;
        RECT 250.950 270.450 253.050 271.050 ;
        RECT 259.950 270.450 262.050 271.050 ;
        RECT 250.950 269.400 262.050 270.450 ;
        RECT 250.950 268.950 253.050 269.400 ;
        RECT 259.950 268.950 262.050 269.400 ;
        RECT 274.950 270.450 277.050 271.050 ;
        RECT 283.950 270.450 286.050 271.050 ;
        RECT 274.950 269.400 286.050 270.450 ;
        RECT 274.950 268.950 277.050 269.400 ;
        RECT 283.950 268.950 286.050 269.400 ;
        RECT 382.950 270.450 385.050 271.050 ;
        RECT 430.950 270.450 433.050 271.050 ;
        RECT 382.950 269.400 433.050 270.450 ;
        RECT 382.950 268.950 385.050 269.400 ;
        RECT 430.950 268.950 433.050 269.400 ;
        RECT 439.950 270.450 442.050 271.050 ;
        RECT 448.950 270.450 451.050 271.050 ;
        RECT 439.950 269.400 451.050 270.450 ;
        RECT 439.950 268.950 442.050 269.400 ;
        RECT 448.950 268.950 451.050 269.400 ;
        RECT 505.950 270.450 508.050 271.050 ;
        RECT 514.950 270.450 517.050 271.050 ;
        RECT 505.950 269.400 517.050 270.450 ;
        RECT 505.950 268.950 508.050 269.400 ;
        RECT 514.950 268.950 517.050 269.400 ;
        RECT 520.950 270.450 523.050 271.050 ;
        RECT 533.400 270.450 534.450 272.400 ;
        RECT 538.950 271.950 541.050 272.400 ;
        RECT 544.950 273.450 547.050 274.050 ;
        RECT 583.950 273.450 586.050 274.050 ;
        RECT 544.950 272.400 586.050 273.450 ;
        RECT 544.950 271.950 547.050 272.400 ;
        RECT 583.950 271.950 586.050 272.400 ;
        RECT 616.950 273.450 619.050 274.050 ;
        RECT 664.950 273.450 667.050 274.050 ;
        RECT 616.950 272.400 667.050 273.450 ;
        RECT 616.950 271.950 619.050 272.400 ;
        RECT 664.950 271.950 667.050 272.400 ;
        RECT 793.950 273.450 796.050 274.050 ;
        RECT 823.950 273.450 826.050 274.050 ;
        RECT 895.950 273.450 898.050 274.050 ;
        RECT 793.950 272.400 898.050 273.450 ;
        RECT 793.950 271.950 796.050 272.400 ;
        RECT 823.950 271.950 826.050 272.400 ;
        RECT 895.950 271.950 898.050 272.400 ;
        RECT 520.950 269.400 534.450 270.450 ;
        RECT 604.950 270.450 607.050 271.050 ;
        RECT 622.950 270.450 625.050 271.050 ;
        RECT 604.950 269.400 625.050 270.450 ;
        RECT 520.950 268.950 523.050 269.400 ;
        RECT 604.950 268.950 607.050 269.400 ;
        RECT 622.950 268.950 625.050 269.400 ;
        RECT 628.950 270.450 631.050 271.050 ;
        RECT 640.950 270.450 643.050 271.050 ;
        RECT 652.950 270.450 655.050 271.050 ;
        RECT 628.950 269.400 655.050 270.450 ;
        RECT 628.950 268.950 631.050 269.400 ;
        RECT 640.950 268.950 643.050 269.400 ;
        RECT 652.950 268.950 655.050 269.400 ;
        RECT 670.950 270.450 673.050 271.050 ;
        RECT 715.950 270.450 718.050 271.050 ;
        RECT 670.950 269.400 718.050 270.450 ;
        RECT 670.950 268.950 673.050 269.400 ;
        RECT 715.950 268.950 718.050 269.400 ;
        RECT 859.950 270.450 862.050 271.050 ;
        RECT 886.950 270.450 889.050 271.050 ;
        RECT 859.950 269.400 889.050 270.450 ;
        RECT 859.950 268.950 862.050 269.400 ;
        RECT 886.950 268.950 889.050 269.400 ;
        RECT 13.950 262.950 16.050 268.050 ;
        RECT 46.950 266.400 49.050 268.500 ;
        RECT 67.950 266.400 70.050 268.500 ;
        RECT 91.950 267.450 94.050 268.050 ;
        RECT 80.400 266.400 94.050 267.450 ;
        RECT 19.950 264.450 22.050 265.050 ;
        RECT 31.950 264.450 34.050 265.050 ;
        RECT 19.950 263.400 34.050 264.450 ;
        RECT 19.950 262.950 22.050 263.400 ;
        RECT 31.950 262.950 34.050 263.400 ;
        RECT 13.950 259.950 16.050 261.750 ;
        RECT 19.950 259.950 22.050 261.750 ;
        RECT 37.950 259.950 40.050 262.050 ;
        RECT 43.950 259.950 46.050 262.050 ;
        RECT 16.950 257.250 19.050 259.050 ;
        RECT 37.950 256.950 40.050 258.750 ;
        RECT 43.950 256.950 46.050 258.750 ;
        RECT 16.950 255.450 19.050 256.050 ;
        RECT 21.000 255.450 25.050 256.050 ;
        RECT 16.950 254.400 25.050 255.450 ;
        RECT 16.950 253.950 19.050 254.400 ;
        RECT 21.000 253.950 25.050 254.400 ;
        RECT 34.950 254.250 37.050 256.050 ;
        RECT 34.950 250.950 37.050 253.050 ;
        RECT 47.850 251.400 49.050 266.400 ;
        RECT 61.950 257.250 64.050 259.050 ;
        RECT 61.950 253.950 64.050 256.050 ;
        RECT 46.950 249.300 49.050 251.400 ;
        RECT 28.950 246.450 31.050 247.050 ;
        RECT 34.950 246.450 37.050 247.050 ;
        RECT 28.950 245.400 37.050 246.450 ;
        RECT 47.850 245.700 49.050 249.300 ;
        RECT 68.100 246.600 69.300 266.400 ;
        RECT 70.950 264.450 73.050 265.050 ;
        RECT 80.400 264.450 81.450 266.400 ;
        RECT 91.950 265.950 94.050 266.400 ;
        RECT 70.950 263.400 81.450 264.450 ;
        RECT 70.950 262.950 73.050 263.400 ;
        RECT 112.950 262.950 115.050 268.050 ;
        RECT 145.950 266.400 148.050 268.500 ;
        RECT 166.950 266.400 169.050 268.500 ;
        RECT 172.950 267.450 175.050 268.050 ;
        RECT 199.950 267.450 202.050 268.050 ;
        RECT 172.950 266.400 202.050 267.450 ;
        RECT 118.950 264.450 121.050 265.050 ;
        RECT 130.950 264.450 133.050 265.050 ;
        RECT 118.950 263.400 133.050 264.450 ;
        RECT 118.950 262.950 121.050 263.400 ;
        RECT 130.950 262.950 133.050 263.400 ;
        RECT 85.950 259.950 88.050 262.050 ;
        RECT 91.950 259.950 94.050 262.050 ;
        RECT 112.950 259.950 115.050 261.750 ;
        RECT 118.950 259.950 121.050 261.750 ;
        RECT 136.950 259.950 139.050 262.050 ;
        RECT 142.950 259.950 145.050 262.050 ;
        RECT 70.950 257.250 73.050 259.050 ;
        RECT 85.950 256.950 88.050 258.750 ;
        RECT 91.950 256.950 94.050 258.750 ;
        RECT 115.950 257.250 118.050 259.050 ;
        RECT 136.950 256.950 139.050 258.750 ;
        RECT 142.950 256.950 145.050 258.750 ;
        RECT 70.950 253.950 73.050 256.050 ;
        RECT 88.950 254.250 91.050 256.050 ;
        RECT 94.950 254.250 97.050 256.050 ;
        RECT 100.950 255.450 103.050 256.050 ;
        RECT 115.950 255.450 118.050 256.050 ;
        RECT 100.950 254.400 118.050 255.450 ;
        RECT 100.950 253.950 103.050 254.400 ;
        RECT 115.950 253.950 118.050 254.400 ;
        RECT 133.950 254.250 136.050 256.050 ;
        RECT 88.950 250.950 91.050 253.050 ;
        RECT 94.950 250.950 97.050 253.050 ;
        RECT 133.950 250.950 136.050 253.050 ;
        RECT 146.850 251.400 148.050 266.400 ;
        RECT 160.950 257.250 163.050 259.050 ;
        RECT 145.950 249.300 148.050 251.400 ;
        RECT 160.950 250.950 163.050 256.050 ;
        RECT 28.950 244.950 31.050 245.400 ;
        RECT 34.950 244.950 37.050 245.400 ;
        RECT 46.950 243.600 49.050 245.700 ;
        RECT 67.950 244.500 70.050 246.600 ;
        RECT 79.950 246.450 82.050 247.050 ;
        RECT 88.950 246.450 91.050 247.050 ;
        RECT 79.950 245.400 91.050 246.450 ;
        RECT 146.850 245.700 148.050 249.300 ;
        RECT 167.100 246.600 168.300 266.400 ;
        RECT 172.950 265.950 175.050 266.400 ;
        RECT 199.950 265.950 202.050 266.400 ;
        RECT 229.950 267.450 232.050 268.050 ;
        RECT 280.950 267.450 283.050 268.050 ;
        RECT 229.950 266.400 283.050 267.450 ;
        RECT 289.950 266.400 292.050 268.500 ;
        RECT 310.950 266.400 313.050 268.500 ;
        RECT 388.950 267.450 391.050 268.050 ;
        RECT 394.950 267.450 397.050 268.050 ;
        RECT 478.950 267.450 481.050 268.050 ;
        RECT 526.950 267.450 529.050 268.050 ;
        RECT 388.950 266.400 397.050 267.450 ;
        RECT 229.950 265.950 232.050 266.400 ;
        RECT 280.950 265.950 283.050 266.400 ;
        RECT 184.950 259.950 187.050 262.050 ;
        RECT 190.950 259.950 193.050 262.050 ;
        RECT 196.950 261.450 199.050 262.050 ;
        RECT 208.950 261.450 211.050 262.050 ;
        RECT 196.950 260.400 211.050 261.450 ;
        RECT 196.950 259.950 199.050 260.400 ;
        RECT 208.950 259.950 211.050 260.400 ;
        RECT 220.950 261.450 223.050 262.050 ;
        RECT 232.950 261.450 235.050 262.050 ;
        RECT 220.950 260.400 235.050 261.450 ;
        RECT 220.950 259.950 223.050 260.400 ;
        RECT 232.950 259.950 235.050 260.400 ;
        RECT 241.950 261.450 244.050 262.050 ;
        RECT 250.950 261.450 253.050 262.050 ;
        RECT 241.950 260.400 253.050 261.450 ;
        RECT 241.950 259.950 244.050 260.400 ;
        RECT 250.950 259.950 253.050 260.400 ;
        RECT 271.950 259.950 277.050 262.050 ;
        RECT 280.950 259.950 283.050 262.050 ;
        RECT 286.950 259.950 289.050 262.050 ;
        RECT 169.950 257.250 172.050 259.050 ;
        RECT 184.950 256.950 187.050 258.750 ;
        RECT 190.950 256.950 193.050 258.750 ;
        RECT 208.950 256.950 211.050 258.750 ;
        RECT 232.950 256.950 235.050 258.750 ;
        RECT 250.950 256.950 253.050 258.750 ;
        RECT 274.950 256.950 277.050 258.750 ;
        RECT 280.950 256.950 283.050 258.750 ;
        RECT 286.950 256.950 289.050 258.750 ;
        RECT 169.950 253.950 172.050 256.050 ;
        RECT 187.950 254.250 190.050 256.050 ;
        RECT 193.950 254.250 196.050 256.050 ;
        RECT 211.950 254.250 214.050 256.050 ;
        RECT 229.950 254.250 232.050 256.050 ;
        RECT 235.950 254.250 238.050 256.050 ;
        RECT 247.950 254.250 250.050 256.050 ;
        RECT 253.950 254.250 256.050 256.050 ;
        RECT 271.950 254.250 274.050 256.050 ;
        RECT 277.950 254.250 280.050 256.050 ;
        RECT 187.950 250.950 190.050 253.050 ;
        RECT 193.950 250.950 199.050 253.050 ;
        RECT 211.950 252.450 214.050 253.050 ;
        RECT 216.000 252.450 220.050 253.050 ;
        RECT 211.950 251.400 220.050 252.450 ;
        RECT 211.950 250.950 214.050 251.400 ;
        RECT 216.000 250.950 220.050 251.400 ;
        RECT 229.950 250.950 232.050 253.050 ;
        RECT 235.950 252.450 238.050 253.050 ;
        RECT 240.000 252.450 244.050 253.050 ;
        RECT 235.950 251.400 244.050 252.450 ;
        RECT 235.950 250.950 238.050 251.400 ;
        RECT 240.000 250.950 244.050 251.400 ;
        RECT 247.950 250.950 250.050 253.050 ;
        RECT 253.950 250.950 256.050 253.050 ;
        RECT 271.950 250.950 274.050 253.050 ;
        RECT 277.950 250.950 280.050 253.050 ;
        RECT 290.850 251.400 292.050 266.400 ;
        RECT 304.950 257.250 307.050 259.050 ;
        RECT 304.950 253.950 307.050 256.050 ;
        RECT 169.950 249.450 172.050 250.050 ;
        RECT 169.950 248.400 186.450 249.450 ;
        RECT 169.950 247.950 172.050 248.400 ;
        RECT 79.950 244.950 82.050 245.400 ;
        RECT 88.950 244.950 91.050 245.400 ;
        RECT 145.950 243.600 148.050 245.700 ;
        RECT 166.950 244.500 169.050 246.600 ;
        RECT 185.400 246.450 186.450 248.400 ;
        RECT 193.800 246.450 195.900 247.050 ;
        RECT 185.400 245.400 195.900 246.450 ;
        RECT 193.800 244.950 195.900 245.400 ;
        RECT 197.100 246.450 199.200 247.050 ;
        RECT 241.950 246.450 244.050 247.050 ;
        RECT 197.100 245.400 244.050 246.450 ;
        RECT 197.100 244.950 199.200 245.400 ;
        RECT 241.950 244.950 244.050 245.400 ;
        RECT 253.950 246.450 256.050 247.050 ;
        RECT 272.400 246.450 273.450 250.950 ;
        RECT 289.950 249.300 292.050 251.400 ;
        RECT 283.950 246.450 286.050 247.050 ;
        RECT 253.950 245.400 286.050 246.450 ;
        RECT 290.850 245.700 292.050 249.300 ;
        RECT 311.100 246.600 312.300 266.400 ;
        RECT 388.950 265.950 391.050 266.400 ;
        RECT 394.950 265.950 397.050 266.400 ;
        RECT 473.400 266.400 529.050 267.450 ;
        RECT 538.950 266.400 541.050 268.500 ;
        RECT 559.950 266.400 562.050 268.500 ;
        RECT 667.950 267.450 670.050 268.050 ;
        RECT 700.950 267.450 703.050 268.050 ;
        RECT 748.950 267.450 751.050 268.050 ;
        RECT 667.950 266.400 703.050 267.450 ;
        RECT 319.950 261.450 322.050 262.050 ;
        RECT 334.950 261.450 337.050 262.050 ;
        RECT 319.950 260.400 337.050 261.450 ;
        RECT 319.950 259.950 322.050 260.400 ;
        RECT 334.950 259.950 337.050 260.400 ;
        RECT 340.950 259.950 343.050 262.050 ;
        RECT 352.950 259.950 355.050 262.050 ;
        RECT 358.950 261.450 361.050 262.050 ;
        RECT 376.950 261.450 379.050 262.050 ;
        RECT 358.950 260.400 379.050 261.450 ;
        RECT 358.950 259.950 361.050 260.400 ;
        RECT 376.950 259.950 379.050 260.400 ;
        RECT 382.950 259.950 385.050 265.050 ;
        RECT 439.950 262.950 442.050 265.050 ;
        RECT 445.950 264.450 448.050 265.050 ;
        RECT 454.950 264.450 457.050 265.050 ;
        RECT 445.950 263.400 457.050 264.450 ;
        RECT 445.950 262.950 448.050 263.400 ;
        RECT 454.950 262.950 457.050 263.400 ;
        RECT 460.950 262.950 463.050 265.050 ;
        RECT 466.950 264.450 469.050 265.050 ;
        RECT 473.400 264.450 474.450 266.400 ;
        RECT 478.950 265.950 481.050 266.400 ;
        RECT 526.950 265.950 529.050 266.400 ;
        RECT 466.950 263.400 474.450 264.450 ;
        RECT 466.950 262.950 469.050 263.400 ;
        RECT 388.950 259.950 391.050 262.050 ;
        RECT 421.950 259.950 424.050 262.050 ;
        RECT 439.950 259.950 442.050 261.750 ;
        RECT 445.950 259.950 448.050 261.750 ;
        RECT 460.950 259.950 463.050 261.750 ;
        RECT 466.950 259.950 469.050 261.750 ;
        RECT 478.950 259.950 481.050 262.050 ;
        RECT 496.950 259.950 499.050 262.050 ;
        RECT 502.950 259.950 505.050 262.050 ;
        RECT 511.950 261.450 514.050 262.050 ;
        RECT 520.950 261.450 523.050 262.050 ;
        RECT 511.950 260.400 523.050 261.450 ;
        RECT 511.950 259.950 514.050 260.400 ;
        RECT 520.950 259.950 523.050 260.400 ;
        RECT 313.950 257.250 316.050 259.050 ;
        RECT 334.950 256.950 337.050 258.750 ;
        RECT 340.950 256.950 343.050 258.750 ;
        RECT 352.950 256.950 355.050 258.750 ;
        RECT 358.950 256.950 361.050 258.750 ;
        RECT 382.950 256.950 385.050 258.750 ;
        RECT 388.950 256.950 391.050 258.750 ;
        RECT 400.950 256.950 403.050 258.750 ;
        RECT 421.950 256.950 424.050 258.750 ;
        RECT 442.950 257.250 445.050 259.050 ;
        RECT 463.950 257.250 466.050 259.050 ;
        RECT 478.950 256.950 481.050 258.750 ;
        RECT 496.950 256.950 499.050 258.750 ;
        RECT 502.950 256.950 505.050 258.750 ;
        RECT 508.950 256.950 514.050 259.050 ;
        RECT 520.950 256.950 523.050 258.750 ;
        RECT 526.950 257.250 529.050 259.050 ;
        RECT 535.950 257.250 538.050 259.050 ;
        RECT 313.950 253.950 316.050 256.050 ;
        RECT 331.950 254.250 334.050 256.050 ;
        RECT 337.950 254.250 340.050 256.050 ;
        RECT 355.950 254.250 358.050 256.050 ;
        RECT 361.950 254.250 364.050 256.050 ;
        RECT 379.950 254.250 382.050 256.050 ;
        RECT 385.950 254.250 388.050 256.050 ;
        RECT 403.950 254.250 406.050 256.050 ;
        RECT 424.950 254.250 427.050 256.050 ;
        RECT 430.950 255.450 433.050 256.050 ;
        RECT 442.950 255.450 445.050 256.050 ;
        RECT 430.950 254.400 445.050 255.450 ;
        RECT 430.950 253.950 433.050 254.400 ;
        RECT 442.950 253.950 445.050 254.400 ;
        RECT 448.950 255.450 451.050 256.050 ;
        RECT 463.950 255.450 466.050 256.050 ;
        RECT 448.950 254.400 466.050 255.450 ;
        RECT 448.950 253.950 451.050 254.400 ;
        RECT 463.950 253.950 466.050 254.400 ;
        RECT 481.950 254.250 484.050 256.050 ;
        RECT 499.950 254.250 502.050 256.050 ;
        RECT 505.950 254.250 508.050 256.050 ;
        RECT 526.950 253.950 532.050 256.050 ;
        RECT 535.950 253.950 538.050 256.050 ;
        RECT 331.950 250.950 334.050 253.050 ;
        RECT 337.950 250.950 340.050 253.050 ;
        RECT 355.950 247.950 358.050 253.050 ;
        RECT 361.950 250.950 364.050 253.050 ;
        RECT 379.950 250.950 382.050 253.050 ;
        RECT 385.950 250.950 388.050 253.050 ;
        RECT 394.950 252.450 397.050 253.050 ;
        RECT 403.950 252.450 406.050 253.050 ;
        RECT 394.950 251.400 406.050 252.450 ;
        RECT 394.950 250.950 397.050 251.400 ;
        RECT 403.950 250.950 406.050 251.400 ;
        RECT 424.950 250.950 427.050 253.050 ;
        RECT 481.950 252.450 484.050 253.050 ;
        RECT 493.950 252.450 496.050 253.050 ;
        RECT 481.950 251.400 496.050 252.450 ;
        RECT 481.950 250.950 484.050 251.400 ;
        RECT 493.950 250.950 496.050 251.400 ;
        RECT 499.950 250.950 502.050 253.050 ;
        RECT 505.950 250.950 508.050 253.050 ;
        RECT 362.400 247.050 363.450 250.950 ;
        RECT 511.950 249.450 514.050 250.050 ;
        RECT 529.950 249.450 532.050 250.050 ;
        RECT 511.950 248.400 532.050 249.450 ;
        RECT 511.950 247.950 514.050 248.400 ;
        RECT 529.950 247.950 532.050 248.400 ;
        RECT 253.950 244.950 256.050 245.400 ;
        RECT 283.950 244.950 286.050 245.400 ;
        RECT 178.950 243.450 181.050 244.050 ;
        RECT 196.950 243.450 199.050 244.050 ;
        RECT 178.950 242.400 199.050 243.450 ;
        RECT 178.950 241.950 181.050 242.400 ;
        RECT 196.950 241.950 199.050 242.400 ;
        RECT 259.950 243.450 262.050 244.050 ;
        RECT 274.950 243.450 277.050 244.050 ;
        RECT 289.950 243.600 292.050 245.700 ;
        RECT 310.950 244.500 313.050 246.600 ;
        RECT 358.950 246.450 363.450 247.050 ;
        RECT 391.950 246.450 394.050 247.050 ;
        RECT 358.950 245.400 394.050 246.450 ;
        RECT 358.950 244.950 363.000 245.400 ;
        RECT 391.950 244.950 394.050 245.400 ;
        RECT 415.950 246.450 418.050 247.050 ;
        RECT 493.950 246.450 496.050 247.050 ;
        RECT 415.950 245.400 496.050 246.450 ;
        RECT 415.950 244.950 418.050 245.400 ;
        RECT 493.950 244.950 496.050 245.400 ;
        RECT 505.950 246.450 508.050 247.050 ;
        RECT 514.950 246.450 517.050 247.050 ;
        RECT 539.700 246.600 540.900 266.400 ;
        RECT 544.950 257.250 547.050 259.050 ;
        RECT 544.950 253.950 547.050 256.050 ;
        RECT 559.950 251.400 561.150 266.400 ;
        RECT 667.950 265.950 670.050 266.400 ;
        RECT 700.950 265.950 703.050 266.400 ;
        RECT 707.400 266.400 751.050 267.450 ;
        RECT 562.950 259.950 565.050 262.050 ;
        RECT 577.950 259.950 580.050 262.050 ;
        RECT 583.950 259.950 586.050 265.050 ;
        RECT 622.950 262.950 625.050 265.050 ;
        RECT 628.950 262.950 631.050 265.050 ;
        RECT 682.950 262.050 685.050 265.050 ;
        RECT 707.400 262.050 708.450 266.400 ;
        RECT 748.950 265.950 751.050 266.400 ;
        RECT 793.950 267.450 796.050 268.050 ;
        RECT 802.950 267.450 805.050 268.050 ;
        RECT 793.950 266.400 805.050 267.450 ;
        RECT 793.950 265.950 796.050 266.400 ;
        RECT 802.950 265.950 805.050 266.400 ;
        RECT 817.950 267.450 820.050 268.050 ;
        RECT 829.950 267.450 832.050 268.050 ;
        RECT 817.950 266.400 832.050 267.450 ;
        RECT 817.950 265.950 820.050 266.400 ;
        RECT 829.950 265.950 832.050 266.400 ;
        RECT 847.950 264.450 852.000 265.050 ;
        RECT 853.950 264.450 856.050 265.050 ;
        RECT 847.950 263.400 856.050 264.450 ;
        RECT 847.950 262.950 852.000 263.400 ;
        RECT 853.950 262.950 856.050 263.400 ;
        RECT 859.950 262.950 862.050 265.050 ;
        RECT 868.950 264.450 873.000 265.050 ;
        RECT 874.950 264.450 877.050 265.050 ;
        RECT 868.950 263.400 877.050 264.450 ;
        RECT 868.950 262.950 873.000 263.400 ;
        RECT 874.950 262.950 877.050 263.400 ;
        RECT 880.950 262.950 883.050 265.050 ;
        RECT 589.950 261.450 592.050 262.050 ;
        RECT 604.950 261.450 607.050 262.050 ;
        RECT 589.950 260.400 607.050 261.450 ;
        RECT 589.950 259.950 592.050 260.400 ;
        RECT 604.950 259.950 607.050 260.400 ;
        RECT 622.950 259.950 625.050 261.750 ;
        RECT 628.950 259.950 631.050 261.750 ;
        RECT 679.950 259.950 685.050 262.050 ;
        RECT 700.950 259.950 703.050 262.050 ;
        RECT 706.950 259.950 709.050 262.050 ;
        RECT 715.950 261.450 718.050 262.050 ;
        RECT 730.950 261.450 733.050 262.050 ;
        RECT 715.950 260.400 733.050 261.450 ;
        RECT 715.950 259.950 718.050 260.400 ;
        RECT 730.950 259.950 733.050 260.400 ;
        RECT 751.950 261.450 754.050 262.050 ;
        RECT 763.950 261.450 766.050 262.050 ;
        RECT 751.950 260.400 766.050 261.450 ;
        RECT 751.950 259.950 754.050 260.400 ;
        RECT 763.950 259.950 766.050 260.400 ;
        RECT 772.950 261.450 775.050 262.050 ;
        RECT 781.950 261.450 784.050 262.050 ;
        RECT 772.950 260.400 784.050 261.450 ;
        RECT 772.950 259.950 775.050 260.400 ;
        RECT 781.950 259.950 784.050 260.400 ;
        RECT 787.950 259.950 790.050 262.050 ;
        RECT 793.950 259.950 796.050 262.050 ;
        RECT 817.950 259.950 820.050 262.050 ;
        RECT 823.950 259.950 826.050 262.050 ;
        RECT 841.950 259.950 844.050 262.050 ;
        RECT 853.950 259.950 856.050 261.750 ;
        RECT 859.950 259.950 862.050 261.750 ;
        RECT 874.950 259.950 877.050 261.750 ;
        RECT 880.950 259.950 883.050 261.750 ;
        RECT 895.950 259.950 898.050 262.050 ;
        RECT 562.950 256.950 565.050 258.750 ;
        RECT 577.950 256.950 580.050 258.750 ;
        RECT 583.950 256.950 586.050 258.750 ;
        RECT 604.950 256.950 607.050 258.750 ;
        RECT 625.950 257.250 628.050 259.050 ;
        RECT 646.950 257.250 649.050 259.050 ;
        RECT 667.950 257.250 670.050 259.050 ;
        RECT 682.950 256.950 685.050 258.750 ;
        RECT 700.950 256.950 703.050 258.750 ;
        RECT 706.950 256.950 709.050 258.750 ;
        RECT 730.950 256.950 733.050 258.750 ;
        RECT 751.950 256.950 754.050 258.750 ;
        RECT 772.950 256.950 775.050 258.750 ;
        RECT 787.950 256.950 790.050 258.750 ;
        RECT 793.950 256.950 796.050 258.750 ;
        RECT 817.950 256.950 820.050 258.750 ;
        RECT 823.950 256.950 826.050 258.750 ;
        RECT 841.950 256.950 844.050 258.750 ;
        RECT 856.950 257.250 859.050 259.050 ;
        RECT 877.950 257.250 880.050 259.050 ;
        RECT 895.950 256.950 898.050 258.750 ;
        RECT 901.950 257.250 904.050 259.050 ;
        RECT 580.950 254.250 583.050 256.050 ;
        RECT 586.950 254.250 589.050 256.050 ;
        RECT 601.950 254.250 604.050 256.050 ;
        RECT 607.950 254.250 610.050 256.050 ;
        RECT 619.950 255.450 624.000 256.050 ;
        RECT 625.950 255.450 628.050 256.050 ;
        RECT 619.950 254.400 628.050 255.450 ;
        RECT 619.950 253.950 624.000 254.400 ;
        RECT 625.950 253.950 628.050 254.400 ;
        RECT 667.950 255.450 670.050 256.050 ;
        RECT 679.950 255.450 682.050 256.050 ;
        RECT 667.950 254.400 682.050 255.450 ;
        RECT 667.950 253.950 670.050 254.400 ;
        RECT 679.950 253.950 682.050 254.400 ;
        RECT 685.950 254.250 688.050 256.050 ;
        RECT 703.950 254.250 706.050 256.050 ;
        RECT 709.950 254.250 712.050 256.050 ;
        RECT 727.950 254.250 730.050 256.050 ;
        RECT 733.950 254.250 736.050 256.050 ;
        RECT 748.950 254.250 751.050 256.050 ;
        RECT 754.950 254.250 757.050 256.050 ;
        RECT 769.950 254.250 772.050 256.050 ;
        RECT 775.950 254.250 778.050 256.050 ;
        RECT 790.950 254.250 793.050 256.050 ;
        RECT 796.950 254.250 799.050 256.050 ;
        RECT 814.950 254.250 817.050 256.050 ;
        RECT 820.950 254.250 823.050 256.050 ;
        RECT 838.950 254.250 841.050 256.050 ;
        RECT 856.950 255.450 859.050 256.050 ;
        RECT 865.950 255.450 868.050 256.050 ;
        RECT 856.950 254.400 868.050 255.450 ;
        RECT 856.950 253.950 859.050 254.400 ;
        RECT 865.950 253.950 868.050 254.400 ;
        RECT 871.950 255.450 876.000 256.050 ;
        RECT 877.950 255.450 880.050 256.050 ;
        RECT 871.950 254.400 880.050 255.450 ;
        RECT 871.950 253.950 876.000 254.400 ;
        RECT 877.950 253.950 880.050 254.400 ;
        RECT 559.950 249.300 562.050 251.400 ;
        RECT 580.950 250.950 583.050 253.050 ;
        RECT 586.950 250.950 589.050 253.050 ;
        RECT 601.950 250.950 604.050 253.050 ;
        RECT 607.950 250.950 610.050 253.050 ;
        RECT 685.950 252.450 691.050 253.050 ;
        RECT 697.950 252.450 700.050 253.050 ;
        RECT 685.950 251.400 700.050 252.450 ;
        RECT 685.950 250.950 691.050 251.400 ;
        RECT 697.950 250.950 700.050 251.400 ;
        RECT 703.950 250.950 706.050 253.050 ;
        RECT 709.950 250.950 712.050 253.050 ;
        RECT 727.950 250.950 730.050 253.050 ;
        RECT 733.950 252.450 736.050 253.050 ;
        RECT 742.950 252.450 745.050 253.050 ;
        RECT 733.950 251.400 745.050 252.450 ;
        RECT 733.950 250.950 736.050 251.400 ;
        RECT 742.950 250.950 745.050 251.400 ;
        RECT 748.950 250.950 751.050 253.050 ;
        RECT 754.950 250.950 757.050 253.050 ;
        RECT 769.950 250.950 772.050 253.050 ;
        RECT 775.950 252.450 778.050 253.050 ;
        RECT 784.950 252.450 787.050 253.050 ;
        RECT 775.950 251.400 787.050 252.450 ;
        RECT 775.950 250.950 778.050 251.400 ;
        RECT 784.950 250.950 787.050 251.400 ;
        RECT 790.950 250.950 793.050 253.050 ;
        RECT 796.950 250.950 799.050 253.050 ;
        RECT 814.950 250.950 817.050 253.050 ;
        RECT 820.950 250.950 823.050 253.050 ;
        RECT 826.950 252.450 829.050 253.050 ;
        RECT 838.950 252.450 841.050 253.050 ;
        RECT 826.950 251.400 841.050 252.450 ;
        RECT 826.950 250.950 829.050 251.400 ;
        RECT 838.950 250.950 841.050 251.400 ;
        RECT 505.950 245.400 517.050 246.450 ;
        RECT 505.950 244.950 508.050 245.400 ;
        RECT 514.950 244.950 517.050 245.400 ;
        RECT 538.950 244.500 541.050 246.600 ;
        RECT 559.950 245.700 561.150 249.300 ;
        RECT 565.950 246.450 568.050 247.050 ;
        RECT 602.400 246.450 603.450 250.950 ;
        RECT 259.950 242.400 277.050 243.450 ;
        RECT 259.950 241.950 262.050 242.400 ;
        RECT 274.950 241.950 277.050 242.400 ;
        RECT 337.950 243.450 340.050 244.050 ;
        RECT 343.950 243.450 346.050 244.050 ;
        RECT 385.950 243.450 388.050 244.050 ;
        RECT 409.950 243.450 412.050 244.050 ;
        RECT 337.950 242.400 388.050 243.450 ;
        RECT 337.950 241.950 340.050 242.400 ;
        RECT 343.950 241.950 346.050 242.400 ;
        RECT 385.950 241.950 388.050 242.400 ;
        RECT 389.400 242.400 412.050 243.450 ;
        RECT 121.950 240.450 124.050 241.050 ;
        RECT 199.950 240.450 202.050 241.050 ;
        RECT 121.950 239.400 202.050 240.450 ;
        RECT 121.950 238.950 124.050 239.400 ;
        RECT 199.950 238.950 202.050 239.400 ;
        RECT 262.950 240.450 265.050 241.050 ;
        RECT 277.950 240.450 280.050 241.050 ;
        RECT 292.950 240.450 295.050 241.050 ;
        RECT 262.950 239.400 295.050 240.450 ;
        RECT 262.950 238.950 265.050 239.400 ;
        RECT 277.950 238.950 280.050 239.400 ;
        RECT 292.950 238.950 295.050 239.400 ;
        RECT 304.950 240.450 307.050 241.050 ;
        RECT 319.950 240.450 322.050 241.050 ;
        RECT 304.950 239.400 322.050 240.450 ;
        RECT 304.950 238.950 307.050 239.400 ;
        RECT 319.950 238.950 322.050 239.400 ;
        RECT 325.950 240.450 328.050 241.050 ;
        RECT 389.400 240.450 390.450 242.400 ;
        RECT 409.950 241.950 412.050 242.400 ;
        RECT 424.950 243.450 427.050 244.050 ;
        RECT 451.800 243.450 453.900 244.050 ;
        RECT 424.950 242.400 453.900 243.450 ;
        RECT 424.950 241.950 427.050 242.400 ;
        RECT 451.800 241.950 453.900 242.400 ;
        RECT 455.100 243.450 457.200 244.050 ;
        RECT 481.950 243.450 484.050 244.050 ;
        RECT 455.100 242.400 484.050 243.450 ;
        RECT 455.100 241.950 457.200 242.400 ;
        RECT 481.950 241.950 484.050 242.400 ;
        RECT 514.950 241.950 520.050 244.050 ;
        RECT 559.950 243.600 562.050 245.700 ;
        RECT 565.950 245.400 675.450 246.450 ;
        RECT 565.950 244.950 568.050 245.400 ;
        RECT 674.400 243.450 675.450 245.400 ;
        RECT 712.950 244.950 718.050 247.050 ;
        RECT 781.950 246.450 784.050 247.050 ;
        RECT 796.950 246.450 799.050 247.050 ;
        RECT 781.950 245.400 799.050 246.450 ;
        RECT 781.950 244.950 784.050 245.400 ;
        RECT 796.950 244.950 799.050 245.400 ;
        RECT 802.950 246.450 805.050 247.050 ;
        RECT 823.950 246.450 826.050 247.050 ;
        RECT 802.950 245.400 826.050 246.450 ;
        RECT 802.950 244.950 805.050 245.400 ;
        RECT 823.950 244.950 826.050 245.400 ;
        RECT 838.950 246.450 841.050 247.050 ;
        RECT 847.950 246.450 850.050 247.050 ;
        RECT 838.950 245.400 850.050 246.450 ;
        RECT 838.950 244.950 841.050 245.400 ;
        RECT 847.950 244.950 850.050 245.400 ;
        RECT 712.950 243.450 715.050 244.050 ;
        RECT 674.400 242.400 715.050 243.450 ;
        RECT 712.950 241.950 715.050 242.400 ;
        RECT 718.950 243.450 721.050 244.050 ;
        RECT 748.950 243.450 751.050 244.050 ;
        RECT 718.950 242.400 751.050 243.450 ;
        RECT 718.950 241.950 721.050 242.400 ;
        RECT 748.950 241.950 751.050 242.400 ;
        RECT 763.950 243.450 766.050 244.050 ;
        RECT 814.950 243.450 817.050 244.050 ;
        RECT 763.950 242.400 817.050 243.450 ;
        RECT 763.950 241.950 766.050 242.400 ;
        RECT 814.950 241.950 817.050 242.400 ;
        RECT 325.950 239.400 390.450 240.450 ;
        RECT 394.950 240.450 397.050 241.050 ;
        RECT 421.950 240.450 424.050 241.050 ;
        RECT 394.950 239.400 424.050 240.450 ;
        RECT 325.950 238.950 328.050 239.400 ;
        RECT 394.950 238.950 397.050 239.400 ;
        RECT 421.950 238.950 424.050 239.400 ;
        RECT 427.950 240.450 430.050 241.050 ;
        RECT 448.950 240.450 451.050 241.050 ;
        RECT 427.950 239.400 451.050 240.450 ;
        RECT 452.400 240.450 453.450 241.950 ;
        RECT 460.950 240.450 463.050 241.050 ;
        RECT 452.400 239.400 463.050 240.450 ;
        RECT 427.950 238.950 430.050 239.400 ;
        RECT 448.950 238.950 451.050 239.400 ;
        RECT 460.950 238.950 463.050 239.400 ;
        RECT 484.950 240.450 487.050 241.050 ;
        RECT 580.950 240.450 583.050 241.050 ;
        RECT 607.950 240.450 610.050 241.050 ;
        RECT 673.950 240.450 676.050 241.050 ;
        RECT 484.950 239.400 579.450 240.450 ;
        RECT 484.950 238.050 487.050 239.400 ;
        RECT 28.950 237.450 31.050 238.050 ;
        RECT 70.950 237.450 73.050 238.050 ;
        RECT 28.950 236.400 73.050 237.450 ;
        RECT 28.950 235.950 31.050 236.400 ;
        RECT 70.950 235.950 73.050 236.400 ;
        RECT 94.950 237.450 97.050 238.050 ;
        RECT 220.950 237.450 223.050 238.050 ;
        RECT 94.950 236.400 223.050 237.450 ;
        RECT 94.950 235.950 97.050 236.400 ;
        RECT 220.950 235.950 223.050 236.400 ;
        RECT 286.950 237.450 289.050 238.050 ;
        RECT 307.950 237.450 310.050 238.050 ;
        RECT 286.950 236.400 310.050 237.450 ;
        RECT 286.950 235.950 289.050 236.400 ;
        RECT 307.950 235.950 310.050 236.400 ;
        RECT 481.950 237.000 487.050 238.050 ;
        RECT 578.400 237.450 579.450 239.400 ;
        RECT 580.950 239.400 676.050 240.450 ;
        RECT 580.950 238.950 583.050 239.400 ;
        RECT 607.950 238.950 610.050 239.400 ;
        RECT 673.950 238.950 676.050 239.400 ;
        RECT 679.950 240.450 682.050 241.050 ;
        RECT 754.950 240.450 757.050 241.050 ;
        RECT 775.950 240.450 778.050 241.050 ;
        RECT 679.950 239.400 711.450 240.450 ;
        RECT 679.950 238.950 682.050 239.400 ;
        RECT 661.950 237.450 664.050 238.050 ;
        RECT 481.950 236.400 486.450 237.000 ;
        RECT 578.400 236.400 664.050 237.450 ;
        RECT 710.400 237.450 711.450 239.400 ;
        RECT 754.950 239.400 778.050 240.450 ;
        RECT 754.950 238.950 757.050 239.400 ;
        RECT 775.950 238.950 778.050 239.400 ;
        RECT 784.950 237.450 787.050 238.050 ;
        RECT 802.950 237.450 805.050 238.050 ;
        RECT 710.400 236.400 805.050 237.450 ;
        RECT 481.950 235.950 486.000 236.400 ;
        RECT 661.950 235.950 664.050 236.400 ;
        RECT 784.950 235.950 787.050 236.400 ;
        RECT 802.950 235.950 805.050 236.400 ;
        RECT 64.950 234.450 67.050 235.050 ;
        RECT 133.950 234.450 136.050 235.050 ;
        RECT 187.950 234.450 190.050 235.050 ;
        RECT 64.950 233.400 190.050 234.450 ;
        RECT 64.950 232.950 67.050 233.400 ;
        RECT 133.950 232.950 136.050 233.400 ;
        RECT 187.950 232.950 190.050 233.400 ;
        RECT 271.950 234.450 274.050 235.050 ;
        RECT 331.950 234.450 334.050 235.050 ;
        RECT 415.950 234.450 418.050 235.050 ;
        RECT 475.950 234.450 478.050 235.050 ;
        RECT 505.950 234.450 508.050 235.050 ;
        RECT 271.950 233.400 334.050 234.450 ;
        RECT 271.950 232.950 274.050 233.400 ;
        RECT 331.950 232.950 334.050 233.400 ;
        RECT 335.400 233.400 418.050 234.450 ;
        RECT 85.950 231.450 88.050 232.050 ;
        RECT 100.950 231.450 103.050 232.050 ;
        RECT 85.950 230.400 103.050 231.450 ;
        RECT 85.950 229.950 88.050 230.400 ;
        RECT 100.950 229.950 103.050 230.400 ;
        RECT 109.950 231.450 112.050 232.050 ;
        RECT 139.950 231.450 142.050 232.050 ;
        RECT 109.950 230.400 142.050 231.450 ;
        RECT 109.950 229.950 112.050 230.400 ;
        RECT 139.950 229.950 142.050 230.400 ;
        RECT 190.950 231.450 193.050 232.050 ;
        RECT 232.950 231.450 235.050 232.050 ;
        RECT 190.950 230.400 235.050 231.450 ;
        RECT 190.950 229.950 193.050 230.400 ;
        RECT 232.950 229.950 235.050 230.400 ;
        RECT 250.950 231.450 253.050 232.050 ;
        RECT 313.950 231.450 316.050 232.050 ;
        RECT 335.400 231.450 336.450 233.400 ;
        RECT 415.950 232.950 418.050 233.400 ;
        RECT 452.400 233.400 478.050 234.450 ;
        RECT 250.950 230.400 336.450 231.450 ;
        RECT 361.950 231.450 364.050 232.050 ;
        RECT 421.950 231.450 424.050 232.050 ;
        RECT 430.950 231.450 433.050 232.050 ;
        RECT 361.950 230.400 399.450 231.450 ;
        RECT 250.950 229.950 253.050 230.400 ;
        RECT 313.950 229.950 316.050 230.400 ;
        RECT 361.950 229.950 364.050 230.400 ;
        RECT 40.950 228.450 43.050 229.050 ;
        RECT 55.950 228.450 58.050 229.050 ;
        RECT 40.950 227.400 58.050 228.450 ;
        RECT 265.950 228.450 268.050 229.050 ;
        RECT 280.950 228.450 283.050 229.050 ;
        RECT 265.950 227.400 283.050 228.450 ;
        RECT 40.950 226.950 43.050 227.400 ;
        RECT 55.950 226.950 58.050 227.400 ;
        RECT 13.950 225.450 16.050 226.050 ;
        RECT 37.950 225.450 40.050 226.050 ;
        RECT 70.950 225.450 73.050 226.050 ;
        RECT 13.950 224.400 73.050 225.450 ;
        RECT 94.950 225.300 97.050 227.400 ;
        RECT 13.950 223.950 16.050 224.400 ;
        RECT 37.950 223.950 40.050 224.400 ;
        RECT 70.950 223.950 73.050 224.400 ;
        RECT 49.950 222.450 52.050 223.050 ;
        RECT 64.950 222.450 67.050 223.050 ;
        RECT 49.950 221.400 67.050 222.450 ;
        RECT 95.850 221.700 97.050 225.300 ;
        RECT 115.950 224.400 118.050 226.500 ;
        RECT 175.950 225.300 178.050 227.400 ;
        RECT 265.950 226.950 268.050 227.400 ;
        RECT 280.950 226.950 283.050 227.400 ;
        RECT 298.950 228.450 301.050 229.050 ;
        RECT 325.950 228.450 328.050 229.050 ;
        RECT 298.950 227.400 328.050 228.450 ;
        RECT 398.400 228.450 399.450 230.400 ;
        RECT 421.950 230.400 433.050 231.450 ;
        RECT 421.950 229.950 424.050 230.400 ;
        RECT 430.950 229.950 433.050 230.400 ;
        RECT 442.950 231.450 445.050 232.050 ;
        RECT 452.400 231.450 453.450 233.400 ;
        RECT 475.950 232.950 478.050 233.400 ;
        RECT 479.400 233.400 508.050 234.450 ;
        RECT 442.950 230.400 453.450 231.450 ;
        RECT 454.950 231.450 457.050 232.050 ;
        RECT 479.400 231.450 480.450 233.400 ;
        RECT 505.950 232.950 508.050 233.400 ;
        RECT 559.950 234.450 562.050 235.050 ;
        RECT 613.950 234.450 616.050 235.050 ;
        RECT 688.950 234.450 691.050 235.050 ;
        RECT 559.950 233.400 691.050 234.450 ;
        RECT 803.400 234.450 804.450 235.950 ;
        RECT 841.950 234.450 844.050 235.050 ;
        RECT 803.400 233.400 844.050 234.450 ;
        RECT 559.950 232.950 562.050 233.400 ;
        RECT 613.950 232.950 616.050 233.400 ;
        RECT 688.950 232.950 691.050 233.400 ;
        RECT 841.950 232.950 844.050 233.400 ;
        RECT 454.950 230.400 480.450 231.450 ;
        RECT 493.950 231.450 496.050 232.050 ;
        RECT 523.950 231.450 526.050 232.050 ;
        RECT 667.800 231.450 669.900 232.050 ;
        RECT 493.950 230.400 669.900 231.450 ;
        RECT 442.950 229.950 445.050 230.400 ;
        RECT 454.950 229.950 457.050 230.400 ;
        RECT 493.950 229.950 496.050 230.400 ;
        RECT 523.950 229.950 526.050 230.400 ;
        RECT 667.800 229.950 669.900 230.400 ;
        RECT 671.100 231.450 673.200 232.050 ;
        RECT 703.950 231.450 706.050 232.050 ;
        RECT 721.950 231.450 724.050 232.050 ;
        RECT 727.950 231.450 730.050 232.050 ;
        RECT 742.950 231.450 745.050 232.050 ;
        RECT 671.100 230.400 745.050 231.450 ;
        RECT 671.100 229.950 673.200 230.400 ;
        RECT 703.950 229.950 706.050 230.400 ;
        RECT 721.950 229.950 724.050 230.400 ;
        RECT 727.950 229.950 730.050 230.400 ;
        RECT 742.950 229.950 745.050 230.400 ;
        RECT 760.950 231.450 763.050 232.050 ;
        RECT 859.950 231.450 862.050 232.050 ;
        RECT 760.950 230.400 862.050 231.450 ;
        RECT 760.950 229.950 763.050 230.400 ;
        RECT 859.950 229.950 862.050 230.400 ;
        RECT 865.950 231.450 868.050 232.050 ;
        RECT 883.950 231.450 886.050 232.050 ;
        RECT 865.950 230.400 886.050 231.450 ;
        RECT 865.950 229.950 868.050 230.400 ;
        RECT 883.950 229.950 886.050 230.400 ;
        RECT 421.950 228.450 424.050 229.050 ;
        RECT 398.400 227.400 424.050 228.450 ;
        RECT 511.950 228.450 514.050 229.050 ;
        RECT 547.950 228.450 550.050 229.050 ;
        RECT 511.950 227.400 550.050 228.450 ;
        RECT 661.950 228.450 664.050 229.050 ;
        RECT 715.950 228.450 718.050 229.050 ;
        RECT 661.950 227.400 718.050 228.450 ;
        RECT 298.950 226.950 301.050 227.400 ;
        RECT 325.950 226.950 328.050 227.400 ;
        RECT 49.950 220.950 52.050 221.400 ;
        RECT 64.950 220.950 67.050 221.400 ;
        RECT 13.950 217.950 16.050 220.050 ;
        RECT 19.950 217.950 22.050 220.050 ;
        RECT 34.950 217.950 37.050 220.050 ;
        RECT 40.950 217.950 43.050 220.050 ;
        RECT 94.950 219.600 97.050 221.700 ;
        RECT 13.950 214.950 16.050 216.750 ;
        RECT 19.950 214.950 22.050 216.750 ;
        RECT 34.950 214.950 37.050 216.750 ;
        RECT 40.950 214.950 43.050 216.750 ;
        RECT 61.950 216.450 64.050 217.050 ;
        RECT 70.950 216.450 73.050 217.050 ;
        RECT 82.950 216.450 85.050 217.050 ;
        RECT 61.950 215.400 69.450 216.450 ;
        RECT 61.950 214.950 64.050 215.400 ;
        RECT 16.950 212.250 19.050 214.050 ;
        RECT 37.950 212.250 40.050 214.050 ;
        RECT 43.950 212.250 46.050 214.050 ;
        RECT 61.950 211.950 64.050 213.750 ;
        RECT 68.400 213.450 69.450 215.400 ;
        RECT 70.950 215.400 85.050 216.450 ;
        RECT 70.950 214.950 73.050 215.400 ;
        RECT 82.950 214.950 85.050 215.400 ;
        RECT 76.950 213.450 79.050 214.050 ;
        RECT 68.400 212.400 79.050 213.450 ;
        RECT 76.950 211.950 79.050 212.400 ;
        RECT 82.950 211.950 85.050 213.750 ;
        RECT 91.950 212.250 94.050 214.050 ;
        RECT 16.950 210.450 19.050 211.050 ;
        RECT 31.950 210.450 34.050 211.050 ;
        RECT 16.950 209.400 34.050 210.450 ;
        RECT 16.950 208.950 19.050 209.400 ;
        RECT 31.950 208.950 34.050 209.400 ;
        RECT 37.950 205.950 40.050 211.050 ;
        RECT 43.950 208.950 46.050 211.050 ;
        RECT 58.950 209.250 61.050 211.050 ;
        RECT 64.950 209.250 67.050 211.050 ;
        RECT 79.950 209.250 82.050 211.050 ;
        RECT 85.950 209.250 88.050 211.050 ;
        RECT 91.950 208.950 94.050 211.050 ;
        RECT 58.950 205.950 61.050 208.050 ;
        RECT 64.950 205.950 67.050 208.050 ;
        RECT 79.950 205.950 82.050 208.050 ;
        RECT 85.950 205.950 88.050 208.050 ;
        RECT 43.950 204.450 46.050 205.050 ;
        RECT 49.950 204.450 52.050 205.050 ;
        RECT 95.850 204.600 97.050 219.600 ;
        RECT 109.950 214.950 112.050 220.050 ;
        RECT 109.950 211.950 112.050 213.750 ;
        RECT 116.100 204.600 117.300 224.400 ;
        RECT 124.950 222.450 127.050 223.050 ;
        RECT 133.950 222.450 136.050 223.050 ;
        RECT 124.950 221.400 136.050 222.450 ;
        RECT 176.850 221.700 178.050 225.300 ;
        RECT 196.950 224.400 199.050 226.500 ;
        RECT 247.950 225.450 250.050 226.050 ;
        RECT 316.950 225.450 319.050 226.050 ;
        RECT 336.000 225.450 340.050 226.050 ;
        RECT 247.950 224.400 340.050 225.450 ;
        RECT 124.950 220.950 127.050 221.400 ;
        RECT 133.950 220.950 136.050 221.400 ;
        RECT 136.950 217.950 139.050 220.050 ;
        RECT 142.950 217.950 145.050 220.050 ;
        RECT 157.950 217.950 160.050 220.050 ;
        RECT 163.950 217.950 166.050 220.050 ;
        RECT 175.950 219.600 178.050 221.700 ;
        RECT 118.950 214.950 121.050 217.050 ;
        RECT 136.950 214.950 139.050 216.750 ;
        RECT 142.950 214.950 145.050 216.750 ;
        RECT 157.950 214.950 160.050 216.750 ;
        RECT 163.950 214.950 166.050 216.750 ;
        RECT 118.950 211.950 121.050 213.750 ;
        RECT 133.950 212.250 136.050 214.050 ;
        RECT 139.950 212.250 142.050 214.050 ;
        RECT 160.950 212.250 163.050 214.050 ;
        RECT 172.950 212.250 175.050 214.050 ;
        RECT 133.950 208.950 136.050 211.050 ;
        RECT 139.950 208.950 142.050 211.050 ;
        RECT 145.950 210.450 148.050 211.050 ;
        RECT 160.950 210.450 163.050 211.050 ;
        RECT 145.950 209.400 163.050 210.450 ;
        RECT 145.950 208.950 148.050 209.400 ;
        RECT 160.950 208.950 163.050 209.400 ;
        RECT 172.950 208.950 175.050 211.050 ;
        RECT 43.950 203.400 52.050 204.450 ;
        RECT 43.950 202.950 46.050 203.400 ;
        RECT 49.950 202.950 52.050 203.400 ;
        RECT 94.950 202.500 97.050 204.600 ;
        RECT 115.950 202.500 118.050 204.600 ;
        RECT 133.950 204.450 136.050 205.050 ;
        RECT 157.950 204.450 160.050 205.050 ;
        RECT 176.850 204.600 178.050 219.600 ;
        RECT 190.950 214.950 193.050 217.050 ;
        RECT 190.950 211.950 193.050 213.750 ;
        RECT 197.100 204.600 198.300 224.400 ;
        RECT 247.950 223.950 250.050 224.400 ;
        RECT 316.950 223.950 319.050 224.400 ;
        RECT 335.400 223.950 340.050 224.400 ;
        RECT 346.950 225.450 349.050 226.050 ;
        RECT 352.950 225.450 355.050 226.050 ;
        RECT 346.950 224.400 355.050 225.450 ;
        RECT 364.950 225.300 367.050 227.400 ;
        RECT 421.950 226.950 424.050 227.400 ;
        RECT 346.950 223.950 349.050 224.400 ;
        RECT 352.950 223.950 355.050 224.400 ;
        RECT 262.950 222.450 267.000 223.050 ;
        RECT 283.950 222.450 286.050 223.050 ;
        RECT 304.950 222.450 307.050 223.050 ;
        RECT 262.950 220.950 268.050 222.450 ;
        RECT 283.950 221.400 307.050 222.450 ;
        RECT 283.950 220.950 286.050 221.400 ;
        RECT 304.950 220.950 307.050 221.400 ;
        RECT 205.950 219.450 208.050 220.050 ;
        RECT 217.950 219.450 220.050 220.050 ;
        RECT 205.950 218.400 220.050 219.450 ;
        RECT 205.950 217.950 208.050 218.400 ;
        RECT 217.950 217.950 220.050 218.400 ;
        RECT 223.950 217.950 226.050 220.050 ;
        RECT 241.950 217.950 244.050 220.050 ;
        RECT 247.950 217.950 250.050 220.050 ;
        RECT 265.950 217.950 268.050 220.950 ;
        RECT 335.400 220.050 336.450 223.950 ;
        RECT 365.850 221.700 367.050 225.300 ;
        RECT 385.950 224.400 388.050 226.500 ;
        RECT 409.950 225.450 412.050 226.050 ;
        RECT 430.800 225.450 432.900 226.050 ;
        RECT 409.950 224.400 432.900 225.450 ;
        RECT 271.950 217.950 274.050 220.050 ;
        RECT 310.950 217.950 313.050 220.050 ;
        RECT 316.950 217.950 319.050 220.050 ;
        RECT 334.950 217.950 337.050 220.050 ;
        RECT 346.950 217.950 349.050 220.050 ;
        RECT 352.950 219.450 355.050 220.050 ;
        RECT 357.000 219.450 361.050 220.050 ;
        RECT 364.950 219.600 367.050 221.700 ;
        RECT 352.950 218.400 361.050 219.450 ;
        RECT 352.950 217.950 355.050 218.400 ;
        RECT 357.000 217.950 361.050 218.400 ;
        RECT 199.950 214.950 202.050 217.050 ;
        RECT 217.950 214.950 220.050 216.750 ;
        RECT 223.950 214.950 226.050 216.750 ;
        RECT 241.950 214.950 244.050 216.750 ;
        RECT 247.950 214.950 250.050 216.750 ;
        RECT 265.950 214.950 268.050 216.750 ;
        RECT 271.950 214.950 274.050 216.750 ;
        RECT 292.950 214.950 295.050 217.050 ;
        RECT 310.950 214.950 313.050 216.750 ;
        RECT 316.950 214.950 319.050 216.750 ;
        RECT 334.950 214.950 337.050 216.750 ;
        RECT 346.950 214.950 349.050 216.750 ;
        RECT 352.950 214.950 355.050 216.750 ;
        RECT 199.950 211.950 202.050 213.750 ;
        RECT 220.950 212.250 223.050 214.050 ;
        RECT 226.950 212.250 229.050 214.050 ;
        RECT 244.950 212.250 247.050 214.050 ;
        RECT 250.950 212.250 253.050 214.050 ;
        RECT 262.950 212.250 265.050 214.050 ;
        RECT 268.950 212.250 271.050 214.050 ;
        RECT 292.950 211.950 295.050 213.750 ;
        RECT 313.950 212.250 316.050 214.050 ;
        RECT 319.950 212.250 322.050 214.050 ;
        RECT 337.950 212.250 340.050 214.050 ;
        RECT 349.950 212.250 352.050 214.050 ;
        RECT 361.950 212.250 364.050 214.050 ;
        RECT 220.950 208.950 223.050 211.050 ;
        RECT 226.950 208.950 229.050 211.050 ;
        RECT 232.950 210.450 235.050 211.050 ;
        RECT 244.950 210.450 247.050 211.050 ;
        RECT 232.950 209.400 247.050 210.450 ;
        RECT 232.950 208.950 235.050 209.400 ;
        RECT 244.950 208.950 247.050 209.400 ;
        RECT 250.950 208.950 253.050 211.050 ;
        RECT 262.950 208.950 265.050 211.050 ;
        RECT 268.950 210.450 271.050 211.050 ;
        RECT 283.950 210.450 286.050 211.050 ;
        RECT 268.950 209.400 286.050 210.450 ;
        RECT 268.950 208.950 271.050 209.400 ;
        RECT 283.950 208.950 286.050 209.400 ;
        RECT 289.950 209.250 292.050 211.050 ;
        RECT 295.950 209.250 298.050 211.050 ;
        RECT 307.950 210.450 312.000 211.050 ;
        RECT 313.950 210.450 316.050 211.050 ;
        RECT 307.950 209.400 316.050 210.450 ;
        RECT 307.950 208.950 312.000 209.400 ;
        RECT 313.950 208.950 316.050 209.400 ;
        RECT 319.950 208.950 322.050 211.050 ;
        RECT 325.950 210.450 328.050 211.050 ;
        RECT 337.950 210.450 340.050 211.050 ;
        RECT 325.950 209.400 340.050 210.450 ;
        RECT 325.950 208.950 328.050 209.400 ;
        RECT 337.950 208.950 340.050 209.400 ;
        RECT 133.950 203.400 160.050 204.450 ;
        RECT 133.950 202.950 136.050 203.400 ;
        RECT 157.950 202.950 160.050 203.400 ;
        RECT 175.950 202.500 178.050 204.600 ;
        RECT 196.950 202.500 199.050 204.600 ;
        RECT 221.400 204.450 222.450 208.950 ;
        RECT 289.950 205.950 292.050 208.050 ;
        RECT 295.950 205.950 298.050 208.050 ;
        RECT 349.950 205.950 352.050 211.050 ;
        RECT 358.950 208.950 364.050 211.050 ;
        RECT 241.950 204.450 244.050 205.050 ;
        RECT 221.400 203.400 244.050 204.450 ;
        RECT 241.950 202.950 244.050 203.400 ;
        RECT 319.950 204.450 322.050 205.050 ;
        RECT 331.950 204.450 334.050 205.050 ;
        RECT 365.850 204.600 367.050 219.600 ;
        RECT 379.950 214.950 382.050 217.050 ;
        RECT 379.950 211.950 382.050 213.750 ;
        RECT 386.100 204.600 387.300 224.400 ;
        RECT 409.950 223.950 412.050 224.400 ;
        RECT 430.800 223.950 432.900 224.400 ;
        RECT 434.100 225.450 436.200 226.050 ;
        RECT 448.950 225.450 451.050 226.050 ;
        RECT 463.950 225.450 466.050 226.050 ;
        RECT 434.100 224.400 466.050 225.450 ;
        RECT 469.950 224.400 472.050 226.500 ;
        RECT 490.950 225.300 493.050 227.400 ;
        RECT 511.950 226.950 514.050 227.400 ;
        RECT 547.950 226.950 550.050 227.400 ;
        RECT 529.950 225.450 532.050 226.050 ;
        RECT 538.950 225.450 541.050 226.050 ;
        RECT 434.100 223.950 436.200 224.400 ;
        RECT 448.950 223.950 451.050 224.400 ;
        RECT 463.950 223.950 466.050 224.400 ;
        RECT 388.950 222.450 391.050 223.050 ;
        RECT 394.950 222.450 397.050 223.050 ;
        RECT 388.950 221.400 397.050 222.450 ;
        RECT 388.950 220.950 391.050 221.400 ;
        RECT 394.950 220.950 397.050 221.400 ;
        RECT 409.950 217.950 412.050 220.050 ;
        RECT 415.950 217.950 418.050 220.050 ;
        RECT 388.950 214.950 391.050 217.050 ;
        RECT 409.950 214.950 412.050 216.750 ;
        RECT 415.950 214.950 418.050 216.750 ;
        RECT 430.950 214.950 433.050 220.050 ;
        RECT 448.950 217.950 451.050 220.050 ;
        RECT 454.950 217.950 457.050 220.050 ;
        RECT 448.950 214.950 451.050 216.750 ;
        RECT 454.950 214.950 457.050 216.750 ;
        RECT 466.950 214.950 469.050 217.050 ;
        RECT 388.950 211.950 391.050 213.750 ;
        RECT 406.950 212.250 409.050 214.050 ;
        RECT 412.950 212.250 415.050 214.050 ;
        RECT 430.950 211.950 433.050 213.750 ;
        RECT 451.950 212.250 454.050 214.050 ;
        RECT 457.950 212.250 460.050 214.050 ;
        RECT 466.950 211.950 469.050 213.750 ;
        RECT 391.950 210.450 394.050 211.050 ;
        RECT 406.950 210.450 409.050 211.050 ;
        RECT 391.950 209.400 409.050 210.450 ;
        RECT 391.950 208.950 394.050 209.400 ;
        RECT 406.950 208.950 409.050 209.400 ;
        RECT 412.950 208.950 415.050 211.050 ;
        RECT 427.950 209.250 430.050 211.050 ;
        RECT 433.950 209.250 436.050 211.050 ;
        RECT 439.950 210.450 442.050 211.050 ;
        RECT 451.950 210.450 454.050 211.050 ;
        RECT 439.950 209.400 454.050 210.450 ;
        RECT 439.950 208.950 442.050 209.400 ;
        RECT 451.950 208.950 454.050 209.400 ;
        RECT 457.950 208.950 460.050 211.050 ;
        RECT 421.950 207.450 426.000 208.050 ;
        RECT 427.950 207.450 430.050 208.050 ;
        RECT 421.950 206.400 430.050 207.450 ;
        RECT 421.950 205.950 426.000 206.400 ;
        RECT 427.950 205.950 430.050 206.400 ;
        RECT 433.950 205.950 436.050 208.050 ;
        RECT 319.950 203.400 334.050 204.450 ;
        RECT 319.950 202.950 322.050 203.400 ;
        RECT 331.950 202.950 334.050 203.400 ;
        RECT 364.950 202.500 367.050 204.600 ;
        RECT 385.950 202.500 388.050 204.600 ;
        RECT 442.950 204.450 445.050 205.050 ;
        RECT 458.400 204.450 459.450 208.950 ;
        RECT 470.700 204.600 471.900 224.400 ;
        RECT 490.950 221.700 492.150 225.300 ;
        RECT 529.950 224.400 541.050 225.450 ;
        RECT 571.950 224.400 574.050 226.500 ;
        RECT 592.950 225.300 595.050 227.400 ;
        RECT 661.950 226.950 664.050 227.400 ;
        RECT 715.950 226.950 718.050 227.400 ;
        RECT 754.950 228.450 757.050 229.050 ;
        RECT 763.950 228.450 766.050 229.050 ;
        RECT 754.950 227.400 766.050 228.450 ;
        RECT 754.950 226.950 757.050 227.400 ;
        RECT 763.950 226.950 766.050 227.400 ;
        RECT 631.950 225.450 634.050 226.050 ;
        RECT 769.950 225.450 772.050 226.050 ;
        RECT 529.950 223.950 532.050 224.400 ;
        RECT 538.950 223.950 541.050 224.400 ;
        RECT 499.950 222.450 502.050 223.050 ;
        RECT 526.950 222.450 529.050 223.050 ;
        RECT 490.950 219.600 493.050 221.700 ;
        RECT 499.950 221.400 529.050 222.450 ;
        RECT 499.950 220.950 502.050 221.400 ;
        RECT 526.950 220.950 529.050 221.400 ;
        RECT 475.950 214.950 478.050 217.050 ;
        RECT 475.950 211.950 478.050 213.750 ;
        RECT 490.950 204.600 492.150 219.600 ;
        RECT 532.950 217.950 535.050 220.050 ;
        RECT 538.950 217.950 541.050 220.050 ;
        RECT 553.950 217.950 556.050 220.050 ;
        RECT 559.950 217.950 562.050 220.050 ;
        RECT 505.950 216.450 510.000 217.050 ;
        RECT 511.950 216.450 514.050 217.050 ;
        RECT 505.950 215.400 514.050 216.450 ;
        RECT 505.950 214.950 510.000 215.400 ;
        RECT 511.950 214.950 514.050 215.400 ;
        RECT 532.950 214.950 535.050 216.750 ;
        RECT 538.950 214.950 541.050 216.750 ;
        RECT 553.950 214.950 556.050 216.750 ;
        RECT 559.950 214.950 562.050 216.750 ;
        RECT 568.950 214.950 571.050 217.050 ;
        RECT 493.950 212.250 496.050 214.050 ;
        RECT 511.950 211.950 514.050 213.750 ;
        RECT 535.950 212.250 538.050 214.050 ;
        RECT 556.950 212.250 559.050 214.050 ;
        RECT 562.950 212.250 565.050 214.050 ;
        RECT 568.950 211.950 571.050 213.750 ;
        RECT 493.950 208.950 496.050 211.050 ;
        RECT 508.950 209.250 511.050 211.050 ;
        RECT 514.950 209.250 517.050 211.050 ;
        RECT 535.950 210.450 538.050 211.050 ;
        RECT 550.950 210.450 553.050 211.050 ;
        RECT 535.950 209.400 553.050 210.450 ;
        RECT 535.950 208.950 538.050 209.400 ;
        RECT 550.950 208.950 553.050 209.400 ;
        RECT 556.950 208.950 559.050 211.050 ;
        RECT 562.950 208.950 565.050 211.050 ;
        RECT 499.950 207.450 502.050 208.050 ;
        RECT 508.950 207.450 511.050 208.050 ;
        RECT 499.950 206.400 511.050 207.450 ;
        RECT 499.950 205.950 502.050 206.400 ;
        RECT 508.950 205.950 511.050 206.400 ;
        RECT 514.950 205.950 517.050 208.050 ;
        RECT 442.950 203.400 459.450 204.450 ;
        RECT 442.950 202.950 445.050 203.400 ;
        RECT 469.950 202.500 472.050 204.600 ;
        RECT 490.950 202.500 493.050 204.600 ;
        RECT 556.950 204.450 559.050 205.050 ;
        RECT 565.950 204.450 568.050 205.050 ;
        RECT 572.700 204.600 573.900 224.400 ;
        RECT 592.950 221.700 594.150 225.300 ;
        RECT 631.950 224.400 699.450 225.450 ;
        RECT 631.950 223.950 634.050 224.400 ;
        RECT 698.400 223.050 699.450 224.400 ;
        RECT 752.400 224.400 772.050 225.450 ;
        RECT 781.950 225.300 784.050 227.400 ;
        RECT 664.950 222.450 667.050 223.050 ;
        RECT 679.950 222.450 682.050 223.050 ;
        RECT 592.950 219.600 595.050 221.700 ;
        RECT 664.950 221.400 682.050 222.450 ;
        RECT 664.950 220.950 667.050 221.400 ;
        RECT 679.950 220.950 682.050 221.400 ;
        RECT 697.950 222.450 700.050 223.050 ;
        RECT 703.950 222.450 706.050 223.050 ;
        RECT 697.950 221.400 706.050 222.450 ;
        RECT 697.950 220.950 700.050 221.400 ;
        RECT 703.950 220.950 706.050 221.400 ;
        RECT 752.400 220.050 753.450 224.400 ;
        RECT 769.950 223.950 772.050 224.400 ;
        RECT 782.850 221.700 784.050 225.300 ;
        RECT 802.950 224.400 805.050 226.500 ;
        RECT 817.950 225.300 820.050 227.400 ;
        RECT 577.950 214.950 580.050 217.050 ;
        RECT 577.950 211.950 580.050 213.750 ;
        RECT 592.950 204.600 594.150 219.600 ;
        RECT 613.950 219.450 616.050 220.050 ;
        RECT 625.950 219.450 628.050 220.050 ;
        RECT 613.950 218.400 628.050 219.450 ;
        RECT 613.950 217.950 616.050 218.400 ;
        RECT 625.950 217.950 628.050 218.400 ;
        RECT 631.950 217.950 634.050 220.050 ;
        RECT 637.950 217.950 640.050 220.050 ;
        RECT 655.950 217.950 658.050 220.050 ;
        RECT 661.950 217.950 664.050 220.050 ;
        RECT 721.950 217.950 724.050 220.050 ;
        RECT 727.950 217.950 730.050 220.050 ;
        RECT 745.950 217.950 748.050 220.050 ;
        RECT 751.950 217.950 754.050 220.050 ;
        RECT 763.950 217.950 766.050 220.050 ;
        RECT 769.950 219.450 772.050 220.050 ;
        RECT 774.000 219.450 778.050 220.050 ;
        RECT 781.950 219.600 784.050 221.700 ;
        RECT 769.950 218.400 778.050 219.450 ;
        RECT 769.950 217.950 772.050 218.400 ;
        RECT 774.000 217.950 778.050 218.400 ;
        RECT 613.950 214.950 616.050 216.750 ;
        RECT 631.950 214.950 634.050 216.750 ;
        RECT 637.950 214.950 640.050 216.750 ;
        RECT 655.950 214.950 658.050 216.750 ;
        RECT 661.950 214.950 664.050 216.750 ;
        RECT 679.950 216.450 682.050 217.050 ;
        RECT 688.950 216.450 691.050 217.050 ;
        RECT 679.950 215.400 691.050 216.450 ;
        RECT 679.950 214.950 682.050 215.400 ;
        RECT 688.950 214.950 691.050 215.400 ;
        RECT 697.950 214.950 703.050 217.050 ;
        RECT 721.950 214.950 724.050 216.750 ;
        RECT 727.950 214.950 730.050 216.750 ;
        RECT 745.950 214.950 748.050 216.750 ;
        RECT 751.950 214.950 754.050 216.750 ;
        RECT 763.950 214.950 766.050 216.750 ;
        RECT 769.950 214.950 772.050 216.750 ;
        RECT 595.950 212.250 598.050 214.050 ;
        RECT 610.950 212.250 613.050 214.050 ;
        RECT 628.950 212.250 631.050 214.050 ;
        RECT 634.950 212.250 637.050 214.050 ;
        RECT 658.950 212.250 661.050 214.050 ;
        RECT 664.950 212.250 667.050 214.050 ;
        RECT 679.950 211.950 682.050 213.750 ;
        RECT 700.950 211.950 703.050 213.750 ;
        RECT 718.950 212.250 721.050 214.050 ;
        RECT 724.950 212.250 727.050 214.050 ;
        RECT 748.950 212.250 751.050 214.050 ;
        RECT 766.950 212.250 769.050 214.050 ;
        RECT 778.950 212.250 781.050 214.050 ;
        RECT 595.950 208.950 598.050 211.050 ;
        RECT 610.950 208.950 613.050 211.050 ;
        RECT 628.950 208.950 631.050 211.050 ;
        RECT 634.950 208.950 637.050 211.050 ;
        RECT 640.950 210.450 643.050 211.050 ;
        RECT 658.950 210.450 661.050 211.050 ;
        RECT 640.950 209.400 661.050 210.450 ;
        RECT 640.950 208.950 643.050 209.400 ;
        RECT 658.950 208.950 661.050 209.400 ;
        RECT 664.950 208.950 667.050 211.050 ;
        RECT 676.950 209.250 679.050 211.050 ;
        RECT 682.950 209.250 685.050 211.050 ;
        RECT 697.950 209.250 700.050 211.050 ;
        RECT 703.950 209.250 706.050 211.050 ;
        RECT 718.950 208.950 721.050 211.050 ;
        RECT 556.950 203.400 568.050 204.450 ;
        RECT 556.950 202.950 559.050 203.400 ;
        RECT 565.950 202.950 568.050 203.400 ;
        RECT 571.950 202.500 574.050 204.600 ;
        RECT 592.950 202.500 595.050 204.600 ;
        RECT 601.950 204.450 604.050 205.050 ;
        RECT 635.400 204.450 636.450 208.950 ;
        RECT 676.950 207.450 679.050 208.050 ;
        RECT 671.400 206.400 679.050 207.450 ;
        RECT 601.950 203.400 636.450 204.450 ;
        RECT 664.950 204.450 667.050 205.050 ;
        RECT 671.400 204.450 672.450 206.400 ;
        RECT 676.950 205.950 679.050 206.400 ;
        RECT 682.950 205.950 685.050 208.050 ;
        RECT 688.950 207.450 691.050 208.050 ;
        RECT 697.950 207.450 700.050 208.050 ;
        RECT 688.950 206.400 700.050 207.450 ;
        RECT 688.950 205.950 691.050 206.400 ;
        RECT 697.950 205.950 700.050 206.400 ;
        RECT 703.950 205.950 706.050 208.050 ;
        RECT 724.950 205.950 727.050 211.050 ;
        RECT 730.950 210.450 733.050 211.050 ;
        RECT 748.950 210.450 751.050 211.050 ;
        RECT 730.950 209.400 751.050 210.450 ;
        RECT 730.950 208.950 733.050 209.400 ;
        RECT 748.950 208.950 751.050 209.400 ;
        RECT 766.950 210.450 769.050 211.050 ;
        RECT 771.000 210.450 775.050 211.050 ;
        RECT 766.950 209.400 775.050 210.450 ;
        RECT 766.950 208.950 769.050 209.400 ;
        RECT 771.000 208.950 775.050 209.400 ;
        RECT 778.950 208.950 781.050 211.050 ;
        RECT 782.850 204.600 784.050 219.600 ;
        RECT 796.950 214.950 799.050 217.050 ;
        RECT 796.950 211.950 799.050 213.750 ;
        RECT 803.100 204.600 804.300 224.400 ;
        RECT 818.850 221.700 820.050 225.300 ;
        RECT 838.950 224.400 841.050 226.500 ;
        RECT 853.950 224.400 856.050 226.500 ;
        RECT 874.950 225.300 877.050 227.400 ;
        RECT 892.950 225.450 895.050 226.050 ;
        RECT 898.950 225.450 901.050 226.050 ;
        RECT 817.950 219.600 820.050 221.700 ;
        RECT 805.950 214.950 808.050 217.050 ;
        RECT 805.950 211.950 808.050 213.750 ;
        RECT 814.950 212.250 817.050 214.050 ;
        RECT 814.950 208.950 817.050 211.050 ;
        RECT 818.850 204.600 820.050 219.600 ;
        RECT 823.950 216.450 826.050 217.050 ;
        RECT 832.950 216.450 835.050 217.050 ;
        RECT 823.950 215.400 835.050 216.450 ;
        RECT 823.950 214.950 826.050 215.400 ;
        RECT 832.950 214.950 835.050 215.400 ;
        RECT 832.950 211.950 835.050 213.750 ;
        RECT 839.100 204.600 840.300 224.400 ;
        RECT 841.950 214.950 844.050 217.050 ;
        RECT 850.950 214.950 853.050 217.050 ;
        RECT 841.950 211.950 844.050 213.750 ;
        RECT 850.950 211.950 853.050 213.750 ;
        RECT 841.950 207.450 844.050 208.050 ;
        RECT 850.950 207.450 853.050 208.050 ;
        RECT 841.950 206.400 853.050 207.450 ;
        RECT 841.950 205.950 844.050 206.400 ;
        RECT 850.950 205.950 853.050 206.400 ;
        RECT 854.700 204.600 855.900 224.400 ;
        RECT 874.950 221.700 876.150 225.300 ;
        RECT 892.950 224.400 901.050 225.450 ;
        RECT 892.950 223.950 895.050 224.400 ;
        RECT 898.950 223.950 901.050 224.400 ;
        RECT 859.950 214.950 862.050 220.050 ;
        RECT 874.950 219.600 877.050 221.700 ;
        RECT 859.950 211.950 862.050 213.750 ;
        RECT 874.950 204.600 876.150 219.600 ;
        RECT 898.950 217.950 901.050 220.050 ;
        RECT 904.950 217.950 907.050 220.050 ;
        RECT 898.950 214.950 901.050 216.750 ;
        RECT 904.950 214.950 907.050 216.750 ;
        RECT 877.950 212.250 880.050 214.050 ;
        RECT 895.950 212.250 898.050 214.050 ;
        RECT 901.950 212.250 904.050 214.050 ;
        RECT 877.950 208.950 880.050 211.050 ;
        RECT 883.950 210.450 886.050 211.050 ;
        RECT 895.950 210.450 898.050 211.050 ;
        RECT 883.950 209.400 898.050 210.450 ;
        RECT 883.950 208.950 886.050 209.400 ;
        RECT 895.950 208.950 898.050 209.400 ;
        RECT 901.950 208.950 904.050 211.050 ;
        RECT 664.950 203.400 672.450 204.450 ;
        RECT 601.950 202.950 604.050 203.400 ;
        RECT 664.950 202.950 667.050 203.400 ;
        RECT 202.950 201.450 205.050 202.050 ;
        RECT 208.950 201.450 211.050 202.050 ;
        RECT 202.950 200.400 211.050 201.450 ;
        RECT 202.950 199.950 205.050 200.400 ;
        RECT 208.950 199.950 211.050 200.400 ;
        RECT 226.950 201.450 229.050 202.050 ;
        RECT 259.950 201.450 262.050 202.050 ;
        RECT 226.950 200.400 262.050 201.450 ;
        RECT 226.950 199.950 229.050 200.400 ;
        RECT 259.950 199.950 262.050 200.400 ;
        RECT 286.950 201.450 289.050 202.050 ;
        RECT 292.950 201.450 295.050 202.050 ;
        RECT 286.950 200.400 295.050 201.450 ;
        RECT 286.950 199.950 289.050 200.400 ;
        RECT 292.950 199.950 295.050 200.400 ;
        RECT 394.950 201.450 397.050 202.050 ;
        RECT 538.950 201.450 541.050 202.050 ;
        RECT 562.950 201.450 565.050 202.050 ;
        RECT 394.950 200.400 438.450 201.450 ;
        RECT 394.950 199.950 397.050 200.400 ;
        RECT 97.950 198.450 100.050 199.050 ;
        RECT 133.950 198.450 136.050 199.050 ;
        RECT 97.950 197.400 136.050 198.450 ;
        RECT 97.950 196.950 100.050 197.400 ;
        RECT 133.950 196.950 136.050 197.400 ;
        RECT 163.950 198.450 166.050 199.050 ;
        RECT 172.950 198.450 175.050 199.050 ;
        RECT 205.950 198.450 208.050 199.050 ;
        RECT 163.950 197.400 208.050 198.450 ;
        RECT 163.950 196.950 166.050 197.400 ;
        RECT 172.950 196.950 175.050 197.400 ;
        RECT 205.950 196.950 208.050 197.400 ;
        RECT 412.950 198.450 415.050 199.050 ;
        RECT 433.950 198.450 436.050 199.050 ;
        RECT 412.950 197.400 436.050 198.450 ;
        RECT 412.950 196.950 415.050 197.400 ;
        RECT 433.950 196.950 436.050 197.400 ;
        RECT 13.950 195.450 16.050 196.050 ;
        RECT 19.950 195.450 22.050 196.050 ;
        RECT 13.950 194.400 22.050 195.450 ;
        RECT 13.950 193.950 16.050 194.400 ;
        RECT 19.950 193.950 22.050 194.400 ;
        RECT 91.950 195.450 94.050 196.050 ;
        RECT 112.950 195.450 115.050 196.050 ;
        RECT 91.950 194.400 115.050 195.450 ;
        RECT 91.950 193.950 94.050 194.400 ;
        RECT 112.950 193.950 115.050 194.400 ;
        RECT 136.950 195.450 139.050 196.050 ;
        RECT 187.950 195.450 190.050 196.050 ;
        RECT 136.950 194.400 190.050 195.450 ;
        RECT 136.950 193.950 139.050 194.400 ;
        RECT 187.950 193.950 190.050 194.400 ;
        RECT 223.950 195.450 226.050 196.050 ;
        RECT 265.950 195.450 268.050 196.050 ;
        RECT 355.950 195.450 358.050 196.050 ;
        RECT 394.950 195.450 397.050 196.050 ;
        RECT 223.950 194.400 397.050 195.450 ;
        RECT 437.400 195.450 438.450 200.400 ;
        RECT 538.950 200.400 565.050 201.450 ;
        RECT 538.950 199.950 541.050 200.400 ;
        RECT 562.950 199.950 565.050 200.400 ;
        RECT 610.950 201.450 613.050 202.050 ;
        RECT 665.400 201.450 666.450 202.950 ;
        RECT 781.950 202.500 784.050 204.600 ;
        RECT 802.950 202.500 805.050 204.600 ;
        RECT 817.950 202.500 820.050 204.600 ;
        RECT 838.950 202.500 841.050 204.600 ;
        RECT 853.950 202.500 856.050 204.600 ;
        RECT 874.950 202.500 877.050 204.600 ;
        RECT 610.950 200.400 666.450 201.450 ;
        RECT 679.950 201.450 682.050 202.050 ;
        RECT 688.950 201.450 691.050 202.050 ;
        RECT 679.950 200.400 691.050 201.450 ;
        RECT 610.950 199.950 613.050 200.400 ;
        RECT 679.950 199.950 682.050 200.400 ;
        RECT 688.950 199.950 691.050 200.400 ;
        RECT 724.950 201.450 727.050 202.050 ;
        RECT 883.950 201.450 886.050 202.050 ;
        RECT 901.950 201.450 904.050 202.050 ;
        RECT 724.950 200.400 777.450 201.450 ;
        RECT 724.950 199.950 727.050 200.400 ;
        RECT 466.950 198.450 469.050 199.050 ;
        RECT 475.950 198.450 478.050 199.050 ;
        RECT 547.950 198.450 550.050 199.050 ;
        RECT 580.950 198.450 583.050 199.050 ;
        RECT 466.950 197.400 543.450 198.450 ;
        RECT 466.950 196.950 469.050 197.400 ;
        RECT 475.950 196.950 478.050 197.400 ;
        RECT 467.400 195.450 468.450 196.950 ;
        RECT 437.400 194.400 468.450 195.450 ;
        RECT 472.950 195.450 475.050 196.050 ;
        RECT 538.950 195.450 541.050 196.050 ;
        RECT 472.950 194.400 541.050 195.450 ;
        RECT 542.400 195.450 543.450 197.400 ;
        RECT 547.950 197.400 583.050 198.450 ;
        RECT 547.950 196.950 550.050 197.400 ;
        RECT 580.950 196.950 583.050 197.400 ;
        RECT 595.950 198.450 598.050 199.050 ;
        RECT 611.400 198.450 612.450 199.950 ;
        RECT 595.950 197.400 612.450 198.450 ;
        RECT 763.950 198.450 766.050 199.050 ;
        RECT 772.950 198.450 775.050 199.050 ;
        RECT 763.950 197.400 775.050 198.450 ;
        RECT 776.400 198.450 777.450 200.400 ;
        RECT 883.950 200.400 904.050 201.450 ;
        RECT 883.950 199.950 886.050 200.400 ;
        RECT 901.950 199.950 904.050 200.400 ;
        RECT 796.950 198.450 799.050 199.050 ;
        RECT 776.400 197.400 799.050 198.450 ;
        RECT 595.950 196.950 598.050 197.400 ;
        RECT 763.950 196.950 766.050 197.400 ;
        RECT 772.950 196.950 775.050 197.400 ;
        RECT 796.950 196.950 799.050 197.400 ;
        RECT 850.950 198.450 853.050 199.050 ;
        RECT 883.950 198.450 886.050 199.050 ;
        RECT 850.950 197.400 886.050 198.450 ;
        RECT 850.950 196.950 853.050 197.400 ;
        RECT 883.950 196.950 886.050 197.400 ;
        RECT 553.950 195.450 556.050 196.050 ;
        RECT 542.400 194.400 556.050 195.450 ;
        RECT 223.950 193.950 226.050 194.400 ;
        RECT 265.950 193.950 268.050 194.400 ;
        RECT 355.950 193.950 358.050 194.400 ;
        RECT 394.950 193.950 397.050 194.400 ;
        RECT 472.950 193.950 475.050 194.400 ;
        RECT 538.950 193.950 541.050 194.400 ;
        RECT 553.950 193.950 556.050 194.400 ;
        RECT 790.950 195.450 793.050 196.050 ;
        RECT 826.950 195.450 829.050 196.050 ;
        RECT 790.950 194.400 829.050 195.450 ;
        RECT 790.950 193.950 793.050 194.400 ;
        RECT 826.950 193.950 829.050 194.400 ;
        RECT 871.950 195.450 874.050 196.050 ;
        RECT 871.950 195.000 885.450 195.450 ;
        RECT 871.950 194.400 886.050 195.000 ;
        RECT 871.950 193.950 874.050 194.400 ;
        RECT 22.950 192.450 25.050 193.050 ;
        RECT 28.950 192.450 31.050 193.050 ;
        RECT 22.950 191.400 31.050 192.450 ;
        RECT 22.950 190.950 25.050 191.400 ;
        RECT 28.950 190.950 31.050 191.400 ;
        RECT 100.950 192.450 103.050 193.050 ;
        RECT 139.950 192.450 142.050 193.050 ;
        RECT 100.950 191.400 142.050 192.450 ;
        RECT 100.950 190.950 103.050 191.400 ;
        RECT 139.950 190.950 142.050 191.400 ;
        RECT 196.950 192.450 199.050 193.050 ;
        RECT 214.950 192.450 217.050 193.050 ;
        RECT 196.950 191.400 217.050 192.450 ;
        RECT 196.950 190.950 199.050 191.400 ;
        RECT 214.950 190.950 217.050 191.400 ;
        RECT 319.950 192.450 322.050 193.050 ;
        RECT 325.950 192.450 328.050 193.050 ;
        RECT 319.950 191.400 328.050 192.450 ;
        RECT 319.950 190.950 322.050 191.400 ;
        RECT 325.950 190.950 328.050 191.400 ;
        RECT 331.950 192.450 334.050 193.050 ;
        RECT 367.950 192.450 370.050 193.050 ;
        RECT 331.950 191.400 370.050 192.450 ;
        RECT 331.950 190.950 334.050 191.400 ;
        RECT 367.950 190.950 370.050 191.400 ;
        RECT 427.950 192.450 430.050 193.050 ;
        RECT 433.950 192.450 436.050 193.050 ;
        RECT 427.950 191.400 436.050 192.450 ;
        RECT 427.950 190.950 430.050 191.400 ;
        RECT 433.950 190.950 436.050 191.400 ;
        RECT 451.950 192.450 454.050 193.050 ;
        RECT 457.950 192.450 460.050 193.050 ;
        RECT 490.950 192.450 493.050 193.050 ;
        RECT 511.950 192.450 514.050 193.050 ;
        RECT 451.950 191.400 514.050 192.450 ;
        RECT 451.950 190.950 454.050 191.400 ;
        RECT 457.950 190.950 460.050 191.400 ;
        RECT 490.950 190.950 493.050 191.400 ;
        RECT 511.950 190.950 514.050 191.400 ;
        RECT 574.950 192.450 577.050 193.050 ;
        RECT 619.950 192.450 622.050 193.050 ;
        RECT 643.950 192.450 646.050 193.050 ;
        RECT 658.950 192.450 661.050 193.050 ;
        RECT 574.950 191.400 661.050 192.450 ;
        RECT 574.950 190.950 577.050 191.400 ;
        RECT 619.950 190.950 622.050 191.400 ;
        RECT 643.950 190.950 646.050 191.400 ;
        RECT 658.950 190.950 661.050 191.400 ;
        RECT 685.950 192.450 688.050 193.050 ;
        RECT 697.950 192.450 700.050 193.050 ;
        RECT 685.950 191.400 700.050 192.450 ;
        RECT 685.950 190.950 688.050 191.400 ;
        RECT 697.950 190.950 700.050 191.400 ;
        RECT 703.950 192.450 706.050 193.050 ;
        RECT 721.950 192.450 724.050 193.050 ;
        RECT 703.950 191.400 724.050 192.450 ;
        RECT 703.950 190.950 706.050 191.400 ;
        RECT 721.950 190.950 724.050 191.400 ;
        RECT 751.950 192.450 754.050 193.050 ;
        RECT 820.950 192.450 823.050 193.050 ;
        RECT 877.950 192.450 880.050 193.050 ;
        RECT 751.950 191.400 880.050 192.450 ;
        RECT 751.950 190.950 754.050 191.400 ;
        RECT 46.950 189.450 49.050 190.050 ;
        RECT 52.950 189.450 55.050 190.050 ;
        RECT 46.950 188.400 55.050 189.450 ;
        RECT 148.950 188.400 151.050 190.500 ;
        RECT 169.950 188.400 172.050 190.500 ;
        RECT 175.950 189.450 178.050 190.050 ;
        RECT 253.950 189.450 256.050 190.050 ;
        RECT 271.950 189.450 274.050 190.050 ;
        RECT 283.950 189.450 286.050 190.050 ;
        RECT 175.950 188.400 195.450 189.450 ;
        RECT 46.950 187.950 49.050 188.400 ;
        RECT 52.950 187.950 55.050 188.400 ;
        RECT 13.950 184.950 16.050 187.050 ;
        RECT 19.950 184.950 22.050 187.050 ;
        RECT 91.950 184.950 97.050 187.050 ;
        RECT 100.950 184.950 103.050 187.050 ;
        RECT 13.950 181.950 16.050 183.750 ;
        RECT 19.950 181.950 22.050 183.750 ;
        RECT 31.950 181.950 34.050 184.050 ;
        RECT 37.950 183.450 40.050 184.050 ;
        RECT 49.950 183.450 52.050 184.050 ;
        RECT 37.950 182.400 52.050 183.450 ;
        RECT 37.950 181.950 40.050 182.400 ;
        RECT 49.950 181.950 52.050 182.400 ;
        RECT 55.950 181.950 58.050 184.050 ;
        RECT 76.950 183.450 79.050 184.050 ;
        RECT 88.950 183.450 91.050 184.050 ;
        RECT 76.950 182.400 91.050 183.450 ;
        RECT 76.950 181.950 79.050 182.400 ;
        RECT 88.950 181.950 91.050 182.400 ;
        RECT 94.950 181.950 97.050 183.750 ;
        RECT 100.950 181.950 103.050 183.750 ;
        RECT 115.950 181.950 118.050 184.050 ;
        RECT 133.950 183.450 136.050 184.050 ;
        RECT 138.000 183.450 142.050 184.050 ;
        RECT 133.950 182.400 142.050 183.450 ;
        RECT 133.950 181.950 136.050 182.400 ;
        RECT 138.000 181.950 142.050 182.400 ;
        RECT 145.950 181.950 148.050 184.050 ;
        RECT 16.950 179.250 19.050 181.050 ;
        RECT 31.950 178.950 34.050 180.750 ;
        RECT 37.950 178.950 40.050 180.750 ;
        RECT 55.950 178.950 58.050 180.750 ;
        RECT 76.950 178.950 79.050 180.750 ;
        RECT 97.950 179.250 100.050 181.050 ;
        RECT 115.950 178.950 118.050 180.750 ;
        RECT 133.950 178.950 136.050 180.750 ;
        RECT 145.950 178.950 148.050 180.750 ;
        RECT 13.950 175.950 19.050 178.050 ;
        RECT 34.950 176.250 37.050 178.050 ;
        RECT 40.950 176.250 43.050 178.050 ;
        RECT 58.950 176.250 61.050 178.050 ;
        RECT 73.950 176.250 76.050 178.050 ;
        RECT 79.950 176.250 82.050 178.050 ;
        RECT 94.950 175.950 100.050 178.050 ;
        RECT 118.950 176.250 121.050 178.050 ;
        RECT 136.950 176.250 139.050 178.050 ;
        RECT 34.950 172.950 37.050 175.050 ;
        RECT 40.950 174.450 43.050 175.050 ;
        RECT 58.950 174.450 61.050 175.050 ;
        RECT 40.950 173.400 61.050 174.450 ;
        RECT 40.950 172.950 43.050 173.400 ;
        RECT 58.950 172.950 61.050 173.400 ;
        RECT 73.950 172.950 76.050 175.050 ;
        RECT 79.950 172.950 82.050 175.050 ;
        RECT 118.950 172.950 121.050 175.050 ;
        RECT 133.950 172.950 139.050 175.050 ;
        RECT 149.850 173.400 151.050 188.400 ;
        RECT 163.950 179.250 166.050 181.050 ;
        RECT 163.950 175.950 166.050 178.050 ;
        RECT 16.950 171.450 19.050 172.050 ;
        RECT 22.950 171.450 25.050 172.050 ;
        RECT 31.950 171.450 34.050 172.050 ;
        RECT 16.950 170.400 34.050 171.450 ;
        RECT 148.950 171.300 151.050 173.400 ;
        RECT 16.950 169.950 19.050 170.400 ;
        RECT 22.950 169.950 25.050 170.400 ;
        RECT 31.950 169.950 34.050 170.400 ;
        RECT 49.950 168.450 52.050 169.050 ;
        RECT 79.950 168.450 82.050 169.050 ;
        RECT 49.950 167.400 82.050 168.450 ;
        RECT 149.850 167.700 151.050 171.300 ;
        RECT 170.100 168.600 171.300 188.400 ;
        RECT 175.950 187.950 178.050 188.400 ;
        RECT 194.400 184.050 195.450 188.400 ;
        RECT 253.950 188.400 286.050 189.450 ;
        RECT 289.950 188.400 292.050 190.500 ;
        RECT 310.950 188.400 313.050 190.500 ;
        RECT 319.950 189.450 322.050 190.050 ;
        RECT 352.950 189.450 355.050 190.050 ;
        RECT 373.950 189.450 376.050 190.050 ;
        RECT 319.950 188.400 336.450 189.450 ;
        RECT 253.950 187.950 256.050 188.400 ;
        RECT 271.950 187.950 274.050 188.400 ;
        RECT 283.950 187.950 286.050 188.400 ;
        RECT 187.950 181.950 190.050 184.050 ;
        RECT 193.950 181.950 196.050 184.050 ;
        RECT 238.950 183.450 241.050 184.050 ;
        RECT 256.950 183.450 259.050 184.050 ;
        RECT 238.950 182.400 259.050 183.450 ;
        RECT 238.950 181.950 241.050 182.400 ;
        RECT 256.950 181.950 259.050 182.400 ;
        RECT 280.950 181.950 283.050 184.050 ;
        RECT 286.950 181.950 289.050 184.050 ;
        RECT 172.950 179.250 175.050 181.050 ;
        RECT 187.950 178.950 190.050 180.750 ;
        RECT 193.950 178.950 196.050 180.750 ;
        RECT 214.950 179.250 217.050 181.050 ;
        RECT 235.950 179.250 238.050 181.050 ;
        RECT 256.950 178.950 259.050 180.750 ;
        RECT 274.950 179.250 277.050 181.050 ;
        RECT 280.950 178.950 283.050 180.750 ;
        RECT 286.950 178.950 289.050 180.750 ;
        RECT 172.950 175.950 175.050 178.050 ;
        RECT 190.950 176.250 193.050 178.050 ;
        RECT 196.950 176.250 199.050 178.050 ;
        RECT 205.950 177.450 208.050 178.050 ;
        RECT 214.950 177.450 217.050 178.050 ;
        RECT 205.950 176.400 217.050 177.450 ;
        RECT 205.950 175.950 208.050 176.400 ;
        RECT 214.950 175.950 217.050 176.400 ;
        RECT 253.950 176.250 256.050 178.050 ;
        RECT 259.950 176.250 262.050 178.050 ;
        RECT 265.950 177.450 268.050 178.050 ;
        RECT 274.950 177.450 277.050 178.050 ;
        RECT 265.950 176.400 277.050 177.450 ;
        RECT 265.950 175.950 268.050 176.400 ;
        RECT 274.950 175.950 277.050 176.400 ;
        RECT 190.950 172.950 193.050 175.050 ;
        RECT 196.950 172.950 199.050 175.050 ;
        RECT 253.950 172.950 256.050 175.050 ;
        RECT 259.950 172.950 262.050 175.050 ;
        RECT 290.850 173.400 292.050 188.400 ;
        RECT 304.950 179.250 307.050 181.050 ;
        RECT 304.950 175.950 307.050 178.050 ;
        RECT 289.950 171.300 292.050 173.400 ;
        RECT 49.950 166.950 52.050 167.400 ;
        RECT 79.950 166.950 82.050 167.400 ;
        RECT 67.950 165.450 70.050 166.050 ;
        RECT 91.950 165.450 94.050 166.050 ;
        RECT 148.950 165.600 151.050 167.700 ;
        RECT 169.950 166.500 172.050 168.600 ;
        RECT 190.950 168.450 193.050 169.050 ;
        RECT 259.950 168.450 262.050 169.050 ;
        RECT 265.950 168.450 268.050 169.050 ;
        RECT 190.950 167.400 268.050 168.450 ;
        RECT 290.850 167.700 292.050 171.300 ;
        RECT 311.100 168.600 312.300 188.400 ;
        RECT 319.950 187.950 322.050 188.400 ;
        RECT 335.400 184.050 336.450 188.400 ;
        RECT 352.950 188.400 376.050 189.450 ;
        RECT 352.950 187.950 355.050 188.400 ;
        RECT 373.950 187.950 376.050 188.400 ;
        RECT 409.950 189.450 412.050 190.050 ;
        RECT 427.950 189.450 430.050 190.050 ;
        RECT 409.950 188.400 430.050 189.450 ;
        RECT 409.950 187.950 412.050 188.400 ;
        RECT 427.950 187.950 430.050 188.400 ;
        RECT 436.950 189.450 439.050 190.050 ;
        RECT 463.950 189.450 466.050 190.050 ;
        RECT 436.950 188.400 466.050 189.450 ;
        RECT 529.950 188.400 532.050 190.500 ;
        RECT 550.950 188.400 553.050 190.500 ;
        RECT 637.950 189.450 640.050 190.050 ;
        RECT 667.950 189.450 670.050 190.050 ;
        RECT 727.950 189.450 730.050 190.050 ;
        RECT 637.950 188.400 670.050 189.450 ;
        RECT 436.950 187.950 439.050 188.400 ;
        RECT 463.950 187.950 466.050 188.400 ;
        RECT 328.950 181.950 331.050 184.050 ;
        RECT 334.950 181.950 337.050 184.050 ;
        RECT 343.950 183.450 346.050 184.050 ;
        RECT 355.950 183.450 358.050 184.050 ;
        RECT 343.950 182.400 358.050 183.450 ;
        RECT 343.950 181.950 346.050 182.400 ;
        RECT 355.950 181.950 358.050 182.400 ;
        RECT 415.950 183.450 418.050 184.050 ;
        RECT 427.950 183.450 430.050 184.050 ;
        RECT 415.950 182.400 430.050 183.450 ;
        RECT 415.950 181.950 418.050 182.400 ;
        RECT 427.950 181.950 430.050 182.400 ;
        RECT 433.950 181.950 436.050 184.050 ;
        RECT 457.950 183.450 460.050 184.050 ;
        RECT 463.950 183.450 466.050 184.050 ;
        RECT 457.950 182.400 466.050 183.450 ;
        RECT 457.950 181.950 460.050 182.400 ;
        RECT 463.950 181.950 466.050 182.400 ;
        RECT 496.950 183.450 499.050 184.050 ;
        RECT 505.950 183.450 508.050 184.050 ;
        RECT 514.950 183.450 517.050 184.050 ;
        RECT 496.950 182.400 504.450 183.450 ;
        RECT 496.950 181.950 499.050 182.400 ;
        RECT 313.950 179.250 316.050 181.050 ;
        RECT 328.950 178.950 331.050 180.750 ;
        RECT 334.950 178.950 337.050 180.750 ;
        RECT 355.950 178.950 358.050 180.750 ;
        RECT 376.950 179.250 379.050 181.050 ;
        RECT 397.950 179.250 400.050 181.050 ;
        RECT 415.950 178.950 418.050 180.750 ;
        RECT 433.950 178.950 436.050 180.750 ;
        RECT 454.950 179.250 457.050 181.050 ;
        RECT 475.950 179.250 478.050 181.050 ;
        RECT 496.950 178.950 499.050 180.750 ;
        RECT 503.400 180.450 504.450 182.400 ;
        RECT 505.950 182.400 517.050 183.450 ;
        RECT 505.950 181.950 508.050 182.400 ;
        RECT 514.950 181.950 517.050 182.400 ;
        RECT 526.950 181.950 529.050 184.050 ;
        RECT 508.950 180.450 511.050 181.050 ;
        RECT 503.400 179.400 511.050 180.450 ;
        RECT 508.950 178.950 511.050 179.400 ;
        RECT 514.950 178.950 517.050 180.750 ;
        RECT 526.950 178.950 529.050 180.750 ;
        RECT 313.950 175.950 316.050 178.050 ;
        RECT 331.950 176.250 334.050 178.050 ;
        RECT 337.950 176.250 340.050 178.050 ;
        RECT 352.950 176.250 355.050 178.050 ;
        RECT 358.950 176.250 361.050 178.050 ;
        RECT 364.950 177.450 367.050 178.050 ;
        RECT 376.950 177.450 379.050 178.050 ;
        RECT 364.950 176.400 379.050 177.450 ;
        RECT 364.950 175.950 367.050 176.400 ;
        RECT 376.950 175.950 379.050 176.400 ;
        RECT 412.950 176.250 415.050 178.050 ;
        RECT 418.950 176.250 421.050 178.050 ;
        RECT 436.950 176.250 439.050 178.050 ;
        RECT 475.950 175.950 478.050 178.050 ;
        RECT 493.950 176.250 496.050 178.050 ;
        RECT 499.950 176.250 502.050 178.050 ;
        RECT 511.950 176.250 514.050 178.050 ;
        RECT 517.950 176.250 520.050 178.050 ;
        RECT 331.950 172.950 334.050 175.050 ;
        RECT 337.950 172.950 340.050 175.050 ;
        RECT 352.950 169.950 355.050 175.050 ;
        RECT 358.950 172.950 361.050 175.050 ;
        RECT 412.950 172.950 415.050 175.050 ;
        RECT 418.950 172.950 421.050 175.050 ;
        RECT 430.950 174.450 435.000 175.050 ;
        RECT 436.950 174.450 439.050 175.050 ;
        RECT 430.950 173.400 439.050 174.450 ;
        RECT 430.950 172.950 435.000 173.400 ;
        RECT 436.950 172.950 439.050 173.400 ;
        RECT 493.950 172.950 496.050 175.050 ;
        RECT 499.950 174.450 502.050 175.050 ;
        RECT 504.000 174.450 508.050 175.050 ;
        RECT 499.950 173.400 508.050 174.450 ;
        RECT 499.950 172.950 502.050 173.400 ;
        RECT 504.000 172.950 508.050 173.400 ;
        RECT 511.950 172.950 514.050 175.050 ;
        RECT 517.950 172.950 520.050 175.050 ;
        RECT 530.850 173.400 532.050 188.400 ;
        RECT 544.950 179.250 547.050 181.050 ;
        RECT 544.950 175.950 547.050 178.050 ;
        RECT 529.950 171.300 532.050 173.400 ;
        RECT 190.950 166.950 193.050 167.400 ;
        RECT 259.950 166.950 262.050 167.400 ;
        RECT 265.950 166.950 268.050 167.400 ;
        RECT 214.950 165.450 217.050 166.050 ;
        RECT 289.950 165.600 292.050 167.700 ;
        RECT 310.950 166.500 313.050 168.600 ;
        RECT 316.950 168.450 319.050 169.050 ;
        RECT 316.950 167.400 336.450 168.450 ;
        RECT 530.850 167.700 532.050 171.300 ;
        RECT 551.100 168.600 552.300 188.400 ;
        RECT 637.950 187.950 640.050 188.400 ;
        RECT 667.950 187.950 670.050 188.400 ;
        RECT 722.400 188.400 730.050 189.450 ;
        RECT 613.950 184.950 616.050 187.050 ;
        RECT 619.950 184.950 622.050 187.050 ;
        RECT 679.950 184.950 682.050 187.050 ;
        RECT 685.950 184.950 688.050 187.050 ;
        RECT 703.950 184.950 706.050 187.050 ;
        RECT 709.950 186.450 712.050 187.050 ;
        RECT 722.400 186.450 723.450 188.400 ;
        RECT 727.950 187.950 730.050 188.400 ;
        RECT 760.950 189.450 763.050 190.050 ;
        RECT 769.950 189.450 772.050 190.050 ;
        RECT 760.950 188.400 772.050 189.450 ;
        RECT 760.950 187.950 763.050 188.400 ;
        RECT 769.950 187.950 772.050 188.400 ;
        RECT 775.950 189.450 778.050 190.050 ;
        RECT 781.950 189.450 784.050 190.050 ;
        RECT 775.950 188.400 784.050 189.450 ;
        RECT 775.950 187.950 778.050 188.400 ;
        RECT 781.950 187.950 784.050 188.400 ;
        RECT 788.400 187.050 789.450 191.400 ;
        RECT 820.950 190.950 823.050 191.400 ;
        RECT 877.950 190.950 880.050 191.400 ;
        RECT 883.950 190.950 886.050 194.400 ;
        RECT 814.950 189.450 817.050 190.050 ;
        RECT 832.950 189.450 835.050 190.050 ;
        RECT 814.950 188.400 835.050 189.450 ;
        RECT 814.950 187.950 817.050 188.400 ;
        RECT 709.950 185.400 723.450 186.450 ;
        RECT 709.950 184.950 712.050 185.400 ;
        RECT 787.950 184.950 790.050 187.050 ;
        RECT 793.950 184.950 796.050 187.050 ;
        RECT 827.400 186.450 828.450 188.400 ;
        RECT 832.950 187.950 835.050 188.400 ;
        RECT 889.950 189.450 892.050 190.050 ;
        RECT 901.950 189.450 904.050 190.050 ;
        RECT 889.950 188.400 904.050 189.450 ;
        RECT 889.950 187.950 892.050 188.400 ;
        RECT 901.950 187.950 904.050 188.400 ;
        RECT 817.950 185.400 828.450 186.450 ;
        RECT 574.950 181.950 577.050 184.050 ;
        RECT 586.950 181.950 592.050 184.050 ;
        RECT 595.950 181.950 598.050 184.050 ;
        RECT 613.950 181.950 616.050 183.750 ;
        RECT 619.950 181.950 622.050 183.750 ;
        RECT 637.950 181.950 640.050 184.050 ;
        RECT 658.950 181.950 661.050 184.050 ;
        RECT 664.950 183.450 667.050 184.050 ;
        RECT 673.950 183.450 676.050 184.050 ;
        RECT 664.950 182.400 676.050 183.450 ;
        RECT 664.950 181.950 667.050 182.400 ;
        RECT 673.950 181.950 676.050 182.400 ;
        RECT 679.950 181.950 682.050 183.750 ;
        RECT 685.950 181.950 688.050 183.750 ;
        RECT 703.950 181.950 706.050 183.750 ;
        RECT 709.950 181.950 712.050 183.750 ;
        RECT 727.950 181.950 730.050 184.050 ;
        RECT 751.950 181.950 754.050 184.050 ;
        RECT 769.950 181.950 772.050 184.050 ;
        RECT 775.950 181.950 778.050 184.050 ;
        RECT 787.950 181.950 790.050 183.750 ;
        RECT 793.950 181.950 796.050 183.750 ;
        RECT 802.950 183.450 805.050 184.050 ;
        RECT 811.950 183.450 814.050 184.050 ;
        RECT 802.950 182.400 814.050 183.450 ;
        RECT 802.950 181.950 805.050 182.400 ;
        RECT 811.950 181.950 814.050 182.400 ;
        RECT 817.950 181.950 820.050 185.400 ;
        RECT 871.950 184.950 874.050 187.050 ;
        RECT 877.950 184.950 880.050 187.050 ;
        RECT 832.950 181.950 835.050 184.050 ;
        RECT 841.950 183.450 844.050 184.050 ;
        RECT 850.950 183.450 853.050 184.050 ;
        RECT 841.950 182.400 853.050 183.450 ;
        RECT 841.950 181.950 844.050 182.400 ;
        RECT 850.950 181.950 853.050 182.400 ;
        RECT 871.950 181.950 874.050 183.750 ;
        RECT 877.950 181.950 880.050 183.750 ;
        RECT 895.950 181.950 898.050 184.050 ;
        RECT 553.950 179.250 556.050 181.050 ;
        RECT 574.950 178.950 577.050 180.750 ;
        RECT 589.950 178.950 592.050 180.750 ;
        RECT 595.950 178.950 598.050 180.750 ;
        RECT 616.950 179.250 619.050 181.050 ;
        RECT 634.950 180.750 636.750 181.050 ;
        RECT 634.950 179.250 637.050 180.750 ;
        RECT 637.950 179.250 640.050 180.750 ;
        RECT 643.950 179.250 646.050 181.050 ;
        RECT 638.250 178.950 640.050 179.250 ;
        RECT 658.950 178.950 661.050 180.750 ;
        RECT 664.950 178.950 667.050 180.750 ;
        RECT 682.950 179.250 685.050 181.050 ;
        RECT 706.950 179.250 709.050 181.050 ;
        RECT 721.950 179.250 724.050 181.050 ;
        RECT 731.250 180.750 733.050 181.050 ;
        RECT 727.950 179.250 730.050 180.750 ;
        RECT 730.950 179.250 733.050 180.750 ;
        RECT 727.950 178.950 729.750 179.250 ;
        RECT 751.950 178.950 754.050 180.750 ;
        RECT 769.950 178.950 772.050 180.750 ;
        RECT 775.950 178.950 778.050 180.750 ;
        RECT 790.950 179.250 793.050 181.050 ;
        RECT 811.950 178.950 814.050 180.750 ;
        RECT 817.950 178.950 820.050 180.750 ;
        RECT 832.950 178.950 835.050 180.750 ;
        RECT 850.950 178.950 853.050 180.750 ;
        RECT 874.950 179.250 877.050 181.050 ;
        RECT 895.950 178.950 898.050 180.750 ;
        RECT 553.950 175.950 556.050 178.050 ;
        RECT 571.950 176.250 574.050 178.050 ;
        RECT 592.950 176.250 595.050 178.050 ;
        RECT 598.950 176.250 601.050 178.050 ;
        RECT 616.950 175.950 621.900 178.050 ;
        RECT 623.100 177.450 625.200 178.050 ;
        RECT 634.950 177.450 637.050 178.050 ;
        RECT 623.100 176.400 637.050 177.450 ;
        RECT 623.100 175.950 625.200 176.400 ;
        RECT 634.950 175.950 637.050 176.400 ;
        RECT 643.950 175.950 646.050 178.050 ;
        RECT 655.950 176.250 658.050 178.050 ;
        RECT 661.950 176.250 664.050 178.050 ;
        RECT 667.950 177.450 670.050 178.050 ;
        RECT 682.950 177.450 685.050 178.050 ;
        RECT 700.950 177.450 703.050 178.050 ;
        RECT 667.950 176.400 703.050 177.450 ;
        RECT 667.950 175.950 670.050 176.400 ;
        RECT 682.950 175.950 685.050 176.400 ;
        RECT 700.950 175.950 703.050 176.400 ;
        RECT 706.950 175.950 712.050 178.050 ;
        RECT 721.950 175.950 724.050 178.050 ;
        RECT 571.950 169.950 574.050 175.050 ;
        RECT 592.950 172.950 595.050 175.050 ;
        RECT 598.950 174.450 601.050 175.050 ;
        RECT 610.950 174.450 613.050 175.050 ;
        RECT 598.950 173.400 613.050 174.450 ;
        RECT 598.950 172.950 601.050 173.400 ;
        RECT 610.950 172.950 613.050 173.400 ;
        RECT 655.950 172.950 658.050 175.050 ;
        RECT 661.950 172.950 664.050 175.050 ;
        RECT 730.950 172.950 733.050 178.050 ;
        RECT 748.950 176.250 751.050 178.050 ;
        RECT 766.950 176.250 769.050 178.050 ;
        RECT 772.950 176.250 775.050 178.050 ;
        RECT 781.950 177.450 784.050 178.050 ;
        RECT 790.950 177.450 793.050 178.050 ;
        RECT 781.950 176.400 793.050 177.450 ;
        RECT 781.950 175.950 784.050 176.400 ;
        RECT 790.950 175.950 793.050 176.400 ;
        RECT 814.950 176.250 817.050 178.050 ;
        RECT 820.950 176.250 823.050 178.050 ;
        RECT 835.950 176.250 838.050 178.050 ;
        RECT 853.950 176.250 856.050 178.050 ;
        RECT 868.950 177.450 873.000 178.050 ;
        RECT 874.950 177.450 877.050 178.050 ;
        RECT 868.950 176.400 877.050 177.450 ;
        RECT 868.950 175.950 873.000 176.400 ;
        RECT 874.950 175.950 877.050 176.400 ;
        RECT 892.950 176.250 895.050 178.050 ;
        RECT 748.950 172.950 751.050 175.050 ;
        RECT 766.950 172.950 769.050 175.050 ;
        RECT 772.950 172.950 775.050 175.050 ;
        RECT 796.950 174.450 799.050 175.050 ;
        RECT 814.950 174.450 817.050 175.050 ;
        RECT 796.950 173.400 817.050 174.450 ;
        RECT 796.950 172.950 799.050 173.400 ;
        RECT 814.950 172.950 817.050 173.400 ;
        RECT 820.950 172.950 823.050 175.050 ;
        RECT 826.950 174.450 829.050 175.050 ;
        RECT 835.950 174.450 838.050 175.050 ;
        RECT 826.950 173.400 838.050 174.450 ;
        RECT 826.950 172.950 829.050 173.400 ;
        RECT 835.950 172.950 838.050 173.400 ;
        RECT 853.950 172.950 856.050 175.050 ;
        RECT 889.950 172.950 895.050 175.050 ;
        RECT 673.950 171.450 676.050 172.050 ;
        RECT 721.950 171.450 724.050 172.050 ;
        RECT 673.950 170.400 724.050 171.450 ;
        RECT 673.950 169.950 676.050 170.400 ;
        RECT 721.950 169.950 724.050 170.400 ;
        RECT 316.950 166.950 319.050 167.400 ;
        RECT 67.950 164.400 94.050 165.450 ;
        RECT 67.950 163.950 70.050 164.400 ;
        RECT 91.950 163.950 94.050 164.400 ;
        RECT 194.400 164.400 217.050 165.450 ;
        RECT 335.400 165.450 336.450 167.400 ;
        RECT 364.950 165.450 367.050 166.050 ;
        RECT 335.400 164.400 367.050 165.450 ;
        RECT 88.950 162.450 91.050 163.050 ;
        RECT 194.400 162.450 195.450 164.400 ;
        RECT 214.950 163.950 217.050 164.400 ;
        RECT 364.950 163.950 367.050 164.400 ;
        RECT 505.950 165.450 508.050 166.050 ;
        RECT 520.950 165.450 523.050 166.050 ;
        RECT 529.950 165.600 532.050 167.700 ;
        RECT 550.950 166.500 553.050 168.600 ;
        RECT 592.950 168.450 595.050 169.050 ;
        RECT 601.950 168.450 604.050 169.050 ;
        RECT 592.950 167.400 604.050 168.450 ;
        RECT 592.950 166.950 595.050 167.400 ;
        RECT 601.950 166.950 604.050 167.400 ;
        RECT 610.950 168.450 613.050 169.050 ;
        RECT 655.950 168.450 658.050 169.050 ;
        RECT 610.950 167.400 658.050 168.450 ;
        RECT 610.950 166.950 613.050 167.400 ;
        RECT 655.950 166.950 658.050 167.400 ;
        RECT 766.950 168.450 769.050 169.050 ;
        RECT 781.950 168.450 784.050 169.050 ;
        RECT 766.950 167.400 784.050 168.450 ;
        RECT 766.950 166.950 769.050 167.400 ;
        RECT 781.950 166.950 784.050 167.400 ;
        RECT 832.950 168.450 835.050 169.050 ;
        RECT 854.400 168.450 855.450 172.950 ;
        RECT 832.950 167.400 855.450 168.450 ;
        RECT 832.950 166.950 835.050 167.400 ;
        RECT 505.950 164.400 523.050 165.450 ;
        RECT 505.950 163.950 508.050 164.400 ;
        RECT 520.950 163.950 523.050 164.400 ;
        RECT 589.950 165.450 592.050 166.050 ;
        RECT 595.950 165.450 598.050 166.050 ;
        RECT 622.950 165.450 625.050 166.050 ;
        RECT 589.950 164.400 625.050 165.450 ;
        RECT 589.950 163.950 592.050 164.400 ;
        RECT 595.950 163.950 598.050 164.400 ;
        RECT 622.950 163.950 625.050 164.400 ;
        RECT 649.950 165.450 652.050 166.050 ;
        RECT 661.950 165.450 664.050 166.050 ;
        RECT 649.950 164.400 664.050 165.450 ;
        RECT 649.950 163.950 652.050 164.400 ;
        RECT 661.950 163.950 664.050 164.400 ;
        RECT 88.950 161.400 195.450 162.450 ;
        RECT 310.950 162.450 313.050 163.050 ;
        RECT 319.950 162.450 322.050 163.050 ;
        RECT 310.950 161.400 322.050 162.450 ;
        RECT 88.950 160.950 91.050 161.400 ;
        RECT 310.950 160.950 313.050 161.400 ;
        RECT 319.950 160.950 322.050 161.400 ;
        RECT 367.950 162.450 370.050 163.050 ;
        RECT 481.950 162.450 484.050 163.050 ;
        RECT 367.950 161.400 484.050 162.450 ;
        RECT 367.950 160.950 370.050 161.400 ;
        RECT 481.950 160.950 484.050 161.400 ;
        RECT 505.950 162.450 508.050 163.050 ;
        RECT 526.950 162.450 529.050 163.050 ;
        RECT 505.950 161.400 529.050 162.450 ;
        RECT 505.950 160.950 508.050 161.400 ;
        RECT 526.950 160.950 529.050 161.400 ;
        RECT 580.950 162.450 583.050 163.050 ;
        RECT 736.950 162.450 739.050 163.050 ;
        RECT 580.950 161.400 739.050 162.450 ;
        RECT 580.950 160.950 583.050 161.400 ;
        RECT 736.950 160.950 739.050 161.400 ;
        RECT 748.950 162.450 751.050 163.050 ;
        RECT 772.950 162.450 775.050 163.050 ;
        RECT 808.950 162.450 811.050 163.050 ;
        RECT 748.950 161.400 811.050 162.450 ;
        RECT 748.950 160.950 751.050 161.400 ;
        RECT 772.950 160.950 775.050 161.400 ;
        RECT 808.950 160.950 811.050 161.400 ;
        RECT 814.950 162.450 817.050 163.050 ;
        RECT 829.950 162.450 832.050 163.050 ;
        RECT 814.950 161.400 832.050 162.450 ;
        RECT 814.950 160.950 817.050 161.400 ;
        RECT 829.950 160.950 832.050 161.400 ;
        RECT 91.950 159.450 94.050 160.050 ;
        RECT 172.950 159.450 175.050 160.050 ;
        RECT 205.950 159.450 208.050 160.050 ;
        RECT 91.950 158.400 208.050 159.450 ;
        RECT 91.950 157.950 94.050 158.400 ;
        RECT 172.950 157.950 175.050 158.400 ;
        RECT 205.950 157.950 208.050 158.400 ;
        RECT 226.950 159.450 229.050 160.050 ;
        RECT 274.950 159.450 277.050 160.050 ;
        RECT 319.800 159.450 321.900 160.200 ;
        RECT 226.950 158.400 267.450 159.450 ;
        RECT 226.950 157.950 229.050 158.400 ;
        RECT 266.400 157.050 267.450 158.400 ;
        RECT 274.950 158.400 321.900 159.450 ;
        RECT 274.950 157.950 277.050 158.400 ;
        RECT 319.800 158.100 321.900 158.400 ;
        RECT 323.100 159.450 325.200 160.050 ;
        RECT 328.950 159.450 331.050 160.050 ;
        RECT 355.950 159.450 358.050 160.050 ;
        RECT 323.100 158.400 358.050 159.450 ;
        RECT 323.100 157.950 325.200 158.400 ;
        RECT 328.950 157.950 331.050 158.400 ;
        RECT 355.950 157.950 358.050 158.400 ;
        RECT 406.950 159.450 409.050 160.050 ;
        RECT 418.950 159.450 421.050 160.050 ;
        RECT 506.400 159.450 507.450 160.950 ;
        RECT 406.950 158.400 507.450 159.450 ;
        RECT 520.950 159.450 523.050 160.050 ;
        RECT 544.950 159.450 547.050 160.050 ;
        RECT 520.950 158.400 547.050 159.450 ;
        RECT 406.950 157.950 409.050 158.400 ;
        RECT 418.950 157.950 421.050 158.400 ;
        RECT 520.950 157.950 523.050 158.400 ;
        RECT 544.950 157.950 547.050 158.400 ;
        RECT 685.950 159.450 688.050 160.050 ;
        RECT 784.950 159.450 787.050 160.050 ;
        RECT 685.950 158.400 787.050 159.450 ;
        RECT 685.950 157.950 688.050 158.400 ;
        RECT 784.950 157.950 787.050 158.400 ;
        RECT 13.950 156.450 16.050 157.050 ;
        RECT 37.950 156.450 40.050 157.050 ;
        RECT 79.950 156.450 82.050 157.050 ;
        RECT 13.950 155.400 30.450 156.450 ;
        RECT 13.950 154.950 16.050 155.400 ;
        RECT 16.950 153.450 19.050 154.050 ;
        RECT 22.950 153.450 25.050 154.050 ;
        RECT 16.950 152.400 25.050 153.450 ;
        RECT 16.950 151.950 19.050 152.400 ;
        RECT 22.950 151.950 25.050 152.400 ;
        RECT 29.400 150.450 30.450 155.400 ;
        RECT 37.950 155.400 82.050 156.450 ;
        RECT 37.950 154.950 40.050 155.400 ;
        RECT 79.950 154.950 82.050 155.400 ;
        RECT 115.950 156.450 118.050 157.050 ;
        RECT 160.950 156.450 163.050 157.050 ;
        RECT 184.950 156.450 187.050 157.050 ;
        RECT 190.950 156.450 193.050 157.050 ;
        RECT 115.950 155.400 193.050 156.450 ;
        RECT 115.950 154.950 118.050 155.400 ;
        RECT 160.950 154.950 163.050 155.400 ;
        RECT 184.950 154.950 187.050 155.400 ;
        RECT 190.950 154.950 193.050 155.400 ;
        RECT 196.950 156.450 199.050 157.050 ;
        RECT 238.950 156.450 241.050 157.050 ;
        RECT 196.950 155.400 241.050 156.450 ;
        RECT 196.950 154.950 199.050 155.400 ;
        RECT 238.950 154.950 241.050 155.400 ;
        RECT 265.950 156.450 268.050 157.050 ;
        RECT 301.950 156.450 304.050 157.050 ;
        RECT 316.800 156.450 318.900 157.050 ;
        RECT 265.950 155.400 318.900 156.450 ;
        RECT 265.950 154.950 268.050 155.400 ;
        RECT 301.950 154.950 304.050 155.400 ;
        RECT 316.800 154.950 318.900 155.400 ;
        RECT 320.100 156.450 322.200 156.900 ;
        RECT 346.950 156.450 349.050 157.050 ;
        RECT 320.100 155.400 349.050 156.450 ;
        RECT 320.100 154.800 322.200 155.400 ;
        RECT 346.950 154.950 349.050 155.400 ;
        RECT 358.950 156.450 361.050 157.050 ;
        RECT 373.950 156.450 376.050 157.050 ;
        RECT 472.950 156.450 475.050 157.050 ;
        RECT 358.950 155.400 475.050 156.450 ;
        RECT 358.950 154.950 361.050 155.400 ;
        RECT 373.950 154.950 376.050 155.400 ;
        RECT 472.950 154.950 475.050 155.400 ;
        RECT 493.950 156.450 496.050 157.050 ;
        RECT 502.950 156.450 505.050 157.050 ;
        RECT 493.950 155.400 505.050 156.450 ;
        RECT 493.950 154.950 496.050 155.400 ;
        RECT 502.950 154.950 505.050 155.400 ;
        RECT 640.950 156.450 643.050 157.050 ;
        RECT 676.950 156.450 679.050 157.050 ;
        RECT 640.950 155.400 679.050 156.450 ;
        RECT 640.950 154.950 643.050 155.400 ;
        RECT 676.950 154.950 679.050 155.400 ;
        RECT 31.950 153.450 34.050 154.050 ;
        RECT 40.950 153.450 43.050 154.050 ;
        RECT 31.950 152.400 43.050 153.450 ;
        RECT 31.950 151.950 34.050 152.400 ;
        RECT 40.950 151.950 43.050 152.400 ;
        RECT 46.950 153.450 49.050 154.050 ;
        RECT 73.950 153.450 76.050 154.050 ;
        RECT 46.950 152.400 76.050 153.450 ;
        RECT 46.950 151.950 49.050 152.400 ;
        RECT 73.950 151.950 76.050 152.400 ;
        RECT 34.950 150.450 37.050 151.050 ;
        RECT 29.400 149.400 37.050 150.450 ;
        RECT 34.950 148.950 37.050 149.400 ;
        RECT 94.950 148.950 97.050 154.050 ;
        RECT 124.950 153.450 127.050 154.050 ;
        RECT 286.950 153.450 289.050 154.050 ;
        RECT 124.950 152.400 289.050 153.450 ;
        RECT 124.950 151.950 127.050 152.400 ;
        RECT 286.950 151.950 289.050 152.400 ;
        RECT 292.950 153.450 295.050 154.050 ;
        RECT 304.950 153.450 307.050 154.050 ;
        RECT 292.950 152.400 307.050 153.450 ;
        RECT 292.950 151.950 295.050 152.400 ;
        RECT 304.950 151.950 307.050 152.400 ;
        RECT 337.950 153.450 340.050 154.050 ;
        RECT 352.950 153.450 355.050 154.050 ;
        RECT 337.950 152.400 355.050 153.450 ;
        RECT 337.950 151.950 340.050 152.400 ;
        RECT 352.950 151.950 355.050 152.400 ;
        RECT 439.950 153.450 442.050 154.050 ;
        RECT 475.950 153.450 478.050 154.050 ;
        RECT 439.950 152.400 478.050 153.450 ;
        RECT 439.950 151.950 442.050 152.400 ;
        RECT 475.950 151.950 478.050 152.400 ;
        RECT 487.950 153.450 490.050 154.050 ;
        RECT 565.950 153.450 568.050 154.050 ;
        RECT 607.950 153.450 610.050 154.050 ;
        RECT 487.950 152.400 610.050 153.450 ;
        RECT 487.950 151.950 490.050 152.400 ;
        RECT 565.950 151.950 568.050 152.400 ;
        RECT 607.950 151.950 610.050 152.400 ;
        RECT 646.950 153.450 649.050 154.050 ;
        RECT 724.950 153.450 727.050 154.050 ;
        RECT 730.950 153.450 733.050 154.050 ;
        RECT 646.950 152.400 705.450 153.450 ;
        RECT 646.950 151.950 649.050 152.400 ;
        RECT 704.400 151.050 705.450 152.400 ;
        RECT 724.950 152.400 733.050 153.450 ;
        RECT 724.950 151.950 727.050 152.400 ;
        RECT 730.950 151.950 733.050 152.400 ;
        RECT 343.950 150.450 346.050 151.050 ;
        RECT 349.950 150.450 352.050 151.050 ;
        RECT 343.950 149.400 352.050 150.450 ;
        RECT 22.950 147.450 25.050 148.050 ;
        RECT 40.950 147.450 43.050 148.050 ;
        RECT 46.800 147.450 48.900 148.050 ;
        RECT 22.950 146.400 48.900 147.450 ;
        RECT 22.950 145.950 25.050 146.400 ;
        RECT 40.950 145.950 43.050 146.400 ;
        RECT 46.800 145.950 48.900 146.400 ;
        RECT 50.100 147.450 52.200 148.050 ;
        RECT 55.950 147.450 58.050 148.050 ;
        RECT 50.100 146.400 58.050 147.450 ;
        RECT 50.100 145.950 52.200 146.400 ;
        RECT 55.950 145.950 58.050 146.400 ;
        RECT 73.950 147.450 76.050 148.050 ;
        RECT 103.950 147.450 106.050 148.050 ;
        RECT 73.950 146.400 106.050 147.450 ;
        RECT 73.950 145.950 76.050 146.400 ;
        RECT 103.950 145.950 106.050 146.400 ;
        RECT 175.950 147.450 178.050 148.050 ;
        RECT 187.950 147.450 190.050 148.050 ;
        RECT 175.950 146.400 190.050 147.450 ;
        RECT 232.950 146.400 235.050 148.500 ;
        RECT 253.950 147.300 256.050 149.400 ;
        RECT 175.950 145.950 178.050 146.400 ;
        RECT 187.950 145.950 190.050 146.400 ;
        RECT 94.950 144.450 97.050 145.050 ;
        RECT 94.950 143.400 132.450 144.450 ;
        RECT 94.950 142.950 97.050 143.400 ;
        RECT 16.950 139.950 19.050 142.050 ;
        RECT 22.950 139.950 25.050 142.050 ;
        RECT 34.950 139.950 37.050 142.050 ;
        RECT 40.950 139.950 43.050 142.050 ;
        RECT 55.950 139.950 58.050 142.050 ;
        RECT 61.950 139.950 64.050 142.050 ;
        RECT 73.950 141.450 78.000 142.050 ;
        RECT 79.950 141.450 82.050 142.050 ;
        RECT 73.950 140.400 82.050 141.450 ;
        RECT 73.950 139.950 78.000 140.400 ;
        RECT 79.950 139.950 82.050 140.400 ;
        RECT 85.950 139.950 88.050 142.050 ;
        RECT 131.400 139.050 132.450 143.400 ;
        RECT 172.950 139.950 175.050 142.050 ;
        RECT 190.950 139.950 193.050 142.050 ;
        RECT 196.950 139.950 199.050 142.050 ;
        RECT 214.950 139.950 217.050 142.050 ;
        RECT 220.950 139.950 223.050 142.050 ;
        RECT 16.950 136.950 19.050 138.750 ;
        RECT 22.950 136.950 25.050 138.750 ;
        RECT 34.950 136.950 37.050 138.750 ;
        RECT 40.950 136.950 43.050 138.750 ;
        RECT 55.950 136.950 58.050 138.750 ;
        RECT 61.950 136.950 64.050 138.750 ;
        RECT 79.950 136.950 82.050 138.750 ;
        RECT 85.950 136.950 88.050 138.750 ;
        RECT 103.950 136.950 106.050 139.050 ;
        RECT 112.950 138.450 115.050 139.050 ;
        RECT 124.950 138.450 127.050 139.050 ;
        RECT 112.950 137.400 127.050 138.450 ;
        RECT 112.950 136.950 115.050 137.400 ;
        RECT 124.950 136.950 127.050 137.400 ;
        RECT 130.950 136.950 133.050 139.050 ;
        RECT 139.950 138.450 142.050 139.050 ;
        RECT 154.950 138.450 157.050 139.050 ;
        RECT 139.950 137.400 157.050 138.450 ;
        RECT 139.950 136.950 142.050 137.400 ;
        RECT 154.950 136.950 157.050 137.400 ;
        RECT 172.950 136.950 175.050 138.750 ;
        RECT 190.950 136.950 193.050 138.750 ;
        RECT 196.950 136.950 199.050 138.750 ;
        RECT 214.950 136.950 217.050 138.750 ;
        RECT 220.950 136.950 223.050 138.750 ;
        RECT 229.950 136.950 232.050 139.050 ;
        RECT 13.950 134.250 16.050 136.050 ;
        RECT 19.950 134.250 22.050 136.050 ;
        RECT 37.950 134.250 40.050 136.050 ;
        RECT 58.950 134.250 61.050 136.050 ;
        RECT 64.950 134.250 67.050 136.050 ;
        RECT 82.950 134.250 85.050 136.050 ;
        RECT 88.950 134.250 91.050 136.050 ;
        RECT 109.950 135.750 111.750 136.050 ;
        RECT 103.950 133.950 106.050 135.750 ;
        RECT 109.950 134.250 112.050 135.750 ;
        RECT 112.950 134.250 115.050 135.750 ;
        RECT 113.250 133.950 115.050 134.250 ;
        RECT 130.950 133.950 133.050 135.750 ;
        RECT 154.950 133.950 157.050 135.750 ;
        RECT 169.950 134.250 172.050 136.050 ;
        RECT 187.950 134.250 190.050 136.050 ;
        RECT 193.950 134.250 196.050 136.050 ;
        RECT 211.950 134.250 214.050 136.050 ;
        RECT 217.950 134.250 220.050 136.050 ;
        RECT 229.950 133.950 232.050 135.750 ;
        RECT 13.950 127.950 16.050 133.050 ;
        RECT 19.950 130.950 22.050 133.050 ;
        RECT 37.950 132.450 40.050 133.050 ;
        RECT 46.950 132.450 49.050 133.050 ;
        RECT 37.950 131.400 49.050 132.450 ;
        RECT 37.950 130.950 40.050 131.400 ;
        RECT 46.950 130.950 49.050 131.400 ;
        RECT 58.950 130.950 61.050 133.050 ;
        RECT 64.950 132.450 67.050 133.050 ;
        RECT 73.950 132.450 76.050 133.050 ;
        RECT 64.950 131.400 76.050 132.450 ;
        RECT 64.950 130.950 67.050 131.400 ;
        RECT 73.950 130.950 76.050 131.400 ;
        RECT 82.950 130.950 85.050 133.050 ;
        RECT 88.950 132.450 91.050 133.050 ;
        RECT 100.950 132.450 103.050 133.050 ;
        RECT 88.950 131.400 103.050 132.450 ;
        RECT 88.950 130.950 91.050 131.400 ;
        RECT 100.950 130.950 103.050 131.400 ;
        RECT 109.950 130.950 112.050 133.050 ;
        RECT 127.950 131.250 130.050 133.050 ;
        RECT 133.950 131.250 136.050 133.050 ;
        RECT 151.950 131.250 154.050 133.050 ;
        RECT 157.950 131.250 160.050 133.050 ;
        RECT 169.950 130.950 172.050 133.050 ;
        RECT 187.950 130.950 190.050 133.050 ;
        RECT 193.950 130.950 196.050 133.050 ;
        RECT 211.950 130.950 214.050 133.050 ;
        RECT 217.950 132.450 220.050 133.050 ;
        RECT 217.950 131.400 228.450 132.450 ;
        RECT 217.950 130.950 220.050 131.400 ;
        RECT 227.400 130.050 228.450 131.400 ;
        RECT 46.950 129.450 49.050 130.050 ;
        RECT 55.950 129.450 58.050 130.050 ;
        RECT 46.950 128.400 58.050 129.450 ;
        RECT 46.950 127.950 49.050 128.400 ;
        RECT 55.950 127.950 58.050 128.400 ;
        RECT 124.950 127.950 130.050 130.050 ;
        RECT 133.950 127.950 136.050 130.050 ;
        RECT 151.950 127.950 154.050 130.050 ;
        RECT 157.950 127.950 163.050 130.050 ;
        RECT 227.400 128.400 232.050 130.050 ;
        RECT 228.000 127.950 232.050 128.400 ;
        RECT 37.950 126.450 40.050 127.050 ;
        RECT 49.950 126.450 52.050 127.050 ;
        RECT 37.950 125.400 52.050 126.450 ;
        RECT 37.950 124.950 40.050 125.400 ;
        RECT 49.950 124.950 52.050 125.400 ;
        RECT 58.950 126.450 61.050 127.050 ;
        RECT 82.950 126.450 85.050 127.050 ;
        RECT 58.950 125.400 85.050 126.450 ;
        RECT 58.950 124.950 61.050 125.400 ;
        RECT 82.950 124.950 85.050 125.400 ;
        RECT 88.950 126.450 91.050 127.050 ;
        RECT 97.950 126.450 100.050 127.050 ;
        RECT 88.950 125.400 100.050 126.450 ;
        RECT 88.950 124.950 91.050 125.400 ;
        RECT 97.950 124.950 100.050 125.400 ;
        RECT 175.950 126.450 178.050 127.050 ;
        RECT 187.950 126.450 190.050 127.050 ;
        RECT 233.700 126.600 234.900 146.400 ;
        RECT 253.950 143.700 255.150 147.300 ;
        RECT 268.950 146.400 271.050 148.500 ;
        RECT 289.950 147.300 292.050 149.400 ;
        RECT 253.950 141.600 256.050 143.700 ;
        RECT 238.950 136.950 241.050 139.050 ;
        RECT 238.950 133.950 241.050 135.750 ;
        RECT 253.950 126.600 255.150 141.600 ;
        RECT 265.950 136.950 268.050 139.050 ;
        RECT 256.950 134.250 259.050 136.050 ;
        RECT 265.950 133.950 268.050 135.750 ;
        RECT 256.950 130.950 259.050 133.050 ;
        RECT 269.700 126.600 270.900 146.400 ;
        RECT 289.950 143.700 291.150 147.300 ;
        RECT 304.950 146.400 307.050 148.500 ;
        RECT 325.950 147.300 328.050 149.400 ;
        RECT 343.950 148.950 346.050 149.400 ;
        RECT 349.950 148.950 352.050 149.400 ;
        RECT 400.950 150.450 403.050 151.050 ;
        RECT 409.950 150.450 412.050 151.050 ;
        RECT 400.950 149.400 412.050 150.450 ;
        RECT 400.950 148.950 403.050 149.400 ;
        RECT 409.950 148.950 412.050 149.400 ;
        RECT 466.950 150.450 469.050 151.050 ;
        RECT 514.950 150.450 517.050 151.050 ;
        RECT 466.950 149.400 517.050 150.450 ;
        RECT 466.950 148.950 469.050 149.400 ;
        RECT 514.950 148.950 517.050 149.400 ;
        RECT 520.950 150.450 523.050 151.050 ;
        RECT 526.950 150.450 529.050 151.050 ;
        RECT 520.950 149.400 529.050 150.450 ;
        RECT 520.950 148.950 523.050 149.400 ;
        RECT 526.950 148.950 529.050 149.400 ;
        RECT 544.950 150.450 547.050 151.050 ;
        RECT 601.950 150.450 604.050 151.050 ;
        RECT 544.950 149.400 604.050 150.450 ;
        RECT 703.950 150.450 706.050 151.050 ;
        RECT 712.950 150.450 715.050 151.050 ;
        RECT 748.950 150.450 751.050 151.050 ;
        RECT 703.950 149.400 751.050 150.450 ;
        RECT 544.950 148.950 547.050 149.400 ;
        RECT 601.950 148.950 604.050 149.400 ;
        RECT 331.950 147.450 334.050 148.050 ;
        RECT 364.950 147.450 367.050 148.050 ;
        RECT 412.950 147.450 415.050 148.050 ;
        RECT 289.950 141.600 292.050 143.700 ;
        RECT 274.950 136.950 277.050 139.050 ;
        RECT 274.950 133.950 277.050 135.750 ;
        RECT 289.950 126.600 291.150 141.600 ;
        RECT 301.950 136.950 304.050 139.050 ;
        RECT 292.950 134.250 295.050 136.050 ;
        RECT 301.950 133.950 304.050 135.750 ;
        RECT 292.950 130.950 295.050 133.050 ;
        RECT 305.700 126.600 306.900 146.400 ;
        RECT 325.950 143.700 327.150 147.300 ;
        RECT 331.950 146.400 415.050 147.450 ;
        RECT 331.950 145.950 334.050 146.400 ;
        RECT 364.950 145.950 367.050 146.400 ;
        RECT 412.950 145.950 415.050 146.400 ;
        RECT 439.950 147.450 442.050 148.050 ;
        RECT 445.950 147.450 448.050 148.050 ;
        RECT 439.950 146.400 448.050 147.450 ;
        RECT 439.950 145.950 442.050 146.400 ;
        RECT 445.950 145.950 448.050 146.400 ;
        RECT 478.950 147.450 481.050 148.050 ;
        RECT 487.950 147.450 490.050 148.050 ;
        RECT 478.950 146.400 490.050 147.450 ;
        RECT 478.950 145.950 481.050 146.400 ;
        RECT 487.950 145.950 490.050 146.400 ;
        RECT 508.950 147.450 511.050 148.050 ;
        RECT 538.950 147.450 541.050 148.050 ;
        RECT 583.950 147.450 586.050 148.050 ;
        RECT 508.950 146.400 586.050 147.450 ;
        RECT 661.950 147.300 664.050 149.400 ;
        RECT 703.950 148.950 706.050 149.400 ;
        RECT 712.950 148.950 715.050 149.400 ;
        RECT 748.950 148.950 751.050 149.400 ;
        RECT 508.950 145.950 511.050 146.400 ;
        RECT 538.950 145.950 541.050 146.400 ;
        RECT 583.950 145.950 586.050 146.400 ;
        RECT 394.950 144.450 397.050 145.050 ;
        RECT 415.800 144.450 417.900 145.050 ;
        RECT 325.950 141.600 328.050 143.700 ;
        RECT 394.950 143.400 417.900 144.450 ;
        RECT 394.950 142.950 397.050 143.400 ;
        RECT 415.800 142.950 417.900 143.400 ;
        RECT 419.100 144.450 421.200 145.050 ;
        RECT 424.950 144.450 427.050 145.050 ;
        RECT 436.950 144.450 439.050 145.050 ;
        RECT 419.100 143.400 439.050 144.450 ;
        RECT 662.850 143.700 664.050 147.300 ;
        RECT 682.950 146.400 685.050 148.500 ;
        RECT 730.950 147.450 733.050 148.050 ;
        RECT 742.950 147.450 745.050 148.050 ;
        RECT 775.950 147.450 778.050 148.050 ;
        RECT 793.950 147.450 796.050 148.050 ;
        RECT 730.950 146.400 796.050 147.450 ;
        RECT 419.100 142.950 421.200 143.400 ;
        RECT 424.950 142.950 427.050 143.400 ;
        RECT 436.950 142.950 439.050 143.400 ;
        RECT 310.950 138.450 313.050 139.050 ;
        RECT 319.950 138.450 322.050 139.050 ;
        RECT 310.950 137.400 322.050 138.450 ;
        RECT 310.950 136.950 313.050 137.400 ;
        RECT 319.950 136.950 322.050 137.400 ;
        RECT 310.950 133.950 313.050 135.750 ;
        RECT 325.950 126.600 327.150 141.600 ;
        RECT 346.950 139.950 349.050 142.050 ;
        RECT 352.950 141.450 355.050 142.050 ;
        RECT 370.950 141.450 373.050 142.050 ;
        RECT 352.950 140.400 373.050 141.450 ;
        RECT 352.950 139.950 355.050 140.400 ;
        RECT 370.950 139.950 373.050 140.400 ;
        RECT 379.950 141.450 382.050 142.050 ;
        RECT 388.950 141.450 391.050 142.050 ;
        RECT 379.950 140.400 391.050 141.450 ;
        RECT 379.950 139.950 382.050 140.400 ;
        RECT 388.950 139.950 391.050 140.400 ;
        RECT 445.950 139.950 448.050 142.050 ;
        RECT 451.950 139.950 454.050 142.050 ;
        RECT 472.950 139.950 475.050 142.050 ;
        RECT 478.950 139.950 481.050 142.050 ;
        RECT 514.950 139.950 517.050 142.050 ;
        RECT 520.950 139.950 523.050 142.050 ;
        RECT 538.950 139.950 541.050 142.050 ;
        RECT 544.950 139.950 547.050 142.050 ;
        RECT 559.950 139.950 562.050 142.050 ;
        RECT 565.950 139.950 568.050 142.050 ;
        RECT 583.950 139.950 586.050 142.050 ;
        RECT 589.950 139.950 592.050 142.050 ;
        RECT 598.950 141.450 603.000 142.050 ;
        RECT 604.950 141.450 607.050 142.050 ;
        RECT 598.950 140.400 607.050 141.450 ;
        RECT 598.950 139.950 603.000 140.400 ;
        RECT 604.950 139.950 607.050 140.400 ;
        RECT 622.950 139.950 625.050 142.050 ;
        RECT 628.950 139.950 631.050 142.050 ;
        RECT 646.950 139.950 649.050 142.050 ;
        RECT 652.950 139.950 658.050 142.050 ;
        RECT 661.950 141.600 664.050 143.700 ;
        RECT 346.950 136.950 349.050 138.750 ;
        RECT 352.950 136.950 355.050 138.750 ;
        RECT 370.950 136.950 373.050 138.750 ;
        RECT 388.950 136.950 391.050 138.750 ;
        RECT 403.950 138.450 408.000 139.050 ;
        RECT 409.950 138.450 412.050 139.050 ;
        RECT 403.950 137.400 412.050 138.450 ;
        RECT 403.950 136.950 408.000 137.400 ;
        RECT 409.950 136.950 412.050 137.400 ;
        RECT 415.950 138.450 418.050 139.050 ;
        RECT 427.950 138.450 430.050 139.050 ;
        RECT 439.950 138.450 442.050 139.050 ;
        RECT 415.950 137.400 442.050 138.450 ;
        RECT 415.950 136.950 418.050 137.400 ;
        RECT 427.950 136.950 430.050 137.400 ;
        RECT 439.950 136.950 442.050 137.400 ;
        RECT 445.950 136.950 448.050 138.750 ;
        RECT 451.950 136.950 454.050 138.750 ;
        RECT 472.950 136.950 475.050 138.750 ;
        RECT 478.950 136.950 481.050 138.750 ;
        RECT 496.950 138.450 499.050 139.050 ;
        RECT 508.950 138.450 511.050 139.050 ;
        RECT 496.950 137.400 511.050 138.450 ;
        RECT 496.950 136.950 499.050 137.400 ;
        RECT 508.950 136.950 511.050 137.400 ;
        RECT 514.950 136.950 517.050 138.750 ;
        RECT 520.950 136.950 523.050 138.750 ;
        RECT 538.950 136.950 541.050 138.750 ;
        RECT 544.950 136.950 547.050 138.750 ;
        RECT 559.950 136.950 562.050 138.750 ;
        RECT 565.950 136.950 568.050 138.750 ;
        RECT 583.950 136.950 586.050 138.750 ;
        RECT 589.950 136.950 592.050 138.750 ;
        RECT 604.950 136.950 607.050 138.750 ;
        RECT 622.950 136.950 625.050 138.750 ;
        RECT 628.950 136.950 631.050 138.750 ;
        RECT 646.950 136.950 649.050 138.750 ;
        RECT 652.950 136.950 655.050 138.750 ;
        RECT 328.950 134.250 331.050 136.050 ;
        RECT 349.950 134.250 352.050 136.050 ;
        RECT 355.950 134.250 358.050 136.050 ;
        RECT 367.950 134.250 370.050 136.050 ;
        RECT 391.950 134.250 394.050 136.050 ;
        RECT 409.950 133.950 412.050 135.750 ;
        RECT 427.950 133.950 430.050 135.750 ;
        RECT 448.950 134.250 451.050 136.050 ;
        RECT 454.950 134.250 457.050 136.050 ;
        RECT 475.950 134.250 478.050 136.050 ;
        RECT 481.950 134.250 484.050 136.050 ;
        RECT 496.950 133.950 499.050 135.750 ;
        RECT 517.950 134.250 520.050 136.050 ;
        RECT 541.950 134.250 544.050 136.050 ;
        RECT 562.950 134.250 565.050 136.050 ;
        RECT 568.950 134.250 571.050 136.050 ;
        RECT 586.950 134.250 589.050 136.050 ;
        RECT 607.950 134.250 610.050 136.050 ;
        RECT 619.950 134.250 622.050 136.050 ;
        RECT 625.950 134.250 628.050 136.050 ;
        RECT 649.950 134.250 652.050 136.050 ;
        RECT 658.950 134.250 661.050 136.050 ;
        RECT 328.950 130.950 331.050 133.050 ;
        RECT 349.950 130.950 352.050 133.050 ;
        RECT 355.950 130.950 358.050 133.050 ;
        RECT 367.950 130.950 370.050 133.050 ;
        RECT 391.950 130.950 394.050 133.050 ;
        RECT 406.950 131.250 409.050 133.050 ;
        RECT 412.950 131.250 415.050 133.050 ;
        RECT 424.950 131.250 427.050 133.050 ;
        RECT 430.950 131.250 433.050 133.050 ;
        RECT 448.950 130.950 451.050 133.050 ;
        RECT 454.950 132.450 457.050 133.050 ;
        RECT 466.800 132.450 468.900 133.050 ;
        RECT 454.950 131.400 468.900 132.450 ;
        RECT 454.950 130.950 457.050 131.400 ;
        RECT 466.800 130.950 468.900 131.400 ;
        RECT 470.100 132.450 474.000 133.050 ;
        RECT 475.950 132.450 478.050 133.050 ;
        RECT 470.100 131.400 478.050 132.450 ;
        RECT 470.100 130.950 474.000 131.400 ;
        RECT 475.950 130.950 478.050 131.400 ;
        RECT 481.950 130.950 484.050 133.050 ;
        RECT 493.950 131.250 496.050 133.050 ;
        RECT 499.950 131.250 502.050 133.050 ;
        RECT 517.950 132.450 520.050 133.050 ;
        RECT 522.000 132.450 525.900 133.050 ;
        RECT 517.950 131.400 525.900 132.450 ;
        RECT 517.950 130.950 520.050 131.400 ;
        RECT 522.000 130.950 525.900 131.400 ;
        RECT 527.100 132.450 529.200 133.050 ;
        RECT 541.950 132.450 544.050 133.050 ;
        RECT 527.100 131.400 544.050 132.450 ;
        RECT 527.100 130.950 529.200 131.400 ;
        RECT 541.950 130.950 544.050 131.400 ;
        RECT 562.950 130.950 565.050 133.050 ;
        RECT 568.950 130.950 571.050 133.050 ;
        RECT 586.950 132.450 589.050 133.050 ;
        RECT 601.950 132.450 604.050 133.050 ;
        RECT 586.950 131.400 604.050 132.450 ;
        RECT 586.950 130.950 589.050 131.400 ;
        RECT 601.950 130.950 604.050 131.400 ;
        RECT 607.950 130.950 610.050 133.050 ;
        RECT 619.950 130.950 622.050 133.050 ;
        RECT 625.950 130.950 628.050 133.050 ;
        RECT 631.950 132.450 634.050 133.050 ;
        RECT 649.950 132.450 652.050 133.050 ;
        RECT 631.950 131.400 652.050 132.450 ;
        RECT 631.950 130.950 634.050 131.400 ;
        RECT 649.950 130.950 652.050 131.400 ;
        RECT 658.950 130.950 661.050 133.050 ;
        RECT 406.950 127.950 409.050 130.050 ;
        RECT 412.950 127.950 415.050 130.050 ;
        RECT 424.950 127.950 427.050 130.050 ;
        RECT 430.950 127.950 433.050 130.050 ;
        RECT 493.950 127.950 496.050 130.050 ;
        RECT 499.950 127.950 502.050 130.050 ;
        RECT 175.950 125.400 190.050 126.450 ;
        RECT 175.950 124.950 178.050 125.400 ;
        RECT 187.950 124.950 190.050 125.400 ;
        RECT 232.950 124.500 235.050 126.600 ;
        RECT 253.950 124.500 256.050 126.600 ;
        RECT 268.950 124.500 271.050 126.600 ;
        RECT 289.950 124.500 292.050 126.600 ;
        RECT 304.950 124.500 307.050 126.600 ;
        RECT 325.950 124.500 328.050 126.600 ;
        RECT 361.950 126.450 364.050 127.050 ;
        RECT 370.950 126.450 373.050 127.200 ;
        RECT 361.950 125.400 373.050 126.450 ;
        RECT 361.950 124.950 364.050 125.400 ;
        RECT 370.950 125.100 373.050 125.400 ;
        RECT 436.950 126.450 439.050 127.050 ;
        RECT 448.950 126.450 451.050 127.050 ;
        RECT 436.950 125.400 451.050 126.450 ;
        RECT 436.950 124.950 439.050 125.400 ;
        RECT 448.950 124.950 451.050 125.400 ;
        RECT 508.950 126.450 511.050 127.050 ;
        RECT 553.950 126.450 556.050 127.050 ;
        RECT 508.950 125.400 556.050 126.450 ;
        RECT 563.400 126.450 564.450 130.950 ;
        RECT 619.950 126.450 622.050 127.050 ;
        RECT 563.400 125.400 622.050 126.450 ;
        RECT 626.400 126.450 627.450 130.950 ;
        RECT 640.950 126.450 643.050 127.050 ;
        RECT 662.850 126.600 664.050 141.600 ;
        RECT 676.950 136.950 679.050 139.050 ;
        RECT 676.950 133.950 679.050 135.750 ;
        RECT 683.100 126.600 684.300 146.400 ;
        RECT 730.950 145.950 733.050 146.400 ;
        RECT 742.950 145.950 745.050 146.400 ;
        RECT 775.950 145.950 778.050 146.400 ;
        RECT 793.950 145.950 796.050 146.400 ;
        RECT 778.950 144.450 781.050 145.050 ;
        RECT 784.950 144.450 787.050 145.050 ;
        RECT 778.950 143.400 787.050 144.450 ;
        RECT 778.950 142.950 781.050 143.400 ;
        RECT 784.950 142.950 787.050 143.400 ;
        RECT 685.950 136.950 688.050 139.050 ;
        RECT 703.950 136.950 706.050 142.050 ;
        RECT 709.950 141.450 712.050 142.050 ;
        RECT 718.950 141.450 721.050 142.050 ;
        RECT 709.950 140.400 721.050 141.450 ;
        RECT 709.950 139.950 712.050 140.400 ;
        RECT 718.950 139.950 721.050 140.400 ;
        RECT 724.950 139.950 727.050 142.050 ;
        RECT 730.950 139.950 733.050 142.050 ;
        RECT 748.950 139.950 751.050 142.050 ;
        RECT 754.950 141.450 757.050 142.050 ;
        RECT 759.000 141.450 763.050 142.050 ;
        RECT 754.950 140.400 763.050 141.450 ;
        RECT 754.950 139.950 757.050 140.400 ;
        RECT 759.000 139.950 763.050 140.400 ;
        RECT 769.950 139.950 772.050 142.050 ;
        RECT 775.950 139.950 778.050 142.050 ;
        RECT 793.950 139.950 796.050 142.050 ;
        RECT 799.950 139.950 802.050 142.050 ;
        RECT 817.950 139.950 820.050 142.050 ;
        RECT 823.950 141.450 826.050 142.050 ;
        RECT 835.950 141.450 838.050 142.050 ;
        RECT 823.950 140.400 838.050 141.450 ;
        RECT 823.950 139.950 826.050 140.400 ;
        RECT 835.950 139.950 838.050 140.400 ;
        RECT 841.950 139.950 844.050 142.050 ;
        RECT 847.950 139.950 850.050 142.050 ;
        RECT 853.950 141.450 856.050 142.050 ;
        RECT 865.950 141.450 868.050 142.050 ;
        RECT 853.950 140.400 868.050 141.450 ;
        RECT 853.950 139.950 856.050 140.400 ;
        RECT 865.950 139.950 868.050 140.400 ;
        RECT 883.950 139.950 886.050 142.050 ;
        RECT 889.950 139.950 892.050 142.050 ;
        RECT 724.950 136.950 727.050 138.750 ;
        RECT 730.950 136.950 733.050 138.750 ;
        RECT 748.950 136.950 751.050 138.750 ;
        RECT 754.950 136.950 757.050 138.750 ;
        RECT 769.950 136.950 772.050 138.750 ;
        RECT 775.950 136.950 778.050 138.750 ;
        RECT 793.950 136.950 796.050 138.750 ;
        RECT 799.950 136.950 802.050 138.750 ;
        RECT 817.950 136.950 820.050 138.750 ;
        RECT 823.950 136.950 826.050 138.750 ;
        RECT 841.950 136.950 844.050 138.750 ;
        RECT 847.950 136.950 850.050 138.750 ;
        RECT 865.950 136.950 868.050 138.750 ;
        RECT 883.950 136.950 886.050 138.750 ;
        RECT 889.950 136.950 892.050 138.750 ;
        RECT 685.950 133.950 688.050 135.750 ;
        RECT 703.950 133.950 706.050 135.750 ;
        RECT 709.950 134.250 712.050 136.050 ;
        RECT 721.950 134.250 724.050 136.050 ;
        RECT 727.950 134.250 730.050 136.050 ;
        RECT 751.950 134.250 754.050 136.050 ;
        RECT 772.950 134.250 775.050 136.050 ;
        RECT 778.950 134.250 781.050 136.050 ;
        RECT 796.950 134.250 799.050 136.050 ;
        RECT 802.950 134.250 805.050 136.050 ;
        RECT 814.950 134.250 817.050 136.050 ;
        RECT 820.950 134.250 823.050 136.050 ;
        RECT 844.950 134.250 847.050 136.050 ;
        RECT 850.950 134.250 853.050 136.050 ;
        RECT 862.950 134.250 865.050 136.050 ;
        RECT 880.950 134.250 883.050 136.050 ;
        RECT 886.950 134.250 889.050 136.050 ;
        RECT 904.950 135.450 907.050 136.050 ;
        RECT 910.950 135.450 913.050 136.050 ;
        RECT 904.950 134.400 913.050 135.450 ;
        RECT 904.950 133.950 907.050 134.400 ;
        RECT 910.950 133.950 913.050 134.400 ;
        RECT 709.950 130.950 715.050 133.050 ;
        RECT 721.950 130.950 724.050 133.050 ;
        RECT 727.950 127.950 730.050 133.050 ;
        RECT 751.950 132.450 754.050 133.050 ;
        RECT 766.950 132.450 769.050 133.050 ;
        RECT 751.950 131.400 769.050 132.450 ;
        RECT 751.950 130.950 754.050 131.400 ;
        RECT 766.950 130.950 769.050 131.400 ;
        RECT 772.950 130.950 775.050 133.050 ;
        RECT 778.950 130.950 781.050 133.050 ;
        RECT 784.950 132.450 787.050 133.050 ;
        RECT 796.950 132.450 799.050 133.050 ;
        RECT 784.950 131.400 799.050 132.450 ;
        RECT 784.950 130.950 787.050 131.400 ;
        RECT 796.950 130.950 799.050 131.400 ;
        RECT 802.950 132.450 805.050 133.050 ;
        RECT 807.000 132.450 811.050 133.050 ;
        RECT 802.950 131.400 811.050 132.450 ;
        RECT 802.950 130.950 805.050 131.400 ;
        RECT 807.000 130.950 811.050 131.400 ;
        RECT 814.950 130.950 817.050 133.050 ;
        RECT 820.950 130.950 823.050 133.050 ;
        RECT 829.950 132.450 832.050 133.050 ;
        RECT 844.950 132.450 847.050 133.050 ;
        RECT 829.950 131.400 847.050 132.450 ;
        RECT 829.950 130.950 832.050 131.400 ;
        RECT 844.950 130.950 847.050 131.400 ;
        RECT 850.950 130.950 853.050 133.050 ;
        RECT 862.950 130.950 865.050 133.050 ;
        RECT 880.950 130.950 883.050 133.050 ;
        RECT 886.950 132.450 892.050 133.050 ;
        RECT 907.950 132.450 910.050 133.050 ;
        RECT 886.950 131.400 910.050 132.450 ;
        RECT 886.950 130.950 892.050 131.400 ;
        RECT 907.950 130.950 910.050 131.400 ;
        RECT 626.400 125.400 643.050 126.450 ;
        RECT 508.950 124.950 511.050 125.400 ;
        RECT 553.950 124.950 556.050 125.400 ;
        RECT 619.950 124.950 622.050 125.400 ;
        RECT 640.950 124.950 643.050 125.400 ;
        RECT 661.950 124.500 664.050 126.600 ;
        RECT 682.950 124.500 685.050 126.600 ;
        RECT 773.400 126.450 774.450 130.950 ;
        RECT 781.950 126.450 784.050 127.050 ;
        RECT 773.400 125.400 784.050 126.450 ;
        RECT 781.950 124.950 784.050 125.400 ;
        RECT 814.950 126.450 817.050 127.050 ;
        RECT 821.400 126.450 822.450 130.950 ;
        RECT 814.950 125.400 822.450 126.450 ;
        RECT 835.950 126.450 838.050 127.050 ;
        RECT 862.950 126.450 865.050 127.050 ;
        RECT 892.950 126.450 895.050 127.050 ;
        RECT 835.950 125.400 895.050 126.450 ;
        RECT 814.950 124.950 817.050 125.400 ;
        RECT 835.950 124.950 838.050 125.400 ;
        RECT 862.950 124.950 865.050 125.400 ;
        RECT 892.950 124.950 895.050 125.400 ;
        RECT 19.950 123.450 22.050 124.050 ;
        RECT 25.950 123.450 28.050 124.050 ;
        RECT 34.950 123.450 37.050 124.050 ;
        RECT 19.950 122.400 37.050 123.450 ;
        RECT 19.950 121.950 22.050 122.400 ;
        RECT 25.950 121.950 28.050 122.400 ;
        RECT 34.950 121.950 37.050 122.400 ;
        RECT 67.950 123.450 70.050 124.050 ;
        RECT 91.950 123.450 97.050 124.050 ;
        RECT 67.950 122.400 97.050 123.450 ;
        RECT 67.950 121.950 70.050 122.400 ;
        RECT 91.950 121.950 97.050 122.400 ;
        RECT 151.950 123.450 154.050 124.050 ;
        RECT 178.950 123.450 181.050 124.050 ;
        RECT 151.950 122.400 181.050 123.450 ;
        RECT 151.950 121.950 154.050 122.400 ;
        RECT 178.950 121.950 181.050 122.400 ;
        RECT 370.950 123.450 373.050 123.900 ;
        RECT 397.950 123.450 400.050 124.050 ;
        RECT 370.950 122.400 400.050 123.450 ;
        RECT 370.950 121.800 373.050 122.400 ;
        RECT 397.950 121.950 400.050 122.400 ;
        RECT 403.950 123.450 406.050 124.050 ;
        RECT 424.950 123.450 427.050 124.050 ;
        RECT 403.950 122.400 427.050 123.450 ;
        RECT 403.950 121.950 406.050 122.400 ;
        RECT 424.950 121.950 427.050 122.400 ;
        RECT 430.950 123.450 433.050 124.050 ;
        RECT 451.950 123.450 454.050 124.050 ;
        RECT 430.950 122.400 454.050 123.450 ;
        RECT 430.950 121.950 433.050 122.400 ;
        RECT 451.950 121.950 454.050 122.400 ;
        RECT 13.950 120.450 16.050 121.050 ;
        RECT 46.950 120.450 49.050 121.050 ;
        RECT 13.950 119.400 49.050 120.450 ;
        RECT 13.950 118.950 16.050 119.400 ;
        RECT 46.950 118.950 49.050 119.400 ;
        RECT 133.950 120.450 136.050 121.050 ;
        RECT 139.950 120.450 142.050 121.050 ;
        RECT 133.950 119.400 142.050 120.450 ;
        RECT 133.950 118.950 136.050 119.400 ;
        RECT 139.950 118.950 142.050 119.400 ;
        RECT 160.950 120.450 163.050 121.050 ;
        RECT 169.950 120.450 172.050 121.050 ;
        RECT 160.950 119.400 172.050 120.450 ;
        RECT 160.950 118.950 163.050 119.400 ;
        RECT 169.950 118.950 172.050 119.400 ;
        RECT 211.950 120.450 214.050 121.050 ;
        RECT 292.950 120.450 295.050 121.050 ;
        RECT 301.950 120.450 304.050 121.050 ;
        RECT 211.950 119.400 246.450 120.450 ;
        RECT 211.950 118.950 214.050 119.400 ;
        RECT 245.400 118.050 246.450 119.400 ;
        RECT 292.950 119.400 304.050 120.450 ;
        RECT 292.950 118.950 295.050 119.400 ;
        RECT 301.950 118.950 304.050 119.400 ;
        RECT 391.950 120.450 394.050 121.050 ;
        RECT 445.950 120.450 448.050 121.050 ;
        RECT 487.950 120.450 490.050 124.050 ;
        RECT 496.950 123.450 499.050 124.050 ;
        RECT 502.950 123.450 505.050 124.050 ;
        RECT 496.950 122.400 505.050 123.450 ;
        RECT 496.950 121.950 499.050 122.400 ;
        RECT 502.950 121.950 505.050 122.400 ;
        RECT 523.950 123.450 526.050 124.050 ;
        RECT 799.950 123.450 802.050 124.050 ;
        RECT 820.950 123.450 823.050 124.050 ;
        RECT 523.950 122.400 657.450 123.450 ;
        RECT 523.950 121.950 526.050 122.400 ;
        RECT 586.950 120.450 589.050 121.050 ;
        RECT 391.950 119.400 589.050 120.450 ;
        RECT 656.400 120.450 657.450 122.400 ;
        RECT 799.950 122.400 823.050 123.450 ;
        RECT 799.950 121.950 802.050 122.400 ;
        RECT 820.950 121.950 823.050 122.400 ;
        RECT 688.950 120.450 691.050 121.050 ;
        RECT 656.400 119.400 691.050 120.450 ;
        RECT 391.950 118.950 394.050 119.400 ;
        RECT 445.950 118.950 448.050 119.400 ;
        RECT 586.950 118.950 589.050 119.400 ;
        RECT 688.950 118.950 691.050 119.400 ;
        RECT 694.950 120.450 697.050 121.050 ;
        RECT 847.950 120.450 850.050 121.050 ;
        RECT 883.950 120.450 886.050 121.050 ;
        RECT 694.950 119.400 886.050 120.450 ;
        RECT 694.950 118.950 697.050 119.400 ;
        RECT 847.950 118.950 850.050 119.400 ;
        RECT 883.950 118.950 886.050 119.400 ;
        RECT 43.950 117.450 46.050 118.050 ;
        RECT 73.950 117.450 76.050 118.050 ;
        RECT 43.950 116.400 76.050 117.450 ;
        RECT 43.950 115.950 46.050 116.400 ;
        RECT 73.950 115.950 76.050 116.400 ;
        RECT 82.950 117.450 85.050 118.050 ;
        RECT 103.950 117.450 106.050 118.050 ;
        RECT 115.950 117.450 118.050 118.050 ;
        RECT 82.950 117.000 99.450 117.450 ;
        RECT 82.950 116.400 100.050 117.000 ;
        RECT 82.950 115.950 85.050 116.400 ;
        RECT 97.950 115.050 100.050 116.400 ;
        RECT 103.950 116.400 118.050 117.450 ;
        RECT 103.950 115.950 106.050 116.400 ;
        RECT 115.950 115.950 118.050 116.400 ;
        RECT 145.950 117.450 148.050 118.050 ;
        RECT 172.950 117.450 175.050 118.050 ;
        RECT 145.950 116.400 175.050 117.450 ;
        RECT 145.950 115.950 148.050 116.400 ;
        RECT 172.950 115.950 175.050 116.400 ;
        RECT 178.950 117.450 181.050 118.050 ;
        RECT 193.950 117.450 196.050 118.050 ;
        RECT 178.950 116.400 196.050 117.450 ;
        RECT 178.950 115.950 181.050 116.400 ;
        RECT 193.950 115.950 196.050 116.400 ;
        RECT 220.950 117.450 223.050 118.050 ;
        RECT 229.950 117.450 232.050 118.050 ;
        RECT 220.950 116.400 232.050 117.450 ;
        RECT 220.950 115.950 223.050 116.400 ;
        RECT 229.950 115.950 232.050 116.400 ;
        RECT 244.950 117.450 247.050 118.050 ;
        RECT 274.950 117.450 277.050 118.050 ;
        RECT 244.950 116.400 277.050 117.450 ;
        RECT 244.950 115.950 247.050 116.400 ;
        RECT 274.950 115.950 277.050 116.400 ;
        RECT 286.950 117.450 289.050 118.050 ;
        RECT 487.950 117.450 490.050 118.050 ;
        RECT 517.950 117.450 520.050 118.050 ;
        RECT 286.950 116.400 490.050 117.450 ;
        RECT 286.950 115.950 289.050 116.400 ;
        RECT 487.950 115.950 490.050 116.400 ;
        RECT 506.400 116.400 520.050 117.450 ;
        RECT 28.950 114.450 31.050 115.050 ;
        RECT 37.950 114.450 40.050 115.050 ;
        RECT 28.950 113.400 40.050 114.450 ;
        RECT 28.950 112.950 31.050 113.400 ;
        RECT 37.950 112.950 40.050 113.400 ;
        RECT 61.950 114.450 64.050 115.050 ;
        RECT 94.800 114.450 96.900 115.050 ;
        RECT 61.950 113.400 96.900 114.450 ;
        RECT 97.950 114.000 100.200 115.050 ;
        RECT 61.950 112.950 64.050 113.400 ;
        RECT 94.800 112.950 96.900 113.400 ;
        RECT 98.100 112.950 100.200 114.000 ;
        RECT 208.950 114.450 211.050 115.050 ;
        RECT 217.950 114.450 220.050 115.050 ;
        RECT 208.950 113.400 220.050 114.450 ;
        RECT 208.950 112.950 211.050 113.400 ;
        RECT 217.950 112.950 220.050 113.400 ;
        RECT 238.950 114.450 241.050 115.050 ;
        RECT 256.950 114.450 259.050 115.050 ;
        RECT 295.950 114.450 298.050 115.050 ;
        RECT 238.950 113.400 298.050 114.450 ;
        RECT 238.950 112.950 241.050 113.400 ;
        RECT 256.950 112.950 259.050 113.400 ;
        RECT 295.950 112.950 298.050 113.400 ;
        RECT 301.950 114.450 304.050 115.050 ;
        RECT 337.950 114.450 340.050 115.050 ;
        RECT 301.950 113.400 340.050 114.450 ;
        RECT 301.950 112.950 304.050 113.400 ;
        RECT 337.950 112.950 340.050 113.400 ;
        RECT 397.950 114.450 400.050 115.050 ;
        RECT 409.950 114.450 412.050 115.050 ;
        RECT 418.950 114.450 421.050 115.050 ;
        RECT 397.950 113.400 421.050 114.450 ;
        RECT 397.950 112.950 400.050 113.400 ;
        RECT 409.950 112.950 412.050 113.400 ;
        RECT 418.950 112.950 421.050 113.400 ;
        RECT 463.950 112.950 469.050 115.050 ;
        RECT 478.950 114.450 481.050 115.050 ;
        RECT 506.400 114.450 507.450 116.400 ;
        RECT 517.950 115.950 520.050 116.400 ;
        RECT 565.950 117.450 568.050 118.050 ;
        RECT 655.950 117.450 658.050 118.050 ;
        RECT 565.950 117.000 606.300 117.450 ;
        RECT 565.950 116.400 607.050 117.000 ;
        RECT 565.950 115.950 568.050 116.400 ;
        RECT 604.950 115.050 607.050 116.400 ;
        RECT 650.400 116.400 658.050 117.450 ;
        RECT 650.400 115.050 651.450 116.400 ;
        RECT 655.950 115.950 658.050 116.400 ;
        RECT 721.950 117.450 724.050 118.050 ;
        RECT 838.950 117.450 841.050 118.050 ;
        RECT 853.950 117.450 856.050 118.050 ;
        RECT 721.950 116.400 856.050 117.450 ;
        RECT 721.950 115.950 724.050 116.400 ;
        RECT 838.950 115.950 841.050 116.400 ;
        RECT 853.950 115.950 856.050 116.400 ;
        RECT 478.950 113.400 507.450 114.450 ;
        RECT 553.950 114.450 556.050 115.050 ;
        RECT 562.950 114.450 565.050 115.050 ;
        RECT 553.950 113.400 565.050 114.450 ;
        RECT 478.950 112.950 481.050 113.400 ;
        RECT 553.950 112.950 556.050 113.400 ;
        RECT 562.950 112.950 565.050 113.400 ;
        RECT 604.800 114.000 607.050 115.050 ;
        RECT 608.100 114.450 610.200 115.050 ;
        RECT 616.950 114.450 619.050 115.050 ;
        RECT 604.800 112.950 606.900 114.000 ;
        RECT 608.100 113.400 619.050 114.450 ;
        RECT 608.100 112.950 610.200 113.400 ;
        RECT 616.950 112.950 619.050 113.400 ;
        RECT 646.950 113.400 651.450 115.050 ;
        RECT 652.950 114.450 655.050 115.050 ;
        RECT 670.950 114.450 673.050 115.050 ;
        RECT 652.950 113.400 673.050 114.450 ;
        RECT 646.950 112.950 651.000 113.400 ;
        RECT 652.950 112.950 655.050 113.400 ;
        RECT 670.950 112.950 673.050 113.400 ;
        RECT 688.950 114.450 691.050 115.050 ;
        RECT 703.950 114.450 706.050 115.050 ;
        RECT 688.950 113.400 706.050 114.450 ;
        RECT 688.950 112.950 691.050 113.400 ;
        RECT 703.950 112.950 706.050 113.400 ;
        RECT 862.950 114.450 865.050 115.050 ;
        RECT 868.950 114.450 871.050 115.050 ;
        RECT 862.950 113.400 871.050 114.450 ;
        RECT 862.950 112.950 865.050 113.400 ;
        RECT 868.950 112.950 871.050 113.400 ;
        RECT 97.950 111.450 100.050 112.050 ;
        RECT 86.400 110.400 100.050 111.450 ;
        RECT 163.950 110.400 166.050 112.500 ;
        RECT 184.950 110.400 187.050 112.500 ;
        RECT 226.950 111.450 229.050 112.050 ;
        RECT 244.950 111.450 247.050 112.050 ;
        RECT 286.950 111.450 289.050 112.050 ;
        RECT 226.950 110.400 247.050 111.450 ;
        RECT 61.950 106.950 64.050 109.050 ;
        RECT 67.950 106.950 70.050 109.050 ;
        RECT 86.400 106.050 87.450 110.400 ;
        RECT 97.950 109.950 100.050 110.400 ;
        RECT 145.950 106.950 148.050 109.050 ;
        RECT 151.950 106.950 154.050 109.050 ;
        RECT 16.950 103.950 19.050 106.050 ;
        RECT 37.950 103.950 40.050 106.050 ;
        RECT 43.950 105.450 46.050 106.050 ;
        RECT 55.950 105.450 58.050 106.050 ;
        RECT 43.950 104.400 58.050 105.450 ;
        RECT 43.950 103.950 46.050 104.400 ;
        RECT 55.950 103.950 58.050 104.400 ;
        RECT 61.950 103.950 64.050 105.750 ;
        RECT 67.950 103.950 70.050 105.750 ;
        RECT 85.950 103.950 88.050 106.050 ;
        RECT 91.950 103.950 94.050 106.050 ;
        RECT 109.950 103.950 112.050 106.050 ;
        RECT 118.950 105.450 121.050 106.050 ;
        RECT 127.950 105.450 130.050 106.050 ;
        RECT 118.950 104.400 130.050 105.450 ;
        RECT 118.950 103.950 121.050 104.400 ;
        RECT 127.950 103.950 130.050 104.400 ;
        RECT 133.950 103.950 136.050 106.050 ;
        RECT 145.950 103.950 148.050 105.750 ;
        RECT 151.950 103.950 154.050 105.750 ;
        RECT 160.950 103.950 163.050 106.050 ;
        RECT 10.950 101.250 13.050 103.050 ;
        RECT 20.250 102.750 22.050 103.050 ;
        RECT 16.950 101.250 19.050 102.750 ;
        RECT 19.950 101.250 22.050 102.750 ;
        RECT 16.950 100.950 18.750 101.250 ;
        RECT 37.950 100.950 40.050 102.750 ;
        RECT 43.950 100.950 46.050 102.750 ;
        RECT 64.950 101.250 67.050 103.050 ;
        RECT 85.950 100.950 88.050 102.750 ;
        RECT 91.950 100.950 94.050 102.750 ;
        RECT 109.950 100.950 112.050 102.750 ;
        RECT 127.950 100.950 130.050 102.750 ;
        RECT 133.950 100.950 136.050 102.750 ;
        RECT 148.950 101.250 151.050 103.050 ;
        RECT 160.950 100.950 163.050 102.750 ;
        RECT 10.950 97.950 13.050 100.050 ;
        RECT 19.950 99.450 22.050 100.050 ;
        RECT 28.950 99.450 31.050 100.050 ;
        RECT 19.950 98.400 31.050 99.450 ;
        RECT 19.950 97.950 22.050 98.400 ;
        RECT 28.950 97.950 31.050 98.400 ;
        RECT 34.950 98.250 37.050 100.050 ;
        RECT 40.950 98.250 43.050 100.050 ;
        RECT 64.950 99.450 67.050 100.050 ;
        RECT 73.950 99.450 76.050 100.050 ;
        RECT 64.950 98.400 76.050 99.450 ;
        RECT 64.950 97.950 67.050 98.400 ;
        RECT 73.950 97.950 76.050 98.400 ;
        RECT 82.950 98.250 85.050 100.050 ;
        RECT 88.950 98.250 91.050 100.050 ;
        RECT 106.950 98.250 109.050 100.050 ;
        RECT 124.950 98.250 127.050 100.050 ;
        RECT 130.950 98.250 133.050 100.050 ;
        RECT 139.950 99.450 142.050 100.050 ;
        RECT 148.950 99.450 151.050 100.050 ;
        RECT 139.950 98.400 151.050 99.450 ;
        RECT 139.950 97.950 142.050 98.400 ;
        RECT 148.950 97.950 151.050 98.400 ;
        RECT 34.950 94.950 37.050 97.050 ;
        RECT 40.950 94.950 43.050 97.050 ;
        RECT 82.950 94.950 85.050 97.050 ;
        RECT 88.950 94.950 91.050 97.050 ;
        RECT 106.950 96.450 109.050 97.050 ;
        RECT 118.950 96.450 121.050 97.050 ;
        RECT 106.950 95.400 121.050 96.450 ;
        RECT 106.950 94.950 109.050 95.400 ;
        RECT 118.950 94.950 121.050 95.400 ;
        RECT 124.950 94.950 127.050 97.050 ;
        RECT 130.950 94.950 133.050 97.050 ;
        RECT 164.850 95.400 166.050 110.400 ;
        RECT 178.950 101.250 181.050 103.050 ;
        RECT 178.950 97.950 181.050 100.050 ;
        RECT 10.950 93.450 13.050 94.050 ;
        RECT 25.950 93.450 28.050 94.050 ;
        RECT 10.950 92.400 28.050 93.450 ;
        RECT 10.950 91.950 13.050 92.400 ;
        RECT 25.950 91.950 28.050 92.400 ;
        RECT 88.950 90.450 91.050 91.050 ;
        RECT 107.400 90.450 108.450 94.950 ;
        RECT 163.950 93.300 166.050 95.400 ;
        RECT 88.950 89.400 108.450 90.450 ;
        RECT 118.950 90.450 121.050 91.050 ;
        RECT 142.950 90.450 145.050 91.050 ;
        RECT 118.950 89.400 145.050 90.450 ;
        RECT 164.850 89.700 166.050 93.300 ;
        RECT 185.100 90.600 186.300 110.400 ;
        RECT 226.950 109.950 229.050 110.400 ;
        RECT 244.950 109.950 247.050 110.400 ;
        RECT 251.400 110.400 289.050 111.450 ;
        RECT 187.950 108.450 190.050 109.050 ;
        RECT 202.950 108.450 205.050 109.050 ;
        RECT 187.950 107.400 205.050 108.450 ;
        RECT 187.950 106.950 190.050 107.400 ;
        RECT 202.950 106.950 205.050 107.400 ;
        RECT 208.950 106.950 211.050 109.050 ;
        RECT 202.950 103.950 205.050 105.750 ;
        RECT 208.950 103.950 211.050 105.750 ;
        RECT 229.950 103.950 232.050 109.050 ;
        RECT 251.400 106.050 252.450 110.400 ;
        RECT 286.950 109.950 289.050 110.400 ;
        RECT 307.950 111.450 310.050 112.050 ;
        RECT 334.950 111.450 337.050 112.050 ;
        RECT 307.950 110.400 337.050 111.450 ;
        RECT 307.950 109.950 310.050 110.400 ;
        RECT 334.950 109.950 337.050 110.400 ;
        RECT 349.950 111.450 352.050 112.050 ;
        RECT 355.950 111.450 358.050 112.050 ;
        RECT 349.950 110.400 358.050 111.450 ;
        RECT 349.950 109.950 352.050 110.400 ;
        RECT 355.950 109.950 358.050 110.400 ;
        RECT 394.950 111.450 397.050 112.050 ;
        RECT 400.950 111.450 403.050 112.050 ;
        RECT 394.950 110.400 403.050 111.450 ;
        RECT 394.950 109.950 397.050 110.400 ;
        RECT 400.950 109.950 403.050 110.400 ;
        RECT 439.950 111.450 442.050 112.050 ;
        RECT 451.950 111.450 454.050 112.050 ;
        RECT 484.950 111.450 487.050 112.050 ;
        RECT 499.950 111.450 502.050 112.050 ;
        RECT 439.950 110.400 502.050 111.450 ;
        RECT 511.950 110.400 514.050 112.500 ;
        RECT 532.950 110.400 535.050 112.500 ;
        RECT 544.950 111.450 547.050 112.050 ;
        RECT 550.950 111.450 553.050 112.050 ;
        RECT 544.950 110.400 553.050 111.450 ;
        RECT 571.950 110.400 574.050 112.500 ;
        RECT 592.950 110.400 595.050 112.500 ;
        RECT 625.950 111.450 628.050 112.050 ;
        RECT 643.950 111.450 646.050 112.050 ;
        RECT 625.950 110.400 646.050 111.450 ;
        RECT 439.950 109.950 442.050 110.400 ;
        RECT 451.950 109.950 454.050 110.400 ;
        RECT 484.950 109.950 487.050 110.400 ;
        RECT 499.950 109.950 502.050 110.400 ;
        RECT 295.950 106.950 298.050 109.050 ;
        RECT 301.950 106.950 304.050 109.050 ;
        RECT 409.950 106.950 412.050 109.050 ;
        RECT 415.950 106.950 418.050 109.050 ;
        RECT 490.950 106.950 496.050 109.050 ;
        RECT 244.950 103.950 247.050 106.050 ;
        RECT 250.950 103.950 253.050 106.050 ;
        RECT 256.950 105.450 259.050 106.050 ;
        RECT 271.950 105.450 274.050 106.050 ;
        RECT 256.950 104.400 274.050 105.450 ;
        RECT 256.950 103.950 259.050 104.400 ;
        RECT 271.950 103.950 274.050 104.400 ;
        RECT 295.950 103.950 298.050 105.750 ;
        RECT 301.950 103.950 304.050 105.750 ;
        RECT 325.950 103.950 328.050 106.050 ;
        RECT 349.950 103.950 352.050 106.050 ;
        RECT 370.950 103.950 373.050 106.050 ;
        RECT 385.950 103.950 391.050 106.050 ;
        RECT 394.950 105.450 397.050 106.050 ;
        RECT 403.950 105.450 406.050 106.050 ;
        RECT 394.950 104.400 406.050 105.450 ;
        RECT 394.950 103.950 397.050 104.400 ;
        RECT 403.950 103.950 406.050 104.400 ;
        RECT 409.950 103.950 412.050 105.750 ;
        RECT 415.950 103.950 418.050 105.750 ;
        RECT 427.950 103.950 430.050 106.050 ;
        RECT 451.950 103.950 454.050 106.050 ;
        RECT 469.950 103.950 472.050 106.050 ;
        RECT 475.950 103.950 480.900 106.050 ;
        RECT 482.100 105.450 484.200 106.050 ;
        RECT 499.950 105.450 502.050 106.050 ;
        RECT 482.100 104.400 502.050 105.450 ;
        RECT 482.100 103.950 484.200 104.400 ;
        RECT 499.950 103.950 502.050 104.400 ;
        RECT 187.950 101.250 190.050 103.050 ;
        RECT 205.950 101.250 208.050 103.050 ;
        RECT 229.950 100.950 232.050 102.750 ;
        RECT 244.950 100.950 247.050 102.750 ;
        RECT 250.950 100.950 253.050 102.750 ;
        RECT 271.950 100.950 274.050 102.750 ;
        RECT 292.950 101.250 295.050 103.050 ;
        RECT 298.950 101.250 301.050 103.050 ;
        RECT 304.950 101.250 307.050 103.050 ;
        RECT 319.950 101.250 322.050 103.050 ;
        RECT 325.950 100.950 328.050 102.750 ;
        RECT 343.950 101.250 346.050 103.050 ;
        RECT 349.950 100.950 352.050 102.750 ;
        RECT 370.950 100.950 373.050 102.750 ;
        RECT 388.950 100.950 391.050 102.750 ;
        RECT 394.950 100.950 397.050 102.750 ;
        RECT 412.950 101.250 415.050 103.050 ;
        RECT 427.950 100.950 430.050 102.750 ;
        RECT 445.950 101.250 448.050 103.050 ;
        RECT 455.250 102.750 457.050 103.050 ;
        RECT 451.950 101.250 454.050 102.750 ;
        RECT 454.950 101.250 457.050 102.750 ;
        RECT 451.950 100.950 453.750 101.250 ;
        RECT 469.950 100.950 472.050 102.750 ;
        RECT 475.950 100.950 478.050 102.750 ;
        RECT 499.950 100.950 502.050 102.750 ;
        RECT 508.950 101.250 511.050 103.050 ;
        RECT 187.950 97.950 190.050 100.050 ;
        RECT 193.950 99.450 196.050 100.050 ;
        RECT 205.950 99.450 208.050 100.050 ;
        RECT 193.950 98.400 208.050 99.450 ;
        RECT 193.950 97.950 196.050 98.400 ;
        RECT 205.950 97.950 208.050 98.400 ;
        RECT 226.950 98.250 229.050 100.050 ;
        RECT 232.950 98.250 235.050 100.050 ;
        RECT 247.950 98.250 250.050 100.050 ;
        RECT 253.950 98.250 256.050 100.050 ;
        RECT 268.950 98.250 271.050 100.050 ;
        RECT 274.950 98.250 277.050 100.050 ;
        RECT 292.950 97.950 295.050 100.050 ;
        RECT 226.950 94.950 229.050 97.050 ;
        RECT 232.950 96.450 235.050 97.050 ;
        RECT 237.000 96.450 241.050 97.050 ;
        RECT 232.950 95.400 241.050 96.450 ;
        RECT 232.950 94.950 235.050 95.400 ;
        RECT 237.000 94.950 241.050 95.400 ;
        RECT 247.950 94.950 250.050 97.050 ;
        RECT 253.950 94.950 256.050 97.050 ;
        RECT 268.950 91.950 271.050 97.050 ;
        RECT 274.950 94.950 277.050 97.050 ;
        RECT 298.950 94.950 301.050 100.050 ;
        RECT 304.950 97.950 307.050 100.050 ;
        RECT 310.950 99.450 313.050 100.050 ;
        RECT 319.950 99.450 325.050 100.050 ;
        RECT 310.950 98.400 325.050 99.450 ;
        RECT 310.950 97.950 313.050 98.400 ;
        RECT 319.950 97.950 325.050 98.400 ;
        RECT 328.950 99.450 331.050 100.050 ;
        RECT 343.950 99.450 346.050 100.050 ;
        RECT 328.950 98.400 346.050 99.450 ;
        RECT 328.950 97.950 331.050 98.400 ;
        RECT 343.950 97.950 346.050 98.400 ;
        RECT 367.950 98.250 370.050 100.050 ;
        RECT 385.950 98.250 388.050 100.050 ;
        RECT 391.950 98.250 394.050 100.050 ;
        RECT 412.950 99.450 415.050 100.050 ;
        RECT 424.950 99.450 427.050 100.050 ;
        RECT 412.950 98.400 427.050 99.450 ;
        RECT 412.950 97.950 415.050 98.400 ;
        RECT 424.950 97.950 427.050 98.400 ;
        RECT 430.950 98.250 433.050 100.050 ;
        RECT 445.950 97.950 448.050 100.050 ;
        RECT 454.950 99.450 457.050 100.050 ;
        RECT 466.950 99.450 469.050 100.050 ;
        RECT 454.950 98.400 469.050 99.450 ;
        RECT 454.950 97.950 457.050 98.400 ;
        RECT 466.950 97.950 469.050 98.400 ;
        RECT 472.950 98.250 475.050 100.050 ;
        RECT 478.950 98.250 481.050 100.050 ;
        RECT 496.950 98.250 499.050 100.050 ;
        RECT 502.950 98.250 505.050 100.050 ;
        RECT 508.950 97.950 511.050 100.050 ;
        RECT 367.950 96.450 370.050 97.050 ;
        RECT 385.950 96.450 388.050 97.050 ;
        RECT 367.950 95.400 388.050 96.450 ;
        RECT 367.950 94.950 370.050 95.400 ;
        RECT 385.950 94.950 388.050 95.400 ;
        RECT 391.950 94.950 394.050 97.050 ;
        RECT 430.950 96.450 433.050 97.050 ;
        RECT 439.950 96.450 442.050 97.050 ;
        RECT 430.950 95.400 442.050 96.450 ;
        RECT 430.950 94.950 433.050 95.400 ;
        RECT 439.950 94.950 442.050 95.400 ;
        RECT 472.950 94.950 475.050 97.050 ;
        RECT 478.950 94.950 481.050 97.050 ;
        RECT 496.950 94.950 499.050 97.050 ;
        RECT 292.950 93.450 295.050 94.050 ;
        RECT 334.950 93.450 337.050 94.050 ;
        RECT 292.950 92.400 337.050 93.450 ;
        RECT 292.950 91.950 295.050 92.400 ;
        RECT 334.950 91.950 337.050 92.400 ;
        RECT 502.950 91.950 505.050 97.050 ;
        RECT 88.950 88.950 91.050 89.400 ;
        RECT 118.950 88.950 121.050 89.400 ;
        RECT 142.950 88.950 145.050 89.400 ;
        RECT 55.950 87.450 58.050 88.050 ;
        RECT 100.950 87.450 103.050 88.050 ;
        RECT 130.950 87.450 133.050 88.050 ;
        RECT 163.950 87.600 166.050 89.700 ;
        RECT 184.950 88.500 187.050 90.600 ;
        RECT 202.950 90.450 205.050 91.050 ;
        RECT 247.950 90.450 250.050 91.050 ;
        RECT 202.950 89.400 250.050 90.450 ;
        RECT 202.950 88.950 205.050 89.400 ;
        RECT 247.950 88.950 250.050 89.400 ;
        RECT 274.950 90.450 277.050 91.050 ;
        RECT 310.950 90.450 313.050 91.050 ;
        RECT 274.950 89.400 313.050 90.450 ;
        RECT 274.950 88.950 277.050 89.400 ;
        RECT 310.950 88.950 313.050 89.400 ;
        RECT 379.950 88.950 384.900 91.050 ;
        RECT 386.100 90.450 388.200 91.050 ;
        RECT 391.950 90.450 394.050 91.050 ;
        RECT 386.100 89.400 394.050 90.450 ;
        RECT 386.100 88.950 388.200 89.400 ;
        RECT 391.950 88.950 394.050 89.400 ;
        RECT 427.950 90.450 430.050 91.050 ;
        RECT 487.950 90.450 490.050 91.050 ;
        RECT 512.700 90.600 513.900 110.400 ;
        RECT 517.950 101.250 520.050 103.050 ;
        RECT 517.950 97.950 520.050 100.050 ;
        RECT 532.950 95.400 534.150 110.400 ;
        RECT 544.950 109.950 547.050 110.400 ;
        RECT 550.950 109.950 553.050 110.400 ;
        RECT 535.950 105.450 538.050 106.050 ;
        RECT 544.950 105.450 547.050 106.050 ;
        RECT 535.950 104.400 547.050 105.450 ;
        RECT 535.950 103.950 538.050 104.400 ;
        RECT 544.950 103.950 547.050 104.400 ;
        RECT 550.950 103.950 553.050 106.050 ;
        RECT 556.950 105.450 559.050 106.050 ;
        RECT 565.950 105.450 568.050 106.050 ;
        RECT 556.950 104.400 568.050 105.450 ;
        RECT 556.950 103.950 559.050 104.400 ;
        RECT 565.950 103.950 568.050 104.400 ;
        RECT 535.950 100.950 538.050 102.750 ;
        RECT 550.950 100.950 553.050 102.750 ;
        RECT 556.950 100.950 559.050 102.750 ;
        RECT 568.950 101.250 571.050 103.050 ;
        RECT 553.950 98.250 556.050 100.050 ;
        RECT 559.950 98.250 562.050 100.050 ;
        RECT 568.950 97.950 571.050 100.050 ;
        RECT 517.950 93.450 520.050 94.050 ;
        RECT 526.950 93.450 529.050 94.050 ;
        RECT 517.950 92.400 529.050 93.450 ;
        RECT 517.950 91.950 520.050 92.400 ;
        RECT 526.950 91.950 529.050 92.400 ;
        RECT 532.950 93.300 535.050 95.400 ;
        RECT 553.950 94.950 556.050 97.050 ;
        RECT 559.950 94.950 562.050 97.050 ;
        RECT 544.950 93.450 547.050 94.050 ;
        RECT 550.950 93.450 553.050 94.050 ;
        RECT 427.950 89.400 490.050 90.450 ;
        RECT 427.950 88.950 430.050 89.400 ;
        RECT 487.950 88.950 490.050 89.400 ;
        RECT 511.950 88.500 514.050 90.600 ;
        RECT 532.950 89.700 534.150 93.300 ;
        RECT 544.950 92.400 553.050 93.450 ;
        RECT 544.950 91.950 547.050 92.400 ;
        RECT 550.950 91.950 553.050 92.400 ;
        RECT 572.700 90.600 573.900 110.400 ;
        RECT 580.950 105.450 583.050 106.050 ;
        RECT 586.950 105.450 589.050 106.050 ;
        RECT 580.950 104.400 589.050 105.450 ;
        RECT 580.950 103.950 583.050 104.400 ;
        RECT 586.950 103.950 589.050 104.400 ;
        RECT 577.950 101.250 580.050 103.050 ;
        RECT 577.950 97.950 580.050 100.050 ;
        RECT 592.950 95.400 594.150 110.400 ;
        RECT 625.950 109.950 628.050 110.400 ;
        RECT 643.950 109.950 646.050 110.400 ;
        RECT 649.950 111.450 652.050 112.050 ;
        RECT 655.950 111.450 658.050 112.050 ;
        RECT 649.950 110.400 658.050 111.450 ;
        RECT 649.950 109.950 652.050 110.400 ;
        RECT 655.950 109.950 658.050 110.400 ;
        RECT 721.950 111.450 724.050 112.050 ;
        RECT 727.950 111.450 730.050 112.050 ;
        RECT 721.950 110.400 730.050 111.450 ;
        RECT 721.950 109.950 724.050 110.400 ;
        RECT 727.950 109.950 730.050 110.400 ;
        RECT 736.950 111.450 739.050 112.050 ;
        RECT 748.950 111.450 751.050 112.050 ;
        RECT 736.950 110.400 751.050 111.450 ;
        RECT 766.950 110.400 769.050 112.500 ;
        RECT 787.950 110.400 790.050 112.500 ;
        RECT 736.950 109.950 739.050 110.400 ;
        RECT 748.950 109.950 751.050 110.400 ;
        RECT 610.950 106.950 613.050 109.050 ;
        RECT 616.950 106.950 619.050 109.050 ;
        RECT 682.950 106.950 685.050 109.050 ;
        RECT 688.950 106.950 691.050 109.050 ;
        RECT 595.950 103.950 598.050 106.050 ;
        RECT 610.950 103.950 613.050 105.750 ;
        RECT 616.950 103.950 619.050 105.750 ;
        RECT 634.950 103.950 637.050 106.050 ;
        RECT 640.950 105.450 643.050 106.050 ;
        RECT 649.950 105.450 652.050 106.050 ;
        RECT 640.950 104.400 652.050 105.450 ;
        RECT 640.950 103.950 643.050 104.400 ;
        RECT 649.950 103.950 652.050 104.400 ;
        RECT 655.950 103.950 658.050 106.050 ;
        RECT 661.950 105.450 664.050 106.050 ;
        RECT 670.950 105.450 673.050 106.050 ;
        RECT 661.950 104.400 673.050 105.450 ;
        RECT 661.950 103.950 664.050 104.400 ;
        RECT 670.950 103.950 673.050 104.400 ;
        RECT 682.950 103.950 685.050 105.750 ;
        RECT 688.950 103.950 691.050 105.750 ;
        RECT 703.950 103.950 706.050 106.050 ;
        RECT 715.950 105.450 718.050 106.050 ;
        RECT 730.950 105.450 733.050 106.050 ;
        RECT 715.950 104.400 733.050 105.450 ;
        RECT 715.950 103.950 718.050 104.400 ;
        RECT 730.950 103.950 733.050 104.400 ;
        RECT 736.950 103.950 739.050 106.050 ;
        RECT 748.950 103.950 751.050 106.050 ;
        RECT 763.950 103.950 766.050 106.050 ;
        RECT 595.950 100.950 598.050 102.750 ;
        RECT 613.950 101.250 616.050 103.050 ;
        RECT 634.950 100.950 637.050 102.750 ;
        RECT 640.950 100.950 643.050 102.750 ;
        RECT 655.950 100.950 658.050 102.750 ;
        RECT 661.950 100.950 664.050 102.750 ;
        RECT 685.950 101.250 688.050 103.050 ;
        RECT 703.950 100.950 706.050 102.750 ;
        RECT 709.950 101.250 712.050 103.050 ;
        RECT 730.950 100.950 733.050 102.750 ;
        RECT 736.950 100.950 739.050 102.750 ;
        RECT 748.950 100.950 751.050 102.750 ;
        RECT 754.950 101.250 757.050 103.050 ;
        RECT 763.950 100.950 766.050 102.750 ;
        RECT 613.950 99.450 616.050 100.050 ;
        RECT 625.950 99.450 628.050 100.050 ;
        RECT 613.950 98.400 628.050 99.450 ;
        RECT 613.950 97.950 616.050 98.400 ;
        RECT 625.950 97.950 628.050 98.400 ;
        RECT 631.950 98.250 634.050 100.050 ;
        RECT 637.950 98.250 640.050 100.050 ;
        RECT 643.950 99.450 646.050 100.050 ;
        RECT 652.950 99.450 655.050 100.050 ;
        RECT 643.950 98.400 655.050 99.450 ;
        RECT 643.950 97.950 646.050 98.400 ;
        RECT 652.950 97.950 655.050 98.400 ;
        RECT 658.950 98.250 661.050 100.050 ;
        RECT 664.950 98.250 667.050 100.050 ;
        RECT 685.950 99.450 688.050 100.050 ;
        RECT 694.950 99.450 697.050 100.050 ;
        RECT 685.950 98.400 697.050 99.450 ;
        RECT 685.950 97.950 688.050 98.400 ;
        RECT 694.950 97.950 697.050 98.400 ;
        RECT 700.950 98.250 703.050 100.050 ;
        RECT 709.950 99.450 712.050 100.050 ;
        RECT 721.950 99.450 724.050 100.050 ;
        RECT 709.950 98.400 724.050 99.450 ;
        RECT 709.950 97.950 712.050 98.400 ;
        RECT 721.950 97.950 724.050 98.400 ;
        RECT 727.950 98.250 730.050 100.050 ;
        RECT 733.950 98.250 736.050 100.050 ;
        RECT 751.950 97.950 757.050 100.050 ;
        RECT 622.950 96.450 625.050 97.050 ;
        RECT 631.950 96.450 634.050 97.050 ;
        RECT 622.950 95.400 634.050 96.450 ;
        RECT 592.950 93.300 595.050 95.400 ;
        RECT 622.950 94.950 625.050 95.400 ;
        RECT 631.950 94.950 634.050 95.400 ;
        RECT 637.950 96.450 640.050 97.050 ;
        RECT 652.950 96.450 655.050 97.050 ;
        RECT 637.950 95.400 655.050 96.450 ;
        RECT 637.950 94.950 640.050 95.400 ;
        RECT 652.950 94.950 655.050 95.400 ;
        RECT 658.950 94.950 661.050 97.050 ;
        RECT 664.950 94.950 667.050 97.050 ;
        RECT 700.950 94.950 703.050 97.050 ;
        RECT 727.950 94.950 730.050 97.050 ;
        RECT 733.950 94.950 736.050 97.050 ;
        RECT 767.850 95.400 769.050 110.400 ;
        RECT 781.950 101.250 784.050 103.050 ;
        RECT 781.950 97.950 784.050 100.050 ;
        RECT 766.950 93.300 769.050 95.400 ;
        RECT 55.950 86.400 133.050 87.450 ;
        RECT 55.950 85.950 58.050 86.400 ;
        RECT 100.950 85.950 103.050 86.400 ;
        RECT 130.950 85.950 133.050 86.400 ;
        RECT 433.950 87.450 436.050 88.050 ;
        RECT 439.800 87.450 441.900 88.050 ;
        RECT 433.950 86.400 441.900 87.450 ;
        RECT 433.950 85.950 436.050 86.400 ;
        RECT 439.800 85.950 441.900 86.400 ;
        RECT 443.100 87.450 445.200 88.050 ;
        RECT 460.800 87.450 462.900 88.050 ;
        RECT 443.100 86.400 462.900 87.450 ;
        RECT 443.100 85.950 445.200 86.400 ;
        RECT 460.800 85.950 462.900 86.400 ;
        RECT 464.100 87.450 466.200 88.050 ;
        RECT 472.950 87.450 475.050 88.050 ;
        RECT 532.950 87.600 535.050 89.700 ;
        RECT 571.950 88.500 574.050 90.600 ;
        RECT 592.950 89.700 594.150 93.300 ;
        RECT 646.950 90.450 649.050 91.050 ;
        RECT 658.950 90.450 661.050 91.050 ;
        RECT 592.950 87.600 595.050 89.700 ;
        RECT 646.950 89.400 661.050 90.450 ;
        RECT 646.950 88.950 649.050 89.400 ;
        RECT 658.950 88.950 661.050 89.400 ;
        RECT 721.950 90.450 724.050 91.050 ;
        RECT 727.950 90.450 730.050 91.050 ;
        RECT 721.950 89.400 730.050 90.450 ;
        RECT 721.950 88.950 724.050 89.400 ;
        RECT 727.950 88.950 730.050 89.400 ;
        RECT 733.950 90.450 736.050 91.050 ;
        RECT 742.950 90.450 745.050 91.050 ;
        RECT 751.950 90.450 754.050 91.050 ;
        RECT 733.950 89.400 754.050 90.450 ;
        RECT 767.850 89.700 769.050 93.300 ;
        RECT 788.100 90.600 789.300 110.400 ;
        RECT 853.950 106.950 856.050 109.050 ;
        RECT 859.950 106.950 862.050 109.050 ;
        RECT 895.950 106.950 898.050 109.050 ;
        RECT 901.950 106.950 904.050 109.050 ;
        RECT 796.950 105.450 799.050 106.050 ;
        RECT 808.950 105.450 811.050 106.050 ;
        RECT 796.950 104.400 811.050 105.450 ;
        RECT 796.950 103.950 799.050 104.400 ;
        RECT 808.950 103.950 811.050 104.400 ;
        RECT 820.950 105.450 823.050 106.050 ;
        RECT 829.950 105.450 832.050 106.050 ;
        RECT 820.950 104.400 832.050 105.450 ;
        RECT 820.950 103.950 823.050 104.400 ;
        RECT 829.950 103.950 832.050 104.400 ;
        RECT 835.950 103.950 838.050 106.050 ;
        RECT 853.950 103.950 856.050 105.750 ;
        RECT 859.950 103.950 862.050 105.750 ;
        RECT 865.950 105.450 868.050 106.050 ;
        RECT 877.950 105.450 880.050 106.050 ;
        RECT 865.950 104.400 880.050 105.450 ;
        RECT 865.950 103.950 868.050 104.400 ;
        RECT 877.950 103.950 880.050 104.400 ;
        RECT 883.950 103.950 886.050 106.050 ;
        RECT 895.950 103.950 898.050 105.750 ;
        RECT 901.950 103.950 904.050 105.750 ;
        RECT 790.950 101.250 793.050 103.050 ;
        RECT 808.950 100.950 811.050 102.750 ;
        RECT 829.950 100.950 832.050 102.750 ;
        RECT 835.950 100.950 838.050 102.750 ;
        RECT 856.950 101.250 859.050 103.050 ;
        RECT 877.950 100.950 880.050 102.750 ;
        RECT 883.950 100.950 886.050 102.750 ;
        RECT 898.950 101.250 901.050 103.050 ;
        RECT 790.950 97.950 793.050 100.050 ;
        RECT 805.950 98.250 808.050 100.050 ;
        RECT 811.950 98.250 814.050 100.050 ;
        RECT 832.950 98.250 835.050 100.050 ;
        RECT 838.950 98.250 841.050 100.050 ;
        RECT 805.950 94.950 808.050 97.050 ;
        RECT 811.950 94.950 814.050 97.050 ;
        RECT 832.950 94.950 835.050 97.050 ;
        RECT 838.950 94.950 841.050 97.050 ;
        RECT 856.950 94.950 859.050 100.050 ;
        RECT 874.950 98.250 877.050 100.050 ;
        RECT 880.950 98.250 883.050 100.050 ;
        RECT 892.950 99.450 897.000 100.050 ;
        RECT 898.950 99.450 901.050 100.050 ;
        RECT 892.950 98.400 901.050 99.450 ;
        RECT 892.950 97.950 897.000 98.400 ;
        RECT 898.950 97.950 901.050 98.400 ;
        RECT 874.950 94.950 877.050 97.050 ;
        RECT 880.950 94.950 883.050 97.050 ;
        RECT 886.950 94.950 892.050 97.050 ;
        RECT 886.950 93.450 889.050 94.050 ;
        RECT 895.950 93.450 898.050 94.050 ;
        RECT 886.950 92.400 898.050 93.450 ;
        RECT 886.950 91.950 889.050 92.400 ;
        RECT 895.950 91.950 898.050 92.400 ;
        RECT 733.950 88.950 736.050 89.400 ;
        RECT 742.950 88.950 745.050 89.400 ;
        RECT 751.950 88.950 754.050 89.400 ;
        RECT 464.100 86.400 475.050 87.450 ;
        RECT 464.100 85.950 466.200 86.400 ;
        RECT 472.950 85.950 475.050 86.400 ;
        RECT 604.950 87.450 607.050 88.050 ;
        RECT 616.950 87.450 619.050 88.050 ;
        RECT 604.950 86.400 619.050 87.450 ;
        RECT 604.950 85.950 607.050 86.400 ;
        RECT 616.950 85.950 619.050 86.400 ;
        RECT 634.950 87.450 637.050 88.050 ;
        RECT 649.800 87.450 651.900 88.050 ;
        RECT 634.950 86.400 651.900 87.450 ;
        RECT 634.950 85.950 637.050 86.400 ;
        RECT 649.800 85.950 651.900 86.400 ;
        RECT 653.100 87.450 655.200 88.050 ;
        RECT 682.950 87.450 685.050 88.050 ;
        RECT 700.950 87.450 703.050 88.050 ;
        RECT 766.950 87.600 769.050 89.700 ;
        RECT 787.950 88.500 790.050 90.600 ;
        RECT 653.100 86.400 703.050 87.450 ;
        RECT 653.100 85.950 655.200 86.400 ;
        RECT 682.950 85.950 685.050 86.400 ;
        RECT 700.950 85.950 703.050 86.400 ;
        RECT 61.950 84.450 64.050 85.050 ;
        RECT 85.950 84.450 88.050 85.050 ;
        RECT 61.950 83.400 88.050 84.450 ;
        RECT 61.950 82.950 64.050 83.400 ;
        RECT 85.950 82.950 88.050 83.400 ;
        RECT 94.950 82.950 100.050 85.050 ;
        RECT 109.950 84.450 112.050 85.050 ;
        RECT 151.950 84.450 154.050 85.050 ;
        RECT 193.950 84.450 196.050 85.050 ;
        RECT 109.950 83.400 196.050 84.450 ;
        RECT 109.950 82.950 112.050 83.400 ;
        RECT 151.950 82.950 154.050 83.400 ;
        RECT 193.950 82.950 196.050 83.400 ;
        RECT 383.100 84.450 388.050 85.050 ;
        RECT 490.800 84.450 492.900 85.050 ;
        RECT 383.100 83.400 492.900 84.450 ;
        RECT 383.100 82.950 388.050 83.400 ;
        RECT 490.800 82.950 492.900 83.400 ;
        RECT 494.100 84.450 496.200 85.050 ;
        RECT 499.950 84.450 502.050 85.050 ;
        RECT 494.100 83.400 502.050 84.450 ;
        RECT 494.100 82.950 496.200 83.400 ;
        RECT 499.950 82.950 502.050 83.400 ;
        RECT 541.950 84.450 547.050 85.050 ;
        RECT 556.950 84.450 559.050 85.050 ;
        RECT 635.400 84.450 636.450 85.950 ;
        RECT 541.950 83.400 636.450 84.450 ;
        RECT 652.950 84.450 655.050 85.050 ;
        RECT 664.950 84.450 667.050 85.050 ;
        RECT 652.950 83.400 667.050 84.450 ;
        RECT 541.950 82.950 547.050 83.400 ;
        RECT 556.950 82.950 559.050 83.400 ;
        RECT 652.950 82.950 655.050 83.400 ;
        RECT 664.950 82.950 667.050 83.400 ;
        RECT 679.950 84.450 682.050 85.050 ;
        RECT 715.950 84.450 718.050 85.050 ;
        RECT 679.950 83.400 718.050 84.450 ;
        RECT 679.950 82.950 682.050 83.400 ;
        RECT 715.950 82.950 718.050 83.400 ;
        RECT 751.950 84.450 754.050 85.050 ;
        RECT 874.950 84.450 877.050 85.050 ;
        RECT 751.950 83.400 877.050 84.450 ;
        RECT 751.950 82.950 754.050 83.400 ;
        RECT 874.950 82.950 877.050 83.400 ;
        RECT 883.950 82.950 889.050 85.050 ;
        RECT 16.950 81.450 19.050 82.050 ;
        RECT 31.950 81.450 34.050 82.050 ;
        RECT 16.950 80.400 34.050 81.450 ;
        RECT 16.950 79.950 19.050 80.400 ;
        RECT 31.950 79.950 34.050 80.400 ;
        RECT 154.950 81.450 157.050 82.050 ;
        RECT 187.950 81.450 190.050 82.050 ;
        RECT 223.950 81.450 226.050 82.050 ;
        RECT 235.950 81.450 238.050 82.050 ;
        RECT 280.950 81.450 283.050 82.050 ;
        RECT 154.950 80.400 283.050 81.450 ;
        RECT 154.950 79.950 157.050 80.400 ;
        RECT 187.950 79.950 190.050 80.400 ;
        RECT 223.950 79.950 226.050 80.400 ;
        RECT 235.950 79.950 238.050 80.400 ;
        RECT 280.950 79.950 283.050 80.400 ;
        RECT 304.950 81.450 307.050 82.050 ;
        RECT 322.950 81.450 325.050 82.050 ;
        RECT 304.950 80.400 325.050 81.450 ;
        RECT 304.950 79.950 307.050 80.400 ;
        RECT 322.950 79.950 325.050 80.400 ;
        RECT 343.950 81.450 346.050 82.050 ;
        RECT 370.950 81.450 373.050 82.050 ;
        RECT 712.950 81.450 715.050 82.050 ;
        RECT 343.950 80.400 715.050 81.450 ;
        RECT 343.950 79.950 346.050 80.400 ;
        RECT 370.950 79.950 373.050 80.400 ;
        RECT 712.950 79.950 715.050 80.400 ;
        RECT 718.950 81.450 721.050 82.050 ;
        RECT 724.950 81.450 727.050 82.050 ;
        RECT 718.950 80.400 727.050 81.450 ;
        RECT 718.950 79.950 721.050 80.400 ;
        RECT 724.950 79.950 727.050 80.400 ;
        RECT 790.950 81.450 793.050 82.050 ;
        RECT 844.950 81.450 847.050 82.050 ;
        RECT 790.950 80.400 847.050 81.450 ;
        RECT 790.950 79.950 793.050 80.400 ;
        RECT 844.950 79.950 847.050 80.400 ;
        RECT 32.400 78.450 33.450 79.950 ;
        RECT 61.950 78.450 64.050 79.050 ;
        RECT 32.400 77.400 64.050 78.450 ;
        RECT 61.950 76.950 64.050 77.400 ;
        RECT 298.950 78.450 301.050 79.050 ;
        RECT 478.950 78.450 481.050 79.050 ;
        RECT 562.950 78.450 565.050 79.050 ;
        RECT 601.950 78.450 604.050 79.050 ;
        RECT 298.950 77.400 477.450 78.450 ;
        RECT 298.950 76.950 301.050 77.400 ;
        RECT 40.950 75.450 43.050 76.050 ;
        RECT 91.950 75.450 94.050 76.050 ;
        RECT 103.950 75.450 106.050 76.050 ;
        RECT 40.950 74.400 106.050 75.450 ;
        RECT 40.950 73.950 43.050 74.400 ;
        RECT 91.950 73.950 94.050 74.400 ;
        RECT 103.950 73.950 106.050 74.400 ;
        RECT 127.950 75.450 130.050 76.050 ;
        RECT 139.800 75.450 141.900 76.050 ;
        RECT 127.950 74.400 141.900 75.450 ;
        RECT 127.950 73.950 130.050 74.400 ;
        RECT 139.800 73.950 141.900 74.400 ;
        RECT 143.100 75.450 145.200 76.050 ;
        RECT 160.950 75.450 163.050 76.050 ;
        RECT 143.100 74.400 163.050 75.450 ;
        RECT 143.100 73.950 145.200 74.400 ;
        RECT 160.950 73.950 163.050 74.400 ;
        RECT 220.950 75.450 223.050 76.050 ;
        RECT 232.950 75.450 235.050 76.050 ;
        RECT 220.950 74.400 235.050 75.450 ;
        RECT 220.950 73.950 223.050 74.400 ;
        RECT 232.950 73.950 235.050 74.400 ;
        RECT 268.950 75.450 271.050 76.050 ;
        RECT 307.950 75.450 310.050 76.050 ;
        RECT 268.950 74.400 310.050 75.450 ;
        RECT 268.950 73.950 271.050 74.400 ;
        RECT 307.950 73.950 310.050 74.400 ;
        RECT 328.950 75.450 331.050 76.050 ;
        RECT 476.400 75.450 477.450 77.400 ;
        RECT 478.950 77.400 604.050 78.450 ;
        RECT 478.950 76.950 481.050 77.400 ;
        RECT 562.950 76.950 565.050 77.400 ;
        RECT 601.950 76.950 604.050 77.400 ;
        RECT 676.950 78.450 679.050 79.050 ;
        RECT 685.950 78.450 688.050 79.050 ;
        RECT 676.950 77.400 688.050 78.450 ;
        RECT 676.950 76.950 679.050 77.400 ;
        RECT 685.950 76.950 688.050 77.400 ;
        RECT 577.950 75.450 580.050 76.050 ;
        RECT 592.950 75.450 595.050 76.050 ;
        RECT 622.950 75.450 625.050 76.050 ;
        RECT 328.950 74.400 474.450 75.450 ;
        RECT 476.400 74.400 576.450 75.450 ;
        RECT 328.950 73.950 331.050 74.400 ;
        RECT 13.950 72.450 16.050 73.050 ;
        RECT 49.950 72.450 52.050 73.050 ;
        RECT 13.950 71.400 52.050 72.450 ;
        RECT 13.950 70.950 16.050 71.400 ;
        RECT 49.950 70.950 52.050 71.400 ;
        RECT 154.950 72.450 157.050 73.050 ;
        RECT 184.950 72.450 187.050 73.050 ;
        RECT 154.950 71.400 187.050 72.450 ;
        RECT 473.400 72.450 474.450 74.400 ;
        RECT 550.950 72.450 553.050 73.050 ;
        RECT 473.400 71.400 553.050 72.450 ;
        RECT 575.400 72.450 576.450 74.400 ;
        RECT 577.950 74.400 625.050 75.450 ;
        RECT 577.950 73.950 580.050 74.400 ;
        RECT 592.950 73.950 595.050 74.400 ;
        RECT 622.950 73.950 625.050 74.400 ;
        RECT 637.950 75.450 640.050 76.050 ;
        RECT 763.950 75.450 766.050 76.050 ;
        RECT 637.950 74.400 766.050 75.450 ;
        RECT 637.950 73.950 640.050 74.400 ;
        RECT 763.950 73.950 766.050 74.400 ;
        RECT 583.950 72.450 586.050 73.050 ;
        RECT 575.400 71.400 586.050 72.450 ;
        RECT 601.950 72.450 604.050 73.050 ;
        RECT 664.950 72.450 667.050 73.050 ;
        RECT 601.950 71.400 667.050 72.450 ;
        RECT 784.950 72.450 787.050 73.050 ;
        RECT 796.950 72.450 799.050 73.050 ;
        RECT 784.950 71.400 799.050 72.450 ;
        RECT 853.950 72.450 856.050 73.050 ;
        RECT 865.950 72.450 868.050 73.050 ;
        RECT 853.950 71.400 868.050 72.450 ;
        RECT 154.950 70.950 157.050 71.400 ;
        RECT 184.950 70.950 187.050 71.400 ;
        RECT 31.950 69.450 34.050 70.050 ;
        RECT 64.950 69.450 67.050 70.050 ;
        RECT 31.950 68.400 67.050 69.450 ;
        RECT 31.950 67.950 34.050 68.400 ;
        RECT 64.950 67.950 67.050 68.400 ;
        RECT 73.950 69.450 76.050 70.050 ;
        RECT 103.950 69.450 106.050 70.050 ;
        RECT 148.950 69.450 151.050 70.050 ;
        RECT 163.950 69.450 166.050 70.050 ;
        RECT 73.950 68.400 166.050 69.450 ;
        RECT 73.950 67.950 76.050 68.400 ;
        RECT 103.950 67.950 106.050 68.400 ;
        RECT 148.950 67.950 151.050 68.400 ;
        RECT 163.950 67.950 166.050 68.400 ;
        RECT 172.950 69.450 175.050 70.050 ;
        RECT 208.950 69.450 211.050 70.050 ;
        RECT 172.950 68.400 211.050 69.450 ;
        RECT 226.950 68.400 229.050 70.500 ;
        RECT 247.950 69.300 250.050 71.400 ;
        RECT 172.950 67.950 175.050 68.400 ;
        RECT 208.950 67.950 211.050 68.400 ;
        RECT 49.950 66.450 52.050 67.050 ;
        RECT 55.950 66.450 58.050 67.050 ;
        RECT 49.950 65.400 58.050 66.450 ;
        RECT 49.950 64.950 52.050 65.400 ;
        RECT 55.950 64.950 58.050 65.400 ;
        RECT 34.950 61.950 37.050 64.050 ;
        RECT 40.950 61.950 43.050 64.050 ;
        RECT 16.950 60.450 19.050 61.050 ;
        RECT 28.950 60.450 31.050 61.050 ;
        RECT 16.950 59.400 31.050 60.450 ;
        RECT 16.950 58.950 19.050 59.400 ;
        RECT 28.950 58.950 31.050 59.400 ;
        RECT 34.950 58.950 37.050 60.750 ;
        RECT 40.950 58.950 43.050 60.750 ;
        RECT 55.950 58.950 58.050 61.050 ;
        RECT 64.950 58.950 67.050 64.050 ;
        RECT 82.950 61.950 85.050 67.050 ;
        RECT 115.950 63.450 118.050 64.050 ;
        RECT 124.950 63.450 127.050 64.050 ;
        RECT 115.950 62.400 127.050 63.450 ;
        RECT 115.950 61.950 118.050 62.400 ;
        RECT 124.950 61.950 127.050 62.400 ;
        RECT 142.950 61.950 145.050 64.050 ;
        RECT 148.950 61.950 151.050 64.050 ;
        RECT 160.950 61.950 163.050 64.050 ;
        RECT 184.950 61.950 187.050 64.050 ;
        RECT 190.950 61.950 193.050 64.050 ;
        RECT 208.950 61.950 211.050 64.050 ;
        RECT 214.950 61.950 217.050 64.050 ;
        RECT 82.950 58.950 85.050 60.750 ;
        RECT 94.950 60.450 99.000 61.050 ;
        RECT 100.950 60.450 103.050 61.050 ;
        RECT 94.950 59.400 103.050 60.450 ;
        RECT 94.950 58.950 99.000 59.400 ;
        RECT 100.950 58.950 103.050 59.400 ;
        RECT 109.950 58.950 112.050 61.050 ;
        RECT 124.950 58.950 127.050 60.750 ;
        RECT 142.950 58.950 145.050 60.750 ;
        RECT 148.950 58.950 151.050 60.750 ;
        RECT 160.950 58.950 163.050 60.750 ;
        RECT 169.950 60.450 172.050 61.050 ;
        RECT 178.950 60.450 181.050 61.050 ;
        RECT 169.950 59.400 181.050 60.450 ;
        RECT 169.950 58.950 172.050 59.400 ;
        RECT 178.950 58.950 181.050 59.400 ;
        RECT 184.950 58.950 187.050 60.750 ;
        RECT 190.950 58.950 193.050 60.750 ;
        RECT 208.950 58.950 211.050 60.750 ;
        RECT 214.950 58.950 217.050 60.750 ;
        RECT 223.950 58.950 226.050 61.050 ;
        RECT 16.950 55.950 19.050 57.750 ;
        RECT 31.950 56.250 34.050 58.050 ;
        RECT 37.950 56.250 40.050 58.050 ;
        RECT 61.950 57.750 63.750 58.050 ;
        RECT 55.950 55.950 58.050 57.750 ;
        RECT 61.950 56.250 64.050 57.750 ;
        RECT 64.950 56.250 67.050 57.750 ;
        RECT 85.950 56.250 88.050 58.050 ;
        RECT 104.250 57.750 106.050 58.050 ;
        RECT 100.950 56.250 103.050 57.750 ;
        RECT 103.950 56.250 106.050 57.750 ;
        RECT 65.250 55.950 67.050 56.250 ;
        RECT 100.950 55.950 102.750 56.250 ;
        RECT 109.950 55.950 112.050 57.750 ;
        RECT 127.950 56.250 130.050 58.050 ;
        RECT 145.950 56.250 148.050 58.050 ;
        RECT 163.950 56.250 166.050 58.050 ;
        RECT 169.950 55.950 172.050 57.750 ;
        RECT 187.950 56.250 190.050 58.050 ;
        RECT 205.950 56.250 208.050 58.050 ;
        RECT 211.950 56.250 214.050 58.050 ;
        RECT 223.950 55.950 226.050 57.750 ;
        RECT 13.950 53.250 16.050 55.050 ;
        RECT 19.950 53.250 22.050 55.050 ;
        RECT 31.950 52.950 34.050 55.050 ;
        RECT 37.950 54.450 40.050 55.050 ;
        RECT 49.950 54.450 52.050 55.050 ;
        RECT 37.950 53.400 52.050 54.450 ;
        RECT 37.950 52.950 40.050 53.400 ;
        RECT 49.950 52.950 52.050 53.400 ;
        RECT 61.950 52.950 64.050 55.050 ;
        RECT 85.950 52.950 88.050 55.050 ;
        RECT 103.950 52.950 106.050 55.050 ;
        RECT 112.950 54.450 115.050 55.050 ;
        RECT 127.950 54.450 130.050 55.050 ;
        RECT 112.950 53.400 130.050 54.450 ;
        RECT 112.950 52.950 115.050 53.400 ;
        RECT 127.950 52.950 130.050 53.400 ;
        RECT 145.950 54.450 148.050 55.050 ;
        RECT 154.950 54.450 157.050 55.050 ;
        RECT 145.950 53.400 157.050 54.450 ;
        RECT 145.950 52.950 148.050 53.400 ;
        RECT 154.950 52.950 157.050 53.400 ;
        RECT 163.950 52.950 166.050 55.050 ;
        RECT 187.950 54.450 190.050 55.050 ;
        RECT 192.000 54.450 196.050 55.050 ;
        RECT 187.950 53.400 196.050 54.450 ;
        RECT 187.950 52.950 190.050 53.400 ;
        RECT 192.000 52.950 196.050 53.400 ;
        RECT 205.950 52.950 208.050 55.050 ;
        RECT 211.950 54.450 214.050 55.050 ;
        RECT 220.950 54.450 223.050 55.050 ;
        RECT 211.950 53.400 223.050 54.450 ;
        RECT 211.950 52.950 214.050 53.400 ;
        RECT 220.950 52.950 223.050 53.400 ;
        RECT 13.950 49.950 16.050 52.050 ;
        RECT 19.950 49.950 22.050 52.050 ;
        RECT 217.950 51.450 220.050 52.050 ;
        RECT 223.950 51.450 226.050 52.050 ;
        RECT 217.950 50.400 226.050 51.450 ;
        RECT 217.950 49.950 220.050 50.400 ;
        RECT 223.950 49.950 226.050 50.400 ;
        RECT 91.950 43.950 94.050 49.050 ;
        RECT 227.700 48.600 228.900 68.400 ;
        RECT 247.950 65.700 249.150 69.300 ;
        RECT 283.950 68.400 286.050 70.500 ;
        RECT 304.950 69.300 307.050 71.400 ;
        RECT 247.950 63.600 250.050 65.700 ;
        RECT 232.950 58.950 235.050 61.050 ;
        RECT 232.950 55.950 235.050 57.750 ;
        RECT 232.950 51.450 235.050 52.050 ;
        RECT 241.950 51.450 244.050 52.050 ;
        RECT 232.950 50.400 244.050 51.450 ;
        RECT 232.950 49.950 235.050 50.400 ;
        RECT 241.950 49.950 244.050 50.400 ;
        RECT 247.950 48.600 249.150 63.600 ;
        RECT 256.950 63.450 259.050 64.050 ;
        RECT 265.950 63.450 268.050 64.050 ;
        RECT 256.950 62.400 268.050 63.450 ;
        RECT 256.950 61.950 259.050 62.400 ;
        RECT 265.950 61.950 268.050 62.400 ;
        RECT 271.950 61.950 274.050 64.050 ;
        RECT 265.950 58.950 268.050 60.750 ;
        RECT 271.950 58.950 274.050 60.750 ;
        RECT 280.950 58.950 283.050 61.050 ;
        RECT 250.950 56.250 253.050 58.050 ;
        RECT 268.950 56.250 271.050 58.050 ;
        RECT 280.950 55.950 283.050 57.750 ;
        RECT 250.950 52.950 253.050 55.050 ;
        RECT 256.950 54.450 259.050 55.050 ;
        RECT 268.950 54.450 271.050 55.050 ;
        RECT 256.950 53.400 271.050 54.450 ;
        RECT 256.950 52.950 259.050 53.400 ;
        RECT 268.950 52.950 271.050 53.400 ;
        RECT 226.950 46.500 229.050 48.600 ;
        RECT 247.950 46.500 250.050 48.600 ;
        RECT 253.950 48.450 259.050 49.050 ;
        RECT 277.950 48.450 280.050 49.050 ;
        RECT 284.700 48.600 285.900 68.400 ;
        RECT 304.950 65.700 306.150 69.300 ;
        RECT 322.950 66.450 325.050 67.050 ;
        RECT 343.950 66.450 346.050 67.050 ;
        RECT 304.950 63.600 307.050 65.700 ;
        RECT 322.950 65.400 346.050 66.450 ;
        RECT 322.950 64.950 325.050 65.400 ;
        RECT 343.950 64.950 346.050 65.400 ;
        RECT 385.950 64.950 388.050 70.050 ;
        RECT 391.950 69.450 394.050 70.050 ;
        RECT 415.950 69.450 418.050 70.050 ;
        RECT 391.950 68.400 418.050 69.450 ;
        RECT 436.950 68.400 439.050 70.500 ;
        RECT 457.950 69.300 460.050 71.400 ;
        RECT 550.950 70.950 553.050 71.400 ;
        RECT 583.950 70.950 586.050 71.400 ;
        RECT 472.950 69.450 475.050 70.050 ;
        RECT 523.950 69.450 526.050 70.050 ;
        RECT 391.950 67.950 394.050 68.400 ;
        RECT 415.950 67.950 418.050 68.400 ;
        RECT 289.950 58.950 292.050 61.050 ;
        RECT 289.950 55.950 292.050 57.750 ;
        RECT 304.950 48.600 306.150 63.600 ;
        RECT 322.950 58.950 325.050 61.050 ;
        RECT 328.950 58.950 331.050 64.050 ;
        RECT 391.950 61.950 394.050 64.050 ;
        RECT 397.950 63.450 400.050 64.050 ;
        RECT 409.950 63.450 412.050 64.050 ;
        RECT 397.950 62.400 412.050 63.450 ;
        RECT 397.950 61.950 400.050 62.400 ;
        RECT 409.950 61.950 412.050 62.400 ;
        RECT 415.950 61.950 418.050 64.050 ;
        RECT 334.950 58.950 337.050 61.050 ;
        RECT 355.950 58.950 358.050 61.050 ;
        RECT 376.950 60.450 379.050 61.050 ;
        RECT 385.950 60.450 388.050 61.050 ;
        RECT 376.950 59.400 388.050 60.450 ;
        RECT 376.950 58.950 379.050 59.400 ;
        RECT 385.950 58.950 388.050 59.400 ;
        RECT 391.950 58.950 394.050 60.750 ;
        RECT 397.950 58.950 400.050 60.750 ;
        RECT 415.950 58.950 418.050 60.750 ;
        RECT 421.950 58.950 427.050 61.050 ;
        RECT 430.950 58.950 436.050 61.050 ;
        RECT 307.950 56.250 310.050 58.050 ;
        RECT 322.950 55.950 325.050 57.750 ;
        RECT 328.950 55.950 331.050 57.750 ;
        RECT 334.950 55.950 337.050 57.750 ;
        RECT 349.950 56.250 352.050 58.050 ;
        RECT 355.950 55.950 358.050 57.750 ;
        RECT 370.950 56.250 373.050 58.050 ;
        RECT 376.950 55.950 379.050 57.750 ;
        RECT 394.950 56.250 397.050 58.050 ;
        RECT 400.950 56.250 403.050 58.050 ;
        RECT 418.950 56.250 421.050 58.050 ;
        RECT 424.950 55.950 427.050 57.750 ;
        RECT 433.950 55.950 436.050 57.750 ;
        RECT 307.950 54.450 310.050 55.050 ;
        RECT 319.950 54.450 322.050 55.050 ;
        RECT 307.950 53.400 322.050 54.450 ;
        RECT 307.950 52.950 310.050 53.400 ;
        RECT 319.950 52.950 322.050 53.400 ;
        RECT 325.950 53.250 328.050 55.050 ;
        RECT 331.950 53.250 334.050 55.050 ;
        RECT 349.950 52.950 352.050 55.050 ;
        RECT 370.950 52.950 373.050 55.050 ;
        RECT 394.950 52.950 397.050 55.050 ;
        RECT 325.950 49.950 328.050 52.050 ;
        RECT 331.950 49.950 334.050 52.050 ;
        RECT 400.950 49.950 403.050 55.050 ;
        RECT 406.950 54.450 409.050 55.050 ;
        RECT 412.950 54.450 415.050 55.050 ;
        RECT 406.950 53.400 415.050 54.450 ;
        RECT 406.950 52.950 409.050 53.400 ;
        RECT 412.950 52.950 415.050 53.400 ;
        RECT 418.950 52.950 421.050 55.050 ;
        RECT 253.950 47.400 280.050 48.450 ;
        RECT 253.950 46.950 259.050 47.400 ;
        RECT 277.950 46.950 280.050 47.400 ;
        RECT 283.950 46.500 286.050 48.600 ;
        RECT 304.950 46.500 307.050 48.600 ;
        RECT 349.950 48.450 352.050 49.050 ;
        RECT 370.950 48.450 373.050 49.050 ;
        RECT 349.950 47.400 373.050 48.450 ;
        RECT 349.950 46.950 352.050 47.400 ;
        RECT 370.950 46.950 373.050 47.400 ;
        RECT 385.950 48.450 388.050 49.050 ;
        RECT 394.950 48.450 397.050 49.050 ;
        RECT 403.950 48.450 406.050 49.050 ;
        RECT 385.950 47.400 406.050 48.450 ;
        RECT 385.950 46.950 388.050 47.400 ;
        RECT 394.950 46.950 397.050 47.400 ;
        RECT 403.950 46.950 406.050 47.400 ;
        RECT 409.950 46.950 415.050 49.050 ;
        RECT 418.950 48.450 421.050 49.050 ;
        RECT 430.950 48.450 433.050 49.050 ;
        RECT 437.700 48.600 438.900 68.400 ;
        RECT 457.950 65.700 459.150 69.300 ;
        RECT 472.950 68.400 526.050 69.450 ;
        RECT 568.950 68.400 571.050 70.500 ;
        RECT 589.950 69.300 592.050 71.400 ;
        RECT 601.950 70.950 604.050 71.400 ;
        RECT 664.950 70.950 667.050 71.400 ;
        RECT 604.950 69.450 607.050 70.050 ;
        RECT 655.950 69.450 658.050 70.050 ;
        RECT 472.950 67.950 475.050 68.400 ;
        RECT 523.950 67.950 526.050 68.400 ;
        RECT 457.950 63.600 460.050 65.700 ;
        RECT 442.950 58.950 445.050 61.050 ;
        RECT 442.950 55.950 445.050 57.750 ;
        RECT 457.950 48.600 459.150 63.600 ;
        RECT 484.950 63.450 487.050 64.050 ;
        RECT 499.950 63.450 502.050 64.050 ;
        RECT 484.950 62.400 502.050 63.450 ;
        RECT 484.950 61.950 487.050 62.400 ;
        RECT 499.950 61.950 502.050 62.400 ;
        RECT 517.950 61.950 523.050 64.050 ;
        RECT 556.950 61.950 559.050 64.050 ;
        RECT 463.950 60.450 466.050 61.050 ;
        RECT 472.950 60.450 475.050 61.050 ;
        RECT 463.950 59.400 475.050 60.450 ;
        RECT 463.950 58.950 466.050 59.400 ;
        RECT 472.950 58.950 475.050 59.400 ;
        RECT 478.950 58.950 481.050 61.050 ;
        RECT 499.950 58.950 502.050 60.750 ;
        RECT 517.950 58.950 520.050 60.750 ;
        RECT 523.950 60.450 526.050 61.050 ;
        RECT 538.950 60.450 541.050 61.050 ;
        RECT 523.950 59.400 541.050 60.450 ;
        RECT 523.950 58.950 526.050 59.400 ;
        RECT 538.950 58.950 541.050 59.400 ;
        RECT 556.950 58.950 559.050 60.750 ;
        RECT 562.950 58.950 568.050 61.050 ;
        RECT 460.950 56.250 463.050 58.050 ;
        RECT 478.950 55.950 481.050 57.750 ;
        RECT 502.950 56.250 505.050 58.050 ;
        RECT 520.950 56.250 523.050 58.050 ;
        RECT 538.950 55.950 541.050 57.750 ;
        RECT 553.950 56.250 556.050 58.050 ;
        RECT 565.950 55.950 568.050 57.750 ;
        RECT 460.950 52.950 466.050 55.050 ;
        RECT 475.950 53.250 478.050 55.050 ;
        RECT 481.950 53.250 484.050 55.050 ;
        RECT 535.950 53.250 538.050 55.050 ;
        RECT 541.950 53.250 544.050 55.050 ;
        RECT 553.950 52.950 556.050 55.050 ;
        RECT 475.950 49.950 478.050 52.050 ;
        RECT 481.950 49.950 484.050 52.050 ;
        RECT 418.950 47.400 433.050 48.450 ;
        RECT 418.950 46.950 421.050 47.400 ;
        RECT 430.950 46.950 433.050 47.400 ;
        RECT 436.950 46.500 439.050 48.600 ;
        RECT 457.950 46.500 460.050 48.600 ;
        RECT 487.950 48.450 490.050 49.050 ;
        RECT 487.950 47.400 525.450 48.450 ;
        RECT 487.950 46.950 490.050 47.400 ;
        RECT 100.950 45.450 103.050 46.050 ;
        RECT 115.950 45.450 118.050 46.050 ;
        RECT 154.950 45.450 157.050 46.050 ;
        RECT 100.950 44.400 118.050 45.450 ;
        RECT 100.950 43.950 103.050 44.400 ;
        RECT 115.950 43.950 118.050 44.400 ;
        RECT 119.400 44.400 157.050 45.450 ;
        RECT 73.950 42.450 76.050 43.050 ;
        RECT 119.400 42.450 120.450 44.400 ;
        RECT 154.950 43.950 157.050 44.400 ;
        RECT 232.950 45.450 235.050 46.050 ;
        RECT 241.950 45.450 244.050 46.050 ;
        RECT 232.950 44.400 244.050 45.450 ;
        RECT 232.950 43.950 235.050 44.400 ;
        RECT 241.950 43.950 244.050 44.400 ;
        RECT 289.950 45.450 292.050 46.050 ;
        RECT 298.950 45.450 301.050 46.050 ;
        RECT 289.950 44.400 301.050 45.450 ;
        RECT 289.950 43.950 292.050 44.400 ;
        RECT 298.950 43.950 301.050 44.400 ;
        RECT 325.950 45.450 328.050 46.050 ;
        RECT 334.950 45.450 337.050 46.050 ;
        RECT 325.950 44.400 337.050 45.450 ;
        RECT 325.950 43.950 328.050 44.400 ;
        RECT 334.950 43.950 337.050 44.400 ;
        RECT 343.950 45.450 346.050 46.050 ;
        RECT 427.950 45.450 430.050 46.050 ;
        RECT 343.950 44.400 430.050 45.450 ;
        RECT 343.950 43.950 346.050 44.400 ;
        RECT 427.950 43.950 430.050 44.400 ;
        RECT 469.950 45.450 472.050 46.050 ;
        RECT 520.950 45.450 523.050 46.050 ;
        RECT 469.950 44.400 523.050 45.450 ;
        RECT 524.400 45.450 525.450 47.400 ;
        RECT 535.950 46.950 538.050 52.050 ;
        RECT 541.950 49.950 544.050 52.050 ;
        RECT 569.700 48.600 570.900 68.400 ;
        RECT 589.950 65.700 591.150 69.300 ;
        RECT 604.950 68.400 658.050 69.450 ;
        RECT 673.950 68.400 676.050 70.500 ;
        RECT 694.950 69.300 697.050 71.400 ;
        RECT 784.950 70.950 787.050 71.400 ;
        RECT 796.950 70.950 799.050 71.400 ;
        RECT 712.950 69.450 715.050 70.050 ;
        RECT 751.950 69.450 754.050 70.050 ;
        RECT 604.950 67.950 607.050 68.400 ;
        RECT 655.950 67.950 658.050 68.400 ;
        RECT 664.950 66.450 667.050 67.050 ;
        RECT 670.950 66.450 673.050 67.050 ;
        RECT 589.950 63.600 592.050 65.700 ;
        RECT 664.950 65.400 673.050 66.450 ;
        RECT 664.950 64.950 667.050 65.400 ;
        RECT 670.950 64.950 673.050 65.400 ;
        RECT 574.950 58.950 577.050 61.050 ;
        RECT 574.950 55.950 577.050 57.750 ;
        RECT 589.950 48.600 591.150 63.600 ;
        RECT 610.950 61.950 613.050 64.050 ;
        RECT 616.950 61.950 619.050 64.050 ;
        RECT 655.950 61.950 658.050 64.050 ;
        RECT 661.950 61.950 664.050 64.050 ;
        RECT 610.950 58.950 613.050 60.750 ;
        RECT 616.950 58.950 619.050 60.750 ;
        RECT 622.950 60.450 625.050 61.050 ;
        RECT 634.950 60.450 637.050 61.050 ;
        RECT 622.950 59.400 637.050 60.450 ;
        RECT 622.950 58.950 625.050 59.400 ;
        RECT 634.950 58.950 637.050 59.400 ;
        RECT 655.950 58.950 658.050 60.750 ;
        RECT 661.950 58.950 664.050 60.750 ;
        RECT 670.950 58.950 673.050 61.050 ;
        RECT 592.950 56.250 595.050 58.050 ;
        RECT 613.950 56.250 616.050 58.050 ;
        RECT 619.950 56.250 622.050 58.050 ;
        RECT 634.950 55.950 637.050 57.750 ;
        RECT 658.950 56.250 661.050 58.050 ;
        RECT 664.950 56.250 667.050 58.050 ;
        RECT 670.950 55.950 673.050 57.750 ;
        RECT 592.950 52.950 595.050 55.050 ;
        RECT 613.950 52.950 616.050 55.050 ;
        RECT 619.950 52.950 622.050 55.050 ;
        RECT 631.950 53.250 634.050 55.050 ;
        RECT 637.950 53.250 640.050 55.050 ;
        RECT 658.950 52.950 661.050 55.050 ;
        RECT 664.950 52.950 667.050 55.050 ;
        RECT 631.950 49.950 634.050 52.050 ;
        RECT 637.950 49.950 640.050 52.050 ;
        RECT 674.700 48.600 675.900 68.400 ;
        RECT 694.950 65.700 696.150 69.300 ;
        RECT 712.950 68.400 754.050 69.450 ;
        RECT 712.950 67.950 715.050 68.400 ;
        RECT 751.950 67.950 754.050 68.400 ;
        RECT 793.950 69.450 796.050 70.050 ;
        RECT 808.950 69.450 811.050 70.050 ;
        RECT 793.950 68.400 811.050 69.450 ;
        RECT 814.950 69.300 817.050 71.400 ;
        RECT 853.950 70.950 856.050 71.400 ;
        RECT 865.950 70.950 868.050 71.400 ;
        RECT 793.950 67.950 796.050 68.400 ;
        RECT 808.950 67.950 811.050 68.400 ;
        RECT 815.850 65.700 817.050 69.300 ;
        RECT 820.950 69.450 823.050 70.050 ;
        RECT 829.950 69.450 832.050 70.050 ;
        RECT 820.950 68.400 832.050 69.450 ;
        RECT 835.950 68.400 838.050 70.500 ;
        RECT 841.950 69.450 844.050 70.050 ;
        RECT 862.950 69.450 865.050 70.050 ;
        RECT 841.950 68.400 865.050 69.450 ;
        RECT 820.950 67.950 823.050 68.400 ;
        RECT 829.950 67.950 832.050 68.400 ;
        RECT 694.950 63.600 697.050 65.700 ;
        RECT 679.950 58.950 682.050 61.050 ;
        RECT 679.950 55.950 682.050 57.750 ;
        RECT 679.950 51.450 682.050 52.050 ;
        RECT 688.950 51.450 691.050 52.050 ;
        RECT 679.950 50.400 691.050 51.450 ;
        RECT 679.950 49.950 682.050 50.400 ;
        RECT 688.950 49.950 691.050 50.400 ;
        RECT 694.950 48.600 696.150 63.600 ;
        RECT 715.950 61.950 718.050 64.050 ;
        RECT 775.950 61.950 778.050 64.050 ;
        RECT 781.950 61.950 784.050 64.050 ;
        RECT 799.950 61.950 802.050 64.050 ;
        RECT 805.950 61.950 811.050 64.050 ;
        RECT 814.950 63.600 817.050 65.700 ;
        RECT 715.950 58.950 718.050 60.750 ;
        RECT 721.950 60.450 724.050 61.050 ;
        RECT 733.950 60.450 736.050 61.050 ;
        RECT 721.950 59.400 736.050 60.450 ;
        RECT 721.950 58.950 724.050 59.400 ;
        RECT 733.950 58.950 736.050 59.400 ;
        RECT 757.950 60.450 760.050 61.050 ;
        RECT 769.950 60.450 772.050 61.050 ;
        RECT 757.950 59.400 772.050 60.450 ;
        RECT 757.950 58.950 760.050 59.400 ;
        RECT 769.950 58.950 772.050 59.400 ;
        RECT 775.950 58.950 778.050 60.750 ;
        RECT 781.950 58.950 784.050 60.750 ;
        RECT 799.950 58.950 802.050 60.750 ;
        RECT 805.950 58.950 808.050 60.750 ;
        RECT 697.950 56.250 700.050 58.050 ;
        RECT 712.950 56.250 715.050 58.050 ;
        RECT 733.950 55.950 736.050 57.750 ;
        RECT 751.950 56.250 754.050 58.050 ;
        RECT 757.950 55.950 760.050 57.750 ;
        RECT 778.950 56.250 781.050 58.050 ;
        RECT 784.950 56.250 787.050 58.050 ;
        RECT 802.950 56.250 805.050 58.050 ;
        RECT 811.950 56.250 814.050 58.050 ;
        RECT 697.950 54.450 700.050 55.050 ;
        RECT 706.950 54.450 709.050 55.050 ;
        RECT 697.950 53.400 709.050 54.450 ;
        RECT 697.950 52.950 700.050 53.400 ;
        RECT 706.950 52.950 709.050 53.400 ;
        RECT 712.950 52.950 715.050 55.050 ;
        RECT 730.950 53.250 733.050 55.050 ;
        RECT 736.950 53.250 739.050 55.050 ;
        RECT 751.950 52.950 754.050 55.050 ;
        RECT 772.950 54.450 777.000 55.050 ;
        RECT 778.950 54.450 781.050 55.050 ;
        RECT 772.950 53.400 781.050 54.450 ;
        RECT 772.950 52.950 777.000 53.400 ;
        RECT 778.950 52.950 781.050 53.400 ;
        RECT 784.950 52.950 787.050 55.050 ;
        RECT 793.950 54.450 796.050 55.050 ;
        RECT 802.950 54.450 805.050 55.050 ;
        RECT 793.950 53.400 805.050 54.450 ;
        RECT 793.950 52.950 796.050 53.400 ;
        RECT 802.950 52.950 805.050 53.400 ;
        RECT 811.950 52.950 814.050 55.050 ;
        RECT 730.950 49.950 733.050 52.050 ;
        RECT 736.950 49.950 739.050 52.050 ;
        RECT 568.950 46.500 571.050 48.600 ;
        RECT 589.950 46.500 592.050 48.600 ;
        RECT 673.950 46.500 676.050 48.600 ;
        RECT 694.950 46.500 697.050 48.600 ;
        RECT 700.950 48.450 703.050 49.050 ;
        RECT 721.950 48.450 724.050 49.050 ;
        RECT 700.950 47.400 724.050 48.450 ;
        RECT 700.950 46.950 703.050 47.400 ;
        RECT 721.950 46.950 724.050 47.400 ;
        RECT 769.950 48.450 772.050 49.050 ;
        RECT 778.950 48.450 781.050 49.050 ;
        RECT 784.950 48.450 787.050 49.050 ;
        RECT 796.950 48.450 799.050 49.050 ;
        RECT 815.850 48.600 817.050 63.600 ;
        RECT 829.950 58.950 832.050 61.050 ;
        RECT 829.950 55.950 832.050 57.750 ;
        RECT 836.100 48.600 837.300 68.400 ;
        RECT 841.950 67.950 844.050 68.400 ;
        RECT 862.950 67.950 865.050 68.400 ;
        RECT 883.950 69.450 886.050 70.050 ;
        RECT 889.950 69.450 892.050 70.050 ;
        RECT 883.950 68.400 892.050 69.450 ;
        RECT 883.950 67.950 886.050 68.400 ;
        RECT 889.950 67.950 892.050 68.400 ;
        RECT 838.950 66.450 841.050 67.050 ;
        RECT 844.950 66.450 847.050 67.050 ;
        RECT 838.950 65.400 847.050 66.450 ;
        RECT 838.950 64.950 841.050 65.400 ;
        RECT 844.950 64.950 847.050 65.400 ;
        RECT 856.950 61.950 859.050 64.050 ;
        RECT 862.950 61.950 865.050 64.050 ;
        RECT 883.950 61.950 886.050 64.050 ;
        RECT 889.950 61.950 892.050 64.050 ;
        RECT 895.950 63.450 900.000 64.050 ;
        RECT 901.950 63.450 904.050 64.050 ;
        RECT 895.950 62.400 904.050 63.450 ;
        RECT 895.950 61.950 900.000 62.400 ;
        RECT 901.950 61.950 904.050 62.400 ;
        RECT 838.950 58.950 841.050 61.050 ;
        RECT 856.950 58.950 859.050 60.750 ;
        RECT 862.950 58.950 865.050 60.750 ;
        RECT 883.950 58.950 886.050 60.750 ;
        RECT 889.950 58.950 892.050 60.750 ;
        RECT 901.950 58.950 904.050 60.750 ;
        RECT 838.950 55.950 841.050 57.750 ;
        RECT 853.950 56.250 856.050 58.050 ;
        RECT 859.950 56.250 862.050 58.050 ;
        RECT 880.950 56.250 883.050 58.050 ;
        RECT 886.950 56.250 889.050 58.050 ;
        RECT 898.950 56.250 901.050 58.050 ;
        RECT 853.950 52.950 856.050 55.050 ;
        RECT 859.950 52.950 862.050 55.050 ;
        RECT 769.950 47.400 799.050 48.450 ;
        RECT 769.950 46.950 772.050 47.400 ;
        RECT 778.950 46.950 781.050 47.400 ;
        RECT 784.950 46.950 787.050 47.400 ;
        RECT 796.950 46.950 799.050 47.400 ;
        RECT 814.950 46.500 817.050 48.600 ;
        RECT 835.950 46.500 838.050 48.600 ;
        RECT 844.950 48.450 847.050 49.050 ;
        RECT 860.400 48.450 861.450 52.950 ;
        RECT 880.950 49.950 883.050 55.050 ;
        RECT 886.950 52.950 889.050 55.050 ;
        RECT 898.950 52.950 901.050 55.050 ;
        RECT 844.950 47.400 861.450 48.450 ;
        RECT 868.950 48.450 871.050 49.050 ;
        RECT 898.950 48.450 901.050 49.050 ;
        RECT 868.950 47.400 901.050 48.450 ;
        RECT 844.950 46.950 847.050 47.400 ;
        RECT 868.950 46.950 871.050 47.400 ;
        RECT 898.950 46.950 901.050 47.400 ;
        RECT 562.950 45.450 565.050 46.050 ;
        RECT 524.400 44.400 565.050 45.450 ;
        RECT 469.950 43.950 472.050 44.400 ;
        RECT 520.950 43.950 523.050 44.400 ;
        RECT 562.950 43.950 565.050 44.400 ;
        RECT 736.950 45.450 739.050 46.050 ;
        RECT 808.950 45.450 811.050 46.050 ;
        RECT 736.950 44.400 811.050 45.450 ;
        RECT 736.950 43.950 739.050 44.400 ;
        RECT 808.950 43.950 811.050 44.400 ;
        RECT 73.950 41.400 120.450 42.450 ;
        RECT 151.950 42.450 154.050 43.050 ;
        RECT 163.950 42.450 166.050 43.050 ;
        RECT 151.950 41.400 166.050 42.450 ;
        RECT 73.950 40.950 76.050 41.400 ;
        RECT 151.950 40.950 154.050 41.400 ;
        RECT 163.950 40.950 166.050 41.400 ;
        RECT 181.950 42.450 184.050 43.050 ;
        RECT 331.950 42.450 334.050 43.050 ;
        RECT 181.950 41.400 334.050 42.450 ;
        RECT 181.950 40.950 184.050 41.400 ;
        RECT 331.950 40.950 334.050 41.400 ;
        RECT 412.950 42.450 415.050 43.050 ;
        RECT 466.950 42.450 469.050 43.050 ;
        RECT 499.950 42.450 502.050 43.050 ;
        RECT 412.950 41.400 502.050 42.450 ;
        RECT 412.950 40.950 415.050 41.400 ;
        RECT 466.950 40.950 469.050 41.400 ;
        RECT 499.950 40.950 502.050 41.400 ;
        RECT 550.950 42.450 553.050 43.050 ;
        RECT 610.800 42.450 612.900 43.050 ;
        RECT 550.950 41.400 612.900 42.450 ;
        RECT 550.950 40.950 553.050 41.400 ;
        RECT 610.800 40.950 612.900 41.400 ;
        RECT 614.100 42.450 616.200 43.050 ;
        RECT 694.950 42.450 697.050 43.050 ;
        RECT 614.100 41.400 697.050 42.450 ;
        RECT 614.100 40.950 616.200 41.400 ;
        RECT 694.950 40.950 697.050 41.400 ;
        RECT 880.950 42.450 883.050 43.050 ;
        RECT 892.950 42.450 895.050 43.050 ;
        RECT 880.950 41.400 895.050 42.450 ;
        RECT 880.950 40.950 883.050 41.400 ;
        RECT 892.950 40.950 895.050 41.400 ;
        RECT 43.950 39.450 46.050 40.050 ;
        RECT 205.950 39.450 208.050 40.050 ;
        RECT 217.950 39.450 220.050 40.050 ;
        RECT 271.950 39.450 274.050 40.050 ;
        RECT 283.950 39.450 286.050 40.050 ;
        RECT 355.950 39.450 358.050 40.050 ;
        RECT 43.950 38.400 204.450 39.450 ;
        RECT 43.950 37.950 46.050 38.400 ;
        RECT 22.950 36.450 25.050 37.050 ;
        RECT 34.950 36.450 37.050 37.050 ;
        RECT 22.950 35.400 37.050 36.450 ;
        RECT 22.950 34.950 25.050 35.400 ;
        RECT 34.950 34.950 37.050 35.400 ;
        RECT 100.950 36.450 103.050 37.050 ;
        RECT 118.950 36.450 121.050 37.050 ;
        RECT 100.950 35.400 121.050 36.450 ;
        RECT 203.400 36.450 204.450 38.400 ;
        RECT 205.950 38.400 358.050 39.450 ;
        RECT 205.950 37.950 208.050 38.400 ;
        RECT 217.950 37.950 220.050 38.400 ;
        RECT 271.950 37.950 274.050 38.400 ;
        RECT 283.950 37.950 286.050 38.400 ;
        RECT 355.950 37.950 358.050 38.400 ;
        RECT 376.950 39.450 379.050 40.050 ;
        RECT 394.950 39.450 397.050 40.050 ;
        RECT 376.950 38.400 397.050 39.450 ;
        RECT 376.950 37.950 379.050 38.400 ;
        RECT 394.950 37.950 397.050 38.400 ;
        RECT 400.950 39.450 403.050 40.050 ;
        RECT 457.950 39.450 460.050 40.050 ;
        RECT 400.950 38.400 460.050 39.450 ;
        RECT 400.950 37.950 403.050 38.400 ;
        RECT 457.950 37.950 460.050 38.400 ;
        RECT 463.950 39.450 466.050 40.050 ;
        RECT 541.950 39.450 544.050 40.050 ;
        RECT 553.950 39.450 556.050 40.050 ;
        RECT 574.950 39.450 577.050 40.050 ;
        RECT 589.950 39.450 592.050 40.050 ;
        RECT 631.950 39.450 634.050 40.050 ;
        RECT 730.950 39.450 733.050 40.050 ;
        RECT 736.950 39.450 739.050 40.050 ;
        RECT 760.950 39.450 763.050 40.050 ;
        RECT 772.950 39.450 775.050 40.050 ;
        RECT 463.950 38.400 763.050 39.450 ;
        RECT 767.250 39.000 775.050 39.450 ;
        RECT 463.950 37.950 466.050 38.400 ;
        RECT 541.950 37.950 544.050 38.400 ;
        RECT 553.950 37.950 556.050 38.400 ;
        RECT 574.950 37.950 577.050 38.400 ;
        RECT 589.950 37.950 592.050 38.400 ;
        RECT 631.950 37.950 634.050 38.400 ;
        RECT 730.950 37.950 733.050 38.400 ;
        RECT 736.950 37.950 739.050 38.400 ;
        RECT 760.950 37.950 763.050 38.400 ;
        RECT 766.950 38.400 775.050 39.000 ;
        RECT 766.950 37.050 769.050 38.400 ;
        RECT 772.950 37.950 775.050 38.400 ;
        RECT 796.950 39.450 799.050 40.050 ;
        RECT 886.950 39.450 889.050 40.050 ;
        RECT 796.950 38.400 889.050 39.450 ;
        RECT 796.950 37.950 799.050 38.400 ;
        RECT 886.950 37.950 889.050 38.400 ;
        RECT 229.950 36.450 232.050 37.050 ;
        RECT 203.400 35.400 232.050 36.450 ;
        RECT 100.950 34.950 103.050 35.400 ;
        RECT 118.950 34.950 121.050 35.400 ;
        RECT 229.950 34.950 232.050 35.400 ;
        RECT 265.950 36.450 268.050 37.050 ;
        RECT 331.950 36.450 334.050 37.050 ;
        RECT 265.950 35.400 334.050 36.450 ;
        RECT 265.950 34.950 268.050 35.400 ;
        RECT 331.950 34.950 334.050 35.400 ;
        RECT 337.950 36.450 340.050 37.050 ;
        RECT 367.950 36.450 370.050 37.050 ;
        RECT 337.950 35.400 370.050 36.450 ;
        RECT 337.950 34.950 340.050 35.400 ;
        RECT 367.950 34.950 370.050 35.400 ;
        RECT 436.950 36.450 439.050 37.050 ;
        RECT 442.950 36.450 445.050 37.050 ;
        RECT 436.950 35.400 445.050 36.450 ;
        RECT 436.950 34.950 439.050 35.400 ;
        RECT 442.950 34.950 445.050 35.400 ;
        RECT 559.950 36.450 562.050 37.050 ;
        RECT 643.950 36.450 646.050 37.050 ;
        RECT 559.950 35.400 646.050 36.450 ;
        RECT 559.950 34.950 562.050 35.400 ;
        RECT 643.950 34.950 646.050 35.400 ;
        RECT 766.800 36.000 769.050 37.050 ;
        RECT 770.100 36.450 772.200 37.050 ;
        RECT 775.950 36.450 778.050 37.050 ;
        RECT 766.800 34.950 768.900 36.000 ;
        RECT 770.100 35.400 778.050 36.450 ;
        RECT 770.100 34.950 772.200 35.400 ;
        RECT 775.950 34.950 778.050 35.400 ;
        RECT 832.950 36.450 835.050 37.050 ;
        RECT 841.950 36.450 844.050 37.050 ;
        RECT 832.950 35.400 844.050 36.450 ;
        RECT 832.950 34.950 835.050 35.400 ;
        RECT 841.950 34.950 844.050 35.400 ;
        RECT 43.950 33.450 46.050 34.050 ;
        RECT 17.400 32.400 46.050 33.450 ;
        RECT 49.950 32.400 52.050 34.500 ;
        RECT 70.950 32.400 73.050 34.500 ;
        RECT 136.950 33.450 139.050 34.050 ;
        RECT 95.400 32.400 139.050 33.450 ;
        RECT 157.950 32.400 160.050 34.500 ;
        RECT 178.950 32.400 181.050 34.500 ;
        RECT 238.950 32.400 241.050 34.500 ;
        RECT 259.950 32.400 262.050 34.500 ;
        RECT 368.400 33.450 369.450 34.950 ;
        RECT 388.950 33.450 391.050 34.050 ;
        RECT 368.400 32.400 391.050 33.450 ;
        RECT 394.950 32.400 397.050 34.500 ;
        RECT 415.950 32.400 418.050 34.500 ;
        RECT 475.950 32.400 478.050 34.500 ;
        RECT 496.950 32.400 499.050 34.500 ;
        RECT 535.950 33.450 538.050 34.050 ;
        RECT 565.950 33.450 568.050 34.050 ;
        RECT 607.950 33.450 610.050 34.050 ;
        RECT 631.950 33.450 634.050 34.050 ;
        RECT 535.950 32.400 634.050 33.450 ;
        RECT 17.400 28.050 18.450 32.400 ;
        RECT 43.950 31.950 46.050 32.400 ;
        RECT 16.950 25.950 19.050 28.050 ;
        RECT 28.950 25.950 31.050 28.050 ;
        RECT 34.950 25.950 37.050 31.050 ;
        RECT 46.950 25.950 49.050 28.050 ;
        RECT 16.950 22.950 19.050 24.750 ;
        RECT 28.950 22.950 31.050 24.750 ;
        RECT 34.950 22.950 37.050 24.750 ;
        RECT 46.950 22.950 49.050 24.750 ;
        RECT 13.950 20.250 16.050 22.050 ;
        RECT 31.950 20.250 34.050 22.050 ;
        RECT 37.950 20.250 40.050 22.050 ;
        RECT 13.950 18.450 16.050 19.050 ;
        RECT 25.950 18.450 28.050 19.050 ;
        RECT 13.950 17.400 28.050 18.450 ;
        RECT 13.950 16.950 16.050 17.400 ;
        RECT 25.950 16.950 28.050 17.400 ;
        RECT 31.950 16.950 34.050 19.050 ;
        RECT 37.950 16.950 40.050 19.050 ;
        RECT 50.850 17.400 52.050 32.400 ;
        RECT 64.950 23.250 67.050 25.050 ;
        RECT 64.950 19.950 67.050 22.050 ;
        RECT 49.950 15.300 52.050 17.400 ;
        RECT 50.850 11.700 52.050 15.300 ;
        RECT 71.100 12.600 72.300 32.400 ;
        RECT 95.400 28.050 96.450 32.400 ;
        RECT 136.950 31.950 139.050 32.400 ;
        RECT 94.950 25.950 97.050 28.050 ;
        RECT 100.950 25.950 103.050 28.050 ;
        RECT 118.950 25.950 121.050 28.050 ;
        RECT 136.950 25.950 139.050 28.050 ;
        RECT 142.950 27.450 145.050 28.050 ;
        RECT 151.950 27.450 154.050 28.050 ;
        RECT 142.950 26.400 154.050 27.450 ;
        RECT 142.950 25.950 145.050 26.400 ;
        RECT 151.950 25.950 154.050 26.400 ;
        RECT 73.950 23.250 76.050 25.050 ;
        RECT 94.950 22.950 97.050 24.750 ;
        RECT 100.950 22.950 103.050 24.750 ;
        RECT 112.950 23.250 115.050 25.050 ;
        RECT 122.250 24.750 124.050 25.050 ;
        RECT 118.950 23.250 121.050 24.750 ;
        RECT 121.950 23.250 124.050 24.750 ;
        RECT 118.950 22.950 120.750 23.250 ;
        RECT 136.950 22.950 139.050 24.750 ;
        RECT 142.950 22.950 145.050 24.750 ;
        RECT 154.950 23.250 157.050 25.050 ;
        RECT 73.950 19.950 76.050 22.050 ;
        RECT 91.950 20.250 94.050 22.050 ;
        RECT 97.950 20.250 100.050 22.050 ;
        RECT 112.950 19.950 115.050 22.050 ;
        RECT 121.950 21.450 124.050 22.050 ;
        RECT 133.950 21.450 136.050 22.050 ;
        RECT 121.950 20.400 136.050 21.450 ;
        RECT 121.950 19.950 124.050 20.400 ;
        RECT 133.950 19.950 136.050 20.400 ;
        RECT 139.950 20.250 142.050 22.050 ;
        RECT 145.950 20.250 148.050 22.050 ;
        RECT 154.950 19.950 157.050 22.050 ;
        RECT 91.950 16.950 94.050 19.050 ;
        RECT 97.950 18.450 100.050 19.050 ;
        RECT 106.950 18.450 109.050 19.050 ;
        RECT 97.950 17.400 109.050 18.450 ;
        RECT 97.950 16.950 100.050 17.400 ;
        RECT 106.950 16.950 109.050 17.400 ;
        RECT 139.950 16.950 142.050 19.050 ;
        RECT 145.950 16.950 148.050 19.050 ;
        RECT 49.950 9.600 52.050 11.700 ;
        RECT 70.950 10.500 73.050 12.600 ;
        RECT 133.950 12.450 136.050 13.050 ;
        RECT 139.950 12.450 142.050 13.050 ;
        RECT 158.700 12.600 159.900 32.400 ;
        RECT 163.950 23.250 166.050 25.050 ;
        RECT 163.950 19.950 166.050 22.050 ;
        RECT 178.950 17.400 180.150 32.400 ;
        RECT 181.950 25.950 184.050 28.050 ;
        RECT 187.950 27.450 190.050 28.050 ;
        RECT 199.950 27.450 202.050 28.050 ;
        RECT 187.950 26.400 202.050 27.450 ;
        RECT 187.950 25.950 190.050 26.400 ;
        RECT 199.950 25.950 202.050 26.400 ;
        RECT 217.950 25.950 220.050 28.050 ;
        RECT 223.950 25.950 229.050 28.050 ;
        RECT 181.950 22.950 184.050 24.750 ;
        RECT 199.950 22.950 202.050 24.750 ;
        RECT 217.950 22.950 220.050 24.750 ;
        RECT 223.950 22.950 226.050 24.750 ;
        RECT 235.950 23.250 238.050 25.050 ;
        RECT 196.950 20.250 199.050 22.050 ;
        RECT 202.950 20.250 205.050 22.050 ;
        RECT 220.950 20.250 223.050 22.050 ;
        RECT 226.950 20.250 229.050 22.050 ;
        RECT 235.950 19.950 238.050 22.050 ;
        RECT 184.950 18.450 187.050 19.050 ;
        RECT 196.950 18.450 199.050 19.050 ;
        RECT 184.950 17.400 199.050 18.450 ;
        RECT 178.950 15.300 181.050 17.400 ;
        RECT 184.950 16.950 187.050 17.400 ;
        RECT 196.950 16.950 199.050 17.400 ;
        RECT 202.950 16.950 205.050 19.050 ;
        RECT 220.950 16.950 223.050 19.050 ;
        RECT 226.950 16.950 229.050 19.050 ;
        RECT 133.950 11.400 142.050 12.450 ;
        RECT 133.950 10.950 136.050 11.400 ;
        RECT 139.950 10.950 142.050 11.400 ;
        RECT 157.950 10.500 160.050 12.600 ;
        RECT 178.950 11.700 180.150 15.300 ;
        RECT 193.950 12.450 196.050 13.050 ;
        RECT 220.950 12.450 223.050 13.050 ;
        RECT 239.700 12.600 240.900 32.400 ;
        RECT 244.950 23.250 247.050 25.050 ;
        RECT 244.950 19.950 247.050 22.050 ;
        RECT 259.950 17.400 261.150 32.400 ;
        RECT 388.950 31.950 391.050 32.400 ;
        RECT 301.950 28.950 304.050 31.050 ;
        RECT 307.950 28.950 310.050 31.050 ;
        RECT 313.950 28.950 319.050 31.050 ;
        RECT 331.950 28.950 334.050 31.050 ;
        RECT 337.950 28.950 340.050 31.050 ;
        RECT 262.950 25.950 265.050 28.050 ;
        RECT 268.950 27.450 271.050 28.050 ;
        RECT 280.950 27.450 283.050 28.050 ;
        RECT 268.950 26.400 283.050 27.450 ;
        RECT 268.950 25.950 271.050 26.400 ;
        RECT 280.950 25.950 283.050 26.400 ;
        RECT 301.950 25.950 304.050 27.750 ;
        RECT 307.950 25.950 310.050 27.750 ;
        RECT 331.950 25.950 334.050 27.750 ;
        RECT 337.950 25.950 340.050 27.750 ;
        RECT 358.950 27.450 361.050 28.050 ;
        RECT 370.950 27.450 373.050 28.050 ;
        RECT 358.950 26.400 373.050 27.450 ;
        RECT 358.950 25.950 361.050 26.400 ;
        RECT 370.950 25.950 373.050 26.400 ;
        RECT 376.950 25.950 382.050 28.050 ;
        RECT 385.950 25.950 388.050 28.050 ;
        RECT 391.950 25.950 394.050 28.050 ;
        RECT 262.950 22.950 265.050 24.750 ;
        RECT 280.950 22.950 283.050 24.750 ;
        RECT 298.950 23.250 301.050 25.050 ;
        RECT 304.950 23.250 307.050 25.050 ;
        RECT 310.950 23.250 313.050 25.050 ;
        RECT 328.950 23.250 331.050 25.050 ;
        RECT 334.950 23.250 337.050 25.050 ;
        RECT 340.950 23.250 343.050 25.050 ;
        RECT 358.950 22.950 361.050 24.750 ;
        RECT 379.950 22.950 382.050 24.750 ;
        RECT 385.950 22.950 388.050 24.750 ;
        RECT 391.950 22.950 394.050 24.750 ;
        RECT 277.950 20.250 280.050 22.050 ;
        RECT 283.950 20.250 286.050 22.050 ;
        RECT 298.950 19.950 301.050 22.050 ;
        RECT 265.950 18.450 268.050 19.050 ;
        RECT 277.950 18.450 280.050 19.050 ;
        RECT 265.950 17.400 280.050 18.450 ;
        RECT 244.950 15.450 247.050 16.050 ;
        RECT 253.950 15.450 256.050 16.050 ;
        RECT 244.950 14.400 256.050 15.450 ;
        RECT 244.950 13.950 247.050 14.400 ;
        RECT 253.950 13.950 256.050 14.400 ;
        RECT 259.950 15.300 262.050 17.400 ;
        RECT 265.950 16.950 268.050 17.400 ;
        RECT 277.950 16.950 280.050 17.400 ;
        RECT 283.950 16.950 286.050 19.050 ;
        RECT 304.950 16.950 307.050 22.050 ;
        RECT 310.950 19.950 313.050 22.050 ;
        RECT 328.950 19.950 331.050 22.050 ;
        RECT 334.950 16.950 337.050 22.050 ;
        RECT 340.950 19.950 343.050 22.050 ;
        RECT 355.950 20.250 358.050 22.050 ;
        RECT 361.950 20.250 364.050 22.050 ;
        RECT 376.950 20.250 379.050 22.050 ;
        RECT 382.950 20.250 385.050 22.050 ;
        RECT 355.950 16.950 358.050 19.050 ;
        RECT 361.950 18.450 364.050 19.050 ;
        RECT 366.000 18.450 370.050 19.050 ;
        RECT 361.950 17.400 370.050 18.450 ;
        RECT 361.950 16.950 364.050 17.400 ;
        RECT 366.000 16.950 370.050 17.400 ;
        RECT 376.950 16.950 379.050 19.050 ;
        RECT 382.950 16.950 385.050 19.050 ;
        RECT 395.850 17.400 397.050 32.400 ;
        RECT 400.950 30.450 403.050 31.050 ;
        RECT 409.950 30.450 412.050 31.050 ;
        RECT 400.950 29.400 412.050 30.450 ;
        RECT 400.950 28.950 403.050 29.400 ;
        RECT 409.950 28.950 412.050 29.400 ;
        RECT 409.950 23.250 412.050 25.050 ;
        RECT 409.950 19.950 412.050 22.050 ;
        RECT 178.950 9.600 181.050 11.700 ;
        RECT 193.950 11.400 223.050 12.450 ;
        RECT 193.950 10.950 196.050 11.400 ;
        RECT 220.950 10.950 223.050 11.400 ;
        RECT 238.950 10.500 241.050 12.600 ;
        RECT 259.950 11.700 261.150 15.300 ;
        RECT 278.400 12.450 279.450 16.950 ;
        RECT 298.950 15.450 301.050 16.050 ;
        RECT 340.950 15.450 343.050 16.050 ;
        RECT 298.950 14.400 343.050 15.450 ;
        RECT 394.950 15.300 397.050 17.400 ;
        RECT 298.950 13.950 301.050 14.400 ;
        RECT 340.950 13.950 343.050 14.400 ;
        RECT 316.950 12.450 319.050 13.050 ;
        RECT 259.950 9.600 262.050 11.700 ;
        RECT 278.400 11.400 319.050 12.450 ;
        RECT 316.950 10.950 319.050 11.400 ;
        RECT 361.950 12.450 364.050 13.050 ;
        RECT 382.950 12.450 385.050 13.050 ;
        RECT 361.950 11.400 385.050 12.450 ;
        RECT 395.850 11.700 397.050 15.300 ;
        RECT 416.100 12.600 417.300 32.400 ;
        RECT 457.950 28.950 460.050 31.050 ;
        RECT 463.950 28.950 466.050 31.050 ;
        RECT 457.950 25.950 460.050 27.750 ;
        RECT 463.950 25.950 466.050 27.750 ;
        RECT 418.950 23.250 421.050 25.050 ;
        RECT 433.950 22.950 436.050 24.750 ;
        RECT 454.950 23.250 457.050 25.050 ;
        RECT 460.950 23.250 463.050 25.050 ;
        RECT 466.950 23.250 469.050 25.050 ;
        RECT 472.950 23.250 475.050 25.050 ;
        RECT 418.950 19.950 421.050 22.050 ;
        RECT 436.950 20.250 439.050 22.050 ;
        RECT 454.950 19.950 457.050 22.050 ;
        RECT 436.950 18.450 439.050 19.050 ;
        RECT 441.000 18.450 445.050 19.050 ;
        RECT 436.950 17.400 445.050 18.450 ;
        RECT 436.950 16.950 439.050 17.400 ;
        RECT 441.000 16.950 445.050 17.400 ;
        RECT 460.950 16.950 463.050 22.050 ;
        RECT 466.950 19.950 469.050 22.050 ;
        RECT 472.950 19.950 475.050 22.050 ;
        RECT 361.950 10.950 364.050 11.400 ;
        RECT 382.950 10.950 385.050 11.400 ;
        RECT 310.950 9.450 313.050 10.050 ;
        RECT 325.950 9.450 328.050 10.050 ;
        RECT 394.950 9.600 397.050 11.700 ;
        RECT 415.950 10.500 418.050 12.600 ;
        RECT 421.950 12.450 424.050 13.050 ;
        RECT 454.950 12.450 457.050 13.050 ;
        RECT 476.700 12.600 477.900 32.400 ;
        RECT 481.950 30.450 484.050 31.050 ;
        RECT 487.950 30.450 490.050 31.050 ;
        RECT 481.950 29.400 490.050 30.450 ;
        RECT 481.950 28.950 484.050 29.400 ;
        RECT 487.950 28.950 490.050 29.400 ;
        RECT 481.950 23.250 484.050 25.050 ;
        RECT 481.950 19.950 484.050 22.050 ;
        RECT 496.950 17.400 498.150 32.400 ;
        RECT 535.950 31.950 538.050 32.400 ;
        RECT 565.950 31.950 568.050 32.400 ;
        RECT 607.950 31.950 610.050 32.400 ;
        RECT 631.950 31.950 634.050 32.400 ;
        RECT 637.950 33.450 640.050 34.050 ;
        RECT 718.950 33.450 721.050 34.050 ;
        RECT 730.950 33.450 733.050 34.050 ;
        RECT 637.950 32.400 687.450 33.450 ;
        RECT 637.950 31.950 640.050 32.400 ;
        RECT 499.950 27.450 502.050 28.050 ;
        RECT 508.950 27.450 511.050 28.050 ;
        RECT 499.950 26.400 511.050 27.450 ;
        RECT 499.950 25.950 502.050 26.400 ;
        RECT 508.950 25.950 511.050 26.400 ;
        RECT 514.950 25.950 517.050 28.050 ;
        RECT 538.950 27.450 541.050 28.050 ;
        RECT 553.950 27.450 556.050 28.050 ;
        RECT 538.950 26.400 556.050 27.450 ;
        RECT 538.950 25.950 541.050 26.400 ;
        RECT 553.950 25.950 556.050 26.400 ;
        RECT 559.950 25.950 562.050 28.050 ;
        RECT 565.950 25.950 568.050 28.050 ;
        RECT 571.950 27.450 574.050 28.050 ;
        RECT 583.950 27.450 586.050 28.050 ;
        RECT 571.950 26.400 586.050 27.450 ;
        RECT 571.950 25.950 574.050 26.400 ;
        RECT 583.950 25.950 586.050 26.400 ;
        RECT 589.950 25.950 592.050 28.050 ;
        RECT 601.950 25.950 604.050 28.050 ;
        RECT 625.950 25.950 628.050 28.050 ;
        RECT 631.950 25.950 634.050 28.050 ;
        RECT 643.950 25.950 646.050 31.050 ;
        RECT 686.400 28.050 687.450 32.400 ;
        RECT 718.950 32.400 733.050 33.450 ;
        RECT 718.950 31.950 721.050 32.400 ;
        RECT 730.950 31.950 733.050 32.400 ;
        RECT 772.950 33.450 775.050 34.050 ;
        RECT 784.950 33.450 787.050 34.050 ;
        RECT 772.950 32.400 787.050 33.450 ;
        RECT 790.950 32.400 793.050 34.500 ;
        RECT 811.950 32.400 814.050 34.500 ;
        RECT 826.950 32.400 829.050 34.500 ;
        RECT 847.950 32.400 850.050 34.500 ;
        RECT 772.950 31.950 775.050 32.400 ;
        RECT 784.950 31.950 787.050 32.400 ;
        RECT 658.950 27.450 663.000 28.050 ;
        RECT 664.950 27.450 667.050 28.050 ;
        RECT 658.950 26.400 667.050 27.450 ;
        RECT 658.950 25.950 663.000 26.400 ;
        RECT 664.950 25.950 667.050 26.400 ;
        RECT 685.950 25.950 688.050 28.050 ;
        RECT 694.950 27.450 697.050 28.050 ;
        RECT 706.950 27.450 709.050 28.050 ;
        RECT 694.950 26.400 709.050 27.450 ;
        RECT 694.950 25.950 697.050 26.400 ;
        RECT 706.950 25.950 709.050 26.400 ;
        RECT 733.950 27.450 736.050 28.050 ;
        RECT 742.950 27.450 745.050 28.050 ;
        RECT 754.950 27.450 757.050 28.050 ;
        RECT 733.950 26.400 741.450 27.450 ;
        RECT 733.950 25.950 736.050 26.400 ;
        RECT 499.950 22.950 502.050 24.750 ;
        RECT 514.950 22.950 517.050 24.750 ;
        RECT 538.950 22.950 541.050 24.750 ;
        RECT 559.950 22.950 562.050 24.750 ;
        RECT 565.950 22.950 568.050 24.750 ;
        RECT 583.950 22.950 586.050 24.750 ;
        RECT 589.950 22.950 592.050 24.750 ;
        RECT 601.950 22.950 604.050 24.750 ;
        RECT 625.950 22.950 628.050 24.750 ;
        RECT 631.950 22.950 634.050 24.750 ;
        RECT 643.950 22.950 646.050 24.750 ;
        RECT 649.950 23.250 652.050 25.050 ;
        RECT 664.950 22.950 667.050 24.750 ;
        RECT 670.950 23.250 673.050 25.050 ;
        RECT 685.950 22.950 688.050 24.750 ;
        RECT 691.950 23.250 694.050 25.050 ;
        RECT 706.950 22.950 709.050 24.750 ;
        RECT 712.950 23.250 715.050 25.050 ;
        RECT 733.950 22.950 736.050 24.750 ;
        RECT 740.400 24.450 741.450 26.400 ;
        RECT 742.950 26.400 757.050 27.450 ;
        RECT 742.950 25.950 745.050 26.400 ;
        RECT 754.950 25.950 757.050 26.400 ;
        RECT 760.950 25.950 763.050 28.050 ;
        RECT 769.950 27.450 774.000 28.050 ;
        RECT 775.950 27.450 778.050 28.050 ;
        RECT 769.950 26.400 778.050 27.450 ;
        RECT 769.950 25.950 774.000 26.400 ;
        RECT 775.950 25.950 778.050 26.400 ;
        RECT 787.950 25.950 790.050 28.050 ;
        RECT 748.950 24.450 751.050 25.050 ;
        RECT 740.400 23.400 751.050 24.450 ;
        RECT 748.950 22.950 751.050 23.400 ;
        RECT 754.950 22.950 757.050 24.750 ;
        RECT 760.950 22.950 763.050 24.750 ;
        RECT 775.950 22.950 778.050 24.750 ;
        RECT 787.950 22.950 790.050 24.750 ;
        RECT 517.950 20.250 520.050 22.050 ;
        RECT 535.950 20.250 538.050 22.050 ;
        RECT 541.950 20.250 544.050 22.050 ;
        RECT 556.950 20.250 559.050 22.050 ;
        RECT 562.950 20.250 565.050 22.050 ;
        RECT 580.950 20.250 583.050 22.050 ;
        RECT 586.950 20.250 589.050 22.050 ;
        RECT 604.950 20.250 607.050 22.050 ;
        RECT 622.950 20.250 625.050 22.050 ;
        RECT 628.950 20.250 631.050 22.050 ;
        RECT 730.950 20.250 733.050 22.050 ;
        RECT 736.950 20.250 739.050 22.050 ;
        RECT 751.950 20.250 754.050 22.050 ;
        RECT 757.950 20.250 760.050 22.050 ;
        RECT 772.950 20.250 775.050 22.050 ;
        RECT 778.950 20.250 781.050 22.050 ;
        RECT 496.950 15.300 499.050 17.400 ;
        RECT 517.950 16.950 520.050 19.050 ;
        RECT 535.950 16.950 538.050 19.050 ;
        RECT 541.950 16.950 544.050 19.050 ;
        RECT 556.950 16.950 559.050 19.050 ;
        RECT 562.950 16.950 565.050 19.050 ;
        RECT 580.950 16.950 583.050 19.050 ;
        RECT 586.950 16.950 589.050 19.050 ;
        RECT 604.950 16.950 607.050 19.050 ;
        RECT 622.950 16.950 625.050 19.050 ;
        RECT 628.950 16.950 631.050 19.050 ;
        RECT 730.950 16.950 733.050 19.050 ;
        RECT 736.950 16.950 739.050 19.050 ;
        RECT 751.950 16.950 754.050 19.050 ;
        RECT 757.950 16.950 760.050 19.050 ;
        RECT 772.950 16.950 775.050 19.050 ;
        RECT 778.950 16.950 781.050 19.050 ;
        RECT 791.850 17.400 793.050 32.400 ;
        RECT 796.950 30.450 799.050 31.050 ;
        RECT 805.950 30.450 808.050 31.050 ;
        RECT 796.950 29.400 808.050 30.450 ;
        RECT 796.950 28.950 799.050 29.400 ;
        RECT 805.950 28.950 808.050 29.400 ;
        RECT 805.950 23.250 808.050 25.050 ;
        RECT 805.950 19.950 808.050 22.050 ;
        RECT 565.950 15.450 568.050 16.050 ;
        RECT 574.950 15.450 577.050 16.050 ;
        RECT 421.950 11.400 457.050 12.450 ;
        RECT 421.950 10.950 424.050 11.400 ;
        RECT 454.950 10.950 457.050 11.400 ;
        RECT 475.950 10.500 478.050 12.600 ;
        RECT 496.950 11.700 498.150 15.300 ;
        RECT 565.950 14.400 577.050 15.450 ;
        RECT 790.950 15.300 793.050 17.400 ;
        RECT 565.950 13.950 568.050 14.400 ;
        RECT 574.950 13.950 577.050 14.400 ;
        RECT 502.950 12.450 505.050 13.050 ;
        RECT 622.950 12.450 625.050 13.050 ;
        RECT 496.950 9.600 499.050 11.700 ;
        RECT 502.950 11.400 625.050 12.450 ;
        RECT 502.950 10.950 505.050 11.400 ;
        RECT 622.950 10.950 625.050 11.400 ;
        RECT 628.950 12.450 631.050 13.050 ;
        RECT 742.950 12.450 745.050 13.050 ;
        RECT 628.950 11.400 745.050 12.450 ;
        RECT 628.950 10.950 631.050 11.400 ;
        RECT 742.950 10.950 745.050 11.400 ;
        RECT 757.950 12.450 760.050 13.050 ;
        RECT 784.950 12.450 787.050 13.050 ;
        RECT 757.950 11.400 787.050 12.450 ;
        RECT 791.850 11.700 793.050 15.300 ;
        RECT 812.100 12.600 813.300 32.400 ;
        RECT 817.950 27.450 822.000 28.050 ;
        RECT 823.950 27.450 826.050 28.050 ;
        RECT 817.950 26.400 826.050 27.450 ;
        RECT 817.950 25.950 822.000 26.400 ;
        RECT 823.950 25.950 826.050 26.400 ;
        RECT 814.950 23.250 817.050 25.050 ;
        RECT 823.950 22.950 826.050 24.750 ;
        RECT 814.950 19.950 817.050 22.050 ;
        RECT 827.850 17.400 829.050 32.400 ;
        RECT 832.950 30.450 835.050 31.050 ;
        RECT 841.950 30.450 844.050 31.050 ;
        RECT 832.950 29.400 844.050 30.450 ;
        RECT 832.950 28.950 835.050 29.400 ;
        RECT 841.950 28.950 844.050 29.400 ;
        RECT 841.950 23.250 844.050 25.050 ;
        RECT 841.950 19.950 844.050 22.050 ;
        RECT 826.950 15.300 829.050 17.400 ;
        RECT 757.950 10.950 760.050 11.400 ;
        RECT 784.950 10.950 787.050 11.400 ;
        RECT 310.950 8.400 328.050 9.450 ;
        RECT 310.950 7.950 313.050 8.400 ;
        RECT 325.950 7.950 328.050 8.400 ;
        RECT 511.950 9.450 514.050 10.050 ;
        RECT 556.950 9.450 559.050 10.050 ;
        RECT 511.950 8.400 559.050 9.450 ;
        RECT 511.950 7.950 514.050 8.400 ;
        RECT 556.950 7.950 559.050 8.400 ;
        RECT 586.950 9.450 589.050 10.050 ;
        RECT 772.950 9.450 775.050 10.050 ;
        RECT 790.950 9.600 793.050 11.700 ;
        RECT 811.950 10.500 814.050 12.600 ;
        RECT 827.850 11.700 829.050 15.300 ;
        RECT 848.100 12.600 849.300 32.400 ;
        RECT 886.950 28.950 889.050 31.050 ;
        RECT 892.950 28.950 895.050 31.050 ;
        RECT 853.950 27.450 856.050 28.050 ;
        RECT 865.950 27.450 868.050 28.050 ;
        RECT 853.950 26.400 868.050 27.450 ;
        RECT 853.950 25.950 856.050 26.400 ;
        RECT 865.950 25.950 868.050 26.400 ;
        RECT 886.950 25.950 889.050 27.750 ;
        RECT 892.950 25.950 895.050 27.750 ;
        RECT 850.950 23.250 853.050 25.050 ;
        RECT 865.950 22.950 868.050 24.750 ;
        RECT 883.950 23.250 886.050 25.050 ;
        RECT 889.950 23.250 892.050 25.050 ;
        RECT 895.950 23.250 898.050 25.050 ;
        RECT 850.950 19.950 853.050 22.050 ;
        RECT 868.950 20.250 871.050 22.050 ;
        RECT 883.950 19.950 886.050 22.050 ;
        RECT 889.950 19.950 892.050 22.050 ;
        RECT 895.950 19.950 898.050 22.050 ;
        RECT 868.950 18.450 871.050 19.050 ;
        RECT 877.950 18.450 880.050 19.050 ;
        RECT 868.950 17.400 880.050 18.450 ;
        RECT 868.950 16.950 871.050 17.400 ;
        RECT 877.950 16.950 880.050 17.400 ;
        RECT 850.950 15.450 853.050 16.050 ;
        RECT 862.950 15.450 865.050 16.050 ;
        RECT 850.950 14.400 865.050 15.450 ;
        RECT 850.950 13.950 853.050 14.400 ;
        RECT 862.950 13.950 865.050 14.400 ;
        RECT 874.950 15.450 877.050 16.050 ;
        RECT 890.400 15.450 891.450 19.950 ;
        RECT 874.950 14.400 891.450 15.450 ;
        RECT 895.950 15.450 898.050 16.050 ;
        RECT 904.950 15.450 907.050 16.050 ;
        RECT 895.950 14.400 907.050 15.450 ;
        RECT 874.950 13.950 877.050 14.400 ;
        RECT 895.950 13.950 898.050 14.400 ;
        RECT 904.950 13.950 907.050 14.400 ;
        RECT 826.950 9.600 829.050 11.700 ;
        RECT 847.950 10.500 850.050 12.600 ;
        RECT 586.950 8.400 775.050 9.450 ;
        RECT 586.950 7.950 589.050 8.400 ;
        RECT 772.950 7.950 775.050 8.400 ;
        RECT 22.950 6.450 25.050 7.050 ;
        RECT 37.950 6.450 40.050 7.050 ;
        RECT 49.950 6.450 52.050 7.050 ;
        RECT 22.950 5.400 30.450 6.450 ;
        RECT 22.950 4.950 25.050 5.400 ;
        RECT 29.400 3.450 30.450 5.400 ;
        RECT 37.950 5.400 52.050 6.450 ;
        RECT 37.950 4.950 40.050 5.400 ;
        RECT 49.950 4.950 52.050 5.400 ;
        RECT 145.950 6.450 148.050 7.050 ;
        RECT 187.950 6.450 190.050 7.050 ;
        RECT 145.950 5.400 190.050 6.450 ;
        RECT 145.950 4.950 148.050 5.400 ;
        RECT 187.950 4.950 190.050 5.400 ;
        RECT 226.950 6.450 229.050 7.050 ;
        RECT 268.950 6.450 271.050 7.050 ;
        RECT 226.950 5.400 271.050 6.450 ;
        RECT 226.950 4.950 229.050 5.400 ;
        RECT 268.950 4.950 271.050 5.400 ;
        RECT 334.950 6.450 337.050 7.050 ;
        RECT 493.950 6.450 496.050 7.050 ;
        RECT 334.950 5.400 496.050 6.450 ;
        RECT 334.950 4.950 337.050 5.400 ;
        RECT 493.950 4.950 496.050 5.400 ;
        RECT 520.950 6.450 523.050 7.050 ;
        RECT 535.950 6.450 538.050 7.050 ;
        RECT 520.950 5.400 538.050 6.450 ;
        RECT 520.950 4.950 523.050 5.400 ;
        RECT 535.950 4.950 538.050 5.400 ;
        RECT 766.950 6.450 769.050 7.050 ;
        RECT 805.950 6.450 808.050 7.050 ;
        RECT 766.950 5.400 808.050 6.450 ;
        RECT 766.950 4.950 769.050 5.400 ;
        RECT 805.950 4.950 808.050 5.400 ;
        RECT 64.950 3.450 67.050 4.050 ;
        RECT 29.400 2.400 67.050 3.450 ;
        RECT 64.950 1.950 67.050 2.400 ;
        RECT 304.950 3.450 307.050 4.050 ;
        RECT 511.950 3.450 514.050 4.050 ;
        RECT 304.950 2.400 514.050 3.450 ;
        RECT 304.950 1.950 307.050 2.400 ;
        RECT 511.950 1.950 514.050 2.400 ;
      LAYER metal3 ;
        RECT 550.950 898.950 553.050 901.050 ;
        RECT 619.950 898.950 622.050 901.050 ;
        RECT 691.950 898.950 694.050 901.050 ;
        RECT 775.950 898.950 778.050 901.050 ;
        RECT 787.950 898.950 790.050 901.050 ;
        RECT 826.950 898.950 829.050 901.050 ;
        RECT 19.950 895.950 22.050 898.050 ;
        RECT 31.950 895.950 34.050 898.050 ;
        RECT 124.950 895.950 127.050 898.050 ;
        RECT 133.950 895.950 136.050 898.050 ;
        RECT 169.950 895.950 172.050 898.050 ;
        RECT 193.950 895.950 196.050 898.050 ;
        RECT 343.950 895.950 346.050 898.050 ;
        RECT 397.950 895.950 400.050 898.050 ;
        RECT 412.950 895.950 415.050 898.050 ;
        RECT 433.950 895.950 436.050 898.050 ;
        RECT 439.950 895.950 442.050 898.050 ;
        RECT 460.950 895.950 463.050 898.050 ;
        RECT 481.950 895.950 484.050 898.050 ;
        RECT 496.950 895.950 499.050 898.050 ;
        RECT 523.950 895.950 526.050 898.050 ;
        RECT 20.400 886.050 21.600 895.950 ;
        RECT 13.950 883.950 16.050 886.050 ;
        RECT 19.950 883.950 22.050 886.050 ;
        RECT 25.950 883.950 28.050 886.050 ;
        RECT 14.400 865.050 15.600 883.950 ;
        RECT 26.400 877.050 27.600 883.950 ;
        RECT 16.950 874.950 19.050 877.050 ;
        RECT 22.950 875.400 27.600 877.050 ;
        RECT 32.400 877.050 33.600 895.950 ;
        RECT 64.950 892.950 67.050 895.050 ;
        RECT 37.950 885.600 40.050 886.050 ;
        RECT 50.100 885.600 52.200 886.050 ;
        RECT 37.950 884.400 52.200 885.600 ;
        RECT 37.950 883.950 40.050 884.400 ;
        RECT 50.100 883.950 52.200 884.400 ;
        RECT 65.400 877.050 66.600 892.950 ;
        RECT 67.950 889.950 70.050 892.050 ;
        RECT 91.950 889.950 94.050 892.050 ;
        RECT 68.400 886.050 69.600 889.950 ;
        RECT 92.400 886.050 93.600 889.950 ;
        RECT 116.400 887.400 123.600 888.600 ;
        RECT 67.950 883.950 70.050 886.050 ;
        RECT 91.950 883.950 94.050 886.050 ;
        RECT 116.400 885.600 117.600 887.400 ;
        RECT 107.400 885.000 117.600 885.600 ;
        RECT 106.950 884.400 117.600 885.000 ;
        RECT 106.950 880.950 109.050 884.400 ;
        RECT 118.950 883.950 121.050 886.050 ;
        RECT 83.400 879.000 102.600 879.600 ;
        RECT 82.950 878.400 103.050 879.000 ;
        RECT 32.400 875.400 37.050 877.050 ;
        RECT 22.950 874.950 27.000 875.400 ;
        RECT 33.000 874.950 37.050 875.400 ;
        RECT 40.950 874.950 43.050 877.050 ;
        RECT 64.950 874.950 67.050 877.050 ;
        RECT 70.950 876.600 73.050 877.050 ;
        RECT 76.950 876.600 79.050 877.050 ;
        RECT 70.950 875.400 79.050 876.600 ;
        RECT 70.950 874.950 73.050 875.400 ;
        RECT 76.950 874.950 79.050 875.400 ;
        RECT 82.950 874.950 85.050 878.400 ;
        RECT 88.950 874.950 91.050 877.050 ;
        RECT 94.950 874.950 97.050 877.050 ;
        RECT 100.950 874.950 103.050 878.400 ;
        RECT 109.950 874.950 112.050 877.050 ;
        RECT 115.950 874.950 118.050 877.050 ;
        RECT 13.950 862.950 16.050 865.050 ;
        RECT 17.400 862.050 18.600 874.950 ;
        RECT 34.950 862.950 37.050 865.050 ;
        RECT 16.950 859.950 19.050 862.050 ;
        RECT 35.400 850.050 36.600 862.950 ;
        RECT 41.400 862.050 42.600 874.950 ;
        RECT 89.400 871.050 90.600 874.950 ;
        RECT 95.400 871.050 96.600 874.950 ;
        RECT 110.400 871.050 111.600 874.950 ;
        RECT 88.950 868.950 91.050 871.050 ;
        RECT 94.950 868.950 97.050 871.050 ;
        RECT 109.950 868.950 112.050 871.050 ;
        RECT 116.400 868.050 117.600 874.950 ;
        RECT 115.950 865.950 118.050 868.050 ;
        RECT 119.400 865.050 120.600 883.950 ;
        RECT 122.400 877.050 123.600 887.400 ;
        RECT 125.400 886.050 126.600 895.950 ;
        RECT 124.950 883.950 127.050 886.050 ;
        RECT 134.400 883.050 135.600 895.950 ;
        RECT 142.950 883.950 145.050 886.050 ;
        RECT 154.950 883.950 157.050 886.050 ;
        RECT 130.950 881.400 135.600 883.050 ;
        RECT 130.950 880.950 135.000 881.400 ;
        RECT 128.400 878.400 141.600 879.600 ;
        RECT 121.950 874.950 124.050 877.050 ;
        RECT 128.400 874.050 129.600 878.400 ;
        RECT 133.950 874.950 136.050 877.050 ;
        RECT 127.950 871.950 130.050 874.050 ;
        RECT 134.400 871.050 135.600 874.950 ;
        RECT 140.400 871.050 141.600 878.400 ;
        RECT 133.950 868.950 136.050 871.050 ;
        RECT 139.950 868.950 142.050 871.050 ;
        RECT 143.400 865.050 144.600 883.950 ;
        RECT 145.950 874.950 148.050 877.050 ;
        RECT 146.400 868.050 147.600 874.950 ;
        RECT 155.400 871.050 156.600 883.950 ;
        RECT 170.400 877.050 171.600 895.950 ;
        RECT 184.950 889.950 187.050 892.050 ;
        RECT 172.950 883.950 175.050 886.050 ;
        RECT 169.950 874.950 172.050 877.050 ;
        RECT 154.950 868.950 157.050 871.050 ;
        RECT 145.950 865.950 148.050 868.050 ;
        RECT 173.400 865.050 174.600 883.950 ;
        RECT 185.400 877.050 186.600 889.950 ;
        RECT 194.400 886.050 195.600 895.950 ;
        RECT 250.950 892.950 253.050 895.050 ;
        RECT 241.950 889.950 244.050 892.050 ;
        RECT 242.400 886.050 243.600 889.950 ;
        RECT 251.400 886.050 252.600 892.950 ;
        RECT 280.950 889.950 283.050 892.050 ;
        RECT 328.950 889.950 331.050 892.050 ;
        RECT 337.950 889.950 340.050 892.050 ;
        RECT 193.950 883.950 196.050 886.050 ;
        RECT 202.950 883.950 205.050 886.050 ;
        RECT 229.950 883.950 232.050 886.050 ;
        RECT 235.950 883.950 238.050 886.050 ;
        RECT 241.950 883.950 244.050 886.050 ;
        RECT 250.950 883.950 253.050 886.050 ;
        RECT 184.950 876.600 187.050 877.050 ;
        RECT 190.950 876.600 193.050 877.050 ;
        RECT 184.950 875.400 193.050 876.600 ;
        RECT 184.950 874.950 187.050 875.400 ;
        RECT 190.950 874.950 193.050 875.400 ;
        RECT 196.950 874.950 199.050 877.050 ;
        RECT 197.400 868.050 198.600 874.950 ;
        RECT 196.950 865.950 199.050 868.050 ;
        RECT 43.950 862.950 46.050 865.050 ;
        RECT 76.950 862.950 79.050 865.050 ;
        RECT 83.100 862.950 85.200 865.050 ;
        RECT 118.950 862.950 121.050 865.050 ;
        RECT 142.950 862.950 145.050 865.050 ;
        RECT 172.950 862.950 175.050 865.050 ;
        RECT 40.950 859.950 43.050 862.050 ;
        RECT 16.950 847.950 19.050 850.050 ;
        RECT 34.950 847.950 37.050 850.050 ;
        RECT 17.400 844.050 18.600 847.950 ;
        RECT 35.400 844.050 36.600 847.950 ;
        RECT 44.400 844.050 45.600 862.950 ;
        RECT 64.950 847.950 67.050 850.050 ;
        RECT 65.400 844.050 66.600 847.950 ;
        RECT 16.950 841.950 19.050 844.050 ;
        RECT 22.950 843.600 27.000 844.050 ;
        RECT 22.950 841.950 27.600 843.600 ;
        RECT 34.950 841.950 37.050 844.050 ;
        RECT 40.950 841.950 45.600 844.050 ;
        RECT 64.950 841.950 67.050 844.050 ;
        RECT 13.950 829.950 16.050 832.050 ;
        RECT 4.950 820.950 7.050 823.050 ;
        RECT 1.950 736.950 4.050 739.050 ;
        RECT 2.400 628.050 3.600 736.950 ;
        RECT 1.950 625.950 4.050 628.050 ;
        RECT 5.400 622.050 6.600 820.950 ;
        RECT 14.400 817.050 15.600 829.950 ;
        RECT 13.950 814.950 16.050 817.050 ;
        RECT 13.950 805.950 16.050 808.050 ;
        RECT 14.400 742.050 15.600 805.950 ;
        RECT 17.400 804.600 18.600 841.950 ;
        RECT 19.950 832.950 22.050 835.050 ;
        RECT 20.400 814.050 21.600 832.950 ;
        RECT 26.400 829.050 27.600 841.950 ;
        RECT 37.950 832.950 40.050 835.050 ;
        RECT 38.400 829.050 39.600 832.950 ;
        RECT 25.950 826.950 28.050 829.050 ;
        RECT 37.950 826.950 40.050 829.050 ;
        RECT 19.950 811.950 22.050 814.050 ;
        RECT 20.400 808.050 21.600 811.950 ;
        RECT 19.950 805.950 22.050 808.050 ;
        RECT 17.400 803.400 21.600 804.600 ;
        RECT 20.400 799.050 21.600 803.400 ;
        RECT 16.950 796.950 19.050 799.050 ;
        RECT 20.400 797.400 25.050 799.050 ;
        RECT 21.000 796.950 25.050 797.400 ;
        RECT 17.400 793.050 18.600 796.950 ;
        RECT 16.950 790.950 19.050 793.050 ;
        RECT 22.950 792.600 25.050 793.050 ;
        RECT 26.400 792.600 27.600 826.950 ;
        RECT 44.400 810.600 45.600 841.950 ;
        RECT 70.950 840.600 73.050 844.050 ;
        RECT 70.950 840.000 75.600 840.600 ;
        RECT 71.400 839.400 75.600 840.000 ;
        RECT 46.950 832.950 49.050 835.050 ;
        RECT 67.950 834.600 72.000 835.050 ;
        RECT 67.950 834.000 72.600 834.600 ;
        RECT 67.950 832.950 73.050 834.000 ;
        RECT 47.400 823.050 48.600 832.950 ;
        RECT 61.950 829.950 64.050 832.050 ;
        RECT 70.950 829.950 73.050 832.950 ;
        RECT 46.950 820.950 49.050 823.050 ;
        RECT 46.950 814.950 49.050 817.050 ;
        RECT 41.400 809.400 45.600 810.600 ;
        RECT 34.950 805.950 37.050 808.050 ;
        RECT 22.950 791.400 27.600 792.600 ;
        RECT 22.950 790.950 25.050 791.400 ;
        RECT 16.950 775.950 19.050 778.050 ;
        RECT 17.400 757.050 18.600 775.950 ;
        RECT 23.400 766.050 24.600 790.950 ;
        RECT 28.950 784.950 31.050 787.050 ;
        RECT 29.400 766.050 30.600 784.950 ;
        RECT 35.400 766.050 36.600 805.950 ;
        RECT 41.400 801.600 42.600 809.400 ;
        RECT 47.400 808.050 48.600 814.950 ;
        RECT 62.400 814.050 63.600 829.950 ;
        RECT 74.400 826.050 75.600 839.400 ;
        RECT 77.400 832.050 78.600 862.950 ;
        RECT 83.400 850.050 84.600 862.950 ;
        RECT 103.950 859.950 106.050 862.050 ;
        RECT 82.950 847.950 85.050 850.050 ;
        RECT 83.400 844.050 84.600 847.950 ;
        RECT 82.950 841.950 85.050 844.050 ;
        RECT 88.950 843.600 91.050 844.050 ;
        RECT 94.950 843.600 97.050 844.050 ;
        RECT 88.950 842.400 97.050 843.600 ;
        RECT 88.950 841.950 91.050 842.400 ;
        RECT 94.950 841.950 97.050 842.400 ;
        RECT 104.400 835.050 105.600 859.950 ;
        RECT 136.950 853.950 139.050 856.050 ;
        RECT 151.950 853.950 154.050 856.050 ;
        RECT 184.950 853.950 187.050 856.050 ;
        RECT 112.950 847.950 115.050 850.050 ;
        RECT 113.400 844.050 114.600 847.950 ;
        RECT 112.950 841.950 115.050 844.050 ;
        RECT 118.950 841.950 121.050 844.050 ;
        RECT 85.950 834.600 88.050 835.050 ;
        RECT 80.400 833.400 88.050 834.600 ;
        RECT 76.950 831.600 79.050 832.050 ;
        RECT 80.400 831.600 81.600 833.400 ;
        RECT 85.950 832.950 88.050 833.400 ;
        RECT 97.950 832.950 100.050 835.050 ;
        RECT 103.950 832.950 106.050 835.050 ;
        RECT 115.950 832.950 118.050 835.050 ;
        RECT 76.950 830.400 81.600 831.600 ;
        RECT 76.950 829.950 79.050 830.400 ;
        RECT 91.950 826.950 94.050 829.050 ;
        RECT 73.950 823.950 76.050 826.050 ;
        RECT 61.950 811.950 64.050 814.050 ;
        RECT 70.950 811.950 73.050 814.050 ;
        RECT 82.950 811.950 85.050 814.050 ;
        RECT 46.950 805.950 49.050 808.050 ;
        RECT 55.950 805.950 58.050 808.050 ;
        RECT 41.400 801.000 45.600 801.600 ;
        RECT 41.400 800.400 46.050 801.000 ;
        RECT 37.950 796.950 40.050 799.050 ;
        RECT 43.950 796.950 46.050 800.400 ;
        RECT 38.400 778.050 39.600 796.950 ;
        RECT 56.400 793.050 57.600 805.950 ;
        RECT 62.400 799.050 63.600 811.950 ;
        RECT 71.400 808.050 72.600 811.950 ;
        RECT 64.950 807.600 69.000 808.050 ;
        RECT 64.950 805.950 69.600 807.600 ;
        RECT 70.950 805.950 73.050 808.050 ;
        RECT 68.400 804.600 69.600 805.950 ;
        RECT 68.400 803.400 75.600 804.600 ;
        RECT 61.950 796.950 64.050 799.050 ;
        RECT 67.950 796.950 70.050 799.050 ;
        RECT 68.400 793.050 69.600 796.950 ;
        RECT 55.950 790.950 58.050 793.050 ;
        RECT 67.950 790.950 70.050 793.050 ;
        RECT 74.400 789.600 75.600 803.400 ;
        RECT 71.400 788.400 75.600 789.600 ;
        RECT 37.950 775.950 40.050 778.050 ;
        RECT 22.950 763.950 25.050 766.050 ;
        RECT 28.950 763.950 31.050 766.050 ;
        RECT 34.950 763.950 37.050 766.050 ;
        RECT 55.950 763.950 58.050 766.050 ;
        RECT 16.950 754.950 19.050 757.050 ;
        RECT 29.400 747.600 30.600 763.950 ;
        RECT 31.950 754.950 34.050 757.050 ;
        RECT 37.950 754.950 40.050 757.050 ;
        RECT 43.950 754.950 46.050 757.050 ;
        RECT 32.400 751.050 33.600 754.950 ;
        RECT 31.950 748.950 34.050 751.050 ;
        RECT 26.400 747.000 30.600 747.600 ;
        RECT 25.950 746.400 30.600 747.000 ;
        RECT 16.950 742.950 19.050 745.050 ;
        RECT 25.950 742.950 28.050 746.400 ;
        RECT 13.950 739.950 16.050 742.050 ;
        RECT 7.950 733.950 10.050 736.050 ;
        RECT 8.400 664.050 9.600 733.950 ;
        RECT 17.400 730.050 18.600 742.950 ;
        RECT 28.950 739.950 31.050 742.050 ;
        RECT 29.400 730.050 30.600 739.950 ;
        RECT 38.400 739.050 39.600 754.950 ;
        RECT 44.400 751.050 45.600 754.950 ;
        RECT 43.950 748.950 46.050 751.050 ;
        RECT 56.400 745.050 57.600 763.950 ;
        RECT 61.950 762.600 64.050 766.050 ;
        RECT 59.400 762.000 64.050 762.600 ;
        RECT 59.400 761.400 63.600 762.000 ;
        RECT 59.400 751.050 60.600 761.400 ;
        RECT 64.950 756.600 69.000 757.050 ;
        RECT 64.950 754.950 69.600 756.600 ;
        RECT 58.950 748.950 61.050 751.050 ;
        RECT 55.950 742.950 58.050 745.050 ;
        RECT 37.950 736.950 40.050 739.050 ;
        RECT 61.950 736.950 64.050 739.050 ;
        RECT 40.950 733.950 43.050 736.050 ;
        RECT 46.950 733.950 49.050 736.050 ;
        RECT 55.950 733.950 58.050 736.050 ;
        RECT 16.950 727.950 19.050 730.050 ;
        RECT 28.950 727.950 31.050 730.050 ;
        RECT 41.400 721.050 42.600 733.950 ;
        RECT 31.950 718.950 34.050 721.050 ;
        RECT 37.950 719.400 42.600 721.050 ;
        RECT 37.950 718.950 42.000 719.400 ;
        RECT 32.400 715.050 33.600 718.950 ;
        RECT 31.950 712.950 34.050 715.050 ;
        RECT 40.950 712.950 43.050 715.050 ;
        RECT 34.950 709.950 37.050 712.050 ;
        RECT 16.950 694.950 19.050 697.050 ;
        RECT 17.400 679.050 18.600 694.950 ;
        RECT 28.950 691.950 31.050 694.050 ;
        RECT 16.950 676.950 19.050 679.050 ;
        RECT 7.950 661.950 10.050 664.050 ;
        RECT 13.950 661.950 16.050 664.050 ;
        RECT 10.950 658.950 13.050 661.050 ;
        RECT 7.950 655.950 10.050 658.050 ;
        RECT 4.950 619.950 7.050 622.050 ;
        RECT 5.400 583.050 6.600 619.950 ;
        RECT 5.100 580.950 7.200 583.050 ;
        RECT 4.950 574.950 7.050 577.050 ;
        RECT 5.400 472.050 6.600 574.950 ;
        RECT 8.400 502.050 9.600 655.950 ;
        RECT 11.400 642.600 12.600 658.950 ;
        RECT 14.400 655.050 15.600 661.950 ;
        RECT 19.950 655.950 22.050 658.050 ;
        RECT 13.950 652.950 16.050 655.050 ;
        RECT 20.400 652.050 21.600 655.950 ;
        RECT 19.950 649.950 22.050 652.050 ;
        RECT 29.400 649.050 30.600 691.950 ;
        RECT 35.400 688.050 36.600 709.950 ;
        RECT 37.950 693.600 40.050 694.050 ;
        RECT 41.400 693.600 42.600 712.950 ;
        RECT 47.400 712.050 48.600 733.950 ;
        RECT 56.400 730.050 57.600 733.950 ;
        RECT 62.400 733.050 63.600 736.950 ;
        RECT 61.950 730.950 64.050 733.050 ;
        RECT 55.950 727.950 58.050 730.050 ;
        RECT 52.950 718.950 55.050 721.050 ;
        RECT 58.950 720.600 61.050 721.050 ;
        RECT 64.950 720.600 67.050 721.050 ;
        RECT 58.950 719.400 67.050 720.600 ;
        RECT 58.950 718.950 61.050 719.400 ;
        RECT 64.950 718.950 67.050 719.400 ;
        RECT 53.400 715.050 54.600 718.950 ;
        RECT 52.950 712.950 55.050 715.050 ;
        RECT 64.950 714.600 67.050 715.050 ;
        RECT 68.400 714.600 69.600 754.950 ;
        RECT 71.400 742.050 72.600 788.400 ;
        RECT 83.400 778.050 84.600 811.950 ;
        RECT 92.400 808.050 93.600 826.950 ;
        RECT 98.400 817.050 99.600 832.950 ;
        RECT 116.400 829.050 117.600 832.950 ;
        RECT 115.950 826.950 118.050 829.050 ;
        RECT 97.950 814.950 100.050 817.050 ;
        RECT 112.950 814.950 115.050 817.050 ;
        RECT 91.950 805.950 94.050 808.050 ;
        RECT 106.950 805.950 109.050 808.050 ;
        RECT 88.950 796.950 91.050 799.050 ;
        RECT 94.950 798.600 97.050 799.050 ;
        RECT 100.950 798.600 103.050 799.050 ;
        RECT 94.950 797.400 103.050 798.600 ;
        RECT 94.950 796.950 97.050 797.400 ;
        RECT 100.950 796.950 103.050 797.400 ;
        RECT 89.400 793.050 90.600 796.950 ;
        RECT 88.950 790.950 91.050 793.050 ;
        RECT 91.950 784.950 94.050 787.050 ;
        RECT 82.950 775.950 85.050 778.050 ;
        RECT 85.950 772.950 88.050 775.050 ;
        RECT 81.000 765.600 85.050 766.050 ;
        RECT 80.400 763.950 85.050 765.600 ;
        RECT 73.950 754.950 76.050 757.050 ;
        RECT 70.950 739.950 73.050 742.050 ;
        RECT 74.400 733.050 75.600 754.950 ;
        RECT 80.400 739.050 81.600 763.950 ;
        RECT 86.400 757.050 87.600 772.950 ;
        RECT 92.400 766.050 93.600 784.950 ;
        RECT 100.950 781.950 103.050 784.050 ;
        RECT 101.400 772.050 102.600 781.950 ;
        RECT 107.400 781.050 108.600 805.950 ;
        RECT 113.400 799.050 114.600 814.950 ;
        RECT 116.400 808.050 117.600 826.950 ;
        RECT 119.400 817.200 120.600 841.950 ;
        RECT 137.400 835.050 138.600 853.950 ;
        RECT 152.400 844.050 153.600 853.950 ;
        RECT 181.950 847.950 184.050 850.050 ;
        RECT 182.400 844.050 183.600 847.950 ;
        RECT 151.950 841.950 154.050 844.050 ;
        RECT 157.950 841.950 160.050 844.050 ;
        RECT 175.950 841.950 178.050 844.050 ;
        RECT 181.950 841.950 184.050 844.050 ;
        RECT 136.950 832.950 139.050 835.050 ;
        RECT 148.950 832.950 151.050 835.050 ;
        RECT 149.400 826.050 150.600 832.950 ;
        RECT 148.950 823.950 151.050 826.050 ;
        RECT 127.950 820.950 130.050 823.050 ;
        RECT 118.950 815.100 121.050 817.200 ;
        RECT 118.950 811.800 121.050 813.900 ;
        RECT 115.950 805.950 118.050 808.050 ;
        RECT 119.400 799.050 120.600 811.800 ;
        RECT 112.950 796.950 115.050 799.050 ;
        RECT 118.950 796.950 121.050 799.050 ;
        RECT 119.400 793.050 120.600 796.950 ;
        RECT 118.950 790.950 121.050 793.050 ;
        RECT 128.400 784.050 129.600 820.950 ;
        RECT 149.400 808.050 150.600 823.950 ;
        RECT 158.400 814.050 159.600 841.950 ;
        RECT 172.950 832.950 175.050 835.050 ;
        RECT 157.950 811.950 160.050 814.050 ;
        RECT 158.400 808.050 159.600 811.950 ;
        RECT 136.950 805.950 139.050 808.050 ;
        RECT 148.950 805.950 151.050 808.050 ;
        RECT 157.950 805.950 160.050 808.050 ;
        RECT 137.400 784.050 138.600 805.950 ;
        RECT 151.950 796.950 154.050 799.050 ;
        RECT 156.000 798.600 160.050 799.050 ;
        RECT 155.400 796.950 160.050 798.600 ;
        RECT 152.400 793.050 153.600 796.950 ;
        RECT 151.950 790.950 154.050 793.050 ;
        RECT 145.950 787.950 148.050 790.050 ;
        RECT 127.950 781.950 130.050 784.050 ;
        RECT 136.950 781.950 139.050 784.050 ;
        RECT 106.950 778.950 109.050 781.050 ;
        RECT 118.950 778.950 121.050 781.050 ;
        RECT 100.950 769.950 103.050 772.050 ;
        RECT 106.950 769.950 109.050 772.050 ;
        RECT 107.400 766.050 108.600 769.950 ;
        RECT 88.950 764.400 93.600 766.050 ;
        RECT 88.950 763.950 93.000 764.400 ;
        RECT 100.950 763.950 103.050 766.050 ;
        RECT 106.950 763.950 109.050 766.050 ;
        RECT 112.950 763.950 115.050 766.050 ;
        RECT 85.950 754.950 88.050 757.050 ;
        RECT 91.950 754.950 94.050 757.050 ;
        RECT 101.400 756.600 102.600 763.950 ;
        RECT 109.950 756.600 112.050 757.050 ;
        RECT 101.400 755.400 112.050 756.600 ;
        RECT 109.950 754.950 112.050 755.400 ;
        RECT 85.950 745.950 88.050 748.050 ;
        RECT 82.950 742.950 85.050 745.050 ;
        RECT 79.950 736.950 82.050 739.050 ;
        RECT 73.950 730.950 76.050 733.050 ;
        RECT 83.400 730.050 84.600 742.950 ;
        RECT 70.950 727.950 73.050 730.050 ;
        RECT 82.950 727.950 85.050 730.050 ;
        RECT 64.950 713.400 69.600 714.600 ;
        RECT 64.950 712.950 67.050 713.400 ;
        RECT 46.950 709.950 49.050 712.050 ;
        RECT 55.950 706.950 58.050 709.050 ;
        RECT 37.950 692.400 42.600 693.600 ;
        RECT 37.950 691.950 40.050 692.400 ;
        RECT 38.400 688.050 39.600 691.950 ;
        RECT 34.950 685.950 37.050 688.050 ;
        RECT 38.400 686.400 43.050 688.050 ;
        RECT 39.000 685.950 43.050 686.400 ;
        RECT 37.950 676.950 40.050 679.050 ;
        RECT 43.950 676.950 46.050 679.050 ;
        RECT 56.400 678.600 57.600 706.950 ;
        RECT 58.950 697.950 61.050 700.050 ;
        RECT 59.400 688.050 60.600 697.950 ;
        RECT 65.400 697.050 66.600 712.950 ;
        RECT 64.950 694.950 67.050 697.050 ;
        RECT 65.400 688.050 66.600 694.950 ;
        RECT 58.950 685.950 61.050 688.050 ;
        RECT 64.950 685.950 67.050 688.050 ;
        RECT 61.950 678.600 64.050 679.050 ;
        RECT 56.400 677.400 64.050 678.600 ;
        RECT 61.950 676.950 64.050 677.400 ;
        RECT 31.950 673.950 34.050 676.050 ;
        RECT 32.400 661.050 33.600 673.950 ;
        RECT 38.400 673.050 39.600 676.950 ;
        RECT 37.950 670.950 40.050 673.050 ;
        RECT 31.950 658.950 34.050 661.050 ;
        RECT 37.950 658.950 40.050 661.050 ;
        RECT 38.400 652.050 39.600 658.950 ;
        RECT 44.400 658.050 45.600 676.950 ;
        RECT 71.400 673.050 72.600 727.950 ;
        RECT 86.400 699.600 87.600 745.950 ;
        RECT 92.400 745.050 93.600 754.950 ;
        RECT 113.400 751.050 114.600 763.950 ;
        RECT 119.400 763.050 120.600 778.950 ;
        RECT 124.950 769.950 127.050 772.050 ;
        RECT 125.400 766.050 126.600 769.950 ;
        RECT 124.950 763.950 127.050 766.050 ;
        RECT 130.950 763.950 133.050 766.050 ;
        RECT 118.950 760.950 121.050 763.050 ;
        RECT 121.950 756.600 124.050 757.050 ;
        RECT 127.950 756.600 130.050 757.050 ;
        RECT 121.950 755.400 130.050 756.600 ;
        RECT 121.950 754.950 124.050 755.400 ;
        RECT 127.950 754.950 130.050 755.400 ;
        RECT 131.400 751.050 132.600 763.950 ;
        RECT 146.400 763.050 147.600 787.950 ;
        RECT 155.400 766.050 156.600 796.950 ;
        RECT 169.950 784.950 172.050 787.050 ;
        RECT 166.950 781.950 169.050 784.050 ;
        RECT 167.400 766.050 168.600 781.950 ;
        RECT 170.400 781.050 171.600 784.950 ;
        RECT 169.950 778.950 172.050 781.050 ;
        RECT 173.400 772.050 174.600 832.950 ;
        RECT 176.400 826.050 177.600 841.950 ;
        RECT 185.400 835.050 186.600 853.950 ;
        RECT 197.400 853.050 198.600 865.950 ;
        RECT 196.950 850.950 199.050 853.050 ;
        RECT 187.950 847.950 190.050 850.050 ;
        RECT 188.400 841.050 189.600 847.950 ;
        RECT 203.400 847.050 204.600 883.950 ;
        RECT 223.950 874.950 226.050 877.050 ;
        RECT 211.950 865.950 214.050 868.050 ;
        RECT 193.950 844.950 196.050 847.050 ;
        RECT 202.950 844.950 205.050 847.050 ;
        RECT 187.950 838.950 190.050 841.050 ;
        RECT 184.950 832.950 187.050 835.050 ;
        RECT 175.950 823.950 178.050 826.050 ;
        RECT 181.950 820.950 184.050 823.050 ;
        RECT 178.950 811.950 181.050 814.050 ;
        RECT 179.400 799.050 180.600 811.950 ;
        RECT 182.400 808.050 183.600 820.950 ;
        RECT 194.400 820.050 195.600 844.950 ;
        RECT 196.950 829.950 199.050 832.050 ;
        RECT 202.950 829.950 205.050 832.050 ;
        RECT 193.950 817.950 196.050 820.050 ;
        RECT 197.400 808.050 198.600 829.950 ;
        RECT 203.400 826.050 204.600 829.950 ;
        RECT 202.950 823.950 205.050 826.050 ;
        RECT 205.950 820.950 208.050 823.050 ;
        RECT 206.400 811.050 207.600 820.950 ;
        RECT 212.400 817.050 213.600 865.950 ;
        RECT 224.400 859.050 225.600 874.950 ;
        RECT 230.400 871.050 231.600 883.950 ;
        RECT 229.950 868.950 232.050 871.050 ;
        RECT 236.400 865.050 237.600 883.950 ;
        RECT 251.400 879.600 252.600 883.950 ;
        RECT 245.400 879.000 252.600 879.600 ;
        RECT 244.950 878.400 252.600 879.000 ;
        RECT 238.950 874.950 241.050 877.050 ;
        RECT 244.950 874.950 247.050 878.400 ;
        RECT 274.950 877.950 277.050 880.050 ;
        RECT 259.950 876.600 264.000 877.050 ;
        RECT 259.950 874.950 264.600 876.600 ;
        RECT 265.950 874.950 268.050 877.050 ;
        RECT 239.400 871.050 240.600 874.950 ;
        RECT 238.950 868.950 241.050 871.050 ;
        RECT 263.400 865.050 264.600 874.950 ;
        RECT 266.400 868.050 267.600 874.950 ;
        RECT 266.100 865.950 268.200 868.050 ;
        RECT 235.950 862.950 238.050 865.050 ;
        RECT 262.950 862.950 265.050 865.050 ;
        RECT 268.950 862.950 271.050 865.050 ;
        RECT 223.950 856.950 226.050 859.050 ;
        RECT 259.950 856.950 262.050 859.050 ;
        RECT 223.950 850.950 226.050 853.050 ;
        RECT 224.400 832.050 225.600 850.950 ;
        RECT 226.950 847.950 229.050 850.050 ;
        RECT 217.950 829.950 220.050 832.050 ;
        RECT 223.950 829.950 226.050 832.050 ;
        RECT 218.400 826.050 219.600 829.950 ;
        RECT 217.950 823.950 220.050 826.050 ;
        RECT 220.950 820.950 223.050 823.050 ;
        RECT 211.950 814.950 214.050 817.050 ;
        RECT 221.400 813.600 222.600 820.950 ;
        RECT 227.400 814.050 228.600 847.950 ;
        RECT 238.950 841.950 241.050 844.050 ;
        RECT 244.950 841.950 247.050 844.050 ;
        RECT 229.950 832.950 232.050 835.050 ;
        RECT 230.400 826.050 231.600 832.950 ;
        RECT 229.950 823.950 232.050 826.050 ;
        RECT 239.400 823.050 240.600 841.950 ;
        RECT 245.400 826.050 246.600 841.950 ;
        RECT 260.400 841.050 261.600 856.950 ;
        RECT 262.950 853.950 265.050 856.050 ;
        RECT 259.950 838.950 262.050 841.050 ;
        RECT 244.950 823.950 247.050 826.050 ;
        RECT 238.950 820.950 241.050 823.050 ;
        RECT 260.400 817.050 261.600 838.950 ;
        RECT 263.400 832.050 264.600 853.950 ;
        RECT 269.400 847.050 270.600 862.950 ;
        RECT 275.400 856.050 276.600 877.950 ;
        RECT 274.950 853.950 277.050 856.050 ;
        RECT 268.950 844.950 271.050 847.050 ;
        RECT 271.950 838.950 274.050 841.050 ;
        RECT 262.950 829.950 265.050 832.050 ;
        RECT 268.950 829.950 271.050 832.050 ;
        RECT 269.400 826.050 270.600 829.950 ;
        RECT 268.950 823.950 271.050 826.050 ;
        RECT 272.400 823.050 273.600 838.950 ;
        RECT 271.950 820.950 274.050 823.050 ;
        RECT 262.950 817.950 265.050 820.050 ;
        RECT 259.950 814.950 262.050 817.050 ;
        RECT 218.400 812.400 222.600 813.600 ;
        RECT 205.950 808.950 208.050 811.050 ;
        RECT 218.400 808.050 219.600 812.400 ;
        RECT 226.950 811.950 229.050 814.050 ;
        RECT 181.950 805.950 184.050 808.050 ;
        RECT 196.950 805.950 199.050 808.050 ;
        RECT 218.400 805.950 223.050 808.050 ;
        RECT 259.950 805.950 262.050 808.050 ;
        RECT 190.950 802.950 193.050 805.050 ;
        RECT 178.950 796.950 181.050 799.050 ;
        RECT 179.400 784.050 180.600 796.950 ;
        RECT 181.950 784.950 184.050 787.050 ;
        RECT 178.950 781.950 181.050 784.050 ;
        RECT 172.950 769.950 175.050 772.050 ;
        RECT 178.950 769.950 181.050 772.050 ;
        RECT 179.400 766.050 180.600 769.950 ;
        RECT 154.950 763.950 157.050 766.050 ;
        RECT 145.950 760.950 148.050 763.050 ;
        RECT 139.950 754.950 142.050 757.050 ;
        RECT 133.950 751.950 136.050 754.050 ;
        RECT 97.950 748.950 100.050 751.050 ;
        RECT 112.950 748.950 115.050 751.050 ;
        RECT 130.950 748.950 133.050 751.050 ;
        RECT 98.400 745.050 99.600 748.950 ;
        RECT 106.950 745.950 109.050 748.050 ;
        RECT 118.950 745.950 121.050 748.050 ;
        RECT 91.950 742.950 94.050 745.050 ;
        RECT 97.950 742.950 100.050 745.050 ;
        RECT 88.950 739.950 91.050 742.050 ;
        RECT 89.400 708.600 90.600 739.950 ;
        RECT 97.950 736.950 100.050 739.050 ;
        RECT 98.400 721.050 99.600 736.950 ;
        RECT 107.400 730.050 108.600 745.950 ;
        RECT 112.950 733.950 115.050 736.050 ;
        RECT 106.950 727.950 109.050 730.050 ;
        RECT 97.950 718.950 100.050 721.050 ;
        RECT 103.950 720.600 108.000 721.050 ;
        RECT 103.950 720.000 108.600 720.600 ;
        RECT 103.950 718.950 109.050 720.000 ;
        RECT 106.950 715.950 109.050 718.950 ;
        RECT 89.400 707.400 93.600 708.600 ;
        RECT 86.400 699.000 90.600 699.600 ;
        RECT 86.400 698.400 91.050 699.000 ;
        RECT 88.950 694.950 91.050 698.400 ;
        RECT 85.950 691.950 88.050 694.050 ;
        RECT 86.400 679.050 87.600 691.950 ;
        RECT 82.950 677.400 87.600 679.050 ;
        RECT 82.950 676.950 87.000 677.400 ;
        RECT 70.950 670.950 73.050 673.050 ;
        RECT 88.950 667.950 91.050 670.050 ;
        RECT 55.950 661.950 58.050 664.050 ;
        RECT 85.950 661.950 88.050 664.050 ;
        RECT 43.950 655.950 46.050 658.050 ;
        RECT 37.950 649.950 40.050 652.050 ;
        RECT 49.950 649.950 52.050 652.050 ;
        RECT 28.950 646.950 31.050 649.050 ;
        RECT 32.400 644.400 42.600 645.600 ;
        RECT 16.950 642.600 19.050 643.050 ;
        RECT 11.400 641.400 19.050 642.600 ;
        RECT 16.950 640.950 19.050 641.400 ;
        RECT 22.950 642.600 25.050 643.050 ;
        RECT 32.400 642.600 33.600 644.400 ;
        RECT 41.400 643.050 42.600 644.400 ;
        RECT 22.950 641.400 33.600 642.600 ;
        RECT 22.950 640.950 25.050 641.400 ;
        RECT 34.950 640.950 37.050 643.050 ;
        RECT 40.950 642.600 43.050 643.050 ;
        RECT 46.950 642.600 49.050 643.050 ;
        RECT 40.950 641.400 49.050 642.600 ;
        RECT 40.950 640.950 43.050 641.400 ;
        RECT 46.950 640.950 49.050 641.400 ;
        RECT 35.400 637.050 36.600 640.950 ;
        RECT 34.950 634.950 37.050 637.050 ;
        RECT 16.950 628.950 19.050 631.050 ;
        RECT 10.950 625.950 13.050 628.050 ;
        RECT 11.400 586.050 12.600 625.950 ;
        RECT 17.400 610.050 18.600 628.950 ;
        RECT 19.950 625.950 22.050 628.050 ;
        RECT 20.400 610.050 21.600 625.950 ;
        RECT 50.400 625.050 51.600 649.950 ;
        RECT 25.950 622.950 28.050 625.050 ;
        RECT 49.950 622.950 52.050 625.050 ;
        RECT 13.950 608.400 18.600 610.050 ;
        RECT 13.950 607.950 18.000 608.400 ;
        RECT 19.950 607.950 22.050 610.050 ;
        RECT 16.950 598.950 19.050 601.050 ;
        RECT 17.400 595.050 18.600 598.950 ;
        RECT 16.950 592.950 19.050 595.050 ;
        RECT 10.950 583.950 13.050 586.050 ;
        RECT 19.950 580.950 22.050 583.050 ;
        RECT 13.950 577.950 16.050 580.050 ;
        RECT 14.400 565.050 15.600 577.950 ;
        RECT 16.950 571.950 19.050 574.050 ;
        RECT 13.950 562.950 16.050 565.050 ;
        RECT 17.400 559.050 18.600 571.950 ;
        RECT 20.400 565.050 21.600 580.950 ;
        RECT 19.950 562.950 22.050 565.050 ;
        RECT 16.950 556.950 19.050 559.050 ;
        RECT 26.400 541.050 27.600 622.950 ;
        RECT 37.950 619.950 40.050 622.050 ;
        RECT 43.950 619.950 46.050 622.050 ;
        RECT 38.400 610.050 39.600 619.950 ;
        RECT 44.400 610.050 45.600 619.950 ;
        RECT 37.950 607.950 40.050 610.050 ;
        RECT 43.950 607.950 46.050 610.050 ;
        RECT 40.950 598.950 43.050 601.050 ;
        RECT 34.950 595.950 37.050 598.050 ;
        RECT 35.400 574.050 36.600 595.950 ;
        RECT 41.400 591.600 42.600 598.950 ;
        RECT 46.950 592.950 49.050 595.050 ;
        RECT 41.400 591.000 45.600 591.600 ;
        RECT 41.400 590.400 46.050 591.000 ;
        RECT 43.950 586.950 46.050 590.400 ;
        RECT 40.950 583.950 43.050 586.050 ;
        RECT 41.400 574.050 42.600 583.950 ;
        RECT 34.950 571.950 37.050 574.050 ;
        RECT 40.950 571.950 43.050 574.050 ;
        RECT 30.000 564.600 34.050 565.050 ;
        RECT 29.400 562.950 34.050 564.600 ;
        RECT 37.950 562.950 40.050 565.050 ;
        RECT 25.950 538.950 28.050 541.050 ;
        RECT 29.400 535.050 30.600 562.950 ;
        RECT 38.400 559.050 39.600 562.950 ;
        RECT 31.950 556.950 34.050 559.050 ;
        RECT 37.950 556.950 40.050 559.050 ;
        RECT 32.400 547.050 33.600 556.950 ;
        RECT 31.950 544.950 34.050 547.050 ;
        RECT 28.950 532.950 31.050 535.050 ;
        RECT 13.950 531.600 16.050 532.050 ;
        RECT 19.950 531.600 22.050 532.050 ;
        RECT 13.950 530.400 22.050 531.600 ;
        RECT 13.950 529.950 16.050 530.400 ;
        RECT 19.950 529.950 22.050 530.400 ;
        RECT 32.400 523.050 33.600 544.950 ;
        RECT 47.400 538.050 48.600 592.950 ;
        RECT 56.400 592.050 57.600 661.950 ;
        RECT 64.950 658.950 67.050 661.050 ;
        RECT 65.400 652.050 66.600 658.950 ;
        RECT 86.400 655.050 87.600 661.950 ;
        RECT 64.950 649.950 67.050 652.050 ;
        RECT 79.950 651.600 82.050 655.050 ;
        RECT 85.950 652.950 88.050 655.050 ;
        RECT 77.400 651.000 82.050 651.600 ;
        RECT 77.400 650.400 81.600 651.000 ;
        RECT 70.950 643.950 73.050 646.050 ;
        RECT 64.950 607.950 67.050 610.050 ;
        RECT 49.950 589.950 52.050 592.050 ;
        RECT 55.950 589.950 58.050 592.050 ;
        RECT 34.950 535.950 37.050 538.050 ;
        RECT 40.950 535.950 43.050 538.050 ;
        RECT 46.950 535.950 49.050 538.050 ;
        RECT 35.400 532.050 36.600 535.950 ;
        RECT 41.400 532.050 42.600 535.950 ;
        RECT 34.950 529.950 37.050 532.050 ;
        RECT 40.950 529.950 43.050 532.050 ;
        RECT 50.400 525.600 51.600 589.950 ;
        RECT 52.950 586.950 55.050 589.050 ;
        RECT 53.400 556.050 54.600 586.950 ;
        RECT 65.400 580.050 66.600 607.950 ;
        RECT 71.400 607.050 72.600 643.950 ;
        RECT 77.400 643.050 78.600 650.400 ;
        RECT 76.950 640.950 79.050 643.050 ;
        RECT 82.950 637.950 85.050 640.050 ;
        RECT 79.950 609.600 82.050 610.050 ;
        RECT 74.400 608.400 82.050 609.600 ;
        RECT 70.950 604.950 73.050 607.050 ;
        RECT 74.400 601.050 75.600 608.400 ;
        RECT 79.950 607.950 82.050 608.400 ;
        RECT 73.800 598.950 75.900 601.050 ;
        RECT 70.950 589.950 73.050 592.050 ;
        RECT 58.950 577.950 61.050 580.050 ;
        RECT 64.950 577.950 67.050 580.050 ;
        RECT 59.400 565.050 60.600 577.950 ;
        RECT 67.950 571.950 70.050 574.050 ;
        RECT 68.400 567.600 69.600 571.950 ;
        RECT 62.400 566.400 69.600 567.600 ;
        RECT 62.400 565.050 63.600 566.400 ;
        RECT 58.950 563.400 63.600 565.050 ;
        RECT 58.950 562.950 63.000 563.400 ;
        RECT 64.950 562.950 67.050 565.050 ;
        RECT 65.400 559.050 66.600 562.950 ;
        RECT 64.950 556.950 67.050 559.050 ;
        RECT 52.950 553.950 55.050 556.050 ;
        RECT 71.400 553.050 72.600 589.950 ;
        RECT 83.400 583.050 84.600 637.950 ;
        RECT 89.400 610.050 90.600 667.950 ;
        RECT 92.400 640.050 93.600 707.400 ;
        RECT 106.950 706.950 109.050 709.050 ;
        RECT 100.950 703.950 103.050 706.050 ;
        RECT 95.100 694.950 97.200 697.050 ;
        RECT 95.400 688.050 96.600 694.950 ;
        RECT 101.400 688.050 102.600 703.950 ;
        RECT 107.400 688.050 108.600 706.950 ;
        RECT 113.400 700.050 114.600 733.950 ;
        RECT 119.400 730.050 120.600 745.950 ;
        RECT 124.950 739.950 127.050 742.050 ;
        RECT 118.950 727.950 121.050 730.050 ;
        RECT 125.400 723.600 126.600 739.950 ;
        RECT 127.950 735.600 130.050 736.050 ;
        RECT 131.400 735.600 132.600 748.950 ;
        RECT 134.400 745.050 135.600 751.950 ;
        RECT 133.950 742.950 136.050 745.050 ;
        RECT 127.950 734.400 132.600 735.600 ;
        RECT 127.950 733.950 130.050 734.400 ;
        RECT 122.400 723.000 126.600 723.600 ;
        RECT 121.950 722.400 126.600 723.000 ;
        RECT 121.950 718.950 124.050 722.400 ;
        RECT 128.400 721.050 129.600 733.950 ;
        RECT 127.950 718.950 130.050 721.050 ;
        RECT 121.950 709.950 124.050 712.050 ;
        RECT 112.950 697.950 115.050 700.050 ;
        RECT 118.950 691.950 121.050 694.050 ;
        RECT 94.950 685.950 97.050 688.050 ;
        RECT 100.950 685.950 103.050 688.050 ;
        RECT 106.950 685.950 109.050 688.050 ;
        RECT 95.400 678.600 96.600 685.950 ;
        RECT 119.400 679.050 120.600 691.950 ;
        RECT 122.400 688.050 123.600 709.950 ;
        RECT 140.400 706.050 141.600 754.950 ;
        RECT 151.950 751.950 154.050 754.050 ;
        RECT 142.950 727.950 145.050 730.050 ;
        RECT 139.950 703.950 142.050 706.050 ;
        RECT 136.950 700.950 139.050 703.050 ;
        RECT 127.950 697.950 130.050 700.050 ;
        RECT 128.400 688.050 129.600 697.950 ;
        RECT 121.950 685.950 124.050 688.050 ;
        RECT 127.950 685.950 130.050 688.050 ;
        RECT 137.400 684.600 138.600 700.950 ;
        RECT 143.400 700.050 144.600 727.950 ;
        RECT 152.400 721.050 153.600 751.950 ;
        RECT 155.400 751.050 156.600 763.950 ;
        RECT 160.950 762.600 163.050 766.050 ;
        RECT 166.950 763.950 169.050 766.050 ;
        RECT 178.950 763.950 181.050 766.050 ;
        RECT 160.950 762.000 165.600 762.600 ;
        RECT 161.400 761.400 166.050 762.000 ;
        RECT 163.950 757.950 166.050 761.400 ;
        RECT 182.400 757.050 183.600 784.950 ;
        RECT 184.800 771.600 189.000 772.050 ;
        RECT 184.800 769.950 189.600 771.600 ;
        RECT 188.400 757.050 189.600 769.950 ;
        RECT 157.950 754.950 160.050 757.050 ;
        RECT 166.950 754.950 169.050 757.050 ;
        RECT 181.950 754.950 184.050 757.050 ;
        RECT 187.950 754.950 190.050 757.050 ;
        RECT 154.950 748.950 157.050 751.050 ;
        RECT 158.400 748.050 159.600 754.950 ;
        RECT 157.950 745.950 160.050 748.050 ;
        RECT 163.950 745.950 166.050 748.050 ;
        RECT 157.950 733.950 160.050 736.050 ;
        RECT 145.950 718.950 148.050 721.050 ;
        RECT 151.950 718.950 154.050 721.050 ;
        RECT 146.400 714.600 147.600 718.950 ;
        RECT 146.400 713.400 150.600 714.600 ;
        RECT 142.950 697.950 145.050 700.050 ;
        RECT 149.400 694.050 150.600 713.400 ;
        RECT 151.950 703.950 154.050 706.050 ;
        RECT 148.950 691.950 151.050 694.050 ;
        RECT 149.400 688.050 150.600 691.950 ;
        RECT 148.950 685.950 151.050 688.050 ;
        RECT 152.400 685.050 153.600 703.950 ;
        RECT 158.400 703.050 159.600 733.950 ;
        RECT 157.950 700.950 160.050 703.050 ;
        RECT 164.400 687.600 165.600 745.950 ;
        RECT 167.400 742.050 168.600 754.950 ;
        RECT 178.950 745.950 181.050 748.050 ;
        RECT 166.950 739.950 169.050 742.050 ;
        RECT 175.950 736.950 178.050 739.050 ;
        RECT 176.400 733.050 177.600 736.950 ;
        RECT 179.400 736.050 180.600 745.950 ;
        RECT 191.400 739.050 192.600 802.950 ;
        RECT 218.400 801.600 219.600 805.950 ;
        RECT 215.400 800.400 219.600 801.600 ;
        RECT 196.950 796.950 199.050 799.050 ;
        RECT 202.950 796.950 205.050 799.050 ;
        RECT 197.400 793.050 198.600 796.950 ;
        RECT 196.950 790.950 199.050 793.050 ;
        RECT 203.400 787.050 204.600 796.950 ;
        RECT 208.950 793.950 211.050 796.050 ;
        RECT 209.400 790.050 210.600 793.950 ;
        RECT 215.400 793.050 216.600 800.400 ;
        RECT 226.950 799.950 229.050 802.050 ;
        RECT 217.950 796.950 220.050 799.050 ;
        RECT 214.950 790.950 217.050 793.050 ;
        RECT 218.400 792.600 219.600 796.950 ;
        RECT 227.400 793.050 228.600 799.950 ;
        RECT 218.400 791.400 222.600 792.600 ;
        RECT 208.800 787.950 210.900 790.050 ;
        RECT 199.800 784.950 201.900 787.050 ;
        RECT 203.100 784.950 205.200 787.050 ;
        RECT 200.400 781.050 201.600 784.950 ;
        RECT 208.950 781.950 211.050 784.050 ;
        RECT 193.950 778.950 196.050 781.050 ;
        RECT 199.950 778.950 202.050 781.050 ;
        RECT 194.400 772.050 195.600 778.950 ;
        RECT 209.400 775.050 210.600 781.950 ;
        RECT 211.950 778.950 214.050 781.050 ;
        RECT 208.950 772.950 211.050 775.050 ;
        RECT 193.950 769.950 196.050 772.050 ;
        RECT 196.950 763.950 199.050 766.050 ;
        RECT 197.400 745.050 198.600 763.950 ;
        RECT 212.400 757.050 213.600 778.950 ;
        RECT 211.950 754.950 214.050 757.050 ;
        RECT 205.950 745.950 208.050 748.050 ;
        RECT 196.950 742.950 199.050 745.050 ;
        RECT 190.950 736.950 193.050 739.050 ;
        RECT 196.800 736.950 198.900 739.050 ;
        RECT 200.100 736.950 202.200 739.050 ;
        RECT 178.950 733.950 181.050 736.050 ;
        RECT 197.400 733.050 198.600 736.950 ;
        RECT 175.950 730.950 178.050 733.050 ;
        RECT 169.950 729.600 172.050 730.050 ;
        RECT 190.950 729.600 193.050 733.050 ;
        RECT 196.950 730.950 199.050 733.050 ;
        RECT 169.950 728.400 180.600 729.600 ;
        RECT 190.950 729.000 195.600 729.600 ;
        RECT 191.400 728.400 195.600 729.000 ;
        RECT 169.950 727.950 172.050 728.400 ;
        RECT 166.950 718.950 169.050 721.050 ;
        RECT 172.950 718.950 175.050 721.050 ;
        RECT 167.400 709.050 168.600 718.950 ;
        RECT 173.400 712.050 174.600 718.950 ;
        RECT 179.400 714.600 180.600 728.400 ;
        RECT 187.950 715.950 190.050 718.050 ;
        RECT 176.400 713.400 180.600 714.600 ;
        RECT 172.950 709.950 175.050 712.050 ;
        RECT 166.950 706.950 169.050 709.050 ;
        RECT 167.400 703.050 168.600 706.950 ;
        RECT 166.950 700.950 169.050 703.050 ;
        RECT 176.400 697.050 177.600 713.400 ;
        RECT 185.100 709.950 187.200 712.050 ;
        RECT 175.800 694.950 177.900 697.050 ;
        RECT 179.100 694.950 181.200 697.050 ;
        RECT 172.950 691.950 175.050 694.050 ;
        RECT 173.400 688.050 174.600 691.950 ;
        RECT 179.400 688.050 180.600 694.950 ;
        RECT 164.400 686.400 168.600 687.600 ;
        RECT 142.950 684.600 145.050 685.050 ;
        RECT 137.400 683.400 145.050 684.600 ;
        RECT 152.400 683.400 157.050 685.050 ;
        RECT 103.950 678.600 106.050 679.050 ;
        RECT 95.400 677.400 106.050 678.600 ;
        RECT 103.950 676.950 106.050 677.400 ;
        RECT 118.950 676.950 121.050 679.050 ;
        RECT 106.950 670.950 109.050 673.050 ;
        RECT 112.950 670.950 115.050 673.050 ;
        RECT 97.950 661.950 100.050 664.050 ;
        RECT 94.950 655.950 97.050 658.050 ;
        RECT 91.950 637.950 94.050 640.050 ;
        RECT 91.950 631.950 94.050 634.050 ;
        RECT 92.400 619.050 93.600 631.950 ;
        RECT 91.950 616.950 94.050 619.050 ;
        RECT 85.950 608.400 90.600 610.050 ;
        RECT 85.950 607.950 90.000 608.400 ;
        RECT 95.400 601.050 96.600 655.950 ;
        RECT 98.400 652.050 99.600 661.950 ;
        RECT 107.400 652.050 108.600 670.950 ;
        RECT 97.950 649.950 100.050 652.050 ;
        RECT 106.950 649.950 109.050 652.050 ;
        RECT 113.400 643.050 114.600 670.950 ;
        RECT 137.400 667.050 138.600 683.400 ;
        RECT 142.950 682.950 145.050 683.400 ;
        RECT 153.000 682.950 157.050 683.400 ;
        RECT 163.950 682.950 166.050 685.050 ;
        RECT 157.950 678.600 160.050 679.050 ;
        RECT 149.400 677.400 160.050 678.600 ;
        RECT 149.400 676.050 150.600 677.400 ;
        RECT 157.950 676.950 160.050 677.400 ;
        RECT 145.950 674.400 150.600 676.050 ;
        RECT 145.950 673.950 150.000 674.400 ;
        RECT 151.950 673.950 154.050 676.050 ;
        RECT 152.400 670.050 153.600 673.950 ;
        RECT 151.950 667.950 154.050 670.050 ;
        RECT 136.950 664.950 139.050 667.050 ;
        RECT 130.950 658.950 133.050 661.050 ;
        RECT 131.400 655.050 132.600 658.950 ;
        RECT 137.400 658.050 138.600 664.950 ;
        RECT 136.950 655.950 139.050 658.050 ;
        RECT 130.950 652.950 133.050 655.050 ;
        RECT 164.400 652.050 165.600 682.950 ;
        RECT 167.400 670.050 168.600 686.400 ;
        RECT 172.950 685.950 175.050 688.050 ;
        RECT 178.950 685.950 181.050 688.050 ;
        RECT 169.950 676.950 172.050 679.050 ;
        RECT 166.950 667.950 169.050 670.050 ;
        RECT 170.400 661.050 171.600 676.950 ;
        RECT 185.400 673.050 186.600 709.950 ;
        RECT 188.400 703.050 189.600 715.950 ;
        RECT 187.950 700.950 190.050 703.050 ;
        RECT 190.950 694.950 193.050 697.050 ;
        RECT 191.400 679.050 192.600 694.950 ;
        RECT 194.400 688.050 195.600 728.400 ;
        RECT 200.400 694.050 201.600 736.950 ;
        RECT 206.400 699.600 207.600 745.950 ;
        RECT 215.400 739.050 216.600 790.950 ;
        RECT 217.950 787.950 220.050 790.050 ;
        RECT 218.400 775.050 219.600 787.950 ;
        RECT 217.950 772.950 220.050 775.050 ;
        RECT 221.400 766.050 222.600 791.400 ;
        RECT 226.950 790.950 229.050 793.050 ;
        RECT 247.950 790.950 250.050 793.050 ;
        RECT 235.950 787.950 238.050 790.050 ;
        RECT 236.400 784.050 237.600 787.950 ;
        RECT 248.400 787.050 249.600 790.950 ;
        RECT 247.950 784.950 250.050 787.050 ;
        RECT 226.950 781.950 229.050 784.050 ;
        RECT 235.950 781.950 238.050 784.050 ;
        RECT 227.400 766.050 228.600 781.950 ;
        RECT 232.950 778.950 235.050 781.050 ;
        RECT 220.950 763.950 223.050 766.050 ;
        RECT 226.950 763.950 229.050 766.050 ;
        RECT 221.400 751.050 222.600 763.950 ;
        RECT 233.400 759.600 234.600 778.950 ;
        RECT 248.400 766.050 249.600 784.950 ;
        RECT 253.950 775.950 256.050 778.050 ;
        RECT 247.950 763.950 250.050 766.050 ;
        RECT 230.400 759.000 234.600 759.600 ;
        RECT 229.950 758.400 234.600 759.000 ;
        RECT 229.950 754.950 232.050 758.400 ;
        RECT 244.950 754.950 247.050 757.050 ;
        RECT 220.950 748.950 223.050 751.050 ;
        RECT 245.400 745.050 246.600 754.950 ;
        RECT 248.400 751.050 249.600 763.950 ;
        RECT 247.950 748.950 250.050 751.050 ;
        RECT 223.950 742.950 226.050 745.050 ;
        RECT 244.950 742.950 247.050 745.050 ;
        RECT 214.950 736.950 217.050 739.050 ;
        RECT 208.950 733.950 211.050 736.050 ;
        RECT 209.400 712.050 210.600 733.950 ;
        RECT 211.950 729.600 214.050 730.050 ;
        RECT 217.950 729.600 220.050 730.050 ;
        RECT 211.950 728.400 220.050 729.600 ;
        RECT 211.950 727.950 214.050 728.400 ;
        RECT 208.950 709.950 211.050 712.050 ;
        RECT 211.950 703.950 214.050 706.050 ;
        RECT 203.400 698.400 207.600 699.600 ;
        RECT 199.950 691.950 202.050 694.050 ;
        RECT 203.400 688.050 204.600 698.400 ;
        RECT 205.950 694.950 208.050 697.050 ;
        RECT 193.950 687.600 198.000 688.050 ;
        RECT 193.950 685.950 198.600 687.600 ;
        RECT 199.950 686.400 204.600 688.050 ;
        RECT 199.950 685.950 204.000 686.400 ;
        RECT 197.400 684.600 198.600 685.950 ;
        RECT 197.400 683.400 201.600 684.600 ;
        RECT 190.950 676.950 193.050 679.050 ;
        RECT 172.950 670.950 175.050 673.050 ;
        RECT 184.950 670.950 187.050 673.050 ;
        RECT 193.950 670.950 196.050 673.050 ;
        RECT 169.950 658.950 172.050 661.050 ;
        RECT 118.950 651.600 121.050 652.050 ;
        RECT 124.950 651.600 127.050 652.050 ;
        RECT 118.950 650.400 127.050 651.600 ;
        RECT 164.400 650.400 169.050 652.050 ;
        RECT 118.950 649.950 121.050 650.400 ;
        RECT 124.950 649.950 127.050 650.400 ;
        RECT 165.000 649.950 169.050 650.400 ;
        RECT 139.950 643.950 142.050 646.050 ;
        RECT 148.950 643.950 151.050 646.050 ;
        RECT 103.950 640.950 106.050 643.050 ;
        RECT 109.950 640.950 114.600 643.050 ;
        RECT 121.950 640.950 124.050 643.050 ;
        RECT 127.950 640.950 130.050 643.050 ;
        RECT 104.400 625.050 105.600 640.950 ;
        RECT 113.400 637.050 114.600 640.950 ;
        RECT 112.950 634.950 115.050 637.050 ;
        RECT 122.400 625.050 123.600 640.950 ;
        RECT 128.400 637.050 129.600 640.950 ;
        RECT 127.950 634.950 130.050 637.050 ;
        RECT 133.950 631.950 136.050 634.050 ;
        RECT 103.950 622.950 106.050 625.050 ;
        RECT 121.950 622.950 124.050 625.050 ;
        RECT 100.950 619.950 103.050 622.050 ;
        RECT 88.950 598.950 91.050 601.050 ;
        RECT 94.950 598.950 97.050 601.050 ;
        RECT 73.950 580.950 76.050 583.050 ;
        RECT 82.950 580.950 85.050 583.050 ;
        RECT 74.400 559.050 75.600 580.950 ;
        RECT 89.400 580.050 90.600 598.950 ;
        RECT 101.400 586.050 102.600 619.950 ;
        RECT 127.950 616.950 130.050 619.050 ;
        RECT 121.950 609.600 124.050 613.050 ;
        RECT 119.400 609.000 124.050 609.600 ;
        RECT 119.400 608.400 123.600 609.000 ;
        RECT 112.950 606.600 115.050 607.050 ;
        RECT 119.400 606.600 120.600 608.400 ;
        RECT 128.400 607.050 129.600 616.950 ;
        RECT 134.400 616.050 135.600 631.950 ;
        RECT 140.400 619.050 141.600 643.950 ;
        RECT 139.950 616.950 142.050 619.050 ;
        RECT 149.400 616.050 150.600 643.950 ;
        RECT 169.950 642.750 172.050 643.200 ;
        RECT 158.400 642.000 172.050 642.750 ;
        RECT 157.950 641.550 172.050 642.000 ;
        RECT 151.950 637.950 154.050 640.050 ;
        RECT 157.950 637.950 160.050 641.550 ;
        RECT 169.950 641.100 172.050 641.550 ;
        RECT 133.950 613.950 136.050 616.050 ;
        RECT 148.950 613.950 151.050 616.050 ;
        RECT 152.400 613.050 153.600 637.950 ;
        RECT 169.950 637.800 172.050 639.900 ;
        RECT 170.400 630.600 171.600 637.800 ;
        RECT 155.400 630.000 171.600 630.600 ;
        RECT 154.950 629.400 171.600 630.000 ;
        RECT 154.950 625.950 157.050 629.400 ;
        RECT 160.950 625.950 163.050 628.050 ;
        RECT 151.950 610.950 154.050 613.050 ;
        RECT 139.950 607.950 142.050 610.050 ;
        RECT 112.950 605.400 120.600 606.600 ;
        RECT 112.950 604.950 115.050 605.400 ;
        RECT 121.950 604.950 124.050 607.050 ;
        RECT 127.950 604.950 130.050 607.050 ;
        RECT 122.400 586.050 123.600 604.950 ;
        RECT 140.400 595.050 141.600 607.950 ;
        RECT 154.950 604.950 157.050 607.050 ;
        RECT 148.950 598.950 151.050 601.050 ;
        RECT 139.950 592.950 142.050 595.050 ;
        RECT 145.950 592.950 148.050 595.050 ;
        RECT 94.950 583.950 97.050 586.050 ;
        RECT 100.950 583.950 103.050 586.050 ;
        RECT 112.950 583.950 115.050 586.050 ;
        RECT 121.950 583.950 124.050 586.050 ;
        RECT 139.950 583.950 142.050 586.050 ;
        RECT 88.950 577.950 91.050 580.050 ;
        RECT 95.400 576.600 96.600 583.950 ;
        RECT 92.400 575.400 96.600 576.600 ;
        RECT 92.400 570.600 93.600 575.400 ;
        RECT 97.950 571.950 100.050 574.050 ;
        RECT 106.950 571.950 109.050 574.050 ;
        RECT 89.400 569.400 93.600 570.600 ;
        RECT 89.400 565.050 90.600 569.400 ;
        RECT 79.950 562.950 82.050 565.050 ;
        RECT 85.950 563.400 90.600 565.050 ;
        RECT 85.950 562.950 90.000 563.400 ;
        RECT 73.950 556.950 76.050 559.050 ;
        RECT 80.400 556.050 81.600 562.950 ;
        RECT 79.950 553.950 82.050 556.050 ;
        RECT 70.950 550.950 73.050 553.050 ;
        RECT 85.950 550.950 88.050 553.050 ;
        RECT 76.950 544.950 79.050 547.050 ;
        RECT 61.950 538.950 64.050 541.050 ;
        RECT 50.400 524.400 54.600 525.600 ;
        RECT 16.950 520.950 19.050 523.050 ;
        RECT 31.950 520.950 34.050 523.050 ;
        RECT 49.950 520.950 52.050 523.050 ;
        RECT 17.400 517.050 18.600 520.950 ;
        RECT 16.950 514.950 19.050 517.050 ;
        RECT 40.950 511.950 43.050 514.050 ;
        RECT 41.400 505.050 42.600 511.950 ;
        RECT 50.400 511.050 51.600 520.950 ;
        RECT 49.950 508.950 52.050 511.050 ;
        RECT 40.950 502.950 43.050 505.050 ;
        RECT 53.400 502.050 54.600 524.400 ;
        RECT 62.400 523.050 63.600 538.950 ;
        RECT 70.950 535.950 73.050 538.050 ;
        RECT 71.400 532.050 72.600 535.950 ;
        RECT 77.400 532.050 78.600 544.950 ;
        RECT 70.950 529.950 73.050 532.050 ;
        RECT 76.950 529.950 79.050 532.050 ;
        RECT 58.950 521.400 63.600 523.050 ;
        RECT 67.950 522.600 70.050 523.050 ;
        RECT 73.950 522.600 76.050 523.050 ;
        RECT 67.950 521.400 76.050 522.600 ;
        RECT 58.950 520.950 63.000 521.400 ;
        RECT 67.950 520.950 70.050 521.400 ;
        RECT 73.950 520.950 76.050 521.400 ;
        RECT 79.950 520.950 82.050 523.050 ;
        RECT 80.400 508.050 81.600 520.950 ;
        RECT 79.950 505.950 82.050 508.050 ;
        RECT 7.950 499.950 10.050 502.050 ;
        RECT 19.950 499.950 22.050 502.050 ;
        RECT 37.950 499.950 40.050 502.050 ;
        RECT 52.950 499.950 55.050 502.050 ;
        RECT 58.950 499.950 61.050 502.050 ;
        RECT 20.400 496.050 21.600 499.950 ;
        RECT 38.400 496.050 39.600 499.950 ;
        RECT 59.400 496.050 60.600 499.950 ;
        RECT 10.950 493.950 13.050 496.050 ;
        RECT 19.950 493.950 22.050 496.050 ;
        RECT 37.950 493.950 40.050 496.050 ;
        RECT 43.950 493.950 46.050 496.050 ;
        RECT 58.950 493.950 61.050 496.050 ;
        RECT 4.950 469.950 7.050 472.050 ;
        RECT 11.400 445.050 12.600 493.950 ;
        RECT 16.950 484.950 19.050 487.050 ;
        RECT 22.950 484.950 25.050 487.050 ;
        RECT 34.950 484.950 37.050 487.050 ;
        RECT 40.950 484.950 43.050 487.050 ;
        RECT 17.400 478.050 18.600 484.950 ;
        RECT 16.950 475.950 19.050 478.050 ;
        RECT 23.400 472.050 24.600 484.950 ;
        RECT 35.400 472.050 36.600 484.950 ;
        RECT 41.400 478.050 42.600 484.950 ;
        RECT 44.400 481.050 45.600 493.950 ;
        RECT 43.950 478.950 46.050 481.050 ;
        RECT 40.950 475.950 43.050 478.050 ;
        RECT 22.950 469.950 25.050 472.050 ;
        RECT 34.950 469.950 37.050 472.050 ;
        RECT 16.950 457.950 19.050 460.050 ;
        RECT 31.950 457.950 34.050 460.050 ;
        RECT 17.400 454.050 18.600 457.950 ;
        RECT 16.950 451.950 19.050 454.050 ;
        RECT 22.950 451.950 25.050 454.050 ;
        RECT 11.400 443.400 16.050 445.050 ;
        RECT 12.000 442.950 16.050 443.400 ;
        RECT 19.950 442.950 22.050 445.050 ;
        RECT 16.950 436.950 19.050 439.050 ;
        RECT 7.950 427.950 10.050 430.050 ;
        RECT 8.400 412.050 9.600 427.950 ;
        RECT 4.950 410.400 9.600 412.050 ;
        RECT 4.950 409.950 9.000 410.400 ;
        RECT 4.950 364.950 7.050 367.050 ;
        RECT 5.400 340.050 6.600 364.950 ;
        RECT 4.950 337.950 7.050 340.050 ;
        RECT 10.950 337.950 13.050 340.050 ;
        RECT 11.400 282.600 12.600 337.950 ;
        RECT 17.400 331.050 18.600 436.950 ;
        RECT 20.400 373.050 21.600 442.950 ;
        RECT 23.400 436.050 24.600 451.950 ;
        RECT 25.950 442.950 28.050 445.050 ;
        RECT 26.400 439.050 27.600 442.950 ;
        RECT 25.950 436.950 28.050 439.050 ;
        RECT 22.950 433.950 25.050 436.050 ;
        RECT 32.400 418.050 33.600 457.950 ;
        RECT 44.400 454.050 45.600 478.950 ;
        RECT 52.950 472.950 55.050 475.050 ;
        RECT 37.950 451.950 40.050 454.050 ;
        RECT 43.950 451.950 46.050 454.050 ;
        RECT 38.400 439.050 39.600 451.950 ;
        RECT 46.950 442.950 49.050 445.050 ;
        RECT 37.950 436.950 40.050 439.050 ;
        RECT 40.950 427.950 43.050 430.050 ;
        RECT 31.950 415.950 34.050 418.050 ;
        RECT 41.400 388.050 42.600 427.950 ;
        RECT 47.400 408.600 48.600 442.950 ;
        RECT 53.400 420.600 54.600 472.950 ;
        RECT 59.400 454.050 60.600 493.950 ;
        RECT 61.950 481.950 64.050 484.050 ;
        RECT 62.400 478.050 63.600 481.950 ;
        RECT 61.950 475.950 64.050 478.050 ;
        RECT 86.400 465.600 87.600 550.950 ;
        RECT 98.400 532.050 99.600 571.950 ;
        RECT 107.400 556.050 108.600 571.950 ;
        RECT 113.400 565.050 114.600 583.950 ;
        RECT 118.800 571.950 120.900 574.050 ;
        RECT 130.950 571.950 133.050 574.050 ;
        RECT 112.800 562.950 114.900 565.050 ;
        RECT 113.400 559.050 114.600 562.950 ;
        RECT 112.950 556.950 115.050 559.050 ;
        RECT 119.400 556.050 120.600 571.950 ;
        RECT 131.400 556.050 132.600 571.950 ;
        RECT 133.950 562.950 136.050 565.050 ;
        RECT 134.400 559.050 135.600 562.950 ;
        RECT 133.950 556.950 136.050 559.050 ;
        RECT 106.950 553.950 109.050 556.050 ;
        RECT 119.100 553.950 121.200 556.050 ;
        RECT 130.950 553.950 133.050 556.050 ;
        RECT 112.950 550.950 115.050 553.050 ;
        RECT 121.950 550.950 124.050 553.050 ;
        RECT 127.950 550.950 130.050 553.050 ;
        RECT 103.950 538.950 106.050 541.050 ;
        RECT 104.400 535.050 105.600 538.950 ;
        RECT 103.950 532.950 106.050 535.050 ;
        RECT 97.950 529.950 100.050 532.050 ;
        RECT 109.950 505.950 112.050 508.050 ;
        RECT 103.950 502.950 106.050 505.050 ;
        RECT 104.400 499.050 105.600 502.950 ;
        RECT 110.400 502.050 111.600 505.950 ;
        RECT 109.950 499.950 112.050 502.050 ;
        RECT 103.950 496.950 106.050 499.050 ;
        RECT 94.950 493.950 97.050 496.050 ;
        RECT 95.400 478.050 96.600 493.950 ;
        RECT 113.400 490.050 114.600 550.950 ;
        RECT 122.400 541.050 123.600 550.950 ;
        RECT 121.950 538.950 124.050 541.050 ;
        RECT 128.400 529.050 129.600 550.950 ;
        RECT 140.400 550.050 141.600 583.950 ;
        RECT 142.950 580.950 145.050 583.050 ;
        RECT 143.400 565.050 144.600 580.950 ;
        RECT 146.400 574.050 147.600 592.950 ;
        RECT 149.400 583.050 150.600 598.950 ;
        RECT 155.400 586.050 156.600 604.950 ;
        RECT 154.950 583.950 157.050 586.050 ;
        RECT 148.950 580.950 151.050 583.050 ;
        RECT 157.950 577.950 160.050 580.050 ;
        RECT 145.950 571.950 148.050 574.050 ;
        RECT 142.950 562.950 145.050 565.050 ;
        RECT 145.950 562.950 148.050 565.050 ;
        RECT 146.400 553.050 147.600 562.950 ;
        RECT 145.950 550.950 148.050 553.050 ;
        RECT 158.400 552.600 159.600 577.950 ;
        RECT 161.400 556.050 162.600 625.950 ;
        RECT 173.400 622.050 174.600 670.950 ;
        RECT 187.950 667.950 190.050 670.050 ;
        RECT 175.950 664.950 178.050 667.050 ;
        RECT 176.400 634.050 177.600 664.950 ;
        RECT 188.400 661.050 189.600 667.950 ;
        RECT 181.950 658.950 184.050 661.050 ;
        RECT 187.950 658.950 190.050 661.050 ;
        RECT 182.400 655.050 183.600 658.950 ;
        RECT 181.950 652.950 184.050 655.050 ;
        RECT 187.950 654.600 192.000 655.050 ;
        RECT 187.950 652.950 192.600 654.600 ;
        RECT 191.400 649.050 192.600 652.950 ;
        RECT 190.950 646.950 193.050 649.050 ;
        RECT 187.950 643.950 190.050 646.050 ;
        RECT 184.950 634.950 187.050 637.050 ;
        RECT 175.950 631.950 178.050 634.050 ;
        RECT 185.400 622.050 186.600 634.950 ;
        RECT 188.400 625.050 189.600 643.950 ;
        RECT 187.950 622.950 190.050 625.050 ;
        RECT 172.950 619.950 175.050 622.050 ;
        RECT 184.950 619.950 187.050 622.050 ;
        RECT 184.950 613.950 187.050 616.050 ;
        RECT 163.950 604.950 166.050 607.050 ;
        RECT 164.400 586.050 165.600 604.950 ;
        RECT 185.400 603.600 186.600 613.950 ;
        RECT 182.400 603.000 186.600 603.600 ;
        RECT 181.950 602.400 186.600 603.000 ;
        RECT 181.950 598.950 184.050 602.400 ;
        RECT 163.950 583.950 166.050 586.050 ;
        RECT 175.950 580.950 178.050 583.050 ;
        RECT 172.950 577.950 175.050 580.050 ;
        RECT 173.400 574.050 174.600 577.950 ;
        RECT 172.950 571.950 175.050 574.050 ;
        RECT 169.950 562.950 172.050 565.050 ;
        RECT 170.400 559.050 171.600 562.950 ;
        RECT 169.950 556.950 172.050 559.050 ;
        RECT 160.950 553.950 163.050 556.050 ;
        RECT 158.400 551.400 162.600 552.600 ;
        RECT 161.400 550.050 162.600 551.400 ;
        RECT 133.950 547.950 136.050 550.050 ;
        RECT 139.950 547.950 142.050 550.050 ;
        RECT 160.950 547.950 163.050 550.050 ;
        RECT 134.400 529.050 135.600 547.950 ;
        RECT 127.950 526.950 130.050 529.050 ;
        RECT 133.950 526.950 136.050 529.050 ;
        RECT 141.000 528.600 145.050 529.050 ;
        RECT 140.400 526.950 145.050 528.600 ;
        RECT 140.400 525.600 141.600 526.950 ;
        RECT 137.400 524.400 141.600 525.600 ;
        RECT 118.950 520.950 121.050 523.050 ;
        RECT 100.950 487.950 103.050 490.050 ;
        RECT 112.950 487.950 115.050 490.050 ;
        RECT 115.950 487.950 118.050 490.050 ;
        RECT 101.400 484.050 102.600 487.950 ;
        RECT 106.950 484.950 109.050 487.050 ;
        RECT 100.950 481.950 103.050 484.050 ;
        RECT 94.950 475.950 97.050 478.050 ;
        RECT 101.400 472.050 102.600 481.950 ;
        RECT 107.400 475.050 108.600 484.950 ;
        RECT 116.400 481.050 117.600 487.950 ;
        RECT 115.950 478.950 118.050 481.050 ;
        RECT 106.950 472.950 109.050 475.050 ;
        RECT 100.950 469.950 103.050 472.050 ;
        RECT 83.400 464.400 87.600 465.600 ;
        RECT 83.400 454.050 84.600 464.400 ;
        RECT 119.400 460.050 120.600 520.950 ;
        RECT 137.400 520.050 138.600 524.400 ;
        RECT 161.400 523.050 162.600 547.950 ;
        RECT 166.950 544.950 169.050 547.050 ;
        RECT 160.950 520.950 163.050 523.050 ;
        RECT 127.950 517.950 130.050 520.050 ;
        RECT 133.950 518.400 138.600 520.050 ;
        RECT 133.950 517.950 138.000 518.400 ;
        RECT 128.400 508.050 129.600 517.950 ;
        RECT 130.950 516.600 133.050 517.050 ;
        RECT 142.950 516.600 145.050 517.050 ;
        RECT 130.950 515.400 145.050 516.600 ;
        RECT 130.950 514.950 133.050 515.400 ;
        RECT 142.950 514.950 145.050 515.400 ;
        RECT 151.950 516.600 154.050 517.050 ;
        RECT 163.950 516.600 166.050 517.050 ;
        RECT 151.950 515.400 166.050 516.600 ;
        RECT 151.950 514.950 154.050 515.400 ;
        RECT 163.950 514.950 166.050 515.400 ;
        RECT 167.400 514.050 168.600 544.950 ;
        RECT 170.400 535.050 171.600 556.950 ;
        RECT 169.950 532.950 172.050 535.050 ;
        RECT 176.400 523.050 177.600 580.950 ;
        RECT 188.400 574.050 189.600 622.950 ;
        RECT 184.950 572.400 189.600 574.050 ;
        RECT 184.950 571.950 189.000 572.400 ;
        RECT 194.400 559.050 195.600 670.950 ;
        RECT 200.400 652.050 201.600 683.400 ;
        RECT 202.950 676.950 205.050 679.050 ;
        RECT 203.400 673.050 204.600 676.950 ;
        RECT 202.950 670.950 205.050 673.050 ;
        RECT 206.400 664.050 207.600 694.950 ;
        RECT 208.950 664.950 211.050 667.050 ;
        RECT 205.950 661.950 208.050 664.050 ;
        RECT 209.400 658.050 210.600 664.950 ;
        RECT 208.950 655.950 211.050 658.050 ;
        RECT 199.950 649.950 202.050 652.050 ;
        RECT 209.400 643.050 210.600 655.950 ;
        RECT 202.950 640.950 205.050 643.050 ;
        RECT 208.950 640.950 211.050 643.050 ;
        RECT 196.950 637.950 199.050 640.050 ;
        RECT 197.400 634.050 198.600 637.950 ;
        RECT 203.400 637.050 204.600 640.950 ;
        RECT 202.950 634.950 205.050 637.050 ;
        RECT 196.950 631.950 199.050 634.050 ;
        RECT 203.400 622.050 204.600 634.950 ;
        RECT 202.950 619.950 205.050 622.050 ;
        RECT 205.950 616.950 208.050 619.050 ;
        RECT 206.400 610.050 207.600 616.950 ;
        RECT 212.400 616.050 213.600 703.950 ;
        RECT 215.400 700.050 216.600 728.400 ;
        RECT 217.950 727.950 220.050 728.400 ;
        RECT 214.950 697.950 217.050 700.050 ;
        RECT 224.400 694.050 225.600 742.950 ;
        RECT 250.950 739.950 253.050 742.050 ;
        RECT 251.400 723.600 252.600 739.950 ;
        RECT 254.400 730.050 255.600 775.950 ;
        RECT 260.400 759.600 261.600 805.950 ;
        RECT 263.400 799.050 264.600 817.950 ;
        RECT 281.400 817.050 282.600 889.950 ;
        RECT 329.400 886.050 330.600 889.950 ;
        RECT 334.950 886.950 337.050 889.050 ;
        RECT 328.950 883.950 331.050 886.050 ;
        RECT 316.950 877.950 319.050 880.050 ;
        RECT 335.400 879.600 336.600 886.950 ;
        RECT 332.400 879.000 336.600 879.600 ;
        RECT 331.950 878.400 336.600 879.000 ;
        RECT 317.400 868.050 318.600 877.950 ;
        RECT 325.950 874.950 328.050 877.050 ;
        RECT 331.950 874.950 334.050 878.400 ;
        RECT 326.400 868.050 327.600 874.950 ;
        RECT 316.950 865.950 319.050 868.050 ;
        RECT 325.950 865.950 328.050 868.050 ;
        RECT 298.950 856.950 301.050 859.050 ;
        RECT 310.950 856.950 313.050 859.050 ;
        RECT 299.400 841.050 300.600 856.950 ;
        RECT 304.950 847.950 307.050 850.050 ;
        RECT 298.950 838.950 301.050 841.050 ;
        RECT 292.950 832.950 295.050 835.050 ;
        RECT 293.400 826.050 294.600 832.950 ;
        RECT 292.950 823.950 295.050 826.050 ;
        RECT 299.400 823.050 300.600 838.950 ;
        RECT 305.400 823.050 306.600 847.950 ;
        RECT 311.400 841.050 312.600 856.950 ;
        RECT 311.400 839.400 316.050 841.050 ;
        RECT 312.000 838.950 316.050 839.400 ;
        RECT 317.400 832.050 318.600 865.950 ;
        RECT 319.950 859.950 322.050 862.050 ;
        RECT 320.400 844.050 321.600 859.950 ;
        RECT 332.400 846.600 333.600 874.950 ;
        RECT 338.400 853.050 339.600 889.950 ;
        RECT 344.400 889.050 345.600 895.950 ;
        RECT 382.950 889.950 385.050 892.050 ;
        RECT 391.950 889.950 394.050 892.050 ;
        RECT 343.950 886.950 346.050 889.050 ;
        RECT 344.400 880.050 345.600 886.950 ;
        RECT 349.950 883.950 352.050 886.050 ;
        RECT 343.950 877.950 346.050 880.050 ;
        RECT 350.400 868.050 351.600 883.950 ;
        RECT 379.950 882.600 382.050 883.050 ;
        RECT 371.400 881.400 382.050 882.600 ;
        RECT 364.950 876.600 367.050 880.050 ;
        RECT 371.400 877.050 372.600 881.400 ;
        RECT 379.950 880.950 382.050 881.400 ;
        RECT 370.950 876.600 373.050 877.050 ;
        RECT 364.950 876.000 373.050 876.600 ;
        RECT 365.400 875.400 373.050 876.000 ;
        RECT 349.950 865.950 352.050 868.050 ;
        RECT 365.400 865.050 366.600 875.400 ;
        RECT 370.950 874.950 373.050 875.400 ;
        RECT 376.950 874.950 379.050 877.050 ;
        RECT 383.400 876.600 384.600 889.950 ;
        RECT 392.400 886.050 393.600 889.950 ;
        RECT 398.400 886.050 399.600 895.950 ;
        RECT 413.400 892.050 414.600 895.950 ;
        RECT 412.950 889.950 415.050 892.050 ;
        RECT 424.950 889.950 427.050 892.050 ;
        RECT 418.950 886.950 421.050 889.050 ;
        RECT 391.950 883.950 394.050 886.050 ;
        RECT 397.950 883.950 400.050 886.050 ;
        RECT 385.950 880.950 388.050 883.050 ;
        RECT 380.400 875.400 384.600 876.600 ;
        RECT 386.400 877.050 387.600 880.950 ;
        RECT 400.950 877.950 403.050 880.050 ;
        RECT 386.400 875.400 391.050 877.050 ;
        RECT 377.400 865.050 378.600 874.950 ;
        RECT 364.950 862.950 367.050 865.050 ;
        RECT 376.950 862.950 379.050 865.050 ;
        RECT 364.950 853.950 367.050 856.050 ;
        RECT 337.950 850.950 340.050 853.050 ;
        RECT 361.950 847.950 364.050 850.050 ;
        RECT 329.400 845.400 333.600 846.600 ;
        RECT 319.950 841.950 322.050 844.050 ;
        RECT 329.400 841.050 330.600 845.400 ;
        RECT 325.950 839.400 330.600 841.050 ;
        RECT 325.950 838.950 330.000 839.400 ;
        RECT 331.950 838.950 334.050 841.050 ;
        RECT 316.950 829.950 319.050 832.050 ;
        RECT 322.950 831.600 327.000 832.050 ;
        RECT 322.950 831.000 327.600 831.600 ;
        RECT 322.950 829.950 328.050 831.000 ;
        RECT 323.400 826.050 324.600 829.950 ;
        RECT 325.950 826.950 328.050 829.950 ;
        RECT 332.400 829.050 333.600 838.950 ;
        RECT 352.950 832.950 355.050 835.050 ;
        RECT 362.400 834.600 363.600 847.950 ;
        RECT 365.400 844.050 366.600 853.950 ;
        RECT 364.950 841.950 367.050 844.050 ;
        RECT 370.950 843.600 375.000 844.050 ;
        RECT 370.950 841.950 375.600 843.600 ;
        RECT 367.950 834.600 370.050 835.050 ;
        RECT 362.400 833.400 370.050 834.600 ;
        RECT 367.950 832.950 370.050 833.400 ;
        RECT 331.950 826.950 334.050 829.050 ;
        RECT 322.950 823.950 325.050 826.050 ;
        RECT 328.950 823.950 331.050 826.050 ;
        RECT 298.950 820.950 301.050 823.050 ;
        RECT 304.950 820.950 307.050 823.050 ;
        RECT 280.950 814.950 283.050 817.050 ;
        RECT 286.950 814.950 289.050 817.050 ;
        RECT 295.950 814.950 298.050 817.050 ;
        RECT 267.000 807.600 271.050 808.050 ;
        RECT 266.400 805.950 271.050 807.600 ;
        RECT 262.950 796.950 265.050 799.050 ;
        RECT 266.400 775.050 267.600 805.950 ;
        RECT 287.400 799.050 288.600 814.950 ;
        RECT 296.400 808.050 297.600 814.950 ;
        RECT 295.950 805.950 298.050 808.050 ;
        RECT 271.950 796.950 274.050 799.050 ;
        RECT 286.950 796.950 289.050 799.050 ;
        RECT 292.950 796.950 295.050 799.050 ;
        RECT 272.400 793.050 273.600 796.950 ;
        RECT 271.950 790.950 274.050 793.050 ;
        RECT 280.950 790.950 283.050 793.050 ;
        RECT 268.950 784.950 271.050 787.050 ;
        RECT 278.100 784.950 280.200 787.050 ;
        RECT 265.950 772.950 268.050 775.050 ;
        RECT 269.400 766.050 270.600 784.950 ;
        RECT 278.400 772.050 279.600 784.950 ;
        RECT 281.400 778.050 282.600 790.950 ;
        RECT 287.400 787.050 288.600 796.950 ;
        RECT 293.400 793.050 294.600 796.950 ;
        RECT 292.950 790.950 295.050 793.050 ;
        RECT 299.400 789.600 300.600 820.950 ;
        RECT 310.950 817.950 313.050 820.050 ;
        RECT 311.400 799.050 312.600 817.950 ;
        RECT 319.950 814.950 322.050 817.050 ;
        RECT 320.400 808.050 321.600 814.950 ;
        RECT 313.950 807.600 318.000 808.050 ;
        RECT 313.950 805.950 318.600 807.600 ;
        RECT 319.950 805.950 322.050 808.050 ;
        RECT 325.950 805.950 328.050 808.050 ;
        RECT 317.400 804.600 318.600 805.950 ;
        RECT 317.400 803.400 321.600 804.600 ;
        RECT 310.950 796.950 313.050 799.050 ;
        RECT 316.950 796.950 319.050 799.050 ;
        RECT 317.400 793.050 318.600 796.950 ;
        RECT 316.950 790.950 319.050 793.050 ;
        RECT 299.400 788.400 303.600 789.600 ;
        RECT 286.950 784.950 289.050 787.050 ;
        RECT 298.950 784.950 301.050 787.050 ;
        RECT 280.950 775.950 283.050 778.050 ;
        RECT 277.950 769.950 280.050 772.050 ;
        RECT 281.400 766.050 282.600 775.950 ;
        RECT 286.950 772.950 289.050 775.050 ;
        RECT 265.950 764.400 270.600 766.050 ;
        RECT 265.950 763.950 270.000 764.400 ;
        RECT 271.950 763.950 274.050 766.050 ;
        RECT 280.950 763.950 283.050 766.050 ;
        RECT 260.400 758.400 267.600 759.600 ;
        RECT 266.400 757.050 267.600 758.400 ;
        RECT 261.000 756.600 265.050 757.050 ;
        RECT 260.400 754.950 265.050 756.600 ;
        RECT 266.400 755.400 271.050 757.050 ;
        RECT 267.000 754.950 271.050 755.400 ;
        RECT 256.950 748.950 259.050 751.050 ;
        RECT 257.400 739.050 258.600 748.950 ;
        RECT 256.950 736.950 259.050 739.050 ;
        RECT 260.400 736.050 261.600 754.950 ;
        RECT 265.950 745.950 268.050 748.050 ;
        RECT 259.800 733.950 261.900 736.050 ;
        RECT 263.100 733.950 265.200 736.050 ;
        RECT 263.400 730.050 264.600 733.950 ;
        RECT 253.950 727.950 256.050 730.050 ;
        RECT 262.950 727.950 265.050 730.050 ;
        RECT 251.400 722.400 258.600 723.600 ;
        RECT 257.400 721.050 258.600 722.400 ;
        RECT 229.950 718.950 232.050 721.050 ;
        RECT 253.950 718.950 256.050 721.050 ;
        RECT 257.400 719.400 262.050 721.050 ;
        RECT 258.000 718.950 262.050 719.400 ;
        RECT 230.400 715.050 231.600 718.950 ;
        RECT 247.950 715.950 250.050 718.050 ;
        RECT 229.950 712.950 232.050 715.050 ;
        RECT 223.950 691.950 226.050 694.050 ;
        RECT 217.950 685.950 220.050 688.050 ;
        RECT 223.950 685.950 226.050 688.050 ;
        RECT 214.950 676.950 217.050 679.050 ;
        RECT 215.400 673.050 216.600 676.950 ;
        RECT 214.950 670.950 217.050 673.050 ;
        RECT 218.400 670.050 219.600 685.950 ;
        RECT 217.950 667.950 220.050 670.050 ;
        RECT 224.400 667.050 225.600 685.950 ;
        RECT 223.950 664.950 226.050 667.050 ;
        RECT 217.950 661.950 220.050 664.050 ;
        RECT 211.950 613.950 214.050 616.050 ;
        RECT 199.950 607.950 202.050 610.050 ;
        RECT 205.950 607.950 208.050 610.050 ;
        RECT 200.400 595.050 201.600 607.950 ;
        RECT 208.950 598.950 211.050 601.050 ;
        RECT 202.950 595.950 205.050 598.050 ;
        RECT 199.950 592.950 202.050 595.050 ;
        RECT 203.400 586.050 204.600 595.950 ;
        RECT 209.400 592.050 210.600 598.950 ;
        RECT 218.400 594.600 219.600 661.950 ;
        RECT 230.400 661.050 231.600 712.950 ;
        RECT 235.950 703.950 238.050 706.050 ;
        RECT 248.400 705.600 249.600 715.950 ;
        RECT 254.400 706.050 255.600 718.950 ;
        RECT 263.400 714.600 264.600 727.950 ;
        RECT 260.400 714.000 264.600 714.600 ;
        RECT 259.950 713.400 264.600 714.000 ;
        RECT 259.950 709.950 262.050 713.400 ;
        RECT 266.400 709.050 267.600 745.950 ;
        RECT 272.400 739.050 273.600 763.950 ;
        RECT 287.400 757.050 288.600 772.950 ;
        RECT 292.950 769.950 295.050 772.050 ;
        RECT 286.950 754.950 289.050 757.050 ;
        RECT 280.950 739.950 283.050 742.050 ;
        RECT 289.950 739.950 292.050 742.050 ;
        RECT 271.950 736.950 274.050 739.050 ;
        RECT 281.400 736.050 282.600 739.950 ;
        RECT 280.950 733.950 283.050 736.050 ;
        RECT 273.000 720.600 277.050 721.050 ;
        RECT 272.400 718.950 277.050 720.600 ;
        RECT 272.400 715.050 273.600 718.950 ;
        RECT 271.800 712.950 273.900 715.050 ;
        RECT 290.400 712.050 291.600 739.950 ;
        RECT 289.950 709.950 292.050 712.050 ;
        RECT 265.950 706.950 268.050 709.050 ;
        RECT 293.400 706.050 294.600 769.950 ;
        RECT 299.400 757.050 300.600 784.950 ;
        RECT 298.950 754.950 301.050 757.050 ;
        RECT 302.400 748.050 303.600 788.400 ;
        RECT 307.950 781.950 310.050 784.050 ;
        RECT 308.400 766.050 309.600 781.950 ;
        RECT 320.400 778.050 321.600 803.400 ;
        RECT 326.400 793.050 327.600 805.950 ;
        RECT 325.950 790.950 328.050 793.050 ;
        RECT 313.950 775.950 316.050 778.050 ;
        RECT 319.950 775.950 322.050 778.050 ;
        RECT 310.950 772.950 313.050 775.050 ;
        RECT 307.950 763.950 310.050 766.050 ;
        RECT 311.400 757.050 312.600 772.950 ;
        RECT 314.400 766.050 315.600 775.950 ;
        RECT 329.400 766.050 330.600 823.950 ;
        RECT 340.950 817.950 343.050 820.050 ;
        RECT 341.400 808.050 342.600 817.950 ;
        RECT 353.400 817.200 354.600 832.950 ;
        RECT 374.400 829.050 375.600 841.950 ;
        RECT 373.950 826.950 376.050 829.050 ;
        RECT 370.950 817.950 373.050 820.050 ;
        RECT 352.950 815.100 355.050 817.200 ;
        RECT 371.400 814.050 372.600 817.950 ;
        RECT 352.950 811.800 355.050 813.900 ;
        RECT 358.950 811.950 361.050 814.050 ;
        RECT 370.950 811.950 373.050 814.050 ;
        RECT 340.950 805.950 343.050 808.050 ;
        RECT 337.950 796.950 340.050 799.050 ;
        RECT 343.950 796.950 346.050 799.050 ;
        RECT 338.400 793.050 339.600 796.950 ;
        RECT 337.950 790.950 340.050 793.050 ;
        RECT 340.950 784.950 343.050 787.050 ;
        RECT 341.400 766.050 342.600 784.950 ;
        RECT 344.400 784.050 345.600 796.950 ;
        RECT 343.950 781.950 346.050 784.050 ;
        RECT 353.400 775.050 354.600 811.800 ;
        RECT 359.400 808.050 360.600 811.950 ;
        RECT 367.950 808.050 370.050 811.050 ;
        RECT 358.950 805.950 361.050 808.050 ;
        RECT 364.950 807.000 370.050 808.050 ;
        RECT 364.950 806.400 369.600 807.000 ;
        RECT 364.950 805.950 369.000 806.400 ;
        RECT 371.400 799.050 372.600 811.950 ;
        RECT 373.950 808.950 376.050 811.050 ;
        RECT 374.400 799.050 375.600 808.950 ;
        RECT 360.000 798.600 364.050 799.050 ;
        RECT 359.400 796.950 364.050 798.600 ;
        RECT 367.950 797.400 372.600 799.050 ;
        RECT 367.950 796.950 372.000 797.400 ;
        RECT 373.950 796.950 376.050 799.050 ;
        RECT 359.400 790.050 360.600 796.950 ;
        RECT 358.950 787.950 361.050 790.050 ;
        RECT 359.400 784.050 360.600 787.950 ;
        RECT 374.400 787.050 375.600 796.950 ;
        RECT 380.400 790.050 381.600 875.400 ;
        RECT 387.000 874.950 391.050 875.400 ;
        RECT 394.950 874.950 397.050 877.050 ;
        RECT 382.950 871.950 385.050 874.050 ;
        RECT 383.400 850.050 384.600 871.950 ;
        RECT 395.400 862.050 396.600 874.950 ;
        RECT 394.950 859.950 397.050 862.050 ;
        RECT 382.950 847.950 385.050 850.050 ;
        RECT 383.400 843.600 384.600 847.950 ;
        RECT 388.950 843.600 391.050 844.050 ;
        RECT 383.400 842.400 391.050 843.600 ;
        RECT 388.950 841.950 391.050 842.400 ;
        RECT 394.950 840.600 397.050 844.050 ;
        RECT 394.950 840.000 399.600 840.600 ;
        RECT 395.400 839.400 399.600 840.000 ;
        RECT 385.950 832.950 388.050 835.050 ;
        RECT 391.950 832.950 394.050 835.050 ;
        RECT 386.400 826.050 387.600 832.950 ;
        RECT 392.400 829.050 393.600 832.950 ;
        RECT 391.950 826.950 394.050 829.050 ;
        RECT 398.400 826.050 399.600 839.400 ;
        RECT 385.950 823.950 388.050 826.050 ;
        RECT 397.950 825.600 400.050 826.050 ;
        RECT 395.400 824.400 400.050 825.600 ;
        RECT 385.950 804.600 388.050 808.050 ;
        RECT 395.400 804.600 396.600 824.400 ;
        RECT 397.950 823.950 400.050 824.400 ;
        RECT 385.950 804.000 396.600 804.600 ;
        RECT 386.400 803.400 396.600 804.000 ;
        RECT 401.400 799.050 402.600 877.950 ;
        RECT 419.400 874.050 420.600 886.950 ;
        RECT 406.950 871.950 409.050 874.050 ;
        RECT 418.950 871.950 421.050 874.050 ;
        RECT 407.400 853.050 408.600 871.950 ;
        RECT 418.800 865.950 420.900 868.050 ;
        RECT 422.100 865.950 424.200 868.050 ;
        RECT 412.950 859.950 415.050 862.050 ;
        RECT 406.950 850.950 409.050 853.050 ;
        RECT 407.400 844.050 408.600 850.950 ;
        RECT 413.400 844.050 414.600 859.950 ;
        RECT 406.950 841.950 409.050 844.050 ;
        RECT 412.950 841.950 415.050 844.050 ;
        RECT 419.400 835.050 420.600 865.950 ;
        RECT 422.400 859.050 423.600 865.950 ;
        RECT 425.400 862.050 426.600 889.950 ;
        RECT 434.400 886.050 435.600 895.950 ;
        RECT 433.950 883.950 436.050 886.050 ;
        RECT 440.400 879.600 441.600 895.950 ;
        RECT 461.400 880.050 462.600 895.950 ;
        RECT 475.950 889.950 478.050 892.050 ;
        RECT 476.400 880.050 477.600 889.950 ;
        RECT 482.400 888.600 483.600 895.950 ;
        RECT 479.400 888.000 483.600 888.600 ;
        RECT 478.950 887.400 483.600 888.000 ;
        RECT 478.950 883.950 481.050 887.400 ;
        RECT 487.950 883.950 490.050 886.050 ;
        RECT 437.400 879.000 441.600 879.600 ;
        RECT 436.950 878.400 441.600 879.000 ;
        RECT 430.950 874.950 433.050 877.050 ;
        RECT 436.950 874.950 439.050 878.400 ;
        RECT 460.950 877.950 463.050 880.050 ;
        RECT 475.950 877.950 478.050 880.050 ;
        RECT 484.950 877.950 487.050 880.050 ;
        RECT 424.950 859.950 427.050 862.050 ;
        RECT 431.400 859.050 432.600 874.950 ;
        RECT 442.950 871.950 445.050 874.050 ;
        RECT 454.950 871.950 457.050 874.050 ;
        RECT 436.950 862.950 439.050 865.050 ;
        RECT 421.950 856.950 424.050 859.050 ;
        RECT 430.950 858.600 433.050 859.050 ;
        RECT 428.400 857.400 433.050 858.600 ;
        RECT 424.950 853.950 427.050 856.050 ;
        RECT 418.950 832.950 421.050 835.050 ;
        RECT 415.950 829.950 418.050 832.050 ;
        RECT 412.950 823.950 415.050 826.050 ;
        RECT 413.400 814.050 414.600 823.950 ;
        RECT 412.950 811.950 415.050 814.050 ;
        RECT 382.950 798.600 385.050 799.050 ;
        RECT 388.950 798.600 391.050 799.050 ;
        RECT 382.950 797.400 391.050 798.600 ;
        RECT 401.400 797.400 406.050 799.050 ;
        RECT 382.950 796.950 385.050 797.400 ;
        RECT 388.950 796.950 391.050 797.400 ;
        RECT 402.000 796.950 406.050 797.400 ;
        RECT 409.950 796.950 412.050 799.050 ;
        RECT 410.400 792.600 411.600 796.950 ;
        RECT 416.400 796.050 417.600 829.950 ;
        RECT 416.400 794.400 421.050 796.050 ;
        RECT 417.000 793.950 421.050 794.400 ;
        RECT 425.400 793.050 426.600 853.950 ;
        RECT 428.400 832.050 429.600 857.400 ;
        RECT 430.950 856.950 433.050 857.400 ;
        RECT 430.950 850.950 433.050 853.050 ;
        RECT 431.400 844.050 432.600 850.950 ;
        RECT 430.950 841.950 433.050 844.050 ;
        RECT 437.400 835.050 438.600 862.950 ;
        RECT 443.400 862.050 444.600 871.950 ;
        RECT 455.400 868.050 456.600 871.950 ;
        RECT 448.950 865.950 451.050 868.050 ;
        RECT 454.950 865.950 457.050 868.050 ;
        RECT 449.400 862.050 450.600 865.950 ;
        RECT 442.950 859.950 445.050 862.050 ;
        RECT 448.950 859.950 451.050 862.050 ;
        RECT 445.950 850.950 448.050 853.050 ;
        RECT 433.950 832.950 436.050 835.050 ;
        RECT 437.400 833.400 442.050 835.050 ;
        RECT 438.000 832.950 442.050 833.400 ;
        RECT 427.950 829.950 430.050 832.050 ;
        RECT 434.400 820.050 435.600 832.950 ;
        RECT 446.400 823.050 447.600 850.950 ;
        RECT 448.950 844.950 451.050 847.050 ;
        RECT 445.950 820.950 448.050 823.050 ;
        RECT 449.400 820.050 450.600 844.950 ;
        RECT 455.400 841.050 456.600 865.950 ;
        RECT 451.950 839.400 456.600 841.050 ;
        RECT 451.950 838.950 456.000 839.400 ;
        RECT 461.400 832.050 462.600 877.950 ;
        RECT 485.400 874.050 486.600 877.950 ;
        RECT 463.950 871.950 466.050 874.050 ;
        RECT 484.950 871.950 487.050 874.050 ;
        RECT 464.400 859.050 465.600 871.950 ;
        RECT 463.950 856.950 466.050 859.050 ;
        RECT 464.400 841.050 465.600 856.950 ;
        RECT 469.950 853.950 472.050 856.050 ;
        RECT 470.400 844.050 471.600 853.950 ;
        RECT 469.950 841.950 472.050 844.050 ;
        RECT 481.950 841.950 484.050 844.050 ;
        RECT 463.950 838.950 466.050 841.050 ;
        RECT 478.950 834.600 481.050 835.050 ;
        RECT 473.400 834.000 481.050 834.600 ;
        RECT 472.950 833.400 481.050 834.000 ;
        RECT 454.950 829.950 457.050 832.050 ;
        RECT 460.950 829.950 463.050 832.050 ;
        RECT 472.950 829.950 475.050 833.400 ;
        RECT 478.950 832.950 481.050 833.400 ;
        RECT 455.400 826.050 456.600 829.950 ;
        RECT 454.950 823.950 457.050 826.050 ;
        RECT 469.950 823.950 472.050 826.050 ;
        RECT 433.800 817.950 435.900 820.050 ;
        RECT 437.100 817.950 439.200 820.050 ;
        RECT 448.950 817.950 451.050 820.050 ;
        RECT 427.950 805.950 430.050 808.050 ;
        RECT 407.400 792.000 411.600 792.600 ;
        RECT 406.950 791.400 411.600 792.000 ;
        RECT 406.950 790.050 409.050 791.400 ;
        RECT 424.950 790.950 427.050 793.050 ;
        RECT 428.400 790.050 429.600 805.950 ;
        RECT 430.950 796.950 433.050 799.050 ;
        RECT 431.400 793.050 432.600 796.950 ;
        RECT 437.400 793.050 438.600 817.950 ;
        RECT 454.950 816.600 457.050 820.050 ;
        RECT 452.400 816.000 457.050 816.600 ;
        RECT 452.400 815.400 456.600 816.000 ;
        RECT 452.400 811.050 453.600 815.400 ;
        RECT 463.800 814.950 465.900 817.050 ;
        RECT 451.950 808.950 454.050 811.050 ;
        RECT 457.950 805.950 460.050 808.050 ;
        RECT 442.950 798.600 445.050 799.050 ;
        RECT 448.950 798.600 451.050 799.050 ;
        RECT 442.950 797.400 451.050 798.600 ;
        RECT 442.950 796.950 445.050 797.400 ;
        RECT 448.950 796.950 451.050 797.400 ;
        RECT 454.950 796.950 457.050 799.050 ;
        RECT 430.950 790.950 433.050 793.050 ;
        RECT 436.950 790.950 439.050 793.050 ;
        RECT 445.950 790.950 448.050 793.050 ;
        RECT 379.950 787.950 382.050 790.050 ;
        RECT 406.800 789.000 409.050 790.050 ;
        RECT 406.800 787.950 408.900 789.000 ;
        RECT 410.100 787.950 412.200 790.050 ;
        RECT 416.100 787.950 418.200 790.050 ;
        RECT 427.950 787.950 430.050 790.050 ;
        RECT 440.100 787.950 442.200 790.050 ;
        RECT 373.950 784.950 376.050 787.050 ;
        RECT 382.950 784.950 385.050 787.050 ;
        RECT 403.950 784.950 406.050 787.050 ;
        RECT 358.950 781.950 361.050 784.050 ;
        RECT 364.950 781.950 367.050 784.050 ;
        RECT 365.400 775.050 366.600 781.950 ;
        RECT 383.400 781.050 384.600 784.950 ;
        RECT 397.950 781.950 400.050 784.050 ;
        RECT 382.950 778.950 385.050 781.050 ;
        RECT 352.950 772.950 355.050 775.050 ;
        RECT 364.800 772.950 366.900 775.050 ;
        RECT 368.100 772.950 370.200 775.050 ;
        RECT 385.950 772.950 388.050 775.050 ;
        RECT 361.950 769.950 364.050 772.050 ;
        RECT 362.400 766.050 363.600 769.950 ;
        RECT 368.400 766.050 369.600 772.950 ;
        RECT 386.400 766.050 387.600 772.950 ;
        RECT 394.950 769.950 397.050 772.050 ;
        RECT 395.400 766.050 396.600 769.950 ;
        RECT 313.950 763.950 316.050 766.050 ;
        RECT 328.950 763.950 331.050 766.050 ;
        RECT 333.000 765.600 337.050 766.050 ;
        RECT 332.400 763.950 337.050 765.600 ;
        RECT 340.950 763.950 343.050 766.050 ;
        RECT 361.950 763.950 364.050 766.050 ;
        RECT 367.950 763.950 370.050 766.050 ;
        RECT 385.950 763.950 388.050 766.050 ;
        RECT 391.950 763.950 396.600 766.050 ;
        RECT 310.950 754.950 313.050 757.050 ;
        RECT 316.950 754.950 319.050 757.050 ;
        RECT 328.950 754.950 331.050 757.050 ;
        RECT 301.950 745.950 304.050 748.050 ;
        RECT 307.950 742.950 310.050 745.050 ;
        RECT 298.950 733.950 301.050 736.050 ;
        RECT 299.400 721.050 300.600 733.950 ;
        RECT 308.400 730.050 309.600 742.950 ;
        RECT 317.400 736.050 318.600 754.950 ;
        RECT 319.950 745.950 322.050 748.050 ;
        RECT 317.100 733.950 319.200 736.050 ;
        RECT 307.950 729.600 310.050 730.050 ;
        RECT 307.950 728.400 315.600 729.600 ;
        RECT 307.950 727.950 310.050 728.400 ;
        RECT 298.950 718.950 301.050 721.050 ;
        RECT 304.950 718.950 307.050 721.050 ;
        RECT 305.400 712.050 306.600 718.950 ;
        RECT 304.950 709.950 307.050 712.050 ;
        RECT 301.950 706.950 304.050 709.050 ;
        RECT 248.400 704.400 252.600 705.600 ;
        RECT 236.400 679.050 237.600 703.950 ;
        RECT 238.950 700.950 241.050 703.050 ;
        RECT 239.400 697.050 240.600 700.950 ;
        RECT 251.400 697.050 252.600 704.400 ;
        RECT 253.950 703.950 256.050 706.050 ;
        RECT 292.950 703.950 295.050 706.050 ;
        RECT 268.950 697.950 271.050 700.050 ;
        RECT 295.950 697.950 298.050 700.050 ;
        RECT 238.950 694.950 241.050 697.050 ;
        RECT 250.950 694.950 253.050 697.050 ;
        RECT 265.950 694.950 268.050 697.050 ;
        RECT 251.400 682.050 252.600 694.950 ;
        RECT 250.950 679.950 253.050 682.050 ;
        RECT 259.950 681.600 264.000 682.050 ;
        RECT 259.950 679.950 264.600 681.600 ;
        RECT 235.950 676.950 238.050 679.050 ;
        RECT 241.950 676.950 244.050 679.050 ;
        RECT 235.950 670.950 238.050 673.050 ;
        RECT 236.400 664.050 237.600 670.950 ;
        RECT 242.400 664.050 243.600 676.950 ;
        RECT 256.950 667.950 259.050 670.050 ;
        RECT 235.950 661.950 238.050 664.050 ;
        RECT 241.950 661.950 244.050 664.050 ;
        RECT 257.400 661.050 258.600 667.950 ;
        RECT 223.950 658.950 226.050 661.050 ;
        RECT 229.950 658.950 232.050 661.050 ;
        RECT 247.950 658.950 250.050 661.050 ;
        RECT 256.800 658.950 258.900 661.050 ;
        RECT 220.950 607.950 223.050 610.050 ;
        RECT 215.400 593.400 219.600 594.600 ;
        RECT 208.950 589.950 211.050 592.050 ;
        RECT 202.950 583.950 205.050 586.050 ;
        RECT 215.400 574.050 216.600 593.400 ;
        RECT 221.400 592.050 222.600 607.950 ;
        RECT 220.950 589.950 223.050 592.050 ;
        RECT 221.400 583.050 222.600 589.950 ;
        RECT 220.950 580.950 223.050 583.050 ;
        RECT 224.400 580.050 225.600 658.950 ;
        RECT 238.950 655.950 241.050 658.050 ;
        RECT 244.950 655.950 247.050 658.050 ;
        RECT 229.950 648.600 232.050 652.050 ;
        RECT 235.950 649.950 238.050 652.050 ;
        RECT 229.950 648.000 234.600 648.600 ;
        RECT 230.400 647.400 235.050 648.000 ;
        RECT 232.950 643.950 235.050 647.400 ;
        RECT 226.950 640.950 229.050 643.050 ;
        RECT 227.400 637.050 228.600 640.950 ;
        RECT 226.950 634.950 229.050 637.050 ;
        RECT 227.400 625.050 228.600 634.950 ;
        RECT 226.950 622.950 229.050 625.050 ;
        RECT 236.400 622.050 237.600 649.950 ;
        RECT 236.100 619.950 238.200 622.050 ;
        RECT 229.950 616.950 232.050 619.050 ;
        RECT 230.400 586.050 231.600 616.950 ;
        RECT 229.950 583.950 232.050 586.050 ;
        RECT 223.950 577.950 226.050 580.050 ;
        RECT 239.400 576.600 240.600 655.950 ;
        RECT 245.400 643.050 246.600 655.950 ;
        RECT 248.400 643.050 249.600 658.950 ;
        RECT 253.950 651.600 258.000 652.050 ;
        RECT 253.950 649.950 258.600 651.600 ;
        RECT 244.950 640.950 247.050 643.050 ;
        RECT 248.400 641.400 253.050 643.050 ;
        RECT 249.000 640.950 253.050 641.400 ;
        RECT 257.400 637.050 258.600 649.950 ;
        RECT 263.400 646.050 264.600 679.950 ;
        RECT 266.400 679.050 267.600 694.950 ;
        RECT 265.950 676.950 268.050 679.050 ;
        RECT 262.950 643.950 265.050 646.050 ;
        RECT 265.950 643.950 268.050 646.050 ;
        RECT 266.400 640.200 267.600 643.950 ;
        RECT 265.950 638.100 268.050 640.200 ;
        RECT 256.950 634.950 259.050 637.050 ;
        RECT 265.950 634.800 268.050 636.900 ;
        RECT 253.950 622.950 256.050 625.050 ;
        RECT 247.950 607.950 250.050 610.050 ;
        RECT 248.400 595.050 249.600 607.950 ;
        RECT 247.950 592.950 250.050 595.050 ;
        RECT 248.400 583.050 249.600 592.950 ;
        RECT 247.950 580.950 250.050 583.050 ;
        RECT 254.400 577.050 255.600 622.950 ;
        RECT 266.400 622.050 267.600 634.800 ;
        RECT 269.400 628.050 270.600 697.950 ;
        RECT 277.950 694.950 280.050 697.050 ;
        RECT 278.400 688.050 279.600 694.950 ;
        RECT 271.950 685.950 274.050 688.050 ;
        RECT 277.950 685.950 280.050 688.050 ;
        RECT 283.950 687.600 288.000 688.050 ;
        RECT 283.950 685.950 288.600 687.600 ;
        RECT 272.400 673.050 273.600 685.950 ;
        RECT 280.950 676.950 283.050 679.050 ;
        RECT 271.950 670.950 274.050 673.050 ;
        RECT 281.400 648.600 282.600 676.950 ;
        RECT 287.400 675.600 288.600 685.950 ;
        RECT 284.400 674.400 288.600 675.600 ;
        RECT 284.400 664.050 285.600 674.400 ;
        RECT 283.950 661.950 286.050 664.050 ;
        RECT 296.400 655.050 297.600 697.950 ;
        RECT 302.400 688.050 303.600 706.950 ;
        RECT 305.400 706.050 306.600 709.950 ;
        RECT 304.950 703.950 307.050 706.050 ;
        RECT 310.950 700.950 313.050 703.050 ;
        RECT 307.950 697.950 310.050 700.050 ;
        RECT 308.400 688.050 309.600 697.950 ;
        RECT 311.400 697.050 312.600 700.950 ;
        RECT 310.950 694.950 313.050 697.050 ;
        RECT 314.400 691.050 315.600 728.400 ;
        RECT 320.400 721.050 321.600 745.950 ;
        RECT 329.400 727.050 330.600 754.950 ;
        RECT 332.400 736.050 333.600 763.950 ;
        RECT 373.950 760.950 376.050 763.050 ;
        RECT 379.950 762.600 382.050 763.050 ;
        RECT 379.950 761.400 390.600 762.600 ;
        RECT 379.950 760.950 382.050 761.400 ;
        RECT 364.950 756.600 367.050 757.050 ;
        RECT 374.400 756.600 375.600 760.950 ;
        RECT 389.400 757.050 390.600 761.400 ;
        RECT 395.400 760.200 396.600 763.950 ;
        RECT 394.950 758.100 397.050 760.200 ;
        RECT 364.950 755.400 375.600 756.600 ;
        RECT 388.950 756.600 391.050 757.050 ;
        RECT 394.950 756.600 397.050 756.900 ;
        RECT 388.950 755.400 397.050 756.600 ;
        RECT 364.950 754.950 367.050 755.400 ;
        RECT 388.950 754.950 391.050 755.400 ;
        RECT 394.950 754.800 397.050 755.400 ;
        RECT 343.950 751.950 346.050 754.050 ;
        RECT 358.950 751.950 361.050 754.050 ;
        RECT 391.950 753.600 396.000 754.050 ;
        RECT 391.950 751.950 396.600 753.600 ;
        RECT 334.950 739.950 337.050 742.050 ;
        RECT 331.950 733.950 334.050 736.050 ;
        RECT 328.950 724.950 331.050 727.050 ;
        RECT 319.950 718.950 322.050 721.050 ;
        RECT 319.950 706.950 322.050 709.050 ;
        RECT 313.950 688.950 316.050 691.050 ;
        RECT 301.950 685.950 304.050 688.050 ;
        RECT 307.950 685.950 310.050 688.050 ;
        RECT 303.000 678.600 307.050 679.050 ;
        RECT 302.400 676.950 307.050 678.600 ;
        RECT 310.950 678.600 313.050 679.050 ;
        RECT 310.950 677.400 318.600 678.600 ;
        RECT 310.950 676.950 313.050 677.400 ;
        RECT 302.400 673.050 303.600 676.950 ;
        RECT 301.950 670.950 304.050 673.050 ;
        RECT 307.950 670.950 310.050 673.050 ;
        RECT 301.800 661.950 303.900 664.050 ;
        RECT 305.100 661.950 307.200 664.050 ;
        RECT 295.950 652.950 298.050 655.050 ;
        RECT 302.400 652.050 303.600 661.950 ;
        RECT 301.950 649.950 304.050 652.050 ;
        RECT 278.400 647.400 282.600 648.600 ;
        RECT 278.400 637.050 279.600 647.400 ;
        RECT 286.950 642.600 289.050 646.050 ;
        RECT 292.950 642.600 295.050 643.050 ;
        RECT 297.000 642.600 301.050 643.050 ;
        RECT 286.950 642.000 295.050 642.600 ;
        RECT 287.400 641.400 295.050 642.000 ;
        RECT 292.950 640.950 295.050 641.400 ;
        RECT 296.400 640.950 301.050 642.600 ;
        RECT 286.950 637.950 289.050 640.050 ;
        RECT 277.950 634.950 280.050 637.050 ;
        RECT 287.400 628.050 288.600 637.950 ;
        RECT 296.400 634.050 297.600 640.950 ;
        RECT 295.950 631.950 298.050 634.050 ;
        RECT 268.950 625.950 271.050 628.050 ;
        RECT 286.950 625.950 289.050 628.050 ;
        RECT 265.950 619.950 268.050 622.050 ;
        RECT 280.950 619.950 283.050 622.050 ;
        RECT 271.950 616.950 274.050 619.050 ;
        RECT 256.950 613.950 259.050 616.050 ;
        RECT 257.400 601.050 258.600 613.950 ;
        RECT 268.950 607.950 271.050 610.050 ;
        RECT 256.950 598.950 259.050 601.050 ;
        RECT 269.400 595.050 270.600 607.950 ;
        RECT 268.950 592.950 271.050 595.050 ;
        RECT 272.400 586.050 273.600 616.950 ;
        RECT 281.400 601.050 282.600 619.950 ;
        RECT 296.400 607.050 297.600 631.950 ;
        RECT 305.400 616.050 306.600 661.950 ;
        RECT 304.950 613.950 307.050 616.050 ;
        RECT 283.950 604.950 286.050 607.050 ;
        RECT 295.950 604.950 298.050 607.050 ;
        RECT 280.950 598.950 283.050 601.050 ;
        RECT 284.400 592.050 285.600 604.950 ;
        RECT 301.950 598.950 304.050 601.050 ;
        RECT 283.950 589.950 286.050 592.050 ;
        RECT 271.950 583.950 274.050 586.050 ;
        RECT 256.950 580.950 259.050 583.050 ;
        RECT 236.400 576.000 240.600 576.600 ;
        RECT 235.950 575.400 240.600 576.000 ;
        RECT 211.950 572.400 216.600 574.050 ;
        RECT 211.950 571.950 216.000 572.400 ;
        RECT 223.950 571.950 226.050 574.050 ;
        RECT 235.950 571.950 238.050 575.400 ;
        RECT 253.950 574.950 256.050 577.050 ;
        RECT 202.950 564.600 205.050 565.050 ;
        RECT 208.950 564.600 211.050 565.050 ;
        RECT 202.950 563.400 211.050 564.600 ;
        RECT 202.950 562.950 205.050 563.400 ;
        RECT 208.950 562.950 211.050 563.400 ;
        RECT 214.950 564.600 217.050 565.050 ;
        RECT 220.950 564.600 223.050 565.050 ;
        RECT 214.950 563.400 223.050 564.600 ;
        RECT 214.950 562.950 217.050 563.400 ;
        RECT 220.950 562.950 223.050 563.400 ;
        RECT 193.950 556.950 196.050 559.050 ;
        RECT 214.950 553.950 217.050 556.050 ;
        RECT 199.950 535.950 202.050 538.050 ;
        RECT 208.950 535.950 211.050 538.050 ;
        RECT 184.950 531.600 189.000 532.050 ;
        RECT 184.950 529.950 189.600 531.600 ;
        RECT 188.400 523.050 189.600 529.950 ;
        RECT 175.950 520.950 178.050 523.050 ;
        RECT 187.950 520.950 190.050 523.050 ;
        RECT 181.950 517.950 184.050 520.050 ;
        RECT 166.950 511.950 169.050 514.050 ;
        RECT 175.950 511.950 178.050 514.050 ;
        RECT 127.950 505.950 130.050 508.050 ;
        RECT 124.950 502.950 127.050 505.050 ;
        RECT 125.400 496.050 126.600 502.950 ;
        RECT 127.950 499.950 130.050 502.050 ;
        RECT 124.950 493.950 127.050 496.050 ;
        RECT 128.400 487.050 129.600 499.950 ;
        RECT 176.400 490.050 177.600 511.950 ;
        RECT 182.400 508.050 183.600 517.950 ;
        RECT 200.400 508.050 201.600 535.950 ;
        RECT 209.400 532.050 210.600 535.950 ;
        RECT 208.950 529.950 211.050 532.050 ;
        RECT 181.950 505.950 184.050 508.050 ;
        RECT 199.950 505.950 202.050 508.050 ;
        RECT 215.400 502.050 216.600 553.950 ;
        RECT 217.950 538.950 220.050 541.050 ;
        RECT 218.400 514.050 219.600 538.950 ;
        RECT 224.400 532.050 225.600 571.950 ;
        RECT 257.400 565.050 258.600 580.950 ;
        RECT 280.950 577.950 283.050 580.050 ;
        RECT 281.400 574.050 282.600 577.950 ;
        RECT 262.950 571.950 265.050 574.050 ;
        RECT 280.950 571.950 283.050 574.050 ;
        RECT 295.950 571.950 298.050 574.050 ;
        RECT 232.950 562.950 235.050 565.050 ;
        RECT 238.950 562.950 241.050 565.050 ;
        RECT 256.950 562.950 259.050 565.050 ;
        RECT 229.950 537.600 232.050 538.050 ;
        RECT 233.400 537.600 234.600 562.950 ;
        RECT 239.400 556.050 240.600 562.950 ;
        RECT 238.950 553.950 241.050 556.050 ;
        RECT 239.400 550.050 240.600 553.950 ;
        RECT 238.950 547.950 241.050 550.050 ;
        RECT 263.400 538.050 264.600 571.950 ;
        RECT 277.950 562.950 280.050 565.050 ;
        RECT 283.950 564.600 286.050 565.050 ;
        RECT 289.950 564.600 292.050 565.050 ;
        RECT 283.950 563.400 292.050 564.600 ;
        RECT 283.950 562.950 286.050 563.400 ;
        RECT 289.950 562.950 292.050 563.400 ;
        RECT 278.400 559.050 279.600 562.950 ;
        RECT 277.950 556.950 280.050 559.050 ;
        RECT 280.950 547.950 283.050 550.050 ;
        RECT 268.950 538.950 271.050 541.050 ;
        RECT 229.950 536.400 234.600 537.600 ;
        RECT 238.950 537.600 243.000 538.050 ;
        RECT 229.950 535.950 232.050 536.400 ;
        RECT 238.950 535.950 243.600 537.600 ;
        RECT 253.950 535.950 256.050 538.050 ;
        RECT 262.950 535.950 265.050 538.050 ;
        RECT 230.400 532.050 231.600 535.950 ;
        RECT 223.950 529.950 226.050 532.050 ;
        RECT 229.950 529.950 232.050 532.050 ;
        RECT 226.950 520.950 229.050 523.050 ;
        RECT 232.950 520.950 235.050 523.050 ;
        RECT 238.950 520.950 241.050 523.050 ;
        RECT 217.950 511.950 220.050 514.050 ;
        RECT 205.950 499.950 208.050 502.050 ;
        RECT 214.950 499.950 217.050 502.050 ;
        RECT 160.950 487.950 163.050 490.050 ;
        RECT 175.950 487.950 178.050 490.050 ;
        RECT 121.950 484.950 124.050 487.050 ;
        RECT 127.950 484.950 130.050 487.050 ;
        RECT 142.950 484.950 145.050 487.050 ;
        RECT 122.400 481.050 123.600 484.950 ;
        RECT 121.950 478.950 124.050 481.050 ;
        RECT 143.400 478.050 144.600 484.950 ;
        RECT 142.950 475.950 145.050 478.050 ;
        RECT 161.400 466.050 162.600 487.950 ;
        RECT 184.950 478.950 187.050 481.050 ;
        RECT 185.400 469.050 186.600 478.950 ;
        RECT 184.950 466.950 187.050 469.050 ;
        RECT 160.950 463.950 163.050 466.050 ;
        RECT 151.950 460.950 154.050 463.050 ;
        RECT 172.950 460.950 175.050 463.050 ;
        RECT 118.950 457.950 121.050 460.050 ;
        RECT 59.400 452.400 64.050 454.050 ;
        RECT 60.000 451.950 64.050 452.400 ;
        RECT 67.950 451.950 70.050 454.050 ;
        RECT 82.950 451.950 85.050 454.050 ;
        RECT 88.950 451.950 91.050 454.050 ;
        RECT 102.000 453.600 106.050 454.050 ;
        RECT 101.400 451.950 106.050 453.600 ;
        RECT 109.950 451.950 112.050 454.050 ;
        RECT 148.950 453.600 151.050 454.050 ;
        RECT 140.400 452.400 151.050 453.600 ;
        RECT 68.400 436.050 69.600 451.950 ;
        RECT 79.950 436.950 82.050 439.050 ;
        RECT 67.950 433.950 70.050 436.050 ;
        RECT 61.950 427.950 64.050 430.050 ;
        RECT 55.950 421.950 58.050 424.050 ;
        RECT 50.400 420.000 54.600 420.600 ;
        RECT 49.950 419.400 54.600 420.000 ;
        RECT 49.950 415.950 52.050 419.400 ;
        RECT 56.400 418.050 57.600 421.950 ;
        RECT 62.400 418.050 63.600 427.950 ;
        RECT 55.950 415.950 58.050 418.050 ;
        RECT 61.950 415.950 64.050 418.050 ;
        RECT 80.400 412.050 81.600 436.950 ;
        RECT 89.400 436.050 90.600 451.950 ;
        RECT 101.400 445.050 102.600 451.950 ;
        RECT 100.950 442.950 103.050 445.050 ;
        RECT 106.950 442.950 109.050 445.050 ;
        RECT 107.400 439.050 108.600 442.950 ;
        RECT 106.950 436.950 109.050 439.050 ;
        RECT 110.400 436.050 111.600 451.950 ;
        RECT 130.950 448.950 133.050 451.050 ;
        RECT 112.950 442.950 115.050 445.050 ;
        RECT 113.400 439.050 114.600 442.950 ;
        RECT 112.950 438.600 115.050 439.050 ;
        RECT 112.950 437.400 117.600 438.600 ;
        RECT 112.950 436.950 115.050 437.400 ;
        RECT 88.950 433.950 91.050 436.050 ;
        RECT 109.950 433.950 112.050 436.050 ;
        RECT 85.950 427.950 88.050 430.050 ;
        RECT 67.950 409.950 70.050 412.050 ;
        RECT 79.950 409.950 82.050 412.050 ;
        RECT 52.950 408.600 55.050 409.050 ;
        RECT 47.400 407.400 55.050 408.600 ;
        RECT 52.950 406.950 55.050 407.400 ;
        RECT 58.950 406.950 61.050 409.050 ;
        RECT 49.950 400.950 52.050 403.050 ;
        RECT 40.950 385.950 43.050 388.050 ;
        RECT 41.400 373.050 42.600 385.950 ;
        RECT 50.400 376.050 51.600 400.950 ;
        RECT 59.400 397.050 60.600 406.950 ;
        RECT 58.950 394.950 61.050 397.050 ;
        RECT 68.400 388.050 69.600 409.950 ;
        RECT 67.950 385.950 70.050 388.050 ;
        RECT 86.400 376.050 87.600 427.950 ;
        RECT 89.400 397.050 90.600 433.950 ;
        RECT 116.400 424.050 117.600 437.400 ;
        RECT 109.950 421.950 112.050 424.050 ;
        RECT 115.950 421.950 118.050 424.050 ;
        RECT 94.950 417.600 97.050 418.050 ;
        RECT 100.950 417.600 103.050 418.050 ;
        RECT 94.950 416.400 103.050 417.600 ;
        RECT 94.950 415.950 97.050 416.400 ;
        RECT 100.950 415.950 103.050 416.400 ;
        RECT 110.400 409.050 111.600 421.950 ;
        RECT 115.950 417.600 118.050 418.050 ;
        RECT 121.950 417.600 124.050 421.050 ;
        RECT 115.950 417.000 124.050 417.600 ;
        RECT 115.950 416.400 123.600 417.000 ;
        RECT 115.950 415.950 118.050 416.400 ;
        RECT 110.400 407.400 115.050 409.050 ;
        RECT 111.000 406.950 115.050 407.400 ;
        RECT 88.950 394.950 91.050 397.050 ;
        RECT 131.400 382.050 132.600 448.950 ;
        RECT 140.400 442.050 141.600 452.400 ;
        RECT 148.950 451.950 151.050 452.400 ;
        RECT 144.000 444.600 148.050 445.050 ;
        RECT 143.400 442.950 148.050 444.600 ;
        RECT 139.950 439.950 142.050 442.050 ;
        RECT 143.400 430.050 144.600 442.950 ;
        RECT 136.950 427.950 139.050 430.050 ;
        RECT 142.950 427.950 145.050 430.050 ;
        RECT 137.400 424.050 138.600 427.950 ;
        RECT 136.950 421.950 139.050 424.050 ;
        RECT 143.400 418.050 144.600 427.950 ;
        RECT 142.950 415.950 145.050 418.050 ;
        RECT 133.950 406.950 136.050 409.050 ;
        RECT 106.950 379.950 109.050 382.050 ;
        RECT 130.950 379.950 133.050 382.050 ;
        RECT 107.400 376.050 108.600 379.950 ;
        RECT 49.950 373.950 52.050 376.050 ;
        RECT 85.950 373.950 88.050 376.050 ;
        RECT 106.950 373.950 109.050 376.050 ;
        RECT 112.950 373.950 115.050 376.050 ;
        RECT 19.950 370.950 22.050 373.050 ;
        RECT 31.950 370.950 34.050 373.050 ;
        RECT 40.950 370.950 43.050 373.050 ;
        RECT 32.400 355.050 33.600 370.950 ;
        RECT 41.400 355.050 42.600 370.950 ;
        RECT 67.950 364.950 70.050 367.050 ;
        RECT 68.400 355.050 69.600 364.950 ;
        RECT 25.950 352.950 28.050 355.050 ;
        RECT 31.950 352.950 34.050 355.050 ;
        RECT 40.950 352.950 43.050 355.050 ;
        RECT 67.950 352.950 70.050 355.050 ;
        RECT 13.950 328.950 16.050 331.050 ;
        RECT 16.950 328.950 19.050 331.050 ;
        RECT 14.400 286.050 15.600 328.950 ;
        RECT 16.950 292.950 19.050 295.050 ;
        RECT 13.950 283.950 16.050 286.050 ;
        RECT 11.400 281.400 15.600 282.600 ;
        RECT 14.400 268.050 15.600 281.400 ;
        RECT 13.950 265.950 16.050 268.050 ;
        RECT 13.950 223.950 16.050 226.050 ;
        RECT 14.400 220.050 15.600 223.950 ;
        RECT 17.400 222.600 18.600 292.950 ;
        RECT 22.950 283.950 25.050 286.050 ;
        RECT 23.400 271.050 24.600 283.950 ;
        RECT 22.950 268.950 25.050 271.050 ;
        RECT 26.400 261.600 27.600 352.950 ;
        RECT 86.400 349.050 87.600 373.950 ;
        RECT 88.950 364.950 91.050 367.050 ;
        RECT 109.950 364.950 112.050 367.050 ;
        RECT 89.400 355.050 90.600 364.950 ;
        RECT 103.950 361.950 106.050 364.050 ;
        RECT 88.950 352.950 91.050 355.050 ;
        RECT 85.950 346.950 88.050 349.050 ;
        RECT 89.400 346.050 90.600 352.950 ;
        RECT 88.950 343.950 91.050 346.050 ;
        RECT 34.950 337.950 37.050 340.050 ;
        RECT 52.950 339.600 57.000 340.050 ;
        RECT 52.950 337.950 57.600 339.600 ;
        RECT 31.950 325.950 34.050 328.050 ;
        RECT 28.950 304.950 31.050 307.050 ;
        RECT 29.400 289.050 30.600 304.950 ;
        RECT 32.400 297.600 33.600 325.950 ;
        RECT 35.400 310.050 36.600 337.950 ;
        RECT 56.400 334.050 57.600 337.950 ;
        RECT 55.950 331.950 58.050 334.050 ;
        RECT 76.950 331.950 79.050 334.050 ;
        RECT 85.950 331.950 88.050 334.050 ;
        RECT 52.950 328.950 55.050 331.050 ;
        RECT 34.950 307.950 37.050 310.050 ;
        RECT 43.950 301.950 46.050 304.050 ;
        RECT 44.400 298.050 45.600 301.950 ;
        RECT 37.950 297.600 40.050 298.050 ;
        RECT 32.400 296.400 40.050 297.600 ;
        RECT 37.950 295.950 40.050 296.400 ;
        RECT 43.950 295.950 46.050 298.050 ;
        RECT 53.400 297.600 54.600 328.950 ;
        RECT 77.400 313.050 78.600 331.950 ;
        RECT 76.950 310.950 79.050 313.050 ;
        RECT 64.950 307.950 67.050 310.050 ;
        RECT 65.400 298.050 66.600 307.950 ;
        RECT 58.950 297.600 61.050 298.050 ;
        RECT 53.400 296.400 61.050 297.600 ;
        RECT 28.950 286.950 31.050 289.050 ;
        RECT 40.950 286.050 43.050 289.050 ;
        RECT 46.950 286.950 49.050 289.050 ;
        RECT 40.950 285.000 46.050 286.050 ;
        RECT 41.400 284.400 46.050 285.000 ;
        RECT 42.000 283.950 46.050 284.400 ;
        RECT 31.950 261.600 34.050 265.050 ;
        RECT 37.950 261.600 40.050 262.050 ;
        RECT 43.950 261.600 46.050 262.050 ;
        RECT 26.400 260.400 30.600 261.600 ;
        RECT 31.950 261.000 46.050 261.600 ;
        RECT 32.400 260.400 46.050 261.000 ;
        RECT 22.950 253.950 25.050 256.050 ;
        RECT 17.400 222.000 21.600 222.600 ;
        RECT 17.400 221.400 22.050 222.000 ;
        RECT 13.950 217.950 16.050 220.050 ;
        RECT 19.950 217.950 22.050 221.400 ;
        RECT 20.400 196.050 21.600 217.950 ;
        RECT 13.950 195.600 16.050 196.050 ;
        RECT 13.950 194.400 18.600 195.600 ;
        RECT 13.950 193.950 16.050 194.400 ;
        RECT 14.400 187.050 15.600 193.950 ;
        RECT 13.950 184.950 16.050 187.050 ;
        RECT 13.950 175.950 16.050 178.050 ;
        RECT 14.400 157.050 15.600 175.950 ;
        RECT 17.400 172.050 18.600 194.400 ;
        RECT 19.950 193.950 22.050 196.050 ;
        RECT 23.400 193.050 24.600 253.950 ;
        RECT 29.400 238.050 30.600 260.400 ;
        RECT 37.950 259.950 40.050 260.400 ;
        RECT 43.950 259.950 46.050 260.400 ;
        RECT 34.950 250.950 37.050 253.050 ;
        RECT 35.400 247.050 36.600 250.950 ;
        RECT 34.950 244.950 37.050 247.050 ;
        RECT 28.950 235.950 31.050 238.050 ;
        RECT 40.950 226.950 43.050 229.050 ;
        RECT 37.950 223.950 40.050 226.050 ;
        RECT 33.000 219.600 37.050 220.050 ;
        RECT 32.400 217.950 37.050 219.600 ;
        RECT 32.400 211.050 33.600 217.950 ;
        RECT 31.950 208.950 34.050 211.050 ;
        RECT 38.400 210.600 39.600 223.950 ;
        RECT 41.400 220.050 42.600 226.950 ;
        RECT 40.950 217.950 43.050 220.050 ;
        RECT 38.400 209.400 42.600 210.600 ;
        RECT 37.950 205.950 40.050 208.050 ;
        RECT 22.950 190.950 25.050 193.050 ;
        RECT 28.950 190.950 31.050 193.050 ;
        RECT 23.400 187.050 24.600 190.950 ;
        RECT 19.950 185.400 24.600 187.050 ;
        RECT 19.950 184.950 24.000 185.400 ;
        RECT 29.400 184.050 30.600 190.950 ;
        RECT 29.400 182.400 34.050 184.050 ;
        RECT 30.000 181.950 34.050 182.400 ;
        RECT 33.000 174.600 37.050 175.050 ;
        RECT 32.400 174.000 37.050 174.600 ;
        RECT 31.950 172.950 37.050 174.000 ;
        RECT 16.950 169.950 19.050 172.050 ;
        RECT 22.950 169.950 25.050 172.050 ;
        RECT 31.950 169.950 34.050 172.950 ;
        RECT 13.950 154.950 16.050 157.050 ;
        RECT 23.400 154.050 24.600 169.950 ;
        RECT 38.400 157.050 39.600 205.950 ;
        RECT 37.950 154.950 40.050 157.050 ;
        RECT 41.400 154.050 42.600 209.400 ;
        RECT 43.950 208.950 46.050 211.050 ;
        RECT 44.400 205.050 45.600 208.950 ;
        RECT 43.950 202.950 46.050 205.050 ;
        RECT 47.400 190.050 48.600 286.950 ;
        RECT 53.400 286.050 54.600 296.400 ;
        RECT 58.950 295.950 61.050 296.400 ;
        RECT 64.950 295.950 67.050 298.050 ;
        RECT 86.400 289.050 87.600 331.950 ;
        RECT 100.950 310.950 103.050 313.050 ;
        RECT 101.400 298.050 102.600 310.950 ;
        RECT 104.400 310.050 105.600 361.950 ;
        RECT 110.400 361.050 111.600 364.950 ;
        RECT 109.950 358.950 112.050 361.050 ;
        RECT 113.400 358.050 114.600 373.950 ;
        RECT 118.950 370.950 121.050 373.050 ;
        RECT 119.400 361.050 120.600 370.950 ;
        RECT 131.400 366.600 132.600 379.950 ;
        RECT 128.400 366.000 132.600 366.600 ;
        RECT 127.950 365.400 132.600 366.000 ;
        RECT 127.950 361.950 130.050 365.400 ;
        RECT 134.400 364.050 135.600 406.950 ;
        RECT 152.400 397.050 153.600 460.950 ;
        RECT 173.400 454.050 174.600 460.950 ;
        RECT 160.950 453.600 163.050 454.050 ;
        RECT 166.950 453.600 169.050 454.050 ;
        RECT 160.950 452.400 169.050 453.600 ;
        RECT 160.950 451.950 163.050 452.400 ;
        RECT 166.950 451.950 169.050 452.400 ;
        RECT 172.950 451.950 175.050 454.050 ;
        RECT 163.950 442.950 166.050 445.050 ;
        RECT 169.950 442.950 172.050 445.050 ;
        RECT 164.400 439.050 165.600 442.950 ;
        RECT 163.950 436.950 166.050 439.050 ;
        RECT 170.400 430.050 171.600 442.950 ;
        RECT 185.400 436.050 186.600 466.950 ;
        RECT 193.950 463.950 196.050 466.050 ;
        RECT 194.400 454.050 195.600 463.950 ;
        RECT 206.400 463.050 207.600 499.950 ;
        RECT 210.000 495.600 214.050 496.050 ;
        RECT 209.400 493.950 214.050 495.600 ;
        RECT 209.400 475.050 210.600 493.950 ;
        RECT 218.400 490.050 219.600 511.950 ;
        RECT 227.400 490.050 228.600 520.950 ;
        RECT 217.950 487.950 220.050 490.050 ;
        RECT 226.950 487.950 229.050 490.050 ;
        RECT 208.950 472.950 211.050 475.050 ;
        RECT 233.400 466.050 234.600 520.950 ;
        RECT 239.400 511.050 240.600 520.950 ;
        RECT 238.950 508.950 241.050 511.050 ;
        RECT 232.950 463.950 235.050 466.050 ;
        RECT 242.400 463.050 243.600 535.950 ;
        RECT 254.400 532.050 255.600 535.950 ;
        RECT 246.000 531.600 250.050 532.050 ;
        RECT 245.400 529.950 250.050 531.600 ;
        RECT 253.950 529.950 256.050 532.050 ;
        RECT 245.400 523.050 246.600 529.950 ;
        RECT 244.950 520.950 247.050 523.050 ;
        RECT 256.950 522.600 259.050 523.050 ;
        RECT 262.950 522.600 265.050 523.050 ;
        RECT 256.950 521.400 265.050 522.600 ;
        RECT 256.950 520.950 259.050 521.400 ;
        RECT 262.950 520.950 265.050 521.400 ;
        RECT 250.950 517.950 253.050 520.050 ;
        RECT 251.400 508.050 252.600 517.950 ;
        RECT 269.400 514.050 270.600 538.950 ;
        RECT 274.800 535.950 276.900 538.050 ;
        RECT 278.100 535.950 280.200 538.050 ;
        RECT 275.400 532.050 276.600 535.950 ;
        RECT 274.950 529.950 277.050 532.050 ;
        RECT 278.400 523.050 279.600 535.950 ;
        RECT 281.400 532.050 282.600 547.950 ;
        RECT 296.400 532.050 297.600 571.950 ;
        RECT 302.400 565.050 303.600 598.950 ;
        RECT 304.950 592.950 307.050 595.050 ;
        RECT 305.400 580.050 306.600 592.950 ;
        RECT 308.400 580.050 309.600 670.950 ;
        RECT 317.400 670.050 318.600 677.400 ;
        RECT 317.100 667.950 319.200 670.050 ;
        RECT 310.950 664.950 313.050 667.050 ;
        RECT 311.400 619.050 312.600 664.950 ;
        RECT 320.400 645.600 321.600 706.950 ;
        RECT 328.950 697.950 331.050 700.050 ;
        RECT 322.950 688.950 325.050 691.050 ;
        RECT 323.400 652.050 324.600 688.950 ;
        RECT 329.400 688.050 330.600 697.950 ;
        RECT 335.400 690.600 336.600 739.950 ;
        RECT 344.400 739.050 345.600 751.950 ;
        RECT 355.950 748.950 358.050 751.050 ;
        RECT 346.950 745.950 349.050 748.050 ;
        RECT 347.400 739.050 348.600 745.950 ;
        RECT 343.800 736.950 345.900 739.050 ;
        RECT 347.100 736.950 349.200 739.050 ;
        RECT 344.400 730.050 345.600 736.950 ;
        RECT 343.950 727.950 346.050 730.050 ;
        RECT 356.400 726.600 357.600 748.950 ;
        RECT 359.400 742.050 360.600 751.950 ;
        RECT 395.400 745.050 396.600 751.950 ;
        RECT 376.950 742.950 379.050 745.050 ;
        RECT 394.950 742.950 397.050 745.050 ;
        RECT 358.950 739.950 361.050 742.050 ;
        RECT 367.950 727.950 370.050 730.050 ;
        RECT 373.950 727.950 376.050 730.050 ;
        RECT 353.400 725.400 357.600 726.600 ;
        RECT 340.950 718.950 343.050 721.050 ;
        RECT 345.000 720.600 349.050 721.050 ;
        RECT 344.400 718.950 349.050 720.600 ;
        RECT 337.950 706.950 340.050 709.050 ;
        RECT 332.400 689.400 336.600 690.600 ;
        RECT 328.950 685.950 331.050 688.050 ;
        RECT 325.950 673.950 328.050 676.050 ;
        RECT 326.400 658.050 327.600 673.950 ;
        RECT 332.400 669.600 333.600 689.400 ;
        RECT 334.950 685.950 337.050 688.050 ;
        RECT 335.400 670.050 336.600 685.950 ;
        RECT 338.400 682.050 339.600 706.950 ;
        RECT 341.400 697.050 342.600 718.950 ;
        RECT 341.100 694.950 343.200 697.050 ;
        RECT 341.400 688.050 342.600 694.950 ;
        RECT 344.400 691.050 345.600 718.950 ;
        RECT 353.400 718.050 354.600 725.400 ;
        RECT 361.950 723.600 364.050 724.050 ;
        RECT 356.400 723.000 364.050 723.600 ;
        RECT 355.950 722.400 364.050 723.000 ;
        RECT 355.950 718.950 358.050 722.400 ;
        RECT 361.950 721.950 364.050 722.400 ;
        RECT 368.400 718.050 369.600 727.950 ;
        RECT 374.400 724.050 375.600 727.950 ;
        RECT 370.950 722.400 375.600 724.050 ;
        RECT 370.950 721.950 375.000 722.400 ;
        RECT 352.950 715.950 355.050 718.050 ;
        RECT 361.950 715.950 364.050 718.050 ;
        RECT 367.950 715.950 370.050 718.050 ;
        RECT 373.950 715.950 376.050 718.050 ;
        RECT 349.950 709.950 352.050 712.050 ;
        RECT 343.950 688.950 346.050 691.050 ;
        RECT 350.400 690.600 351.600 709.950 ;
        RECT 355.950 706.950 358.050 709.050 ;
        RECT 356.400 694.050 357.600 706.950 ;
        RECT 362.400 703.200 363.600 715.950 ;
        RECT 358.800 700.950 360.900 703.050 ;
        RECT 362.100 701.100 364.200 703.200 ;
        RECT 355.950 691.950 358.050 694.050 ;
        RECT 350.400 689.400 354.600 690.600 ;
        RECT 340.950 685.950 343.050 688.050 ;
        RECT 349.950 685.950 352.050 688.050 ;
        RECT 337.950 679.950 340.050 682.050 ;
        RECT 346.950 679.950 349.050 682.050 ;
        RECT 340.950 670.950 343.050 673.050 ;
        RECT 329.400 668.400 333.600 669.600 ;
        RECT 325.800 655.950 327.900 658.050 ;
        RECT 322.950 651.600 327.000 652.050 ;
        RECT 322.950 649.950 327.600 651.600 ;
        RECT 326.400 646.050 327.600 649.950 ;
        RECT 317.400 644.400 321.600 645.600 ;
        RECT 313.950 640.950 316.050 643.050 ;
        RECT 314.400 637.050 315.600 640.950 ;
        RECT 313.950 634.950 316.050 637.050 ;
        RECT 317.400 621.600 318.600 644.400 ;
        RECT 325.950 643.950 328.050 646.050 ;
        RECT 319.950 640.050 322.050 643.050 ;
        RECT 319.950 639.000 325.050 640.050 ;
        RECT 320.400 638.400 325.050 639.000 ;
        RECT 321.000 637.950 325.050 638.400 ;
        RECT 322.950 631.950 325.050 634.050 ;
        RECT 323.400 628.050 324.600 631.950 ;
        RECT 322.950 625.950 325.050 628.050 ;
        RECT 317.400 620.400 321.600 621.600 ;
        RECT 310.800 616.950 312.900 619.050 ;
        RECT 314.100 616.950 316.200 619.050 ;
        RECT 314.400 610.050 315.600 616.950 ;
        RECT 320.400 616.050 321.600 620.400 ;
        RECT 329.400 616.050 330.600 668.400 ;
        RECT 334.950 667.950 337.050 670.050 ;
        RECT 331.950 664.950 334.050 667.050 ;
        RECT 332.400 652.050 333.600 664.950 ;
        RECT 332.400 650.400 337.050 652.050 ;
        RECT 333.000 649.950 337.050 650.400 ;
        RECT 341.400 643.050 342.600 670.950 ;
        RECT 343.950 667.950 346.050 670.050 ;
        RECT 344.400 643.050 345.600 667.950 ;
        RECT 337.950 641.400 342.600 643.050 ;
        RECT 337.950 640.950 342.000 641.400 ;
        RECT 343.950 640.950 346.050 643.050 ;
        RECT 347.400 628.050 348.600 679.950 ;
        RECT 350.400 661.050 351.600 685.950 ;
        RECT 353.400 673.050 354.600 689.400 ;
        RECT 359.400 679.050 360.600 700.950 ;
        RECT 370.950 697.950 373.050 700.050 ;
        RECT 371.400 688.050 372.600 697.950 ;
        RECT 374.400 697.050 375.600 715.950 ;
        RECT 377.400 700.050 378.600 742.950 ;
        RECT 385.950 739.950 388.050 742.050 ;
        RECT 386.400 733.050 387.600 739.950 ;
        RECT 398.400 739.050 399.600 781.950 ;
        RECT 400.950 772.950 403.050 775.050 ;
        RECT 401.400 748.050 402.600 772.950 ;
        RECT 400.950 745.950 403.050 748.050 ;
        RECT 397.950 736.950 400.050 739.050 ;
        RECT 385.950 730.950 388.050 733.050 ;
        RECT 379.950 724.950 382.050 727.050 ;
        RECT 376.950 697.950 379.050 700.050 ;
        RECT 380.400 697.050 381.600 724.950 ;
        RECT 386.400 721.050 387.600 730.950 ;
        RECT 388.950 729.600 393.000 730.050 ;
        RECT 394.950 729.600 397.050 730.050 ;
        RECT 388.950 727.950 393.600 729.600 ;
        RECT 394.950 728.400 402.600 729.600 ;
        RECT 394.950 727.950 397.050 728.400 ;
        RECT 392.400 726.600 393.600 727.950 ;
        RECT 392.400 725.400 399.600 726.600 ;
        RECT 398.400 721.050 399.600 725.400 ;
        RECT 385.950 718.950 388.050 721.050 ;
        RECT 391.950 718.950 394.050 721.050 ;
        RECT 397.950 718.950 400.050 721.050 ;
        RECT 392.400 715.050 393.600 718.950 ;
        RECT 401.400 717.600 402.600 728.400 ;
        RECT 398.400 716.400 402.600 717.600 ;
        RECT 391.950 712.950 394.050 715.050 ;
        RECT 391.950 706.950 394.050 709.050 ;
        RECT 388.950 700.950 391.050 703.050 ;
        RECT 373.950 694.950 376.050 697.050 ;
        RECT 379.950 694.950 382.050 697.050 ;
        RECT 370.950 685.950 373.050 688.050 ;
        RECT 358.950 676.950 361.050 679.050 ;
        RECT 389.400 678.600 390.600 700.950 ;
        RECT 392.400 691.050 393.600 706.950 ;
        RECT 398.400 706.050 399.600 716.400 ;
        RECT 404.400 706.050 405.600 784.950 ;
        RECT 406.950 775.950 409.050 778.050 ;
        RECT 407.400 748.050 408.600 775.950 ;
        RECT 410.400 772.050 411.600 787.950 ;
        RECT 416.400 781.050 417.600 787.950 ;
        RECT 424.950 784.950 427.050 787.050 ;
        RECT 415.800 778.950 417.900 781.050 ;
        RECT 419.100 778.950 421.200 781.050 ;
        RECT 409.950 769.950 412.050 772.050 ;
        RECT 410.400 766.050 411.600 769.950 ;
        RECT 419.400 766.050 420.600 778.950 ;
        RECT 409.950 763.950 412.050 766.050 ;
        RECT 415.950 764.400 420.600 766.050 ;
        RECT 415.950 763.950 420.000 764.400 ;
        RECT 412.950 756.600 417.000 757.050 ;
        RECT 425.400 756.600 426.600 784.950 ;
        RECT 428.400 766.050 429.600 787.950 ;
        RECT 440.400 778.050 441.600 787.950 ;
        RECT 442.950 781.950 445.050 784.050 ;
        RECT 443.400 778.050 444.600 781.950 ;
        RECT 433.950 775.950 436.050 778.050 ;
        RECT 439.800 775.950 441.900 778.050 ;
        RECT 443.100 775.950 445.200 778.050 ;
        RECT 434.400 766.050 435.600 775.950 ;
        RECT 446.400 769.050 447.600 790.950 ;
        RECT 449.400 787.050 450.600 796.950 ;
        RECT 455.400 793.050 456.600 796.950 ;
        RECT 454.950 790.950 457.050 793.050 ;
        RECT 448.950 784.950 451.050 787.050 ;
        RECT 458.400 784.050 459.600 805.950 ;
        RECT 457.950 781.950 460.050 784.050 ;
        RECT 448.950 778.950 451.050 781.050 ;
        RECT 445.950 766.950 448.050 769.050 ;
        RECT 427.950 763.950 430.050 766.050 ;
        RECT 433.950 763.950 436.050 766.050 ;
        RECT 449.400 757.050 450.600 778.950 ;
        RECT 460.950 769.950 463.050 772.050 ;
        RECT 451.950 766.050 454.050 769.050 ;
        RECT 461.400 766.050 462.600 769.950 ;
        RECT 451.950 765.000 457.050 766.050 ;
        RECT 452.400 764.400 457.050 765.000 ;
        RECT 453.000 763.950 457.050 764.400 ;
        RECT 460.950 763.950 463.050 766.050 ;
        RECT 464.400 757.050 465.600 814.950 ;
        RECT 466.950 793.950 469.050 796.050 ;
        RECT 467.400 760.050 468.600 793.950 ;
        RECT 470.400 790.050 471.600 823.950 ;
        RECT 482.400 823.050 483.600 841.950 ;
        RECT 472.950 820.950 475.050 823.050 ;
        RECT 481.950 820.950 484.050 823.050 ;
        RECT 473.400 817.050 474.600 820.950 ;
        RECT 478.950 817.950 481.050 820.050 ;
        RECT 472.950 814.950 475.050 817.050 ;
        RECT 475.950 811.950 478.050 814.050 ;
        RECT 476.400 799.050 477.600 811.950 ;
        RECT 479.400 808.050 480.600 817.950 ;
        RECT 481.950 808.950 484.050 811.050 ;
        RECT 478.950 805.950 481.050 808.050 ;
        RECT 482.400 799.050 483.600 808.950 ;
        RECT 475.950 796.950 478.050 799.050 ;
        RECT 481.950 796.950 484.050 799.050 ;
        RECT 488.400 793.050 489.600 883.950 ;
        RECT 490.950 871.950 493.050 874.050 ;
        RECT 491.400 862.200 492.600 871.950 ;
        RECT 497.400 867.600 498.600 895.950 ;
        RECT 524.400 889.050 525.600 895.950 ;
        RECT 551.400 892.050 552.600 898.950 ;
        RECT 562.950 895.950 565.050 898.050 ;
        RECT 574.950 895.950 577.050 898.050 ;
        RECT 550.950 889.950 553.050 892.050 ;
        RECT 523.950 886.950 526.050 889.050 ;
        RECT 531.000 888.600 535.050 889.050 ;
        RECT 530.400 888.000 535.050 888.600 ;
        RECT 529.950 886.950 535.050 888.000 ;
        RECT 541.950 888.600 544.050 889.050 ;
        RECT 541.950 888.000 555.600 888.600 ;
        RECT 541.950 887.400 556.050 888.000 ;
        RECT 541.950 886.950 544.050 887.400 ;
        RECT 505.950 885.600 508.050 886.050 ;
        RECT 511.950 885.600 514.050 886.050 ;
        RECT 505.950 884.400 514.050 885.600 ;
        RECT 505.950 883.950 508.050 884.400 ;
        RECT 511.950 883.950 514.050 884.400 ;
        RECT 517.950 885.600 520.050 886.050 ;
        RECT 529.950 885.600 532.050 886.950 ;
        RECT 517.950 884.400 532.050 885.600 ;
        RECT 517.950 883.950 520.050 884.400 ;
        RECT 529.950 883.950 532.050 884.400 ;
        RECT 535.950 883.950 538.050 886.050 ;
        RECT 553.950 883.950 556.050 887.400 ;
        RECT 506.400 878.400 519.600 879.600 ;
        RECT 506.400 877.050 507.600 878.400 ;
        RECT 502.950 875.400 507.600 877.050 ;
        RECT 502.950 874.950 507.000 875.400 ;
        RECT 508.950 874.950 511.050 877.050 ;
        RECT 509.400 868.050 510.600 874.950 ;
        RECT 514.950 871.950 517.050 874.050 ;
        RECT 494.400 866.400 498.600 867.600 ;
        RECT 490.950 860.100 493.050 862.200 ;
        RECT 490.950 856.800 493.050 858.900 ;
        RECT 491.400 843.600 492.600 856.800 ;
        RECT 494.400 856.050 495.600 866.400 ;
        RECT 508.950 865.950 511.050 868.050 ;
        RECT 496.950 862.950 499.050 865.050 ;
        RECT 497.400 859.050 498.600 862.950 ;
        RECT 496.950 856.950 499.050 859.050 ;
        RECT 493.950 853.950 496.050 856.050 ;
        RECT 515.400 853.050 516.600 871.950 ;
        RECT 508.950 850.950 511.050 853.050 ;
        RECT 514.950 850.950 517.050 853.050 ;
        RECT 496.950 843.600 499.050 844.050 ;
        RECT 491.400 842.400 499.050 843.600 ;
        RECT 487.950 790.950 490.050 793.050 ;
        RECT 469.950 787.950 472.050 790.050 ;
        RECT 470.400 765.600 471.600 787.950 ;
        RECT 491.400 787.050 492.600 842.400 ;
        RECT 496.950 841.950 499.050 842.400 ;
        RECT 499.950 832.950 502.050 835.050 ;
        RECT 505.950 832.950 508.050 835.050 ;
        RECT 500.400 829.050 501.600 832.950 ;
        RECT 499.950 826.950 502.050 829.050 ;
        RECT 506.400 828.600 507.600 832.950 ;
        RECT 503.400 827.400 507.600 828.600 ;
        RECT 493.950 820.950 496.050 823.050 ;
        RECT 494.400 814.200 495.600 820.950 ;
        RECT 499.950 817.950 502.050 820.050 ;
        RECT 493.950 812.100 496.050 814.200 ;
        RECT 500.400 811.050 501.600 817.950 ;
        RECT 493.950 808.800 496.050 810.900 ;
        RECT 499.950 808.950 502.050 811.050 ;
        RECT 494.400 802.050 495.600 808.800 ;
        RECT 493.950 799.950 496.050 802.050 ;
        RECT 496.950 799.950 499.050 802.050 ;
        RECT 503.400 801.600 504.600 827.400 ;
        RECT 505.950 823.950 508.050 826.050 ;
        RECT 506.400 811.050 507.600 823.950 ;
        RECT 505.950 808.950 508.050 811.050 ;
        RECT 509.400 802.050 510.600 850.950 ;
        RECT 518.400 817.050 519.600 878.400 ;
        RECT 536.400 877.050 537.600 883.950 ;
        RECT 526.950 874.950 529.050 877.050 ;
        RECT 532.950 875.400 537.600 877.050 ;
        RECT 532.950 874.950 537.000 875.400 ;
        RECT 527.400 868.050 528.600 874.950 ;
        RECT 526.950 865.950 529.050 868.050 ;
        RECT 523.950 841.950 526.050 844.050 ;
        RECT 529.950 841.950 532.050 844.050 ;
        RECT 524.400 829.050 525.600 841.950 ;
        RECT 523.950 826.950 526.050 829.050 ;
        RECT 524.400 820.050 525.600 826.950 ;
        RECT 530.400 823.050 531.600 841.950 ;
        RECT 533.400 829.050 534.600 874.950 ;
        RECT 539.100 862.950 541.200 865.050 ;
        RECT 533.400 826.950 538.200 829.050 ;
        RECT 529.950 822.600 532.050 823.050 ;
        RECT 527.400 821.400 532.050 822.600 ;
        RECT 523.950 817.950 526.050 820.050 ;
        RECT 511.950 813.600 514.050 817.050 ;
        RECT 517.950 814.950 520.050 817.050 ;
        RECT 511.950 813.000 516.600 813.600 ;
        RECT 512.400 812.400 516.600 813.000 ;
        RECT 500.400 800.400 504.600 801.600 ;
        RECT 497.400 796.200 498.600 799.950 ;
        RECT 496.950 794.100 499.050 796.200 ;
        RECT 496.950 790.800 499.050 792.900 ;
        RECT 478.950 784.950 481.050 787.050 ;
        RECT 484.950 784.950 487.050 787.050 ;
        RECT 490.950 784.950 493.050 787.050 ;
        RECT 479.400 768.600 480.600 784.950 ;
        RECT 485.400 772.050 486.600 784.950 ;
        RECT 497.400 772.050 498.600 790.800 ;
        RECT 500.400 784.050 501.600 800.400 ;
        RECT 508.950 799.950 511.050 802.050 ;
        RECT 502.950 796.950 505.050 799.050 ;
        RECT 503.400 784.050 504.600 796.950 ;
        RECT 505.950 784.950 508.050 787.050 ;
        RECT 499.800 781.950 501.900 784.050 ;
        RECT 503.100 781.950 505.200 784.050 ;
        RECT 506.400 772.050 507.600 784.950 ;
        RECT 484.950 769.950 487.050 772.050 ;
        RECT 496.950 769.950 499.050 772.050 ;
        RECT 502.800 769.950 504.900 772.050 ;
        RECT 506.100 769.950 508.200 772.050 ;
        RECT 479.400 768.000 483.600 768.600 ;
        RECT 479.400 767.400 484.050 768.000 ;
        RECT 475.950 765.600 478.050 766.050 ;
        RECT 470.400 764.400 478.050 765.600 ;
        RECT 475.950 763.950 478.050 764.400 ;
        RECT 481.950 763.950 484.050 767.400 ;
        RECT 503.400 766.050 504.600 769.950 ;
        RECT 515.400 769.050 516.600 812.400 ;
        RECT 527.400 801.600 528.600 821.400 ;
        RECT 529.950 820.950 532.050 821.400 ;
        RECT 533.400 817.050 534.600 826.950 ;
        RECT 539.400 820.050 540.600 862.950 ;
        RECT 544.950 859.950 547.050 862.050 ;
        RECT 545.400 850.050 546.600 859.950 ;
        RECT 563.400 856.050 564.600 895.950 ;
        RECT 575.400 886.050 576.600 895.950 ;
        RECT 574.950 883.950 577.050 886.050 ;
        RECT 580.950 885.600 583.050 886.050 ;
        RECT 580.950 884.400 585.600 885.600 ;
        RECT 580.950 883.950 583.050 884.400 ;
        RECT 571.950 876.600 574.050 877.050 ;
        RECT 581.400 876.600 582.600 883.950 ;
        RECT 571.950 875.400 582.600 876.600 ;
        RECT 571.950 874.950 574.050 875.400 ;
        RECT 568.950 856.950 571.050 859.050 ;
        RECT 580.950 856.950 583.050 859.050 ;
        RECT 557.100 853.950 559.200 856.050 ;
        RECT 562.950 853.950 565.050 856.050 ;
        RECT 550.950 850.800 553.050 852.900 ;
        RECT 544.950 847.950 547.050 850.050 ;
        RECT 551.400 844.050 552.600 850.800 ;
        RECT 550.950 841.950 553.050 844.050 ;
        RECT 541.950 832.950 544.050 835.050 ;
        RECT 547.950 832.950 550.050 835.050 ;
        RECT 553.950 832.950 556.050 835.050 ;
        RECT 538.950 817.950 541.050 820.050 ;
        RECT 532.950 814.950 535.050 817.050 ;
        RECT 533.400 808.050 534.600 814.950 ;
        RECT 532.950 805.950 535.050 808.050 ;
        RECT 524.400 801.000 528.600 801.600 ;
        RECT 523.950 800.400 528.600 801.000 ;
        RECT 523.950 796.950 526.050 800.400 ;
        RECT 535.950 799.950 538.050 802.050 ;
        RECT 529.950 798.600 534.000 799.050 ;
        RECT 529.950 798.000 534.600 798.600 ;
        RECT 529.950 796.950 535.050 798.000 ;
        RECT 532.950 793.950 535.050 796.950 ;
        RECT 536.400 787.050 537.600 799.950 ;
        RECT 542.400 790.050 543.600 832.950 ;
        RECT 548.400 829.050 549.600 832.950 ;
        RECT 547.950 826.950 550.050 829.050 ;
        RECT 554.400 823.050 555.600 832.950 ;
        RECT 553.950 820.950 556.050 823.050 ;
        RECT 550.950 814.950 553.050 817.050 ;
        RECT 551.400 811.050 552.600 814.950 ;
        RECT 557.400 811.050 558.600 853.950 ;
        RECT 565.950 847.950 568.050 850.050 ;
        RECT 566.400 844.050 567.600 847.950 ;
        RECT 565.950 841.950 568.050 844.050 ;
        RECT 569.400 835.050 570.600 856.950 ;
        RECT 571.950 850.950 574.050 853.050 ;
        RECT 568.950 832.950 571.050 835.050 ;
        RECT 559.950 817.950 562.050 820.050 ;
        RECT 550.950 808.950 553.050 811.050 ;
        RECT 556.950 808.950 559.050 811.050 ;
        RECT 560.400 802.050 561.600 817.950 ;
        RECT 572.400 817.050 573.600 850.950 ;
        RECT 581.400 850.050 582.600 856.950 ;
        RECT 577.800 847.950 579.900 850.050 ;
        RECT 581.100 847.950 583.200 850.050 ;
        RECT 578.400 826.050 579.600 847.950 ;
        RECT 581.400 844.050 582.600 847.950 ;
        RECT 584.400 846.600 585.600 884.400 ;
        RECT 613.950 877.950 616.050 880.050 ;
        RECT 592.950 874.950 595.050 877.050 ;
        RECT 598.950 874.950 601.050 877.050 ;
        RECT 593.400 865.050 594.600 874.950 ;
        RECT 592.950 862.950 595.050 865.050 ;
        RECT 593.400 853.050 594.600 862.950 ;
        RECT 599.400 859.050 600.600 874.950 ;
        RECT 610.950 865.800 613.050 867.900 ;
        RECT 598.950 856.950 601.050 859.050 ;
        RECT 592.950 850.950 595.050 853.050 ;
        RECT 584.400 846.000 591.600 846.600 ;
        RECT 584.400 845.400 592.050 846.000 ;
        RECT 581.400 842.400 586.050 844.050 ;
        RECT 582.000 841.950 586.050 842.400 ;
        RECT 589.950 841.950 592.050 845.400 ;
        RECT 601.950 841.950 604.050 844.050 ;
        RECT 580.950 832.950 583.050 835.050 ;
        RECT 581.400 829.050 582.600 832.950 ;
        RECT 586.950 829.950 589.050 832.050 ;
        RECT 580.950 826.950 583.050 829.050 ;
        RECT 577.950 823.950 580.050 826.050 ;
        RECT 578.400 820.200 579.600 823.950 ;
        RECT 577.950 818.100 580.050 820.200 ;
        RECT 571.950 814.950 574.050 817.050 ;
        RECT 577.950 814.800 580.050 816.900 ;
        RECT 565.950 811.950 568.050 814.050 ;
        RECT 547.950 798.600 550.050 802.050 ;
        RECT 559.950 799.950 562.050 802.050 ;
        RECT 547.950 798.000 552.600 798.600 ;
        RECT 548.400 797.400 552.600 798.000 ;
        RECT 551.400 793.050 552.600 797.400 ;
        RECT 550.950 790.950 553.050 793.050 ;
        RECT 566.400 790.050 567.600 811.950 ;
        RECT 578.400 808.050 579.600 814.800 ;
        RECT 587.400 814.050 588.600 829.950 ;
        RECT 602.400 814.050 603.600 841.950 ;
        RECT 611.400 835.050 612.600 865.800 ;
        RECT 614.400 865.050 615.600 877.950 ;
        RECT 620.400 871.050 621.600 898.950 ;
        RECT 643.950 895.950 646.050 898.050 ;
        RECT 658.950 895.950 661.050 898.050 ;
        RECT 644.400 889.050 645.600 895.950 ;
        RECT 637.950 888.600 640.050 889.050 ;
        RECT 629.400 887.400 640.050 888.600 ;
        RECT 629.400 880.050 630.600 887.400 ;
        RECT 637.950 886.950 640.050 887.400 ;
        RECT 643.950 886.950 646.050 889.050 ;
        RECT 659.400 880.050 660.600 895.950 ;
        RECT 685.950 885.600 690.000 886.050 ;
        RECT 685.950 883.950 690.600 885.600 ;
        RECT 628.950 877.950 631.050 880.050 ;
        RECT 634.950 877.950 637.050 880.050 ;
        RECT 645.000 879.600 649.050 880.050 ;
        RECT 644.400 877.950 649.050 879.600 ;
        RECT 658.950 877.950 661.050 880.050 ;
        RECT 635.400 874.050 636.600 877.950 ;
        RECT 640.950 874.950 643.050 877.050 ;
        RECT 634.950 871.950 637.050 874.050 ;
        RECT 619.950 868.950 622.050 871.050 ;
        RECT 628.950 868.950 631.050 871.050 ;
        RECT 625.950 865.950 628.050 868.050 ;
        RECT 613.950 862.950 616.050 865.050 ;
        RECT 619.950 850.950 622.050 853.050 ;
        RECT 613.950 843.600 616.050 844.050 ;
        RECT 620.400 843.600 621.600 850.950 ;
        RECT 613.950 843.000 621.600 843.600 ;
        RECT 613.950 842.400 622.050 843.000 ;
        RECT 613.950 841.950 616.050 842.400 ;
        RECT 619.950 838.950 622.050 842.400 ;
        RECT 610.950 832.950 613.050 835.050 ;
        RECT 607.950 817.950 610.050 820.050 ;
        RECT 586.950 811.950 589.050 814.050 ;
        RECT 601.950 811.950 604.050 814.050 ;
        RECT 577.950 805.950 580.050 808.050 ;
        RECT 592.950 799.950 595.050 802.050 ;
        RECT 571.950 796.950 574.050 799.050 ;
        RECT 593.400 798.600 594.600 799.950 ;
        RECT 608.400 799.050 609.600 817.950 ;
        RECT 622.950 814.950 625.050 817.050 ;
        RECT 610.800 811.950 612.900 814.050 ;
        RECT 598.950 798.600 601.050 799.050 ;
        RECT 593.400 797.400 601.050 798.600 ;
        RECT 572.400 790.200 573.600 796.950 ;
        RECT 541.950 787.950 544.050 790.050 ;
        RECT 565.950 787.950 568.050 790.050 ;
        RECT 571.950 788.100 574.050 790.200 ;
        RECT 529.950 784.950 532.050 787.050 ;
        RECT 535.950 784.950 538.050 787.050 ;
        RECT 550.950 784.950 553.050 787.050 ;
        RECT 556.950 784.950 559.050 787.050 ;
        RECT 514.950 766.950 517.050 769.050 ;
        RECT 530.400 766.050 531.600 784.950 ;
        RECT 547.950 772.950 550.050 775.050 ;
        RECT 532.950 769.950 535.050 772.050 ;
        RECT 502.950 763.950 505.050 766.050 ;
        RECT 529.950 763.950 532.050 766.050 ;
        RECT 466.950 757.950 469.050 760.050 ;
        RECT 430.950 756.600 433.050 757.050 ;
        RECT 412.950 756.000 417.600 756.600 ;
        RECT 412.950 754.950 418.050 756.000 ;
        RECT 425.400 755.400 433.050 756.600 ;
        RECT 415.950 751.950 418.050 754.950 ;
        RECT 406.950 745.950 409.050 748.050 ;
        RECT 412.950 745.950 415.050 748.050 ;
        RECT 406.950 736.950 409.050 739.050 ;
        RECT 397.950 703.950 400.050 706.050 ;
        RECT 403.950 703.950 406.050 706.050 ;
        RECT 400.950 700.950 403.050 703.050 ;
        RECT 391.950 688.950 394.050 691.050 ;
        RECT 401.400 688.050 402.600 700.950 ;
        RECT 407.400 694.050 408.600 736.950 ;
        RECT 413.400 733.050 414.600 745.950 ;
        RECT 428.400 739.050 429.600 755.400 ;
        RECT 430.950 754.950 433.050 755.400 ;
        RECT 439.950 754.950 442.050 757.050 ;
        RECT 449.400 755.400 454.050 757.050 ;
        RECT 450.000 754.950 454.050 755.400 ;
        RECT 460.800 754.950 462.900 757.050 ;
        RECT 464.100 754.950 466.200 757.050 ;
        RECT 472.950 754.950 475.050 757.050 ;
        RECT 478.950 754.950 481.050 757.050 ;
        RECT 490.950 754.950 493.050 757.050 ;
        RECT 526.950 754.950 529.050 757.050 ;
        RECT 436.950 742.950 439.050 745.050 ;
        RECT 430.800 739.950 432.900 742.050 ;
        RECT 427.950 736.950 430.050 739.050 ;
        RECT 412.950 730.950 415.050 733.050 ;
        RECT 431.400 730.050 432.600 739.950 ;
        RECT 430.950 727.950 433.050 730.050 ;
        RECT 415.950 718.950 418.050 721.050 ;
        RECT 421.950 718.950 424.050 721.050 ;
        RECT 416.400 715.050 417.600 718.950 ;
        RECT 422.400 715.050 423.600 718.950 ;
        RECT 437.400 715.050 438.600 742.950 ;
        RECT 415.950 712.950 418.050 715.050 ;
        RECT 421.950 712.950 424.050 715.050 ;
        RECT 436.950 712.950 439.050 715.050 ;
        RECT 440.400 709.050 441.600 754.950 ;
        RECT 451.950 745.950 454.050 748.050 ;
        RECT 452.400 721.050 453.600 745.950 ;
        RECT 454.950 733.950 457.050 736.050 ;
        RECT 455.400 730.050 456.600 733.950 ;
        RECT 454.950 727.950 457.050 730.050 ;
        RECT 451.950 718.950 454.050 721.050 ;
        RECT 424.950 706.950 427.050 709.050 ;
        RECT 439.950 706.950 442.050 709.050 ;
        RECT 409.800 703.950 411.900 706.050 ;
        RECT 413.100 703.950 415.200 706.050 ;
        RECT 410.400 697.050 411.600 703.950 ;
        RECT 409.950 694.950 412.050 697.050 ;
        RECT 406.800 691.950 408.900 694.050 ;
        RECT 400.950 685.950 403.050 688.050 ;
        RECT 409.950 685.950 412.050 688.050 ;
        RECT 389.400 677.400 396.600 678.600 ;
        RECT 379.950 673.950 382.050 676.050 ;
        RECT 385.950 673.950 388.050 676.050 ;
        RECT 391.950 673.950 394.050 676.050 ;
        RECT 352.950 670.950 355.050 673.050 ;
        RECT 370.950 667.950 373.050 670.050 ;
        RECT 380.400 669.600 381.600 673.950 ;
        RECT 374.400 668.400 381.600 669.600 ;
        RECT 386.400 669.600 387.600 673.950 ;
        RECT 386.400 669.000 390.600 669.600 ;
        RECT 386.400 668.400 391.050 669.000 ;
        RECT 364.950 664.950 367.050 667.050 ;
        RECT 349.950 658.950 352.050 661.050 ;
        RECT 350.400 634.050 351.600 658.950 ;
        RECT 365.400 652.050 366.600 664.950 ;
        RECT 371.400 652.050 372.600 667.950 ;
        RECT 374.400 661.050 375.600 668.400 ;
        RECT 388.950 667.050 391.050 668.400 ;
        RECT 385.800 664.950 387.900 667.050 ;
        RECT 388.950 666.000 391.200 667.050 ;
        RECT 389.100 664.950 391.200 666.000 ;
        RECT 373.950 658.950 376.050 661.050 ;
        RECT 355.950 649.950 358.050 652.050 ;
        RECT 364.950 649.950 367.050 652.050 ;
        RECT 370.950 649.950 373.050 652.050 ;
        RECT 356.400 634.050 357.600 649.950 ;
        RECT 386.400 646.050 387.600 664.950 ;
        RECT 376.950 643.950 379.050 646.050 ;
        RECT 385.950 643.950 388.050 646.050 ;
        RECT 361.950 640.950 364.050 643.050 ;
        RECT 367.950 640.950 370.050 643.050 ;
        RECT 349.950 631.950 352.050 634.050 ;
        RECT 355.950 631.950 358.050 634.050 ;
        RECT 334.950 625.950 337.050 628.050 ;
        RECT 346.950 625.950 349.050 628.050 ;
        RECT 335.400 619.050 336.600 625.950 ;
        RECT 362.400 625.050 363.600 640.950 ;
        RECT 368.400 628.050 369.600 640.950 ;
        RECT 373.950 631.950 376.050 634.050 ;
        RECT 367.950 625.950 370.050 628.050 ;
        RECT 361.800 622.950 363.900 625.050 ;
        RECT 334.950 616.950 337.050 619.050 ;
        RECT 343.950 616.950 346.050 619.050 ;
        RECT 358.950 616.950 361.050 619.050 ;
        RECT 319.950 613.950 322.050 616.050 ;
        RECT 329.100 613.950 331.200 616.050 ;
        RECT 335.400 610.050 336.600 616.950 ;
        RECT 340.950 613.950 343.050 616.050 ;
        RECT 341.400 610.050 342.600 613.950 ;
        RECT 313.950 607.950 316.050 610.050 ;
        RECT 319.950 609.600 322.050 610.050 ;
        RECT 319.950 608.400 327.600 609.600 ;
        RECT 319.950 607.950 322.050 608.400 ;
        RECT 316.950 598.950 319.050 601.050 ;
        RECT 317.400 589.050 318.600 598.950 ;
        RECT 316.950 586.950 319.050 589.050 ;
        RECT 326.400 583.200 327.600 608.400 ;
        RECT 334.950 607.950 337.050 610.050 ;
        RECT 340.950 607.950 343.050 610.050 ;
        RECT 344.400 601.050 345.600 616.950 ;
        RECT 359.400 610.050 360.600 616.950 ;
        RECT 358.950 607.950 361.050 610.050 ;
        RECT 364.950 607.950 367.050 610.050 ;
        RECT 343.950 598.950 346.050 601.050 ;
        RECT 349.950 600.600 352.050 601.050 ;
        RECT 355.950 600.600 358.050 601.050 ;
        RECT 349.950 599.400 358.050 600.600 ;
        RECT 349.950 598.950 352.050 599.400 ;
        RECT 355.950 598.950 358.050 599.400 ;
        RECT 337.950 595.950 340.050 598.050 ;
        RECT 325.950 581.100 328.050 583.200 ;
        RECT 304.800 577.950 306.900 580.050 ;
        RECT 308.100 577.950 310.200 580.050 ;
        RECT 316.950 577.950 319.050 580.050 ;
        RECT 305.400 574.050 306.600 577.950 ;
        RECT 304.950 571.950 307.050 574.050 ;
        RECT 301.950 562.950 304.050 565.050 ;
        RECT 307.950 562.950 310.050 565.050 ;
        RECT 308.400 559.050 309.600 562.950 ;
        RECT 307.950 556.950 310.050 559.050 ;
        RECT 317.400 541.050 318.600 577.950 ;
        RECT 325.950 577.800 328.050 579.900 ;
        RECT 326.400 574.050 327.600 577.800 ;
        RECT 325.950 571.950 328.050 574.050 ;
        RECT 334.950 571.950 337.050 574.050 ;
        RECT 328.950 553.950 331.050 556.050 ;
        RECT 322.950 547.950 325.050 550.050 ;
        RECT 316.950 538.950 319.050 541.050 ;
        RECT 317.400 532.050 318.600 538.950 ;
        RECT 319.950 535.950 322.050 538.050 ;
        RECT 280.950 529.950 283.050 532.050 ;
        RECT 296.400 530.400 301.050 532.050 ;
        RECT 297.000 529.950 301.050 530.400 ;
        RECT 304.950 531.600 309.000 532.050 ;
        RECT 304.950 529.950 309.600 531.600 ;
        RECT 316.950 529.950 319.050 532.050 ;
        RECT 277.950 520.950 280.050 523.050 ;
        RECT 301.950 522.600 304.050 523.050 ;
        RECT 293.400 521.400 304.050 522.600 ;
        RECT 293.400 517.050 294.600 521.400 ;
        RECT 301.950 520.950 304.050 521.400 ;
        RECT 292.950 514.950 295.050 517.050 ;
        RECT 308.400 514.050 309.600 529.950 ;
        RECT 320.400 523.050 321.600 535.950 ;
        RECT 323.400 532.050 324.600 547.950 ;
        RECT 329.400 541.050 330.600 553.950 ;
        RECT 335.400 553.050 336.600 571.950 ;
        RECT 334.950 550.950 337.050 553.050 ;
        RECT 338.400 550.050 339.600 595.950 ;
        RECT 365.400 592.050 366.600 607.950 ;
        RECT 340.950 589.950 343.050 592.050 ;
        RECT 364.950 589.950 367.050 592.050 ;
        RECT 341.400 565.050 342.600 589.950 ;
        RECT 349.950 586.950 352.050 589.050 ;
        RECT 346.950 580.950 349.050 583.050 ;
        RECT 347.400 574.050 348.600 580.950 ;
        RECT 350.400 580.050 351.600 586.950 ;
        RECT 355.950 580.950 358.050 583.050 ;
        RECT 349.950 577.950 352.050 580.050 ;
        RECT 346.950 571.950 349.050 574.050 ;
        RECT 350.400 565.050 351.600 577.950 ;
        RECT 341.400 563.400 346.050 565.050 ;
        RECT 342.000 562.950 346.050 563.400 ;
        RECT 349.950 562.950 352.050 565.050 ;
        RECT 356.400 559.050 357.600 580.950 ;
        RECT 365.400 565.050 366.600 589.950 ;
        RECT 368.400 583.050 369.600 625.950 ;
        RECT 374.400 625.050 375.600 631.950 ;
        RECT 373.950 622.950 376.050 625.050 ;
        RECT 373.950 613.950 376.050 616.050 ;
        RECT 370.950 598.950 373.050 601.050 ;
        RECT 367.950 580.950 370.050 583.050 ;
        RECT 371.400 580.050 372.600 598.950 ;
        RECT 374.400 589.050 375.600 613.950 ;
        RECT 377.400 592.050 378.600 643.950 ;
        RECT 392.400 631.050 393.600 673.950 ;
        RECT 391.950 628.950 394.050 631.050 ;
        RECT 385.950 619.950 388.050 622.050 ;
        RECT 386.400 610.050 387.600 619.950 ;
        RECT 391.950 613.950 394.050 616.050 ;
        RECT 392.400 610.050 393.600 613.950 ;
        RECT 385.950 607.950 388.050 610.050 ;
        RECT 391.950 607.950 394.050 610.050 ;
        RECT 388.950 598.950 391.050 601.050 ;
        RECT 376.950 589.950 379.050 592.050 ;
        RECT 373.950 586.950 376.050 589.050 ;
        RECT 389.400 586.050 390.600 598.950 ;
        RECT 388.950 583.950 391.050 586.050 ;
        RECT 395.400 580.050 396.600 677.400 ;
        RECT 403.950 667.950 406.050 670.050 ;
        RECT 404.400 652.050 405.600 667.950 ;
        RECT 406.950 664.950 409.050 667.050 ;
        RECT 407.400 661.050 408.600 664.950 ;
        RECT 406.950 658.950 409.050 661.050 ;
        RECT 410.400 658.050 411.600 685.950 ;
        RECT 409.950 655.950 412.050 658.050 ;
        RECT 403.950 649.950 406.050 652.050 ;
        RECT 413.400 637.050 414.600 703.950 ;
        RECT 425.400 685.050 426.600 706.950 ;
        RECT 461.400 706.050 462.600 754.950 ;
        RECT 467.100 751.950 469.200 754.050 ;
        RECT 467.400 736.050 468.600 751.950 ;
        RECT 473.400 739.050 474.600 754.950 ;
        RECT 479.400 751.050 480.600 754.950 ;
        RECT 478.950 748.950 481.050 751.050 ;
        RECT 484.950 748.950 487.050 751.050 ;
        RECT 481.950 745.950 484.050 748.050 ;
        RECT 472.950 736.950 475.050 739.050 ;
        RECT 466.950 733.950 469.050 736.050 ;
        RECT 468.000 729.600 472.050 730.050 ;
        RECT 467.400 727.950 472.050 729.600 ;
        RECT 475.950 727.950 478.050 730.050 ;
        RECT 467.400 715.050 468.600 727.950 ;
        RECT 472.950 718.950 475.050 721.050 ;
        RECT 466.950 712.950 469.050 715.050 ;
        RECT 460.950 703.950 463.050 706.050 ;
        RECT 430.950 694.950 433.050 697.050 ;
        RECT 460.950 694.950 463.050 697.050 ;
        RECT 424.950 682.950 427.050 685.050 ;
        RECT 421.950 678.600 424.050 679.050 ;
        RECT 427.950 678.600 430.050 679.200 ;
        RECT 421.950 677.400 430.050 678.600 ;
        RECT 421.950 676.950 424.050 677.400 ;
        RECT 427.950 677.100 430.050 677.400 ;
        RECT 427.950 673.800 430.050 675.900 ;
        RECT 424.950 670.950 427.050 673.050 ;
        RECT 421.950 655.950 424.050 658.050 ;
        RECT 422.400 652.050 423.600 655.950 ;
        RECT 421.950 649.950 424.050 652.050 ;
        RECT 425.400 643.050 426.600 670.950 ;
        RECT 428.400 658.050 429.600 673.800 ;
        RECT 431.400 661.050 432.600 694.950 ;
        RECT 461.400 688.050 462.600 694.950 ;
        RECT 454.950 684.600 457.050 688.050 ;
        RECT 460.950 685.950 463.050 688.050 ;
        RECT 452.400 684.000 457.050 684.600 ;
        RECT 452.400 683.400 456.600 684.000 ;
        RECT 452.400 679.200 453.600 683.400 ;
        RECT 451.950 677.100 454.050 679.200 ;
        RECT 457.950 676.950 460.050 679.050 ;
        RECT 442.950 673.950 445.050 676.050 ;
        RECT 443.400 670.050 444.600 673.950 ;
        RECT 451.950 673.800 454.050 675.900 ;
        RECT 442.950 667.950 445.050 670.050 ;
        RECT 442.800 661.950 444.900 664.050 ;
        RECT 446.100 661.950 448.200 664.050 ;
        RECT 430.950 658.950 433.050 661.050 ;
        RECT 427.950 655.950 430.050 658.050 ;
        RECT 418.950 640.950 421.050 643.050 ;
        RECT 424.950 640.950 427.050 643.050 ;
        RECT 427.950 640.950 430.050 643.050 ;
        RECT 412.950 634.950 415.050 637.050 ;
        RECT 409.950 631.950 412.050 634.050 ;
        RECT 410.400 616.050 411.600 631.950 ;
        RECT 415.950 628.950 418.050 631.050 ;
        RECT 416.400 622.050 417.600 628.950 ;
        RECT 419.400 625.050 420.600 640.950 ;
        RECT 418.950 622.950 421.050 625.050 ;
        RECT 415.950 619.950 418.050 622.050 ;
        RECT 409.950 613.950 412.050 616.050 ;
        RECT 406.950 607.950 409.050 610.050 ;
        RECT 407.400 586.050 408.600 607.950 ;
        RECT 410.400 601.050 411.600 613.950 ;
        RECT 416.400 610.050 417.600 619.950 ;
        RECT 415.950 607.950 418.050 610.050 ;
        RECT 420.000 606.600 424.050 607.050 ;
        RECT 419.400 604.950 424.050 606.600 ;
        RECT 410.400 599.400 415.050 601.050 ;
        RECT 411.000 598.950 415.050 599.400 ;
        RECT 419.400 592.050 420.600 604.950 ;
        RECT 418.950 589.950 421.050 592.050 ;
        RECT 406.950 583.950 409.050 586.050 ;
        RECT 412.950 580.950 415.050 583.050 ;
        RECT 370.950 577.950 373.050 580.050 ;
        RECT 394.950 577.950 397.050 580.050 ;
        RECT 371.400 574.050 372.600 577.950 ;
        RECT 370.950 571.950 373.050 574.050 ;
        RECT 413.400 565.050 414.600 580.950 ;
        RECT 365.400 563.400 370.050 565.050 ;
        RECT 366.000 562.950 370.050 563.400 ;
        RECT 373.950 562.950 376.050 565.050 ;
        RECT 388.950 562.950 391.050 565.050 ;
        RECT 394.950 562.950 397.050 565.050 ;
        RECT 412.950 562.950 415.050 565.050 ;
        RECT 374.400 559.050 375.600 562.950 ;
        RECT 340.950 556.950 343.050 559.050 ;
        RECT 355.950 556.950 358.050 559.050 ;
        RECT 373.950 556.950 376.050 559.050 ;
        RECT 337.950 547.950 340.050 550.050 ;
        RECT 328.950 538.950 331.050 541.050 ;
        RECT 322.950 529.950 325.050 532.050 ;
        RECT 341.400 523.050 342.600 556.950 ;
        RECT 343.950 550.950 346.050 553.050 ;
        RECT 349.950 550.950 352.050 553.050 ;
        RECT 367.950 550.950 370.050 553.050 ;
        RECT 344.400 532.050 345.600 550.950 ;
        RECT 350.400 538.050 351.600 550.950 ;
        RECT 355.950 541.950 358.050 544.050 ;
        RECT 349.950 535.950 352.050 538.050 ;
        RECT 350.400 532.050 351.600 535.950 ;
        RECT 343.950 529.950 346.050 532.050 ;
        RECT 349.950 529.950 352.050 532.050 ;
        RECT 319.950 520.950 322.050 523.050 ;
        RECT 340.950 520.950 343.050 523.050 ;
        RECT 325.950 517.950 328.050 520.050 ;
        RECT 326.400 514.050 327.600 517.950 ;
        RECT 337.950 514.950 340.050 517.050 ;
        RECT 268.950 511.950 271.050 514.050 ;
        RECT 307.950 511.950 310.050 514.050 ;
        RECT 325.950 511.950 328.050 514.050 ;
        RECT 298.950 508.950 301.050 511.050 ;
        RECT 316.950 508.950 319.050 511.050 ;
        RECT 250.950 505.950 253.050 508.050 ;
        RECT 253.950 495.600 256.050 496.050 ;
        RECT 259.950 495.600 262.050 496.050 ;
        RECT 253.950 494.400 262.050 495.600 ;
        RECT 253.950 493.950 256.050 494.400 ;
        RECT 259.950 493.950 262.050 494.400 ;
        RECT 262.950 484.950 265.050 487.050 ;
        RECT 280.950 484.950 283.050 487.050 ;
        RECT 263.400 481.050 264.600 484.950 ;
        RECT 281.400 481.050 282.600 484.950 ;
        RECT 262.950 478.950 265.050 481.050 ;
        RECT 271.950 478.950 274.050 481.050 ;
        RECT 280.950 478.950 283.050 481.050 ;
        RECT 286.950 478.950 289.050 481.050 ;
        RECT 272.400 466.050 273.600 478.950 ;
        RECT 287.400 475.050 288.600 478.950 ;
        RECT 280.950 472.950 283.050 475.050 ;
        RECT 286.950 472.950 289.050 475.050 ;
        RECT 281.400 466.050 282.600 472.950 ;
        RECT 289.950 469.950 292.050 472.050 ;
        RECT 271.950 463.950 274.050 466.050 ;
        RECT 280.950 463.950 283.050 466.050 ;
        RECT 205.950 460.950 208.050 463.050 ;
        RECT 214.950 460.950 217.050 463.050 ;
        RECT 241.950 460.950 244.050 463.050 ;
        RECT 259.950 460.950 262.050 463.050 ;
        RECT 215.400 454.050 216.600 460.950 ;
        RECT 260.400 454.050 261.600 460.950 ;
        RECT 272.400 457.050 273.600 463.950 ;
        RECT 271.950 454.950 274.050 457.050 ;
        RECT 193.950 451.950 196.050 454.050 ;
        RECT 199.950 451.950 202.050 454.050 ;
        RECT 214.950 451.950 217.050 454.050 ;
        RECT 196.950 442.950 199.050 445.050 ;
        RECT 190.950 439.950 193.050 442.050 ;
        RECT 184.950 433.950 187.050 436.050 ;
        RECT 160.950 427.950 163.050 430.050 ;
        RECT 169.950 427.950 172.050 430.050 ;
        RECT 161.400 412.050 162.600 427.950 ;
        RECT 178.950 415.950 181.050 418.050 ;
        RECT 160.950 409.950 163.050 412.050 ;
        RECT 169.950 409.950 172.050 412.050 ;
        RECT 151.950 394.950 154.050 397.050 ;
        RECT 160.950 391.950 163.050 394.050 ;
        RECT 145.950 373.950 148.050 376.050 ;
        RECT 139.950 370.950 142.050 373.050 ;
        RECT 133.950 361.950 136.050 364.050 ;
        RECT 140.400 361.050 141.600 370.950 ;
        RECT 118.950 358.950 121.050 361.050 ;
        RECT 139.950 358.950 142.050 361.050 ;
        RECT 146.400 358.050 147.600 373.950 ;
        RECT 161.400 373.050 162.600 391.950 ;
        RECT 170.400 388.050 171.600 409.950 ;
        RECT 179.400 388.050 180.600 415.950 ;
        RECT 169.950 385.950 172.050 388.050 ;
        RECT 178.950 385.950 181.050 388.050 ;
        RECT 191.400 382.050 192.600 439.950 ;
        RECT 197.400 436.200 198.600 442.950 ;
        RECT 200.400 439.050 201.600 451.950 ;
        RECT 220.950 450.600 223.050 454.050 ;
        RECT 259.950 451.950 262.050 454.050 ;
        RECT 264.000 453.600 268.050 454.050 ;
        RECT 263.400 451.950 268.050 453.600 ;
        RECT 226.950 450.600 229.050 451.050 ;
        RECT 220.950 450.000 229.050 450.600 ;
        RECT 221.400 449.400 229.050 450.000 ;
        RECT 216.000 444.600 220.050 445.050 ;
        RECT 215.400 442.950 220.050 444.600 ;
        RECT 199.950 436.950 202.050 439.050 ;
        RECT 196.950 434.100 199.050 436.200 ;
        RECT 196.950 430.800 199.050 432.900 ;
        RECT 197.400 412.050 198.600 430.800 ;
        RECT 215.400 430.050 216.600 442.950 ;
        RECT 221.400 439.050 222.600 449.400 ;
        RECT 226.950 448.950 229.050 449.400 ;
        RECT 223.950 444.600 228.000 445.050 ;
        RECT 223.950 442.950 228.600 444.600 ;
        RECT 244.950 442.950 247.050 445.050 ;
        RECT 256.950 442.950 259.050 445.050 ;
        RECT 220.950 436.950 223.050 439.050 ;
        RECT 227.400 435.600 228.600 442.950 ;
        RECT 232.950 436.950 235.050 439.050 ;
        RECT 227.400 434.400 231.600 435.600 ;
        RECT 214.950 427.950 217.050 430.050 ;
        RECT 223.950 427.950 226.050 430.050 ;
        RECT 224.400 412.050 225.600 427.950 ;
        RECT 196.950 409.950 199.050 412.050 ;
        RECT 205.950 409.950 208.050 412.050 ;
        RECT 214.950 409.950 217.050 412.050 ;
        RECT 223.950 409.950 226.050 412.050 ;
        RECT 206.400 406.050 207.600 409.950 ;
        RECT 215.400 406.050 216.600 409.950 ;
        RECT 205.950 403.950 208.050 406.050 ;
        RECT 214.950 403.950 217.050 406.050 ;
        RECT 196.950 391.950 199.050 394.050 ;
        RECT 190.950 379.950 193.050 382.050 ;
        RECT 197.400 376.050 198.600 391.950 ;
        RECT 215.400 391.050 216.600 403.950 ;
        RECT 214.950 388.950 217.050 391.050 ;
        RECT 230.400 379.050 231.600 434.400 ;
        RECT 233.400 433.050 234.600 436.950 ;
        RECT 238.950 433.950 241.050 436.050 ;
        RECT 232.950 430.950 235.050 433.050 ;
        RECT 223.950 376.050 226.050 379.050 ;
        RECT 229.950 376.950 232.050 379.050 ;
        RECT 168.000 375.600 172.050 376.050 ;
        RECT 167.400 373.950 172.050 375.600 ;
        RECT 175.950 373.950 178.050 376.050 ;
        RECT 184.950 375.600 187.050 376.050 ;
        RECT 190.950 375.600 193.050 376.050 ;
        RECT 184.950 374.400 193.050 375.600 ;
        RECT 184.950 373.950 187.050 374.400 ;
        RECT 190.950 373.950 193.050 374.400 ;
        RECT 196.950 373.950 199.050 376.050 ;
        RECT 214.950 373.950 217.050 376.050 ;
        RECT 220.950 375.000 226.050 376.050 ;
        RECT 220.950 374.400 225.600 375.000 ;
        RECT 220.950 373.950 225.000 374.400 ;
        RECT 160.950 370.950 163.050 373.050 ;
        RECT 148.950 364.950 151.050 367.050 ;
        RECT 149.400 361.050 150.600 364.950 ;
        RECT 167.400 361.050 168.600 373.950 ;
        RECT 148.950 358.950 151.050 361.050 ;
        RECT 166.950 358.950 169.050 361.050 ;
        RECT 112.950 355.950 115.050 358.050 ;
        RECT 145.950 355.950 148.050 358.050 ;
        RECT 176.400 355.050 177.600 373.950 ;
        RECT 185.100 364.950 187.200 367.050 ;
        RECT 199.950 364.950 202.050 367.050 ;
        RECT 205.950 364.950 208.050 367.050 ;
        RECT 175.950 352.950 178.050 355.050 ;
        RECT 112.950 345.600 115.050 346.050 ;
        RECT 112.950 344.400 117.600 345.600 ;
        RECT 112.950 343.950 115.050 344.400 ;
        RECT 113.400 340.050 114.600 343.950 ;
        RECT 116.400 340.050 117.600 344.400 ;
        RECT 145.950 342.600 148.050 343.050 ;
        RECT 137.400 341.400 148.050 342.600 ;
        RECT 112.950 337.950 115.050 340.050 ;
        RECT 116.400 338.400 121.050 340.050 ;
        RECT 117.000 337.950 121.050 338.400 ;
        RECT 137.400 334.050 138.600 341.400 ;
        RECT 145.950 340.950 148.050 341.400 ;
        RECT 160.950 339.600 163.050 343.050 ;
        RECT 166.950 339.600 169.050 340.050 ;
        RECT 160.950 339.000 169.050 339.600 ;
        RECT 161.400 338.400 169.050 339.000 ;
        RECT 166.950 337.950 169.050 338.400 ;
        RECT 172.950 337.950 175.050 340.050 ;
        RECT 136.950 331.950 139.050 334.050 ;
        RECT 145.950 331.950 148.050 334.050 ;
        RECT 109.950 328.950 112.050 331.050 ;
        RECT 110.400 325.050 111.600 328.950 ;
        RECT 109.950 322.950 112.050 325.050 ;
        RECT 110.400 319.050 111.600 322.950 ;
        RECT 109.950 316.950 112.050 319.050 ;
        RECT 146.400 316.050 147.600 331.950 ;
        RECT 163.950 328.950 166.050 331.050 ;
        RECT 169.950 328.950 172.050 331.050 ;
        RECT 145.950 313.950 148.050 316.050 ;
        RECT 164.400 313.050 165.600 328.950 ;
        RECT 170.400 319.050 171.600 328.950 ;
        RECT 169.950 316.950 172.050 319.050 ;
        RECT 163.950 310.950 166.050 313.050 ;
        RECT 173.400 310.050 174.600 337.950 ;
        RECT 178.950 333.600 183.000 334.050 ;
        RECT 178.950 331.950 183.600 333.600 ;
        RECT 178.950 316.950 181.050 319.050 ;
        RECT 103.950 307.950 106.050 310.050 ;
        RECT 172.950 307.950 175.050 310.050 ;
        RECT 104.400 298.050 105.600 307.950 ;
        RECT 127.950 304.950 130.050 307.050 ;
        RECT 128.400 298.050 129.600 304.950 ;
        RECT 100.950 295.950 103.050 298.050 ;
        RECT 104.400 296.400 109.050 298.050 ;
        RECT 120.000 297.600 124.050 298.050 ;
        RECT 105.000 295.950 109.050 296.400 ;
        RECT 119.400 295.950 124.050 297.600 ;
        RECT 127.950 295.950 130.050 298.050 ;
        RECT 145.950 295.950 148.050 298.050 ;
        RECT 119.400 289.050 120.600 295.950 ;
        RECT 67.950 288.600 70.050 289.050 ;
        RECT 73.950 288.600 76.050 289.050 ;
        RECT 67.950 287.400 76.050 288.600 ;
        RECT 67.950 286.950 70.050 287.400 ;
        RECT 73.950 286.950 76.050 287.400 ;
        RECT 85.950 286.950 88.050 289.050 ;
        RECT 91.950 288.600 94.050 289.050 ;
        RECT 97.950 288.600 100.050 289.050 ;
        RECT 91.950 287.400 100.050 288.600 ;
        RECT 91.950 286.950 94.050 287.400 ;
        RECT 97.950 286.950 100.050 287.400 ;
        RECT 118.950 286.950 121.050 289.050 ;
        RECT 136.950 286.950 139.050 289.050 ;
        RECT 142.950 286.950 145.050 289.050 ;
        RECT 52.950 283.950 55.050 286.050 ;
        RECT 112.950 280.950 115.050 283.050 ;
        RECT 55.950 274.950 58.050 277.050 ;
        RECT 56.400 229.050 57.600 274.950 ;
        RECT 79.950 271.950 82.050 274.050 ;
        RECT 70.950 264.600 73.050 265.050 ;
        RECT 62.400 263.400 73.050 264.600 ;
        RECT 62.400 256.050 63.600 263.400 ;
        RECT 70.950 262.950 73.050 263.400 ;
        RECT 61.950 253.950 64.050 256.050 ;
        RECT 70.950 253.950 73.050 256.050 ;
        RECT 71.400 238.050 72.600 253.950 ;
        RECT 80.400 247.050 81.600 271.950 ;
        RECT 85.950 268.950 88.050 271.050 ;
        RECT 97.950 268.950 100.050 271.050 ;
        RECT 86.400 262.050 87.600 268.950 ;
        RECT 91.950 265.950 94.050 268.050 ;
        RECT 92.400 262.050 93.600 265.950 ;
        RECT 85.950 259.950 88.050 262.050 ;
        RECT 91.950 259.950 94.050 262.050 ;
        RECT 88.950 250.950 91.050 253.050 ;
        RECT 94.950 250.950 97.050 253.050 ;
        RECT 89.400 247.050 90.600 250.950 ;
        RECT 79.950 244.950 82.050 247.050 ;
        RECT 88.950 244.950 91.050 247.050 ;
        RECT 95.400 238.050 96.600 250.950 ;
        RECT 70.950 235.950 73.050 238.050 ;
        RECT 94.950 235.950 97.050 238.050 ;
        RECT 64.950 232.950 67.050 235.050 ;
        RECT 55.950 226.950 58.050 229.050 ;
        RECT 49.950 220.950 52.050 223.050 ;
        RECT 50.400 205.050 51.600 220.950 ;
        RECT 56.400 208.050 57.600 226.950 ;
        RECT 65.400 223.050 66.600 232.950 ;
        RECT 64.950 220.950 67.050 223.050 ;
        RECT 65.400 208.050 66.600 220.950 ;
        RECT 56.400 206.400 61.050 208.050 ;
        RECT 57.000 205.950 61.050 206.400 ;
        RECT 64.950 205.950 67.050 208.050 ;
        RECT 49.950 202.950 52.050 205.050 ;
        RECT 71.400 204.600 72.600 235.950 ;
        RECT 85.950 229.950 88.050 232.050 ;
        RECT 76.950 211.950 79.050 214.050 ;
        RECT 77.400 208.050 78.600 211.950 ;
        RECT 86.400 208.050 87.600 229.950 ;
        RECT 91.950 208.950 94.050 211.050 ;
        RECT 77.400 206.400 82.050 208.050 ;
        RECT 78.000 205.950 82.050 206.400 ;
        RECT 85.950 205.950 88.050 208.050 ;
        RECT 68.400 203.400 72.600 204.600 ;
        RECT 46.950 187.950 49.050 190.050 ;
        RECT 52.950 187.950 55.050 190.050 ;
        RECT 16.950 151.950 19.050 154.050 ;
        RECT 22.950 151.950 25.050 154.050 ;
        RECT 31.950 151.950 34.050 154.050 ;
        RECT 40.950 151.950 43.050 154.050 ;
        RECT 17.400 142.050 18.600 151.950 ;
        RECT 22.950 145.950 25.050 148.050 ;
        RECT 23.400 142.050 24.600 145.950 ;
        RECT 16.950 139.950 19.050 142.050 ;
        RECT 22.950 139.950 25.050 142.050 ;
        RECT 19.950 130.950 22.050 133.050 ;
        RECT 13.950 127.950 16.050 130.050 ;
        RECT 14.400 121.050 15.600 127.950 ;
        RECT 20.400 124.050 21.600 130.950 ;
        RECT 19.950 121.950 22.050 124.050 ;
        RECT 25.950 121.950 28.050 124.050 ;
        RECT 13.950 118.950 16.050 121.050 ;
        RECT 16.950 103.950 19.050 106.050 ;
        RECT 10.950 97.950 13.050 100.050 ;
        RECT 11.400 94.050 12.600 97.950 ;
        RECT 10.950 91.950 13.050 94.050 ;
        RECT 17.400 82.050 18.600 103.950 ;
        RECT 26.400 94.050 27.600 121.950 ;
        RECT 28.950 112.950 31.050 115.050 ;
        RECT 29.400 100.050 30.600 112.950 ;
        RECT 28.950 97.950 31.050 100.050 ;
        RECT 25.950 91.950 28.050 94.050 ;
        RECT 32.400 82.050 33.600 151.950 ;
        RECT 34.950 148.950 37.050 151.050 ;
        RECT 35.400 142.050 36.600 148.950 ;
        RECT 47.400 148.050 48.600 187.950 ;
        RECT 53.400 184.050 54.600 187.950 ;
        RECT 49.950 181.950 52.050 184.050 ;
        RECT 53.400 182.400 58.050 184.050 ;
        RECT 54.000 181.950 58.050 182.400 ;
        RECT 50.400 169.050 51.600 181.950 ;
        RECT 49.950 166.950 52.050 169.050 ;
        RECT 68.400 166.050 69.600 203.400 ;
        RECT 92.400 196.050 93.600 208.950 ;
        RECT 98.400 199.050 99.600 268.950 ;
        RECT 113.400 268.050 114.600 280.950 ;
        RECT 137.400 274.050 138.600 286.950 ;
        RECT 143.400 283.050 144.600 286.950 ;
        RECT 142.950 280.950 145.050 283.050 ;
        RECT 146.400 277.050 147.600 295.950 ;
        RECT 172.950 292.950 175.050 295.050 ;
        RECT 153.000 288.600 157.050 289.050 ;
        RECT 152.400 286.950 157.050 288.600 ;
        RECT 152.400 283.050 153.600 286.950 ;
        RECT 151.950 280.950 154.050 283.050 ;
        RECT 145.950 274.950 148.050 277.050 ;
        RECT 173.400 274.050 174.600 292.950 ;
        RECT 136.950 271.950 139.050 274.050 ;
        RECT 148.950 271.950 151.050 274.050 ;
        RECT 172.950 271.950 175.050 274.050 ;
        RECT 112.950 265.950 115.050 268.050 ;
        RECT 130.950 261.600 133.050 265.050 ;
        RECT 136.950 261.600 139.050 262.050 ;
        RECT 142.950 261.600 145.050 262.050 ;
        RECT 130.950 261.000 145.050 261.600 ;
        RECT 131.400 260.400 145.050 261.000 ;
        RECT 136.950 259.950 139.050 260.400 ;
        RECT 142.950 259.950 145.050 260.400 ;
        RECT 100.950 253.950 103.050 256.050 ;
        RECT 101.400 232.050 102.600 253.950 ;
        RECT 133.950 250.950 136.050 253.050 ;
        RECT 121.950 238.950 124.050 241.050 ;
        RECT 100.950 229.950 103.050 232.050 ;
        RECT 109.950 229.950 112.050 232.050 ;
        RECT 110.400 220.050 111.600 229.950 ;
        RECT 109.950 217.950 112.050 220.050 ;
        RECT 122.400 219.600 123.600 238.950 ;
        RECT 134.400 235.050 135.600 250.950 ;
        RECT 133.950 232.950 136.050 235.050 ;
        RECT 139.950 229.950 142.050 232.050 ;
        RECT 124.950 220.950 127.050 223.050 ;
        RECT 119.400 219.000 123.600 219.600 ;
        RECT 118.950 218.400 123.600 219.000 ;
        RECT 118.950 214.950 121.050 218.400 ;
        RECT 97.950 196.950 100.050 199.050 ;
        RECT 91.950 193.950 94.050 196.050 ;
        RECT 112.950 193.950 115.050 196.050 ;
        RECT 92.400 187.050 93.600 193.950 ;
        RECT 100.950 190.950 103.050 193.050 ;
        RECT 101.400 187.050 102.600 190.950 ;
        RECT 91.950 184.950 94.050 187.050 ;
        RECT 100.950 184.950 103.050 187.050 ;
        RECT 113.400 184.050 114.600 193.950 ;
        RECT 113.400 182.400 118.050 184.050 ;
        RECT 114.000 181.950 118.050 182.400 ;
        RECT 94.950 175.950 97.050 178.050 ;
        RECT 73.950 172.950 76.050 175.050 ;
        RECT 79.950 172.950 82.050 175.050 ;
        RECT 67.950 163.950 70.050 166.050 ;
        RECT 74.400 154.050 75.600 172.950 ;
        RECT 80.400 169.050 81.600 172.950 ;
        RECT 79.950 166.950 82.050 169.050 ;
        RECT 91.950 163.950 94.050 166.050 ;
        RECT 92.400 160.050 93.600 163.950 ;
        RECT 91.950 157.950 94.050 160.050 ;
        RECT 79.950 154.950 82.050 157.050 ;
        RECT 73.950 151.950 76.050 154.050 ;
        RECT 40.950 145.950 43.050 148.050 ;
        RECT 46.800 145.950 48.900 148.050 ;
        RECT 55.950 145.950 58.050 148.050 ;
        RECT 41.400 142.050 42.600 145.950 ;
        RECT 34.950 139.950 37.050 142.050 ;
        RECT 40.950 139.950 43.050 142.050 ;
        RECT 35.400 124.050 36.600 139.950 ;
        RECT 37.950 124.950 40.050 127.050 ;
        RECT 34.950 121.950 37.050 124.050 ;
        RECT 38.400 115.050 39.600 124.950 ;
        RECT 37.950 112.950 40.050 115.050 ;
        RECT 38.400 106.050 39.600 112.950 ;
        RECT 37.950 103.950 40.050 106.050 ;
        RECT 41.400 99.600 42.600 139.950 ;
        RECT 47.400 130.050 48.600 145.950 ;
        RECT 56.400 142.050 57.600 145.950 ;
        RECT 80.400 142.050 81.600 154.950 ;
        RECT 95.400 154.050 96.600 175.950 ;
        RECT 118.950 174.600 121.050 175.050 ;
        RECT 125.400 174.600 126.600 220.950 ;
        RECT 133.950 220.050 136.050 223.050 ;
        RECT 133.950 219.000 139.050 220.050 ;
        RECT 134.400 218.400 139.050 219.000 ;
        RECT 135.000 217.950 139.050 218.400 ;
        RECT 140.400 211.050 141.600 229.950 ;
        RECT 142.950 219.600 147.000 220.050 ;
        RECT 142.950 217.950 147.600 219.600 ;
        RECT 146.400 211.050 147.600 217.950 ;
        RECT 133.950 208.950 136.050 211.050 ;
        RECT 139.950 208.950 142.050 211.050 ;
        RECT 145.950 208.950 148.050 211.050 ;
        RECT 134.400 205.050 135.600 208.950 ;
        RECT 133.950 202.950 136.050 205.050 ;
        RECT 134.400 199.050 135.600 202.950 ;
        RECT 133.950 196.950 136.050 199.050 ;
        RECT 136.950 193.950 139.050 196.050 ;
        RECT 137.400 175.050 138.600 193.950 ;
        RECT 139.950 190.950 142.050 193.050 ;
        RECT 140.400 184.050 141.600 190.950 ;
        RECT 139.950 183.600 142.050 184.050 ;
        RECT 145.950 183.600 148.050 184.050 ;
        RECT 139.950 182.400 148.050 183.600 ;
        RECT 139.950 181.950 142.050 182.400 ;
        RECT 145.950 181.950 148.050 182.400 ;
        RECT 118.950 173.400 126.600 174.600 ;
        RECT 118.950 172.950 121.050 173.400 ;
        RECT 115.950 154.950 118.050 157.050 ;
        RECT 94.950 151.950 97.050 154.050 ;
        RECT 103.950 145.950 106.050 148.050 ;
        RECT 94.950 142.950 97.050 145.050 ;
        RECT 55.950 139.950 58.050 142.050 ;
        RECT 60.000 141.600 64.050 142.050 ;
        RECT 59.400 139.950 64.050 141.600 ;
        RECT 73.950 139.950 76.050 142.050 ;
        RECT 79.950 139.950 82.050 142.050 ;
        RECT 85.950 141.600 90.000 142.050 ;
        RECT 85.950 139.950 90.600 141.600 ;
        RECT 59.400 138.600 60.600 139.950 ;
        RECT 56.400 137.400 60.600 138.600 ;
        RECT 56.400 130.050 57.600 137.400 ;
        RECT 58.950 130.950 61.050 133.050 ;
        RECT 46.950 127.950 49.050 130.050 ;
        RECT 55.950 127.950 58.050 130.050 ;
        RECT 59.400 127.050 60.600 130.950 ;
        RECT 58.950 124.950 61.050 127.050 ;
        RECT 67.950 121.950 70.050 124.050 ;
        RECT 46.950 120.600 51.000 121.050 ;
        RECT 46.950 118.950 51.600 120.600 ;
        RECT 43.950 115.950 46.050 118.050 ;
        RECT 38.400 98.400 42.600 99.600 ;
        RECT 38.400 97.050 39.600 98.400 ;
        RECT 44.400 97.050 45.600 115.950 ;
        RECT 34.950 95.400 39.600 97.050 ;
        RECT 40.950 95.400 45.600 97.050 ;
        RECT 34.950 94.950 39.000 95.400 ;
        RECT 40.950 94.950 45.000 95.400 ;
        RECT 16.950 81.600 19.050 82.050 ;
        RECT 16.950 80.400 21.600 81.600 ;
        RECT 16.950 79.950 19.050 80.400 ;
        RECT 13.950 70.950 16.050 73.050 ;
        RECT 14.400 52.050 15.600 70.950 ;
        RECT 20.400 52.050 21.600 80.400 ;
        RECT 31.950 79.950 34.050 82.050 ;
        RECT 40.950 73.950 43.050 76.050 ;
        RECT 31.950 67.950 34.050 70.050 ;
        RECT 32.400 64.050 33.600 67.950 ;
        RECT 41.400 64.050 42.600 73.950 ;
        RECT 50.400 73.050 51.600 118.950 ;
        RECT 61.950 112.950 64.050 115.050 ;
        RECT 62.400 109.050 63.600 112.950 ;
        RECT 68.400 109.050 69.600 121.950 ;
        RECT 74.400 118.050 75.600 139.950 ;
        RECT 82.950 130.950 85.050 133.050 ;
        RECT 83.400 127.050 84.600 130.950 ;
        RECT 89.400 127.050 90.600 139.950 ;
        RECT 82.950 124.950 85.050 127.050 ;
        RECT 88.950 124.950 91.050 127.050 ;
        RECT 83.400 118.050 84.600 124.950 ;
        RECT 91.950 121.950 94.050 124.050 ;
        RECT 73.950 115.950 76.050 118.050 ;
        RECT 82.950 115.950 85.050 118.050 ;
        RECT 61.950 106.950 64.050 109.050 ;
        RECT 67.950 106.950 70.050 109.050 ;
        RECT 55.950 103.950 58.050 106.050 ;
        RECT 56.400 88.050 57.600 103.950 ;
        RECT 55.950 85.950 58.050 88.050 ;
        RECT 62.400 85.050 63.600 106.950 ;
        RECT 92.400 106.050 93.600 121.950 ;
        RECT 95.400 115.050 96.600 142.950 ;
        RECT 104.400 139.050 105.600 145.950 ;
        RECT 103.950 136.950 106.050 139.050 ;
        RECT 100.950 132.600 103.050 133.050 ;
        RECT 109.950 132.600 112.050 133.050 ;
        RECT 100.950 131.400 112.050 132.600 ;
        RECT 100.950 130.950 103.050 131.400 ;
        RECT 109.950 130.950 112.050 131.400 ;
        RECT 97.950 124.950 100.050 127.050 ;
        RECT 94.800 112.950 96.900 115.050 ;
        RECT 98.400 112.050 99.600 124.950 ;
        RECT 116.400 118.050 117.600 154.950 ;
        RECT 125.400 130.050 126.600 173.400 ;
        RECT 133.950 172.950 136.050 175.050 ;
        RECT 136.950 172.950 139.050 175.050 ;
        RECT 134.400 130.050 135.600 172.950 ;
        RECT 139.950 136.950 142.050 139.050 ;
        RECT 124.950 127.950 127.050 130.050 ;
        RECT 133.950 127.950 136.050 130.050 ;
        RECT 140.400 121.050 141.600 136.950 ;
        RECT 149.400 132.600 150.600 271.950 ;
        RECT 172.950 265.950 175.050 268.050 ;
        RECT 173.400 258.600 174.600 265.950 ;
        RECT 170.400 258.000 174.600 258.600 ;
        RECT 169.950 257.400 174.600 258.000 ;
        RECT 169.950 253.950 172.050 257.400 ;
        RECT 160.950 249.600 163.050 253.050 ;
        RECT 169.950 249.600 172.050 250.050 ;
        RECT 160.950 249.000 172.050 249.600 ;
        RECT 161.400 248.400 172.050 249.000 ;
        RECT 169.950 247.950 172.050 248.400 ;
        RECT 179.400 244.050 180.600 316.950 ;
        RECT 182.400 316.050 183.600 331.950 ;
        RECT 185.400 319.050 186.600 364.950 ;
        RECT 193.950 355.950 196.050 358.050 ;
        RECT 184.950 316.950 187.050 319.050 ;
        RECT 181.950 313.950 184.050 316.050 ;
        RECT 182.400 301.050 183.600 313.950 ;
        RECT 194.400 304.050 195.600 355.950 ;
        RECT 196.950 349.950 199.050 352.050 ;
        RECT 197.400 334.050 198.600 349.950 ;
        RECT 196.950 331.950 199.050 334.050 ;
        RECT 200.400 315.600 201.600 364.950 ;
        RECT 206.400 355.050 207.600 364.950 ;
        RECT 205.950 352.950 208.050 355.050 ;
        RECT 215.400 352.050 216.600 373.950 ;
        RECT 223.950 364.950 226.050 367.050 ;
        RECT 224.400 361.050 225.600 364.950 ;
        RECT 223.950 358.950 226.050 361.050 ;
        RECT 220.950 352.950 223.050 355.050 ;
        RECT 208.950 349.950 211.050 352.050 ;
        RECT 214.950 349.950 217.050 352.050 ;
        RECT 209.400 346.050 210.600 349.950 ;
        RECT 217.950 346.950 220.050 349.050 ;
        RECT 208.950 343.950 211.050 346.050 ;
        RECT 205.950 339.600 208.050 340.050 ;
        RECT 211.950 339.600 214.050 340.050 ;
        RECT 205.950 338.400 214.050 339.600 ;
        RECT 205.950 337.950 208.050 338.400 ;
        RECT 211.950 337.950 214.050 338.400 ;
        RECT 197.400 314.400 201.600 315.600 ;
        RECT 197.400 307.050 198.600 314.400 ;
        RECT 211.950 313.950 214.050 316.050 ;
        RECT 199.950 307.950 202.050 310.050 ;
        RECT 196.950 304.950 199.050 307.050 ;
        RECT 193.950 301.950 196.050 304.050 ;
        RECT 181.950 298.950 184.050 301.050 ;
        RECT 196.950 298.950 199.050 301.050 ;
        RECT 182.400 295.050 183.600 298.950 ;
        RECT 187.950 295.950 190.050 298.050 ;
        RECT 181.950 292.950 184.050 295.050 ;
        RECT 184.950 286.950 187.050 289.050 ;
        RECT 185.400 277.050 186.600 286.950 ;
        RECT 184.950 274.950 187.050 277.050 ;
        RECT 188.400 262.050 189.600 295.950 ;
        RECT 197.400 273.600 198.600 298.950 ;
        RECT 200.400 298.050 201.600 307.950 ;
        RECT 205.950 301.950 208.050 304.050 ;
        RECT 206.400 298.050 207.600 301.950 ;
        RECT 199.950 295.950 202.050 298.050 ;
        RECT 205.950 295.950 208.050 298.050 ;
        RECT 202.950 283.950 205.050 286.050 ;
        RECT 203.400 277.050 204.600 283.950 ;
        RECT 208.950 277.950 211.050 280.050 ;
        RECT 202.950 274.950 205.050 277.050 ;
        RECT 199.950 273.600 202.050 274.050 ;
        RECT 197.400 272.400 202.050 273.600 ;
        RECT 199.950 271.950 202.050 272.400 ;
        RECT 200.400 268.050 201.600 271.950 ;
        RECT 199.950 265.950 202.050 268.050 ;
        RECT 184.950 260.400 189.600 262.050 ;
        RECT 190.950 261.600 195.000 262.050 ;
        RECT 184.950 259.950 189.000 260.400 ;
        RECT 190.950 259.950 195.600 261.600 ;
        RECT 196.950 259.950 199.050 262.050 ;
        RECT 187.950 250.950 190.050 253.050 ;
        RECT 178.950 241.950 181.050 244.050 ;
        RECT 157.950 217.950 160.050 220.050 ;
        RECT 163.950 217.950 166.050 220.050 ;
        RECT 158.400 205.050 159.600 217.950 ;
        RECT 157.950 202.950 160.050 205.050 ;
        RECT 158.400 174.600 159.600 202.950 ;
        RECT 164.400 199.050 165.600 217.950 ;
        RECT 172.950 208.950 175.050 211.050 ;
        RECT 173.400 199.050 174.600 208.950 ;
        RECT 163.950 196.950 166.050 199.050 ;
        RECT 172.950 196.950 175.050 199.050 ;
        RECT 175.950 187.950 178.050 190.050 ;
        RECT 176.400 183.600 177.600 187.950 ;
        RECT 170.400 182.400 177.600 183.600 ;
        RECT 163.950 177.600 166.050 178.050 ;
        RECT 170.400 177.600 171.600 182.400 ;
        RECT 163.950 176.400 171.600 177.600 ;
        RECT 163.950 175.950 166.050 176.400 ;
        RECT 172.950 175.950 175.050 178.050 ;
        RECT 158.400 173.400 162.600 174.600 ;
        RECT 161.400 157.050 162.600 173.400 ;
        RECT 173.400 160.050 174.600 175.950 ;
        RECT 172.950 157.950 175.050 160.050 ;
        RECT 160.950 154.950 163.050 157.050 ;
        RECT 175.950 145.950 178.050 148.050 ;
        RECT 176.400 142.050 177.600 145.950 ;
        RECT 172.950 139.950 177.600 142.050 ;
        RECT 146.400 131.400 150.600 132.600 ;
        RECT 133.950 118.950 136.050 121.050 ;
        RECT 139.950 118.950 142.050 121.050 ;
        RECT 103.950 115.950 106.050 118.050 ;
        RECT 115.950 115.950 118.050 118.050 ;
        RECT 97.950 109.950 100.050 112.050 ;
        RECT 91.950 103.950 94.050 106.050 ;
        RECT 73.950 97.950 76.050 100.050 ;
        RECT 61.950 82.950 64.050 85.050 ;
        RECT 61.950 76.950 64.050 79.050 ;
        RECT 49.950 70.950 52.050 73.050 ;
        RECT 50.400 67.050 51.600 70.950 ;
        RECT 49.950 64.950 52.050 67.050 ;
        RECT 55.950 64.950 58.050 67.050 ;
        RECT 32.400 62.400 37.050 64.050 ;
        RECT 33.000 61.950 37.050 62.400 ;
        RECT 40.950 61.950 43.050 64.050 ;
        RECT 28.950 58.950 31.050 61.050 ;
        RECT 29.400 55.050 30.600 58.950 ;
        RECT 29.400 53.400 34.050 55.050 ;
        RECT 30.000 52.950 34.050 53.400 ;
        RECT 13.950 49.950 16.050 52.050 ;
        RECT 19.950 49.950 22.050 52.050 ;
        RECT 34.950 34.950 37.050 37.050 ;
        RECT 35.400 31.050 36.600 34.950 ;
        RECT 34.950 28.950 37.050 31.050 ;
        RECT 27.000 27.600 31.050 28.050 ;
        RECT 26.400 25.950 31.050 27.600 ;
        RECT 26.400 19.050 27.600 25.950 ;
        RECT 41.400 21.600 42.600 61.950 ;
        RECT 56.400 61.050 57.600 64.950 ;
        RECT 55.950 58.950 58.050 61.050 ;
        RECT 62.400 55.050 63.600 76.950 ;
        RECT 74.400 70.050 75.600 97.950 ;
        RECT 82.950 94.950 85.050 97.050 ;
        RECT 88.950 94.950 91.050 97.050 ;
        RECT 64.950 67.950 67.050 70.050 ;
        RECT 73.950 67.950 76.050 70.050 ;
        RECT 65.400 64.050 66.600 67.950 ;
        RECT 83.400 67.050 84.600 94.950 ;
        RECT 89.400 91.050 90.600 94.950 ;
        RECT 88.950 88.950 91.050 91.050 ;
        RECT 100.950 85.950 103.050 88.050 ;
        RECT 85.950 82.950 88.050 85.050 ;
        RECT 94.950 82.950 97.050 85.050 ;
        RECT 82.950 64.950 85.050 67.050 ;
        RECT 64.950 61.950 67.050 64.050 ;
        RECT 86.400 55.050 87.600 82.950 ;
        RECT 95.400 61.050 96.600 82.950 ;
        RECT 94.950 58.950 97.050 61.050 ;
        RECT 49.950 52.950 52.050 55.050 ;
        RECT 61.950 52.950 64.050 55.050 ;
        RECT 85.950 52.950 88.050 55.050 ;
        RECT 43.950 37.950 46.050 40.050 ;
        RECT 44.400 34.050 45.600 37.950 ;
        RECT 43.950 31.950 46.050 34.050 ;
        RECT 44.400 28.050 45.600 31.950 ;
        RECT 44.400 26.400 49.050 28.050 ;
        RECT 45.000 25.950 49.050 26.400 ;
        RECT 35.400 20.400 42.600 21.600 ;
        RECT 35.400 19.050 36.600 20.400 ;
        RECT 25.950 16.950 28.050 19.050 ;
        RECT 31.950 17.400 36.600 19.050 ;
        RECT 31.950 16.950 36.000 17.400 ;
        RECT 37.950 16.950 40.050 19.050 ;
        RECT 38.400 7.050 39.600 16.950 ;
        RECT 50.400 7.050 51.600 52.950 ;
        RECT 101.400 48.600 102.600 85.950 ;
        RECT 104.400 76.050 105.600 115.950 ;
        RECT 134.400 106.050 135.600 118.950 ;
        RECT 140.400 108.600 141.600 118.950 ;
        RECT 146.400 118.050 147.600 131.400 ;
        RECT 169.950 130.950 172.050 133.050 ;
        RECT 151.950 127.950 154.050 130.050 ;
        RECT 160.950 127.950 163.050 130.050 ;
        RECT 152.400 124.050 153.600 127.950 ;
        RECT 151.950 121.950 154.050 124.050 ;
        RECT 161.400 121.050 162.600 127.950 ;
        RECT 170.400 121.050 171.600 130.950 ;
        RECT 176.400 127.050 177.600 139.950 ;
        RECT 175.950 124.950 178.050 127.050 ;
        RECT 179.400 124.050 180.600 241.950 ;
        RECT 188.400 235.050 189.600 250.950 ;
        RECT 194.400 247.050 195.600 259.950 ;
        RECT 193.800 244.950 195.900 247.050 ;
        RECT 197.400 244.050 198.600 259.950 ;
        RECT 196.950 241.950 199.050 244.050 ;
        RECT 200.400 241.050 201.600 265.950 ;
        RECT 199.950 238.950 202.050 241.050 ;
        RECT 187.950 232.950 190.050 235.050 ;
        RECT 190.950 229.950 193.050 232.050 ;
        RECT 191.400 217.050 192.600 229.950 ;
        RECT 200.400 217.050 201.600 238.950 ;
        RECT 205.950 217.950 208.050 220.050 ;
        RECT 190.950 214.950 193.050 217.050 ;
        RECT 199.950 214.950 202.050 217.050 ;
        RECT 202.950 199.950 205.050 202.050 ;
        RECT 187.950 193.950 190.050 196.050 ;
        RECT 188.400 184.050 189.600 193.950 ;
        RECT 196.950 190.950 199.050 193.050 ;
        RECT 187.950 181.950 190.050 184.050 ;
        RECT 197.400 175.050 198.600 190.950 ;
        RECT 190.950 172.950 193.050 175.050 ;
        RECT 196.950 172.950 199.050 175.050 ;
        RECT 191.400 169.050 192.600 172.950 ;
        RECT 190.950 166.950 193.050 169.050 ;
        RECT 191.400 157.050 192.600 166.950 ;
        RECT 184.950 154.950 187.050 157.050 ;
        RECT 190.950 154.950 193.050 157.050 ;
        RECT 196.950 154.950 199.050 157.050 ;
        RECT 185.400 133.050 186.600 154.950 ;
        RECT 187.950 145.950 190.050 148.050 ;
        RECT 188.400 142.050 189.600 145.950 ;
        RECT 197.400 142.050 198.600 154.950 ;
        RECT 188.400 140.400 193.050 142.050 ;
        RECT 189.000 139.950 193.050 140.400 ;
        RECT 196.950 139.950 199.050 142.050 ;
        RECT 185.400 131.400 190.050 133.050 ;
        RECT 186.000 130.950 190.050 131.400 ;
        RECT 193.950 130.950 196.050 133.050 ;
        RECT 187.950 124.950 190.050 127.050 ;
        RECT 178.950 121.950 181.050 124.050 ;
        RECT 160.950 118.950 163.050 121.050 ;
        RECT 169.950 118.950 172.050 121.050 ;
        RECT 145.950 115.950 148.050 118.050 ;
        RECT 145.950 108.600 148.050 109.050 ;
        RECT 140.400 107.400 148.050 108.600 ;
        RECT 145.950 106.950 148.050 107.400 ;
        RECT 151.950 106.950 154.050 109.050 ;
        RECT 109.950 103.950 112.050 106.050 ;
        RECT 133.950 103.950 136.050 106.050 ;
        RECT 110.400 85.050 111.600 103.950 ;
        RECT 139.950 97.950 142.050 100.050 ;
        RECT 118.950 96.600 121.050 97.050 ;
        RECT 124.950 96.600 127.050 97.050 ;
        RECT 118.950 95.400 127.050 96.600 ;
        RECT 118.950 94.950 121.050 95.400 ;
        RECT 124.950 94.950 127.050 95.400 ;
        RECT 130.950 94.950 133.050 97.050 ;
        RECT 131.400 88.050 132.600 94.950 ;
        RECT 130.950 85.950 133.050 88.050 ;
        RECT 109.950 82.950 112.050 85.050 ;
        RECT 140.400 76.050 141.600 97.950 ;
        RECT 142.950 88.950 145.050 91.050 ;
        RECT 143.400 76.050 144.600 88.950 ;
        RECT 152.400 85.050 153.600 106.950 ;
        RECT 161.400 106.050 162.600 118.950 ;
        RECT 172.950 115.950 175.050 118.050 ;
        RECT 178.950 115.950 181.050 118.050 ;
        RECT 160.950 103.950 163.050 106.050 ;
        RECT 151.950 82.950 154.050 85.050 ;
        RECT 154.950 79.950 157.050 82.050 ;
        RECT 103.950 73.950 106.050 76.050 ;
        RECT 127.950 73.950 130.050 76.050 ;
        RECT 139.800 73.950 141.900 76.050 ;
        RECT 143.100 73.950 145.200 76.050 ;
        RECT 103.950 67.950 106.050 70.050 ;
        RECT 104.400 55.050 105.600 67.950 ;
        RECT 109.950 60.600 114.000 61.050 ;
        RECT 109.950 58.950 114.600 60.600 ;
        RECT 113.400 55.050 114.600 58.950 ;
        RECT 128.400 55.050 129.600 73.950 ;
        RECT 143.400 64.050 144.600 73.950 ;
        RECT 148.950 67.950 151.050 70.050 ;
        RECT 149.400 64.050 150.600 67.950 ;
        RECT 142.950 61.950 145.050 64.050 ;
        RECT 148.950 61.950 151.050 64.050 ;
        RECT 103.950 52.950 106.050 55.050 ;
        RECT 112.950 52.950 115.050 55.050 ;
        RECT 127.950 52.950 130.050 55.050 ;
        RECT 98.400 47.400 102.600 48.600 ;
        RECT 91.950 43.950 94.050 46.050 ;
        RECT 73.950 40.950 76.050 43.050 ;
        RECT 74.400 22.050 75.600 40.950 ;
        RECT 64.950 19.950 67.050 22.050 ;
        RECT 73.950 19.950 76.050 22.050 ;
        RECT 37.950 4.950 40.050 7.050 ;
        RECT 49.950 4.950 52.050 7.050 ;
        RECT 65.400 4.050 66.600 19.950 ;
        RECT 92.400 19.050 93.600 43.950 ;
        RECT 98.400 19.050 99.600 47.400 ;
        RECT 155.400 46.050 156.600 79.950 ;
        RECT 160.950 73.950 163.050 76.050 ;
        RECT 161.400 64.050 162.600 73.950 ;
        RECT 173.400 70.050 174.600 115.950 ;
        RECT 179.400 100.050 180.600 115.950 ;
        RECT 188.400 109.050 189.600 124.950 ;
        RECT 194.400 118.050 195.600 130.950 ;
        RECT 193.950 115.950 196.050 118.050 ;
        RECT 187.950 106.950 190.050 109.050 ;
        RECT 178.950 97.950 181.050 100.050 ;
        RECT 187.950 97.950 190.050 100.050 ;
        RECT 188.400 82.050 189.600 97.950 ;
        RECT 203.400 91.050 204.600 199.950 ;
        RECT 206.400 199.050 207.600 217.950 ;
        RECT 209.400 202.050 210.600 277.950 ;
        RECT 212.400 231.600 213.600 313.950 ;
        RECT 218.400 253.050 219.600 346.950 ;
        RECT 221.400 340.050 222.600 352.950 ;
        RECT 220.950 337.950 223.050 340.050 ;
        RECT 224.400 331.050 225.600 358.950 ;
        RECT 229.950 355.950 232.050 358.050 ;
        RECT 223.950 328.950 226.050 331.050 ;
        RECT 220.950 322.950 223.050 325.050 ;
        RECT 221.400 310.050 222.600 322.950 ;
        RECT 230.400 316.050 231.600 355.950 ;
        RECT 239.400 349.050 240.600 433.950 ;
        RECT 245.400 433.050 246.600 442.950 ;
        RECT 257.400 436.050 258.600 442.950 ;
        RECT 263.400 436.050 264.600 451.950 ;
        RECT 271.950 448.950 274.050 451.050 ;
        RECT 272.400 445.050 273.600 448.950 ;
        RECT 268.950 443.400 273.600 445.050 ;
        RECT 268.950 442.950 273.000 443.400 ;
        RECT 281.400 442.050 282.600 463.950 ;
        RECT 290.400 442.050 291.600 469.950 ;
        RECT 295.950 451.950 298.050 454.050 ;
        RECT 281.400 440.400 286.050 442.050 ;
        RECT 282.000 439.950 286.050 440.400 ;
        RECT 289.950 439.950 292.050 442.050 ;
        RECT 296.400 438.600 297.600 451.950 ;
        RECT 299.400 450.600 300.600 508.950 ;
        RECT 317.400 490.050 318.600 508.950 ;
        RECT 338.400 496.050 339.600 514.950 ;
        RECT 356.400 511.050 357.600 541.950 ;
        RECT 364.950 528.600 367.050 529.050 ;
        RECT 359.400 527.400 367.050 528.600 ;
        RECT 359.400 514.050 360.600 527.400 ;
        RECT 364.950 526.950 367.050 527.400 ;
        RECT 368.400 520.050 369.600 550.950 ;
        RECT 389.400 541.050 390.600 562.950 ;
        RECT 388.950 538.950 391.050 541.050 ;
        RECT 382.950 532.950 385.050 535.050 ;
        RECT 376.950 526.950 379.050 529.050 ;
        RECT 367.950 517.950 370.050 520.050 ;
        RECT 373.950 517.950 376.050 520.050 ;
        RECT 358.800 511.950 360.900 514.050 ;
        RECT 355.950 508.950 358.050 511.050 ;
        RECT 374.400 508.050 375.600 517.950 ;
        RECT 377.400 511.050 378.600 526.950 ;
        RECT 376.950 508.950 379.050 511.050 ;
        RECT 343.950 505.950 346.050 508.050 ;
        RECT 373.950 505.950 376.050 508.050 ;
        RECT 337.950 493.950 340.050 496.050 ;
        RECT 316.950 487.950 319.050 490.050 ;
        RECT 322.950 487.950 325.050 490.050 ;
        RECT 307.950 484.950 310.050 487.050 ;
        RECT 308.400 477.600 309.600 484.950 ;
        RECT 308.400 476.400 318.600 477.600 ;
        RECT 310.950 472.950 313.050 475.050 ;
        RECT 311.400 454.050 312.600 472.950 ;
        RECT 301.950 453.600 304.050 454.050 ;
        RECT 307.950 453.600 310.050 454.050 ;
        RECT 301.950 452.400 310.050 453.600 ;
        RECT 301.950 451.950 304.050 452.400 ;
        RECT 307.950 451.950 310.050 452.400 ;
        RECT 311.400 451.950 316.050 454.050 ;
        RECT 311.400 450.600 312.600 451.950 ;
        RECT 299.400 449.400 303.600 450.600 ;
        RECT 293.400 437.400 297.600 438.600 ;
        RECT 256.950 433.950 259.050 436.050 ;
        RECT 262.950 433.950 265.050 436.050 ;
        RECT 244.950 430.950 247.050 433.050 ;
        RECT 259.950 424.950 262.050 427.050 ;
        RECT 260.400 418.050 261.600 424.950 ;
        RECT 293.400 421.050 294.600 437.400 ;
        RECT 302.400 427.050 303.600 449.400 ;
        RECT 305.400 449.400 312.600 450.600 ;
        RECT 301.950 424.950 304.050 427.050 ;
        RECT 305.400 424.050 306.600 449.400 ;
        RECT 310.950 439.950 313.050 442.050 ;
        RECT 311.400 424.050 312.600 439.950 ;
        RECT 317.400 439.050 318.600 476.400 ;
        RECT 323.400 472.050 324.600 487.950 ;
        RECT 338.400 478.050 339.600 493.950 ;
        RECT 344.400 490.050 345.600 505.950 ;
        RECT 349.950 499.950 352.050 502.050 ;
        RECT 358.950 499.950 361.050 502.050 ;
        RECT 343.950 487.950 346.050 490.050 ;
        RECT 344.400 481.050 345.600 487.950 ;
        RECT 343.950 478.950 346.050 481.050 ;
        RECT 337.950 475.950 340.050 478.050 ;
        RECT 322.950 469.950 325.050 472.050 ;
        RECT 350.400 466.050 351.600 499.950 ;
        RECT 359.400 496.050 360.600 499.950 ;
        RECT 383.400 499.050 384.600 532.950 ;
        RECT 388.950 502.950 391.050 505.050 ;
        RECT 389.400 499.050 390.600 502.950 ;
        RECT 382.950 496.950 385.050 499.050 ;
        RECT 388.950 496.950 391.050 499.050 ;
        RECT 358.950 493.950 361.050 496.050 ;
        RECT 376.950 493.950 379.050 496.050 ;
        RECT 355.950 484.950 358.050 487.050 ;
        RECT 361.950 484.950 364.050 487.050 ;
        RECT 356.400 478.050 357.600 484.950 ;
        RECT 362.400 481.050 363.600 484.950 ;
        RECT 361.950 478.950 364.050 481.050 ;
        RECT 355.950 475.950 358.050 478.050 ;
        RECT 370.950 469.950 373.050 472.050 ;
        RECT 361.950 466.950 364.050 469.050 ;
        RECT 349.950 463.950 352.050 466.050 ;
        RECT 319.950 460.950 322.050 463.050 ;
        RECT 358.950 460.950 361.050 463.050 ;
        RECT 320.400 445.050 321.600 460.950 ;
        RECT 359.400 454.050 360.600 460.950 ;
        RECT 322.950 453.600 325.050 454.050 ;
        RECT 328.950 453.600 331.050 454.050 ;
        RECT 322.950 452.400 331.050 453.600 ;
        RECT 322.950 451.950 325.050 452.400 ;
        RECT 328.950 451.950 331.050 452.400 ;
        RECT 334.950 453.600 337.050 454.050 ;
        RECT 352.950 453.600 357.000 454.050 ;
        RECT 334.950 452.400 345.600 453.600 ;
        RECT 334.950 451.950 337.050 452.400 ;
        RECT 319.950 442.950 322.050 445.050 ;
        RECT 325.950 442.950 328.050 445.050 ;
        RECT 331.950 442.950 334.050 445.050 ;
        RECT 337.950 442.950 340.050 445.050 ;
        RECT 316.950 436.950 319.050 439.050 ;
        RECT 326.400 435.600 327.600 442.950 ;
        RECT 332.400 439.050 333.600 442.950 ;
        RECT 331.950 436.950 334.050 439.050 ;
        RECT 338.400 436.050 339.600 442.950 ;
        RECT 323.400 434.400 327.600 435.600 ;
        RECT 323.400 424.050 324.600 434.400 ;
        RECT 337.950 433.950 340.050 436.050 ;
        RECT 334.950 430.950 337.050 433.050 ;
        RECT 304.950 421.950 307.050 424.050 ;
        RECT 310.950 421.950 313.050 424.050 ;
        RECT 322.950 421.950 325.050 424.050 ;
        RECT 292.950 418.950 295.050 421.050 ;
        RECT 335.400 418.050 336.600 430.950 ;
        RECT 344.400 418.050 345.600 452.400 ;
        RECT 352.950 451.950 357.600 453.600 ;
        RECT 358.950 451.950 361.050 454.050 ;
        RECT 356.400 424.050 357.600 451.950 ;
        RECT 362.400 445.050 363.600 466.950 ;
        RECT 364.950 460.950 367.050 463.050 ;
        RECT 365.400 454.050 366.600 460.950 ;
        RECT 364.950 451.950 367.050 454.050 ;
        RECT 371.400 445.050 372.600 469.950 ;
        RECT 377.400 463.050 378.600 493.950 ;
        RECT 391.950 487.950 394.050 490.050 ;
        RECT 392.400 463.050 393.600 487.950 ;
        RECT 395.400 474.600 396.600 562.950 ;
        RECT 413.400 559.050 414.600 562.950 ;
        RECT 412.950 556.950 415.050 559.050 ;
        RECT 419.400 553.050 420.600 589.950 ;
        RECT 428.400 580.050 429.600 640.950 ;
        RECT 436.950 637.950 439.050 640.050 ;
        RECT 433.950 604.950 436.050 607.050 ;
        RECT 427.950 577.950 430.050 580.050 ;
        RECT 434.400 574.050 435.600 604.950 ;
        RECT 437.400 586.050 438.600 637.950 ;
        RECT 439.950 628.950 442.050 631.050 ;
        RECT 436.950 583.950 439.050 586.050 ;
        RECT 440.400 574.050 441.600 628.950 ;
        RECT 443.400 628.050 444.600 661.950 ;
        RECT 446.400 634.050 447.600 661.950 ;
        RECT 452.400 661.050 453.600 673.800 ;
        RECT 458.400 667.050 459.600 676.950 ;
        RECT 463.950 673.950 466.050 676.050 ;
        RECT 457.950 664.950 460.050 667.050 ;
        RECT 448.800 658.950 450.900 661.050 ;
        RECT 452.100 658.950 454.200 661.050 ;
        RECT 449.400 652.050 450.600 658.950 ;
        RECT 464.400 655.050 465.600 673.950 ;
        RECT 454.950 652.950 457.050 655.050 ;
        RECT 463.950 652.950 466.050 655.050 ;
        RECT 448.950 649.950 451.050 652.050 ;
        RECT 449.400 634.050 450.600 649.950 ;
        RECT 455.400 646.050 456.600 652.950 ;
        RECT 454.950 643.950 457.050 646.050 ;
        RECT 464.400 645.600 465.600 652.950 ;
        RECT 467.400 652.050 468.600 712.950 ;
        RECT 473.400 712.200 474.600 718.950 ;
        RECT 472.950 710.100 475.050 712.200 ;
        RECT 472.950 706.800 475.050 708.900 ;
        RECT 469.950 676.950 472.050 679.050 ;
        RECT 470.400 661.050 471.600 676.950 ;
        RECT 473.400 664.050 474.600 706.800 ;
        RECT 472.950 661.950 475.050 664.050 ;
        RECT 469.950 658.950 472.050 661.050 ;
        RECT 466.950 649.950 469.050 652.050 ;
        RECT 476.400 649.050 477.600 727.950 ;
        RECT 478.950 718.950 481.050 721.050 ;
        RECT 479.400 709.050 480.600 718.950 ;
        RECT 478.950 706.950 481.050 709.050 ;
        RECT 482.400 706.050 483.600 745.950 ;
        RECT 485.400 736.050 486.600 748.950 ;
        RECT 484.950 733.950 487.050 736.050 ;
        RECT 487.950 727.950 490.050 730.050 ;
        RECT 481.950 703.950 484.050 706.050 ;
        RECT 481.950 691.950 484.050 694.050 ;
        RECT 482.400 679.050 483.600 691.950 ;
        RECT 484.950 685.950 487.050 688.050 ;
        RECT 481.950 676.950 484.050 679.050 ;
        RECT 485.400 670.050 486.600 685.950 ;
        RECT 488.400 673.050 489.600 727.950 ;
        RECT 491.400 712.050 492.600 754.950 ;
        RECT 495.000 753.600 499.050 754.050 ;
        RECT 494.400 751.950 499.050 753.600 ;
        RECT 494.400 736.050 495.600 751.950 ;
        RECT 511.950 750.600 514.050 754.050 ;
        RECT 503.400 750.000 514.050 750.600 ;
        RECT 502.950 749.400 513.600 750.000 ;
        RECT 502.950 748.050 505.050 749.400 ;
        RECT 502.800 747.000 505.050 748.050 ;
        RECT 502.800 745.950 504.900 747.000 ;
        RECT 511.950 739.950 514.050 742.050 ;
        RECT 493.950 733.950 496.050 736.050 ;
        RECT 493.950 720.600 498.000 721.050 ;
        RECT 493.950 718.950 498.600 720.600 ;
        RECT 499.950 718.950 502.050 721.050 ;
        RECT 497.400 715.050 498.600 718.950 ;
        RECT 496.950 712.950 499.050 715.050 ;
        RECT 500.400 712.050 501.600 718.950 ;
        RECT 490.950 709.950 493.050 712.050 ;
        RECT 499.950 709.950 502.050 712.050 ;
        RECT 505.950 709.950 508.050 712.050 ;
        RECT 493.950 703.950 496.050 706.050 ;
        RECT 487.950 670.950 490.050 673.050 ;
        RECT 484.950 667.950 487.050 670.050 ;
        RECT 490.950 667.950 493.050 670.050 ;
        RECT 478.950 664.950 481.050 667.050 ;
        RECT 479.400 658.050 480.600 664.950 ;
        RECT 478.800 655.950 480.900 658.050 ;
        RECT 475.950 646.950 478.050 649.050 ;
        RECT 481.950 646.950 484.050 649.050 ;
        RECT 464.400 645.000 474.600 645.600 ;
        RECT 464.400 644.400 475.050 645.000 ;
        RECT 466.950 640.950 469.050 643.050 ;
        RECT 472.950 640.950 475.050 644.400 ;
        RECT 478.950 640.950 481.050 643.050 ;
        RECT 454.950 637.950 457.050 640.050 ;
        RECT 451.950 634.950 454.050 637.050 ;
        RECT 445.800 631.950 447.900 634.050 ;
        RECT 449.100 631.950 451.200 634.050 ;
        RECT 442.950 625.950 445.050 628.050 ;
        RECT 452.400 618.600 453.600 634.950 ;
        RECT 449.400 617.400 453.600 618.600 ;
        RECT 449.400 606.600 450.600 617.400 ;
        RECT 455.400 616.050 456.600 637.950 ;
        RECT 467.400 634.050 468.600 640.950 ;
        RECT 457.950 631.950 460.050 634.050 ;
        RECT 466.950 631.950 469.050 634.050 ;
        RECT 454.950 613.950 457.050 616.050 ;
        RECT 446.400 605.400 450.600 606.600 ;
        RECT 446.400 601.050 447.600 605.400 ;
        RECT 446.400 599.400 451.050 601.050 ;
        RECT 447.000 598.950 451.050 599.400 ;
        RECT 427.950 571.950 430.050 574.050 ;
        RECT 433.950 571.950 436.050 574.050 ;
        RECT 439.950 571.950 442.050 574.050 ;
        RECT 428.400 565.050 429.600 571.950 ;
        RECT 458.400 567.600 459.600 631.950 ;
        RECT 479.400 616.050 480.600 640.950 ;
        RECT 463.950 613.950 466.050 616.050 ;
        RECT 469.950 613.950 472.050 616.050 ;
        RECT 478.950 613.950 481.050 616.050 ;
        RECT 464.400 610.050 465.600 613.950 ;
        RECT 470.400 610.050 471.600 613.950 ;
        RECT 463.950 607.950 466.050 610.050 ;
        RECT 469.950 607.950 472.050 610.050 ;
        RECT 466.950 598.950 469.050 601.050 ;
        RECT 475.950 598.950 478.050 601.050 ;
        RECT 467.400 595.050 468.600 598.950 ;
        RECT 466.950 592.950 469.050 595.050 ;
        RECT 460.950 577.950 463.050 580.050 ;
        RECT 455.400 567.000 459.600 567.600 ;
        RECT 454.950 566.400 459.600 567.000 ;
        RECT 428.400 563.400 433.050 565.050 ;
        RECT 429.000 562.950 433.050 563.400 ;
        RECT 436.950 562.950 439.050 565.050 ;
        RECT 454.950 562.950 457.050 566.400 ;
        RECT 461.400 565.050 462.600 577.950 ;
        RECT 466.800 571.950 468.900 574.050 ;
        RECT 470.100 571.950 472.200 574.050 ;
        RECT 460.950 562.950 463.050 565.050 ;
        RECT 437.400 559.050 438.600 562.950 ;
        RECT 427.950 556.950 430.050 559.050 ;
        RECT 436.950 556.950 439.050 559.050 ;
        RECT 463.950 556.950 466.050 559.050 ;
        RECT 412.950 550.950 415.050 553.050 ;
        RECT 418.950 550.950 421.050 553.050 ;
        RECT 413.400 544.050 414.600 550.950 ;
        RECT 418.950 544.950 421.050 547.050 ;
        RECT 412.950 541.950 415.050 544.050 ;
        RECT 397.950 538.950 400.050 541.050 ;
        RECT 398.400 529.050 399.600 538.950 ;
        RECT 419.400 532.050 420.600 544.950 ;
        RECT 424.950 535.950 427.050 538.050 ;
        RECT 425.400 532.050 426.600 535.950 ;
        RECT 418.950 529.950 421.050 532.050 ;
        RECT 424.950 529.950 427.050 532.050 ;
        RECT 397.950 526.950 400.050 529.050 ;
        RECT 400.950 520.950 403.050 523.050 ;
        RECT 409.950 520.950 412.050 523.050 ;
        RECT 421.950 522.600 426.000 523.050 ;
        RECT 421.950 520.950 426.600 522.600 ;
        RECT 395.400 473.400 399.600 474.600 ;
        RECT 376.950 460.950 379.050 463.050 ;
        RECT 391.950 460.950 394.050 463.050 ;
        RECT 388.950 450.600 391.050 454.050 ;
        RECT 394.950 450.600 397.050 454.050 ;
        RECT 388.950 450.000 397.050 450.600 ;
        RECT 389.400 449.400 396.600 450.000 ;
        RECT 361.950 442.950 364.050 445.050 ;
        RECT 371.400 443.400 376.050 445.050 ;
        RECT 372.000 442.950 376.050 443.400 ;
        RECT 391.950 442.950 394.050 445.050 ;
        RECT 362.400 436.050 363.600 442.950 ;
        RECT 392.400 436.050 393.600 442.950 ;
        RECT 361.950 433.950 364.050 436.050 ;
        RECT 391.950 433.950 394.050 436.050 ;
        RECT 398.400 427.050 399.600 473.400 ;
        RECT 401.400 460.050 402.600 520.950 ;
        RECT 410.400 496.050 411.600 520.950 ;
        RECT 418.950 511.950 421.050 514.050 ;
        RECT 409.950 493.950 412.050 496.050 ;
        RECT 406.950 484.950 409.050 487.050 ;
        RECT 412.950 484.950 415.050 487.050 ;
        RECT 407.400 481.050 408.600 484.950 ;
        RECT 406.950 478.950 409.050 481.050 ;
        RECT 413.400 478.050 414.600 484.950 ;
        RECT 419.400 481.050 420.600 511.950 ;
        RECT 425.400 502.050 426.600 520.950 ;
        RECT 424.950 499.950 427.050 502.050 ;
        RECT 424.950 484.950 427.050 487.050 ;
        RECT 425.400 481.050 426.600 484.950 ;
        RECT 418.950 478.950 421.050 481.050 ;
        RECT 424.950 478.950 427.050 481.050 ;
        RECT 403.950 475.950 406.050 478.050 ;
        RECT 412.950 475.950 415.050 478.050 ;
        RECT 404.400 472.050 405.600 475.950 ;
        RECT 428.400 475.050 429.600 556.950 ;
        RECT 464.400 553.050 465.600 556.950 ;
        RECT 463.800 550.950 465.900 553.050 ;
        RECT 460.950 547.950 463.050 550.050 ;
        RECT 442.950 544.950 445.050 547.050 ;
        RECT 443.400 541.050 444.600 544.950 ;
        RECT 442.950 538.950 445.050 541.050 ;
        RECT 448.950 535.950 451.050 538.050 ;
        RECT 449.400 532.050 450.600 535.950 ;
        RECT 442.950 529.950 445.050 532.050 ;
        RECT 448.950 529.950 451.050 532.050 ;
        RECT 461.400 531.600 462.600 547.950 ;
        RECT 463.950 544.950 466.050 547.050 ;
        RECT 464.400 541.050 465.600 544.950 ;
        RECT 463.950 538.950 466.050 541.050 ;
        RECT 467.400 538.050 468.600 571.950 ;
        RECT 470.400 547.200 471.600 571.950 ;
        RECT 476.400 565.050 477.600 598.950 ;
        RECT 482.400 588.600 483.600 646.950 ;
        RECT 484.950 631.950 487.050 634.050 ;
        RECT 485.400 619.050 486.600 631.950 ;
        RECT 491.400 631.050 492.600 667.950 ;
        RECT 494.400 661.050 495.600 703.950 ;
        RECT 506.400 703.050 507.600 709.950 ;
        RECT 505.950 700.950 508.050 703.050 ;
        RECT 496.950 697.950 499.050 700.050 ;
        RECT 497.400 673.050 498.600 697.950 ;
        RECT 512.400 694.050 513.600 739.950 ;
        RECT 517.950 736.950 520.050 739.050 ;
        RECT 518.400 721.050 519.600 736.950 ;
        RECT 527.400 736.050 528.600 754.950 ;
        RECT 526.950 733.950 529.050 736.050 ;
        RECT 529.950 721.950 532.050 724.050 ;
        RECT 517.950 718.950 520.050 721.050 ;
        RECT 523.950 718.950 526.050 721.050 ;
        RECT 524.400 715.200 525.600 718.950 ;
        RECT 523.950 713.100 526.050 715.200 ;
        RECT 523.950 709.800 526.050 711.900 ;
        RECT 520.950 706.950 523.050 709.050 ;
        RECT 521.400 700.050 522.600 706.950 ;
        RECT 524.400 700.050 525.600 709.800 ;
        RECT 530.400 703.050 531.600 721.950 ;
        RECT 529.950 700.950 532.050 703.050 ;
        RECT 533.400 700.050 534.600 769.950 ;
        RECT 548.400 766.050 549.600 772.950 ;
        RECT 551.400 772.050 552.600 784.950 ;
        RECT 550.950 769.950 553.050 772.050 ;
        RECT 557.400 766.050 558.600 784.950 ;
        RECT 571.950 784.800 574.050 786.900 ;
        RECT 559.950 769.950 562.050 772.050 ;
        RECT 535.950 763.950 538.050 766.050 ;
        RECT 544.950 763.950 547.050 766.050 ;
        RECT 547.950 763.950 550.050 766.050 ;
        RECT 553.950 764.400 558.600 766.050 ;
        RECT 553.950 763.950 558.000 764.400 ;
        RECT 520.800 697.950 522.900 700.050 ;
        RECT 524.100 697.950 526.200 700.050 ;
        RECT 532.950 697.950 535.050 700.050 ;
        RECT 511.950 693.600 514.050 694.050 ;
        RECT 509.400 692.400 514.050 693.600 ;
        RECT 499.950 676.950 502.050 679.050 ;
        RECT 496.950 670.950 499.050 673.050 ;
        RECT 500.400 667.050 501.600 676.950 ;
        RECT 499.950 664.950 502.050 667.050 ;
        RECT 496.800 661.950 498.900 664.050 ;
        RECT 493.950 658.950 496.050 661.050 ;
        RECT 497.400 652.050 498.600 661.950 ;
        RECT 509.400 658.050 510.600 692.400 ;
        RECT 511.950 691.950 514.050 692.400 ;
        RECT 520.950 691.950 523.050 694.050 ;
        RECT 529.950 691.950 532.050 694.050 ;
        RECT 521.400 688.050 522.600 691.950 ;
        RECT 520.950 685.950 523.050 688.050 ;
        RECT 530.400 682.050 531.600 691.950 ;
        RECT 529.950 679.950 532.050 682.050 ;
        RECT 517.950 676.950 520.050 679.050 ;
        RECT 536.400 678.600 537.600 763.950 ;
        RECT 538.950 754.950 541.050 757.050 ;
        RECT 539.400 706.050 540.600 754.950 ;
        RECT 545.400 751.050 546.600 763.950 ;
        RECT 550.950 756.600 555.000 757.050 ;
        RECT 550.950 756.000 555.600 756.600 ;
        RECT 550.950 754.950 556.050 756.000 ;
        RECT 553.950 751.950 556.050 754.950 ;
        RECT 544.950 748.950 547.050 751.050 ;
        RECT 553.950 721.950 556.050 724.050 ;
        RECT 550.950 712.950 553.050 715.050 ;
        RECT 544.950 706.950 547.050 709.050 ;
        RECT 539.400 703.950 544.050 706.050 ;
        RECT 539.400 688.050 540.600 703.950 ;
        RECT 545.400 688.050 546.600 706.950 ;
        RECT 551.400 694.050 552.600 712.950 ;
        RECT 554.400 700.050 555.600 721.950 ;
        RECT 560.400 712.050 561.600 769.950 ;
        RECT 572.400 766.050 573.600 784.800 ;
        RECT 589.950 781.950 592.050 784.050 ;
        RECT 565.950 765.600 570.000 766.050 ;
        RECT 565.950 763.950 570.600 765.600 ;
        RECT 571.950 763.950 574.050 766.050 ;
        RECT 569.400 762.600 570.600 763.950 ;
        RECT 569.400 761.400 582.600 762.600 ;
        RECT 581.400 757.050 582.600 761.400 ;
        RECT 568.950 754.950 571.050 757.050 ;
        RECT 577.800 754.950 579.900 757.050 ;
        RECT 581.100 754.950 583.200 757.050 ;
        RECT 569.400 751.050 570.600 754.950 ;
        RECT 568.950 748.950 571.050 751.050 ;
        RECT 578.400 748.050 579.600 754.950 ;
        RECT 587.100 748.950 589.200 751.050 ;
        RECT 577.950 745.950 580.050 748.050 ;
        RECT 587.400 735.600 588.600 748.950 ;
        RECT 590.400 742.050 591.600 781.950 ;
        RECT 593.400 766.050 594.600 797.400 ;
        RECT 598.950 796.950 601.050 797.400 ;
        RECT 604.950 797.400 609.600 799.050 ;
        RECT 604.950 796.950 609.000 797.400 ;
        RECT 611.400 784.050 612.600 811.950 ;
        RECT 616.950 805.950 619.050 808.050 ;
        RECT 617.400 784.050 618.600 805.950 ;
        RECT 623.400 799.050 624.600 814.950 ;
        RECT 626.400 814.050 627.600 865.950 ;
        RECT 625.950 811.950 628.050 814.050 ;
        RECT 629.400 811.050 630.600 868.950 ;
        RECT 635.400 868.200 636.600 871.950 ;
        RECT 634.950 866.100 637.050 868.200 ;
        RECT 641.400 868.050 642.600 874.950 ;
        RECT 644.400 871.050 645.600 877.950 ;
        RECT 643.950 868.950 646.050 871.050 ;
        RECT 640.950 865.950 643.050 868.050 ;
        RECT 634.950 862.800 637.050 864.900 ;
        RECT 631.950 847.950 634.050 850.050 ;
        RECT 632.400 831.600 633.600 847.950 ;
        RECT 635.400 835.050 636.600 862.800 ;
        RECT 644.400 859.050 645.600 868.950 ;
        RECT 643.950 856.950 646.050 859.050 ;
        RECT 644.400 841.050 645.600 856.950 ;
        RECT 655.950 847.950 658.050 850.050 ;
        RECT 637.950 838.950 640.050 841.050 ;
        RECT 643.950 838.950 646.050 841.050 ;
        RECT 634.950 832.950 637.050 835.050 ;
        RECT 632.400 830.400 636.600 831.600 ;
        RECT 631.950 826.950 634.050 829.050 ;
        RECT 628.950 808.950 631.050 811.050 ;
        RECT 625.950 807.600 628.050 808.050 ;
        RECT 632.400 807.600 633.600 826.950 ;
        RECT 625.950 806.400 633.600 807.600 ;
        RECT 625.950 805.950 628.050 806.400 ;
        RECT 635.400 802.200 636.600 830.400 ;
        RECT 634.950 800.100 637.050 802.200 ;
        RECT 622.950 796.950 625.050 799.050 ;
        RECT 628.950 798.600 631.050 799.050 ;
        RECT 634.950 798.600 637.050 798.900 ;
        RECT 628.950 797.400 637.050 798.600 ;
        RECT 628.950 796.950 631.050 797.400 ;
        RECT 634.950 796.800 637.050 797.400 ;
        RECT 638.400 793.050 639.600 838.950 ;
        RECT 656.400 835.050 657.600 847.950 ;
        RECT 659.400 844.050 660.600 877.950 ;
        RECT 685.950 874.950 688.050 877.050 ;
        RECT 670.950 871.950 673.050 874.050 ;
        RECT 671.400 859.050 672.600 871.950 ;
        RECT 679.950 865.950 682.050 868.050 ;
        RECT 670.950 856.950 673.050 859.050 ;
        RECT 661.950 847.950 664.050 850.050 ;
        RECT 658.950 841.950 661.050 844.050 ;
        RECT 655.950 832.950 658.050 835.050 ;
        RECT 649.950 826.950 652.050 829.050 ;
        RECT 646.950 811.950 649.050 814.050 ;
        RECT 640.950 805.950 643.050 808.050 ;
        RECT 637.950 790.950 640.050 793.050 ;
        RECT 598.950 781.950 601.050 784.050 ;
        RECT 610.950 781.950 613.050 784.050 ;
        RECT 616.950 781.950 619.050 784.050 ;
        RECT 628.950 781.950 631.050 784.050 ;
        RECT 599.400 766.050 600.600 781.950 ;
        RECT 610.950 772.950 613.050 775.050 ;
        RECT 592.950 763.950 595.050 766.050 ;
        RECT 598.950 763.950 601.050 766.050 ;
        RECT 601.950 751.950 604.050 754.050 ;
        RECT 595.950 745.950 598.050 748.050 ;
        RECT 589.950 739.950 592.050 742.050 ;
        RECT 584.400 734.400 588.600 735.600 ;
        RECT 584.400 724.050 585.600 734.400 ;
        RECT 574.950 723.600 577.050 724.050 ;
        RECT 569.400 722.400 577.050 723.600 ;
        RECT 569.400 715.050 570.600 722.400 ;
        RECT 574.950 721.950 577.050 722.400 ;
        RECT 583.950 721.950 586.050 724.050 ;
        RECT 596.400 721.050 597.600 745.950 ;
        RECT 602.400 736.050 603.600 751.950 ;
        RECT 601.800 733.950 603.900 736.050 ;
        RECT 611.400 730.050 612.600 772.950 ;
        RECT 613.950 769.950 616.050 772.050 ;
        RECT 614.400 757.050 615.600 769.950 ;
        RECT 616.950 763.950 619.050 766.050 ;
        RECT 622.950 763.950 625.050 766.050 ;
        RECT 613.950 754.950 616.050 757.050 ;
        RECT 617.400 751.050 618.600 763.950 ;
        RECT 623.400 751.050 624.600 763.950 ;
        RECT 616.950 748.950 619.050 751.050 ;
        RECT 622.950 748.950 625.050 751.050 ;
        RECT 629.400 750.600 630.600 781.950 ;
        RECT 641.400 775.200 642.600 805.950 ;
        RECT 647.400 799.050 648.600 811.950 ;
        RECT 650.400 808.050 651.600 826.950 ;
        RECT 658.950 823.950 661.050 826.050 ;
        RECT 655.950 814.950 658.050 817.050 ;
        RECT 649.950 805.950 652.050 808.050 ;
        RECT 656.400 799.050 657.600 814.950 ;
        RECT 646.950 796.950 649.050 799.050 ;
        RECT 652.950 797.400 657.600 799.050 ;
        RECT 652.950 796.950 657.000 797.400 ;
        RECT 649.950 787.950 652.050 790.050 ;
        RECT 640.950 773.100 643.050 775.200 ;
        RECT 640.950 769.800 643.050 771.900 ;
        RECT 641.400 766.050 642.600 769.800 ;
        RECT 636.000 765.600 640.050 766.050 ;
        RECT 635.400 763.950 640.050 765.600 ;
        RECT 641.400 764.400 646.050 766.050 ;
        RECT 642.000 763.950 646.050 764.400 ;
        RECT 635.400 757.050 636.600 763.950 ;
        RECT 634.950 754.950 637.050 757.050 ;
        RECT 640.950 754.950 643.050 757.050 ;
        RECT 645.000 756.600 649.050 757.050 ;
        RECT 644.400 754.950 649.050 756.600 ;
        RECT 629.400 749.400 633.600 750.600 ;
        RECT 619.950 739.950 622.050 742.050 ;
        RECT 598.950 729.600 601.050 730.050 ;
        RECT 604.950 729.600 607.050 730.050 ;
        RECT 598.950 728.400 607.050 729.600 ;
        RECT 598.950 727.950 601.050 728.400 ;
        RECT 604.950 727.950 607.050 728.400 ;
        RECT 610.950 727.950 613.050 730.050 ;
        RECT 620.400 721.050 621.600 739.950 ;
        RECT 589.950 718.950 592.050 721.050 ;
        RECT 595.950 718.950 598.050 721.050 ;
        RECT 607.950 720.600 610.050 721.050 ;
        RECT 613.950 720.600 616.050 721.050 ;
        RECT 607.950 719.400 616.050 720.600 ;
        RECT 607.950 718.950 610.050 719.400 ;
        RECT 613.950 718.950 616.050 719.400 ;
        RECT 619.950 718.950 622.050 721.050 ;
        RECT 568.950 712.950 571.050 715.050 ;
        RECT 590.400 712.050 591.600 718.950 ;
        RECT 607.950 712.950 610.050 715.050 ;
        RECT 613.950 712.950 616.050 715.050 ;
        RECT 559.950 709.950 562.050 712.050 ;
        RECT 577.950 709.950 580.050 712.050 ;
        RECT 589.950 709.950 592.050 712.050 ;
        RECT 568.950 703.950 571.050 706.050 ;
        RECT 553.950 697.950 556.050 700.050 ;
        RECT 559.950 696.600 562.050 700.050 ;
        RECT 557.400 696.000 562.050 696.600 ;
        RECT 557.400 695.400 561.600 696.000 ;
        RECT 550.950 691.950 553.050 694.050 ;
        RECT 557.400 688.050 558.600 695.400 ;
        RECT 538.950 685.950 541.050 688.050 ;
        RECT 544.950 685.950 547.050 688.050 ;
        RECT 550.950 685.950 553.050 688.050 ;
        RECT 556.950 685.950 559.050 688.050 ;
        RECT 562.950 687.600 565.050 688.050 ;
        RECT 569.400 687.600 570.600 703.950 ;
        RECT 578.400 690.600 579.600 709.950 ;
        RECT 592.800 706.950 594.900 709.050 ;
        RECT 596.100 706.950 598.200 709.050 ;
        RECT 586.950 700.950 589.050 703.050 ;
        RECT 587.400 697.050 588.600 700.950 ;
        RECT 586.950 694.950 589.050 697.050 ;
        RECT 578.400 689.400 585.600 690.600 ;
        RECT 584.400 688.050 585.600 689.400 ;
        RECT 562.950 686.400 570.600 687.600 ;
        RECT 574.950 687.600 577.050 688.050 ;
        RECT 580.950 687.600 583.050 688.050 ;
        RECT 574.950 686.400 583.050 687.600 ;
        RECT 584.400 686.400 589.050 688.050 ;
        RECT 562.950 685.950 565.050 686.400 ;
        RECT 574.950 685.950 577.050 686.400 ;
        RECT 580.950 685.950 583.050 686.400 ;
        RECT 585.000 685.950 589.050 686.400 ;
        RECT 533.400 677.400 537.600 678.600 ;
        RECT 518.400 670.050 519.600 676.950 ;
        RECT 533.400 673.050 534.600 677.400 ;
        RECT 541.950 676.950 544.050 679.050 ;
        RECT 535.950 673.950 538.050 676.050 ;
        RECT 527.100 670.950 529.200 673.050 ;
        RECT 532.950 670.950 535.050 673.050 ;
        RECT 517.950 667.950 520.050 670.050 ;
        RECT 511.950 664.950 514.050 667.050 ;
        RECT 508.950 655.950 511.050 658.050 ;
        RECT 512.400 652.050 513.600 664.950 ;
        RECT 517.950 658.950 520.050 661.050 ;
        RECT 518.400 652.050 519.600 658.950 ;
        RECT 493.950 650.400 498.600 652.050 ;
        RECT 493.950 649.950 498.000 650.400 ;
        RECT 511.950 649.950 514.050 652.050 ;
        RECT 517.950 649.950 520.050 652.050 ;
        RECT 508.950 640.950 511.050 643.050 ;
        RECT 514.950 640.950 517.050 643.050 ;
        RECT 509.400 637.050 510.600 640.950 ;
        RECT 502.950 634.950 505.050 637.050 ;
        RECT 508.950 634.950 511.050 637.050 ;
        RECT 490.950 628.950 493.050 631.050 ;
        RECT 503.400 628.050 504.600 634.950 ;
        RECT 502.800 625.950 504.900 628.050 ;
        RECT 506.100 625.950 508.200 628.050 ;
        RECT 506.400 622.050 507.600 625.950 ;
        RECT 515.400 625.050 516.600 640.950 ;
        RECT 518.400 625.050 519.600 649.950 ;
        RECT 523.950 643.950 526.050 646.050 ;
        RECT 524.400 628.050 525.600 643.950 ;
        RECT 527.400 631.050 528.600 670.950 ;
        RECT 529.950 666.600 534.000 667.050 ;
        RECT 529.950 664.950 534.600 666.600 ;
        RECT 533.400 646.050 534.600 664.950 ;
        RECT 532.950 643.950 535.050 646.050 ;
        RECT 526.950 628.950 529.050 631.050 ;
        RECT 536.400 628.050 537.600 673.950 ;
        RECT 542.400 670.050 543.600 676.950 ;
        RECT 544.950 670.950 547.050 673.050 ;
        RECT 541.950 667.950 544.050 670.050 ;
        RECT 523.950 625.950 526.050 628.050 ;
        RECT 529.950 625.950 532.050 628.050 ;
        RECT 535.950 625.950 538.050 628.050 ;
        RECT 514.800 622.950 516.900 625.050 ;
        RECT 518.100 622.950 520.200 625.050 ;
        RECT 496.950 619.950 499.050 622.050 ;
        RECT 505.950 619.950 508.050 622.050 ;
        RECT 520.950 619.950 523.050 622.050 ;
        RECT 484.950 616.950 487.050 619.050 ;
        RECT 497.400 610.050 498.600 619.950 ;
        RECT 499.950 616.950 502.050 619.050 ;
        RECT 489.000 609.600 493.050 610.050 ;
        RECT 488.400 607.950 493.050 609.600 ;
        RECT 496.950 607.950 499.050 610.050 ;
        RECT 488.400 589.050 489.600 607.950 ;
        RECT 500.400 601.050 501.600 616.950 ;
        RECT 506.400 607.050 507.600 619.950 ;
        RECT 505.950 604.950 508.050 607.050 ;
        RECT 514.950 604.950 517.050 607.050 ;
        RECT 493.950 598.950 496.050 601.050 ;
        RECT 499.950 598.950 502.050 601.050 ;
        RECT 494.400 595.050 495.600 598.950 ;
        RECT 515.400 597.600 516.600 604.950 ;
        RECT 509.400 596.400 516.600 597.600 ;
        RECT 493.950 592.950 496.050 595.050 ;
        RECT 502.950 594.600 505.050 595.050 ;
        RECT 509.400 594.600 510.600 596.400 ;
        RECT 502.950 593.400 510.600 594.600 ;
        RECT 502.950 592.950 505.050 593.400 ;
        RECT 482.400 587.400 486.600 588.600 ;
        RECT 481.950 583.950 484.050 586.050 ;
        RECT 482.400 565.050 483.600 583.950 ;
        RECT 485.400 580.050 486.600 587.400 ;
        RECT 487.950 586.950 490.050 589.050 ;
        RECT 496.950 580.950 499.050 583.050 ;
        RECT 514.950 580.950 517.050 583.050 ;
        RECT 484.950 577.950 487.050 580.050 ;
        RECT 497.400 574.050 498.600 580.950 ;
        RECT 505.950 577.950 508.050 580.050 ;
        RECT 484.950 573.600 487.050 574.050 ;
        RECT 490.950 573.600 493.050 574.050 ;
        RECT 484.950 572.400 493.050 573.600 ;
        RECT 484.950 571.950 487.050 572.400 ;
        RECT 490.950 571.950 493.050 572.400 ;
        RECT 496.950 571.950 499.050 574.050 ;
        RECT 506.400 565.050 507.600 577.950 ;
        RECT 515.400 574.050 516.600 580.950 ;
        RECT 515.100 571.950 517.200 574.050 ;
        RECT 475.950 562.950 478.050 565.050 ;
        RECT 481.950 562.950 484.050 565.050 ;
        RECT 498.000 564.600 502.050 565.050 ;
        RECT 497.400 564.000 502.050 564.600 ;
        RECT 496.950 562.950 502.050 564.000 ;
        RECT 505.950 562.950 508.050 565.050 ;
        RECT 517.950 562.950 520.050 565.050 ;
        RECT 496.950 559.950 499.050 562.950 ;
        RECT 502.950 550.950 505.050 553.050 ;
        RECT 469.950 545.100 472.050 547.200 ;
        RECT 478.950 544.950 481.050 547.050 ;
        RECT 496.950 544.950 499.050 547.050 ;
        RECT 469.950 541.800 472.050 543.900 ;
        RECT 466.950 535.950 469.050 538.050 ;
        RECT 466.950 531.600 469.050 532.050 ;
        RECT 461.400 530.400 469.050 531.600 ;
        RECT 466.950 529.950 469.050 530.400 ;
        RECT 430.950 520.950 433.050 523.050 ;
        RECT 431.400 511.050 432.600 520.950 ;
        RECT 443.400 517.050 444.600 529.950 ;
        RECT 470.400 523.050 471.600 541.800 ;
        RECT 472.950 538.950 475.050 541.050 ;
        RECT 473.400 532.050 474.600 538.950 ;
        RECT 472.950 529.950 475.050 532.050 ;
        RECT 445.950 520.950 448.050 523.050 ;
        RECT 469.950 520.950 472.050 523.050 ;
        RECT 442.950 514.950 445.050 517.050 ;
        RECT 446.400 511.050 447.600 520.950 ;
        RECT 454.800 511.950 456.900 514.050 ;
        RECT 430.950 508.950 433.050 511.050 ;
        RECT 445.950 508.950 448.050 511.050 ;
        RECT 431.400 505.050 432.600 508.950 ;
        RECT 430.950 502.950 433.050 505.050 ;
        RECT 455.400 496.050 456.600 511.950 ;
        RECT 469.950 505.950 472.050 508.050 ;
        RECT 470.400 496.050 471.600 505.950 ;
        RECT 479.400 505.050 480.600 544.950 ;
        RECT 484.950 541.950 487.050 544.050 ;
        RECT 485.400 532.050 486.600 541.950 ;
        RECT 490.950 538.950 493.050 541.050 ;
        RECT 484.950 529.950 487.050 532.050 ;
        RECT 491.400 523.050 492.600 538.950 ;
        RECT 497.400 532.050 498.600 544.950 ;
        RECT 496.950 529.950 499.050 532.050 ;
        RECT 491.400 521.400 496.050 523.050 ;
        RECT 492.000 520.950 496.050 521.400 ;
        RECT 487.950 517.950 490.050 520.050 ;
        RECT 478.950 502.950 481.050 505.050 ;
        RECT 488.400 502.050 489.600 517.950 ;
        RECT 496.950 514.950 499.050 517.050 ;
        RECT 487.950 499.950 490.050 502.050 ;
        RECT 439.950 493.950 442.050 496.050 ;
        RECT 454.950 493.950 457.050 496.050 ;
        RECT 469.950 493.950 472.050 496.050 ;
        RECT 484.800 493.950 486.900 496.050 ;
        RECT 430.950 484.950 433.050 487.050 ;
        RECT 431.400 481.050 432.600 484.950 ;
        RECT 430.950 478.950 433.050 481.050 ;
        RECT 409.950 472.950 412.050 475.050 ;
        RECT 427.950 472.950 430.050 475.050 ;
        RECT 403.950 469.950 406.050 472.050 ;
        RECT 400.950 457.950 403.050 460.050 ;
        RECT 404.400 454.050 405.600 469.950 ;
        RECT 400.950 452.400 405.600 454.050 ;
        RECT 400.950 451.950 405.000 452.400 ;
        RECT 400.950 442.950 403.050 445.050 ;
        RECT 397.950 424.950 400.050 427.050 ;
        RECT 355.950 421.950 358.050 424.050 ;
        RECT 376.950 421.950 379.050 424.050 ;
        RECT 241.950 417.600 244.050 418.050 ;
        RECT 247.950 417.600 250.050 418.050 ;
        RECT 241.950 416.400 250.050 417.600 ;
        RECT 241.950 415.950 244.050 416.400 ;
        RECT 247.950 415.950 250.050 416.400 ;
        RECT 256.950 416.400 261.600 418.050 ;
        RECT 316.950 417.600 319.050 418.050 ;
        RECT 311.400 416.400 319.050 417.600 ;
        RECT 256.950 415.950 261.000 416.400 ;
        RECT 311.400 412.050 312.600 416.400 ;
        RECT 316.950 415.950 319.050 416.400 ;
        RECT 334.950 415.950 337.050 418.050 ;
        RECT 343.950 415.950 346.050 418.050 ;
        RECT 289.950 409.950 292.050 412.050 ;
        RECT 310.950 409.950 313.050 412.050 ;
        RECT 259.950 406.950 262.050 409.050 ;
        RECT 244.950 397.950 247.050 400.050 ;
        RECT 245.400 355.050 246.600 397.950 ;
        RECT 260.400 394.050 261.600 406.950 ;
        RECT 247.950 391.950 250.050 394.050 ;
        RECT 259.950 391.950 262.050 394.050 ;
        RECT 248.400 379.050 249.600 391.950 ;
        RECT 274.950 379.950 277.050 382.050 ;
        RECT 280.950 379.950 283.050 382.050 ;
        RECT 247.950 376.950 250.050 379.050 ;
        RECT 248.400 364.050 249.600 376.950 ;
        RECT 275.400 373.050 276.600 379.950 ;
        RECT 281.400 376.050 282.600 379.950 ;
        RECT 290.400 376.050 291.600 409.950 ;
        RECT 313.950 406.950 316.050 409.050 ;
        RECT 298.950 403.950 301.050 406.050 ;
        RECT 280.950 373.950 283.050 376.050 ;
        RECT 286.950 374.400 291.600 376.050 ;
        RECT 299.400 376.050 300.600 403.950 ;
        RECT 299.400 374.400 304.050 376.050 ;
        RECT 286.950 373.950 291.000 374.400 ;
        RECT 300.000 373.950 304.050 374.400 ;
        RECT 307.950 375.600 310.050 376.050 ;
        RECT 314.400 375.600 315.600 406.950 ;
        RECT 335.400 400.050 336.600 415.950 ;
        RECT 352.950 408.600 355.050 412.050 ;
        RECT 356.400 408.600 357.600 421.950 ;
        RECT 370.950 415.950 373.050 418.050 ;
        RECT 358.950 408.600 361.050 409.050 ;
        RECT 352.950 408.000 361.050 408.600 ;
        RECT 353.400 407.400 361.050 408.000 ;
        RECT 358.950 406.950 361.050 407.400 ;
        RECT 364.950 406.950 367.050 409.050 ;
        RECT 334.950 397.950 337.050 400.050 ;
        RECT 322.950 394.950 325.050 397.050 ;
        RECT 331.950 394.950 334.050 397.050 ;
        RECT 323.400 376.050 324.600 394.950 ;
        RECT 307.950 374.400 315.600 375.600 ;
        RECT 307.950 373.950 310.050 374.400 ;
        RECT 256.950 370.950 259.050 373.050 ;
        RECT 274.950 370.950 277.050 373.050 ;
        RECT 316.950 372.600 319.050 376.050 ;
        RECT 322.950 373.950 325.050 376.050 ;
        RECT 327.000 375.600 331.050 376.050 ;
        RECT 326.400 373.950 331.050 375.600 ;
        RECT 326.400 372.600 327.600 373.950 ;
        RECT 316.950 372.000 327.600 372.600 ;
        RECT 317.400 371.400 327.600 372.000 ;
        RECT 257.400 364.050 258.600 370.950 ;
        RECT 268.950 369.600 271.050 370.050 ;
        RECT 260.400 368.400 271.050 369.600 ;
        RECT 260.400 364.050 261.600 368.400 ;
        RECT 268.950 367.950 271.050 368.400 ;
        RECT 277.950 366.600 280.050 370.050 ;
        RECT 298.950 366.600 301.050 367.050 ;
        RECT 277.950 366.000 301.050 366.600 ;
        RECT 278.400 365.400 301.050 366.000 ;
        RECT 298.950 364.950 301.050 365.400 ;
        RECT 247.950 361.950 250.050 364.050 ;
        RECT 257.400 362.400 262.050 364.050 ;
        RECT 258.000 361.950 262.050 362.400 ;
        RECT 265.950 361.950 268.050 364.050 ;
        RECT 325.950 361.950 328.050 364.050 ;
        RECT 266.400 358.050 267.600 361.950 ;
        RECT 271.950 358.950 274.050 361.050 ;
        RECT 265.950 355.950 268.050 358.050 ;
        RECT 244.950 352.950 247.050 355.050 ;
        RECT 272.400 352.050 273.600 358.950 ;
        RECT 295.950 352.950 298.050 355.050 ;
        RECT 271.950 349.950 274.050 352.050 ;
        RECT 238.950 346.950 241.050 349.050 ;
        RECT 296.400 346.050 297.600 352.950 ;
        RECT 244.950 343.950 247.050 346.050 ;
        RECT 262.950 343.950 265.050 346.050 ;
        RECT 295.950 343.950 298.050 346.050 ;
        RECT 316.950 343.950 319.050 346.050 ;
        RECT 245.400 340.050 246.600 343.950 ;
        RECT 263.400 340.050 264.600 343.950 ;
        RECT 237.000 339.600 241.050 340.050 ;
        RECT 236.400 337.950 241.050 339.600 ;
        RECT 244.950 337.950 247.050 340.050 ;
        RECT 262.950 337.950 265.050 340.050 ;
        RECT 236.400 325.050 237.600 337.950 ;
        RECT 271.950 336.600 274.050 340.050 ;
        RECT 269.400 336.000 274.050 336.600 ;
        RECT 269.400 335.400 273.600 336.000 ;
        RECT 240.000 330.600 244.050 331.050 ;
        RECT 239.400 330.000 244.050 330.600 ;
        RECT 238.950 328.950 244.050 330.000 ;
        RECT 247.950 330.600 250.050 331.050 ;
        RECT 253.950 330.600 256.050 331.050 ;
        RECT 247.950 329.400 256.050 330.600 ;
        RECT 247.950 328.950 250.050 329.400 ;
        RECT 253.950 328.950 256.050 329.400 ;
        RECT 262.950 330.600 265.050 331.050 ;
        RECT 269.400 330.600 270.600 335.400 ;
        RECT 271.950 331.950 274.050 334.050 ;
        RECT 262.950 329.400 270.600 330.600 ;
        RECT 262.950 328.950 265.050 329.400 ;
        RECT 238.950 325.950 241.050 328.950 ;
        RECT 272.400 325.050 273.600 331.950 ;
        RECT 283.950 328.950 286.050 331.050 ;
        RECT 289.950 328.950 292.050 331.050 ;
        RECT 284.400 325.050 285.600 328.950 ;
        RECT 290.400 325.050 291.600 328.950 ;
        RECT 235.950 322.950 238.050 325.050 ;
        RECT 271.950 322.950 274.050 325.050 ;
        RECT 283.950 322.950 286.050 325.050 ;
        RECT 289.950 322.950 292.050 325.050 ;
        RECT 229.950 313.950 232.050 316.050 ;
        RECT 232.950 310.950 235.050 313.050 ;
        RECT 220.950 307.950 223.050 310.050 ;
        RECT 221.400 298.050 222.600 307.950 ;
        RECT 220.950 295.950 223.050 298.050 ;
        RECT 226.950 297.600 231.000 298.050 ;
        RECT 226.950 295.950 231.600 297.600 ;
        RECT 230.400 286.050 231.600 295.950 ;
        RECT 233.400 289.050 234.600 310.950 ;
        RECT 232.950 286.950 235.050 289.050 ;
        RECT 229.950 283.950 232.050 286.050 ;
        RECT 229.950 265.950 232.050 268.050 ;
        RECT 220.950 259.950 223.050 262.050 ;
        RECT 217.950 250.950 220.050 253.050 ;
        RECT 212.400 230.400 216.600 231.600 ;
        RECT 208.950 199.950 211.050 202.050 ;
        RECT 205.950 196.950 208.050 199.050 ;
        RECT 215.400 193.050 216.600 230.400 ;
        RECT 214.950 190.950 217.050 193.050 ;
        RECT 205.950 175.950 208.050 178.050 ;
        RECT 206.400 160.050 207.600 175.950 ;
        RECT 214.950 163.950 217.050 166.050 ;
        RECT 205.950 157.950 208.050 160.050 ;
        RECT 215.400 142.050 216.600 163.950 ;
        RECT 214.950 139.950 217.050 142.050 ;
        RECT 211.950 130.950 214.050 133.050 ;
        RECT 212.400 121.050 213.600 130.950 ;
        RECT 211.950 118.950 214.050 121.050 ;
        RECT 218.400 115.050 219.600 250.950 ;
        RECT 221.400 238.050 222.600 259.950 ;
        RECT 230.400 253.050 231.600 265.950 ;
        RECT 236.400 253.050 237.600 322.950 ;
        RECT 296.400 321.600 297.600 343.950 ;
        RECT 317.400 340.050 318.600 343.950 ;
        RECT 313.950 338.400 318.600 340.050 ;
        RECT 313.950 337.950 318.000 338.400 ;
        RECT 310.950 331.950 313.050 334.050 ;
        RECT 316.950 331.950 319.050 334.050 ;
        RECT 293.400 320.400 297.600 321.600 ;
        RECT 241.950 310.950 244.050 313.050 ;
        RECT 242.400 280.050 243.600 310.950 ;
        RECT 265.950 300.600 268.050 301.050 ;
        RECT 254.400 299.400 268.050 300.600 ;
        RECT 254.400 295.050 255.600 299.400 ;
        RECT 265.950 298.950 268.050 299.400 ;
        RECT 274.950 300.600 277.050 301.050 ;
        RECT 283.950 300.600 286.050 301.050 ;
        RECT 274.950 299.400 286.050 300.600 ;
        RECT 274.950 298.950 277.050 299.400 ;
        RECT 283.950 298.950 286.050 299.400 ;
        RECT 253.950 292.950 256.050 295.050 ;
        RECT 274.950 292.950 277.050 295.050 ;
        RECT 256.950 288.600 259.050 289.050 ;
        RECT 245.400 288.000 259.050 288.600 ;
        RECT 244.950 287.400 259.050 288.000 ;
        RECT 244.950 283.950 247.050 287.400 ;
        RECT 256.950 286.950 259.050 287.400 ;
        RECT 250.950 283.950 253.050 286.050 ;
        RECT 251.400 280.050 252.600 283.950 ;
        RECT 241.950 277.950 244.050 280.050 ;
        RECT 250.950 277.950 253.050 280.050 ;
        RECT 251.400 271.050 252.600 277.950 ;
        RECT 265.950 274.950 268.050 277.050 ;
        RECT 250.950 268.950 253.050 271.050 ;
        RECT 259.950 268.950 262.050 271.050 ;
        RECT 229.950 250.950 232.050 253.050 ;
        RECT 235.950 250.950 238.050 253.050 ;
        RECT 241.950 252.600 244.050 253.050 ;
        RECT 247.950 252.600 250.050 253.050 ;
        RECT 241.950 251.400 250.050 252.600 ;
        RECT 241.950 250.950 244.050 251.400 ;
        RECT 247.950 250.950 250.050 251.400 ;
        RECT 253.950 250.950 256.050 253.050 ;
        RECT 254.400 247.050 255.600 250.950 ;
        RECT 253.950 244.950 256.050 247.050 ;
        RECT 260.400 244.050 261.600 268.950 ;
        RECT 259.950 241.950 262.050 244.050 ;
        RECT 220.950 235.950 223.050 238.050 ;
        RECT 232.950 229.950 235.050 232.050 ;
        RECT 250.950 229.950 253.050 232.050 ;
        RECT 223.950 217.950 226.050 220.050 ;
        RECT 224.400 196.050 225.600 217.950 ;
        RECT 233.400 211.050 234.600 229.950 ;
        RECT 247.950 223.950 250.050 226.050 ;
        RECT 248.400 220.050 249.600 223.950 ;
        RECT 241.950 217.950 244.050 220.050 ;
        RECT 247.950 217.950 250.050 220.050 ;
        RECT 226.950 208.950 229.050 211.050 ;
        RECT 232.950 208.950 235.050 211.050 ;
        RECT 227.400 202.050 228.600 208.950 ;
        RECT 242.400 205.050 243.600 217.950 ;
        RECT 251.400 211.050 252.600 229.950 ;
        RECT 260.400 211.050 261.600 241.950 ;
        RECT 262.950 238.950 265.050 241.050 ;
        RECT 263.400 223.050 264.600 238.950 ;
        RECT 266.400 229.050 267.600 274.950 ;
        RECT 275.400 271.050 276.600 292.950 ;
        RECT 283.950 291.600 286.050 295.050 ;
        RECT 283.950 291.000 288.600 291.600 ;
        RECT 284.400 290.400 288.600 291.000 ;
        RECT 283.950 283.950 286.050 286.050 ;
        RECT 284.400 273.600 285.600 283.950 ;
        RECT 287.400 280.050 288.600 290.400 ;
        RECT 286.950 277.950 289.050 280.050 ;
        RECT 287.400 274.050 288.600 277.950 ;
        RECT 293.400 277.050 294.600 320.400 ;
        RECT 311.400 319.050 312.600 331.950 ;
        RECT 310.950 316.950 313.050 319.050 ;
        RECT 317.400 313.050 318.600 331.950 ;
        RECT 319.950 316.950 322.050 319.050 ;
        RECT 316.950 310.950 319.050 313.050 ;
        RECT 298.950 297.600 301.050 301.050 ;
        RECT 304.950 297.600 307.050 298.050 ;
        RECT 298.950 297.000 307.050 297.600 ;
        RECT 299.400 296.400 307.050 297.000 ;
        RECT 304.950 295.950 307.050 296.400 ;
        RECT 310.950 297.600 313.050 298.050 ;
        RECT 317.400 297.600 318.600 310.950 ;
        RECT 310.950 296.400 318.600 297.600 ;
        RECT 310.950 295.950 313.050 296.400 ;
        RECT 295.950 286.950 298.050 289.050 ;
        RECT 307.950 288.600 312.000 289.050 ;
        RECT 307.950 286.950 312.600 288.600 ;
        RECT 292.950 274.950 295.050 277.050 ;
        RECT 281.400 272.400 285.600 273.600 ;
        RECT 274.950 268.950 277.050 271.050 ;
        RECT 281.400 268.050 282.600 272.400 ;
        RECT 286.950 271.950 289.050 274.050 ;
        RECT 280.950 265.950 283.050 268.050 ;
        RECT 283.950 267.600 286.050 271.050 ;
        RECT 296.400 267.600 297.600 286.950 ;
        RECT 307.950 271.950 310.050 274.050 ;
        RECT 283.950 267.000 297.600 267.600 ;
        RECT 284.400 266.400 297.600 267.000 ;
        RECT 271.950 259.950 274.050 262.050 ;
        RECT 280.950 261.600 283.050 262.050 ;
        RECT 285.000 261.600 289.050 262.050 ;
        RECT 275.400 260.400 283.050 261.600 ;
        RECT 272.400 235.050 273.600 259.950 ;
        RECT 275.400 244.050 276.600 260.400 ;
        RECT 280.950 259.950 283.050 260.400 ;
        RECT 284.400 259.950 289.050 261.600 ;
        RECT 277.950 250.950 280.050 253.050 ;
        RECT 274.950 241.950 277.050 244.050 ;
        RECT 278.400 241.050 279.600 250.950 ;
        RECT 284.400 247.050 285.600 259.950 ;
        RECT 304.950 253.950 307.050 256.050 ;
        RECT 283.950 244.950 286.050 247.050 ;
        RECT 305.400 241.050 306.600 253.950 ;
        RECT 277.950 238.950 280.050 241.050 ;
        RECT 292.950 238.950 295.050 241.050 ;
        RECT 304.950 238.950 307.050 241.050 ;
        RECT 286.950 235.950 289.050 238.050 ;
        RECT 271.950 232.950 274.050 235.050 ;
        RECT 265.950 226.950 268.050 229.050 ;
        RECT 280.950 226.950 283.050 229.050 ;
        RECT 262.950 220.950 265.050 223.050 ;
        RECT 265.950 217.950 268.050 220.050 ;
        RECT 271.950 217.950 274.050 220.050 ;
        RECT 250.950 208.950 253.050 211.050 ;
        RECT 260.400 208.950 265.050 211.050 ;
        RECT 241.950 202.950 244.050 205.050 ;
        RECT 260.400 202.050 261.600 208.950 ;
        RECT 226.950 199.950 229.050 202.050 ;
        RECT 259.950 199.950 262.050 202.050 ;
        RECT 266.400 196.050 267.600 217.950 ;
        RECT 223.950 193.950 226.050 196.050 ;
        RECT 265.950 193.950 268.050 196.050 ;
        RECT 272.400 190.050 273.600 217.950 ;
        RECT 253.950 187.950 256.050 190.050 ;
        RECT 271.950 187.950 274.050 190.050 ;
        RECT 238.950 181.950 241.050 184.050 ;
        RECT 226.950 157.950 229.050 160.050 ;
        RECT 220.950 139.950 223.050 142.050 ;
        RECT 221.400 118.050 222.600 139.950 ;
        RECT 227.400 139.050 228.600 157.950 ;
        RECT 239.400 157.050 240.600 181.950 ;
        RECT 254.400 175.050 255.600 187.950 ;
        RECT 281.400 184.050 282.600 226.950 ;
        RECT 283.950 220.950 286.050 223.050 ;
        RECT 284.400 211.050 285.600 220.950 ;
        RECT 283.950 208.950 286.050 211.050 ;
        RECT 287.400 202.050 288.600 235.950 ;
        RECT 293.400 222.600 294.600 238.950 ;
        RECT 308.400 238.050 309.600 271.950 ;
        RECT 311.400 252.600 312.600 286.950 ;
        RECT 314.400 286.050 315.600 296.400 ;
        RECT 316.950 292.950 319.050 295.050 ;
        RECT 313.950 283.950 316.050 286.050 ;
        RECT 317.400 280.050 318.600 292.950 ;
        RECT 316.950 277.950 319.050 280.050 ;
        RECT 317.400 261.600 318.600 277.950 ;
        RECT 320.400 274.050 321.600 316.950 ;
        RECT 319.950 271.950 322.050 274.050 ;
        RECT 326.400 273.600 327.600 361.950 ;
        RECT 332.400 360.600 333.600 394.950 ;
        RECT 329.400 359.400 333.600 360.600 ;
        RECT 329.400 346.050 330.600 359.400 ;
        RECT 335.400 355.050 336.600 397.950 ;
        RECT 352.950 379.950 355.050 382.050 ;
        RECT 353.400 376.050 354.600 379.950 ;
        RECT 346.950 373.950 349.050 376.050 ;
        RECT 352.950 373.950 355.050 376.050 ;
        RECT 347.400 361.050 348.600 373.950 ;
        RECT 365.400 364.050 366.600 406.950 ;
        RECT 371.400 403.050 372.600 415.950 ;
        RECT 377.400 409.050 378.600 421.950 ;
        RECT 376.950 406.950 379.050 409.050 ;
        RECT 382.950 406.950 385.050 409.050 ;
        RECT 370.950 400.950 373.050 403.050 ;
        RECT 383.400 394.050 384.600 406.950 ;
        RECT 382.950 391.950 385.050 394.050 ;
        RECT 398.400 391.050 399.600 424.950 ;
        RECT 401.400 421.050 402.600 442.950 ;
        RECT 406.950 424.950 409.050 427.050 ;
        RECT 407.400 421.050 408.600 424.950 ;
        RECT 400.950 418.950 403.050 421.050 ;
        RECT 406.950 418.950 409.050 421.050 ;
        RECT 403.950 391.950 406.050 394.050 ;
        RECT 397.950 388.950 400.050 391.050 ;
        RECT 398.400 376.050 399.600 388.950 ;
        RECT 391.950 375.600 394.050 376.050 ;
        RECT 386.400 375.000 394.050 375.600 ;
        RECT 385.950 374.400 394.050 375.000 ;
        RECT 385.950 370.950 388.050 374.400 ;
        RECT 391.950 373.950 394.050 374.400 ;
        RECT 397.950 373.950 400.050 376.050 ;
        RECT 404.400 367.050 405.600 391.950 ;
        RECT 379.950 364.950 382.050 367.050 ;
        RECT 394.950 364.950 397.050 367.050 ;
        RECT 403.950 364.950 406.050 367.050 ;
        RECT 349.950 361.950 352.050 364.050 ;
        RECT 364.950 363.600 367.050 364.050 ;
        RECT 362.400 362.400 367.050 363.600 ;
        RECT 346.950 358.950 349.050 361.050 ;
        RECT 334.950 352.950 337.050 355.050 ;
        RECT 328.950 343.950 331.050 346.050 ;
        RECT 340.950 340.950 343.050 343.050 ;
        RECT 341.400 325.050 342.600 340.950 ;
        RECT 340.950 322.950 343.050 325.050 ;
        RECT 341.400 310.050 342.600 322.950 ;
        RECT 340.950 307.950 343.050 310.050 ;
        RECT 350.400 307.050 351.600 361.950 ;
        RECT 355.950 352.950 358.050 355.050 ;
        RECT 356.400 343.050 357.600 352.950 ;
        RECT 355.950 340.950 358.050 343.050 ;
        RECT 362.400 340.050 363.600 362.400 ;
        RECT 364.950 361.950 367.050 362.400 ;
        RECT 373.950 361.950 376.050 364.050 ;
        RECT 374.400 355.050 375.600 361.950 ;
        RECT 373.950 352.950 376.050 355.050 ;
        RECT 361.950 337.950 364.050 340.050 ;
        RECT 380.400 334.050 381.600 364.950 ;
        RECT 388.950 349.950 391.050 352.050 ;
        RECT 389.400 334.050 390.600 349.950 ;
        RECT 355.950 331.950 358.050 334.050 ;
        RECT 379.950 331.950 382.050 334.050 ;
        RECT 388.950 331.950 391.050 334.050 ;
        RECT 349.950 304.950 352.050 307.050 ;
        RECT 356.400 304.050 357.600 331.950 ;
        RECT 395.400 313.050 396.600 364.950 ;
        RECT 404.400 343.050 405.600 364.950 ;
        RECT 403.950 340.950 406.050 343.050 ;
        RECT 394.950 310.950 397.050 313.050 ;
        RECT 395.400 309.600 396.600 310.950 ;
        RECT 395.400 308.400 399.600 309.600 ;
        RECT 373.950 304.950 376.050 307.050 ;
        RECT 355.950 301.950 358.050 304.050 ;
        RECT 367.950 301.950 370.050 304.050 ;
        RECT 368.400 298.050 369.600 301.950 ;
        RECT 360.000 297.600 364.050 298.050 ;
        RECT 359.400 295.950 364.050 297.600 ;
        RECT 367.950 295.950 370.050 298.050 ;
        RECT 359.400 286.050 360.600 295.950 ;
        RECT 364.950 286.950 367.050 289.050 ;
        RECT 352.950 283.950 355.050 286.050 ;
        RECT 358.950 283.950 361.050 286.050 ;
        RECT 340.950 274.950 343.050 277.050 ;
        RECT 326.400 272.400 330.600 273.600 ;
        RECT 314.400 260.400 318.600 261.600 ;
        RECT 314.400 256.050 315.600 260.400 ;
        RECT 319.950 259.950 322.050 262.050 ;
        RECT 313.950 253.950 316.050 256.050 ;
        RECT 311.400 251.400 315.600 252.600 ;
        RECT 307.950 235.950 310.050 238.050 ;
        RECT 314.400 232.050 315.600 251.400 ;
        RECT 320.400 241.050 321.600 259.950 ;
        RECT 319.950 238.950 322.050 241.050 ;
        RECT 325.950 238.950 328.050 241.050 ;
        RECT 313.950 229.950 316.050 232.050 ;
        RECT 326.400 229.050 327.600 238.950 ;
        RECT 298.950 225.600 301.050 229.050 ;
        RECT 325.950 226.950 328.050 229.050 ;
        RECT 290.400 221.400 294.600 222.600 ;
        RECT 296.400 225.000 301.050 225.600 ;
        RECT 296.400 224.400 300.600 225.000 ;
        RECT 290.400 208.050 291.600 221.400 ;
        RECT 296.400 217.050 297.600 224.400 ;
        RECT 316.950 223.950 319.050 226.050 ;
        RECT 304.950 219.600 307.050 223.050 ;
        RECT 317.400 220.050 318.600 223.950 ;
        RECT 310.950 219.600 313.050 220.050 ;
        RECT 304.950 219.000 313.050 219.600 ;
        RECT 305.400 218.400 313.050 219.000 ;
        RECT 310.950 217.950 313.050 218.400 ;
        RECT 316.950 217.950 319.050 220.050 ;
        RECT 292.950 215.400 297.600 217.050 ;
        RECT 292.950 214.950 297.000 215.400 ;
        RECT 326.400 211.050 327.600 226.950 ;
        RECT 307.950 208.950 310.050 211.050 ;
        RECT 319.950 208.950 322.050 211.050 ;
        RECT 325.950 208.950 328.050 211.050 ;
        RECT 289.950 205.950 292.050 208.050 ;
        RECT 294.000 207.600 298.050 208.050 ;
        RECT 293.400 205.950 298.050 207.600 ;
        RECT 293.400 202.050 294.600 205.950 ;
        RECT 286.950 199.950 289.050 202.050 ;
        RECT 292.950 199.950 295.050 202.050 ;
        RECT 283.950 187.950 286.050 190.050 ;
        RECT 284.400 184.050 285.600 187.950 ;
        RECT 280.950 181.950 283.050 184.050 ;
        RECT 284.400 182.400 289.050 184.050 ;
        RECT 285.000 181.950 289.050 182.400 ;
        RECT 265.950 175.950 268.050 178.050 ;
        RECT 253.950 172.950 256.050 175.050 ;
        RECT 259.950 172.950 262.050 175.050 ;
        RECT 260.400 169.050 261.600 172.950 ;
        RECT 266.400 169.050 267.600 175.950 ;
        RECT 259.950 166.950 262.050 169.050 ;
        RECT 265.950 166.950 268.050 169.050 ;
        RECT 274.950 157.950 277.050 160.050 ;
        RECT 238.950 154.950 241.050 157.050 ;
        RECT 265.950 154.950 268.050 157.050 ;
        RECT 266.400 139.050 267.600 154.950 ;
        RECT 275.400 139.050 276.600 157.950 ;
        RECT 293.400 154.050 294.600 199.950 ;
        RECT 308.400 178.050 309.600 208.950 ;
        RECT 320.400 205.050 321.600 208.950 ;
        RECT 319.950 202.950 322.050 205.050 ;
        RECT 326.400 193.050 327.600 208.950 ;
        RECT 325.950 190.950 328.050 193.050 ;
        RECT 319.950 187.950 322.050 190.050 ;
        RECT 304.950 176.400 309.600 178.050 ;
        RECT 304.950 175.950 309.000 176.400 ;
        RECT 313.950 174.600 316.050 178.050 ;
        RECT 313.950 174.000 318.600 174.600 ;
        RECT 314.400 173.400 318.600 174.000 ;
        RECT 317.400 169.050 318.600 173.400 ;
        RECT 316.950 166.950 319.050 169.050 ;
        RECT 310.950 160.950 313.050 163.050 ;
        RECT 301.950 154.950 304.050 157.050 ;
        RECT 286.950 151.950 289.050 154.050 ;
        RECT 292.950 151.950 295.050 154.050 ;
        RECT 227.400 136.950 232.050 139.050 ;
        RECT 238.950 138.600 241.050 139.050 ;
        RECT 233.400 137.400 241.050 138.600 ;
        RECT 220.950 115.950 223.050 118.050 ;
        RECT 208.950 112.950 211.050 115.050 ;
        RECT 217.950 112.950 220.050 115.050 ;
        RECT 227.400 114.600 228.600 136.950 ;
        RECT 233.400 135.600 234.600 137.400 ;
        RECT 238.950 136.950 241.050 137.400 ;
        RECT 265.950 136.950 268.050 139.050 ;
        RECT 274.950 136.950 277.050 139.050 ;
        RECT 230.400 134.400 234.600 135.600 ;
        RECT 230.400 130.050 231.600 134.400 ;
        RECT 256.950 130.950 259.050 133.050 ;
        RECT 229.950 127.950 232.050 130.050 ;
        RECT 229.950 115.950 232.050 118.050 ;
        RECT 244.950 115.950 247.050 118.050 ;
        RECT 224.400 113.400 228.600 114.600 ;
        RECT 209.400 109.050 210.600 112.950 ;
        RECT 208.950 106.950 211.050 109.050 ;
        RECT 202.950 88.950 205.050 91.050 ;
        RECT 224.400 82.050 225.600 113.400 ;
        RECT 226.950 109.950 229.050 112.050 ;
        RECT 227.400 97.050 228.600 109.950 ;
        RECT 230.400 109.050 231.600 115.950 ;
        RECT 245.400 112.050 246.600 115.950 ;
        RECT 257.400 115.050 258.600 130.950 ;
        RECT 287.400 118.050 288.600 151.950 ;
        RECT 302.400 139.050 303.600 154.950 ;
        RECT 304.950 151.950 307.050 154.050 ;
        RECT 301.950 136.950 304.050 139.050 ;
        RECT 292.950 130.950 295.050 133.050 ;
        RECT 293.400 121.050 294.600 130.950 ;
        RECT 292.950 118.950 295.050 121.050 ;
        RECT 301.950 118.950 304.050 121.050 ;
        RECT 274.950 115.950 277.050 118.050 ;
        RECT 286.950 115.950 289.050 118.050 ;
        RECT 256.950 112.950 259.050 115.050 ;
        RECT 244.950 109.950 247.050 112.050 ;
        RECT 229.950 106.950 232.050 109.050 ;
        RECT 245.400 106.050 246.600 109.950 ;
        RECT 244.950 103.950 247.050 106.050 ;
        RECT 256.950 103.950 259.050 106.050 ;
        RECT 257.400 97.050 258.600 103.950 ;
        RECT 275.400 97.050 276.600 115.950 ;
        RECT 302.400 115.050 303.600 118.950 ;
        RECT 295.950 112.950 298.050 115.050 ;
        RECT 301.950 112.950 304.050 115.050 ;
        RECT 286.950 109.950 289.050 112.050 ;
        RECT 226.950 94.950 229.050 97.050 ;
        RECT 247.950 94.950 250.050 97.050 ;
        RECT 253.950 95.400 258.600 97.050 ;
        RECT 253.950 94.950 258.000 95.400 ;
        RECT 274.950 94.950 277.050 97.050 ;
        RECT 248.400 91.050 249.600 94.950 ;
        RECT 268.950 91.950 271.050 94.050 ;
        RECT 247.950 88.950 250.050 91.050 ;
        RECT 187.950 79.950 190.050 82.050 ;
        RECT 223.950 79.950 226.050 82.050 ;
        RECT 235.950 79.950 238.050 82.050 ;
        RECT 220.950 73.950 223.050 76.050 ;
        RECT 184.950 70.950 187.050 73.050 ;
        RECT 163.950 67.950 166.050 70.050 ;
        RECT 172.950 67.950 175.050 70.050 ;
        RECT 160.950 61.950 163.050 64.050 ;
        RECT 164.400 55.050 165.600 67.950 ;
        RECT 185.400 64.050 186.600 70.950 ;
        RECT 208.950 67.950 211.050 70.050 ;
        RECT 209.400 64.050 210.600 67.950 ;
        RECT 184.950 61.950 187.050 64.050 ;
        RECT 178.950 60.600 181.050 61.050 ;
        RECT 190.950 60.600 193.050 64.050 ;
        RECT 208.950 61.950 211.050 64.050 ;
        RECT 214.950 63.600 219.000 64.050 ;
        RECT 214.950 61.950 219.600 63.600 ;
        RECT 178.950 60.000 193.050 60.600 ;
        RECT 178.950 59.400 192.600 60.000 ;
        RECT 178.950 58.950 181.050 59.400 ;
        RECT 163.950 52.950 166.050 55.050 ;
        RECT 193.950 52.950 196.050 55.050 ;
        RECT 205.950 52.950 208.050 55.050 ;
        RECT 100.950 43.950 103.050 46.050 ;
        RECT 154.950 43.950 157.050 46.050 ;
        RECT 101.400 37.050 102.600 43.950 ;
        RECT 151.950 40.950 154.050 43.050 ;
        RECT 100.950 34.950 103.050 37.050 ;
        RECT 118.950 34.950 121.050 37.050 ;
        RECT 101.400 28.050 102.600 34.950 ;
        RECT 119.400 28.050 120.600 34.950 ;
        RECT 136.950 31.950 139.050 34.050 ;
        RECT 137.400 28.050 138.600 31.950 ;
        RECT 152.400 28.050 153.600 40.950 ;
        RECT 100.950 25.950 103.050 28.050 ;
        RECT 118.950 25.950 121.050 28.050 ;
        RECT 136.950 25.950 139.050 28.050 ;
        RECT 151.950 25.950 154.050 28.050 ;
        RECT 155.400 22.050 156.600 43.950 ;
        RECT 163.950 40.950 166.050 43.050 ;
        RECT 181.950 40.950 184.050 43.050 ;
        RECT 164.400 22.050 165.600 40.950 ;
        RECT 182.400 28.050 183.600 40.950 ;
        RECT 181.950 24.600 184.050 28.050 ;
        RECT 187.950 25.950 190.050 28.050 ;
        RECT 181.950 24.000 186.600 24.600 ;
        RECT 182.400 23.400 186.600 24.000 ;
        RECT 112.950 21.600 115.050 22.050 ;
        RECT 107.400 21.000 115.050 21.600 ;
        RECT 106.950 20.400 115.050 21.000 ;
        RECT 91.950 16.950 94.050 19.050 ;
        RECT 97.950 16.950 100.050 19.050 ;
        RECT 106.950 16.950 109.050 20.400 ;
        RECT 112.950 19.950 115.050 20.400 ;
        RECT 133.950 19.950 136.050 22.050 ;
        RECT 154.950 19.950 157.050 22.050 ;
        RECT 163.950 19.950 166.050 22.050 ;
        RECT 134.400 13.050 135.600 19.950 ;
        RECT 185.400 19.050 186.600 23.400 ;
        RECT 139.950 16.950 142.050 19.050 ;
        RECT 145.950 16.950 148.050 19.050 ;
        RECT 184.950 16.950 187.050 19.050 ;
        RECT 140.400 13.050 141.600 16.950 ;
        RECT 133.950 10.950 136.050 13.050 ;
        RECT 139.950 10.950 142.050 13.050 ;
        RECT 146.400 7.050 147.600 16.950 ;
        RECT 188.400 7.050 189.600 25.950 ;
        RECT 194.400 13.050 195.600 52.950 ;
        RECT 206.400 40.050 207.600 52.950 ;
        RECT 218.400 52.050 219.600 61.950 ;
        RECT 221.400 55.050 222.600 73.950 ;
        RECT 224.400 61.050 225.600 79.950 ;
        RECT 232.950 73.950 235.050 76.050 ;
        RECT 233.400 61.050 234.600 73.950 ;
        RECT 223.950 58.950 226.050 61.050 ;
        RECT 232.950 58.950 235.050 61.050 ;
        RECT 220.950 52.950 223.050 55.050 ;
        RECT 217.950 49.950 220.050 52.050 ;
        RECT 223.950 51.600 226.050 52.050 ;
        RECT 232.950 51.600 235.050 52.050 ;
        RECT 223.950 50.400 235.050 51.600 ;
        RECT 223.950 49.950 226.050 50.400 ;
        RECT 232.950 49.950 235.050 50.400 ;
        RECT 232.950 45.600 235.050 46.050 ;
        RECT 227.400 44.400 235.050 45.600 ;
        RECT 205.950 37.950 208.050 40.050 ;
        RECT 217.950 37.950 220.050 40.050 ;
        RECT 206.400 19.050 207.600 37.950 ;
        RECT 218.400 28.050 219.600 37.950 ;
        RECT 227.400 28.050 228.600 44.400 ;
        RECT 232.950 43.950 235.050 44.400 ;
        RECT 229.950 34.950 232.050 37.050 ;
        RECT 217.950 25.950 220.050 28.050 ;
        RECT 226.950 25.950 229.050 28.050 ;
        RECT 202.950 17.400 207.600 19.050 ;
        RECT 202.950 16.950 207.000 17.400 ;
        RECT 220.950 16.950 223.050 19.050 ;
        RECT 226.950 16.950 229.050 19.050 ;
        RECT 221.400 13.050 222.600 16.950 ;
        RECT 193.950 10.950 196.050 13.050 ;
        RECT 220.950 10.950 223.050 13.050 ;
        RECT 227.400 7.050 228.600 16.950 ;
        RECT 230.400 15.600 231.600 34.950 ;
        RECT 236.400 22.050 237.600 79.950 ;
        RECT 269.400 76.050 270.600 91.950 ;
        RECT 275.400 91.050 276.600 94.950 ;
        RECT 274.950 88.950 277.050 91.050 ;
        RECT 280.950 79.950 283.050 82.050 ;
        RECT 268.950 73.950 271.050 76.050 ;
        RECT 271.950 61.950 274.050 64.050 ;
        RECT 248.400 57.000 258.600 57.600 ;
        RECT 248.400 56.400 259.050 57.000 ;
        RECT 241.950 51.600 244.050 52.050 ;
        RECT 248.400 51.600 249.600 56.400 ;
        RECT 250.950 54.600 255.000 55.050 ;
        RECT 250.950 52.950 255.600 54.600 ;
        RECT 256.950 52.950 259.050 56.400 ;
        RECT 241.950 50.400 249.600 51.600 ;
        RECT 241.950 49.950 244.050 50.400 ;
        RECT 254.400 49.050 255.600 52.950 ;
        RECT 253.950 46.950 256.050 49.050 ;
        RECT 241.950 43.950 244.050 46.050 ;
        RECT 242.400 22.050 243.600 43.950 ;
        RECT 272.400 40.050 273.600 61.950 ;
        RECT 281.400 61.050 282.600 79.950 ;
        RECT 287.400 61.050 288.600 109.950 ;
        RECT 296.400 109.050 297.600 112.950 ;
        RECT 302.400 109.050 303.600 112.950 ;
        RECT 295.950 106.950 298.050 109.050 ;
        RECT 301.950 106.950 304.050 109.050 ;
        RECT 305.400 100.050 306.600 151.950 ;
        RECT 311.400 123.600 312.600 160.950 ;
        RECT 317.400 157.050 318.600 166.950 ;
        RECT 320.400 160.200 321.600 187.950 ;
        RECT 329.400 186.600 330.600 272.400 ;
        RECT 341.400 262.050 342.600 274.950 ;
        RECT 353.400 262.050 354.600 283.950 ;
        RECT 355.950 279.600 358.050 283.050 ;
        RECT 355.950 279.000 360.600 279.600 ;
        RECT 356.400 278.400 360.600 279.000 ;
        RECT 340.950 259.950 343.050 262.050 ;
        RECT 352.950 259.950 355.050 262.050 ;
        RECT 331.950 250.950 334.050 253.050 ;
        RECT 337.950 252.600 340.050 253.050 ;
        RECT 337.950 251.400 345.600 252.600 ;
        RECT 337.950 250.950 340.050 251.400 ;
        RECT 332.400 235.050 333.600 250.950 ;
        RECT 344.400 244.050 345.600 251.400 ;
        RECT 355.950 247.950 358.050 250.050 ;
        RECT 337.950 241.950 340.050 244.050 ;
        RECT 343.950 241.950 346.050 244.050 ;
        RECT 331.950 232.950 334.050 235.050 ;
        RECT 338.400 226.050 339.600 241.950 ;
        RECT 337.950 223.950 340.050 226.050 ;
        RECT 346.950 223.950 349.050 226.050 ;
        RECT 352.950 223.950 355.050 226.050 ;
        RECT 347.400 220.050 348.600 223.950 ;
        RECT 346.950 217.950 349.050 220.050 ;
        RECT 349.950 205.950 352.050 208.050 ;
        RECT 331.950 202.950 334.050 205.050 ;
        RECT 332.400 193.050 333.600 202.950 ;
        RECT 331.950 190.950 334.050 193.050 ;
        RECT 329.400 185.400 333.600 186.600 ;
        RECT 328.950 181.950 331.050 184.050 ;
        RECT 319.800 158.100 321.900 160.200 ;
        RECT 329.400 160.050 330.600 181.950 ;
        RECT 332.400 175.050 333.600 185.400 ;
        RECT 343.950 181.950 346.050 184.050 ;
        RECT 331.950 172.950 334.050 175.050 ;
        RECT 337.950 174.600 340.050 175.050 ;
        RECT 344.400 174.600 345.600 181.950 ;
        RECT 350.400 174.600 351.600 205.950 ;
        RECT 353.400 190.050 354.600 223.950 ;
        RECT 356.400 196.050 357.600 247.950 ;
        RECT 359.400 247.050 360.600 278.400 ;
        RECT 365.400 277.050 366.600 286.950 ;
        RECT 370.950 283.950 373.050 286.050 ;
        RECT 364.950 274.950 367.050 277.050 ;
        RECT 371.400 274.050 372.600 283.950 ;
        RECT 370.950 271.950 373.050 274.050 ;
        RECT 358.950 244.950 361.050 247.050 ;
        RECT 361.950 229.950 364.050 232.050 ;
        RECT 358.950 217.950 361.050 220.050 ;
        RECT 359.400 211.050 360.600 217.950 ;
        RECT 362.400 211.050 363.600 229.950 ;
        RECT 358.950 208.950 361.050 211.050 ;
        RECT 361.950 208.950 364.050 211.050 ;
        RECT 355.950 193.950 358.050 196.050 ;
        RECT 374.400 195.600 375.600 304.950 ;
        RECT 378.000 294.600 382.050 295.050 ;
        RECT 377.400 292.950 382.050 294.600 ;
        RECT 388.950 292.950 391.050 295.050 ;
        RECT 377.400 280.050 378.600 292.950 ;
        RECT 389.400 282.600 390.600 292.950 ;
        RECT 386.400 281.400 390.600 282.600 ;
        RECT 376.950 277.950 379.050 280.050 ;
        RECT 386.400 274.050 387.600 281.400 ;
        RECT 391.950 274.950 394.050 277.050 ;
        RECT 385.950 271.950 388.050 274.050 ;
        RECT 382.950 268.950 385.050 271.050 ;
        RECT 383.400 265.050 384.600 268.950 ;
        RECT 388.950 265.950 391.050 268.050 ;
        RECT 382.950 262.950 385.050 265.050 ;
        RECT 389.400 262.050 390.600 265.950 ;
        RECT 376.950 259.950 379.050 262.050 ;
        RECT 388.950 259.950 391.050 262.050 ;
        RECT 377.400 253.050 378.600 259.950 ;
        RECT 377.400 251.400 382.050 253.050 ;
        RECT 378.000 250.950 382.050 251.400 ;
        RECT 385.950 250.950 388.050 253.050 ;
        RECT 386.400 244.050 387.600 250.950 ;
        RECT 392.400 247.050 393.600 274.950 ;
        RECT 394.950 267.600 397.050 268.050 ;
        RECT 398.400 267.600 399.600 308.400 ;
        RECT 406.950 307.950 409.050 310.050 ;
        RECT 407.400 289.050 408.600 307.950 ;
        RECT 406.950 286.950 409.050 289.050 ;
        RECT 394.950 266.400 399.600 267.600 ;
        RECT 394.950 265.950 397.050 266.400 ;
        RECT 395.400 253.050 396.600 265.950 ;
        RECT 394.950 250.950 397.050 253.050 ;
        RECT 391.950 244.950 394.050 247.050 ;
        RECT 410.400 244.050 411.600 472.950 ;
        RECT 421.950 469.950 424.050 472.050 ;
        RECT 418.950 460.950 421.050 463.050 ;
        RECT 412.950 457.950 415.050 460.050 ;
        RECT 413.400 397.050 414.600 457.950 ;
        RECT 419.400 454.050 420.600 460.950 ;
        RECT 418.950 451.950 421.050 454.050 ;
        RECT 422.400 445.050 423.600 469.950 ;
        RECT 436.950 463.950 439.050 466.050 ;
        RECT 437.400 454.050 438.600 463.950 ;
        RECT 440.400 460.050 441.600 493.950 ;
        RECT 464.400 488.400 477.600 489.600 ;
        RECT 464.400 483.600 465.600 488.400 ;
        RECT 466.950 484.950 469.050 487.050 ;
        RECT 472.950 484.950 475.050 487.050 ;
        RECT 461.400 482.400 465.600 483.600 ;
        RECT 454.950 480.600 457.050 481.050 ;
        RECT 461.400 480.600 462.600 482.400 ;
        RECT 467.400 481.050 468.600 484.950 ;
        RECT 454.950 479.400 462.600 480.600 ;
        RECT 454.950 478.950 457.050 479.400 ;
        RECT 466.950 478.950 469.050 481.050 ;
        RECT 473.400 478.050 474.600 484.950 ;
        RECT 476.400 478.050 477.600 488.400 ;
        RECT 472.800 475.950 474.900 478.050 ;
        RECT 476.100 475.950 478.200 478.050 ;
        RECT 463.950 469.950 466.050 472.050 ;
        RECT 442.950 466.950 445.050 469.050 ;
        RECT 439.950 457.950 442.050 460.050 ;
        RECT 443.400 454.050 444.600 466.950 ;
        RECT 457.950 460.950 460.050 463.050 ;
        RECT 424.950 453.600 429.000 454.050 ;
        RECT 424.950 451.950 429.600 453.600 ;
        RECT 436.950 451.950 439.050 454.050 ;
        RECT 442.950 451.950 445.050 454.050 ;
        RECT 421.950 442.950 424.050 445.050 ;
        RECT 415.950 439.950 418.050 442.050 ;
        RECT 416.400 418.050 417.600 439.950 ;
        RECT 428.400 439.050 429.600 451.950 ;
        RECT 458.400 445.050 459.600 460.950 ;
        RECT 464.400 454.050 465.600 469.950 ;
        RECT 469.950 463.950 472.050 466.050 ;
        RECT 481.950 463.950 484.050 466.050 ;
        RECT 470.400 460.050 471.600 463.950 ;
        RECT 469.950 457.950 472.050 460.050 ;
        RECT 470.400 454.050 471.600 457.950 ;
        RECT 482.400 454.050 483.600 463.950 ;
        RECT 485.400 454.050 486.600 493.950 ;
        RECT 497.400 487.050 498.600 514.950 ;
        RECT 503.400 511.050 504.600 550.950 ;
        RECT 518.400 547.050 519.600 562.950 ;
        RECT 521.400 559.050 522.600 619.950 ;
        RECT 530.400 583.050 531.600 625.950 ;
        RECT 545.400 622.050 546.600 670.950 ;
        RECT 551.400 670.050 552.600 685.950 ;
        RECT 559.950 676.950 562.050 679.050 ;
        RECT 577.950 678.600 580.050 679.050 ;
        RECT 583.950 678.600 586.050 679.050 ;
        RECT 577.950 677.400 586.050 678.600 ;
        RECT 577.950 676.950 580.050 677.400 ;
        RECT 583.950 676.950 586.050 677.400 ;
        RECT 560.400 670.050 561.600 676.950 ;
        RECT 565.950 673.950 568.050 676.050 ;
        RECT 589.950 673.950 592.050 676.050 ;
        RECT 550.950 667.950 553.050 670.050 ;
        RECT 559.950 667.950 562.050 670.050 ;
        RECT 553.950 664.950 556.050 667.050 ;
        RECT 554.400 661.050 555.600 664.950 ;
        RECT 553.950 658.950 556.050 661.050 ;
        RECT 566.400 655.050 567.600 673.950 ;
        RECT 568.950 670.950 571.050 673.050 ;
        RECT 559.950 652.950 562.050 655.050 ;
        RECT 565.950 652.950 568.050 655.050 ;
        RECT 550.950 649.950 553.050 652.050 ;
        RECT 551.400 628.050 552.600 649.950 ;
        RECT 550.950 625.950 553.050 628.050 ;
        RECT 532.950 619.950 535.050 622.050 ;
        RECT 544.950 619.950 547.050 622.050 ;
        RECT 533.400 601.050 534.600 619.950 ;
        RECT 560.400 616.050 561.600 652.950 ;
        RECT 569.400 646.050 570.600 670.950 ;
        RECT 577.800 658.950 579.900 661.050 ;
        RECT 565.950 644.400 570.600 646.050 ;
        RECT 565.950 643.950 570.000 644.400 ;
        RECT 562.950 634.950 565.050 637.050 ;
        RECT 563.400 619.050 564.600 634.950 ;
        RECT 568.950 628.950 571.050 631.050 ;
        RECT 569.400 625.050 570.600 628.950 ;
        RECT 578.400 628.050 579.600 658.950 ;
        RECT 590.400 658.050 591.600 673.950 ;
        RECT 593.400 661.050 594.600 706.950 ;
        RECT 596.400 670.050 597.600 706.950 ;
        RECT 601.950 694.950 604.050 697.050 ;
        RECT 602.400 673.050 603.600 694.950 ;
        RECT 608.400 681.600 609.600 712.950 ;
        RECT 614.400 694.050 615.600 712.950 ;
        RECT 620.400 709.050 621.600 718.950 ;
        RECT 625.950 709.950 628.050 712.050 ;
        RECT 619.800 706.950 621.900 709.050 ;
        RECT 623.100 706.950 625.200 709.050 ;
        RECT 623.400 700.050 624.600 706.950 ;
        RECT 622.950 697.950 625.050 700.050 ;
        RECT 626.400 697.050 627.600 709.950 ;
        RECT 632.400 709.050 633.600 749.400 ;
        RECT 641.400 748.050 642.600 754.950 ;
        RECT 644.400 751.050 645.600 754.950 ;
        RECT 643.800 748.950 645.900 751.050 ;
        RECT 647.100 748.950 649.200 751.050 ;
        RECT 640.950 745.950 643.050 748.050 ;
        RECT 634.950 736.950 637.050 739.050 ;
        RECT 631.950 706.950 634.050 709.050 ;
        RECT 625.950 694.950 628.050 697.050 ;
        RECT 614.100 691.950 616.200 694.050 ;
        RECT 622.950 685.950 625.050 688.050 ;
        RECT 605.400 680.400 609.600 681.600 ;
        RECT 601.950 670.950 604.050 673.050 ;
        RECT 605.400 670.050 606.600 680.400 ;
        RECT 607.950 676.950 610.050 679.050 ;
        RECT 608.400 673.050 609.600 676.950 ;
        RECT 607.950 670.950 610.050 673.050 ;
        RECT 613.950 670.950 616.050 673.050 ;
        RECT 595.800 667.950 597.900 670.050 ;
        RECT 604.950 667.950 607.050 670.050 ;
        RECT 592.950 658.950 595.050 661.050 ;
        RECT 604.950 658.950 607.050 661.050 ;
        RECT 589.950 655.950 592.050 658.050 ;
        RECT 598.950 655.950 601.050 658.050 ;
        RECT 586.950 642.600 589.050 646.050 ;
        RECT 599.400 643.050 600.600 655.950 ;
        RECT 592.950 642.600 595.050 643.050 ;
        RECT 586.950 642.000 595.050 642.600 ;
        RECT 587.400 641.400 595.050 642.000 ;
        RECT 592.950 640.950 595.050 641.400 ;
        RECT 598.950 640.950 601.050 643.050 ;
        RECT 577.950 625.950 580.050 628.050 ;
        RECT 568.950 622.950 571.050 625.050 ;
        RECT 593.400 619.050 594.600 640.950 ;
        RECT 562.950 616.950 565.050 619.050 ;
        RECT 577.950 616.950 580.050 619.050 ;
        RECT 592.950 616.950 595.050 619.050 ;
        RECT 559.950 613.950 562.050 616.050 ;
        RECT 563.400 610.050 564.600 616.950 ;
        RECT 578.400 610.050 579.600 616.950 ;
        RECT 605.400 610.050 606.600 658.950 ;
        RECT 614.400 658.050 615.600 670.950 ;
        RECT 623.400 670.050 624.600 685.950 ;
        RECT 625.950 673.950 628.050 676.050 ;
        RECT 622.950 667.950 625.050 670.050 ;
        RECT 626.400 661.050 627.600 673.950 ;
        RECT 635.400 673.050 636.600 736.950 ;
        RECT 644.400 721.050 645.600 748.950 ;
        RECT 647.400 739.050 648.600 748.950 ;
        RECT 650.400 745.050 651.600 787.950 ;
        RECT 652.950 763.950 655.050 766.050 ;
        RECT 653.400 745.050 654.600 763.950 ;
        RECT 659.400 759.600 660.600 823.950 ;
        RECT 662.400 820.050 663.600 847.950 ;
        RECT 680.400 844.050 681.600 865.950 ;
        RECT 686.400 856.050 687.600 874.950 ;
        RECT 689.400 868.050 690.600 883.950 ;
        RECT 688.950 865.950 691.050 868.050 ;
        RECT 692.400 864.600 693.600 898.950 ;
        RECT 719.400 896.400 729.600 897.600 ;
        RECT 719.400 892.050 720.600 896.400 ;
        RECT 724.950 892.950 727.050 895.050 ;
        RECT 728.400 894.600 729.600 896.400 ;
        RECT 736.950 895.950 739.050 898.050 ;
        RECT 728.400 893.400 732.600 894.600 ;
        RECT 718.950 889.950 721.050 892.050 ;
        RECT 725.400 886.050 726.600 892.950 ;
        RECT 724.950 885.600 727.050 886.050 ;
        RECT 716.400 884.400 727.050 885.600 ;
        RECT 716.400 880.050 717.600 884.400 ;
        RECT 724.950 883.950 727.050 884.400 ;
        RECT 731.400 880.050 732.600 893.400 ;
        RECT 715.800 877.950 717.900 880.050 ;
        RECT 719.100 877.950 721.200 880.050 ;
        RECT 730.950 877.950 733.050 880.050 ;
        RECT 737.400 879.600 738.600 895.950 ;
        RECT 776.400 894.600 777.600 898.950 ;
        RECT 788.400 895.050 789.600 898.950 ;
        RECT 776.400 893.400 780.600 894.600 ;
        RECT 769.950 885.600 772.050 889.050 ;
        RECT 775.950 885.600 778.050 886.050 ;
        RECT 769.950 885.000 778.050 885.600 ;
        RECT 770.400 884.400 778.050 885.000 ;
        RECT 775.950 883.950 778.050 884.400 ;
        RECT 779.400 880.050 780.600 893.400 ;
        RECT 787.800 892.950 789.900 895.050 ;
        RECT 788.400 889.050 789.600 892.950 ;
        RECT 808.950 889.950 811.050 892.050 ;
        RECT 787.950 886.950 790.050 889.050 ;
        RECT 809.400 885.600 810.600 889.950 ;
        RECT 803.400 884.400 810.600 885.600 ;
        RECT 803.400 880.050 804.600 884.400 ;
        RECT 742.950 879.600 745.050 880.050 ;
        RECT 737.400 878.400 745.050 879.600 ;
        RECT 742.950 877.950 745.050 878.400 ;
        RECT 754.950 877.950 757.050 880.050 ;
        RECT 768.000 879.600 772.050 880.050 ;
        RECT 767.400 877.950 772.050 879.600 ;
        RECT 778.950 877.950 781.050 880.050 ;
        RECT 784.950 877.950 787.050 880.050 ;
        RECT 796.950 877.950 799.050 880.050 ;
        RECT 802.950 877.950 805.050 880.050 ;
        RECT 808.950 877.950 811.050 880.050 ;
        RECT 709.950 871.950 712.050 874.050 ;
        RECT 697.950 865.950 700.050 868.050 ;
        RECT 689.400 863.400 693.600 864.600 ;
        RECT 685.950 853.950 688.050 856.050 ;
        RECT 689.400 850.050 690.600 863.400 ;
        RECT 691.950 859.950 694.050 862.050 ;
        RECT 688.950 847.950 691.050 850.050 ;
        RECT 672.000 843.600 676.050 844.050 ;
        RECT 671.400 841.950 676.050 843.600 ;
        RECT 679.950 841.950 682.050 844.050 ;
        RECT 667.950 826.950 670.050 829.050 ;
        RECT 661.950 817.950 664.050 820.050 ;
        RECT 661.950 781.950 664.050 784.050 ;
        RECT 662.400 769.050 663.600 781.950 ;
        RECT 668.400 772.050 669.600 826.950 ;
        RECT 671.400 817.050 672.600 841.950 ;
        RECT 682.950 834.600 685.050 835.050 ;
        RECT 688.950 834.600 691.050 835.050 ;
        RECT 682.950 833.400 691.050 834.600 ;
        RECT 682.950 832.950 685.050 833.400 ;
        RECT 688.950 832.950 691.050 833.400 ;
        RECT 676.950 829.950 679.050 832.050 ;
        RECT 677.400 820.050 678.600 829.950 ;
        RECT 676.950 817.950 679.050 820.050 ;
        RECT 670.950 814.950 673.050 817.050 ;
        RECT 683.400 811.050 684.600 832.950 ;
        RECT 692.400 814.050 693.600 859.950 ;
        RECT 698.400 859.050 699.600 865.950 ;
        RECT 703.950 862.950 706.050 865.050 ;
        RECT 697.950 856.950 700.050 859.050 ;
        RECT 704.400 844.050 705.600 862.950 ;
        RECT 703.950 841.950 706.050 844.050 ;
        RECT 706.950 835.950 709.050 838.050 ;
        RECT 707.400 826.050 708.600 835.950 ;
        RECT 700.950 823.950 703.050 826.050 ;
        RECT 706.950 823.950 709.050 826.050 ;
        RECT 691.950 811.950 694.050 814.050 ;
        RECT 697.950 811.950 700.050 814.050 ;
        RECT 670.950 807.600 673.050 808.050 ;
        RECT 676.950 807.600 679.050 811.050 ;
        RECT 682.950 808.950 685.050 811.050 ;
        RECT 670.950 807.000 679.050 807.600 ;
        RECT 688.950 807.600 691.050 808.050 ;
        RECT 694.950 807.600 697.050 808.050 ;
        RECT 670.950 806.400 678.600 807.000 ;
        RECT 688.950 806.400 697.050 807.600 ;
        RECT 670.950 805.950 673.050 806.400 ;
        RECT 688.950 805.950 691.050 806.400 ;
        RECT 694.950 805.950 697.050 806.400 ;
        RECT 671.400 787.200 672.600 805.950 ;
        RECT 682.950 799.950 685.050 802.050 ;
        RECT 683.400 790.050 684.600 799.950 ;
        RECT 695.400 796.050 696.600 805.950 ;
        RECT 698.400 802.050 699.600 811.950 ;
        RECT 697.950 799.950 700.050 802.050 ;
        RECT 701.400 799.050 702.600 823.950 ;
        RECT 703.950 820.950 706.050 823.050 ;
        RECT 704.400 811.050 705.600 820.950 ;
        RECT 710.400 817.050 711.600 871.950 ;
        RECT 719.400 856.050 720.600 877.950 ;
        RECT 724.950 859.950 727.050 862.050 ;
        RECT 718.800 853.950 720.900 856.050 ;
        RECT 722.100 853.950 724.200 856.050 ;
        RECT 715.950 850.950 718.050 853.050 ;
        RECT 716.400 841.050 717.600 850.950 ;
        RECT 722.400 847.050 723.600 853.950 ;
        RECT 718.950 845.400 723.600 847.050 ;
        RECT 718.950 844.950 723.000 845.400 ;
        RECT 715.950 838.950 718.050 841.050 ;
        RECT 725.400 832.050 726.600 859.950 ;
        RECT 731.400 859.050 732.600 877.950 ;
        RECT 736.950 868.950 739.050 871.050 ;
        RECT 727.800 856.950 729.900 859.050 ;
        RECT 731.100 856.950 733.200 859.050 ;
        RECT 728.400 841.050 729.600 856.950 ;
        RECT 727.950 838.950 730.050 841.050 ;
        RECT 724.950 829.950 727.050 832.050 ;
        RECT 715.950 828.600 720.000 829.050 ;
        RECT 715.950 826.950 720.600 828.600 ;
        RECT 719.400 817.050 720.600 826.950 ;
        RECT 737.400 826.200 738.600 868.950 ;
        RECT 743.400 844.050 744.600 877.950 ;
        RECT 755.400 865.050 756.600 877.950 ;
        RECT 767.400 871.050 768.600 877.950 ;
        RECT 766.950 868.950 769.050 871.050 ;
        RECT 754.950 862.950 757.050 865.050 ;
        RECT 749.100 850.950 751.200 853.050 ;
        RECT 749.400 844.050 750.600 850.950 ;
        RECT 742.950 841.950 745.050 844.050 ;
        RECT 748.950 841.950 751.050 844.050 ;
        RECT 737.100 824.100 739.200 826.200 ;
        RECT 755.400 826.050 756.600 862.950 ;
        RECT 763.950 853.950 766.050 856.050 ;
        RECT 764.400 829.050 765.600 853.950 ;
        RECT 775.950 850.950 778.050 853.050 ;
        RECT 776.400 844.050 777.600 850.950 ;
        RECT 775.950 841.950 778.050 844.050 ;
        RECT 766.950 838.950 769.050 841.050 ;
        RECT 763.800 826.950 765.900 829.050 ;
        RECT 767.400 826.050 768.600 838.950 ;
        RECT 785.400 829.050 786.600 877.950 ;
        RECT 797.400 858.600 798.600 877.950 ;
        RECT 809.400 874.050 810.600 877.950 ;
        RECT 827.400 877.050 828.600 898.950 ;
        RECT 832.950 889.950 835.050 892.050 ;
        RECT 865.950 889.950 868.050 892.050 ;
        RECT 820.950 874.950 823.050 877.050 ;
        RECT 826.950 874.950 829.050 877.050 ;
        RECT 808.950 871.950 811.050 874.050 ;
        RECT 821.400 868.050 822.600 874.950 ;
        RECT 826.950 868.950 829.050 871.050 ;
        RECT 820.950 865.950 823.050 868.050 ;
        RECT 799.950 858.600 802.050 859.050 ;
        RECT 797.400 857.400 802.050 858.600 ;
        RECT 799.950 856.950 802.050 857.400 ;
        RECT 800.400 844.050 801.600 856.950 ;
        RECT 805.950 853.950 808.050 856.050 ;
        RECT 817.950 853.950 820.050 856.050 ;
        RECT 799.950 841.950 802.050 844.050 ;
        RECT 787.950 838.950 790.050 841.050 ;
        RECT 788.400 834.600 789.600 838.950 ;
        RECT 788.400 833.400 795.600 834.600 ;
        RECT 790.950 829.950 793.050 832.050 ;
        RECT 784.950 826.950 787.050 829.050 ;
        RECT 745.950 823.950 748.050 826.050 ;
        RECT 754.950 823.950 757.050 826.050 ;
        RECT 766.950 823.950 769.050 826.050 ;
        RECT 736.950 820.800 739.050 822.900 ;
        RECT 709.950 814.950 712.050 817.050 ;
        RECT 718.950 814.950 721.050 817.050 ;
        RECT 703.950 808.950 706.050 811.050 ;
        RECT 715.950 807.600 718.050 808.050 ;
        RECT 704.400 806.400 718.050 807.600 ;
        RECT 700.950 796.950 703.050 799.050 ;
        RECT 694.950 793.950 697.050 796.050 ;
        RECT 682.950 787.950 685.050 790.050 ;
        RECT 694.950 787.950 697.050 790.050 ;
        RECT 670.950 785.100 673.050 787.200 ;
        RECT 670.950 781.800 673.050 783.900 ;
        RECT 667.950 769.950 670.050 772.050 ;
        RECT 661.950 766.950 664.050 769.050 ;
        RECT 656.400 758.400 660.600 759.600 ;
        RECT 649.800 742.950 651.900 745.050 ;
        RECT 653.100 742.950 655.200 745.050 ;
        RECT 646.950 736.950 649.050 739.050 ;
        RECT 650.400 733.050 651.600 742.950 ;
        RECT 656.400 739.050 657.600 758.400 ;
        RECT 662.400 756.600 663.600 766.950 ;
        RECT 671.400 763.050 672.600 781.800 ;
        RECT 676.950 775.950 679.050 778.050 ;
        RECT 670.950 760.950 673.050 763.050 ;
        RECT 659.400 756.000 663.600 756.600 ;
        RECT 658.950 755.400 663.600 756.000 ;
        RECT 658.950 751.950 661.050 755.400 ;
        RECT 664.950 751.950 667.050 754.050 ;
        RECT 665.400 748.050 666.600 751.950 ;
        RECT 664.950 745.950 667.050 748.050 ;
        RECT 677.400 747.600 678.600 775.950 ;
        RECT 688.950 769.950 691.050 772.050 ;
        RECT 689.400 766.050 690.600 769.950 ;
        RECT 682.950 762.600 685.050 766.050 ;
        RECT 688.950 763.950 691.050 766.050 ;
        RECT 695.400 762.600 696.600 787.950 ;
        RECT 704.400 784.050 705.600 806.400 ;
        RECT 715.950 805.950 718.050 806.400 ;
        RECT 706.950 798.600 709.050 799.200 ;
        RECT 737.400 799.050 738.600 820.800 ;
        RECT 712.950 798.600 715.050 799.050 ;
        RECT 706.950 797.400 715.050 798.600 ;
        RECT 706.950 797.100 709.050 797.400 ;
        RECT 712.950 796.950 715.050 797.400 ;
        RECT 718.950 796.950 721.050 799.050 ;
        RECT 729.000 798.600 733.050 799.050 ;
        RECT 728.400 796.950 733.050 798.600 ;
        RECT 736.950 796.950 739.050 799.050 ;
        RECT 706.950 793.800 709.050 795.900 ;
        RECT 707.400 786.600 708.600 793.800 ;
        RECT 707.400 786.000 711.600 786.600 ;
        RECT 707.400 785.400 712.050 786.000 ;
        RECT 703.950 781.950 706.050 784.050 ;
        RECT 709.950 781.950 712.050 785.400 ;
        RECT 712.950 784.950 715.050 787.050 ;
        RECT 704.400 772.050 705.600 781.950 ;
        RECT 706.950 778.950 709.050 781.050 ;
        RECT 703.950 769.950 706.050 772.050 ;
        RECT 700.950 766.950 703.050 769.050 ;
        RECT 682.950 762.000 687.600 762.600 ;
        RECT 683.400 761.400 687.600 762.000 ;
        RECT 679.950 754.950 682.050 757.050 ;
        RECT 680.400 751.200 681.600 754.950 ;
        RECT 679.950 749.100 682.050 751.200 ;
        RECT 686.400 748.050 687.600 761.400 ;
        RECT 692.400 761.400 696.600 762.600 ;
        RECT 692.400 759.600 693.600 761.400 ;
        RECT 689.400 758.400 693.600 759.600 ;
        RECT 689.400 751.050 690.600 758.400 ;
        RECT 691.950 756.600 694.050 757.050 ;
        RECT 697.950 756.600 700.050 757.050 ;
        RECT 691.950 755.400 700.050 756.600 ;
        RECT 691.950 754.950 694.050 755.400 ;
        RECT 697.950 754.950 700.050 755.400 ;
        RECT 688.950 748.950 691.050 751.050 ;
        RECT 674.400 746.400 678.600 747.600 ;
        RECT 655.950 736.950 658.050 739.050 ;
        RECT 674.400 736.050 675.600 746.400 ;
        RECT 679.950 745.800 682.050 747.900 ;
        RECT 685.950 745.950 688.050 748.050 ;
        RECT 661.950 733.950 664.050 736.050 ;
        RECT 673.950 733.950 676.050 736.050 ;
        RECT 649.950 730.950 652.050 733.050 ;
        RECT 655.950 730.950 658.050 733.050 ;
        RECT 652.950 727.950 655.050 730.050 ;
        RECT 653.400 721.050 654.600 727.950 ;
        RECT 637.950 718.950 640.050 721.050 ;
        RECT 643.950 718.950 646.050 721.050 ;
        RECT 652.950 718.950 655.050 721.050 ;
        RECT 638.400 712.050 639.600 718.950 ;
        RECT 637.950 709.950 640.050 712.050 ;
        RECT 644.400 709.050 645.600 718.950 ;
        RECT 649.950 709.950 652.050 712.050 ;
        RECT 643.950 706.950 646.050 709.050 ;
        RECT 644.400 700.050 645.600 706.950 ;
        RECT 650.400 700.050 651.600 709.950 ;
        RECT 643.950 697.950 646.050 700.050 ;
        RECT 649.950 697.950 652.050 700.050 ;
        RECT 652.950 691.950 655.050 694.050 ;
        RECT 653.400 688.050 654.600 691.950 ;
        RECT 646.950 687.600 651.000 688.050 ;
        RECT 646.950 685.950 651.600 687.600 ;
        RECT 652.950 685.950 655.050 688.050 ;
        RECT 650.400 684.600 651.600 685.950 ;
        RECT 650.400 683.400 654.600 684.600 ;
        RECT 643.950 676.950 646.050 679.050 ;
        RECT 644.400 673.050 645.600 676.950 ;
        RECT 649.950 673.950 652.050 676.050 ;
        RECT 634.950 670.950 637.050 673.050 ;
        RECT 643.800 670.950 645.900 673.050 ;
        RECT 647.100 670.950 649.200 673.050 ;
        RECT 631.950 667.950 634.050 670.050 ;
        RECT 625.950 658.950 628.050 661.050 ;
        RECT 613.950 655.950 616.050 658.050 ;
        RECT 622.950 655.950 625.050 658.050 ;
        RECT 623.400 652.050 624.600 655.950 ;
        RECT 610.950 649.950 613.050 652.050 ;
        RECT 616.950 649.950 619.050 652.050 ;
        RECT 622.950 649.950 625.050 652.050 ;
        RECT 611.400 628.050 612.600 649.950 ;
        RECT 610.950 625.950 613.050 628.050 ;
        RECT 617.400 616.050 618.600 649.950 ;
        RECT 626.400 643.050 627.600 658.950 ;
        RECT 619.950 640.950 622.050 643.050 ;
        RECT 625.950 640.950 628.050 643.050 ;
        RECT 620.400 637.050 621.600 640.950 ;
        RECT 632.400 637.050 633.600 667.950 ;
        RECT 644.400 661.050 645.600 670.950 ;
        RECT 637.950 658.950 640.050 661.050 ;
        RECT 643.950 658.950 646.050 661.050 ;
        RECT 638.400 652.050 639.600 658.950 ;
        RECT 637.950 649.950 640.050 652.050 ;
        RECT 643.950 640.950 646.050 643.050 ;
        RECT 619.950 634.950 622.050 637.050 ;
        RECT 631.950 634.950 634.050 637.050 ;
        RECT 637.950 634.950 640.050 637.050 ;
        RECT 616.950 613.950 619.050 616.050 ;
        RECT 622.950 613.950 625.050 616.050 ;
        RECT 623.400 610.050 624.600 613.950 ;
        RECT 553.950 607.950 556.050 610.050 ;
        RECT 559.950 608.400 564.600 610.050 ;
        RECT 559.950 607.950 564.000 608.400 ;
        RECT 577.950 607.950 580.050 610.050 ;
        RECT 583.950 609.600 588.000 610.050 ;
        RECT 583.950 607.950 588.600 609.600 ;
        RECT 598.950 607.950 601.050 610.050 ;
        RECT 604.950 607.950 607.050 610.050 ;
        RECT 622.950 607.950 625.050 610.050 ;
        RECT 532.950 598.950 535.050 601.050 ;
        RECT 538.950 598.950 541.050 601.050 ;
        RECT 539.400 586.050 540.600 598.950 ;
        RECT 554.400 595.050 555.600 607.950 ;
        RECT 556.950 600.600 561.000 601.050 ;
        RECT 556.950 598.950 561.600 600.600 ;
        RECT 580.950 598.950 583.050 601.050 ;
        RECT 553.950 592.950 556.050 595.050 ;
        RECT 560.400 592.050 561.600 598.950 ;
        RECT 574.950 595.950 577.050 598.050 ;
        RECT 559.950 589.950 562.050 592.050 ;
        RECT 556.950 586.950 559.050 589.050 ;
        RECT 538.950 583.950 541.050 586.050 ;
        RECT 544.950 583.950 547.050 586.050 ;
        RECT 529.950 580.950 532.050 583.050 ;
        RECT 530.400 574.050 531.600 580.950 ;
        RECT 529.950 571.950 532.050 574.050 ;
        RECT 538.950 571.950 541.050 574.050 ;
        RECT 526.950 562.950 529.050 565.050 ;
        RECT 532.950 562.950 535.050 565.050 ;
        RECT 527.400 559.050 528.600 562.950 ;
        RECT 520.950 556.950 523.050 559.050 ;
        RECT 526.950 556.950 529.050 559.050 ;
        RECT 533.400 550.050 534.600 562.950 ;
        RECT 532.950 547.950 535.050 550.050 ;
        RECT 517.950 544.950 520.050 547.050 ;
        RECT 508.950 538.950 511.050 541.050 ;
        RECT 509.400 532.050 510.600 538.950 ;
        RECT 518.400 532.050 519.600 544.950 ;
        RECT 539.400 544.050 540.600 571.950 ;
        RECT 545.400 556.050 546.600 583.950 ;
        RECT 557.400 583.050 558.600 586.950 ;
        RECT 556.950 580.950 559.050 583.050 ;
        RECT 553.950 577.950 556.050 580.050 ;
        RECT 554.400 574.050 555.600 577.950 ;
        RECT 553.950 571.950 556.050 574.050 ;
        RECT 557.400 565.050 558.600 580.950 ;
        RECT 575.400 580.050 576.600 595.950 ;
        RECT 581.400 592.050 582.600 598.950 ;
        RECT 587.400 595.050 588.600 607.950 ;
        RECT 586.950 592.950 589.050 595.050 ;
        RECT 580.950 589.950 583.050 592.050 ;
        RECT 589.950 589.950 592.050 592.050 ;
        RECT 574.950 577.950 577.050 580.050 ;
        RECT 580.950 577.950 583.050 580.050 ;
        RECT 574.950 571.950 577.050 574.050 ;
        RECT 550.950 562.950 553.050 565.050 ;
        RECT 556.950 562.950 559.050 565.050 ;
        RECT 565.950 562.950 568.050 565.050 ;
        RECT 544.950 553.950 547.050 556.050 ;
        RECT 551.400 550.050 552.600 562.950 ;
        RECT 566.400 553.050 567.600 562.950 ;
        RECT 568.950 553.950 571.050 556.050 ;
        RECT 565.950 550.950 568.050 553.050 ;
        RECT 550.950 547.950 553.050 550.050 ;
        RECT 538.950 541.950 541.050 544.050 ;
        RECT 559.950 541.950 562.050 544.050 ;
        RECT 538.950 535.950 541.050 538.050 ;
        RECT 508.950 529.950 511.050 532.050 ;
        RECT 514.950 530.400 519.600 532.050 ;
        RECT 514.950 529.950 519.000 530.400 ;
        RECT 535.950 529.950 538.050 532.050 ;
        RECT 511.950 520.950 514.050 523.050 ;
        RECT 532.950 520.950 535.050 523.050 ;
        RECT 512.400 517.050 513.600 520.950 ;
        RECT 511.950 514.950 514.050 517.050 ;
        RECT 502.950 508.950 505.050 511.050 ;
        RECT 503.400 496.050 504.600 508.950 ;
        RECT 533.400 508.050 534.600 520.950 ;
        RECT 505.950 505.950 508.050 508.050 ;
        RECT 532.950 505.950 535.050 508.050 ;
        RECT 506.400 496.050 507.600 505.950 ;
        RECT 536.400 505.050 537.600 529.950 ;
        RECT 535.950 502.950 538.050 505.050 ;
        RECT 523.950 499.950 526.050 502.050 ;
        RECT 524.400 496.050 525.600 499.950 ;
        RECT 539.400 496.050 540.600 535.950 ;
        RECT 544.950 532.050 547.050 535.050 ;
        RECT 553.950 532.950 556.050 535.050 ;
        RECT 541.950 531.000 547.050 532.050 ;
        RECT 541.950 530.400 546.600 531.000 ;
        RECT 541.950 529.950 546.000 530.400 ;
        RECT 544.950 522.600 547.050 523.050 ;
        RECT 550.950 522.600 553.050 523.050 ;
        RECT 544.950 521.400 553.050 522.600 ;
        RECT 544.950 520.950 547.050 521.400 ;
        RECT 550.950 520.950 553.050 521.400 ;
        RECT 554.400 511.050 555.600 532.950 ;
        RECT 560.400 532.050 561.600 541.950 ;
        RECT 565.950 535.950 568.050 538.050 ;
        RECT 560.400 530.400 565.050 532.050 ;
        RECT 561.000 529.950 565.050 530.400 ;
        RECT 566.400 523.050 567.600 535.950 ;
        RECT 569.400 532.050 570.600 553.950 ;
        RECT 575.400 553.050 576.600 571.950 ;
        RECT 577.950 559.950 580.050 562.050 ;
        RECT 574.800 550.950 576.900 553.050 ;
        RECT 578.400 550.050 579.600 559.950 ;
        RECT 577.950 547.950 580.050 550.050 ;
        RECT 577.950 541.950 580.050 544.050 ;
        RECT 578.400 532.050 579.600 541.950 ;
        RECT 581.400 541.050 582.600 577.950 ;
        RECT 590.400 574.050 591.600 589.950 ;
        RECT 599.400 589.050 600.600 607.950 ;
        RECT 607.950 598.950 610.050 601.050 ;
        RECT 601.950 595.950 604.050 598.050 ;
        RECT 598.950 586.950 601.050 589.050 ;
        RECT 602.400 586.050 603.600 595.950 ;
        RECT 608.400 595.050 609.600 598.950 ;
        RECT 607.950 592.950 610.050 595.050 ;
        RECT 610.950 586.950 613.050 589.050 ;
        RECT 601.950 583.950 604.050 586.050 ;
        RECT 607.950 580.950 610.050 583.050 ;
        RECT 589.950 571.950 592.050 574.050 ;
        RECT 598.950 565.950 601.050 568.050 ;
        RECT 586.950 562.950 589.050 565.050 ;
        RECT 592.950 562.950 595.050 565.050 ;
        RECT 587.400 559.050 588.600 562.950 ;
        RECT 586.950 556.950 589.050 559.050 ;
        RECT 589.950 553.950 592.050 556.050 ;
        RECT 580.950 538.950 583.050 541.050 ;
        RECT 583.950 535.950 586.050 538.050 ;
        RECT 568.950 529.950 571.050 532.050 ;
        RECT 578.400 530.400 583.050 532.050 ;
        RECT 579.000 529.950 583.050 530.400 ;
        RECT 584.400 523.050 585.600 535.950 ;
        RECT 590.400 532.050 591.600 553.950 ;
        RECT 593.400 553.050 594.600 562.950 ;
        RECT 599.400 559.050 600.600 565.950 ;
        RECT 598.950 556.950 601.050 559.050 ;
        RECT 592.950 550.950 595.050 553.050 ;
        RECT 608.400 550.050 609.600 580.950 ;
        RECT 611.400 574.050 612.600 586.950 ;
        RECT 623.400 583.050 624.600 607.950 ;
        RECT 628.950 606.600 631.050 610.050 ;
        RECT 628.950 606.000 633.600 606.600 ;
        RECT 629.400 605.400 633.600 606.000 ;
        RECT 632.400 601.050 633.600 605.400 ;
        RECT 631.950 598.950 634.050 601.050 ;
        RECT 622.950 580.950 625.050 583.050 ;
        RECT 632.400 580.050 633.600 598.950 ;
        RECT 638.400 583.050 639.600 634.950 ;
        RECT 644.400 592.050 645.600 640.950 ;
        RECT 647.400 631.050 648.600 670.950 ;
        RECT 646.950 628.950 649.050 631.050 ;
        RECT 650.400 610.050 651.600 673.950 ;
        RECT 653.400 667.050 654.600 683.400 ;
        RECT 656.400 670.050 657.600 730.950 ;
        RECT 662.400 730.050 663.600 733.950 ;
        RECT 661.950 727.950 664.050 730.050 ;
        RECT 667.950 729.600 672.000 730.050 ;
        RECT 667.950 727.950 672.600 729.600 ;
        RECT 664.950 720.600 667.050 721.050 ;
        RECT 659.400 719.400 667.050 720.600 ;
        RECT 659.400 700.200 660.600 719.400 ;
        RECT 664.950 718.950 667.050 719.400 ;
        RECT 661.950 712.950 664.050 715.050 ;
        RECT 659.100 698.100 661.200 700.200 ;
        RECT 662.400 694.050 663.600 712.950 ;
        RECT 671.400 712.050 672.600 727.950 ;
        RECT 670.950 709.950 673.050 712.050 ;
        RECT 658.800 691.950 660.900 694.050 ;
        RECT 662.100 691.950 664.200 694.050 ;
        RECT 659.400 679.200 660.600 691.950 ;
        RECT 680.400 691.050 681.600 745.800 ;
        RECT 701.400 739.050 702.600 766.950 ;
        RECT 700.950 736.950 703.050 739.050 ;
        RECT 707.400 736.050 708.600 778.950 ;
        RECT 713.400 757.050 714.600 784.950 ;
        RECT 719.400 766.050 720.600 796.950 ;
        RECT 728.400 784.050 729.600 796.950 ;
        RECT 736.950 790.950 739.050 793.050 ;
        RECT 733.950 784.950 736.050 787.050 ;
        RECT 727.950 781.950 730.050 784.050 ;
        RECT 730.950 772.950 733.050 775.050 ;
        RECT 724.950 769.950 727.050 772.050 ;
        RECT 725.400 766.050 726.600 769.950 ;
        RECT 731.400 766.050 732.600 772.950 ;
        RECT 718.950 763.950 721.050 766.050 ;
        RECT 724.950 763.950 727.050 766.050 ;
        RECT 730.950 763.950 733.050 766.050 ;
        RECT 719.400 759.600 720.600 763.950 ;
        RECT 719.400 758.400 726.600 759.600 ;
        RECT 725.400 757.050 726.600 758.400 ;
        RECT 712.950 754.950 715.050 757.050 ;
        RECT 725.400 755.400 730.050 757.050 ;
        RECT 726.000 754.950 730.050 755.400 ;
        RECT 734.400 753.600 735.600 784.950 ;
        RECT 737.400 784.050 738.600 790.950 ;
        RECT 736.950 781.950 739.050 784.050 ;
        RECT 739.950 769.800 742.050 771.900 ;
        RECT 731.400 752.400 735.600 753.600 ;
        RECT 727.950 748.950 730.050 751.050 ;
        RECT 722.100 739.950 724.200 742.050 ;
        RECT 719.100 736.800 721.200 738.900 ;
        RECT 682.950 733.950 685.050 736.050 ;
        RECT 706.950 733.950 709.050 736.050 ;
        RECT 683.400 721.050 684.600 733.950 ;
        RECT 694.950 727.950 697.050 730.050 ;
        RECT 699.000 729.600 703.050 730.050 ;
        RECT 698.400 727.950 703.050 729.600 ;
        RECT 682.950 718.950 685.050 721.050 ;
        RECT 688.950 718.950 691.050 721.050 ;
        RECT 682.950 712.950 685.050 715.050 ;
        RECT 683.400 703.050 684.600 712.950 ;
        RECT 689.400 712.050 690.600 718.950 ;
        RECT 695.400 712.050 696.600 727.950 ;
        RECT 698.400 721.050 699.600 727.950 ;
        RECT 706.950 726.600 709.050 730.050 ;
        RECT 706.950 726.000 714.600 726.600 ;
        RECT 707.400 725.400 714.600 726.000 ;
        RECT 697.950 718.950 700.050 721.050 ;
        RECT 703.950 718.950 706.050 721.050 ;
        RECT 709.950 718.950 712.050 721.050 ;
        RECT 704.400 715.050 705.600 718.950 ;
        RECT 703.950 712.950 706.050 715.050 ;
        RECT 710.400 712.050 711.600 718.950 ;
        RECT 713.400 718.050 714.600 725.400 ;
        RECT 713.400 716.400 718.050 718.050 ;
        RECT 714.000 715.950 718.050 716.400 ;
        RECT 688.950 709.950 691.050 712.050 ;
        RECT 694.950 709.950 697.050 712.050 ;
        RECT 709.950 709.950 712.050 712.050 ;
        RECT 719.400 708.600 720.600 736.800 ;
        RECT 716.400 707.400 720.600 708.600 ;
        RECT 685.950 703.950 688.050 706.050 ;
        RECT 682.950 700.950 685.050 703.050 ;
        RECT 679.950 688.950 682.050 691.050 ;
        RECT 667.950 685.950 670.050 688.050 ;
        RECT 658.950 677.100 661.050 679.200 ;
        RECT 658.950 673.800 661.050 675.900 ;
        RECT 655.950 667.950 658.050 670.050 ;
        RECT 652.950 664.950 655.050 667.050 ;
        RECT 653.400 637.050 654.600 664.950 ;
        RECT 655.950 658.950 658.050 661.050 ;
        RECT 656.400 652.050 657.600 658.950 ;
        RECT 655.950 649.950 658.050 652.050 ;
        RECT 659.400 645.600 660.600 673.800 ;
        RECT 668.400 670.050 669.600 685.950 ;
        RECT 667.950 667.950 670.050 670.050 ;
        RECT 679.950 667.950 682.050 670.050 ;
        RECT 680.400 646.050 681.600 667.950 ;
        RECT 686.400 664.200 687.600 703.950 ;
        RECT 716.400 697.050 717.600 707.400 ;
        RECT 722.400 697.050 723.600 739.950 ;
        RECT 728.400 739.050 729.600 748.950 ;
        RECT 731.400 742.050 732.600 752.400 ;
        RECT 733.950 748.950 736.050 751.050 ;
        RECT 730.950 739.950 733.050 742.050 ;
        RECT 724.800 736.950 726.900 739.050 ;
        RECT 728.100 736.950 730.200 739.050 ;
        RECT 725.400 733.050 726.600 736.950 ;
        RECT 724.950 730.950 727.050 733.050 ;
        RECT 730.950 730.950 733.050 733.050 ;
        RECT 731.400 715.200 732.600 730.950 ;
        RECT 724.950 712.950 727.050 715.050 ;
        RECT 730.950 713.100 733.050 715.200 ;
        RECT 725.400 700.050 726.600 712.950 ;
        RECT 730.950 709.800 733.050 711.900 ;
        RECT 727.950 706.950 730.050 709.050 ;
        RECT 724.950 697.950 727.050 700.050 ;
        RECT 715.950 694.950 718.050 697.050 ;
        RECT 721.950 694.950 724.050 697.050 ;
        RECT 691.950 688.950 694.050 691.050 ;
        RECT 692.400 676.050 693.600 688.950 ;
        RECT 709.950 688.050 712.050 691.050 ;
        RECT 709.950 687.000 715.050 688.050 ;
        RECT 710.400 686.400 715.050 687.000 ;
        RECT 711.000 685.950 715.050 686.400 ;
        RECT 718.950 687.600 721.050 688.050 ;
        RECT 718.950 686.400 726.600 687.600 ;
        RECT 718.950 685.950 721.050 686.400 ;
        RECT 703.950 682.950 706.050 685.050 ;
        RECT 691.950 673.950 694.050 676.050 ;
        RECT 697.950 673.950 700.050 676.050 ;
        RECT 685.950 662.100 688.050 664.200 ;
        RECT 656.400 644.400 660.600 645.600 ;
        RECT 652.950 634.950 655.050 637.050 ;
        RECT 656.400 616.050 657.600 644.400 ;
        RECT 679.950 643.950 682.050 646.050 ;
        RECT 658.950 640.950 661.050 643.050 ;
        RECT 664.950 640.950 667.050 643.050 ;
        RECT 659.400 637.050 660.600 640.950 ;
        RECT 665.400 637.050 666.600 640.950 ;
        RECT 692.400 640.050 693.600 673.950 ;
        RECT 698.400 670.050 699.600 673.950 ;
        RECT 704.400 673.050 705.600 682.950 ;
        RECT 709.950 676.950 712.050 679.050 ;
        RECT 703.950 670.950 706.050 673.050 ;
        RECT 710.400 670.050 711.600 676.950 ;
        RECT 697.950 667.950 700.050 670.050 ;
        RECT 709.950 667.950 712.050 670.050 ;
        RECT 718.950 667.950 721.050 670.050 ;
        RECT 691.950 637.950 694.050 640.050 ;
        RECT 658.950 634.950 661.050 637.050 ;
        RECT 664.950 634.950 667.050 637.050 ;
        RECT 673.950 634.950 676.050 637.050 ;
        RECT 667.950 625.950 670.050 628.050 ;
        RECT 664.950 616.950 667.050 619.050 ;
        RECT 655.950 613.950 658.050 616.050 ;
        RECT 665.400 610.050 666.600 616.950 ;
        RECT 646.950 607.950 649.050 610.050 ;
        RECT 650.400 608.400 655.050 610.050 ;
        RECT 651.000 607.950 655.050 608.400 ;
        RECT 664.950 607.950 667.050 610.050 ;
        RECT 647.400 595.050 648.600 607.950 ;
        RECT 649.950 598.950 652.050 601.050 ;
        RECT 646.950 592.950 649.050 595.050 ;
        RECT 643.950 589.950 646.050 592.050 ;
        RECT 637.950 580.950 640.050 583.050 ;
        RECT 619.950 577.950 622.050 580.050 ;
        RECT 631.950 577.950 634.050 580.050 ;
        RECT 640.950 577.950 643.050 580.050 ;
        RECT 620.400 574.050 621.600 577.950 ;
        RECT 622.950 574.950 625.050 577.050 ;
        RECT 610.950 571.950 613.050 574.050 ;
        RECT 616.950 572.400 621.600 574.050 ;
        RECT 616.950 571.950 621.000 572.400 ;
        RECT 623.400 568.050 624.600 574.950 ;
        RECT 625.950 571.950 628.050 574.050 ;
        RECT 622.950 565.950 625.050 568.050 ;
        RECT 607.950 547.950 610.050 550.050 ;
        RECT 626.400 541.050 627.600 571.950 ;
        RECT 641.400 565.050 642.600 577.950 ;
        RECT 634.950 562.950 637.050 565.050 ;
        RECT 640.950 562.950 643.050 565.050 ;
        RECT 635.400 559.050 636.600 562.950 ;
        RECT 647.400 559.050 648.600 592.950 ;
        RECT 650.400 592.050 651.600 598.950 ;
        RECT 649.950 589.950 652.050 592.050 ;
        RECT 661.950 589.950 664.050 592.050 ;
        RECT 652.950 577.950 655.050 580.050 ;
        RECT 634.950 556.950 637.050 559.050 ;
        RECT 646.950 556.950 649.050 559.050 ;
        RECT 653.400 553.050 654.600 577.950 ;
        RECT 662.400 574.050 663.600 589.950 ;
        RECT 668.400 585.600 669.600 625.950 ;
        RECT 674.400 610.050 675.600 634.950 ;
        RECT 698.400 628.050 699.600 667.950 ;
        RECT 715.950 664.950 718.050 667.050 ;
        RECT 709.950 661.950 712.050 664.050 ;
        RECT 703.950 658.950 706.050 661.050 ;
        RECT 704.400 655.050 705.600 658.950 ;
        RECT 710.400 655.050 711.600 661.950 ;
        RECT 703.950 652.950 706.050 655.050 ;
        RECT 709.950 652.950 712.050 655.050 ;
        RECT 700.950 634.950 703.050 637.050 ;
        RECT 701.400 631.050 702.600 634.950 ;
        RECT 700.950 628.950 703.050 631.050 ;
        RECT 704.400 628.050 705.600 652.950 ;
        RECT 709.950 643.950 712.050 646.050 ;
        RECT 697.950 625.950 700.050 628.050 ;
        RECT 703.950 625.950 706.050 628.050 ;
        RECT 706.950 616.950 709.050 619.050 ;
        RECT 697.950 610.050 700.050 613.050 ;
        RECT 670.950 608.400 675.600 610.050 ;
        RECT 670.950 607.950 675.000 608.400 ;
        RECT 688.950 607.950 691.050 610.050 ;
        RECT 694.950 609.000 700.050 610.050 ;
        RECT 694.950 608.400 699.600 609.000 ;
        RECT 694.950 607.950 699.000 608.400 ;
        RECT 673.950 598.950 676.050 601.050 ;
        RECT 665.400 584.400 669.600 585.600 ;
        RECT 661.950 571.950 664.050 574.050 ;
        RECT 665.400 565.050 666.600 584.400 ;
        RECT 667.950 580.950 670.050 583.050 ;
        RECT 668.400 574.050 669.600 580.950 ;
        RECT 667.950 571.950 670.050 574.050 ;
        RECT 658.950 562.950 661.050 565.050 ;
        RECT 664.950 562.950 667.050 565.050 ;
        RECT 634.950 550.950 637.050 553.050 ;
        RECT 652.950 550.950 655.050 553.050 ;
        RECT 607.950 538.950 610.050 541.050 ;
        RECT 625.950 538.950 628.050 541.050 ;
        RECT 586.950 530.400 591.600 532.050 ;
        RECT 586.950 529.950 591.000 530.400 ;
        RECT 608.400 525.600 609.600 538.950 ;
        RECT 635.400 532.050 636.600 550.950 ;
        RECT 653.400 532.050 654.600 550.950 ;
        RECT 659.400 550.050 660.600 562.950 ;
        RECT 668.400 561.600 669.600 571.950 ;
        RECT 665.400 560.400 669.600 561.600 ;
        RECT 658.950 547.950 661.050 550.050 ;
        RECT 622.950 531.600 625.050 532.050 ;
        RECT 628.950 531.600 631.050 532.050 ;
        RECT 622.950 530.400 633.600 531.600 ;
        RECT 622.950 529.950 625.050 530.400 ;
        RECT 628.950 529.950 631.050 530.400 ;
        RECT 605.400 525.000 609.600 525.600 ;
        RECT 604.950 524.400 609.600 525.000 ;
        RECT 632.400 525.600 633.600 530.400 ;
        RECT 634.950 529.950 637.050 532.050 ;
        RECT 652.950 529.950 655.050 532.050 ;
        RECT 657.000 531.600 661.050 532.050 ;
        RECT 656.400 529.950 661.050 531.600 ;
        RECT 646.950 528.600 649.050 529.050 ;
        RECT 656.400 528.600 657.600 529.950 ;
        RECT 646.950 527.400 657.600 528.600 ;
        RECT 646.950 526.950 649.050 527.400 ;
        RECT 637.950 525.600 640.050 526.050 ;
        RECT 632.400 524.400 640.050 525.600 ;
        RECT 565.950 520.950 568.050 523.050 ;
        RECT 583.950 520.950 586.050 523.050 ;
        RECT 598.950 520.950 601.050 523.050 ;
        RECT 604.950 520.950 607.050 524.400 ;
        RECT 637.950 523.950 640.050 524.400 ;
        RECT 610.950 520.950 613.050 523.050 ;
        RECT 631.950 522.600 636.000 523.050 ;
        RECT 631.950 520.950 636.600 522.600 ;
        RECT 646.950 520.950 649.050 523.050 ;
        RECT 655.950 522.600 660.000 523.050 ;
        RECT 655.950 522.000 660.600 522.600 ;
        RECT 655.950 520.950 661.050 522.000 ;
        RECT 599.400 517.050 600.600 520.950 ;
        RECT 592.950 514.950 595.050 517.050 ;
        RECT 598.950 514.950 601.050 517.050 ;
        RECT 553.950 508.950 556.050 511.050 ;
        RECT 544.950 505.950 547.050 508.050 ;
        RECT 499.950 494.400 504.600 496.050 ;
        RECT 499.950 493.950 504.000 494.400 ;
        RECT 505.950 493.950 508.050 496.050 ;
        RECT 523.950 493.950 526.050 496.050 ;
        RECT 538.950 493.950 541.050 496.050 ;
        RECT 515.400 489.000 528.600 489.600 ;
        RECT 514.950 488.400 528.600 489.000 ;
        RECT 496.950 484.950 499.050 487.050 ;
        RECT 502.950 486.600 505.050 487.050 ;
        RECT 508.950 486.600 511.050 487.050 ;
        RECT 502.950 485.400 511.050 486.600 ;
        RECT 502.950 484.950 505.050 485.400 ;
        RECT 508.950 484.950 511.050 485.400 ;
        RECT 514.950 484.950 517.050 488.400 ;
        RECT 527.400 487.050 528.600 488.400 ;
        RECT 520.950 484.950 523.050 487.050 ;
        RECT 526.950 486.600 529.050 487.050 ;
        RECT 532.950 486.600 535.050 487.050 ;
        RECT 526.950 485.400 535.050 486.600 ;
        RECT 526.950 484.950 529.050 485.400 ;
        RECT 532.950 484.950 535.050 485.400 ;
        RECT 521.400 481.050 522.600 484.950 ;
        RECT 545.400 481.050 546.600 505.950 ;
        RECT 593.400 502.050 594.600 514.950 ;
        RECT 565.950 499.950 568.050 502.050 ;
        RECT 592.950 499.950 595.050 502.050 ;
        RECT 555.000 495.600 559.050 496.050 ;
        RECT 554.400 493.950 559.050 495.600 ;
        RECT 554.400 487.050 555.600 493.950 ;
        RECT 566.400 487.050 567.600 499.950 ;
        RECT 599.400 498.600 600.600 514.950 ;
        RECT 611.400 511.050 612.600 520.950 ;
        RECT 635.400 520.050 636.600 520.950 ;
        RECT 635.400 518.400 640.050 520.050 ;
        RECT 636.000 517.950 640.050 518.400 ;
        RECT 610.950 508.950 613.050 511.050 ;
        RECT 647.400 505.050 648.600 520.950 ;
        RECT 658.950 517.950 661.050 520.950 ;
        RECT 665.400 514.050 666.600 560.400 ;
        RECT 674.400 556.050 675.600 598.950 ;
        RECT 689.400 589.050 690.600 607.950 ;
        RECT 707.400 601.050 708.600 616.950 ;
        RECT 710.400 610.050 711.600 643.950 ;
        RECT 716.400 619.050 717.600 664.950 ;
        RECT 719.400 651.600 720.600 667.950 ;
        RECT 725.400 664.050 726.600 686.400 ;
        RECT 728.400 667.050 729.600 706.950 ;
        RECT 731.400 694.050 732.600 709.800 ;
        RECT 730.950 691.950 733.050 694.050 ;
        RECT 730.950 682.950 733.050 685.050 ;
        RECT 727.950 664.950 730.050 667.050 ;
        RECT 724.950 661.950 727.050 664.050 ;
        RECT 731.400 661.050 732.600 682.950 ;
        RECT 734.400 661.200 735.600 748.950 ;
        RECT 736.950 742.950 739.050 745.050 ;
        RECT 737.400 706.200 738.600 742.950 ;
        RECT 740.400 720.600 741.600 769.800 ;
        RECT 742.950 739.950 745.050 742.050 ;
        RECT 743.400 730.050 744.600 739.950 ;
        RECT 746.400 736.050 747.600 823.950 ;
        RECT 778.950 817.950 781.050 820.050 ;
        RECT 784.950 817.950 787.050 820.050 ;
        RECT 748.950 811.950 751.050 814.050 ;
        RECT 757.950 811.950 760.050 814.050 ;
        RECT 749.400 808.050 750.600 811.950 ;
        RECT 748.950 805.950 751.050 808.050 ;
        RECT 754.950 805.950 757.050 808.050 ;
        RECT 755.400 789.600 756.600 805.950 ;
        RECT 758.400 799.050 759.600 811.950 ;
        RECT 760.950 807.600 763.050 808.050 ;
        RECT 766.950 807.600 769.050 808.050 ;
        RECT 760.950 806.400 769.050 807.600 ;
        RECT 760.950 805.950 763.050 806.400 ;
        RECT 766.950 805.950 769.050 806.400 ;
        RECT 775.950 805.950 778.050 808.050 ;
        RECT 757.950 796.950 760.050 799.050 ;
        RECT 763.950 796.950 766.050 799.050 ;
        RECT 764.400 790.050 765.600 796.950 ;
        RECT 752.400 788.400 756.600 789.600 ;
        RECT 752.400 772.050 753.600 788.400 ;
        RECT 763.950 787.950 766.050 790.050 ;
        RECT 772.950 787.950 775.050 790.050 ;
        RECT 754.950 781.950 757.050 784.050 ;
        RECT 755.400 778.050 756.600 781.950 ;
        RECT 754.950 775.950 757.050 778.050 ;
        RECT 751.950 769.950 754.050 772.050 ;
        RECT 766.950 769.950 769.050 772.050 ;
        RECT 767.400 766.050 768.600 769.950 ;
        RECT 773.400 766.050 774.600 787.950 ;
        RECT 776.400 772.050 777.600 805.950 ;
        RECT 779.400 799.050 780.600 817.950 ;
        RECT 785.400 799.050 786.600 817.950 ;
        RECT 778.950 796.950 781.050 799.050 ;
        RECT 784.950 796.950 787.050 799.050 ;
        RECT 791.400 796.050 792.600 829.950 ;
        RECT 794.400 802.050 795.600 833.400 ;
        RECT 799.950 832.950 802.050 835.050 ;
        RECT 800.400 820.050 801.600 832.950 ;
        RECT 806.400 820.050 807.600 853.950 ;
        RECT 818.400 844.050 819.600 853.950 ;
        RECT 811.950 841.950 814.050 844.050 ;
        RECT 817.950 841.950 820.050 844.050 ;
        RECT 812.400 828.600 813.600 841.950 ;
        RECT 823.950 838.950 826.050 841.050 ;
        RECT 814.950 832.950 817.050 835.050 ;
        RECT 815.400 829.050 816.600 832.950 ;
        RECT 809.400 827.400 813.600 828.600 ;
        RECT 799.950 817.950 802.050 820.050 ;
        RECT 805.950 817.950 808.050 820.050 ;
        RECT 796.950 814.950 799.050 817.050 ;
        RECT 802.950 814.950 805.050 817.050 ;
        RECT 793.800 799.950 795.900 802.050 ;
        RECT 797.400 801.600 798.600 814.950 ;
        RECT 803.400 808.050 804.600 814.950 ;
        RECT 802.950 805.950 805.050 808.050 ;
        RECT 797.400 800.400 801.600 801.600 ;
        RECT 797.100 796.950 799.200 799.050 ;
        RECT 800.400 798.600 801.600 800.400 ;
        RECT 809.400 799.050 810.600 827.400 ;
        RECT 814.950 826.950 817.050 829.050 ;
        RECT 815.400 823.050 816.600 826.950 ;
        RECT 824.400 826.050 825.600 838.950 ;
        RECT 817.950 823.950 820.050 826.050 ;
        RECT 823.950 823.950 826.050 826.050 ;
        RECT 814.950 820.950 817.050 823.050 ;
        RECT 818.400 810.600 819.600 823.950 ;
        RECT 827.400 817.050 828.600 868.950 ;
        RECT 833.400 856.050 834.600 889.950 ;
        RECT 866.400 886.050 867.600 889.950 ;
        RECT 835.950 885.600 838.050 886.050 ;
        RECT 841.950 885.600 844.050 886.050 ;
        RECT 835.950 884.400 844.050 885.600 ;
        RECT 835.950 883.950 838.050 884.400 ;
        RECT 841.950 883.950 844.050 884.400 ;
        RECT 859.950 883.950 862.050 886.050 ;
        RECT 865.950 883.950 868.050 886.050 ;
        RECT 844.950 874.950 847.050 877.050 ;
        RECT 845.400 871.050 846.600 874.950 ;
        RECT 844.950 868.950 847.050 871.050 ;
        RECT 832.950 853.950 835.050 856.050 ;
        RECT 835.950 850.950 838.050 853.050 ;
        RECT 829.950 831.600 832.050 835.050 ;
        RECT 836.400 832.050 837.600 850.950 ;
        RECT 860.400 850.050 861.600 883.950 ;
        RECT 886.950 882.600 889.050 886.050 ;
        RECT 886.950 882.000 891.600 882.600 ;
        RECT 887.400 881.400 891.600 882.000 ;
        RECT 883.950 874.950 886.050 877.050 ;
        RECT 884.400 871.050 885.600 874.950 ;
        RECT 883.950 868.950 886.050 871.050 ;
        RECT 865.950 850.950 868.050 853.050 ;
        RECT 859.950 847.950 862.050 850.050 ;
        RECT 866.400 844.050 867.600 850.950 ;
        RECT 871.950 847.950 874.050 850.050 ;
        RECT 858.000 843.600 862.050 844.050 ;
        RECT 857.400 841.950 862.050 843.600 ;
        RECT 865.950 841.950 868.050 844.050 ;
        RECT 844.950 838.950 847.050 841.050 ;
        RECT 835.950 831.600 838.050 832.050 ;
        RECT 829.950 831.000 838.050 831.600 ;
        RECT 830.400 830.400 838.050 831.000 ;
        RECT 835.950 829.950 838.050 830.400 ;
        RECT 841.950 829.950 844.050 832.050 ;
        RECT 842.400 826.050 843.600 829.950 ;
        RECT 835.950 823.950 838.050 826.050 ;
        RECT 841.950 823.950 844.050 826.050 ;
        RECT 826.950 814.950 829.050 817.050 ;
        RECT 823.950 811.950 826.050 814.050 ;
        RECT 815.400 810.000 819.600 810.600 ;
        RECT 814.950 809.400 819.600 810.000 ;
        RECT 814.950 805.950 817.050 809.400 ;
        RECT 820.950 805.950 823.050 808.050 ;
        RECT 800.400 797.400 804.600 798.600 ;
        RECT 790.950 793.950 793.050 796.050 ;
        RECT 778.950 790.950 781.050 793.050 ;
        RECT 779.400 778.050 780.600 790.950 ;
        RECT 793.950 784.950 796.050 787.050 ;
        RECT 790.950 778.950 793.050 781.050 ;
        RECT 778.950 775.950 781.050 778.050 ;
        RECT 775.950 769.950 778.050 772.050 ;
        RECT 784.950 769.950 787.050 772.050 ;
        RECT 766.950 763.950 769.050 766.050 ;
        RECT 772.950 763.950 775.050 766.050 ;
        RECT 748.950 754.950 751.050 757.050 ;
        RECT 757.950 754.950 760.050 757.050 ;
        RECT 749.400 739.050 750.600 754.950 ;
        RECT 758.400 745.050 759.600 754.950 ;
        RECT 757.950 742.950 760.050 745.050 ;
        RECT 772.950 739.950 775.050 742.050 ;
        RECT 748.950 736.950 751.050 739.050 ;
        RECT 745.950 733.950 748.050 736.050 ;
        RECT 763.950 733.950 766.050 736.050 ;
        RECT 769.950 733.950 772.050 736.050 ;
        RECT 743.400 728.400 748.050 730.050 ;
        RECT 744.000 727.950 748.050 728.400 ;
        RECT 757.950 724.950 760.050 727.050 ;
        RECT 758.400 721.050 759.600 724.950 ;
        RECT 740.400 719.400 744.600 720.600 ;
        RECT 739.950 715.950 742.050 718.050 ;
        RECT 736.800 704.100 738.900 706.200 ;
        RECT 740.400 706.050 741.600 715.950 ;
        RECT 743.400 709.050 744.600 719.400 ;
        RECT 748.950 718.950 751.050 721.050 ;
        RECT 754.950 719.400 759.600 721.050 ;
        RECT 754.950 718.950 759.000 719.400 ;
        RECT 749.400 712.050 750.600 718.950 ;
        RECT 755.400 715.050 756.600 718.950 ;
        RECT 754.950 712.950 757.050 715.050 ;
        RECT 748.950 709.950 751.050 712.050 ;
        RECT 757.950 709.950 760.050 712.050 ;
        RECT 742.950 706.950 745.050 709.050 ;
        RECT 754.950 706.950 757.050 709.050 ;
        RECT 740.100 703.950 742.200 706.050 ;
        RECT 755.400 697.050 756.600 706.950 ;
        RECT 758.400 700.050 759.600 709.950 ;
        RECT 764.400 700.050 765.600 733.950 ;
        RECT 770.400 721.050 771.600 733.950 ;
        RECT 769.950 718.950 772.050 721.050 ;
        RECT 766.950 709.950 769.050 712.050 ;
        RECT 767.400 706.050 768.600 709.950 ;
        RECT 766.950 703.950 769.050 706.050 ;
        RECT 773.400 703.050 774.600 739.950 ;
        RECT 785.400 723.600 786.600 769.950 ;
        RECT 791.400 766.050 792.600 778.950 ;
        RECT 794.400 772.050 795.600 784.950 ;
        RECT 793.950 769.950 796.050 772.050 ;
        RECT 797.400 766.050 798.600 796.950 ;
        RECT 803.400 796.050 804.600 797.400 ;
        RECT 808.950 796.950 811.050 799.050 ;
        RECT 817.950 796.950 820.050 799.050 ;
        RECT 803.400 794.400 808.050 796.050 ;
        RECT 804.000 793.950 808.050 794.400 ;
        RECT 802.950 790.950 805.050 793.050 ;
        RECT 790.950 763.950 793.050 766.050 ;
        RECT 796.950 763.950 799.050 766.050 ;
        RECT 787.950 754.950 790.050 757.050 ;
        RECT 788.400 742.050 789.600 754.950 ;
        RECT 787.950 739.950 790.050 742.050 ;
        RECT 803.400 736.050 804.600 790.950 ;
        RECT 818.400 790.050 819.600 796.950 ;
        RECT 817.950 787.950 820.050 790.050 ;
        RECT 821.400 772.050 822.600 805.950 ;
        RECT 824.400 799.050 825.600 811.950 ;
        RECT 823.950 796.950 826.050 799.050 ;
        RECT 836.400 793.050 837.600 823.950 ;
        RECT 838.950 811.950 841.050 814.050 ;
        RECT 839.400 808.050 840.600 811.950 ;
        RECT 838.950 805.950 841.050 808.050 ;
        RECT 845.400 801.600 846.600 838.950 ;
        RECT 847.950 832.950 850.050 835.050 ;
        RECT 842.400 801.000 846.600 801.600 ;
        RECT 841.950 800.400 846.600 801.000 ;
        RECT 841.950 796.950 844.050 800.400 ;
        RECT 848.400 799.050 849.600 832.950 ;
        RECT 857.400 832.050 858.600 841.950 ;
        RECT 856.950 829.950 859.050 832.050 ;
        RECT 865.950 826.950 868.050 829.050 ;
        RECT 850.950 823.950 853.050 826.050 ;
        RECT 847.950 796.950 850.050 799.050 ;
        RECT 835.950 790.950 838.050 793.050 ;
        RECT 820.950 769.950 823.050 772.050 ;
        RECT 808.950 765.600 811.050 766.050 ;
        RECT 814.950 765.600 817.050 766.050 ;
        RECT 808.950 764.400 817.050 765.600 ;
        RECT 808.950 763.950 811.050 764.400 ;
        RECT 814.950 763.950 817.050 764.400 ;
        RECT 820.950 765.600 823.050 766.050 ;
        RECT 826.950 765.600 829.050 769.050 ;
        RECT 820.950 765.000 829.050 765.600 ;
        RECT 820.950 764.400 828.600 765.000 ;
        RECT 820.950 763.950 823.050 764.400 ;
        RECT 811.950 754.950 814.050 757.050 ;
        RECT 823.800 754.950 825.900 757.050 ;
        RECT 808.950 739.950 811.050 742.050 ;
        RECT 802.950 733.950 805.050 736.050 ;
        RECT 793.950 727.950 796.050 730.050 ;
        RECT 785.400 722.400 789.600 723.600 ;
        RECT 788.400 721.050 789.600 722.400 ;
        RECT 788.400 719.400 793.050 721.050 ;
        RECT 789.000 718.950 793.050 719.400 ;
        RECT 787.950 706.950 790.050 709.050 ;
        RECT 772.950 700.950 775.050 703.050 ;
        RECT 757.950 697.950 760.050 700.050 ;
        RECT 763.950 697.950 766.050 700.050 ;
        RECT 742.950 694.950 745.050 697.050 ;
        RECT 754.950 694.950 757.050 697.050 ;
        RECT 743.400 688.050 744.600 694.950 ;
        RECT 748.950 691.950 751.050 694.050 ;
        RECT 757.950 691.950 760.050 694.050 ;
        RECT 784.950 691.950 787.050 694.050 ;
        RECT 742.950 685.950 745.050 688.050 ;
        RECT 745.950 679.950 748.050 682.050 ;
        RECT 730.800 658.950 732.900 661.050 ;
        RECT 734.100 659.100 736.200 661.200 ;
        RECT 733.950 655.800 736.050 657.900 ;
        RECT 724.950 651.600 727.050 652.050 ;
        RECT 719.400 650.400 727.050 651.600 ;
        RECT 724.950 649.950 727.050 650.400 ;
        RECT 734.400 643.050 735.600 655.800 ;
        RECT 746.400 652.050 747.600 679.950 ;
        RECT 749.400 654.600 750.600 691.950 ;
        RECT 758.400 688.050 759.600 691.950 ;
        RECT 785.400 688.050 786.600 691.950 ;
        RECT 757.950 685.950 760.050 688.050 ;
        RECT 762.000 687.600 766.050 688.050 ;
        RECT 761.400 685.950 766.050 687.600 ;
        RECT 761.400 681.600 762.600 685.950 ;
        RECT 778.950 684.600 781.050 688.050 ;
        RECT 784.950 685.950 787.050 688.050 ;
        RECT 788.400 684.600 789.600 706.950 ;
        RECT 794.400 694.050 795.600 727.950 ;
        RECT 796.950 720.600 801.000 721.050 ;
        RECT 796.950 718.950 801.600 720.600 ;
        RECT 796.950 706.950 799.050 709.050 ;
        RECT 793.950 691.950 796.050 694.050 ;
        RECT 778.950 684.000 789.600 684.600 ;
        RECT 779.400 683.400 789.600 684.000 ;
        RECT 758.400 680.400 762.600 681.600 ;
        RECT 754.950 676.950 757.050 679.050 ;
        RECT 755.400 670.050 756.600 676.950 ;
        RECT 754.950 667.950 757.050 670.050 ;
        RECT 749.400 653.400 753.600 654.600 ;
        RECT 742.950 649.950 745.050 652.050 ;
        RECT 746.400 649.950 751.050 652.050 ;
        RECT 726.000 642.600 730.050 643.050 ;
        RECT 725.400 642.000 730.050 642.600 ;
        RECT 724.950 640.950 730.050 642.000 ;
        RECT 733.950 640.950 736.050 643.050 ;
        RECT 724.950 637.950 727.050 640.950 ;
        RECT 725.400 625.050 726.600 637.950 ;
        RECT 743.400 634.050 744.600 649.950 ;
        RECT 746.400 646.050 747.600 649.950 ;
        RECT 745.950 643.950 748.050 646.050 ;
        RECT 752.400 643.050 753.600 653.400 ;
        RECT 758.400 643.050 759.600 680.400 ;
        RECT 766.950 676.950 769.050 679.050 ;
        RECT 781.950 676.950 784.050 679.050 ;
        RECT 760.950 673.950 763.050 676.050 ;
        RECT 761.400 664.050 762.600 673.950 ;
        RECT 767.400 670.050 768.600 676.950 ;
        RECT 782.400 673.050 783.600 676.950 ;
        RECT 781.950 670.950 784.050 673.050 ;
        RECT 787.950 670.950 790.050 673.050 ;
        RECT 766.800 667.950 768.900 670.050 ;
        RECT 772.800 667.950 774.900 670.050 ;
        RECT 760.950 661.950 763.050 664.050 ;
        RECT 763.950 655.950 766.050 658.050 ;
        RECT 764.400 652.050 765.600 655.950 ;
        RECT 763.950 649.950 766.050 652.050 ;
        RECT 751.950 640.950 754.050 643.050 ;
        RECT 757.950 640.950 760.050 643.050 ;
        RECT 745.950 637.950 748.050 640.050 ;
        RECT 742.950 631.950 745.050 634.050 ;
        RECT 739.950 628.950 742.050 631.050 ;
        RECT 733.950 625.950 736.050 628.050 ;
        RECT 724.950 622.950 727.050 625.050 ;
        RECT 715.950 616.950 718.050 619.050 ;
        RECT 710.400 608.400 715.050 610.050 ;
        RECT 711.000 607.950 715.050 608.400 ;
        RECT 718.950 607.950 721.050 610.050 ;
        RECT 697.950 598.950 700.050 601.050 ;
        RECT 707.400 598.950 712.050 601.050 ;
        RECT 698.400 595.050 699.600 598.950 ;
        RECT 707.400 595.050 708.600 598.950 ;
        RECT 715.950 595.950 718.050 598.050 ;
        RECT 697.950 592.950 700.050 595.050 ;
        RECT 706.950 592.950 709.050 595.050 ;
        RECT 688.950 588.600 691.050 589.050 ;
        RECT 686.400 587.400 691.050 588.600 ;
        RECT 679.950 571.950 682.050 574.050 ;
        RECT 673.950 553.950 676.050 556.050 ;
        RECT 680.400 544.050 681.600 571.950 ;
        RECT 686.400 565.050 687.600 587.400 ;
        RECT 688.950 586.950 691.050 587.400 ;
        RECT 691.950 580.950 694.050 583.050 ;
        RECT 716.400 582.600 717.600 595.950 ;
        RECT 719.400 586.050 720.600 607.950 ;
        RECT 725.400 589.050 726.600 622.950 ;
        RECT 734.400 610.050 735.600 625.950 ;
        RECT 740.400 610.050 741.600 628.950 ;
        RECT 733.950 607.950 736.050 610.050 ;
        RECT 739.950 607.950 742.050 610.050 ;
        RECT 736.950 595.950 739.050 598.050 ;
        RECT 724.950 586.950 727.050 589.050 ;
        RECT 718.950 583.950 721.050 586.050 ;
        RECT 713.400 582.000 717.600 582.600 ;
        RECT 712.950 581.400 717.600 582.000 ;
        RECT 692.400 574.050 693.600 580.950 ;
        RECT 712.950 580.050 715.050 581.400 ;
        RECT 737.400 580.050 738.600 595.950 ;
        RECT 742.950 589.950 745.050 592.050 ;
        RECT 712.800 579.000 715.050 580.050 ;
        RECT 712.800 577.950 714.900 579.000 ;
        RECT 716.100 577.950 718.200 580.050 ;
        RECT 736.950 577.950 739.050 580.050 ;
        RECT 688.950 572.400 693.600 574.050 ;
        RECT 688.950 571.950 693.000 572.400 ;
        RECT 697.950 571.950 700.050 574.050 ;
        RECT 712.950 573.600 715.050 574.050 ;
        RECT 707.400 572.400 715.050 573.600 ;
        RECT 685.950 562.950 688.050 565.050 ;
        RECT 691.950 562.950 694.050 565.050 ;
        RECT 692.400 556.050 693.600 562.950 ;
        RECT 691.950 553.950 694.050 556.050 ;
        RECT 679.950 541.950 682.050 544.050 ;
        RECT 676.950 538.950 679.050 541.050 ;
        RECT 677.400 532.050 678.600 538.950 ;
        RECT 682.950 535.950 685.050 538.050 ;
        RECT 683.400 532.050 684.600 535.950 ;
        RECT 698.400 532.050 699.600 571.950 ;
        RECT 707.400 556.050 708.600 572.400 ;
        RECT 712.950 571.950 715.050 572.400 ;
        RECT 716.400 565.050 717.600 577.950 ;
        RECT 721.950 574.950 724.050 577.050 ;
        RECT 709.950 562.950 712.050 565.050 ;
        RECT 715.950 562.950 718.050 565.050 ;
        RECT 710.400 559.050 711.600 562.950 ;
        RECT 709.950 556.950 712.050 559.050 ;
        RECT 722.400 556.050 723.600 574.950 ;
        RECT 727.950 574.050 730.050 577.050 ;
        RECT 727.950 573.000 733.050 574.050 ;
        RECT 728.400 572.400 733.050 573.000 ;
        RECT 729.000 571.950 733.050 572.400 ;
        RECT 737.400 565.050 738.600 577.950 ;
        RECT 739.950 571.950 742.050 574.050 ;
        RECT 727.950 562.950 730.050 565.050 ;
        RECT 733.950 563.400 738.600 565.050 ;
        RECT 733.950 562.950 738.000 563.400 ;
        RECT 728.400 559.050 729.600 562.950 ;
        RECT 727.950 556.950 730.050 559.050 ;
        RECT 706.950 553.950 709.050 556.050 ;
        RECT 721.950 553.950 724.050 556.050 ;
        RECT 724.950 541.950 727.050 544.050 ;
        RECT 709.950 538.950 712.050 541.050 ;
        RECT 703.950 535.950 706.050 538.050 ;
        RECT 704.400 532.050 705.600 535.950 ;
        RECT 670.950 529.950 673.050 532.050 ;
        RECT 676.950 529.950 679.050 532.050 ;
        RECT 682.950 529.950 685.050 532.050 ;
        RECT 697.950 529.950 700.050 532.050 ;
        RECT 703.950 529.950 706.050 532.050 ;
        RECT 671.400 525.600 672.600 529.950 ;
        RECT 671.400 524.400 684.600 525.600 ;
        RECT 670.950 520.950 673.050 523.050 ;
        RECT 679.950 520.950 682.050 523.050 ;
        RECT 683.400 522.600 684.600 524.400 ;
        RECT 710.400 523.050 711.600 538.950 ;
        RECT 725.400 532.050 726.600 541.950 ;
        RECT 740.400 535.050 741.600 571.950 ;
        RECT 743.400 550.050 744.600 589.950 ;
        RECT 742.950 547.950 745.050 550.050 ;
        RECT 746.400 538.200 747.600 637.950 ;
        RECT 748.950 634.950 751.050 637.050 ;
        RECT 749.400 577.050 750.600 634.950 ;
        RECT 754.950 607.950 757.050 610.050 ;
        RECT 755.400 595.050 756.600 607.950 ;
        RECT 758.400 601.050 759.600 640.950 ;
        RECT 767.400 619.050 768.600 667.950 ;
        RECT 773.400 658.200 774.600 667.950 ;
        RECT 772.950 656.100 775.050 658.200 ;
        RECT 784.950 649.950 787.050 652.050 ;
        RECT 772.950 646.950 775.050 649.050 ;
        RECT 773.400 643.050 774.600 646.950 ;
        RECT 773.400 641.400 778.050 643.050 ;
        RECT 774.000 640.950 778.050 641.400 ;
        RECT 781.950 640.950 784.050 643.050 ;
        RECT 769.950 634.950 772.050 637.050 ;
        RECT 770.400 622.050 771.600 634.950 ;
        RECT 782.400 628.050 783.600 640.950 ;
        RECT 785.400 640.050 786.600 649.950 ;
        RECT 784.950 637.950 787.050 640.050 ;
        RECT 781.950 625.950 784.050 628.050 ;
        RECT 769.950 619.950 772.050 622.050 ;
        RECT 766.950 616.950 769.050 619.050 ;
        RECT 772.950 616.950 775.050 619.050 ;
        RECT 766.950 610.950 769.050 613.050 ;
        RECT 757.950 598.950 760.050 601.050 ;
        RECT 754.950 592.950 757.050 595.050 ;
        RECT 757.950 586.950 760.050 589.050 ;
        RECT 758.400 577.050 759.600 586.950 ;
        RECT 749.400 575.400 754.050 577.050 ;
        RECT 750.000 574.950 754.050 575.400 ;
        RECT 757.950 574.950 760.050 577.050 ;
        RECT 767.400 565.050 768.600 610.950 ;
        RECT 773.400 601.050 774.600 616.950 ;
        RECT 788.400 610.050 789.600 670.950 ;
        RECT 797.400 664.050 798.600 706.950 ;
        RECT 800.400 706.050 801.600 718.950 ;
        RECT 799.950 703.950 802.050 706.050 ;
        RECT 803.400 688.050 804.600 733.950 ;
        RECT 809.400 729.600 810.600 739.950 ;
        RECT 812.400 736.050 813.600 754.950 ;
        RECT 814.950 745.950 817.050 748.050 ;
        RECT 820.950 745.950 823.050 748.050 ;
        RECT 815.400 739.050 816.600 745.950 ;
        RECT 814.950 736.950 817.050 739.050 ;
        RECT 811.950 733.950 814.050 736.050 ;
        RECT 814.950 729.600 817.050 730.050 ;
        RECT 809.400 728.400 817.050 729.600 ;
        RECT 814.950 727.950 817.050 728.400 ;
        RECT 821.400 721.050 822.600 745.950 ;
        RECT 817.950 719.400 822.600 721.050 ;
        RECT 817.950 718.950 822.000 719.400 ;
        RECT 814.950 703.950 817.050 706.050 ;
        RECT 811.950 700.950 814.050 703.050 ;
        RECT 802.950 685.950 805.050 688.050 ;
        RECT 790.950 661.950 793.050 664.050 ;
        RECT 796.950 661.950 799.050 664.050 ;
        RECT 778.950 607.950 781.050 610.050 ;
        RECT 784.950 608.400 789.600 610.050 ;
        RECT 784.950 607.950 789.000 608.400 ;
        RECT 769.950 598.950 772.050 601.050 ;
        RECT 773.400 599.400 778.050 601.050 ;
        RECT 774.000 598.950 778.050 599.400 ;
        RECT 770.400 595.050 771.600 598.950 ;
        RECT 779.400 595.050 780.600 607.950 ;
        RECT 791.400 604.050 792.600 661.950 ;
        RECT 796.950 655.950 799.050 658.050 ;
        RECT 797.400 643.050 798.600 655.950 ;
        RECT 793.950 640.950 796.050 643.050 ;
        RECT 796.950 640.950 799.050 643.050 ;
        RECT 790.950 601.950 793.050 604.050 ;
        RECT 794.400 598.050 795.600 640.950 ;
        RECT 808.950 634.800 811.050 636.900 ;
        RECT 809.400 616.050 810.600 634.800 ;
        RECT 812.400 622.050 813.600 700.950 ;
        RECT 811.950 619.950 814.050 622.050 ;
        RECT 815.400 619.050 816.600 703.950 ;
        RECT 818.400 658.050 819.600 718.950 ;
        RECT 824.400 717.600 825.600 754.950 ;
        RECT 851.400 748.050 852.600 823.950 ;
        RECT 853.950 820.950 856.050 823.050 ;
        RECT 854.400 769.050 855.600 820.950 ;
        RECT 866.400 820.050 867.600 826.950 ;
        RECT 865.950 817.950 868.050 820.050 ;
        RECT 856.800 814.950 858.900 817.050 ;
        RECT 853.950 766.950 856.050 769.050 ;
        RECT 854.400 757.050 855.600 766.950 ;
        RECT 857.400 766.050 858.600 814.950 ;
        RECT 866.400 811.050 867.600 817.950 ;
        RECT 872.400 811.050 873.600 847.950 ;
        RECT 876.000 843.600 880.050 844.050 ;
        RECT 875.400 841.950 880.050 843.600 ;
        RECT 883.950 841.950 886.050 844.050 ;
        RECT 875.400 838.200 876.600 841.950 ;
        RECT 874.950 836.100 877.050 838.200 ;
        RECT 874.950 832.800 877.050 834.900 ;
        RECT 875.400 817.050 876.600 832.800 ;
        RECT 884.400 829.050 885.600 841.950 ;
        RECT 883.950 826.950 886.050 829.050 ;
        RECT 890.400 817.050 891.600 881.400 ;
        RECT 910.950 877.950 913.050 880.050 ;
        RECT 895.950 868.950 898.050 871.050 ;
        RECT 892.950 832.950 895.050 835.050 ;
        RECT 893.400 820.050 894.600 832.950 ;
        RECT 892.950 817.950 895.050 820.050 ;
        RECT 874.950 814.950 877.050 817.050 ;
        RECT 889.950 814.950 892.050 817.050 ;
        RECT 886.950 811.950 889.050 814.050 ;
        RECT 865.950 808.950 868.050 811.050 ;
        RECT 871.950 808.950 874.050 811.050 ;
        RECT 887.400 808.050 888.600 811.950 ;
        RECT 859.950 805.950 862.050 808.050 ;
        RECT 886.950 805.950 889.050 808.050 ;
        RECT 856.950 763.950 859.050 766.050 ;
        RECT 853.950 754.950 856.050 757.050 ;
        RECT 850.950 745.950 853.050 748.050 ;
        RECT 847.950 742.950 850.050 745.050 ;
        RECT 826.950 733.950 829.050 736.050 ;
        RECT 827.400 730.050 828.600 733.950 ;
        RECT 827.400 728.400 832.050 730.050 ;
        RECT 828.000 727.950 832.050 728.400 ;
        RECT 835.950 727.950 838.050 730.050 ;
        RECT 829.950 718.950 832.050 721.050 ;
        RECT 821.400 716.400 825.600 717.600 ;
        RECT 821.400 706.050 822.600 716.400 ;
        RECT 826.950 712.950 829.050 715.050 ;
        RECT 820.950 703.950 823.050 706.050 ;
        RECT 823.950 700.950 826.050 703.050 ;
        RECT 824.400 688.050 825.600 700.950 ;
        RECT 823.950 685.950 826.050 688.050 ;
        RECT 820.950 676.950 823.050 679.050 ;
        RECT 821.400 670.050 822.600 676.950 ;
        RECT 820.950 667.950 823.050 670.050 ;
        RECT 824.400 667.050 825.600 685.950 ;
        RECT 827.400 679.050 828.600 712.950 ;
        RECT 830.400 688.050 831.600 718.950 ;
        RECT 836.400 712.050 837.600 727.950 ;
        RECT 844.950 718.950 847.050 721.050 ;
        RECT 845.400 712.050 846.600 718.950 ;
        RECT 835.950 709.950 838.050 712.050 ;
        RECT 844.950 709.950 847.050 712.050 ;
        RECT 848.400 708.600 849.600 742.950 ;
        RECT 860.400 736.050 861.600 805.950 ;
        RECT 896.400 802.050 897.600 868.950 ;
        RECT 898.950 847.950 901.050 850.050 ;
        RECT 899.400 844.050 900.600 847.950 ;
        RECT 898.950 841.950 901.050 844.050 ;
        RECT 904.950 840.600 907.050 844.050 ;
        RECT 902.400 840.000 907.050 840.600 ;
        RECT 902.400 839.400 906.600 840.000 ;
        RECT 902.400 829.050 903.600 839.400 ;
        RECT 911.400 832.050 912.600 877.950 ;
        RECT 910.950 829.950 913.050 832.050 ;
        RECT 901.950 826.950 904.050 829.050 ;
        RECT 910.950 823.950 913.050 826.050 ;
        RECT 898.950 817.950 901.050 820.050 ;
        RECT 899.400 814.050 900.600 817.950 ;
        RECT 898.950 811.950 901.050 814.050 ;
        RECT 895.950 799.950 898.050 802.050 ;
        RECT 904.950 799.950 907.050 802.050 ;
        RECT 868.950 796.950 871.050 799.050 ;
        RECT 883.950 796.950 886.050 799.050 ;
        RECT 889.950 796.950 892.050 799.050 ;
        RECT 869.400 793.050 870.600 796.950 ;
        RECT 868.950 790.950 871.050 793.050 ;
        RECT 884.400 784.050 885.600 796.950 ;
        RECT 890.400 793.050 891.600 796.950 ;
        RECT 889.800 790.950 891.900 793.050 ;
        RECT 893.100 790.950 895.200 793.050 ;
        RECT 889.950 784.950 892.050 787.050 ;
        RECT 883.950 781.950 886.050 784.050 ;
        RECT 886.950 766.950 889.050 769.050 ;
        RECT 862.950 762.600 865.050 766.050 ;
        RECT 862.950 762.000 870.600 762.600 ;
        RECT 863.400 761.400 870.600 762.000 ;
        RECT 865.950 754.950 868.050 757.050 ;
        RECT 850.950 733.950 853.050 736.050 ;
        RECT 859.950 733.950 862.050 736.050 ;
        RECT 845.400 707.400 849.600 708.600 ;
        RECT 841.950 703.950 844.050 706.050 ;
        RECT 829.950 685.950 832.050 688.050 ;
        RECT 826.950 676.950 829.050 679.050 ;
        RECT 827.400 673.050 828.600 676.950 ;
        RECT 826.950 670.950 829.050 673.050 ;
        RECT 832.950 667.950 835.050 670.050 ;
        RECT 823.950 664.950 826.050 667.050 ;
        RECT 817.950 655.950 820.050 658.050 ;
        RECT 823.950 655.950 826.050 658.050 ;
        RECT 817.950 649.950 820.050 652.050 ;
        RECT 818.400 625.050 819.600 649.950 ;
        RECT 824.400 643.050 825.600 655.950 ;
        RECT 824.400 640.950 829.050 643.050 ;
        RECT 824.400 634.050 825.600 640.950 ;
        RECT 823.950 631.950 826.050 634.050 ;
        RECT 817.950 622.950 820.050 625.050 ;
        RECT 826.950 622.950 829.050 625.050 ;
        RECT 814.950 616.950 817.050 619.050 ;
        RECT 808.950 613.950 811.050 616.050 ;
        RECT 799.950 610.050 802.050 613.050 ;
        RECT 827.400 610.050 828.600 622.950 ;
        RECT 833.400 612.600 834.600 667.950 ;
        RECT 842.400 667.050 843.600 703.950 ;
        RECT 845.400 684.600 846.600 707.400 ;
        RECT 851.400 688.050 852.600 733.950 ;
        RECT 862.950 697.950 865.050 700.050 ;
        RECT 859.950 688.050 862.050 691.050 ;
        RECT 850.950 685.950 853.050 688.050 ;
        RECT 856.950 687.000 862.050 688.050 ;
        RECT 856.950 686.400 861.600 687.000 ;
        RECT 856.950 685.950 861.000 686.400 ;
        RECT 845.400 683.400 849.600 684.600 ;
        RECT 848.400 669.600 849.600 683.400 ;
        RECT 851.400 673.050 852.600 685.950 ;
        RECT 863.400 679.050 864.600 697.950 ;
        RECT 859.950 677.400 864.600 679.050 ;
        RECT 859.950 676.950 864.000 677.400 ;
        RECT 853.950 673.950 856.050 676.050 ;
        RECT 850.950 670.950 853.050 673.050 ;
        RECT 848.400 668.400 852.600 669.600 ;
        RECT 838.800 664.950 840.900 667.050 ;
        RECT 842.100 664.950 844.200 667.050 ;
        RECT 835.950 658.950 838.050 661.050 ;
        RECT 836.400 643.050 837.600 658.950 ;
        RECT 839.400 652.050 840.600 664.950 ;
        RECT 839.400 650.400 844.050 652.050 ;
        RECT 840.000 649.950 844.050 650.400 ;
        RECT 836.400 641.400 841.050 643.050 ;
        RECT 837.000 640.950 841.050 641.400 ;
        RECT 847.950 640.950 850.050 643.050 ;
        RECT 838.950 634.950 841.050 637.050 ;
        RECT 835.950 622.950 838.050 625.050 ;
        RECT 830.400 611.400 834.600 612.600 ;
        RECT 799.950 609.000 805.050 610.050 ;
        RECT 800.400 608.400 805.050 609.000 ;
        RECT 801.000 607.950 805.050 608.400 ;
        RECT 808.950 606.600 811.050 610.050 ;
        RECT 814.950 606.600 817.050 610.050 ;
        RECT 826.950 607.950 829.050 610.050 ;
        RECT 808.950 606.000 817.050 606.600 ;
        RECT 809.400 605.400 816.600 606.000 ;
        RECT 799.950 598.950 802.050 601.050 ;
        RECT 808.950 598.950 811.050 601.050 ;
        RECT 823.950 598.950 826.050 601.050 ;
        RECT 769.950 592.950 772.050 595.050 ;
        RECT 778.950 592.950 781.050 595.050 ;
        RECT 787.950 594.600 790.050 598.050 ;
        RECT 793.950 595.950 796.050 598.050 ;
        RECT 800.400 595.050 801.600 598.950 ;
        RECT 785.400 594.000 790.050 594.600 ;
        RECT 785.400 593.400 789.600 594.000 ;
        RECT 779.400 580.050 780.600 592.950 ;
        RECT 785.400 592.050 786.600 593.400 ;
        RECT 799.950 592.950 802.050 595.050 ;
        RECT 781.950 590.400 786.600 592.050 ;
        RECT 781.950 589.950 786.000 590.400 ;
        RECT 787.950 589.950 790.050 592.050 ;
        RECT 784.950 586.950 787.050 589.050 ;
        RECT 772.950 577.950 775.050 580.050 ;
        RECT 778.800 577.950 780.900 580.050 ;
        RECT 773.400 574.050 774.600 577.950 ;
        RECT 772.950 571.950 775.050 574.050 ;
        RECT 778.950 571.950 781.050 574.050 ;
        RECT 760.950 562.950 763.050 565.050 ;
        RECT 766.950 562.950 769.050 565.050 ;
        RECT 754.950 550.950 757.050 553.050 ;
        RECT 745.950 536.100 748.050 538.200 ;
        RECT 739.950 532.950 742.050 535.050 ;
        RECT 745.950 532.800 748.050 534.900 ;
        RECT 718.950 529.950 721.050 532.050 ;
        RECT 724.950 529.950 727.050 532.050 ;
        RECT 730.950 529.950 733.050 532.050 ;
        RECT 694.950 522.600 697.050 523.050 ;
        RECT 683.400 521.400 697.050 522.600 ;
        RECT 694.950 520.950 697.050 521.400 ;
        RECT 709.950 520.950 712.050 523.050 ;
        RECT 664.950 511.950 667.050 514.050 ;
        RECT 607.950 502.950 610.050 505.050 ;
        RECT 646.950 502.950 649.050 505.050 ;
        RECT 652.950 502.950 655.050 505.050 ;
        RECT 658.950 502.950 661.050 505.050 ;
        RECT 599.400 498.000 603.600 498.600 ;
        RECT 599.400 497.400 604.050 498.000 ;
        RECT 580.950 495.600 583.050 496.050 ;
        RECT 586.950 495.600 589.050 496.050 ;
        RECT 580.950 494.400 589.050 495.600 ;
        RECT 580.950 493.950 583.050 494.400 ;
        RECT 586.950 493.950 589.050 494.400 ;
        RECT 595.950 493.950 598.050 496.050 ;
        RECT 601.950 493.950 604.050 497.400 ;
        RECT 596.400 487.050 597.600 493.950 ;
        RECT 608.400 487.050 609.600 502.950 ;
        RECT 625.950 499.950 628.050 502.050 ;
        RECT 626.400 487.050 627.600 499.950 ;
        RECT 653.400 499.050 654.600 502.950 ;
        RECT 640.950 495.600 643.050 496.050 ;
        RECT 646.950 495.600 649.050 499.050 ;
        RECT 652.950 496.950 655.050 499.050 ;
        RECT 659.400 496.050 660.600 502.950 ;
        RECT 638.400 495.000 649.050 495.600 ;
        RECT 638.400 494.400 648.600 495.000 ;
        RECT 553.950 484.950 556.050 487.050 ;
        RECT 559.950 484.950 562.050 487.050 ;
        RECT 565.950 484.950 568.050 487.050 ;
        RECT 596.400 485.400 601.050 487.050 ;
        RECT 597.000 484.950 601.050 485.400 ;
        RECT 604.950 485.400 609.600 487.050 ;
        RECT 604.950 484.950 609.000 485.400 ;
        RECT 625.950 484.950 628.050 487.050 ;
        RECT 631.950 484.950 634.050 487.050 ;
        RECT 560.400 481.050 561.600 484.950 ;
        RECT 520.950 478.950 523.050 481.050 ;
        RECT 544.950 478.950 547.050 481.050 ;
        RECT 559.950 478.950 562.050 481.050 ;
        RECT 626.400 472.050 627.600 484.950 ;
        RECT 632.400 481.050 633.600 484.950 ;
        RECT 631.950 478.950 634.050 481.050 ;
        RECT 625.950 469.950 628.050 472.050 ;
        RECT 634.950 466.950 637.050 469.050 ;
        RECT 592.950 463.950 595.050 466.050 ;
        RECT 523.950 460.950 526.050 463.050 ;
        RECT 550.950 460.950 553.050 463.050 ;
        RECT 571.950 460.950 574.050 463.050 ;
        RECT 508.950 457.950 511.050 460.050 ;
        RECT 509.400 454.050 510.600 457.950 ;
        RECT 524.400 454.050 525.600 460.950 ;
        RECT 551.400 454.050 552.600 460.950 ;
        RECT 572.400 454.050 573.600 460.950 ;
        RECT 577.950 457.950 580.050 460.050 ;
        RECT 589.950 457.950 592.050 460.050 ;
        RECT 578.400 454.050 579.600 457.950 ;
        RECT 463.950 451.950 466.050 454.050 ;
        RECT 469.950 451.950 472.050 454.050 ;
        RECT 481.950 451.950 484.050 454.050 ;
        RECT 485.400 452.400 490.050 454.050 ;
        RECT 486.000 451.950 490.050 452.400 ;
        RECT 496.950 453.600 499.050 454.050 ;
        RECT 502.950 453.600 505.050 454.050 ;
        RECT 496.950 452.400 505.050 453.600 ;
        RECT 496.950 451.950 499.050 452.400 ;
        RECT 502.950 451.950 505.050 452.400 ;
        RECT 508.950 451.950 511.050 454.050 ;
        RECT 523.950 451.950 526.050 454.050 ;
        RECT 529.950 451.950 532.050 454.050 ;
        RECT 550.950 451.950 553.050 454.050 ;
        RECT 556.950 453.600 561.000 454.050 ;
        RECT 556.950 451.950 561.600 453.600 ;
        RECT 571.950 451.950 574.050 454.050 ;
        RECT 577.950 451.950 580.050 454.050 ;
        RECT 439.950 442.950 442.050 445.050 ;
        RECT 457.950 442.950 460.050 445.050 ;
        RECT 479.100 442.950 481.200 445.050 ;
        RECT 496.950 442.950 499.050 445.050 ;
        RECT 520.950 444.600 523.050 445.050 ;
        RECT 526.950 444.600 529.050 445.050 ;
        RECT 520.950 443.400 529.050 444.600 ;
        RECT 520.950 442.950 523.050 443.400 ;
        RECT 526.950 442.950 529.050 443.400 ;
        RECT 440.400 439.050 441.600 442.950 ;
        RECT 427.800 436.950 429.900 439.050 ;
        RECT 439.950 436.950 442.050 439.050 ;
        RECT 428.400 430.050 429.600 436.950 ;
        RECT 427.950 427.950 430.050 430.050 ;
        RECT 479.400 427.050 480.600 442.950 ;
        RECT 487.950 427.950 490.050 430.050 ;
        RECT 478.950 424.950 481.050 427.050 ;
        RECT 484.950 424.950 487.050 427.050 ;
        RECT 460.950 421.950 463.050 424.050 ;
        RECT 416.400 416.400 421.050 418.050 ;
        RECT 417.000 415.950 421.050 416.400 ;
        RECT 433.950 415.950 436.050 418.050 ;
        RECT 442.950 415.950 445.050 418.050 ;
        RECT 415.950 408.600 418.050 412.050 ;
        RECT 421.950 408.600 424.050 409.050 ;
        RECT 415.950 408.000 424.050 408.600 ;
        RECT 416.400 407.400 424.050 408.000 ;
        RECT 421.950 406.950 424.050 407.400 ;
        RECT 427.950 406.950 430.050 409.050 ;
        RECT 428.400 403.050 429.600 406.950 ;
        RECT 427.950 400.950 430.050 403.050 ;
        RECT 412.950 394.950 415.050 397.050 ;
        RECT 412.950 388.950 415.050 391.050 ;
        RECT 413.400 355.050 414.600 388.950 ;
        RECT 434.400 388.050 435.600 415.950 ;
        RECT 443.400 397.050 444.600 415.950 ;
        RECT 454.950 409.950 457.050 412.050 ;
        RECT 448.950 403.950 451.050 406.050 ;
        RECT 442.950 394.950 445.050 397.050 ;
        RECT 433.950 385.950 436.050 388.050 ;
        RECT 449.400 376.050 450.600 403.950 ;
        RECT 455.400 391.050 456.600 409.950 ;
        RECT 454.950 388.950 457.050 391.050 ;
        RECT 461.400 382.050 462.600 421.950 ;
        RECT 485.400 418.050 486.600 424.950 ;
        RECT 472.950 415.950 475.050 418.050 ;
        RECT 484.950 415.950 487.050 418.050 ;
        RECT 473.400 400.050 474.600 415.950 ;
        RECT 488.400 409.050 489.600 427.950 ;
        RECT 497.400 409.050 498.600 442.950 ;
        RECT 520.950 436.950 523.050 439.050 ;
        RECT 514.950 421.950 517.050 424.050 ;
        RECT 515.400 409.050 516.600 421.950 ;
        RECT 521.400 418.050 522.600 436.950 ;
        RECT 530.400 427.050 531.600 451.950 ;
        RECT 560.400 445.050 561.600 451.950 ;
        RECT 547.950 442.950 550.050 445.050 ;
        RECT 559.950 442.950 562.050 445.050 ;
        RECT 568.950 444.600 571.050 445.050 ;
        RECT 568.950 443.400 579.600 444.600 ;
        RECT 568.950 442.950 571.050 443.400 ;
        RECT 548.400 436.050 549.600 442.950 ;
        RECT 578.400 439.050 579.600 443.400 ;
        RECT 562.950 436.950 565.050 439.050 ;
        RECT 577.950 436.950 580.050 439.050 ;
        RECT 547.950 433.950 550.050 436.050 ;
        RECT 529.950 424.950 532.050 427.050 ;
        RECT 517.950 416.400 522.600 418.050 ;
        RECT 517.950 415.950 522.000 416.400 ;
        RECT 526.950 415.950 529.050 418.050 ;
        RECT 541.950 417.600 544.050 418.050 ;
        RECT 547.950 417.600 550.050 418.050 ;
        RECT 541.950 416.400 550.050 417.600 ;
        RECT 541.950 415.950 544.050 416.400 ;
        RECT 547.950 415.950 550.050 416.400 ;
        RECT 487.950 406.950 490.050 409.050 ;
        RECT 493.950 407.400 498.600 409.050 ;
        RECT 493.950 406.950 498.000 407.400 ;
        RECT 514.950 406.950 517.050 409.050 ;
        RECT 520.950 406.950 523.050 409.050 ;
        RECT 521.400 403.050 522.600 406.950 ;
        RECT 508.950 400.950 511.050 403.050 ;
        RECT 520.950 400.950 523.050 403.050 ;
        RECT 472.950 397.950 475.050 400.050 ;
        RECT 473.400 394.050 474.600 397.950 ;
        RECT 466.950 391.950 469.050 394.050 ;
        RECT 472.950 391.950 475.050 394.050 ;
        RECT 454.950 379.950 457.050 382.050 ;
        RECT 460.950 379.950 463.050 382.050 ;
        RECT 455.400 376.050 456.600 379.950 ;
        RECT 448.950 373.950 451.050 376.050 ;
        RECT 454.950 373.950 457.050 376.050 ;
        RECT 421.950 370.950 424.050 373.050 ;
        RECT 430.950 370.950 433.050 373.050 ;
        RECT 412.950 352.950 415.050 355.050 ;
        RECT 413.400 349.050 414.600 352.950 ;
        RECT 412.950 346.950 415.050 349.050 ;
        RECT 413.400 343.050 414.600 346.950 ;
        RECT 412.950 340.950 415.050 343.050 ;
        RECT 422.400 340.050 423.600 370.950 ;
        RECT 424.950 352.950 427.050 355.050 ;
        RECT 425.400 346.050 426.600 352.950 ;
        RECT 431.400 352.050 432.600 370.950 ;
        RECT 445.950 364.950 448.050 367.050 ;
        RECT 446.400 357.600 447.600 364.950 ;
        RECT 451.950 361.950 454.050 364.050 ;
        RECT 446.400 356.400 450.600 357.600 ;
        RECT 430.950 349.950 433.050 352.050 ;
        RECT 442.950 349.950 445.050 352.050 ;
        RECT 436.950 346.950 439.050 349.050 ;
        RECT 424.950 343.950 427.050 346.050 ;
        RECT 433.950 343.950 436.050 346.050 ;
        RECT 434.400 340.050 435.600 343.950 ;
        RECT 421.950 337.950 424.050 340.050 ;
        RECT 433.950 337.950 436.050 340.050 ;
        RECT 421.950 330.600 424.050 334.050 ;
        RECT 437.400 331.050 438.600 346.950 ;
        RECT 443.400 334.050 444.600 349.950 ;
        RECT 442.950 331.950 445.050 334.050 ;
        RECT 430.950 330.600 433.050 331.050 ;
        RECT 421.950 330.000 433.050 330.600 ;
        RECT 422.400 329.400 433.050 330.000 ;
        RECT 430.950 328.950 433.050 329.400 ;
        RECT 436.950 328.950 439.050 331.050 ;
        RECT 443.400 310.050 444.600 331.950 ;
        RECT 442.950 307.950 445.050 310.050 ;
        RECT 443.400 295.050 444.600 307.950 ;
        RECT 449.400 298.050 450.600 356.400 ;
        RECT 452.400 334.050 453.600 361.950 ;
        RECT 460.950 349.950 463.050 352.050 ;
        RECT 451.950 331.950 454.050 334.050 ;
        RECT 448.950 295.950 451.050 298.050 ;
        RECT 432.000 294.600 436.050 295.050 ;
        RECT 431.400 292.950 436.050 294.600 ;
        RECT 442.950 292.950 445.050 295.050 ;
        RECT 415.950 286.950 418.050 289.050 ;
        RECT 416.400 277.050 417.600 286.950 ;
        RECT 415.950 274.950 418.050 277.050 ;
        RECT 431.400 271.050 432.600 292.950 ;
        RECT 433.950 271.950 436.050 274.050 ;
        RECT 430.950 268.950 433.050 271.050 ;
        RECT 421.950 259.950 424.050 262.050 ;
        RECT 415.950 244.950 418.050 247.050 ;
        RECT 385.950 241.950 388.050 244.050 ;
        RECT 409.950 241.950 412.050 244.050 ;
        RECT 394.950 238.950 397.050 241.050 ;
        RECT 388.950 220.950 391.050 223.050 ;
        RECT 389.400 217.050 390.600 220.950 ;
        RECT 379.950 216.600 382.050 217.050 ;
        RECT 379.950 215.400 387.600 216.600 ;
        RECT 379.950 214.950 382.050 215.400 ;
        RECT 386.400 213.600 387.600 215.400 ;
        RECT 388.950 214.950 391.050 217.050 ;
        RECT 386.400 213.000 393.600 213.600 ;
        RECT 386.400 212.400 394.050 213.000 ;
        RECT 391.950 208.950 394.050 212.400 ;
        RECT 395.400 196.050 396.600 238.950 ;
        RECT 416.400 235.050 417.600 244.950 ;
        RECT 422.400 241.050 423.600 259.950 ;
        RECT 430.950 253.950 433.050 256.050 ;
        RECT 424.950 250.950 427.050 253.050 ;
        RECT 425.400 244.050 426.600 250.950 ;
        RECT 424.950 241.950 427.050 244.050 ;
        RECT 421.950 238.950 424.050 241.050 ;
        RECT 427.950 238.950 430.050 241.050 ;
        RECT 415.950 232.950 418.050 235.050 ;
        RECT 409.950 223.950 412.050 226.050 ;
        RECT 410.400 220.050 411.600 223.950 ;
        RECT 416.400 220.050 417.600 232.950 ;
        RECT 421.950 229.950 424.050 232.050 ;
        RECT 409.950 217.950 412.050 220.050 ;
        RECT 415.950 217.950 418.050 220.050 ;
        RECT 412.950 208.950 415.050 211.050 ;
        RECT 413.400 199.050 414.600 208.950 ;
        RECT 412.950 196.950 415.050 199.050 ;
        RECT 371.400 194.400 375.600 195.600 ;
        RECT 352.950 187.950 355.050 190.050 ;
        RECT 357.000 174.600 361.050 175.050 ;
        RECT 337.950 173.400 345.600 174.600 ;
        RECT 347.400 173.400 351.600 174.600 ;
        RECT 337.950 172.950 340.050 173.400 ;
        RECT 323.100 157.950 325.200 160.050 ;
        RECT 328.950 157.950 331.050 160.050 ;
        RECT 347.400 159.600 348.600 173.400 ;
        RECT 356.400 172.950 361.050 174.600 ;
        RECT 352.950 169.950 355.050 172.050 ;
        RECT 347.400 158.400 351.600 159.600 ;
        RECT 316.800 154.950 318.900 157.050 ;
        RECT 320.100 154.800 322.200 156.900 ;
        RECT 320.400 139.050 321.600 154.800 ;
        RECT 319.950 136.950 322.050 139.050 ;
        RECT 308.400 122.400 312.600 123.600 ;
        RECT 308.400 112.050 309.600 122.400 ;
        RECT 307.950 109.950 310.050 112.050 ;
        RECT 323.400 100.050 324.600 157.950 ;
        RECT 346.950 154.950 349.050 157.050 ;
        RECT 337.950 151.950 340.050 154.050 ;
        RECT 331.950 145.950 334.050 148.050 ;
        RECT 332.400 133.050 333.600 145.950 ;
        RECT 328.950 131.400 333.600 133.050 ;
        RECT 328.950 130.950 333.000 131.400 ;
        RECT 338.400 115.050 339.600 151.950 ;
        RECT 343.950 148.950 346.050 151.050 ;
        RECT 344.400 142.050 345.600 148.950 ;
        RECT 347.400 144.600 348.600 154.950 ;
        RECT 350.400 151.050 351.600 158.400 ;
        RECT 353.400 154.050 354.600 169.950 ;
        RECT 356.400 160.050 357.600 172.950 ;
        RECT 355.950 157.950 358.050 160.050 ;
        RECT 358.950 154.950 361.050 157.050 ;
        RECT 352.950 151.950 355.050 154.050 ;
        RECT 349.950 148.950 352.050 151.050 ;
        RECT 347.400 143.400 351.600 144.600 ;
        RECT 344.400 140.400 349.050 142.050 ;
        RECT 345.000 139.950 349.050 140.400 ;
        RECT 350.400 133.050 351.600 143.400 ;
        RECT 359.400 133.050 360.600 154.950 ;
        RECT 364.950 145.950 367.050 148.050 ;
        RECT 349.950 130.950 352.050 133.050 ;
        RECT 355.950 131.400 360.600 133.050 ;
        RECT 365.400 133.050 366.600 145.950 ;
        RECT 365.400 131.400 370.050 133.050 ;
        RECT 355.950 130.950 360.000 131.400 ;
        RECT 366.000 130.950 370.050 131.400 ;
        RECT 337.950 112.950 340.050 115.050 ;
        RECT 356.400 112.050 357.600 130.950 ;
        RECT 371.400 127.200 372.600 194.400 ;
        RECT 394.950 193.950 397.050 196.050 ;
        RECT 373.950 187.950 376.050 190.050 ;
        RECT 409.950 187.950 412.050 190.050 ;
        RECT 374.400 157.050 375.600 187.950 ;
        RECT 406.950 157.950 409.050 160.050 ;
        RECT 373.950 154.950 376.050 157.050 ;
        RECT 400.950 148.950 403.050 151.050 ;
        RECT 394.950 142.950 397.050 145.050 ;
        RECT 379.950 139.950 382.050 142.050 ;
        RECT 361.950 124.950 364.050 127.050 ;
        RECT 370.950 125.100 373.050 127.200 ;
        RECT 334.950 109.950 337.050 112.050 ;
        RECT 349.950 109.950 352.050 112.050 ;
        RECT 355.950 109.950 358.050 112.050 ;
        RECT 325.950 105.600 330.000 106.050 ;
        RECT 325.950 103.950 330.600 105.600 ;
        RECT 329.400 100.050 330.600 103.950 ;
        RECT 292.950 97.950 295.050 100.050 ;
        RECT 304.950 97.950 307.050 100.050 ;
        RECT 310.950 97.950 313.050 100.050 ;
        RECT 322.950 97.950 325.050 100.050 ;
        RECT 328.950 97.950 331.050 100.050 ;
        RECT 293.400 94.050 294.600 97.950 ;
        RECT 298.950 94.950 301.050 97.050 ;
        RECT 292.950 91.950 295.050 94.050 ;
        RECT 299.400 79.050 300.600 94.950 ;
        RECT 305.400 82.050 306.600 97.950 ;
        RECT 311.400 91.050 312.600 97.950 ;
        RECT 335.400 94.050 336.600 109.950 ;
        RECT 350.400 106.050 351.600 109.950 ;
        RECT 349.950 103.950 352.050 106.050 ;
        RECT 343.950 97.950 346.050 100.050 ;
        RECT 334.950 91.950 337.050 94.050 ;
        RECT 310.950 88.950 313.050 91.050 ;
        RECT 304.950 79.950 307.050 82.050 ;
        RECT 322.950 79.950 325.050 82.050 ;
        RECT 298.950 76.950 301.050 79.050 ;
        RECT 307.950 73.950 310.050 76.050 ;
        RECT 280.950 58.950 283.050 61.050 ;
        RECT 287.400 59.400 292.050 61.050 ;
        RECT 288.000 58.950 292.050 59.400 ;
        RECT 308.400 55.050 309.600 73.950 ;
        RECT 323.400 67.050 324.600 79.950 ;
        RECT 328.950 73.950 331.050 76.050 ;
        RECT 322.950 64.950 325.050 67.050 ;
        RECT 323.400 61.050 324.600 64.950 ;
        RECT 329.400 64.050 330.600 73.950 ;
        RECT 328.950 61.950 331.050 64.050 ;
        RECT 335.400 61.050 336.600 91.950 ;
        RECT 344.400 82.050 345.600 97.950 ;
        RECT 343.950 79.950 346.050 82.050 ;
        RECT 343.950 64.950 346.050 67.050 ;
        RECT 322.950 58.950 325.050 61.050 ;
        RECT 334.950 58.950 337.050 61.050 ;
        RECT 307.950 52.950 310.050 55.050 ;
        RECT 319.950 51.600 322.050 55.050 ;
        RECT 325.950 51.600 328.050 52.050 ;
        RECT 319.950 51.000 328.050 51.600 ;
        RECT 320.400 50.400 328.050 51.000 ;
        RECT 325.950 49.950 328.050 50.400 ;
        RECT 331.950 49.950 334.050 52.050 ;
        RECT 277.950 45.600 280.050 49.050 ;
        RECT 289.950 45.600 292.050 46.050 ;
        RECT 277.950 45.000 292.050 45.600 ;
        RECT 278.400 44.400 292.050 45.000 ;
        RECT 289.950 43.950 292.050 44.400 ;
        RECT 298.950 43.950 301.050 46.050 ;
        RECT 325.950 43.950 328.050 46.050 ;
        RECT 271.950 37.950 274.050 40.050 ;
        RECT 283.950 37.950 286.050 40.050 ;
        RECT 265.950 36.600 268.050 37.050 ;
        RECT 254.400 35.400 268.050 36.600 ;
        RECT 235.950 19.950 238.050 22.050 ;
        RECT 242.400 20.400 247.050 22.050 ;
        RECT 243.000 19.950 247.050 20.400 ;
        RECT 254.400 16.050 255.600 35.400 ;
        RECT 265.950 34.950 268.050 35.400 ;
        RECT 262.950 27.600 267.000 28.050 ;
        RECT 262.950 25.950 267.600 27.600 ;
        RECT 266.400 19.050 267.600 25.950 ;
        RECT 284.400 19.050 285.600 37.950 ;
        RECT 299.400 31.050 300.600 43.950 ;
        RECT 299.400 29.400 304.050 31.050 ;
        RECT 300.000 28.950 304.050 29.400 ;
        RECT 307.950 30.600 310.050 31.050 ;
        RECT 313.950 30.600 316.050 31.050 ;
        RECT 307.950 29.400 316.050 30.600 ;
        RECT 307.950 28.950 310.050 29.400 ;
        RECT 313.950 28.950 316.050 29.400 ;
        RECT 326.400 22.050 327.600 43.950 ;
        RECT 332.400 43.050 333.600 49.950 ;
        RECT 335.400 46.050 336.600 58.950 ;
        RECT 344.400 46.050 345.600 64.950 ;
        RECT 355.950 58.950 358.050 61.050 ;
        RECT 349.950 52.950 352.050 55.050 ;
        RECT 350.400 49.050 351.600 52.950 ;
        RECT 349.950 46.950 352.050 49.050 ;
        RECT 334.950 43.950 337.050 46.050 ;
        RECT 343.950 43.950 346.050 46.050 ;
        RECT 331.950 40.950 334.050 43.050 ;
        RECT 331.950 34.950 334.050 37.050 ;
        RECT 337.950 34.950 340.050 37.050 ;
        RECT 332.400 31.050 333.600 34.950 ;
        RECT 338.400 31.050 339.600 34.950 ;
        RECT 331.950 28.950 334.050 31.050 ;
        RECT 337.950 28.950 340.050 31.050 ;
        RECT 344.400 22.050 345.600 43.950 ;
        RECT 356.400 40.050 357.600 58.950 ;
        RECT 355.950 37.950 358.050 40.050 ;
        RECT 298.950 19.950 301.050 22.050 ;
        RECT 310.950 19.950 313.050 22.050 ;
        RECT 326.400 19.950 331.050 22.050 ;
        RECT 340.950 20.400 345.600 22.050 ;
        RECT 340.950 19.950 345.000 20.400 ;
        RECT 265.950 16.950 268.050 19.050 ;
        RECT 283.950 16.950 286.050 19.050 ;
        RECT 299.400 16.050 300.600 19.950 ;
        RECT 304.950 16.950 307.050 19.050 ;
        RECT 244.950 15.600 247.050 16.050 ;
        RECT 230.400 14.400 247.050 15.600 ;
        RECT 244.950 13.950 247.050 14.400 ;
        RECT 253.950 13.950 256.050 16.050 ;
        RECT 298.950 13.950 301.050 16.050 ;
        RECT 145.950 4.950 148.050 7.050 ;
        RECT 187.950 4.950 190.050 7.050 ;
        RECT 226.950 4.950 229.050 7.050 ;
        RECT 305.400 4.050 306.600 16.950 ;
        RECT 311.400 10.050 312.600 19.950 ;
        RECT 326.400 10.050 327.600 19.950 ;
        RECT 334.950 16.950 337.050 19.050 ;
        RECT 310.950 7.950 313.050 10.050 ;
        RECT 325.950 7.950 328.050 10.050 ;
        RECT 335.400 7.050 336.600 16.950 ;
        RECT 341.400 16.050 342.600 19.950 ;
        RECT 356.400 19.050 357.600 37.950 ;
        RECT 362.400 36.600 363.600 124.950 ;
        RECT 370.950 121.800 373.050 123.900 ;
        RECT 371.400 106.050 372.600 121.800 ;
        RECT 370.950 103.950 373.050 106.050 ;
        RECT 380.400 91.050 381.600 139.950 ;
        RECT 395.400 133.050 396.600 142.950 ;
        RECT 391.950 131.400 396.600 133.050 ;
        RECT 391.950 130.950 396.000 131.400 ;
        RECT 397.950 121.950 400.050 124.050 ;
        RECT 391.950 118.950 394.050 121.050 ;
        RECT 385.950 103.950 388.050 106.050 ;
        RECT 386.400 91.050 387.600 103.950 ;
        RECT 392.400 97.050 393.600 118.950 ;
        RECT 398.400 115.050 399.600 121.950 ;
        RECT 397.950 112.950 400.050 115.050 ;
        RECT 401.400 112.050 402.600 148.950 ;
        RECT 403.950 136.950 406.050 139.050 ;
        RECT 404.400 124.050 405.600 136.950 ;
        RECT 407.400 130.050 408.600 157.950 ;
        RECT 410.400 151.050 411.600 187.950 ;
        RECT 422.400 177.600 423.600 229.950 ;
        RECT 428.400 190.050 429.600 238.950 ;
        RECT 431.400 232.050 432.600 253.950 ;
        RECT 430.950 229.950 433.050 232.050 ;
        RECT 434.400 226.050 435.600 271.950 ;
        RECT 449.400 271.050 450.600 295.950 ;
        RECT 461.400 289.050 462.600 349.950 ;
        RECT 467.400 316.050 468.600 391.950 ;
        RECT 475.950 385.950 478.050 388.050 ;
        RECT 476.400 376.050 477.600 385.950 ;
        RECT 469.950 373.950 472.050 376.050 ;
        RECT 475.950 373.950 478.050 376.050 ;
        RECT 470.400 363.600 471.600 373.950 ;
        RECT 487.950 370.950 490.050 373.050 ;
        RECT 496.950 370.950 499.050 373.050 ;
        RECT 472.950 366.600 477.000 367.050 ;
        RECT 472.950 364.950 477.600 366.600 ;
        RECT 481.950 364.950 484.050 367.050 ;
        RECT 470.400 362.400 474.600 363.600 ;
        RECT 469.950 349.950 472.050 352.050 ;
        RECT 470.400 340.050 471.600 349.950 ;
        RECT 469.950 337.950 472.050 340.050 ;
        RECT 466.950 313.950 469.050 316.050 ;
        RECT 473.400 313.050 474.600 362.400 ;
        RECT 476.400 361.050 477.600 364.950 ;
        RECT 475.950 358.950 478.050 361.050 ;
        RECT 482.400 355.050 483.600 364.950 ;
        RECT 484.950 358.950 487.050 361.050 ;
        RECT 475.950 352.950 478.050 355.050 ;
        RECT 481.950 352.950 484.050 355.050 ;
        RECT 476.400 331.050 477.600 352.950 ;
        RECT 485.400 348.600 486.600 358.950 ;
        RECT 488.400 352.200 489.600 370.950 ;
        RECT 497.400 355.050 498.600 370.950 ;
        RECT 496.950 352.950 499.050 355.050 ;
        RECT 505.950 352.950 508.050 355.050 ;
        RECT 487.950 350.100 490.050 352.200 ;
        RECT 502.950 349.950 505.050 352.050 ;
        RECT 487.950 348.600 490.050 348.900 ;
        RECT 485.400 347.400 490.050 348.600 ;
        RECT 487.950 346.800 490.050 347.400 ;
        RECT 488.400 340.050 489.600 346.800 ;
        RECT 487.950 337.950 490.050 340.050 ;
        RECT 475.950 328.950 478.050 331.050 ;
        RECT 484.950 328.950 487.050 331.050 ;
        RECT 481.950 322.950 484.050 325.050 ;
        RECT 472.950 310.950 475.050 313.050 ;
        RECT 460.950 286.950 463.050 289.050 ;
        RECT 451.950 280.950 454.050 283.050 ;
        RECT 439.950 268.950 442.050 271.050 ;
        RECT 448.950 268.950 451.050 271.050 ;
        RECT 440.400 265.050 441.600 268.950 ;
        RECT 439.950 262.950 442.050 265.050 ;
        RECT 452.400 244.050 453.600 280.950 ;
        RECT 461.400 265.050 462.600 286.950 ;
        RECT 468.000 285.600 472.050 286.050 ;
        RECT 467.400 285.000 472.050 285.600 ;
        RECT 466.950 283.950 472.050 285.000 ;
        RECT 466.950 280.950 469.050 283.950 ;
        RECT 482.400 277.050 483.600 322.950 ;
        RECT 481.950 274.950 484.050 277.050 ;
        RECT 478.950 265.950 481.050 268.050 ;
        RECT 460.950 262.950 463.050 265.050 ;
        RECT 479.400 262.050 480.600 265.950 ;
        RECT 478.950 259.950 481.050 262.050 ;
        RECT 481.950 250.950 484.050 253.050 ;
        RECT 482.400 244.050 483.600 250.950 ;
        RECT 451.800 241.950 453.900 244.050 ;
        RECT 481.950 241.950 484.050 244.050 ;
        RECT 485.400 241.050 486.600 328.950 ;
        RECT 488.400 325.050 489.600 337.950 ;
        RECT 490.950 330.600 493.050 331.050 ;
        RECT 496.950 330.600 499.050 334.050 ;
        RECT 490.950 330.000 499.050 330.600 ;
        RECT 490.950 329.400 498.600 330.000 ;
        RECT 490.950 328.950 493.050 329.400 ;
        RECT 487.950 322.950 490.050 325.050 ;
        RECT 487.950 316.950 490.050 319.050 ;
        RECT 488.400 295.050 489.600 316.950 ;
        RECT 503.400 310.050 504.600 349.950 ;
        RECT 496.950 307.950 499.050 310.050 ;
        RECT 502.950 307.950 505.050 310.050 ;
        RECT 497.400 295.050 498.600 307.950 ;
        RECT 487.950 292.950 490.050 295.050 ;
        RECT 496.950 292.950 499.050 295.050 ;
        RECT 490.950 274.950 493.050 277.050 ;
        RECT 502.950 274.950 505.050 277.050 ;
        RECT 460.950 238.950 463.050 241.050 ;
        RECT 484.950 238.950 487.050 241.050 ;
        RECT 454.950 229.950 457.050 232.050 ;
        RECT 430.800 223.950 432.900 226.050 ;
        RECT 434.100 223.950 436.200 226.050 ;
        RECT 448.950 223.950 451.050 226.050 ;
        RECT 431.400 220.050 432.600 223.950 ;
        RECT 449.400 220.050 450.600 223.950 ;
        RECT 455.400 220.050 456.600 229.950 ;
        RECT 430.950 217.950 433.050 220.050 ;
        RECT 448.950 217.950 451.050 220.050 ;
        RECT 454.950 217.950 457.050 220.050 ;
        RECT 433.950 207.600 436.050 208.050 ;
        RECT 439.950 207.600 442.050 211.050 ;
        RECT 451.950 208.950 454.050 211.050 ;
        RECT 433.950 207.000 442.050 207.600 ;
        RECT 433.950 206.400 441.600 207.000 ;
        RECT 433.950 205.950 436.050 206.400 ;
        RECT 434.400 199.050 435.600 205.950 ;
        RECT 433.950 196.950 436.050 199.050 ;
        RECT 452.400 193.050 453.600 208.950 ;
        RECT 433.950 190.950 436.050 193.050 ;
        RECT 451.950 190.950 454.050 193.050 ;
        RECT 457.950 190.950 460.050 193.050 ;
        RECT 427.950 187.950 430.050 190.050 ;
        RECT 434.400 184.050 435.600 190.950 ;
        RECT 436.950 187.950 439.050 190.050 ;
        RECT 433.950 181.950 436.050 184.050 ;
        RECT 422.400 176.400 426.600 177.600 ;
        RECT 412.950 172.950 415.050 175.050 ;
        RECT 418.950 172.950 421.050 175.050 ;
        RECT 409.950 148.950 412.050 151.050 ;
        RECT 413.400 148.050 414.600 172.950 ;
        RECT 419.400 160.050 420.600 172.950 ;
        RECT 418.950 157.950 421.050 160.050 ;
        RECT 412.950 145.950 415.050 148.050 ;
        RECT 413.400 130.050 414.600 145.950 ;
        RECT 425.400 145.050 426.600 176.400 ;
        RECT 430.950 172.950 433.050 175.050 ;
        RECT 415.800 142.950 417.900 145.050 ;
        RECT 419.100 142.950 421.200 145.050 ;
        RECT 424.950 142.950 427.050 145.050 ;
        RECT 416.400 139.050 417.600 142.950 ;
        RECT 415.950 136.950 418.050 139.050 ;
        RECT 406.950 127.950 409.050 130.050 ;
        RECT 412.950 127.950 415.050 130.050 ;
        RECT 403.950 121.950 406.050 124.050 ;
        RECT 419.400 115.050 420.600 142.950 ;
        RECT 431.400 130.050 432.600 172.950 ;
        RECT 424.950 127.950 427.050 130.050 ;
        RECT 430.950 127.950 433.050 130.050 ;
        RECT 425.400 124.050 426.600 127.950 ;
        RECT 431.400 124.050 432.600 127.950 ;
        RECT 424.950 121.950 427.050 124.050 ;
        RECT 430.950 121.950 433.050 124.050 ;
        RECT 409.950 112.950 412.050 115.050 ;
        RECT 418.950 112.950 421.050 115.050 ;
        RECT 394.950 109.950 397.050 112.050 ;
        RECT 400.950 109.950 403.050 112.050 ;
        RECT 395.400 106.050 396.600 109.950 ;
        RECT 410.400 109.050 411.600 112.950 ;
        RECT 409.950 106.950 412.050 109.050 ;
        RECT 394.950 103.950 397.050 106.050 ;
        RECT 403.950 105.600 406.050 106.050 ;
        RECT 415.950 105.600 418.050 109.050 ;
        RECT 426.000 105.600 430.050 106.050 ;
        RECT 403.950 105.000 418.050 105.600 ;
        RECT 403.950 104.400 417.600 105.000 ;
        RECT 403.950 103.950 406.050 104.400 ;
        RECT 425.400 103.950 430.050 105.600 ;
        RECT 425.400 100.050 426.600 103.950 ;
        RECT 424.950 97.950 427.050 100.050 ;
        RECT 391.950 94.950 394.050 97.050 ;
        RECT 379.950 88.950 382.050 91.050 ;
        RECT 386.100 88.950 388.200 91.050 ;
        RECT 391.950 88.950 394.050 91.050 ;
        RECT 427.950 88.950 430.050 91.050 ;
        RECT 385.950 82.950 388.050 85.050 ;
        RECT 370.950 79.950 373.050 82.050 ;
        RECT 371.400 55.050 372.600 79.950 ;
        RECT 386.400 70.050 387.600 82.950 ;
        RECT 392.400 70.050 393.600 88.950 ;
        RECT 385.950 67.950 388.050 70.050 ;
        RECT 391.950 67.950 394.050 70.050 ;
        RECT 415.950 67.950 418.050 70.050 ;
        RECT 392.400 64.050 393.600 67.950 ;
        RECT 416.400 64.050 417.600 67.950 ;
        RECT 391.950 61.950 394.050 64.050 ;
        RECT 396.000 63.600 400.050 64.050 ;
        RECT 395.400 61.950 400.050 63.600 ;
        RECT 415.950 61.950 418.050 64.050 ;
        RECT 385.950 60.600 388.050 61.050 ;
        RECT 395.400 60.600 396.600 61.950 ;
        RECT 385.950 59.400 396.600 60.600 ;
        RECT 385.950 58.950 388.050 59.400 ;
        RECT 421.950 58.950 424.050 61.050 ;
        RECT 370.950 52.950 373.050 55.050 ;
        RECT 371.400 49.050 372.600 52.950 ;
        RECT 370.950 46.950 373.050 49.050 ;
        RECT 376.950 37.950 379.050 40.050 ;
        RECT 359.400 35.400 363.600 36.600 ;
        RECT 359.400 21.600 360.600 35.400 ;
        RECT 367.950 34.950 370.050 37.050 ;
        RECT 359.400 20.400 363.600 21.600 ;
        RECT 355.950 16.950 358.050 19.050 ;
        RECT 340.950 13.950 343.050 16.050 ;
        RECT 362.400 13.050 363.600 20.400 ;
        RECT 368.400 19.050 369.600 34.950 ;
        RECT 377.400 28.050 378.600 37.950 ;
        RECT 386.400 28.050 387.600 58.950 ;
        RECT 394.950 52.950 397.050 55.050 ;
        RECT 406.950 52.950 409.050 55.050 ;
        RECT 412.950 54.600 415.050 55.050 ;
        RECT 418.950 54.600 421.050 55.050 ;
        RECT 412.950 53.400 421.050 54.600 ;
        RECT 412.950 52.950 415.050 53.400 ;
        RECT 418.950 52.950 421.050 53.400 ;
        RECT 395.400 49.050 396.600 52.950 ;
        RECT 400.950 49.950 403.050 52.050 ;
        RECT 394.950 46.950 397.050 49.050 ;
        RECT 401.400 40.050 402.600 49.950 ;
        RECT 407.400 49.050 408.600 52.950 ;
        RECT 403.950 47.400 408.600 49.050 ;
        RECT 403.950 46.950 408.000 47.400 ;
        RECT 412.950 46.950 415.050 49.050 ;
        RECT 418.950 46.950 421.050 49.050 ;
        RECT 413.400 43.050 414.600 46.950 ;
        RECT 412.950 40.950 415.050 43.050 ;
        RECT 394.950 37.950 397.050 40.050 ;
        RECT 400.950 37.950 403.050 40.050 ;
        RECT 388.950 30.600 391.050 34.050 ;
        RECT 395.400 30.600 396.600 37.950 ;
        RECT 400.950 30.600 403.050 31.050 ;
        RECT 388.950 30.000 393.600 30.600 ;
        RECT 389.400 29.400 394.050 30.000 ;
        RECT 395.400 29.400 403.050 30.600 ;
        RECT 370.950 25.950 373.050 28.050 ;
        RECT 376.950 25.950 379.050 28.050 ;
        RECT 385.950 25.950 388.050 28.050 ;
        RECT 391.950 25.950 394.050 29.400 ;
        RECT 400.950 28.950 403.050 29.400 ;
        RECT 409.950 28.950 412.050 31.050 ;
        RECT 367.950 16.950 370.050 19.050 ;
        RECT 371.400 18.600 372.600 25.950 ;
        RECT 410.400 22.050 411.600 28.950 ;
        RECT 419.400 22.050 420.600 46.950 ;
        RECT 409.950 19.950 412.050 22.050 ;
        RECT 418.950 19.950 421.050 22.050 ;
        RECT 376.950 18.600 379.050 19.050 ;
        RECT 371.400 17.400 379.050 18.600 ;
        RECT 376.950 16.950 379.050 17.400 ;
        RECT 382.950 16.950 385.050 19.050 ;
        RECT 383.400 13.050 384.600 16.950 ;
        RECT 422.400 13.050 423.600 58.950 ;
        RECT 428.400 46.050 429.600 88.950 ;
        RECT 433.950 85.950 436.050 88.050 ;
        RECT 434.400 61.050 435.600 85.950 ;
        RECT 430.950 58.950 433.050 61.050 ;
        RECT 433.950 58.950 436.050 61.050 ;
        RECT 431.400 49.050 432.600 58.950 ;
        RECT 430.950 46.950 433.050 49.050 ;
        RECT 427.950 43.950 430.050 46.050 ;
        RECT 437.400 37.050 438.600 187.950 ;
        RECT 458.400 184.050 459.600 190.950 ;
        RECT 457.950 181.950 460.050 184.050 ;
        RECT 439.950 151.950 442.050 154.050 ;
        RECT 440.400 88.050 441.600 151.950 ;
        RECT 445.950 145.950 448.050 148.050 ;
        RECT 446.400 142.050 447.600 145.950 ;
        RECT 445.950 139.950 448.050 142.050 ;
        RECT 451.950 139.950 454.050 142.050 ;
        RECT 448.950 130.950 451.050 133.050 ;
        RECT 449.400 127.050 450.600 130.950 ;
        RECT 448.950 124.950 451.050 127.050 ;
        RECT 452.400 124.050 453.600 139.950 ;
        RECT 451.950 121.950 454.050 124.050 ;
        RECT 445.950 118.950 448.050 121.050 ;
        RECT 446.400 100.050 447.600 118.950 ;
        RECT 451.950 109.950 454.050 112.050 ;
        RECT 452.400 106.050 453.600 109.950 ;
        RECT 451.950 103.950 454.050 106.050 ;
        RECT 445.950 97.950 448.050 100.050 ;
        RECT 461.400 88.050 462.600 238.950 ;
        RECT 481.950 235.950 484.050 238.050 ;
        RECT 475.950 232.950 478.050 235.050 ;
        RECT 463.950 223.950 466.050 226.050 ;
        RECT 464.400 190.050 465.600 223.950 ;
        RECT 476.400 217.050 477.600 232.950 ;
        RECT 466.950 214.950 469.050 217.050 ;
        RECT 475.950 214.950 478.050 217.050 ;
        RECT 467.400 199.050 468.600 214.950 ;
        RECT 466.950 196.950 469.050 199.050 ;
        RECT 475.950 196.950 478.050 199.050 ;
        RECT 472.950 193.950 475.050 196.050 ;
        RECT 463.950 187.950 466.050 190.050 ;
        RECT 463.950 181.950 466.050 184.050 ;
        RECT 464.400 115.050 465.600 181.950 ;
        RECT 473.400 157.050 474.600 193.950 ;
        RECT 476.400 178.050 477.600 196.950 ;
        RECT 475.950 175.950 478.050 178.050 ;
        RECT 472.950 154.950 475.050 157.050 ;
        RECT 473.400 142.050 474.600 154.950 ;
        RECT 476.400 154.050 477.600 175.950 ;
        RECT 482.400 163.050 483.600 235.950 ;
        RECT 491.400 193.050 492.600 274.950 ;
        RECT 503.400 262.050 504.600 274.950 ;
        RECT 506.400 271.050 507.600 352.950 ;
        RECT 509.400 319.050 510.600 400.950 ;
        RECT 517.950 376.950 520.050 379.050 ;
        RECT 514.950 366.600 517.050 367.050 ;
        RECT 518.400 366.600 519.600 376.950 ;
        RECT 514.950 366.000 522.600 366.600 ;
        RECT 514.950 365.400 523.050 366.000 ;
        RECT 514.950 364.950 517.050 365.400 ;
        RECT 520.950 361.950 523.050 365.400 ;
        RECT 527.400 355.050 528.600 415.950 ;
        RECT 563.400 411.600 564.600 436.950 ;
        RECT 565.950 427.950 568.050 430.050 ;
        RECT 560.400 411.000 564.600 411.600 ;
        RECT 559.950 410.400 564.600 411.000 ;
        RECT 538.950 406.950 541.050 409.050 ;
        RECT 544.950 406.950 547.050 409.050 ;
        RECT 559.950 406.950 562.050 410.400 ;
        RECT 566.400 409.050 567.600 427.950 ;
        RECT 590.400 426.600 591.600 457.950 ;
        RECT 593.400 445.050 594.600 463.950 ;
        RECT 622.950 460.950 625.050 463.050 ;
        RECT 595.950 453.600 600.000 454.050 ;
        RECT 601.950 453.600 604.050 454.050 ;
        RECT 607.950 453.600 610.050 454.050 ;
        RECT 595.950 451.950 600.600 453.600 ;
        RECT 601.950 452.400 610.050 453.600 ;
        RECT 601.950 451.950 604.050 452.400 ;
        RECT 607.950 451.950 610.050 452.400 ;
        RECT 599.400 450.600 600.600 451.950 ;
        RECT 599.400 449.400 606.600 450.600 ;
        RECT 592.950 442.950 595.050 445.050 ;
        RECT 598.950 439.950 601.050 442.050 ;
        RECT 590.400 425.400 594.600 426.600 ;
        RECT 589.950 418.950 592.050 421.050 ;
        RECT 568.950 415.950 571.050 418.050 ;
        RECT 586.950 417.600 589.050 418.050 ;
        RECT 578.400 416.400 589.050 417.600 ;
        RECT 565.950 406.950 568.050 409.050 ;
        RECT 539.400 397.050 540.600 406.950 ;
        RECT 545.400 403.050 546.600 406.950 ;
        RECT 544.950 400.950 547.050 403.050 ;
        RECT 559.950 400.950 562.050 403.050 ;
        RECT 538.950 394.950 541.050 397.050 ;
        RECT 547.950 375.600 550.050 379.050 ;
        RECT 560.400 376.050 561.600 400.950 ;
        RECT 569.400 397.050 570.600 415.950 ;
        RECT 578.400 397.050 579.600 416.400 ;
        RECT 586.950 415.950 589.050 416.400 ;
        RECT 590.400 414.600 591.600 418.950 ;
        RECT 587.400 413.400 591.600 414.600 ;
        RECT 587.400 411.600 588.600 413.400 ;
        RECT 584.400 411.000 588.600 411.600 ;
        RECT 583.950 410.400 588.600 411.000 ;
        RECT 583.950 406.950 586.050 410.400 ;
        RECT 593.400 409.050 594.600 425.400 ;
        RECT 599.400 421.050 600.600 439.950 ;
        RECT 605.400 436.050 606.600 449.400 ;
        RECT 623.400 445.050 624.600 460.950 ;
        RECT 616.950 442.950 619.050 445.050 ;
        RECT 622.950 442.950 625.050 445.050 ;
        RECT 617.400 439.050 618.600 442.950 ;
        RECT 616.950 436.950 619.050 439.050 ;
        RECT 635.400 436.050 636.600 466.950 ;
        RECT 604.950 433.950 607.050 436.050 ;
        RECT 634.950 433.950 637.050 436.050 ;
        RECT 628.950 430.950 631.050 433.050 ;
        RECT 604.950 427.950 607.050 430.050 ;
        RECT 598.950 418.950 601.050 421.050 ;
        RECT 605.400 418.050 606.600 427.950 ;
        RECT 629.400 418.050 630.600 430.950 ;
        RECT 638.400 424.050 639.600 494.400 ;
        RECT 640.950 493.950 643.050 494.400 ;
        RECT 658.950 493.950 661.050 496.050 ;
        RECT 640.950 487.950 643.050 490.050 ;
        RECT 671.400 489.600 672.600 520.950 ;
        RECT 680.400 517.050 681.600 520.950 ;
        RECT 712.950 517.950 715.050 520.050 ;
        RECT 679.950 514.950 682.050 517.050 ;
        RECT 684.000 495.600 688.050 496.050 ;
        RECT 668.400 489.000 672.600 489.600 ;
        RECT 667.950 488.400 672.600 489.000 ;
        RECT 683.400 493.950 688.050 495.600 ;
        RECT 700.800 495.000 702.900 496.050 ;
        RECT 700.800 493.950 703.050 495.000 ;
        RECT 641.400 469.200 642.600 487.950 ;
        RECT 667.950 484.950 670.050 488.400 ;
        RECT 673.950 484.950 676.050 487.050 ;
        RECT 655.950 478.950 658.050 481.050 ;
        RECT 652.950 469.950 655.050 472.050 ;
        RECT 640.950 467.100 643.050 469.200 ;
        RECT 640.950 463.800 643.050 465.900 ;
        RECT 641.400 454.050 642.600 463.800 ;
        RECT 640.950 451.950 643.050 454.050 ;
        RECT 646.950 451.950 649.050 454.050 ;
        RECT 643.950 442.950 646.050 445.050 ;
        RECT 644.400 436.050 645.600 442.950 ;
        RECT 643.950 433.950 646.050 436.050 ;
        RECT 647.400 433.050 648.600 451.950 ;
        RECT 653.400 436.050 654.600 469.950 ;
        RECT 656.400 454.050 657.600 478.950 ;
        RECT 674.400 475.050 675.600 484.950 ;
        RECT 683.400 481.050 684.600 493.950 ;
        RECT 700.950 492.600 703.050 493.950 ;
        RECT 700.950 492.000 705.600 492.600 ;
        RECT 701.400 491.400 705.600 492.000 ;
        RECT 688.950 484.950 691.050 487.050 ;
        RECT 694.950 484.950 697.050 487.050 ;
        RECT 682.950 478.950 685.050 481.050 ;
        RECT 689.400 478.050 690.600 484.950 ;
        RECT 695.400 481.050 696.600 484.950 ;
        RECT 694.950 478.950 697.050 481.050 ;
        RECT 688.950 475.950 691.050 478.050 ;
        RECT 695.400 475.050 696.600 478.950 ;
        RECT 673.950 472.950 676.050 475.050 ;
        RECT 694.950 472.950 697.050 475.050 ;
        RECT 704.400 466.050 705.600 491.400 ;
        RECT 713.400 487.050 714.600 517.950 ;
        RECT 719.400 514.050 720.600 529.950 ;
        RECT 718.950 511.950 721.050 514.050 ;
        RECT 724.950 511.950 727.050 514.050 ;
        RECT 725.400 505.050 726.600 511.950 ;
        RECT 724.950 502.950 727.050 505.050 ;
        RECT 721.950 496.050 724.050 499.050 ;
        RECT 718.950 495.000 724.050 496.050 ;
        RECT 718.950 494.400 723.600 495.000 ;
        RECT 718.950 493.950 723.000 494.400 ;
        RECT 725.400 487.050 726.600 502.950 ;
        RECT 731.400 499.050 732.600 529.950 ;
        RECT 741.000 528.600 745.050 529.050 ;
        RECT 740.400 526.950 745.050 528.600 ;
        RECT 740.400 517.050 741.600 526.950 ;
        RECT 746.400 520.050 747.600 532.800 ;
        RECT 755.400 529.050 756.600 550.950 ;
        RECT 757.950 541.950 760.050 544.050 ;
        RECT 748.950 526.950 751.050 529.050 ;
        RECT 754.950 526.950 757.050 529.050 ;
        RECT 745.950 517.950 748.050 520.050 ;
        RECT 739.950 514.950 742.050 517.050 ;
        RECT 749.400 508.050 750.600 526.950 ;
        RECT 739.950 505.950 742.050 508.050 ;
        RECT 748.950 505.950 751.050 508.050 ;
        RECT 740.400 499.050 741.600 505.950 ;
        RECT 758.400 502.050 759.600 541.950 ;
        RECT 761.400 508.050 762.600 562.950 ;
        RECT 763.950 559.950 766.050 562.050 ;
        RECT 764.400 514.050 765.600 559.950 ;
        RECT 773.400 547.050 774.600 571.950 ;
        RECT 772.950 544.950 775.050 547.050 ;
        RECT 779.400 544.050 780.600 571.950 ;
        RECT 785.400 556.050 786.600 586.950 ;
        RECT 788.400 583.050 789.600 589.950 ;
        RECT 787.950 580.950 790.050 583.050 ;
        RECT 802.950 574.050 805.050 577.050 ;
        RECT 799.950 573.000 805.050 574.050 ;
        RECT 799.950 572.400 804.600 573.000 ;
        RECT 799.950 571.950 804.000 572.400 ;
        RECT 794.400 566.400 801.600 567.600 ;
        RECT 784.950 553.950 787.050 556.050 ;
        RECT 784.950 544.950 787.050 547.050 ;
        RECT 778.950 541.950 781.050 544.050 ;
        RECT 772.950 538.950 775.050 541.050 ;
        RECT 773.400 532.050 774.600 538.950 ;
        RECT 778.950 535.950 781.050 538.050 ;
        RECT 779.400 532.050 780.600 535.950 ;
        RECT 772.950 529.950 775.050 532.050 ;
        RECT 778.950 529.950 781.050 532.050 ;
        RECT 775.950 520.950 778.050 523.050 ;
        RECT 763.950 511.950 766.050 514.050 ;
        RECT 776.400 511.050 777.600 520.950 ;
        RECT 781.950 511.950 784.050 514.050 ;
        RECT 775.950 508.950 778.050 511.050 ;
        RECT 760.950 505.950 763.050 508.050 ;
        RECT 757.950 499.950 760.050 502.050 ;
        RECT 763.950 499.950 766.050 502.050 ;
        RECT 769.950 499.950 772.050 502.050 ;
        RECT 727.950 497.400 732.600 499.050 ;
        RECT 727.950 496.950 732.000 497.400 ;
        RECT 733.950 496.950 736.050 499.050 ;
        RECT 739.950 496.950 742.050 499.050 ;
        RECT 727.950 487.950 730.050 490.050 ;
        RECT 713.400 485.400 718.050 487.050 ;
        RECT 714.000 484.950 718.050 485.400 ;
        RECT 721.950 485.400 726.600 487.050 ;
        RECT 721.950 484.950 726.000 485.400 ;
        RECT 716.400 481.050 717.600 484.950 ;
        RECT 715.950 478.950 718.050 481.050 ;
        RECT 703.950 463.950 706.050 466.050 ;
        RECT 664.950 460.950 667.050 463.050 ;
        RECT 694.950 460.950 697.050 463.050 ;
        RECT 665.400 454.050 666.600 460.950 ;
        RECT 656.400 451.950 661.050 454.050 ;
        RECT 664.950 451.950 667.050 454.050 ;
        RECT 652.950 433.950 655.050 436.050 ;
        RECT 656.400 433.050 657.600 451.950 ;
        RECT 685.950 448.950 688.050 451.050 ;
        RECT 661.950 442.950 664.050 445.050 ;
        RECT 676.950 442.950 679.050 445.050 ;
        RECT 662.400 436.050 663.600 442.950 ;
        RECT 661.950 433.950 664.050 436.050 ;
        RECT 646.950 430.950 649.050 433.050 ;
        RECT 655.950 430.950 658.050 433.050 ;
        RECT 677.400 427.050 678.600 442.950 ;
        RECT 686.400 436.050 687.600 448.950 ;
        RECT 688.950 442.950 691.050 445.050 ;
        RECT 685.950 433.950 688.050 436.050 ;
        RECT 682.950 430.950 685.050 433.050 ;
        RECT 676.950 424.950 679.050 427.050 ;
        RECT 637.950 421.950 640.050 424.050 ;
        RECT 658.950 421.950 661.050 424.050 ;
        RECT 638.400 418.050 639.600 421.950 ;
        RECT 659.400 418.050 660.600 421.950 ;
        RECT 683.400 418.050 684.600 430.950 ;
        RECT 604.950 415.950 607.050 418.050 ;
        RECT 622.950 415.950 625.050 418.050 ;
        RECT 628.950 415.950 631.050 418.050 ;
        RECT 634.950 416.400 639.600 418.050 ;
        RECT 634.950 415.950 639.000 416.400 ;
        RECT 649.950 415.950 652.050 418.050 ;
        RECT 658.950 415.950 661.050 418.050 ;
        RECT 682.950 415.950 685.050 418.050 ;
        RECT 589.950 407.400 594.600 409.050 ;
        RECT 589.950 406.950 594.000 407.400 ;
        RECT 595.950 406.950 598.050 409.050 ;
        RECT 583.950 400.950 586.050 403.050 ;
        RECT 568.950 394.950 571.050 397.050 ;
        RECT 577.950 394.950 580.050 397.050 ;
        RECT 553.950 375.600 556.050 376.050 ;
        RECT 547.950 375.000 556.050 375.600 ;
        RECT 548.400 374.400 556.050 375.000 ;
        RECT 553.950 373.950 556.050 374.400 ;
        RECT 559.950 373.950 562.050 376.050 ;
        RECT 573.000 375.600 577.050 376.050 ;
        RECT 579.000 375.600 583.050 376.050 ;
        RECT 572.400 373.950 577.050 375.600 ;
        RECT 578.400 373.950 583.050 375.600 ;
        RECT 572.400 367.050 573.600 373.950 ;
        RECT 578.400 372.600 579.600 373.950 ;
        RECT 575.400 371.400 579.600 372.600 ;
        RECT 571.950 364.950 574.050 367.050 ;
        RECT 535.950 361.950 538.050 364.050 ;
        RECT 526.950 352.950 529.050 355.050 ;
        RECT 536.400 352.050 537.600 361.950 ;
        RECT 571.950 358.950 574.050 361.050 ;
        RECT 535.950 349.950 538.050 352.050 ;
        RECT 511.950 346.950 514.050 349.050 ;
        RECT 512.400 343.050 513.600 346.950 ;
        RECT 511.950 340.950 514.050 343.050 ;
        RECT 517.950 340.950 520.050 343.050 ;
        RECT 518.400 339.600 519.600 340.950 ;
        RECT 523.950 339.600 526.050 340.050 ;
        RECT 518.400 338.400 526.050 339.600 ;
        RECT 508.950 316.950 511.050 319.050 ;
        RECT 509.400 298.050 510.600 316.950 ;
        RECT 518.400 298.050 519.600 338.400 ;
        RECT 523.950 337.950 526.050 338.400 ;
        RECT 572.400 334.050 573.600 358.950 ;
        RECT 575.400 355.050 576.600 371.400 ;
        RECT 584.400 367.050 585.600 400.950 ;
        RECT 596.400 397.050 597.600 406.950 ;
        RECT 623.400 400.050 624.600 415.950 ;
        RECT 631.950 408.600 634.050 409.050 ;
        RECT 637.950 408.600 640.050 409.050 ;
        RECT 631.950 407.400 640.050 408.600 ;
        RECT 631.950 406.950 634.050 407.400 ;
        RECT 637.950 406.950 640.050 407.400 ;
        RECT 643.950 406.950 646.050 409.050 ;
        RECT 622.950 397.950 625.050 400.050 ;
        RECT 595.950 394.950 598.050 397.050 ;
        RECT 644.400 385.050 645.600 406.950 ;
        RECT 643.950 382.950 646.050 385.050 ;
        RECT 650.400 382.050 651.600 415.950 ;
        RECT 673.950 406.950 676.050 409.050 ;
        RECT 652.950 382.950 655.050 385.050 ;
        RECT 649.950 379.950 652.050 382.050 ;
        RECT 598.950 372.600 601.050 376.050 ;
        RECT 634.950 375.600 637.050 379.050 ;
        RECT 653.400 376.050 654.600 382.950 ;
        RECT 658.950 379.950 661.050 382.050 ;
        RECT 659.400 376.050 660.600 379.950 ;
        RECT 674.400 379.050 675.600 406.950 ;
        RECT 686.400 385.050 687.600 433.950 ;
        RECT 689.400 397.050 690.600 442.950 ;
        RECT 688.950 394.950 691.050 397.050 ;
        RECT 685.950 382.950 688.050 385.050 ;
        RECT 673.950 376.950 676.050 379.050 ;
        RECT 632.400 375.000 637.050 375.600 ;
        RECT 632.400 374.400 636.600 375.000 ;
        RECT 625.950 372.600 628.050 373.050 ;
        RECT 632.400 372.600 633.600 374.400 ;
        RECT 652.950 373.950 655.050 376.050 ;
        RECT 658.950 373.950 661.050 376.050 ;
        RECT 598.950 372.000 603.600 372.600 ;
        RECT 599.400 371.400 603.600 372.000 ;
        RECT 577.950 364.950 580.050 367.050 ;
        RECT 583.950 364.950 586.050 367.050 ;
        RECT 595.950 364.950 598.050 367.050 ;
        RECT 578.400 361.050 579.600 364.950 ;
        RECT 577.950 358.950 580.050 361.050 ;
        RECT 574.950 352.950 577.050 355.050 ;
        RECT 596.400 352.050 597.600 364.950 ;
        RECT 602.400 355.050 603.600 371.400 ;
        RECT 625.950 371.400 633.600 372.600 ;
        RECT 625.950 370.950 628.050 371.400 ;
        RECT 634.950 370.950 637.050 373.050 ;
        RECT 664.950 370.950 667.050 373.050 ;
        RECT 607.950 364.950 610.050 367.050 ;
        RECT 601.950 352.950 604.050 355.050 ;
        RECT 586.950 349.950 589.050 352.050 ;
        RECT 595.950 349.950 598.050 352.050 ;
        RECT 587.400 340.050 588.600 349.950 ;
        RECT 596.400 343.050 597.600 349.950 ;
        RECT 608.400 349.050 609.600 364.950 ;
        RECT 607.950 346.950 610.050 349.050 ;
        RECT 631.950 346.950 634.050 349.050 ;
        RECT 608.400 343.050 609.600 346.950 ;
        RECT 595.950 340.950 598.050 343.050 ;
        RECT 607.950 340.950 610.050 343.050 ;
        RECT 586.950 337.950 589.050 340.050 ;
        RECT 541.950 331.950 544.050 334.050 ;
        RECT 542.400 328.050 543.600 331.950 ;
        RECT 550.950 330.600 553.050 334.050 ;
        RECT 559.950 331.950 562.050 334.050 ;
        RECT 571.950 331.950 574.050 334.050 ;
        RECT 550.950 330.000 555.600 330.600 ;
        RECT 551.400 329.400 555.600 330.000 ;
        RECT 520.950 327.600 523.050 328.050 ;
        RECT 532.950 327.600 535.050 328.050 ;
        RECT 520.950 326.400 535.050 327.600 ;
        RECT 520.950 325.950 523.050 326.400 ;
        RECT 532.950 325.950 535.050 326.400 ;
        RECT 541.950 325.950 544.050 328.050 ;
        RECT 523.950 313.950 526.050 316.050 ;
        RECT 509.400 296.400 514.050 298.050 ;
        RECT 510.000 295.950 514.050 296.400 ;
        RECT 517.950 295.950 520.050 298.050 ;
        RECT 514.950 283.950 517.050 286.050 ;
        RECT 505.950 268.950 508.050 271.050 ;
        RECT 496.950 258.600 499.050 262.050 ;
        RECT 502.950 259.950 505.050 262.050 ;
        RECT 511.950 259.950 514.050 262.050 ;
        RECT 508.950 258.600 511.050 259.050 ;
        RECT 496.950 258.000 511.050 258.600 ;
        RECT 497.400 257.400 511.050 258.000 ;
        RECT 508.950 256.950 511.050 257.400 ;
        RECT 493.950 252.600 496.050 253.050 ;
        RECT 499.950 252.600 502.050 253.050 ;
        RECT 493.950 251.400 502.050 252.600 ;
        RECT 493.950 250.950 496.050 251.400 ;
        RECT 499.950 250.950 502.050 251.400 ;
        RECT 505.950 250.950 508.050 253.050 ;
        RECT 506.400 247.050 507.600 250.950 ;
        RECT 493.950 244.950 496.050 247.050 ;
        RECT 505.950 244.950 508.050 247.050 ;
        RECT 494.400 232.050 495.600 244.950 ;
        RECT 505.950 232.950 508.050 235.050 ;
        RECT 493.950 229.950 496.050 232.050 ;
        RECT 499.950 220.950 502.050 223.050 ;
        RECT 493.950 210.600 496.050 211.050 ;
        RECT 500.400 210.600 501.600 220.950 ;
        RECT 506.400 217.050 507.600 232.950 ;
        RECT 512.400 229.050 513.600 259.950 ;
        RECT 515.400 247.050 516.600 283.950 ;
        RECT 524.400 280.050 525.600 313.950 ;
        RECT 554.400 310.050 555.600 329.400 ;
        RECT 560.400 316.050 561.600 331.950 ;
        RECT 632.400 331.050 633.600 346.950 ;
        RECT 604.950 328.950 607.050 331.050 ;
        RECT 631.950 328.950 634.050 331.050 ;
        RECT 559.950 313.950 562.050 316.050 ;
        RECT 577.950 310.950 580.050 313.050 ;
        RECT 535.950 307.950 538.050 310.050 ;
        RECT 553.950 307.950 556.050 310.050 ;
        RECT 526.950 286.950 529.050 289.050 ;
        RECT 517.950 277.950 520.050 280.050 ;
        RECT 523.950 277.950 526.050 280.050 ;
        RECT 518.400 262.050 519.600 277.950 ;
        RECT 520.950 274.950 523.050 277.050 ;
        RECT 521.400 271.050 522.600 274.950 ;
        RECT 520.950 268.950 523.050 271.050 ;
        RECT 527.400 268.050 528.600 286.950 ;
        RECT 526.950 265.950 529.050 268.050 ;
        RECT 518.400 260.400 523.050 262.050 ;
        RECT 519.000 259.950 523.050 260.400 ;
        RECT 536.400 256.050 537.600 307.950 ;
        RECT 554.400 301.050 555.600 307.950 ;
        RECT 553.950 298.950 556.050 301.050 ;
        RECT 554.400 295.050 555.600 298.950 ;
        RECT 538.950 292.950 541.050 295.050 ;
        RECT 553.950 292.950 556.050 295.050 ;
        RECT 539.400 274.050 540.600 292.950 ;
        RECT 538.950 271.950 541.050 274.050 ;
        RECT 544.950 271.950 547.050 274.050 ;
        RECT 545.400 256.050 546.600 271.950 ;
        RECT 578.400 262.050 579.600 310.950 ;
        RECT 583.950 271.950 586.050 274.050 ;
        RECT 584.400 265.050 585.600 271.950 ;
        RECT 605.400 271.050 606.600 328.950 ;
        RECT 635.400 316.050 636.600 370.950 ;
        RECT 665.400 367.050 666.600 370.950 ;
        RECT 649.950 364.950 652.050 367.050 ;
        RECT 661.950 365.400 666.600 367.050 ;
        RECT 661.950 364.950 666.000 365.400 ;
        RECT 637.950 352.950 640.050 355.050 ;
        RECT 638.400 343.050 639.600 352.950 ;
        RECT 646.950 348.600 649.050 349.050 ;
        RECT 650.400 348.600 651.600 364.950 ;
        RECT 674.400 364.050 675.600 376.950 ;
        RECT 685.950 373.950 688.050 376.050 ;
        RECT 686.400 364.050 687.600 373.950 ;
        RECT 674.400 362.400 679.050 364.050 ;
        RECT 675.000 361.950 679.050 362.400 ;
        RECT 682.950 362.400 687.600 364.050 ;
        RECT 682.950 361.950 687.000 362.400 ;
        RECT 695.400 358.050 696.600 460.950 ;
        RECT 704.400 445.050 705.600 463.950 ;
        RECT 728.400 463.050 729.600 487.950 ;
        RECT 734.400 484.050 735.600 496.950 ;
        RECT 764.400 496.050 765.600 499.950 ;
        RECT 745.950 493.950 748.050 496.050 ;
        RECT 763.950 493.950 766.050 496.050 ;
        RECT 746.400 484.050 747.600 493.950 ;
        RECT 770.400 487.050 771.600 499.950 ;
        RECT 782.400 487.050 783.600 511.950 ;
        RECT 760.950 484.950 763.050 487.050 ;
        RECT 766.950 485.400 771.600 487.050 ;
        RECT 766.950 484.950 771.000 485.400 ;
        RECT 781.950 484.950 784.050 487.050 ;
        RECT 733.950 481.950 736.050 484.050 ;
        RECT 745.950 481.950 748.050 484.050 ;
        RECT 734.400 478.050 735.600 481.950 ;
        RECT 761.400 481.050 762.600 484.950 ;
        RECT 760.950 478.950 763.050 481.050 ;
        RECT 733.950 475.950 736.050 478.050 ;
        RECT 782.400 472.050 783.600 484.950 ;
        RECT 781.950 469.950 784.050 472.050 ;
        RECT 727.950 460.950 730.050 463.050 ;
        RECT 751.950 460.950 754.050 463.050 ;
        RECT 733.950 457.950 736.050 460.050 ;
        RECT 745.950 457.950 748.050 460.050 ;
        RECT 734.400 454.050 735.600 457.950 ;
        RECT 746.400 454.050 747.600 457.950 ;
        RECT 752.400 454.050 753.600 460.950 ;
        RECT 778.950 454.050 781.050 457.050 ;
        RECT 709.950 451.950 712.050 454.050 ;
        RECT 727.950 451.950 730.050 454.050 ;
        RECT 733.950 451.950 736.050 454.050 ;
        RECT 745.950 451.950 748.050 454.050 ;
        RECT 751.950 451.950 754.050 454.050 ;
        RECT 769.950 451.950 772.050 454.050 ;
        RECT 775.950 453.000 781.050 454.050 ;
        RECT 775.950 452.400 780.600 453.000 ;
        RECT 775.950 451.950 780.000 452.400 ;
        RECT 703.950 442.950 706.050 445.050 ;
        RECT 697.950 424.950 700.050 427.050 ;
        RECT 703.950 424.950 706.050 427.050 ;
        RECT 698.400 421.050 699.600 424.950 ;
        RECT 704.400 421.050 705.600 424.950 ;
        RECT 710.400 421.050 711.600 451.950 ;
        RECT 715.950 442.950 718.050 445.050 ;
        RECT 716.400 427.050 717.600 442.950 ;
        RECT 728.400 430.050 729.600 451.950 ;
        RECT 730.950 442.950 733.050 445.050 ;
        RECT 731.400 436.050 732.600 442.950 ;
        RECT 752.400 436.050 753.600 451.950 ;
        RECT 766.950 442.950 769.050 445.050 ;
        RECT 730.950 433.950 733.050 436.050 ;
        RECT 751.950 433.950 754.050 436.050 ;
        RECT 727.950 427.950 730.050 430.050 ;
        RECT 715.950 424.950 718.050 427.050 ;
        RECT 697.950 418.950 700.050 421.050 ;
        RECT 703.950 418.950 706.050 421.050 ;
        RECT 709.950 418.950 712.050 421.050 ;
        RECT 716.400 418.050 717.600 424.950 ;
        RECT 767.400 421.050 768.600 442.950 ;
        RECT 770.400 433.050 771.600 451.950 ;
        RECT 782.400 451.050 783.600 469.950 ;
        RECT 781.950 448.950 784.050 451.050 ;
        RECT 778.950 444.600 781.050 445.050 ;
        RECT 785.400 444.600 786.600 544.950 ;
        RECT 794.400 537.600 795.600 566.400 ;
        RECT 800.400 565.050 801.600 566.400 ;
        RECT 796.950 562.950 799.050 565.050 ;
        RECT 800.400 563.400 805.050 565.050 ;
        RECT 801.000 562.950 805.050 563.400 ;
        RECT 797.400 553.050 798.600 562.950 ;
        RECT 796.950 550.950 799.050 553.050 ;
        RECT 809.400 552.600 810.600 598.950 ;
        RECT 824.400 595.050 825.600 598.950 ;
        RECT 823.950 592.950 826.050 595.050 ;
        RECT 826.950 589.950 829.050 592.050 ;
        RECT 823.950 586.950 826.050 589.050 ;
        RECT 820.950 583.950 823.050 586.050 ;
        RECT 817.950 580.950 820.050 583.050 ;
        RECT 818.400 574.050 819.600 580.950 ;
        RECT 817.950 571.950 820.050 574.050 ;
        RECT 821.400 565.050 822.600 583.950 ;
        RECT 814.950 562.950 817.050 565.050 ;
        RECT 820.950 562.950 823.050 565.050 ;
        RECT 806.400 551.400 810.600 552.600 ;
        RECT 806.400 544.050 807.600 551.400 ;
        RECT 815.400 547.050 816.600 562.950 ;
        RECT 821.400 553.050 822.600 562.950 ;
        RECT 820.950 550.950 823.050 553.050 ;
        RECT 808.950 544.950 811.050 547.050 ;
        RECT 814.950 544.950 817.050 547.050 ;
        RECT 805.950 541.950 808.050 544.050 ;
        RECT 809.400 538.050 810.600 544.950 ;
        RECT 796.950 537.600 799.050 538.050 ;
        RECT 794.400 536.400 799.050 537.600 ;
        RECT 796.950 535.950 799.050 536.400 ;
        RECT 802.950 535.950 805.050 538.050 ;
        RECT 808.950 535.950 811.050 538.050 ;
        RECT 814.950 535.950 817.050 538.050 ;
        RECT 797.400 523.050 798.600 535.950 ;
        RECT 803.400 532.050 804.600 535.950 ;
        RECT 809.400 532.050 810.600 535.950 ;
        RECT 815.400 532.050 816.600 535.950 ;
        RECT 802.950 529.950 805.050 532.050 ;
        RECT 808.950 529.950 811.050 532.050 ;
        RECT 814.950 529.950 817.050 532.050 ;
        RECT 796.950 520.950 799.050 523.050 ;
        RECT 811.950 520.950 814.050 523.050 ;
        RECT 812.400 517.050 813.600 520.950 ;
        RECT 811.950 514.950 814.050 517.050 ;
        RECT 805.950 511.950 808.050 514.050 ;
        RECT 787.950 505.950 790.050 508.050 ;
        RECT 788.400 487.050 789.600 505.950 ;
        RECT 806.400 496.050 807.600 511.950 ;
        RECT 812.400 511.050 813.600 514.950 ;
        RECT 811.950 508.950 814.050 511.050 ;
        RECT 796.950 493.950 799.050 496.050 ;
        RECT 805.950 493.950 808.050 496.050 ;
        RECT 797.400 490.050 798.600 493.950 ;
        RECT 797.400 488.400 802.050 490.050 ;
        RECT 798.000 487.950 802.050 488.400 ;
        RECT 787.950 484.950 790.050 487.050 ;
        RECT 788.400 466.050 789.600 484.950 ;
        RECT 787.950 463.950 790.050 466.050 ;
        RECT 800.400 451.050 801.600 487.950 ;
        RECT 812.400 481.050 813.600 508.950 ;
        RECT 824.400 505.050 825.600 586.950 ;
        RECT 827.400 517.050 828.600 589.950 ;
        RECT 830.400 538.050 831.600 611.400 ;
        RECT 836.400 610.050 837.600 622.950 ;
        RECT 839.400 622.050 840.600 634.950 ;
        RECT 844.950 628.950 847.050 631.050 ;
        RECT 841.950 625.950 844.050 628.050 ;
        RECT 838.950 619.950 841.050 622.050 ;
        RECT 832.950 608.400 837.600 610.050 ;
        RECT 832.950 607.950 837.000 608.400 ;
        RECT 842.400 606.600 843.600 625.950 ;
        RECT 845.400 610.050 846.600 628.950 ;
        RECT 848.400 625.050 849.600 640.950 ;
        RECT 851.400 625.050 852.600 668.400 ;
        RECT 847.800 622.950 849.900 625.050 ;
        RECT 851.100 622.950 853.200 625.050 ;
        RECT 848.400 619.050 849.600 622.950 ;
        RECT 854.400 621.600 855.600 673.950 ;
        RECT 859.800 670.950 861.900 673.050 ;
        RECT 863.100 670.950 865.200 673.050 ;
        RECT 856.950 664.950 859.050 667.050 ;
        RECT 857.400 628.050 858.600 664.950 ;
        RECT 860.400 651.600 861.600 670.950 ;
        RECT 863.400 661.050 864.600 670.950 ;
        RECT 866.400 661.050 867.600 754.950 ;
        RECT 869.400 730.050 870.600 761.400 ;
        RECT 880.950 745.950 883.050 748.050 ;
        RECT 868.950 727.950 871.050 730.050 ;
        RECT 868.950 718.950 871.050 721.050 ;
        RECT 874.950 720.600 879.000 721.050 ;
        RECT 874.950 718.950 879.600 720.600 ;
        RECT 869.400 715.050 870.600 718.950 ;
        RECT 868.950 712.950 871.050 715.050 ;
        RECT 878.400 703.050 879.600 718.950 ;
        RECT 877.950 700.950 880.050 703.050 ;
        RECT 871.950 697.950 874.050 700.050 ;
        RECT 872.400 679.050 873.600 697.950 ;
        RECT 881.400 697.050 882.600 745.950 ;
        RECT 887.400 736.050 888.600 766.950 ;
        RECT 890.400 742.050 891.600 784.950 ;
        RECT 889.950 739.950 892.050 742.050 ;
        RECT 893.400 739.050 894.600 790.950 ;
        RECT 905.400 772.050 906.600 799.950 ;
        RECT 904.950 769.950 907.050 772.050 ;
        RECT 911.400 769.050 912.600 823.950 ;
        RECT 910.950 766.950 913.050 769.050 ;
        RECT 910.950 760.950 913.050 763.050 ;
        RECT 895.950 757.800 898.050 759.900 ;
        RECT 896.400 741.600 897.600 757.800 ;
        RECT 898.950 751.950 901.050 754.050 ;
        RECT 904.950 751.950 907.050 754.050 ;
        RECT 899.400 748.050 900.600 751.950 ;
        RECT 905.400 748.050 906.600 751.950 ;
        RECT 898.950 745.950 901.050 748.050 ;
        RECT 904.950 745.950 907.050 748.050 ;
        RECT 896.400 741.000 900.600 741.600 ;
        RECT 896.400 740.400 901.050 741.000 ;
        RECT 892.950 736.950 895.050 739.050 ;
        RECT 898.950 736.950 901.050 740.400 ;
        RECT 904.950 739.950 907.050 742.050 ;
        RECT 886.950 733.950 889.050 736.050 ;
        RECT 889.950 730.050 892.050 733.050 ;
        RECT 886.950 727.950 889.050 730.050 ;
        RECT 889.950 729.000 895.050 730.050 ;
        RECT 890.400 728.400 895.050 729.000 ;
        RECT 891.000 727.950 895.050 728.400 ;
        RECT 898.950 727.950 901.050 730.050 ;
        RECT 887.400 700.050 888.600 727.950 ;
        RECT 899.400 723.600 900.600 727.950 ;
        RECT 893.400 722.400 900.600 723.600 ;
        RECT 889.950 718.950 892.050 721.050 ;
        RECT 890.400 715.050 891.600 718.950 ;
        RECT 889.950 712.950 892.050 715.050 ;
        RECT 886.950 697.950 889.050 700.050 ;
        RECT 893.400 699.600 894.600 722.400 ;
        RECT 901.950 721.950 904.050 724.050 ;
        RECT 895.950 718.950 898.050 721.050 ;
        RECT 896.400 703.050 897.600 718.950 ;
        RECT 895.950 700.950 898.050 703.050 ;
        RECT 890.400 698.400 894.600 699.600 ;
        RECT 880.950 694.950 883.050 697.050 ;
        RECT 883.950 691.950 886.050 694.050 ;
        RECT 884.400 688.050 885.600 691.950 ;
        RECT 874.950 687.600 879.000 688.050 ;
        RECT 880.950 687.600 885.600 688.050 ;
        RECT 874.950 685.950 879.600 687.600 ;
        RECT 880.950 686.400 888.600 687.600 ;
        RECT 880.950 685.950 885.000 686.400 ;
        RECT 878.400 684.600 879.600 685.950 ;
        RECT 878.400 684.000 885.600 684.600 ;
        RECT 878.400 683.400 886.050 684.000 ;
        RECT 883.950 679.950 886.050 683.400 ;
        RECT 871.950 676.950 874.050 679.050 ;
        RECT 877.950 673.950 880.050 676.050 ;
        RECT 878.400 670.050 879.600 673.950 ;
        RECT 877.950 667.950 880.050 670.050 ;
        RECT 862.800 658.950 864.900 661.050 ;
        RECT 866.100 658.950 868.200 661.050 ;
        RECT 880.950 658.950 883.050 661.050 ;
        RECT 874.950 652.050 877.050 655.050 ;
        RECT 860.400 650.400 867.600 651.600 ;
        RECT 866.400 645.600 867.600 650.400 ;
        RECT 871.950 651.000 877.050 652.050 ;
        RECT 871.950 650.400 876.600 651.000 ;
        RECT 871.950 649.950 876.000 650.400 ;
        RECT 866.400 644.400 873.600 645.600 ;
        RECT 872.400 643.050 873.600 644.400 ;
        RECT 868.950 640.950 871.050 643.050 ;
        RECT 872.400 641.400 877.050 643.050 ;
        RECT 873.000 640.950 877.050 641.400 ;
        RECT 869.400 637.050 870.600 640.950 ;
        RECT 881.400 637.050 882.600 658.950 ;
        RECT 887.400 658.050 888.600 686.400 ;
        RECT 890.400 678.600 891.600 698.400 ;
        RECT 902.400 682.050 903.600 721.950 ;
        RECT 905.400 694.050 906.600 739.950 ;
        RECT 908.100 706.950 910.200 709.050 ;
        RECT 908.400 703.050 909.600 706.950 ;
        RECT 907.950 700.950 910.050 703.050 ;
        RECT 911.400 700.050 912.600 760.950 ;
        RECT 910.950 697.950 913.050 700.050 ;
        RECT 904.950 691.950 907.050 694.050 ;
        RECT 910.950 691.950 913.050 694.050 ;
        RECT 901.950 679.950 904.050 682.050 ;
        RECT 907.950 679.950 910.050 682.050 ;
        RECT 895.950 678.600 898.050 679.050 ;
        RECT 890.400 677.400 898.050 678.600 ;
        RECT 886.950 655.950 889.050 658.050 ;
        RECT 890.400 652.050 891.600 677.400 ;
        RECT 895.950 676.950 898.050 677.400 ;
        RECT 898.950 670.950 901.050 673.050 ;
        RECT 895.950 655.950 898.050 658.050 ;
        RECT 889.950 649.950 892.050 652.050 ;
        RECT 886.950 640.950 889.050 643.050 ;
        RECT 887.400 637.050 888.600 640.950 ;
        RECT 868.950 634.950 871.050 637.050 ;
        RECT 880.950 634.950 883.050 637.050 ;
        RECT 886.950 634.950 889.050 637.050 ;
        RECT 856.950 625.950 859.050 628.050 ;
        RECT 880.950 625.950 883.050 628.050 ;
        RECT 859.950 622.950 862.050 625.050 ;
        RECT 854.400 620.400 858.600 621.600 ;
        RECT 847.950 616.950 850.050 619.050 ;
        RECT 853.950 616.950 856.050 619.050 ;
        RECT 854.400 610.050 855.600 616.950 ;
        RECT 845.400 608.400 850.050 610.050 ;
        RECT 846.000 607.950 850.050 608.400 ;
        RECT 853.950 607.950 856.050 610.050 ;
        RECT 842.400 605.400 846.600 606.600 ;
        RECT 835.950 598.950 838.050 601.050 ;
        RECT 836.400 541.050 837.600 598.950 ;
        RECT 845.400 589.050 846.600 605.400 ;
        RECT 850.950 592.950 853.050 595.050 ;
        RECT 844.950 586.950 847.050 589.050 ;
        RECT 844.950 571.950 847.050 574.050 ;
        RECT 845.400 556.050 846.600 571.950 ;
        RECT 844.950 553.950 847.050 556.050 ;
        RECT 835.950 538.950 838.050 541.050 ;
        RECT 844.950 538.950 847.050 541.050 ;
        RECT 829.950 535.950 832.050 538.050 ;
        RECT 838.950 535.950 841.050 538.050 ;
        RECT 839.400 523.050 840.600 535.950 ;
        RECT 832.950 520.950 835.050 523.050 ;
        RECT 838.950 520.950 841.050 523.050 ;
        RECT 826.950 514.950 829.050 517.050 ;
        RECT 823.950 502.950 826.050 505.050 ;
        RECT 833.400 502.050 834.600 520.950 ;
        RECT 841.950 514.950 844.050 517.050 ;
        RECT 832.950 499.950 835.050 502.050 ;
        RECT 833.400 496.050 834.600 499.950 ;
        RECT 820.950 493.950 823.050 496.050 ;
        RECT 832.950 493.950 835.050 496.050 ;
        RECT 811.950 478.950 814.050 481.050 ;
        RECT 808.950 469.950 811.050 472.050 ;
        RECT 809.400 466.050 810.600 469.950 ;
        RECT 814.950 466.950 817.050 469.050 ;
        RECT 808.950 463.950 811.050 466.050 ;
        RECT 815.400 454.050 816.600 466.950 ;
        RECT 817.950 463.950 820.050 466.050 ;
        RECT 818.400 454.050 819.600 463.950 ;
        RECT 821.400 463.050 822.600 493.950 ;
        RECT 823.950 487.950 826.050 490.050 ;
        RECT 824.400 466.050 825.600 487.950 ;
        RECT 829.950 484.950 832.050 487.050 ;
        RECT 835.950 484.950 838.050 487.050 ;
        RECT 830.400 478.050 831.600 484.950 ;
        RECT 836.400 481.050 837.600 484.950 ;
        RECT 835.950 478.950 838.050 481.050 ;
        RECT 829.950 475.950 832.050 478.050 ;
        RECT 835.950 472.950 838.050 475.050 ;
        RECT 826.950 466.950 829.050 469.050 ;
        RECT 823.950 463.950 826.050 466.050 ;
        RECT 820.950 460.950 823.050 463.050 ;
        RECT 827.400 454.050 828.600 466.950 ;
        RECT 814.950 451.950 817.050 454.050 ;
        RECT 818.400 452.400 823.050 454.050 ;
        RECT 819.000 451.950 823.050 452.400 ;
        RECT 826.950 451.950 829.050 454.050 ;
        RECT 787.950 448.950 790.050 451.050 ;
        RECT 799.950 448.950 802.050 451.050 ;
        RECT 808.950 450.600 813.000 451.050 ;
        RECT 808.950 448.950 813.600 450.600 ;
        RECT 778.950 443.400 786.600 444.600 ;
        RECT 788.400 445.050 789.600 448.950 ;
        RECT 788.400 443.400 793.050 445.050 ;
        RECT 778.950 442.950 781.050 443.400 ;
        RECT 789.000 442.950 793.050 443.400 ;
        RECT 796.950 441.600 799.050 445.050 ;
        RECT 812.400 444.600 813.600 448.950 ;
        RECT 817.950 444.600 820.050 445.050 ;
        RECT 812.400 443.400 820.050 444.600 ;
        RECT 817.950 442.950 820.050 443.400 ;
        RECT 832.950 442.950 835.050 445.050 ;
        RECT 794.400 441.000 799.050 441.600 ;
        RECT 794.400 440.400 798.600 441.000 ;
        RECT 769.950 430.950 772.050 433.050 ;
        RECT 772.950 427.950 775.050 430.050 ;
        RECT 759.000 420.600 763.050 421.050 ;
        RECT 758.400 418.950 763.050 420.600 ;
        RECT 766.950 418.950 769.050 421.050 ;
        RECT 715.950 415.950 718.050 418.050 ;
        RECT 745.950 415.950 748.050 418.050 ;
        RECT 709.950 409.950 712.050 412.050 ;
        RECT 703.950 400.950 706.050 403.050 ;
        RECT 697.950 397.950 700.050 400.050 ;
        RECT 698.400 376.050 699.600 397.950 ;
        RECT 704.400 376.050 705.600 400.950 ;
        RECT 710.400 382.050 711.600 409.950 ;
        RECT 717.000 408.600 721.050 409.050 ;
        RECT 716.400 408.000 721.050 408.600 ;
        RECT 715.950 406.950 721.050 408.000 ;
        RECT 724.950 408.600 729.000 409.050 ;
        RECT 724.950 406.950 729.600 408.600 ;
        RECT 715.950 403.950 718.050 406.950 ;
        RECT 728.400 403.050 729.600 406.950 ;
        RECT 727.950 400.950 730.050 403.050 ;
        RECT 733.950 400.950 736.050 403.050 ;
        RECT 724.950 397.950 727.050 400.050 ;
        RECT 709.950 379.950 712.050 382.050 ;
        RECT 721.950 379.950 724.050 382.050 ;
        RECT 722.400 376.050 723.600 379.950 ;
        RECT 697.950 373.950 700.050 376.050 ;
        RECT 703.950 373.950 706.050 376.050 ;
        RECT 721.950 373.950 724.050 376.050 ;
        RECT 725.400 367.050 726.600 397.950 ;
        RECT 727.950 394.950 730.050 397.050 ;
        RECT 728.400 376.050 729.600 394.950 ;
        RECT 734.400 394.050 735.600 400.950 ;
        RECT 746.400 400.050 747.600 415.950 ;
        RECT 758.400 409.050 759.600 418.950 ;
        RECT 773.400 412.050 774.600 427.950 ;
        RECT 781.950 424.950 784.050 427.050 ;
        RECT 782.400 421.050 783.600 424.950 ;
        RECT 781.950 418.950 784.050 421.050 ;
        RECT 787.950 418.950 790.050 421.050 ;
        RECT 769.800 409.950 771.900 412.050 ;
        RECT 773.100 409.950 775.200 412.050 ;
        RECT 757.950 406.950 760.050 409.050 ;
        RECT 745.950 397.950 748.050 400.050 ;
        RECT 733.950 391.950 736.050 394.050 ;
        RECT 770.400 382.200 771.600 409.950 ;
        RECT 788.400 403.050 789.600 418.950 ;
        RECT 787.950 400.950 790.050 403.050 ;
        RECT 794.400 400.050 795.600 440.400 ;
        RECT 833.400 439.050 834.600 442.950 ;
        RECT 808.950 436.950 811.050 439.050 ;
        RECT 832.950 436.950 835.050 439.050 ;
        RECT 799.800 433.950 801.900 436.050 ;
        RECT 796.950 430.950 799.050 433.050 ;
        RECT 797.400 420.600 798.600 430.950 ;
        RECT 800.400 423.600 801.600 433.950 ;
        RECT 800.400 422.400 804.600 423.600 ;
        RECT 797.400 420.000 801.600 420.600 ;
        RECT 797.400 419.400 802.050 420.000 ;
        RECT 799.950 415.950 802.050 419.400 ;
        RECT 803.400 409.050 804.600 422.400 ;
        RECT 809.400 409.050 810.600 436.950 ;
        RECT 823.950 417.600 826.050 421.050 ;
        RECT 829.950 420.600 834.000 421.050 ;
        RECT 829.950 418.950 834.600 420.600 ;
        RECT 823.950 417.000 828.600 417.600 ;
        RECT 824.400 416.400 828.600 417.000 ;
        RECT 814.950 409.950 817.050 412.050 ;
        RECT 802.950 406.950 805.050 409.050 ;
        RECT 808.950 406.950 811.050 409.050 ;
        RECT 793.950 397.950 796.050 400.050 ;
        RECT 769.950 380.100 772.050 382.200 ;
        RECT 794.400 382.050 795.600 397.950 ;
        RECT 808.950 394.950 811.050 397.050 ;
        RECT 802.950 388.950 805.050 391.050 ;
        RECT 787.950 379.950 790.050 382.050 ;
        RECT 793.950 379.950 796.050 382.050 ;
        RECT 748.950 376.950 751.050 379.050 ;
        RECT 757.950 378.600 760.050 379.050 ;
        RECT 769.950 378.600 772.050 378.900 ;
        RECT 757.950 377.400 772.050 378.600 ;
        RECT 757.950 376.950 760.050 377.400 ;
        RECT 727.950 373.950 730.050 376.050 ;
        RECT 749.400 373.050 750.600 376.950 ;
        RECT 769.950 376.800 772.050 377.400 ;
        RECT 739.950 370.950 742.050 373.050 ;
        RECT 748.950 370.950 751.050 373.050 ;
        RECT 780.000 372.600 784.050 373.050 ;
        RECT 779.400 370.950 784.050 372.600 ;
        RECT 700.950 364.950 703.050 367.050 ;
        RECT 709.950 364.950 712.050 367.050 ;
        RECT 724.950 364.950 727.050 367.050 ;
        RECT 736.950 364.950 739.050 367.050 ;
        RECT 701.400 361.050 702.600 364.950 ;
        RECT 700.950 358.950 703.050 361.050 ;
        RECT 664.950 355.950 667.050 358.050 ;
        RECT 694.950 355.950 697.050 358.050 ;
        RECT 646.950 347.400 651.600 348.600 ;
        RECT 646.950 346.950 649.050 347.400 ;
        RECT 647.400 343.050 648.600 346.950 ;
        RECT 637.950 340.950 640.050 343.050 ;
        RECT 646.950 340.950 649.050 343.050 ;
        RECT 665.400 340.050 666.600 355.950 ;
        RECT 685.950 349.950 688.050 352.050 ;
        RECT 686.400 346.050 687.600 349.950 ;
        RECT 676.950 343.950 679.050 346.050 ;
        RECT 664.950 337.950 667.050 340.050 ;
        RECT 640.950 331.950 643.050 334.050 ;
        RECT 625.950 313.950 628.050 316.050 ;
        RECT 634.950 313.950 637.050 316.050 ;
        RECT 610.950 295.950 613.050 298.050 ;
        RECT 616.950 295.950 619.050 298.050 ;
        RECT 607.950 286.950 610.050 289.050 ;
        RECT 608.400 277.050 609.600 286.950 ;
        RECT 607.950 274.950 610.050 277.050 ;
        RECT 611.400 273.600 612.600 295.950 ;
        RECT 617.400 274.050 618.600 295.950 ;
        RECT 626.400 295.050 627.600 313.950 ;
        RECT 625.950 292.950 628.050 295.050 ;
        RECT 634.950 294.600 637.050 295.050 ;
        RECT 629.400 293.400 637.050 294.600 ;
        RECT 629.400 291.600 630.600 293.400 ;
        RECT 634.950 292.950 637.050 293.400 ;
        RECT 623.400 291.000 630.600 291.600 ;
        RECT 622.950 290.400 630.600 291.000 ;
        RECT 622.950 286.950 625.050 290.400 ;
        RECT 608.400 272.400 612.600 273.600 ;
        RECT 604.950 268.950 607.050 271.050 ;
        RECT 583.950 262.950 586.050 265.050 ;
        RECT 562.950 261.600 567.000 262.050 ;
        RECT 562.950 259.950 567.600 261.600 ;
        RECT 577.950 259.950 580.050 262.050 ;
        RECT 589.950 259.950 592.050 262.050 ;
        RECT 529.950 253.950 532.050 256.050 ;
        RECT 535.950 253.950 538.050 256.050 ;
        RECT 544.950 253.950 547.050 256.050 ;
        RECT 530.400 250.050 531.600 253.950 ;
        RECT 529.950 247.950 532.050 250.050 ;
        RECT 514.950 244.950 517.050 247.050 ;
        RECT 517.950 241.950 520.050 244.050 ;
        RECT 511.950 226.950 514.050 229.050 ;
        RECT 518.400 219.600 519.600 241.950 ;
        RECT 523.950 229.950 526.050 232.050 ;
        RECT 518.400 218.400 522.600 219.600 ;
        RECT 505.950 214.950 508.050 217.050 ;
        RECT 493.950 210.000 501.600 210.600 ;
        RECT 493.950 209.400 502.050 210.000 ;
        RECT 493.950 208.950 496.050 209.400 ;
        RECT 499.950 205.950 502.050 209.400 ;
        RECT 513.000 207.600 517.050 208.050 ;
        RECT 512.400 205.950 517.050 207.600 ;
        RECT 512.400 193.050 513.600 205.950 ;
        RECT 490.950 190.950 493.050 193.050 ;
        RECT 511.950 190.950 514.050 193.050 ;
        RECT 508.950 178.950 511.050 181.050 ;
        RECT 509.400 175.050 510.600 178.950 ;
        RECT 521.400 175.050 522.600 218.400 ;
        RECT 493.950 172.950 496.050 175.050 ;
        RECT 505.950 172.950 508.050 175.050 ;
        RECT 509.400 173.400 514.050 175.050 ;
        RECT 510.000 172.950 514.050 173.400 ;
        RECT 517.950 173.400 522.600 175.050 ;
        RECT 517.950 172.950 522.000 173.400 ;
        RECT 481.950 160.950 484.050 163.050 ;
        RECT 475.950 151.950 478.050 154.050 ;
        RECT 478.950 145.950 481.050 148.050 ;
        RECT 479.400 142.050 480.600 145.950 ;
        RECT 472.950 139.950 475.050 142.050 ;
        RECT 478.950 139.950 481.050 142.050 ;
        RECT 482.400 138.600 483.600 160.950 ;
        RECT 494.400 157.050 495.600 172.950 ;
        RECT 506.400 163.050 507.600 172.950 ;
        RECT 520.950 163.950 523.050 166.050 ;
        RECT 505.950 160.950 508.050 163.050 ;
        RECT 521.400 160.050 522.600 163.950 ;
        RECT 520.950 157.950 523.050 160.050 ;
        RECT 493.950 154.950 496.050 157.050 ;
        RECT 502.950 154.950 505.050 157.050 ;
        RECT 487.950 151.950 490.050 154.050 ;
        RECT 479.400 137.400 483.600 138.600 ;
        RECT 470.100 130.950 472.200 133.050 ;
        RECT 463.950 112.950 466.050 115.050 ;
        RECT 470.400 106.050 471.600 130.950 ;
        RECT 479.400 129.600 480.600 137.400 ;
        RECT 481.950 132.600 486.000 133.050 ;
        RECT 481.950 130.950 486.600 132.600 ;
        RECT 479.400 128.400 483.600 129.600 ;
        RECT 478.950 112.950 481.050 115.050 ;
        RECT 479.400 106.050 480.600 112.950 ;
        RECT 482.400 108.600 483.600 128.400 ;
        RECT 485.400 112.050 486.600 130.950 ;
        RECT 488.400 118.050 489.600 151.950 ;
        RECT 493.950 127.950 496.050 130.050 ;
        RECT 499.950 127.950 502.050 130.050 ;
        RECT 487.950 115.950 490.050 118.050 ;
        RECT 484.950 109.950 487.050 112.050 ;
        RECT 494.400 109.050 495.600 127.950 ;
        RECT 496.950 121.950 499.050 124.050 ;
        RECT 482.400 107.400 486.600 108.600 ;
        RECT 469.950 103.950 472.050 106.050 ;
        RECT 478.800 103.950 480.900 106.050 ;
        RECT 482.100 103.950 484.200 106.050 ;
        RECT 466.950 96.600 469.050 100.050 ;
        RECT 482.400 97.050 483.600 103.950 ;
        RECT 472.950 96.600 475.050 97.050 ;
        RECT 466.950 96.000 475.050 96.600 ;
        RECT 467.400 95.400 475.050 96.000 ;
        RECT 472.950 94.950 475.050 95.400 ;
        RECT 478.950 95.400 483.600 97.050 ;
        RECT 478.950 94.950 483.000 95.400 ;
        RECT 439.800 85.950 441.900 88.050 ;
        RECT 443.100 85.950 445.200 88.050 ;
        RECT 460.800 85.950 462.900 88.050 ;
        RECT 472.950 85.950 475.050 88.050 ;
        RECT 443.400 61.050 444.600 85.950 ;
        RECT 461.400 61.050 462.600 85.950 ;
        RECT 473.400 70.050 474.600 85.950 ;
        RECT 478.950 76.950 481.050 79.050 ;
        RECT 472.950 67.950 475.050 70.050 ;
        RECT 479.400 61.050 480.600 76.950 ;
        RECT 485.400 64.050 486.600 107.400 ;
        RECT 493.950 106.950 496.050 109.050 ;
        RECT 497.400 97.050 498.600 121.950 ;
        RECT 500.400 112.050 501.600 127.950 ;
        RECT 503.400 124.050 504.600 154.950 ;
        RECT 514.950 148.950 517.050 151.050 ;
        RECT 520.950 148.950 523.050 151.050 ;
        RECT 508.950 145.950 511.050 148.050 ;
        RECT 509.400 139.050 510.600 145.950 ;
        RECT 515.400 142.050 516.600 148.950 ;
        RECT 521.400 142.050 522.600 148.950 ;
        RECT 514.950 139.950 517.050 142.050 ;
        RECT 520.950 139.950 523.050 142.050 ;
        RECT 508.950 136.950 511.050 139.050 ;
        RECT 524.400 138.600 525.600 229.950 ;
        RECT 530.400 226.050 531.600 247.950 ;
        RECT 566.400 247.050 567.600 259.950 ;
        RECT 590.400 253.050 591.600 259.950 ;
        RECT 608.400 253.050 609.600 272.400 ;
        RECT 616.950 271.950 619.050 274.050 ;
        RECT 641.400 271.050 642.600 331.950 ;
        RECT 677.400 331.050 678.600 343.950 ;
        RECT 685.950 343.050 688.050 346.050 ;
        RECT 685.950 342.000 691.050 343.050 ;
        RECT 693.000 342.600 697.050 343.050 ;
        RECT 686.400 341.400 691.050 342.000 ;
        RECT 687.000 340.950 691.050 341.400 ;
        RECT 692.400 340.950 697.050 342.600 ;
        RECT 682.950 339.600 685.050 340.050 ;
        RECT 692.400 339.600 693.600 340.950 ;
        RECT 682.950 338.400 693.600 339.600 ;
        RECT 682.950 337.950 685.050 338.400 ;
        RECT 685.950 331.950 688.050 334.050 ;
        RECT 697.950 331.950 700.050 334.050 ;
        RECT 661.950 328.950 664.050 331.050 ;
        RECT 667.950 328.950 670.050 331.050 ;
        RECT 676.950 328.950 679.050 331.050 ;
        RECT 662.400 325.050 663.600 328.950 ;
        RECT 661.950 322.950 664.050 325.050 ;
        RECT 655.950 295.950 658.050 298.050 ;
        RECT 656.400 289.050 657.600 295.950 ;
        RECT 668.400 294.600 669.600 328.950 ;
        RECT 686.400 321.600 687.600 331.950 ;
        RECT 691.950 328.950 694.050 331.050 ;
        RECT 686.400 320.400 690.600 321.600 ;
        RECT 673.950 295.950 676.050 298.050 ;
        RECT 668.400 293.400 672.600 294.600 ;
        RECT 652.950 286.950 657.600 289.050 ;
        RECT 664.950 286.950 667.050 289.050 ;
        RECT 656.400 277.050 657.600 286.950 ;
        RECT 655.950 274.950 658.050 277.050 ;
        RECT 665.400 274.050 666.600 286.950 ;
        RECT 664.950 271.950 667.050 274.050 ;
        RECT 671.400 271.050 672.600 293.400 ;
        RECT 622.950 268.950 625.050 271.050 ;
        RECT 628.950 268.950 631.050 271.050 ;
        RECT 640.950 268.950 643.050 271.050 ;
        RECT 652.950 268.950 655.050 271.050 ;
        RECT 670.950 268.950 673.050 271.050 ;
        RECT 623.400 265.050 624.600 268.950 ;
        RECT 629.400 265.050 630.600 268.950 ;
        RECT 622.950 262.950 625.050 265.050 ;
        RECT 628.950 262.950 631.050 265.050 ;
        RECT 619.950 253.950 622.050 256.050 ;
        RECT 580.950 250.950 583.050 253.050 ;
        RECT 586.950 251.400 591.600 253.050 ;
        RECT 586.950 250.950 591.000 251.400 ;
        RECT 607.950 250.950 610.050 253.050 ;
        RECT 565.950 244.950 568.050 247.050 ;
        RECT 581.400 241.050 582.600 250.950 ;
        RECT 608.400 241.050 609.600 250.950 ;
        RECT 580.950 238.950 583.050 241.050 ;
        RECT 607.950 238.950 610.050 241.050 ;
        RECT 559.950 232.950 562.050 235.050 ;
        RECT 613.950 232.950 616.050 235.050 ;
        RECT 547.950 226.950 550.050 229.050 ;
        RECT 529.950 223.950 532.050 226.050 ;
        RECT 538.950 223.950 541.050 226.050 ;
        RECT 526.950 219.600 529.050 223.050 ;
        RECT 539.400 220.050 540.600 223.950 ;
        RECT 532.950 219.600 535.050 220.050 ;
        RECT 526.950 219.000 535.050 219.600 ;
        RECT 527.400 218.400 535.050 219.000 ;
        RECT 532.950 217.950 535.050 218.400 ;
        RECT 538.950 217.950 541.050 220.050 ;
        RECT 539.400 202.050 540.600 217.950 ;
        RECT 538.950 199.950 541.050 202.050 ;
        RECT 539.400 196.050 540.600 199.950 ;
        RECT 548.400 199.050 549.600 226.950 ;
        RECT 560.400 220.050 561.600 232.950 ;
        RECT 614.400 220.050 615.600 232.950 ;
        RECT 552.000 219.600 556.050 220.050 ;
        RECT 551.400 217.950 556.050 219.600 ;
        RECT 559.950 217.950 562.050 220.050 ;
        RECT 613.950 217.950 616.050 220.050 ;
        RECT 551.400 211.050 552.600 217.950 ;
        RECT 568.950 216.600 571.050 217.050 ;
        RECT 554.400 215.400 571.050 216.600 ;
        RECT 550.950 208.950 553.050 211.050 ;
        RECT 547.950 196.950 550.050 199.050 ;
        RECT 554.400 196.050 555.600 215.400 ;
        RECT 568.950 214.950 571.050 215.400 ;
        RECT 577.950 214.950 580.050 217.050 ;
        RECT 556.950 208.950 559.050 211.050 ;
        RECT 562.950 208.950 565.050 211.050 ;
        RECT 557.400 205.050 558.600 208.950 ;
        RECT 556.950 202.950 559.050 205.050 ;
        RECT 563.400 202.050 564.600 208.950 ;
        RECT 578.400 207.600 579.600 214.950 ;
        RECT 595.950 208.950 598.050 211.050 ;
        RECT 610.950 208.950 613.050 211.050 ;
        RECT 572.400 206.400 579.600 207.600 ;
        RECT 565.950 204.600 568.050 205.050 ;
        RECT 572.400 204.600 573.600 206.400 ;
        RECT 565.950 203.400 573.600 204.600 ;
        RECT 565.950 202.950 568.050 203.400 ;
        RECT 562.950 201.600 565.050 202.050 ;
        RECT 560.400 200.400 565.050 201.600 ;
        RECT 538.950 193.950 541.050 196.050 ;
        RECT 553.950 193.950 556.050 196.050 ;
        RECT 526.950 181.950 529.050 184.050 ;
        RECT 527.400 163.050 528.600 181.950 ;
        RECT 554.400 178.050 555.600 193.950 ;
        RECT 544.950 175.950 547.050 178.050 ;
        RECT 553.950 175.950 556.050 178.050 ;
        RECT 526.950 160.950 529.050 163.050 ;
        RECT 545.400 160.050 546.600 175.950 ;
        RECT 544.950 157.950 547.050 160.050 ;
        RECT 526.950 148.950 529.050 151.050 ;
        RECT 544.950 148.950 547.050 151.050 ;
        RECT 521.400 137.400 525.600 138.600 ;
        RECT 508.950 124.950 511.050 127.050 ;
        RECT 502.950 121.950 505.050 124.050 ;
        RECT 499.950 109.950 502.050 112.050 ;
        RECT 509.400 100.050 510.600 124.950 ;
        RECT 517.950 115.950 520.050 118.050 ;
        RECT 518.400 100.050 519.600 115.950 ;
        RECT 508.950 97.950 511.050 100.050 ;
        RECT 517.950 97.950 520.050 100.050 ;
        RECT 495.000 96.600 499.050 97.050 ;
        RECT 494.400 94.950 499.050 96.600 ;
        RECT 487.950 88.950 490.050 91.050 ;
        RECT 484.950 61.950 487.050 64.050 ;
        RECT 442.950 58.950 445.050 61.050 ;
        RECT 461.400 59.400 466.050 61.050 ;
        RECT 462.000 58.950 466.050 59.400 ;
        RECT 472.950 58.950 475.050 61.050 ;
        RECT 478.950 58.950 481.050 61.050 ;
        RECT 463.950 52.950 466.050 55.050 ;
        RECT 464.400 40.050 465.600 52.950 ;
        RECT 473.400 52.050 474.600 58.950 ;
        RECT 488.400 54.600 489.600 88.950 ;
        RECT 494.400 85.050 495.600 94.950 ;
        RECT 502.950 93.600 505.050 94.050 ;
        RECT 517.950 93.600 520.050 94.050 ;
        RECT 502.950 92.400 520.050 93.600 ;
        RECT 502.950 91.950 505.050 92.400 ;
        RECT 517.950 91.950 520.050 92.400 ;
        RECT 494.100 82.950 496.200 85.050 ;
        RECT 499.950 82.950 502.050 85.050 ;
        RECT 482.400 54.000 489.600 54.600 ;
        RECT 481.950 53.400 489.600 54.000 ;
        RECT 473.400 50.400 478.050 52.050 ;
        RECT 474.000 49.950 478.050 50.400 ;
        RECT 481.950 49.950 484.050 53.400 ;
        RECT 487.950 46.950 490.050 49.050 ;
        RECT 469.950 43.950 472.050 46.050 ;
        RECT 466.950 40.950 469.050 43.050 ;
        RECT 457.950 37.950 460.050 40.050 ;
        RECT 463.950 37.950 466.050 40.050 ;
        RECT 436.950 34.950 439.050 37.050 ;
        RECT 458.400 31.050 459.600 37.950 ;
        RECT 467.400 31.050 468.600 40.950 ;
        RECT 457.950 28.950 460.050 31.050 ;
        RECT 463.950 29.400 468.600 31.050 ;
        RECT 463.950 28.950 468.000 29.400 ;
        RECT 470.400 27.600 471.600 43.950 ;
        RECT 488.400 31.050 489.600 46.950 ;
        RECT 500.400 43.050 501.600 82.950 ;
        RECT 521.400 64.050 522.600 137.400 ;
        RECT 527.400 133.050 528.600 148.950 ;
        RECT 538.950 145.950 541.050 148.050 ;
        RECT 539.400 142.050 540.600 145.950 ;
        RECT 545.400 142.050 546.600 148.950 ;
        RECT 538.950 139.950 541.050 142.050 ;
        RECT 544.950 139.950 547.050 142.050 ;
        RECT 523.800 130.950 525.900 133.050 ;
        RECT 527.100 130.950 529.200 133.050 ;
        RECT 524.400 124.050 525.600 130.950 ;
        RECT 554.400 127.050 555.600 175.950 ;
        RECT 560.400 142.050 561.600 200.400 ;
        RECT 562.950 199.950 565.050 200.400 ;
        RECT 596.400 199.050 597.600 208.950 ;
        RECT 601.950 202.950 604.050 205.050 ;
        RECT 580.950 196.950 583.050 199.050 ;
        RECT 595.950 196.950 598.050 199.050 ;
        RECT 574.950 190.950 577.050 193.050 ;
        RECT 575.400 184.050 576.600 190.950 ;
        RECT 574.950 181.950 577.050 184.050 ;
        RECT 571.950 169.950 574.050 172.050 ;
        RECT 565.950 151.950 568.050 154.050 ;
        RECT 566.400 142.050 567.600 151.950 ;
        RECT 559.950 139.950 562.050 142.050 ;
        RECT 565.950 139.950 568.050 142.050 ;
        RECT 572.400 133.050 573.600 169.950 ;
        RECT 581.400 163.050 582.600 196.950 ;
        RECT 586.950 181.950 589.050 184.050 ;
        RECT 595.950 181.950 598.050 184.050 ;
        RECT 580.950 160.950 583.050 163.050 ;
        RECT 568.950 131.400 573.600 133.050 ;
        RECT 568.950 130.950 573.000 131.400 ;
        RECT 553.950 124.950 556.050 127.050 ;
        RECT 523.950 121.950 526.050 124.050 ;
        RECT 554.400 115.050 555.600 124.950 ;
        RECT 565.950 115.950 568.050 118.050 ;
        RECT 553.950 112.950 556.050 115.050 ;
        RECT 562.950 112.950 565.050 115.050 ;
        RECT 550.950 109.950 553.050 112.050 ;
        RECT 551.400 106.050 552.600 109.950 ;
        RECT 535.950 105.600 538.050 106.050 ;
        RECT 527.400 104.400 538.050 105.600 ;
        RECT 527.400 94.050 528.600 104.400 ;
        RECT 535.950 103.950 538.050 104.400 ;
        RECT 544.950 103.950 547.050 106.050 ;
        RECT 550.950 103.950 553.050 106.050 ;
        RECT 545.400 94.050 546.600 103.950 ;
        RECT 563.400 99.600 564.600 112.950 ;
        RECT 566.400 106.050 567.600 115.950 ;
        RECT 581.400 106.050 582.600 160.950 ;
        RECT 583.950 145.950 586.050 148.050 ;
        RECT 584.400 142.050 585.600 145.950 ;
        RECT 583.950 139.950 586.050 142.050 ;
        RECT 587.400 121.050 588.600 181.950 ;
        RECT 592.950 172.950 595.050 175.050 ;
        RECT 593.400 169.050 594.600 172.950 ;
        RECT 592.950 166.950 595.050 169.050 ;
        RECT 596.400 166.050 597.600 181.950 ;
        RECT 598.950 172.950 601.050 175.050 ;
        RECT 589.950 163.950 592.050 166.050 ;
        RECT 595.950 163.950 598.050 166.050 ;
        RECT 590.400 142.050 591.600 163.950 ;
        RECT 599.400 142.050 600.600 172.950 ;
        RECT 602.400 169.050 603.600 202.950 ;
        RECT 611.400 202.050 612.600 208.950 ;
        RECT 610.950 199.950 613.050 202.050 ;
        RECT 620.400 193.050 621.600 253.950 ;
        RECT 631.950 223.950 634.050 226.050 ;
        RECT 632.400 220.050 633.600 223.950 ;
        RECT 653.400 220.050 654.600 268.950 ;
        RECT 667.950 265.950 670.050 268.050 ;
        RECT 661.950 235.950 664.050 238.050 ;
        RECT 662.400 229.050 663.600 235.950 ;
        RECT 668.400 232.050 669.600 265.950 ;
        RECT 674.400 241.050 675.600 295.950 ;
        RECT 682.950 286.950 685.050 289.050 ;
        RECT 683.400 265.050 684.600 286.950 ;
        RECT 682.950 262.950 685.050 265.050 ;
        RECT 679.950 259.950 682.050 262.050 ;
        RECT 673.950 238.950 676.050 241.050 ;
        RECT 667.800 229.950 669.900 232.050 ;
        RECT 671.100 231.600 673.200 232.050 ;
        RECT 674.400 231.600 675.600 238.950 ;
        RECT 671.100 230.400 675.600 231.600 ;
        RECT 671.100 229.950 673.200 230.400 ;
        RECT 661.950 226.950 664.050 229.050 ;
        RECT 664.950 220.050 667.050 223.050 ;
        RECT 625.950 217.950 628.050 220.050 ;
        RECT 631.950 217.950 634.050 220.050 ;
        RECT 637.950 219.600 642.000 220.050 ;
        RECT 653.400 219.600 658.050 220.050 ;
        RECT 637.950 217.950 642.600 219.600 ;
        RECT 626.400 211.050 627.600 217.950 ;
        RECT 641.400 211.050 642.600 217.950 ;
        RECT 650.400 218.400 658.050 219.600 ;
        RECT 626.400 209.400 631.050 211.050 ;
        RECT 627.000 208.950 631.050 209.400 ;
        RECT 640.950 208.950 643.050 211.050 ;
        RECT 619.950 190.950 622.050 193.050 ;
        RECT 643.950 190.950 646.050 193.050 ;
        RECT 620.400 187.050 621.600 190.950 ;
        RECT 637.950 187.950 640.050 190.050 ;
        RECT 613.950 183.600 616.050 187.050 ;
        RECT 619.950 184.950 622.050 187.050 ;
        RECT 638.400 184.050 639.600 187.950 ;
        RECT 611.400 183.000 616.050 183.600 ;
        RECT 611.400 182.400 615.600 183.000 ;
        RECT 611.400 175.050 612.600 182.400 ;
        RECT 637.950 181.950 640.050 184.050 ;
        RECT 644.400 178.050 645.600 190.950 ;
        RECT 619.800 175.950 621.900 178.050 ;
        RECT 643.950 175.950 646.050 178.050 ;
        RECT 610.950 172.950 613.050 175.050 ;
        RECT 611.400 169.050 612.600 172.950 ;
        RECT 601.950 166.950 604.050 169.050 ;
        RECT 610.950 166.950 613.050 169.050 ;
        RECT 602.400 151.050 603.600 166.950 ;
        RECT 607.950 151.950 610.050 154.050 ;
        RECT 601.950 148.950 604.050 151.050 ;
        RECT 589.950 139.950 592.050 142.050 ;
        RECT 598.950 139.950 601.050 142.050 ;
        RECT 608.400 133.050 609.600 151.950 ;
        RECT 620.400 142.050 621.600 175.950 ;
        RECT 650.400 166.050 651.600 218.400 ;
        RECT 654.000 217.950 658.050 218.400 ;
        RECT 661.950 219.000 667.050 220.050 ;
        RECT 661.950 218.400 666.600 219.000 ;
        RECT 661.950 217.950 666.000 218.400 ;
        RECT 664.950 208.950 667.050 211.050 ;
        RECT 665.400 205.050 666.600 208.950 ;
        RECT 664.950 202.950 667.050 205.050 ;
        RECT 658.950 190.950 661.050 193.050 ;
        RECT 659.400 184.050 660.600 190.950 ;
        RECT 667.950 187.950 670.050 190.050 ;
        RECT 658.950 181.950 661.050 184.050 ;
        RECT 668.400 178.050 669.600 187.950 ;
        RECT 667.950 175.950 670.050 178.050 ;
        RECT 655.950 172.950 658.050 175.050 ;
        RECT 661.950 172.950 664.050 175.050 ;
        RECT 656.400 169.050 657.600 172.950 ;
        RECT 655.950 166.950 658.050 169.050 ;
        RECT 662.400 166.050 663.600 172.950 ;
        RECT 649.950 163.950 652.050 166.050 ;
        RECT 661.950 163.950 664.050 166.050 ;
        RECT 640.950 154.950 643.050 157.050 ;
        RECT 620.400 140.400 625.050 142.050 ;
        RECT 621.000 139.950 625.050 140.400 ;
        RECT 628.950 141.600 633.000 142.050 ;
        RECT 628.950 139.950 633.600 141.600 ;
        RECT 632.400 133.050 633.600 139.950 ;
        RECT 601.950 130.950 604.050 133.050 ;
        RECT 607.950 130.950 610.050 133.050 ;
        RECT 619.950 130.950 622.050 133.050 ;
        RECT 631.950 130.950 634.050 133.050 ;
        RECT 586.950 118.950 589.050 121.050 ;
        RECT 602.400 108.600 603.600 130.950 ;
        RECT 608.400 115.050 609.600 130.950 ;
        RECT 620.400 127.050 621.600 130.950 ;
        RECT 641.400 127.050 642.600 154.950 ;
        RECT 646.950 151.950 649.050 154.050 ;
        RECT 647.400 142.050 648.600 151.950 ;
        RECT 646.950 139.950 649.050 142.050 ;
        RECT 655.950 139.950 658.050 142.050 ;
        RECT 656.400 133.050 657.600 139.950 ;
        RECT 656.400 130.950 661.050 133.050 ;
        RECT 619.950 124.950 622.050 127.050 ;
        RECT 640.950 124.950 643.050 127.050 ;
        RECT 656.400 118.050 657.600 130.950 ;
        RECT 655.950 115.950 658.050 118.050 ;
        RECT 671.400 115.050 672.600 229.950 ;
        RECT 680.400 223.050 681.600 259.950 ;
        RECT 689.400 253.050 690.600 320.400 ;
        RECT 692.400 301.050 693.600 328.950 ;
        RECT 698.400 322.050 699.600 331.950 ;
        RECT 710.400 331.050 711.600 364.950 ;
        RECT 715.950 355.950 718.050 358.050 ;
        RECT 716.400 340.050 717.600 355.950 ;
        RECT 737.400 355.050 738.600 364.950 ;
        RECT 736.950 352.950 739.050 355.050 ;
        RECT 715.950 337.950 718.050 340.050 ;
        RECT 718.950 331.950 721.050 334.050 ;
        RECT 730.950 331.950 733.050 334.050 ;
        RECT 710.400 329.400 715.050 331.050 ;
        RECT 711.000 328.950 715.050 329.400 ;
        RECT 713.400 325.050 714.600 328.950 ;
        RECT 712.950 322.950 715.050 325.050 ;
        RECT 719.400 322.050 720.600 331.950 ;
        RECT 697.950 319.950 700.050 322.050 ;
        RECT 718.950 319.950 721.050 322.050 ;
        RECT 724.950 316.950 727.050 319.050 ;
        RECT 709.950 313.950 712.050 316.050 ;
        RECT 691.950 298.950 694.050 301.050 ;
        RECT 700.950 298.950 703.050 301.050 ;
        RECT 701.400 295.050 702.600 298.950 ;
        RECT 710.400 295.050 711.600 313.950 ;
        RECT 721.950 307.950 724.050 310.050 ;
        RECT 700.950 292.950 703.050 295.050 ;
        RECT 709.950 292.950 712.050 295.050 ;
        RECT 722.400 289.050 723.600 307.950 ;
        RECT 725.400 298.050 726.600 316.950 ;
        RECT 731.400 316.050 732.600 331.950 ;
        RECT 740.400 316.050 741.600 370.950 ;
        RECT 766.950 364.950 769.050 367.050 ;
        RECT 760.950 343.950 763.050 346.050 ;
        RECT 761.400 340.050 762.600 343.950 ;
        RECT 767.400 340.050 768.600 364.950 ;
        RECT 757.950 338.400 762.600 340.050 ;
        RECT 757.950 337.950 762.000 338.400 ;
        RECT 766.950 337.950 769.050 340.050 ;
        RECT 748.950 331.950 751.050 334.050 ;
        RECT 749.400 319.050 750.600 331.950 ;
        RECT 779.400 331.050 780.600 370.950 ;
        RECT 788.400 364.050 789.600 379.950 ;
        RECT 793.950 372.600 798.000 373.050 ;
        RECT 793.950 370.950 798.600 372.600 ;
        RECT 784.950 361.950 787.050 364.050 ;
        RECT 788.400 362.400 793.050 364.050 ;
        RECT 789.000 361.950 793.050 362.400 ;
        RECT 785.400 352.050 786.600 361.950 ;
        RECT 797.400 361.050 798.600 370.950 ;
        RECT 796.950 358.950 799.050 361.050 ;
        RECT 784.950 349.950 787.050 352.050 ;
        RECT 793.950 342.600 796.050 343.050 ;
        RECT 788.400 342.000 796.050 342.600 ;
        RECT 787.950 341.400 796.050 342.000 ;
        RECT 787.950 337.950 790.050 341.400 ;
        RECT 793.950 340.950 796.050 341.400 ;
        RECT 799.950 340.950 802.050 343.050 ;
        RECT 790.950 336.600 793.050 337.050 ;
        RECT 800.400 336.600 801.600 340.950 ;
        RECT 790.950 335.400 801.600 336.600 ;
        RECT 790.950 334.950 793.050 335.400 ;
        RECT 803.400 334.050 804.600 388.950 ;
        RECT 809.400 376.050 810.600 394.950 ;
        RECT 815.400 394.050 816.600 409.950 ;
        RECT 827.400 403.050 828.600 416.400 ;
        RECT 833.400 412.050 834.600 418.950 ;
        RECT 832.950 409.950 835.050 412.050 ;
        RECT 826.950 400.950 829.050 403.050 ;
        RECT 814.950 391.950 817.050 394.050 ;
        RECT 836.400 391.050 837.600 472.950 ;
        RECT 842.400 399.600 843.600 514.950 ;
        RECT 845.400 463.050 846.600 538.950 ;
        RECT 851.400 537.600 852.600 592.950 ;
        RECT 857.400 583.050 858.600 620.400 ;
        RECT 860.400 595.050 861.600 622.950 ;
        RECT 874.950 613.950 877.050 616.050 ;
        RECT 875.400 610.050 876.600 613.950 ;
        RECT 881.400 610.050 882.600 625.950 ;
        RECT 890.400 612.600 891.600 649.950 ;
        RECT 896.400 643.050 897.600 655.950 ;
        RECT 892.950 641.400 897.600 643.050 ;
        RECT 892.950 640.950 897.000 641.400 ;
        RECT 895.950 622.950 898.050 625.050 ;
        RECT 887.400 611.400 891.600 612.600 ;
        RECT 874.950 607.950 877.050 610.050 ;
        RECT 880.950 607.950 883.050 610.050 ;
        RECT 883.950 607.950 886.050 610.050 ;
        RECT 884.400 604.050 885.600 607.950 ;
        RECT 883.950 601.950 886.050 604.050 ;
        RECT 869.100 598.950 871.200 601.050 ;
        RECT 877.950 600.600 880.050 601.050 ;
        RECT 877.950 599.400 885.600 600.600 ;
        RECT 877.950 598.950 880.050 599.400 ;
        RECT 859.950 592.950 862.050 595.050 ;
        RECT 856.950 580.950 859.050 583.050 ;
        RECT 869.400 574.050 870.600 598.950 ;
        RECT 884.400 597.600 885.600 599.400 ;
        RECT 887.400 598.050 888.600 611.400 ;
        RECT 891.000 609.600 895.050 610.050 ;
        RECT 890.400 607.950 895.050 609.600 ;
        RECT 890.400 604.050 891.600 607.950 ;
        RECT 896.400 606.600 897.600 622.950 ;
        RECT 899.400 622.050 900.600 670.950 ;
        RECT 904.950 667.950 907.050 670.050 ;
        RECT 901.950 649.950 904.050 652.050 ;
        RECT 902.400 625.050 903.600 649.950 ;
        RECT 901.950 622.950 904.050 625.050 ;
        RECT 905.400 622.200 906.600 667.950 ;
        RECT 898.950 619.950 901.050 622.050 ;
        RECT 904.950 620.100 907.050 622.200 ;
        RECT 904.950 616.800 907.050 618.900 ;
        RECT 898.950 613.950 901.050 616.050 ;
        RECT 899.400 610.050 900.600 613.950 ;
        RECT 898.950 607.950 901.050 610.050 ;
        RECT 896.400 605.400 900.600 606.600 ;
        RECT 889.950 601.950 892.050 604.050 ;
        RECT 894.000 600.600 898.050 601.050 ;
        RECT 893.400 600.000 898.050 600.600 ;
        RECT 892.950 598.950 898.050 600.000 ;
        RECT 886.950 597.600 889.050 598.050 ;
        RECT 884.400 596.400 889.050 597.600 ;
        RECT 886.950 595.950 889.050 596.400 ;
        RECT 892.950 595.950 895.050 598.950 ;
        RECT 880.950 592.950 883.050 595.050 ;
        RECT 881.400 574.050 882.600 592.950 ;
        RECT 889.950 589.950 892.050 592.050 ;
        RECT 868.950 571.950 871.050 574.050 ;
        RECT 880.950 571.950 883.050 574.050 ;
        RECT 886.950 571.950 889.050 574.050 ;
        RECT 859.950 562.950 862.050 565.050 ;
        RECT 865.950 562.950 868.050 565.050 ;
        RECT 860.400 559.050 861.600 562.950 ;
        RECT 866.400 559.050 867.600 562.950 ;
        RECT 859.950 556.950 862.050 559.050 ;
        RECT 865.950 556.950 868.050 559.050 ;
        RECT 862.950 553.950 865.050 556.050 ;
        RECT 848.400 536.400 852.600 537.600 ;
        RECT 848.400 517.050 849.600 536.400 ;
        RECT 863.400 532.050 864.600 553.950 ;
        RECT 869.400 538.050 870.600 571.950 ;
        RECT 874.950 553.950 877.050 556.050 ;
        RECT 868.950 535.950 871.050 538.050 ;
        RECT 875.400 532.050 876.600 553.950 ;
        RECT 881.400 541.200 882.600 571.950 ;
        RECT 887.400 550.050 888.600 571.950 ;
        RECT 886.950 547.950 889.050 550.050 ;
        RECT 880.950 539.100 883.050 541.200 ;
        RECT 886.950 538.950 889.050 541.050 ;
        RECT 880.950 535.800 883.050 537.900 ;
        RECT 881.400 532.050 882.600 535.800 ;
        RECT 850.950 531.600 853.050 532.050 ;
        RECT 856.950 531.600 859.050 532.050 ;
        RECT 850.950 530.400 859.050 531.600 ;
        RECT 850.950 529.950 853.050 530.400 ;
        RECT 856.950 529.950 859.050 530.400 ;
        RECT 862.950 529.950 865.050 532.050 ;
        RECT 874.950 529.950 877.050 532.050 ;
        RECT 880.950 529.950 883.050 532.050 ;
        RECT 859.950 522.600 862.050 523.050 ;
        RECT 865.950 522.600 868.050 523.050 ;
        RECT 859.950 521.400 868.050 522.600 ;
        RECT 859.950 520.950 862.050 521.400 ;
        RECT 865.950 520.950 868.050 521.400 ;
        RECT 877.950 522.600 880.050 523.050 ;
        RECT 887.400 522.600 888.600 538.950 ;
        RECT 890.400 532.050 891.600 589.950 ;
        RECT 899.400 586.050 900.600 605.400 ;
        RECT 898.950 583.950 901.050 586.050 ;
        RECT 892.950 577.950 895.050 580.050 ;
        RECT 893.400 538.050 894.600 577.950 ;
        RECT 892.950 535.950 895.050 538.050 ;
        RECT 898.950 535.950 901.050 538.050 ;
        RECT 889.950 529.950 892.050 532.050 ;
        RECT 877.950 521.400 888.600 522.600 ;
        RECT 877.950 520.950 880.050 521.400 ;
        RECT 853.950 517.950 856.050 520.050 ;
        RECT 847.950 514.950 850.050 517.050 ;
        RECT 854.400 502.050 855.600 517.950 ;
        RECT 883.950 516.600 886.050 520.050 ;
        RECT 883.950 516.000 888.600 516.600 ;
        RECT 884.400 515.400 888.600 516.000 ;
        RECT 880.950 511.950 883.050 514.050 ;
        RECT 853.950 499.950 856.050 502.050 ;
        RECT 877.950 499.950 880.050 502.050 ;
        RECT 878.400 496.050 879.600 499.950 ;
        RECT 847.950 493.950 850.050 496.050 ;
        RECT 866.100 493.950 868.200 496.050 ;
        RECT 877.950 493.950 880.050 496.050 ;
        RECT 848.400 489.600 849.600 493.950 ;
        RECT 848.400 489.000 852.600 489.600 ;
        RECT 848.400 488.400 853.050 489.000 ;
        RECT 850.950 484.950 853.050 488.400 ;
        RECT 856.950 484.950 859.050 487.050 ;
        RECT 857.400 481.050 858.600 484.950 ;
        RECT 856.950 478.950 859.050 481.050 ;
        RECT 847.950 463.950 850.050 466.050 ;
        RECT 844.950 460.950 847.050 463.050 ;
        RECT 848.400 454.050 849.600 463.950 ;
        RECT 859.950 460.950 862.050 463.050 ;
        RECT 853.950 457.950 856.050 460.050 ;
        RECT 848.400 452.400 853.050 454.050 ;
        RECT 849.000 451.950 853.050 452.400 ;
        RECT 844.950 424.950 847.050 427.050 ;
        RECT 845.400 421.050 846.600 424.950 ;
        RECT 854.400 421.050 855.600 457.950 ;
        RECT 860.400 454.050 861.600 460.950 ;
        RECT 866.400 460.050 867.600 493.950 ;
        RECT 881.400 487.050 882.600 511.950 ;
        RECT 887.400 510.600 888.600 515.400 ;
        RECT 884.400 509.400 888.600 510.600 ;
        RECT 884.400 492.600 885.600 509.400 ;
        RECT 884.400 491.400 888.600 492.600 ;
        RECT 874.950 484.950 877.050 487.050 ;
        RECT 880.950 484.950 883.050 487.050 ;
        RECT 875.400 481.050 876.600 484.950 ;
        RECT 874.950 478.950 877.050 481.050 ;
        RECT 874.950 463.950 877.050 466.050 ;
        RECT 887.400 465.600 888.600 491.400 ;
        RECT 884.400 464.400 888.600 465.600 ;
        RECT 865.950 457.950 868.050 460.050 ;
        RECT 856.950 452.400 861.600 454.050 ;
        RECT 865.950 453.600 868.050 454.050 ;
        RECT 871.950 453.600 874.050 454.050 ;
        RECT 865.950 452.400 874.050 453.600 ;
        RECT 856.950 451.950 861.000 452.400 ;
        RECT 865.950 451.950 868.050 452.400 ;
        RECT 871.950 451.950 874.050 452.400 ;
        RECT 875.400 445.050 876.600 463.950 ;
        RECT 874.950 442.950 877.050 445.050 ;
        RECT 859.950 427.950 862.050 430.050 ;
        RECT 844.950 418.950 847.050 421.050 ;
        RECT 850.950 419.400 855.600 421.050 ;
        RECT 850.950 418.950 855.000 419.400 ;
        RECT 845.400 406.050 846.600 418.950 ;
        RECT 844.950 403.950 847.050 406.050 ;
        RECT 842.400 398.400 846.600 399.600 ;
        RECT 835.950 388.950 838.050 391.050 ;
        RECT 845.400 388.050 846.600 398.400 ;
        RECT 844.950 385.950 847.050 388.050 ;
        RECT 814.950 379.950 817.050 382.050 ;
        RECT 815.400 376.050 816.600 379.950 ;
        RECT 860.400 376.050 861.600 427.950 ;
        RECT 884.400 427.050 885.600 464.400 ;
        RECT 890.400 462.600 891.600 529.950 ;
        RECT 899.400 523.050 900.600 535.950 ;
        RECT 898.950 520.950 901.050 523.050 ;
        RECT 892.950 511.950 895.050 514.050 ;
        RECT 893.400 487.050 894.600 511.950 ;
        RECT 899.400 505.050 900.600 520.950 ;
        RECT 905.400 508.200 906.600 616.800 ;
        RECT 904.950 506.100 907.050 508.200 ;
        RECT 898.950 502.950 901.050 505.050 ;
        RECT 904.950 502.800 907.050 504.900 ;
        RECT 895.950 499.950 898.050 502.050 ;
        RECT 896.400 487.050 897.600 499.950 ;
        RECT 892.950 484.950 895.050 487.050 ;
        RECT 896.400 485.400 901.050 487.050 ;
        RECT 897.000 484.950 901.050 485.400 ;
        RECT 887.400 461.400 891.600 462.600 ;
        RECT 874.950 424.950 877.050 427.050 ;
        RECT 883.950 424.950 886.050 427.050 ;
        RECT 875.400 418.050 876.600 424.950 ;
        RECT 871.950 416.400 876.600 418.050 ;
        RECT 871.950 415.950 876.000 416.400 ;
        RECT 877.950 409.950 880.050 412.050 ;
        RECT 883.950 409.950 886.050 412.050 ;
        RECT 878.400 406.050 879.600 409.950 ;
        RECT 877.950 403.950 880.050 406.050 ;
        RECT 884.400 403.050 885.600 409.950 ;
        RECT 883.950 400.950 886.050 403.050 ;
        RECT 808.950 373.950 811.050 376.050 ;
        RECT 814.950 373.950 817.050 376.050 ;
        RECT 841.950 373.950 844.050 376.050 ;
        RECT 856.950 373.950 859.050 376.050 ;
        RECT 860.400 373.950 865.050 376.050 ;
        RECT 820.950 370.950 823.050 373.050 ;
        RECT 821.400 361.050 822.600 370.950 ;
        RECT 829.950 364.950 832.050 367.050 ;
        RECT 838.950 364.950 841.050 367.050 ;
        RECT 830.400 361.050 831.600 364.950 ;
        RECT 839.400 361.050 840.600 364.950 ;
        RECT 842.400 361.050 843.600 373.950 ;
        RECT 847.950 366.600 850.050 367.050 ;
        RECT 853.950 366.600 856.050 367.050 ;
        RECT 847.950 365.400 856.050 366.600 ;
        RECT 847.950 364.950 850.050 365.400 ;
        RECT 853.950 364.950 856.050 365.400 ;
        RECT 857.400 361.050 858.600 373.950 ;
        RECT 820.950 358.950 823.050 361.050 ;
        RECT 829.950 358.950 832.050 361.050 ;
        RECT 838.800 358.950 840.900 361.050 ;
        RECT 842.100 358.950 844.200 361.050 ;
        RECT 856.950 358.950 859.050 361.050 ;
        RECT 823.950 357.600 828.000 358.050 ;
        RECT 823.950 355.950 828.600 357.600 ;
        RECT 811.950 343.950 814.050 346.050 ;
        RECT 812.400 340.050 813.600 343.950 ;
        RECT 811.950 337.950 814.050 340.050 ;
        RECT 802.950 331.950 805.050 334.050 ;
        RECT 778.950 328.950 781.050 331.050 ;
        RECT 814.950 328.950 817.050 331.050 ;
        RECT 815.400 325.050 816.600 328.950 ;
        RECT 802.950 322.950 805.050 325.050 ;
        RECT 808.950 322.950 811.050 325.050 ;
        RECT 814.950 322.950 817.050 325.050 ;
        RECT 748.950 316.950 751.050 319.050 ;
        RECT 778.950 316.950 781.050 319.050 ;
        RECT 730.950 313.950 733.050 316.050 ;
        RECT 739.950 313.950 742.050 316.050 ;
        RECT 724.950 295.950 727.050 298.050 ;
        RECT 730.950 295.950 733.050 298.050 ;
        RECT 721.950 286.950 724.050 289.050 ;
        RECT 731.400 277.050 732.600 295.950 ;
        RECT 740.400 295.050 741.600 313.950 ;
        RECT 739.950 292.950 742.050 295.050 ;
        RECT 748.950 292.950 751.050 295.050 ;
        RECT 730.950 274.950 733.050 277.050 ;
        RECT 742.950 274.950 745.050 277.050 ;
        RECT 700.950 265.950 703.050 268.050 ;
        RECT 701.400 262.050 702.600 265.950 ;
        RECT 700.950 259.950 703.050 262.050 ;
        RECT 715.950 259.950 718.050 262.050 ;
        RECT 688.950 250.950 691.050 253.050 ;
        RECT 697.950 250.950 700.050 253.050 ;
        RECT 703.950 250.950 706.050 253.050 ;
        RECT 709.950 252.600 712.050 253.050 ;
        RECT 716.400 252.600 717.600 259.950 ;
        RECT 743.400 253.050 744.600 274.950 ;
        RECT 749.400 268.050 750.600 292.950 ;
        RECT 766.950 286.950 769.050 289.050 ;
        RECT 767.400 277.050 768.600 286.950 ;
        RECT 779.400 283.050 780.600 316.950 ;
        RECT 784.950 307.950 787.050 310.050 ;
        RECT 785.400 298.050 786.600 307.950 ;
        RECT 790.950 301.950 793.050 304.050 ;
        RECT 791.400 298.050 792.600 301.950 ;
        RECT 784.950 295.950 787.050 298.050 ;
        RECT 790.950 295.950 793.050 298.050 ;
        RECT 787.950 286.950 790.050 289.050 ;
        RECT 793.950 286.950 796.050 289.050 ;
        RECT 788.400 283.050 789.600 286.950 ;
        RECT 778.950 280.950 781.050 283.050 ;
        RECT 787.950 280.950 790.050 283.050 ;
        RECT 766.950 276.600 769.050 277.050 ;
        RECT 766.950 275.400 771.600 276.600 ;
        RECT 766.950 274.950 769.050 275.400 ;
        RECT 748.950 265.950 751.050 268.050 ;
        RECT 763.950 259.950 766.050 262.050 ;
        RECT 709.950 251.400 717.600 252.600 ;
        RECT 709.950 250.950 712.050 251.400 ;
        RECT 727.950 250.950 730.050 253.050 ;
        RECT 742.950 250.950 745.050 253.050 ;
        RECT 748.950 250.950 751.050 253.050 ;
        RECT 754.950 250.950 757.050 253.050 ;
        RECT 688.950 232.950 691.050 235.050 ;
        RECT 679.950 220.950 682.050 223.050 ;
        RECT 680.400 208.050 681.600 220.950 ;
        RECT 689.400 208.050 690.600 232.950 ;
        RECT 698.400 223.050 699.600 250.950 ;
        RECT 704.400 232.050 705.600 250.950 ;
        RECT 712.950 244.950 715.050 247.050 ;
        RECT 703.950 229.950 706.050 232.050 ;
        RECT 697.950 220.950 700.050 223.050 ;
        RECT 703.950 220.950 706.050 223.050 ;
        RECT 697.950 214.950 700.050 217.050 ;
        RECT 680.400 206.400 685.050 208.050 ;
        RECT 681.000 205.950 685.050 206.400 ;
        RECT 688.950 205.950 691.050 208.050 ;
        RECT 679.950 199.950 682.050 202.050 ;
        RECT 680.400 187.050 681.600 199.950 ;
        RECT 698.400 193.050 699.600 214.950 ;
        RECT 704.400 208.050 705.600 220.950 ;
        RECT 703.950 205.950 706.050 208.050 ;
        RECT 685.950 190.950 688.050 193.050 ;
        RECT 697.950 190.950 700.050 193.050 ;
        RECT 703.950 190.950 706.050 193.050 ;
        RECT 686.400 187.050 687.600 190.950 ;
        RECT 704.400 187.050 705.600 190.950 ;
        RECT 679.950 184.950 682.050 187.050 ;
        RECT 685.950 184.950 688.050 187.050 ;
        RECT 703.950 184.950 706.050 187.050 ;
        RECT 708.000 186.600 712.050 187.050 ;
        RECT 707.400 184.950 712.050 186.600 ;
        RECT 673.950 181.950 676.050 184.050 ;
        RECT 707.400 183.600 708.600 184.950 ;
        RECT 701.400 182.400 708.600 183.600 ;
        RECT 674.400 172.050 675.600 181.950 ;
        RECT 701.400 178.050 702.600 182.400 ;
        RECT 700.950 175.950 703.050 178.050 ;
        RECT 709.950 175.950 712.050 178.050 ;
        RECT 673.950 169.950 676.050 172.050 ;
        RECT 685.950 157.950 688.050 160.050 ;
        RECT 676.950 154.950 679.050 157.050 ;
        RECT 677.400 139.050 678.600 154.950 ;
        RECT 686.400 139.050 687.600 157.950 ;
        RECT 703.950 148.950 706.050 151.050 ;
        RECT 704.400 142.050 705.600 148.950 ;
        RECT 710.400 142.050 711.600 175.950 ;
        RECT 713.400 151.050 714.600 244.950 ;
        RECT 728.400 232.050 729.600 250.950 ;
        RECT 749.400 244.050 750.600 250.950 ;
        RECT 748.950 241.950 751.050 244.050 ;
        RECT 755.400 241.050 756.600 250.950 ;
        RECT 764.400 244.050 765.600 259.950 ;
        RECT 770.400 253.050 771.600 275.400 ;
        RECT 794.400 274.050 795.600 286.950 ;
        RECT 803.400 280.050 804.600 322.950 ;
        RECT 809.400 304.050 810.600 322.950 ;
        RECT 820.950 313.950 823.050 316.050 ;
        RECT 814.950 307.950 817.050 310.050 ;
        RECT 808.950 301.950 811.050 304.050 ;
        RECT 809.400 291.600 810.600 301.950 ;
        RECT 815.400 295.050 816.600 307.950 ;
        RECT 821.400 295.050 822.600 313.950 ;
        RECT 827.400 310.050 828.600 355.950 ;
        RECT 832.950 349.950 835.050 352.050 ;
        RECT 833.400 331.050 834.600 349.950 ;
        RECT 839.400 331.050 840.600 358.950 ;
        RECT 857.400 355.050 858.600 358.950 ;
        RECT 856.950 352.950 859.050 355.050 ;
        RECT 860.400 346.050 861.600 373.950 ;
        RECT 871.950 370.950 874.050 373.050 ;
        RECT 879.000 372.600 883.050 373.050 ;
        RECT 878.400 370.950 883.050 372.600 ;
        RECT 862.950 364.950 865.050 367.050 ;
        RECT 863.400 349.050 864.600 364.950 ;
        RECT 872.400 355.050 873.600 370.950 ;
        RECT 865.950 352.950 868.050 355.050 ;
        RECT 871.950 352.950 874.050 355.050 ;
        RECT 862.950 346.950 865.050 349.050 ;
        RECT 859.950 343.950 862.050 346.050 ;
        RECT 844.950 339.600 847.050 340.050 ;
        RECT 850.950 339.600 853.050 340.050 ;
        RECT 844.950 338.400 853.050 339.600 ;
        RECT 844.950 337.950 847.050 338.400 ;
        RECT 850.950 337.950 853.050 338.400 ;
        RECT 832.950 328.950 835.050 331.050 ;
        RECT 838.950 328.950 841.050 331.050 ;
        RECT 866.400 316.050 867.600 352.950 ;
        RECT 871.950 346.950 874.050 349.050 ;
        RECT 872.400 340.050 873.600 346.950 ;
        RECT 878.400 343.050 879.600 370.950 ;
        RECT 887.400 346.050 888.600 461.400 ;
        RECT 889.950 457.950 892.050 460.050 ;
        RECT 901.950 457.950 904.050 460.050 ;
        RECT 890.400 451.050 891.600 457.950 ;
        RECT 902.400 454.050 903.600 457.950 ;
        RECT 894.000 453.600 898.050 454.050 ;
        RECT 893.400 451.950 898.050 453.600 ;
        RECT 901.950 451.950 904.050 454.050 ;
        RECT 889.950 448.950 892.050 451.050 ;
        RECT 893.400 439.050 894.600 451.950 ;
        RECT 892.950 436.950 895.050 439.050 ;
        RECT 895.950 433.950 898.050 436.050 ;
        RECT 889.950 424.950 892.050 427.050 ;
        RECT 890.400 421.050 891.600 424.950 ;
        RECT 896.400 421.050 897.600 433.950 ;
        RECT 889.950 418.950 892.050 421.050 ;
        RECT 895.950 418.950 898.050 421.050 ;
        RECT 896.400 406.050 897.600 418.950 ;
        RECT 895.950 403.950 898.050 406.050 ;
        RECT 898.950 364.950 901.050 367.050 ;
        RECT 880.950 343.950 883.050 346.050 ;
        RECT 886.950 343.950 889.050 346.050 ;
        RECT 892.950 343.950 895.050 346.050 ;
        RECT 877.950 340.950 880.050 343.050 ;
        RECT 871.950 337.950 874.050 340.050 ;
        RECT 881.400 331.050 882.600 343.950 ;
        RECT 883.950 339.600 888.000 340.050 ;
        RECT 883.950 337.950 888.600 339.600 ;
        RECT 887.400 331.050 888.600 337.950 ;
        RECT 868.950 330.600 871.050 331.050 ;
        RECT 874.950 330.600 877.050 331.050 ;
        RECT 868.950 329.400 877.050 330.600 ;
        RECT 868.950 328.950 871.050 329.400 ;
        RECT 874.950 328.950 877.050 329.400 ;
        RECT 880.950 328.950 883.050 331.050 ;
        RECT 886.950 328.950 889.050 331.050 ;
        RECT 881.400 325.050 882.600 328.950 ;
        RECT 880.950 322.950 883.050 325.050 ;
        RECT 880.950 316.950 883.050 319.050 ;
        RECT 865.950 313.950 868.050 316.050 ;
        RECT 871.950 313.950 874.050 316.050 ;
        RECT 826.950 307.950 829.050 310.050 ;
        RECT 872.400 295.050 873.600 313.950 ;
        RECT 814.950 292.950 817.050 295.050 ;
        RECT 820.950 292.950 823.050 295.050 ;
        RECT 829.950 292.950 832.050 295.050 ;
        RECT 871.950 292.950 874.050 295.050 ;
        RECT 809.400 290.400 816.600 291.600 ;
        RECT 815.400 286.050 816.600 290.400 ;
        RECT 808.950 283.950 811.050 286.050 ;
        RECT 814.950 283.950 817.050 286.050 ;
        RECT 809.400 280.050 810.600 283.950 ;
        RECT 802.950 277.950 805.050 280.050 ;
        RECT 808.950 277.950 811.050 280.050 ;
        RECT 793.950 271.950 796.050 274.050 ;
        RECT 823.950 271.950 826.050 274.050 ;
        RECT 793.950 265.950 796.050 268.050 ;
        RECT 817.950 265.950 820.050 268.050 ;
        RECT 794.400 262.050 795.600 265.950 ;
        RECT 818.400 262.050 819.600 265.950 ;
        RECT 824.400 262.050 825.600 271.950 ;
        RECT 830.400 268.050 831.600 292.950 ;
        RECT 847.950 286.950 850.050 289.050 ;
        RECT 848.400 277.050 849.600 286.950 ;
        RECT 841.950 274.950 844.050 277.050 ;
        RECT 847.950 274.950 850.050 277.050 ;
        RECT 868.950 274.950 871.050 277.050 ;
        RECT 829.950 265.950 832.050 268.050 ;
        RECT 842.400 262.050 843.600 274.950 ;
        RECT 859.950 268.950 862.050 271.050 ;
        RECT 860.400 265.050 861.600 268.950 ;
        RECT 869.400 265.050 870.600 274.950 ;
        RECT 881.400 265.050 882.600 316.950 ;
        RECT 887.400 271.050 888.600 328.950 ;
        RECT 893.400 327.600 894.600 343.950 ;
        RECT 899.400 340.050 900.600 364.950 ;
        RECT 898.950 337.950 901.050 340.050 ;
        RECT 890.400 326.400 894.600 327.600 ;
        RECT 886.950 268.950 889.050 271.050 ;
        RECT 859.950 262.950 862.050 265.050 ;
        RECT 868.950 262.950 871.050 265.050 ;
        RECT 880.950 262.950 883.050 265.050 ;
        RECT 781.950 259.950 784.050 262.050 ;
        RECT 769.950 250.950 772.050 253.050 ;
        RECT 775.950 250.950 778.050 253.050 ;
        RECT 763.950 241.950 766.050 244.050 ;
        RECT 776.400 241.050 777.600 250.950 ;
        RECT 782.400 247.050 783.600 259.950 ;
        RECT 787.950 258.600 790.050 262.050 ;
        RECT 793.950 259.950 796.050 262.050 ;
        RECT 817.950 259.950 820.050 262.050 ;
        RECT 823.950 259.950 826.050 262.050 ;
        RECT 841.950 259.950 844.050 262.050 ;
        RECT 785.400 258.000 790.050 258.600 ;
        RECT 785.400 257.400 789.600 258.000 ;
        RECT 785.400 253.050 786.600 257.400 ;
        RECT 865.950 253.950 868.050 256.050 ;
        RECT 871.950 253.950 874.050 256.050 ;
        RECT 784.950 250.950 787.050 253.050 ;
        RECT 790.950 250.950 793.050 253.050 ;
        RECT 796.950 250.950 799.050 253.050 ;
        RECT 814.950 250.950 817.050 253.050 ;
        RECT 820.950 252.600 823.050 253.050 ;
        RECT 826.950 252.600 829.050 253.050 ;
        RECT 820.950 251.400 829.050 252.600 ;
        RECT 820.950 250.950 823.050 251.400 ;
        RECT 826.950 250.950 829.050 251.400 ;
        RECT 838.950 250.950 841.050 253.050 ;
        RECT 781.950 244.950 784.050 247.050 ;
        RECT 754.950 238.950 757.050 241.050 ;
        RECT 775.950 238.950 778.050 241.050 ;
        RECT 721.950 229.950 724.050 232.050 ;
        RECT 727.950 229.950 730.050 232.050 ;
        RECT 742.950 229.950 745.050 232.050 ;
        RECT 715.950 226.950 718.050 229.050 ;
        RECT 716.400 211.050 717.600 226.950 ;
        RECT 722.400 220.050 723.600 229.950 ;
        RECT 743.400 220.050 744.600 229.950 ;
        RECT 755.400 229.050 756.600 238.950 ;
        RECT 784.950 235.950 787.050 238.050 ;
        RECT 760.950 229.950 763.050 232.050 ;
        RECT 754.950 226.950 757.050 229.050 ;
        RECT 721.950 217.950 724.050 220.050 ;
        RECT 727.950 219.600 732.000 220.050 ;
        RECT 727.950 217.950 732.600 219.600 ;
        RECT 743.400 218.400 748.050 220.050 ;
        RECT 744.000 217.950 748.050 218.400 ;
        RECT 731.400 211.050 732.600 217.950 ;
        RECT 716.400 209.400 721.050 211.050 ;
        RECT 717.000 208.950 721.050 209.400 ;
        RECT 730.950 208.950 733.050 211.050 ;
        RECT 724.950 205.950 727.050 208.050 ;
        RECT 725.400 202.050 726.600 205.950 ;
        RECT 724.950 199.950 727.050 202.050 ;
        RECT 721.950 190.950 724.050 193.050 ;
        RECT 751.950 190.950 754.050 193.050 ;
        RECT 722.400 178.050 723.600 190.950 ;
        RECT 727.950 187.950 730.050 190.050 ;
        RECT 728.400 184.050 729.600 187.950 ;
        RECT 752.400 184.050 753.600 190.950 ;
        RECT 761.400 190.050 762.600 229.950 ;
        RECT 763.950 226.950 766.050 229.050 ;
        RECT 764.400 220.050 765.600 226.950 ;
        RECT 769.950 223.950 772.050 226.050 ;
        RECT 770.400 220.050 771.600 223.950 ;
        RECT 763.950 217.950 766.050 220.050 ;
        RECT 769.950 217.950 772.050 220.050 ;
        RECT 775.950 217.950 778.050 220.050 ;
        RECT 764.400 199.050 765.600 217.950 ;
        RECT 776.400 211.050 777.600 217.950 ;
        RECT 772.950 208.950 775.050 211.050 ;
        RECT 776.400 209.400 781.050 211.050 ;
        RECT 777.000 208.950 781.050 209.400 ;
        RECT 773.400 201.600 774.600 208.950 ;
        RECT 773.400 200.400 777.600 201.600 ;
        RECT 763.950 196.950 766.050 199.050 ;
        RECT 772.950 196.950 775.050 199.050 ;
        RECT 760.950 187.950 763.050 190.050 ;
        RECT 769.950 187.950 772.050 190.050 ;
        RECT 770.400 184.050 771.600 187.950 ;
        RECT 727.950 181.950 730.050 184.050 ;
        RECT 751.950 181.950 754.050 184.050 ;
        RECT 769.950 181.950 772.050 184.050 ;
        RECT 773.400 183.600 774.600 196.950 ;
        RECT 776.400 190.050 777.600 200.400 ;
        RECT 775.950 187.950 778.050 190.050 ;
        RECT 775.950 183.600 778.050 184.050 ;
        RECT 773.400 182.400 778.050 183.600 ;
        RECT 775.950 181.950 778.050 182.400 ;
        RECT 721.950 175.950 724.050 178.050 ;
        RECT 722.400 172.050 723.600 175.950 ;
        RECT 730.950 172.950 733.050 175.050 ;
        RECT 748.950 172.950 751.050 175.050 ;
        RECT 766.950 172.950 769.050 175.050 ;
        RECT 772.950 172.950 775.050 175.050 ;
        RECT 721.950 169.950 724.050 172.050 ;
        RECT 731.400 154.050 732.600 172.950 ;
        RECT 749.400 163.050 750.600 172.950 ;
        RECT 767.400 169.050 768.600 172.950 ;
        RECT 766.950 166.950 769.050 169.050 ;
        RECT 773.400 163.050 774.600 172.950 ;
        RECT 736.950 160.950 739.050 163.050 ;
        RECT 748.950 160.950 751.050 163.050 ;
        RECT 772.950 160.950 775.050 163.050 ;
        RECT 724.950 151.950 727.050 154.050 ;
        RECT 730.950 151.950 733.050 154.050 ;
        RECT 712.950 148.950 715.050 151.050 ;
        RECT 725.400 142.050 726.600 151.950 ;
        RECT 730.950 145.950 733.050 148.050 ;
        RECT 731.400 142.050 732.600 145.950 ;
        RECT 703.950 139.950 706.050 142.050 ;
        RECT 709.950 139.950 712.050 142.050 ;
        RECT 718.950 139.950 721.050 142.050 ;
        RECT 724.950 139.950 727.050 142.050 ;
        RECT 730.950 139.950 733.050 142.050 ;
        RECT 676.950 136.950 679.050 139.050 ;
        RECT 685.950 136.950 688.050 139.050 ;
        RECT 608.100 112.950 610.200 115.050 ;
        RECT 616.950 112.950 619.050 115.050 ;
        RECT 651.000 114.600 655.050 115.050 ;
        RECT 650.400 112.950 655.050 114.600 ;
        RECT 670.950 112.950 673.050 115.050 ;
        RECT 617.400 109.050 618.600 112.950 ;
        RECT 625.950 109.950 628.050 112.050 ;
        RECT 643.950 109.950 646.050 112.050 ;
        RECT 610.950 108.600 613.050 109.050 ;
        RECT 602.400 107.400 613.050 108.600 ;
        RECT 610.950 106.950 613.050 107.400 ;
        RECT 616.950 106.950 619.050 109.050 ;
        RECT 565.950 103.950 568.050 106.050 ;
        RECT 580.950 103.950 583.050 106.050 ;
        RECT 586.950 105.600 589.050 106.050 ;
        RECT 595.950 105.600 598.050 106.050 ;
        RECT 586.950 104.400 598.050 105.600 ;
        RECT 586.950 103.950 589.050 104.400 ;
        RECT 595.950 103.950 598.050 104.400 ;
        RECT 626.400 100.050 627.600 109.950 ;
        RECT 634.950 103.950 637.050 106.050 ;
        RECT 568.950 99.600 571.050 100.050 ;
        RECT 563.400 98.400 571.050 99.600 ;
        RECT 552.000 96.600 556.050 97.050 ;
        RECT 551.400 96.000 556.050 96.600 ;
        RECT 550.950 94.950 556.050 96.000 ;
        RECT 559.950 96.600 564.000 97.050 ;
        RECT 559.950 94.950 564.600 96.600 ;
        RECT 526.950 91.950 529.050 94.050 ;
        RECT 544.950 91.950 547.050 94.050 ;
        RECT 550.950 91.950 553.050 94.950 ;
        RECT 541.950 82.950 544.050 85.050 ;
        RECT 556.950 82.950 559.050 85.050 ;
        RECT 520.950 61.950 523.050 64.050 ;
        RECT 542.400 52.050 543.600 82.950 ;
        RECT 550.950 70.950 553.050 73.050 ;
        RECT 541.950 49.950 544.050 52.050 ;
        RECT 535.950 46.950 538.050 49.050 ;
        RECT 520.950 43.950 523.050 46.050 ;
        RECT 499.950 40.950 502.050 43.050 ;
        RECT 481.950 28.950 484.050 31.050 ;
        RECT 487.950 28.950 490.050 31.050 ;
        RECT 467.400 26.400 471.600 27.600 ;
        RECT 467.400 22.050 468.600 26.400 ;
        RECT 482.400 24.600 483.600 28.950 ;
        RECT 508.950 27.600 511.050 28.050 ;
        RECT 514.950 27.600 517.050 28.050 ;
        RECT 508.950 26.400 517.050 27.600 ;
        RECT 508.950 25.950 511.050 26.400 ;
        RECT 514.950 25.950 517.050 26.400 ;
        RECT 473.400 24.000 483.600 24.600 ;
        RECT 472.950 23.400 483.600 24.000 ;
        RECT 454.950 19.950 457.050 22.050 ;
        RECT 466.950 19.950 469.050 22.050 ;
        RECT 472.950 19.950 475.050 23.400 ;
        RECT 481.950 21.600 484.050 22.050 ;
        RECT 476.400 20.400 484.050 21.600 ;
        RECT 455.400 13.050 456.600 19.950 ;
        RECT 460.950 18.600 463.050 19.050 ;
        RECT 476.400 18.600 477.600 20.400 ;
        RECT 481.950 19.950 484.050 20.400 ;
        RECT 521.400 19.050 522.600 43.950 ;
        RECT 536.400 34.050 537.600 46.950 ;
        RECT 551.400 43.050 552.600 70.950 ;
        RECT 557.400 64.050 558.600 82.950 ;
        RECT 563.400 79.050 564.600 94.950 ;
        RECT 562.950 76.950 565.050 79.050 ;
        RECT 556.950 61.950 559.050 64.050 ;
        RECT 566.400 61.050 567.600 98.400 ;
        RECT 568.950 97.950 571.050 98.400 ;
        RECT 577.950 97.950 580.050 100.050 ;
        RECT 625.950 97.950 628.050 100.050 ;
        RECT 578.400 76.050 579.600 97.950 ;
        RECT 622.950 94.950 625.050 97.050 ;
        RECT 616.950 85.950 619.050 88.050 ;
        RECT 584.400 80.400 606.600 81.600 ;
        RECT 577.950 73.950 580.050 76.050 ;
        RECT 584.400 73.050 585.600 80.400 ;
        RECT 601.950 76.950 604.050 79.050 ;
        RECT 592.950 73.950 595.050 76.050 ;
        RECT 583.950 70.950 586.050 73.050 ;
        RECT 562.950 58.950 565.050 61.050 ;
        RECT 565.950 58.950 568.050 61.050 ;
        RECT 574.950 58.950 577.050 61.050 ;
        RECT 553.950 52.950 556.050 55.050 ;
        RECT 550.950 40.950 553.050 43.050 ;
        RECT 554.400 40.050 555.600 52.950 ;
        RECT 563.400 46.050 564.600 58.950 ;
        RECT 562.950 43.950 565.050 46.050 ;
        RECT 575.400 40.050 576.600 58.950 ;
        RECT 593.400 55.050 594.600 73.950 ;
        RECT 602.400 73.050 603.600 76.950 ;
        RECT 601.950 70.950 604.050 73.050 ;
        RECT 592.950 52.950 595.050 55.050 ;
        RECT 541.950 37.950 544.050 40.050 ;
        RECT 553.950 37.950 556.050 40.050 ;
        RECT 574.950 37.950 577.050 40.050 ;
        RECT 589.950 37.950 592.050 40.050 ;
        RECT 535.950 31.950 538.050 34.050 ;
        RECT 542.400 19.050 543.600 37.950 ;
        RECT 559.950 34.950 562.050 37.050 ;
        RECT 560.400 28.050 561.600 34.950 ;
        RECT 565.950 31.950 568.050 34.050 ;
        RECT 566.400 28.050 567.600 31.950 ;
        RECT 590.400 28.050 591.600 37.950 ;
        RECT 602.400 28.050 603.600 70.950 ;
        RECT 605.400 70.050 606.600 80.400 ;
        RECT 604.950 67.950 607.050 70.050 ;
        RECT 617.400 64.050 618.600 85.950 ;
        RECT 623.400 76.050 624.600 94.950 ;
        RECT 635.400 88.050 636.600 103.950 ;
        RECT 644.400 100.050 645.600 109.950 ;
        RECT 650.400 106.050 651.600 112.950 ;
        RECT 655.950 109.950 658.050 112.050 ;
        RECT 656.400 106.050 657.600 109.950 ;
        RECT 682.950 106.950 685.050 109.050 ;
        RECT 649.950 103.950 652.050 106.050 ;
        RECT 655.950 103.950 658.050 106.050 ;
        RECT 670.950 103.950 673.050 106.050 ;
        RECT 643.950 97.950 646.050 100.050 ;
        RECT 652.950 97.950 655.050 100.050 ;
        RECT 653.400 88.050 654.600 97.950 ;
        RECT 658.950 94.950 661.050 97.050 ;
        RECT 664.950 94.950 667.050 97.050 ;
        RECT 659.400 91.050 660.600 94.950 ;
        RECT 658.950 88.950 661.050 91.050 ;
        RECT 634.950 85.950 637.050 88.050 ;
        RECT 653.100 85.950 655.200 88.050 ;
        RECT 665.400 85.050 666.600 94.950 ;
        RECT 664.950 82.950 667.050 85.050 ;
        RECT 622.950 73.950 625.050 76.050 ;
        RECT 637.950 73.950 640.050 76.050 ;
        RECT 610.950 61.950 613.050 64.050 ;
        RECT 616.950 61.950 619.050 64.050 ;
        RECT 611.400 43.050 612.600 61.950 ;
        RECT 622.950 58.950 625.050 61.050 ;
        RECT 623.400 55.050 624.600 58.950 ;
        RECT 613.950 52.950 616.050 55.050 ;
        RECT 619.950 53.400 624.600 55.050 ;
        RECT 619.950 52.950 624.000 53.400 ;
        RECT 614.400 43.050 615.600 52.950 ;
        RECT 638.400 52.050 639.600 73.950 ;
        RECT 665.400 73.050 666.600 82.950 ;
        RECT 664.950 70.950 667.050 73.050 ;
        RECT 655.950 67.950 658.050 70.050 ;
        RECT 656.400 64.050 657.600 67.950 ;
        RECT 671.400 67.050 672.600 103.950 ;
        RECT 683.400 88.050 684.600 106.950 ;
        RECT 682.950 85.950 685.050 88.050 ;
        RECT 679.950 82.950 682.050 85.050 ;
        RECT 676.950 76.950 679.050 79.050 ;
        RECT 664.950 64.050 667.050 67.050 ;
        RECT 670.950 64.950 673.050 67.050 ;
        RECT 655.950 61.950 658.050 64.050 ;
        RECT 661.950 63.000 667.050 64.050 ;
        RECT 661.950 62.400 666.600 63.000 ;
        RECT 661.950 61.950 666.000 62.400 ;
        RECT 670.950 60.600 673.050 61.050 ;
        RECT 677.400 60.600 678.600 76.950 ;
        RECT 680.400 61.050 681.600 82.950 ;
        RECT 686.400 79.050 687.600 136.950 ;
        RECT 719.400 133.050 720.600 139.950 ;
        RECT 712.950 130.950 715.050 133.050 ;
        RECT 719.400 131.400 724.050 133.050 ;
        RECT 720.000 130.950 724.050 131.400 ;
        RECT 688.950 118.950 691.050 121.050 ;
        RECT 694.950 118.950 697.050 121.050 ;
        RECT 689.400 115.050 690.600 118.950 ;
        RECT 688.950 112.950 691.050 115.050 ;
        RECT 689.400 109.050 690.600 112.950 ;
        RECT 688.950 106.950 691.050 109.050 ;
        RECT 695.400 100.050 696.600 118.950 ;
        RECT 703.950 112.950 706.050 115.050 ;
        RECT 704.400 106.050 705.600 112.950 ;
        RECT 703.950 103.950 706.050 106.050 ;
        RECT 694.950 97.950 697.050 100.050 ;
        RECT 700.950 94.950 703.050 97.050 ;
        RECT 701.400 88.050 702.600 94.950 ;
        RECT 700.950 85.950 703.050 88.050 ;
        RECT 713.400 82.050 714.600 130.950 ;
        RECT 727.950 127.950 730.050 130.050 ;
        RECT 721.950 115.950 724.050 118.050 ;
        RECT 715.950 103.950 718.050 106.050 ;
        RECT 716.400 85.050 717.600 103.950 ;
        RECT 722.400 100.050 723.600 115.950 ;
        RECT 728.400 112.050 729.600 127.950 ;
        RECT 737.400 112.050 738.600 160.950 ;
        RECT 748.950 148.950 751.050 151.050 ;
        RECT 742.950 145.950 745.050 148.050 ;
        RECT 727.950 109.950 730.050 112.050 ;
        RECT 736.950 109.950 739.050 112.050 ;
        RECT 736.950 103.950 739.050 106.050 ;
        RECT 721.950 97.950 724.050 100.050 ;
        RECT 737.400 99.600 738.600 103.950 ;
        RECT 725.400 98.400 738.600 99.600 ;
        RECT 715.950 82.950 718.050 85.050 ;
        RECT 725.400 82.050 726.600 98.400 ;
        RECT 727.950 94.950 730.050 97.050 ;
        RECT 733.950 94.950 736.050 97.050 ;
        RECT 728.400 91.050 729.600 94.950 ;
        RECT 734.400 91.050 735.600 94.950 ;
        RECT 743.400 91.050 744.600 145.950 ;
        RECT 749.400 142.050 750.600 148.950 ;
        RECT 776.400 148.050 777.600 181.950 ;
        RECT 781.950 175.950 784.050 178.050 ;
        RECT 775.950 145.950 778.050 148.050 ;
        RECT 778.950 142.050 781.050 145.050 ;
        RECT 748.950 139.950 751.050 142.050 ;
        RECT 760.950 139.950 763.050 142.050 ;
        RECT 768.000 141.600 772.050 142.050 ;
        RECT 767.400 139.950 772.050 141.600 ;
        RECT 775.950 141.000 781.050 142.050 ;
        RECT 775.950 140.400 780.600 141.000 ;
        RECT 775.950 139.950 780.000 140.400 ;
        RECT 748.950 109.950 751.050 112.050 ;
        RECT 749.400 106.050 750.600 109.950 ;
        RECT 761.400 106.050 762.600 139.950 ;
        RECT 767.400 133.050 768.600 139.950 ;
        RECT 782.400 133.050 783.600 175.950 ;
        RECT 785.400 160.050 786.600 235.950 ;
        RECT 791.400 196.050 792.600 250.950 ;
        RECT 797.400 247.050 798.600 250.950 ;
        RECT 796.950 244.950 799.050 247.050 ;
        RECT 815.400 244.050 816.600 250.950 ;
        RECT 839.400 247.050 840.600 250.950 ;
        RECT 823.950 244.950 826.050 247.050 ;
        RECT 838.950 244.950 841.050 247.050 ;
        RECT 814.950 241.950 817.050 244.050 ;
        RECT 802.950 235.950 805.050 238.050 ;
        RECT 803.400 217.050 804.600 235.950 ;
        RECT 824.400 217.050 825.600 244.950 ;
        RECT 841.950 232.950 844.050 235.050 ;
        RECT 842.400 217.050 843.600 232.950 ;
        RECT 866.400 232.050 867.600 253.950 ;
        RECT 859.950 229.950 862.050 232.050 ;
        RECT 865.950 229.950 868.050 232.050 ;
        RECT 860.400 220.050 861.600 229.950 ;
        RECT 859.950 217.950 862.050 220.050 ;
        RECT 796.950 214.950 799.050 217.050 ;
        RECT 803.400 215.400 808.050 217.050 ;
        RECT 804.000 214.950 808.050 215.400 ;
        RECT 823.950 214.950 826.050 217.050 ;
        RECT 841.950 214.950 844.050 217.050 ;
        RECT 850.950 214.950 853.050 217.050 ;
        RECT 797.400 199.050 798.600 214.950 ;
        RECT 814.950 208.950 817.050 211.050 ;
        RECT 796.950 196.950 799.050 199.050 ;
        RECT 790.950 193.950 793.050 196.050 ;
        RECT 815.400 190.050 816.600 208.950 ;
        RECT 842.400 208.050 843.600 214.950 ;
        RECT 851.400 208.050 852.600 214.950 ;
        RECT 841.950 205.950 844.050 208.050 ;
        RECT 850.950 205.950 853.050 208.050 ;
        RECT 850.950 196.950 853.050 199.050 ;
        RECT 826.950 193.950 829.050 196.050 ;
        RECT 820.950 190.950 823.050 193.050 ;
        RECT 814.950 187.950 817.050 190.050 ;
        RECT 793.950 183.600 796.050 187.050 ;
        RECT 793.950 183.000 798.600 183.600 ;
        RECT 794.400 182.400 798.600 183.000 ;
        RECT 797.400 175.050 798.600 182.400 ;
        RECT 802.950 181.950 805.050 184.050 ;
        RECT 796.950 172.950 799.050 175.050 ;
        RECT 784.950 157.950 787.050 160.050 ;
        RECT 766.950 130.950 769.050 133.050 ;
        RECT 778.950 131.400 783.600 133.050 ;
        RECT 778.950 130.950 783.000 131.400 ;
        RECT 781.950 124.950 784.050 127.050 ;
        RECT 748.950 103.950 751.050 106.050 ;
        RECT 761.400 104.400 766.050 106.050 ;
        RECT 762.000 103.950 766.050 104.400 ;
        RECT 751.950 97.950 754.050 100.050 ;
        RECT 752.400 91.050 753.600 97.950 ;
        RECT 727.950 88.950 730.050 91.050 ;
        RECT 733.950 88.950 736.050 91.050 ;
        RECT 742.950 88.950 745.050 91.050 ;
        RECT 751.950 88.950 754.050 91.050 ;
        RECT 752.400 85.050 753.600 88.950 ;
        RECT 751.950 82.950 754.050 85.050 ;
        RECT 712.950 79.950 715.050 82.050 ;
        RECT 718.950 79.950 721.050 82.050 ;
        RECT 724.950 79.950 727.050 82.050 ;
        RECT 685.950 76.950 688.050 79.050 ;
        RECT 713.400 70.050 714.600 79.950 ;
        RECT 712.950 67.950 715.050 70.050 ;
        RECT 719.400 64.050 720.600 79.950 ;
        RECT 764.400 76.050 765.600 103.950 ;
        RECT 782.400 100.050 783.600 124.950 ;
        RECT 781.950 97.950 784.050 100.050 ;
        RECT 785.400 99.600 786.600 157.950 ;
        RECT 793.950 145.950 796.050 148.050 ;
        RECT 794.400 142.050 795.600 145.950 ;
        RECT 793.950 139.950 796.050 142.050 ;
        RECT 799.950 139.950 802.050 142.050 ;
        RECT 800.400 124.050 801.600 139.950 ;
        RECT 799.950 121.950 802.050 124.050 ;
        RECT 796.950 103.950 799.050 106.050 ;
        RECT 790.950 99.600 793.050 100.050 ;
        RECT 785.400 98.400 793.050 99.600 ;
        RECT 790.950 97.950 793.050 98.400 ;
        RECT 791.400 82.050 792.600 97.950 ;
        RECT 790.950 79.950 793.050 82.050 ;
        RECT 763.950 73.950 766.050 76.050 ;
        RECT 797.400 73.050 798.600 103.950 ;
        RECT 803.400 97.050 804.600 181.950 ;
        RECT 821.400 175.050 822.600 190.950 ;
        RECT 827.400 175.050 828.600 193.950 ;
        RECT 832.950 187.950 835.050 190.050 ;
        RECT 833.400 184.050 834.600 187.950 ;
        RECT 851.400 184.050 852.600 196.950 ;
        RECT 866.400 186.600 867.600 229.950 ;
        RECT 872.400 196.050 873.600 253.950 ;
        RECT 877.950 208.950 880.050 211.050 ;
        RECT 883.950 208.950 886.050 211.050 ;
        RECT 871.950 193.950 874.050 196.050 ;
        RECT 878.400 193.050 879.600 208.950 ;
        RECT 884.400 199.050 885.600 208.950 ;
        RECT 883.950 196.950 886.050 199.050 ;
        RECT 877.950 190.950 880.050 193.050 ;
        RECT 883.950 190.950 886.050 193.050 ;
        RECT 871.950 186.600 874.050 187.050 ;
        RECT 866.400 185.400 874.050 186.600 ;
        RECT 871.950 184.950 874.050 185.400 ;
        RECT 877.950 186.600 880.050 187.050 ;
        RECT 884.400 186.600 885.600 190.950 ;
        RECT 890.400 190.050 891.600 326.400 ;
        RECT 895.950 322.950 898.050 325.050 ;
        RECT 892.950 307.950 895.050 310.050 ;
        RECT 893.400 226.050 894.600 307.950 ;
        RECT 896.400 274.050 897.600 322.950 ;
        RECT 895.950 271.950 898.050 274.050 ;
        RECT 896.400 262.050 897.600 271.950 ;
        RECT 895.950 259.950 898.050 262.050 ;
        RECT 892.950 223.950 895.050 226.050 ;
        RECT 898.950 223.950 901.050 226.050 ;
        RECT 899.400 220.050 900.600 223.950 ;
        RECT 905.400 220.050 906.600 502.800 ;
        RECT 898.950 217.950 901.050 220.050 ;
        RECT 904.950 217.950 907.050 220.050 ;
        RECT 901.950 208.950 904.050 211.050 ;
        RECT 902.400 202.050 903.600 208.950 ;
        RECT 901.950 201.600 904.050 202.050 ;
        RECT 899.400 200.400 904.050 201.600 ;
        RECT 889.950 187.950 892.050 190.050 ;
        RECT 877.950 185.400 885.600 186.600 ;
        RECT 877.950 184.950 880.050 185.400 ;
        RECT 832.950 181.950 835.050 184.050 ;
        RECT 841.950 181.950 844.050 184.050 ;
        RECT 850.950 181.950 853.050 184.050 ;
        RECT 814.950 172.950 817.050 175.050 ;
        RECT 820.950 172.950 823.050 175.050 ;
        RECT 826.950 172.950 829.050 175.050 ;
        RECT 835.950 172.950 838.050 175.050 ;
        RECT 815.400 163.050 816.600 172.950 ;
        RECT 832.950 166.950 835.050 169.050 ;
        RECT 808.950 160.950 811.050 163.050 ;
        RECT 814.950 160.950 817.050 163.050 ;
        RECT 829.950 160.950 832.050 163.050 ;
        RECT 809.400 133.050 810.600 160.950 ;
        RECT 817.950 141.600 822.000 142.050 ;
        RECT 817.950 139.950 822.600 141.600 ;
        RECT 808.950 132.600 811.050 133.050 ;
        RECT 814.950 132.600 817.050 133.050 ;
        RECT 808.950 131.400 817.050 132.600 ;
        RECT 808.950 130.950 811.050 131.400 ;
        RECT 814.950 130.950 817.050 131.400 ;
        RECT 814.950 124.950 817.050 127.050 ;
        RECT 815.400 97.050 816.600 124.950 ;
        RECT 821.400 124.050 822.600 139.950 ;
        RECT 830.400 133.050 831.600 160.950 ;
        RECT 829.950 130.950 832.050 133.050 ;
        RECT 820.950 121.950 823.050 124.050 ;
        RECT 821.400 106.050 822.600 121.950 ;
        RECT 820.950 103.950 823.050 106.050 ;
        RECT 833.400 97.050 834.600 166.950 ;
        RECT 836.400 142.050 837.600 172.950 ;
        RECT 842.400 142.050 843.600 181.950 ;
        RECT 868.950 175.950 871.050 178.050 ;
        RECT 835.950 139.950 838.050 142.050 ;
        RECT 841.950 139.950 844.050 142.050 ;
        RECT 847.950 139.950 850.050 142.050 ;
        RECT 853.950 139.950 856.050 142.050 ;
        RECT 835.950 124.950 838.050 127.050 ;
        RECT 836.400 106.050 837.600 124.950 ;
        RECT 848.400 121.050 849.600 139.950 ;
        RECT 854.400 133.050 855.600 139.950 ;
        RECT 850.950 131.400 855.600 133.050 ;
        RECT 850.950 130.950 855.000 131.400 ;
        RECT 862.950 130.950 865.050 133.050 ;
        RECT 863.400 127.050 864.600 130.950 ;
        RECT 862.950 124.950 865.050 127.050 ;
        RECT 847.950 118.950 850.050 121.050 ;
        RECT 838.950 115.950 841.050 118.050 ;
        RECT 853.950 115.950 856.050 118.050 ;
        RECT 835.950 103.950 838.050 106.050 ;
        RECT 839.400 97.050 840.600 115.950 ;
        RECT 854.400 109.050 855.600 115.950 ;
        RECT 869.400 115.050 870.600 175.950 ;
        RECT 878.400 133.050 879.600 184.950 ;
        RECT 899.400 184.050 900.600 200.400 ;
        RECT 901.950 199.950 904.050 200.400 ;
        RECT 901.950 187.950 904.050 190.050 ;
        RECT 895.950 182.400 900.600 184.050 ;
        RECT 895.950 181.950 900.000 182.400 ;
        RECT 889.950 172.950 892.050 175.050 ;
        RECT 890.400 142.050 891.600 172.950 ;
        RECT 883.950 139.950 886.050 142.050 ;
        RECT 889.950 139.950 892.050 142.050 ;
        RECT 878.400 131.400 883.050 133.050 ;
        RECT 879.000 130.950 883.050 131.400 ;
        RECT 884.400 121.050 885.600 139.950 ;
        RECT 902.400 138.600 903.600 187.950 ;
        RECT 899.400 137.400 903.600 138.600 ;
        RECT 889.950 130.950 892.050 133.050 ;
        RECT 883.950 120.600 886.050 121.050 ;
        RECT 881.400 119.400 886.050 120.600 ;
        RECT 862.950 112.950 865.050 115.050 ;
        RECT 868.950 112.950 871.050 115.050 ;
        RECT 863.400 109.050 864.600 112.950 ;
        RECT 853.950 106.950 856.050 109.050 ;
        RECT 859.950 107.400 864.600 109.050 ;
        RECT 859.950 106.950 864.000 107.400 ;
        RECT 865.950 103.950 868.050 106.050 ;
        RECT 803.400 95.400 808.050 97.050 ;
        RECT 804.000 94.950 808.050 95.400 ;
        RECT 811.950 95.400 816.600 97.050 ;
        RECT 811.950 94.950 816.000 95.400 ;
        RECT 832.950 94.950 835.050 97.050 ;
        RECT 838.950 94.950 841.050 97.050 ;
        RECT 856.950 94.950 859.050 97.050 ;
        RECT 844.950 79.950 847.050 82.050 ;
        RECT 784.950 70.950 787.050 73.050 ;
        RECT 796.950 70.950 799.050 73.050 ;
        RECT 751.950 67.950 754.050 70.050 ;
        RECT 715.950 61.950 720.600 64.050 ;
        RECT 670.950 59.400 678.600 60.600 ;
        RECT 670.950 58.950 673.050 59.400 ;
        RECT 679.950 58.950 682.050 61.050 ;
        RECT 658.950 52.950 661.050 55.050 ;
        RECT 664.950 54.600 667.050 55.050 ;
        RECT 706.950 54.600 709.050 55.050 ;
        RECT 712.950 54.600 715.050 55.050 ;
        RECT 664.950 53.400 675.600 54.600 ;
        RECT 664.950 52.950 667.050 53.400 ;
        RECT 631.950 49.950 634.050 52.050 ;
        RECT 637.950 49.950 640.050 52.050 ;
        RECT 610.800 40.950 612.900 43.050 ;
        RECT 614.100 40.950 616.200 43.050 ;
        RECT 632.400 40.050 633.600 49.950 ;
        RECT 631.950 37.950 634.050 40.050 ;
        RECT 643.950 34.950 646.050 37.050 ;
        RECT 607.950 31.950 610.050 34.050 ;
        RECT 631.950 31.950 634.050 34.050 ;
        RECT 637.950 31.950 640.050 34.050 ;
        RECT 553.950 25.950 556.050 28.050 ;
        RECT 559.950 25.950 562.050 28.050 ;
        RECT 565.950 25.950 568.050 28.050 ;
        RECT 571.950 25.950 574.050 28.050 ;
        RECT 589.950 25.950 592.050 28.050 ;
        RECT 601.950 25.950 604.050 28.050 ;
        RECT 554.400 21.600 555.600 25.950 ;
        RECT 554.400 20.400 561.600 21.600 ;
        RECT 460.950 17.400 477.600 18.600 ;
        RECT 460.950 16.950 463.050 17.400 ;
        RECT 517.950 16.950 522.600 19.050 ;
        RECT 535.950 16.950 538.050 19.050 ;
        RECT 541.950 16.950 544.050 19.050 ;
        RECT 556.950 16.950 559.050 19.050 ;
        RECT 361.950 10.950 364.050 13.050 ;
        RECT 382.950 10.950 385.050 13.050 ;
        RECT 421.950 10.950 424.050 13.050 ;
        RECT 454.950 10.950 457.050 13.050 ;
        RECT 502.950 12.600 505.050 13.050 ;
        RECT 494.400 11.400 505.050 12.600 ;
        RECT 494.400 7.050 495.600 11.400 ;
        RECT 502.950 10.950 505.050 11.400 ;
        RECT 511.950 7.950 514.050 10.050 ;
        RECT 334.950 4.950 337.050 7.050 ;
        RECT 493.950 4.950 496.050 7.050 ;
        RECT 512.400 4.050 513.600 7.950 ;
        RECT 521.400 7.050 522.600 16.950 ;
        RECT 536.400 7.050 537.600 16.950 ;
        RECT 557.400 10.050 558.600 16.950 ;
        RECT 560.400 15.600 561.600 20.400 ;
        RECT 562.950 18.600 565.050 19.050 ;
        RECT 572.400 18.600 573.600 25.950 ;
        RECT 608.400 19.050 609.600 31.950 ;
        RECT 632.400 28.050 633.600 31.950 ;
        RECT 625.950 24.600 628.050 28.050 ;
        RECT 631.950 25.950 634.050 28.050 ;
        RECT 638.400 24.600 639.600 31.950 ;
        RECT 644.400 31.050 645.600 34.950 ;
        RECT 643.950 28.950 646.050 31.050 ;
        RECT 659.400 28.050 660.600 52.950 ;
        RECT 674.400 51.600 675.600 53.400 ;
        RECT 706.950 53.400 715.050 54.600 ;
        RECT 706.950 52.950 709.050 53.400 ;
        RECT 712.950 52.950 715.050 53.400 ;
        RECT 679.950 51.600 682.050 52.050 ;
        RECT 674.400 50.400 682.050 51.600 ;
        RECT 679.950 49.950 682.050 50.400 ;
        RECT 688.950 51.600 691.050 52.050 ;
        RECT 688.950 51.000 702.600 51.600 ;
        RECT 688.950 50.400 703.050 51.000 ;
        RECT 688.950 49.950 691.050 50.400 ;
        RECT 700.950 46.950 703.050 50.400 ;
        RECT 694.950 40.950 697.050 43.050 ;
        RECT 695.400 28.050 696.600 40.950 ;
        RECT 719.400 34.050 720.600 61.950 ;
        RECT 721.950 58.950 724.050 61.050 ;
        RECT 722.400 49.050 723.600 58.950 ;
        RECT 752.400 55.050 753.600 67.950 ;
        RECT 785.400 66.600 786.600 70.950 ;
        RECT 793.950 67.950 796.050 70.050 ;
        RECT 808.950 69.600 811.050 70.050 ;
        RECT 820.950 69.600 823.050 70.050 ;
        RECT 808.950 68.400 823.050 69.600 ;
        RECT 808.950 67.950 811.050 68.400 ;
        RECT 820.950 67.950 823.050 68.400 ;
        RECT 829.950 69.600 832.050 70.050 ;
        RECT 841.950 69.600 844.050 70.050 ;
        RECT 829.950 68.400 844.050 69.600 ;
        RECT 829.950 67.950 832.050 68.400 ;
        RECT 841.950 67.950 844.050 68.400 ;
        RECT 782.400 66.000 786.600 66.600 ;
        RECT 781.950 65.400 786.600 66.000 ;
        RECT 775.950 61.950 778.050 64.050 ;
        RECT 781.950 61.950 784.050 65.400 ;
        RECT 769.950 58.950 772.050 61.050 ;
        RECT 751.950 52.950 754.050 55.050 ;
        RECT 730.950 49.950 733.050 52.050 ;
        RECT 736.950 49.950 739.050 52.050 ;
        RECT 721.950 46.950 724.050 49.050 ;
        RECT 731.400 40.050 732.600 49.950 ;
        RECT 737.400 46.050 738.600 49.950 ;
        RECT 770.400 49.050 771.600 58.950 ;
        RECT 772.950 52.950 775.050 55.050 ;
        RECT 769.950 46.950 772.050 49.050 ;
        RECT 736.950 43.950 739.050 46.050 ;
        RECT 773.400 40.050 774.600 52.950 ;
        RECT 730.950 37.950 733.050 40.050 ;
        RECT 736.950 37.950 739.050 40.050 ;
        RECT 760.950 37.950 763.050 40.050 ;
        RECT 772.950 37.950 775.050 40.050 ;
        RECT 718.950 31.950 721.050 34.050 ;
        RECT 730.950 31.950 733.050 34.050 ;
        RECT 658.950 25.950 661.050 28.050 ;
        RECT 694.950 25.950 697.050 28.050 ;
        RECT 625.950 24.000 639.600 24.600 ;
        RECT 626.400 23.400 639.600 24.000 ;
        RECT 731.400 19.050 732.600 31.950 ;
        RECT 737.400 19.050 738.600 37.950 ;
        RECT 761.400 28.050 762.600 37.950 ;
        RECT 776.400 37.050 777.600 61.950 ;
        RECT 794.400 55.050 795.600 67.950 ;
        RECT 798.000 63.600 802.050 64.050 ;
        RECT 797.400 61.950 802.050 63.600 ;
        RECT 808.950 61.950 811.050 64.050 ;
        RECT 838.950 63.600 841.050 67.050 ;
        RECT 836.400 63.000 841.050 63.600 ;
        RECT 836.400 62.400 840.600 63.000 ;
        RECT 784.950 52.950 787.050 55.050 ;
        RECT 793.950 52.950 796.050 55.050 ;
        RECT 785.400 49.050 786.600 52.950 ;
        RECT 797.400 49.050 798.600 61.950 ;
        RECT 809.400 55.050 810.600 61.950 ;
        RECT 829.950 60.600 832.050 61.050 ;
        RECT 836.400 60.600 837.600 62.400 ;
        RECT 829.950 59.400 837.600 60.600 ;
        RECT 838.950 60.600 841.050 61.050 ;
        RECT 845.400 60.600 846.600 79.950 ;
        RECT 853.950 70.950 856.050 73.050 ;
        RECT 838.950 59.400 846.600 60.600 ;
        RECT 829.950 58.950 832.050 59.400 ;
        RECT 838.950 58.950 841.050 59.400 ;
        RECT 809.400 52.950 814.050 55.050 ;
        RECT 778.950 46.950 781.050 49.050 ;
        RECT 784.950 46.950 787.050 49.050 ;
        RECT 796.950 46.950 799.050 49.050 ;
        RECT 770.100 34.950 772.200 37.050 ;
        RECT 775.950 34.950 778.050 37.050 ;
        RECT 770.400 28.050 771.600 34.950 ;
        RECT 772.950 31.950 775.050 34.050 ;
        RECT 742.950 25.950 745.050 28.050 ;
        RECT 760.950 25.950 763.050 28.050 ;
        RECT 769.950 25.950 772.050 28.050 ;
        RECT 580.950 18.600 583.050 19.050 ;
        RECT 562.950 17.400 573.600 18.600 ;
        RECT 575.400 18.000 583.050 18.600 ;
        RECT 574.950 17.400 583.050 18.000 ;
        RECT 562.950 16.950 565.050 17.400 ;
        RECT 565.950 15.600 568.050 16.050 ;
        RECT 560.400 14.400 568.050 15.600 ;
        RECT 565.950 13.950 568.050 14.400 ;
        RECT 574.950 13.950 577.050 17.400 ;
        RECT 580.950 16.950 583.050 17.400 ;
        RECT 586.950 16.950 589.050 19.050 ;
        RECT 604.950 17.400 609.600 19.050 ;
        RECT 604.950 16.950 609.000 17.400 ;
        RECT 622.950 16.950 625.050 19.050 ;
        RECT 628.950 16.950 631.050 19.050 ;
        RECT 730.950 16.950 733.050 19.050 ;
        RECT 736.950 16.950 739.050 19.050 ;
        RECT 587.400 10.050 588.600 16.950 ;
        RECT 623.400 13.050 624.600 16.950 ;
        RECT 629.400 13.050 630.600 16.950 ;
        RECT 743.400 13.050 744.600 25.950 ;
        RECT 748.950 22.950 751.050 25.050 ;
        RECT 749.400 19.050 750.600 22.950 ;
        RECT 773.400 19.050 774.600 31.950 ;
        RECT 779.400 19.050 780.600 46.950 ;
        RECT 797.400 40.050 798.600 46.950 ;
        RECT 809.400 46.050 810.600 52.950 ;
        RECT 808.950 43.950 811.050 46.050 ;
        RECT 796.950 37.950 799.050 40.050 ;
        RECT 784.950 31.950 787.050 34.050 ;
        RECT 832.950 33.600 835.050 37.050 ;
        RECT 830.400 33.000 835.050 33.600 ;
        RECT 839.400 33.600 840.600 58.950 ;
        RECT 854.400 55.050 855.600 70.950 ;
        RECT 857.400 64.050 858.600 94.950 ;
        RECT 866.400 73.050 867.600 103.950 ;
        RECT 865.950 70.950 868.050 73.050 ;
        RECT 862.950 67.950 865.050 70.050 ;
        RECT 863.400 64.050 864.600 67.950 ;
        RECT 856.950 61.950 859.050 64.050 ;
        RECT 862.950 61.950 865.050 64.050 ;
        RECT 853.950 52.950 856.050 55.050 ;
        RECT 869.400 49.050 870.600 112.950 ;
        RECT 881.400 97.050 882.600 119.400 ;
        RECT 883.950 118.950 886.050 119.400 ;
        RECT 883.950 105.600 888.000 106.050 ;
        RECT 883.950 103.950 888.600 105.600 ;
        RECT 874.950 94.950 877.050 97.050 ;
        RECT 880.950 94.950 883.050 97.050 ;
        RECT 875.400 85.050 876.600 94.950 ;
        RECT 887.400 94.050 888.600 103.950 ;
        RECT 890.400 97.050 891.600 130.950 ;
        RECT 892.950 124.950 895.050 127.050 ;
        RECT 893.400 100.050 894.600 124.950 ;
        RECT 899.400 109.050 900.600 137.400 ;
        RECT 904.950 133.950 907.050 136.050 ;
        RECT 895.950 106.950 898.050 109.050 ;
        RECT 899.400 106.950 904.050 109.050 ;
        RECT 892.950 97.950 895.050 100.050 ;
        RECT 889.950 94.950 892.050 97.050 ;
        RECT 896.400 94.050 897.600 106.950 ;
        RECT 886.950 91.950 889.050 94.050 ;
        RECT 895.950 91.950 898.050 94.050 ;
        RECT 874.950 82.950 877.050 85.050 ;
        RECT 883.950 82.950 886.050 85.050 ;
        RECT 884.400 70.050 885.600 82.950 ;
        RECT 883.950 67.950 886.050 70.050 ;
        RECT 889.950 67.950 892.050 70.050 ;
        RECT 890.400 64.050 891.600 67.950 ;
        RECT 896.400 64.050 897.600 91.950 ;
        RECT 883.950 61.950 886.050 64.050 ;
        RECT 889.950 61.950 892.050 64.050 ;
        RECT 895.950 61.950 898.050 64.050 ;
        RECT 880.950 49.950 883.050 52.050 ;
        RECT 868.950 46.950 871.050 49.050 ;
        RECT 881.400 43.050 882.600 49.950 ;
        RECT 880.950 40.950 883.050 43.050 ;
        RECT 884.400 39.600 885.600 61.950 ;
        RECT 899.400 57.600 900.600 106.950 ;
        RECT 896.400 56.400 900.600 57.600 ;
        RECT 886.950 54.600 889.050 55.050 ;
        RECT 896.400 54.600 897.600 56.400 ;
        RECT 886.950 53.400 897.600 54.600 ;
        RECT 886.950 52.950 889.050 53.400 ;
        RECT 898.950 52.950 901.050 55.050 ;
        RECT 899.400 49.050 900.600 52.950 ;
        RECT 898.950 46.950 901.050 49.050 ;
        RECT 892.950 40.950 895.050 43.050 ;
        RECT 886.950 39.600 889.050 40.050 ;
        RECT 884.400 38.400 889.050 39.600 ;
        RECT 886.950 37.950 889.050 38.400 ;
        RECT 841.950 36.600 844.050 37.050 ;
        RECT 841.950 35.400 855.600 36.600 ;
        RECT 841.950 34.950 844.050 35.400 ;
        RECT 830.400 32.400 834.600 33.000 ;
        RECT 839.400 32.400 843.600 33.600 ;
        RECT 785.400 28.050 786.600 31.950 ;
        RECT 796.950 28.950 799.050 31.050 ;
        RECT 805.950 30.600 808.050 31.050 ;
        RECT 805.950 30.000 819.600 30.600 ;
        RECT 805.950 29.400 820.050 30.000 ;
        RECT 805.950 28.950 808.050 29.400 ;
        RECT 785.400 26.400 790.050 28.050 ;
        RECT 786.000 25.950 790.050 26.400 ;
        RECT 749.400 17.400 754.050 19.050 ;
        RECT 750.000 16.950 754.050 17.400 ;
        RECT 757.950 16.950 760.050 19.050 ;
        RECT 772.950 16.950 775.050 19.050 ;
        RECT 778.950 16.950 781.050 19.050 ;
        RECT 758.400 13.050 759.600 16.950 ;
        RECT 622.950 10.950 625.050 13.050 ;
        RECT 628.950 10.950 631.050 13.050 ;
        RECT 742.950 10.950 745.050 13.050 ;
        RECT 757.950 10.950 760.050 13.050 ;
        RECT 773.400 10.050 774.600 16.950 ;
        RECT 784.950 12.600 787.050 13.050 ;
        RECT 797.400 12.600 798.600 28.950 ;
        RECT 817.950 25.950 820.050 29.400 ;
        RECT 823.950 27.600 826.050 28.050 ;
        RECT 830.400 27.600 831.600 32.400 ;
        RECT 842.400 31.050 843.600 32.400 ;
        RECT 832.950 28.950 835.050 31.050 ;
        RECT 841.950 28.950 844.050 31.050 ;
        RECT 823.950 26.400 831.600 27.600 ;
        RECT 823.950 25.950 826.050 26.400 ;
        RECT 805.950 19.950 808.050 22.050 ;
        RECT 814.950 21.600 817.050 22.050 ;
        RECT 833.400 21.600 834.600 28.950 ;
        RECT 842.400 24.600 843.600 28.950 ;
        RECT 854.400 28.050 855.600 35.400 ;
        RECT 887.400 31.050 888.600 37.950 ;
        RECT 893.400 31.050 894.600 40.950 ;
        RECT 886.950 28.950 889.050 31.050 ;
        RECT 892.950 28.950 895.050 31.050 ;
        RECT 853.950 25.950 856.050 28.050 ;
        RECT 842.400 23.400 846.600 24.600 ;
        RECT 814.950 20.400 834.600 21.600 ;
        RECT 814.950 19.950 817.050 20.400 ;
        RECT 784.950 11.400 798.600 12.600 ;
        RECT 784.950 10.950 787.050 11.400 ;
        RECT 556.950 7.950 559.050 10.050 ;
        RECT 586.950 7.950 589.050 10.050 ;
        RECT 772.950 7.950 775.050 10.050 ;
        RECT 806.400 7.050 807.600 19.950 ;
        RECT 841.950 18.600 844.050 22.050 ;
        RECT 845.400 21.600 846.600 23.400 ;
        RECT 850.950 21.600 853.050 22.050 ;
        RECT 883.950 21.600 886.050 22.050 ;
        RECT 845.400 20.400 853.050 21.600 ;
        RECT 878.400 21.000 886.050 21.600 ;
        RECT 850.950 19.950 853.050 20.400 ;
        RECT 877.950 20.400 886.050 21.000 ;
        RECT 841.950 18.000 849.600 18.600 ;
        RECT 842.400 17.400 849.600 18.000 ;
        RECT 848.400 16.050 849.600 17.400 ;
        RECT 877.950 16.950 880.050 20.400 ;
        RECT 883.950 19.950 886.050 20.400 ;
        RECT 895.950 19.950 898.050 22.050 ;
        RECT 896.400 16.050 897.600 19.950 ;
        RECT 905.400 16.050 906.600 133.950 ;
        RECT 908.400 133.050 909.600 679.950 ;
        RECT 911.400 625.200 912.600 691.950 ;
        RECT 910.950 623.100 913.050 625.200 ;
        RECT 910.950 619.800 913.050 621.900 ;
        RECT 911.400 538.050 912.600 619.800 ;
        RECT 910.950 535.950 913.050 538.050 ;
        RECT 910.950 505.950 913.050 508.050 ;
        RECT 911.400 136.050 912.600 505.950 ;
        RECT 910.950 133.950 913.050 136.050 ;
        RECT 907.950 130.950 910.050 133.050 ;
        RECT 848.400 14.400 853.050 16.050 ;
        RECT 849.000 13.950 853.050 14.400 ;
        RECT 862.950 15.600 865.050 16.050 ;
        RECT 874.950 15.600 877.050 16.050 ;
        RECT 862.950 14.400 877.050 15.600 ;
        RECT 862.950 13.950 865.050 14.400 ;
        RECT 874.950 13.950 877.050 14.400 ;
        RECT 895.950 13.950 898.050 16.050 ;
        RECT 904.950 13.950 907.050 16.050 ;
        RECT 520.950 4.950 523.050 7.050 ;
        RECT 535.950 4.950 538.050 7.050 ;
        RECT 805.950 4.950 808.050 7.050 ;
        RECT 64.950 1.950 67.050 4.050 ;
        RECT 304.950 1.950 307.050 4.050 ;
        RECT 511.950 1.950 514.050 4.050 ;
  END
END fir_pe
END LIBRARY

