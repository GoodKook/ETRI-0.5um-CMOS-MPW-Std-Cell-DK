magic
tech scmos
magscale 1 2
timestamp 1702308830
<< nwell >>
rect -13 154 53 272
<< ntransistor >>
rect 18 14 22 54
<< ptransistor >>
rect 18 166 22 246
<< ndiffusion >>
rect 16 14 18 54
rect 22 14 24 54
<< pdiffusion >>
rect 16 166 18 246
rect 22 166 24 246
<< ndcontact >>
rect 4 14 16 54
rect 24 14 36 54
<< pdcontact >>
rect 4 166 16 246
rect 24 166 36 246
<< psubstratepcontact >>
rect -6 -6 46 6
<< nsubstratencontact >>
rect -6 254 46 266
<< polysilicon >>
rect 18 246 22 250
rect 18 117 22 166
rect 17 105 22 117
rect 18 54 22 105
rect 18 10 22 14
<< polycontact >>
rect 5 105 17 117
<< metal1 >>
rect -6 266 46 268
rect -6 252 46 254
rect 4 246 16 252
rect 3 123 17 137
rect 5 117 17 123
rect 26 117 34 166
rect 23 103 37 117
rect 26 54 34 103
rect 4 8 16 14
rect -6 6 46 8
rect -6 -8 46 -6
<< m1p >>
rect -6 252 46 268
rect 3 123 17 137
rect 23 103 37 117
rect -6 -8 46 8
<< labels >>
rlabel nsubstratencontact 20 260 20 260 0 vdd
port 3 nsew power bidirectional abutment
rlabel psubstratepcontact 20 0 20 0 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 10 127 10 127 0 A
port 1 nsew signal input
rlabel metal1 30 111 30 111 0 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 40 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
