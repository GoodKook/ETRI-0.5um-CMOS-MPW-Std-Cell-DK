magic
tech scmos
timestamp 1702508443
<< nwell >>
rect -6 77 66 136
<< ntransistor >>
rect 9 7 11 27
rect 19 7 21 27
rect 24 7 26 27
rect 34 7 36 27
rect 39 7 41 27
rect 49 7 51 27
<< ptransistor >>
rect 9 83 11 123
rect 19 83 21 123
rect 24 83 26 123
rect 34 83 36 123
rect 39 83 41 123
rect 49 83 51 123
<< ndiffusion >>
rect 8 7 9 27
rect 11 24 19 27
rect 11 7 12 24
rect 18 7 19 24
rect 21 7 24 27
rect 26 7 27 27
rect 33 7 34 27
rect 36 7 39 27
rect 41 24 49 27
rect 41 7 42 24
rect 48 7 49 24
rect 51 7 52 27
<< pdiffusion >>
rect 8 83 9 123
rect 11 90 12 123
rect 18 90 19 123
rect 11 83 19 90
rect 21 83 24 123
rect 26 83 27 123
rect 33 83 34 123
rect 36 83 39 123
rect 41 90 42 123
rect 48 90 49 123
rect 41 83 49 90
rect 51 83 52 123
<< ndcontact >>
rect 2 7 8 27
rect 12 7 18 24
rect 27 7 33 27
rect 42 7 48 24
rect 52 7 58 27
<< pdcontact >>
rect 2 83 8 123
rect 12 90 18 123
rect 27 83 33 123
rect 42 90 48 123
rect 52 83 58 123
<< psubstratepcontact >>
rect -3 -3 63 3
<< nsubstratencontact >>
rect -3 127 63 133
<< polysilicon >>
rect 9 123 11 125
rect 19 123 21 125
rect 24 123 26 125
rect 34 123 36 125
rect 39 123 41 125
rect 49 123 51 125
rect 9 27 11 83
rect 19 80 21 83
rect 13 78 21 80
rect 13 31 15 78
rect 24 76 26 83
rect 34 77 36 83
rect 39 82 41 83
rect 49 82 51 83
rect 39 79 51 82
rect 24 74 27 76
rect 34 75 42 77
rect 25 57 27 74
rect 25 54 32 57
rect 40 55 42 75
rect 25 43 26 49
rect 13 29 21 31
rect 19 27 21 29
rect 24 27 26 43
rect 30 41 32 54
rect 30 39 36 41
rect 34 27 36 39
rect 49 37 51 79
rect 39 34 51 37
rect 39 27 41 34
rect 49 27 51 34
rect 9 5 11 7
rect 19 5 21 7
rect 24 5 26 7
rect 34 5 36 7
rect 39 5 41 7
rect 49 5 51 7
<< polycontact >>
rect 3 45 9 51
rect 15 64 21 70
rect 19 54 25 60
rect 19 43 25 49
rect 36 49 42 55
rect 51 58 57 64
<< metal1 >>
rect -3 133 63 134
rect -3 126 63 127
rect 12 123 18 126
rect 42 123 48 126
rect 8 83 17 86
rect 29 78 33 83
rect 49 83 52 87
rect 29 75 34 78
rect 31 68 34 75
rect 9 54 19 58
rect 28 58 36 61
rect 4 33 25 36
rect 28 39 32 58
rect 4 27 8 33
rect 28 32 31 39
rect 28 27 32 32
rect 49 27 58 30
rect 12 4 18 7
rect 42 4 48 7
rect -3 3 63 4
rect -3 -4 63 -3
<< m2contact >>
rect 10 76 17 83
rect 42 80 49 87
rect 21 64 28 71
rect 31 61 38 68
rect 2 51 9 58
rect 18 36 25 43
rect 51 51 58 58
rect 35 42 42 49
rect 31 32 38 39
rect 42 27 49 34
<< metal2 >>
rect 3 58 7 67
rect 13 46 16 76
rect 33 68 37 77
rect 25 56 28 64
rect 44 56 48 80
rect 25 52 48 56
rect 13 43 35 46
rect 13 42 18 43
rect 25 42 35 43
rect 45 34 48 52
rect 53 43 57 51
rect 33 23 37 32
<< m1p >>
rect -3 126 63 134
rect -3 -4 63 4
<< m2p >>
rect 33 69 37 77
rect 3 59 7 67
rect 53 43 57 50
rect 33 23 37 31
<< labels >>
rlabel metal2 5 65 5 65 1 A
port 1 n signal input
rlabel metal2 55 45 55 45 5 B
port 2 n signal input
rlabel metal2 35 76 35 76 5 Y
port 3 n signal output
rlabel metal1 -3 126 63 134 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 -3 -4 63 4 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal2 35 25 35 25 1 Y
port 3 n signal output
<< properties >>
string FIXED_BBOX 0 0 60 130
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
