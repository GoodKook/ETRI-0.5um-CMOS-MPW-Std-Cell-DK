magic
tech scmos
magscale 1 3
timestamp 1555596690
<< checkpaint >>
rect -55 -58 136 194
use nmos4_CDNS_723012252917  nmos4_CDNS_723012252917_0
timestamp 1555596690
transform 1 0 0 0 1 0
box 5 2 76 134
<< end >>
