magic
tech scmos
magscale 1 2
timestamp 1728304496
<< nwell >>
rect -12 134 292 252
<< ntransistor >>
rect 21 14 25 54
rect 41 14 45 54
rect 61 14 65 54
rect 81 14 85 54
rect 101 14 105 54
rect 121 14 125 54
rect 141 14 145 54
rect 161 14 165 54
rect 181 14 185 54
rect 201 14 205 54
rect 221 14 225 54
rect 241 14 245 54
<< ptransistor >>
rect 21 146 25 226
rect 41 146 45 226
rect 61 146 65 226
rect 81 146 85 226
rect 101 146 105 226
rect 121 146 125 226
rect 141 146 145 226
rect 161 146 165 226
rect 181 146 185 226
rect 201 146 205 226
rect 221 146 225 226
rect 241 146 245 226
<< ndiffusion >>
rect 19 14 21 54
rect 25 14 27 54
rect 39 14 41 54
rect 45 14 47 54
rect 59 14 61 54
rect 65 14 67 54
rect 79 14 81 54
rect 85 14 87 54
rect 99 14 101 54
rect 105 14 107 54
rect 119 14 121 54
rect 125 14 127 54
rect 139 14 141 54
rect 145 14 147 54
rect 159 14 161 54
rect 165 14 167 54
rect 179 14 181 54
rect 185 14 187 54
rect 199 14 201 54
rect 205 14 207 54
rect 219 14 221 54
rect 225 14 227 54
rect 239 14 241 54
rect 245 14 247 54
<< pdiffusion >>
rect 19 146 21 226
rect 25 146 27 226
rect 39 146 41 226
rect 45 146 47 226
rect 59 146 61 226
rect 65 146 67 226
rect 79 146 81 226
rect 85 146 87 226
rect 99 146 101 226
rect 105 146 107 226
rect 119 146 121 226
rect 125 146 127 226
rect 139 146 141 226
rect 145 146 147 226
rect 159 146 161 226
rect 165 146 167 226
rect 179 146 181 226
rect 185 146 187 226
rect 199 146 201 226
rect 205 146 207 226
rect 219 146 221 226
rect 225 146 227 226
rect 239 146 241 226
rect 245 146 247 226
<< ndcontact >>
rect 7 14 19 54
rect 27 14 39 54
rect 47 14 59 54
rect 67 14 79 54
rect 87 14 99 54
rect 107 14 119 54
rect 127 14 139 54
rect 147 14 159 54
rect 167 14 179 54
rect 187 14 199 54
rect 207 14 219 54
rect 227 14 239 54
rect 247 14 259 54
<< pdcontact >>
rect 7 146 19 226
rect 27 146 39 226
rect 47 146 59 226
rect 67 146 79 226
rect 87 146 99 226
rect 107 146 119 226
rect 127 146 139 226
rect 147 146 159 226
rect 167 146 179 226
rect 187 146 199 226
rect 207 146 219 226
rect 227 146 239 226
rect 247 146 259 226
<< psubstratepcontact >>
rect -6 -6 286 6
<< nsubstratencontact >>
rect -6 234 286 246
<< polysilicon >>
rect 21 226 25 230
rect 41 226 45 230
rect 61 226 65 230
rect 81 226 85 230
rect 101 226 105 230
rect 121 226 125 230
rect 141 226 145 230
rect 161 226 165 230
rect 181 226 185 230
rect 201 226 205 230
rect 221 226 225 230
rect 241 226 245 230
rect 21 89 25 146
rect 41 89 45 146
rect 21 77 24 89
rect 36 77 45 89
rect 61 86 65 146
rect 81 86 85 146
rect 101 86 105 146
rect 121 86 125 146
rect 141 86 145 146
rect 161 86 165 146
rect 181 86 185 146
rect 201 86 205 146
rect 221 86 225 146
rect 241 86 245 146
rect 21 54 25 77
rect 41 54 45 77
rect 72 74 85 86
rect 112 74 125 86
rect 152 74 165 86
rect 192 74 205 86
rect 232 74 245 86
rect 61 54 65 74
rect 81 54 85 74
rect 101 54 105 74
rect 121 54 125 74
rect 141 54 145 74
rect 161 54 165 74
rect 181 54 185 74
rect 201 54 205 74
rect 221 54 225 74
rect 241 54 245 74
rect 21 10 25 14
rect 41 10 45 14
rect 61 10 65 14
rect 81 10 85 14
rect 101 10 105 14
rect 121 10 125 14
rect 141 10 145 14
rect 161 10 165 14
rect 181 10 185 14
rect 201 10 205 14
rect 221 10 225 14
rect 241 10 245 14
<< polycontact >>
rect 24 77 36 89
rect 60 74 72 86
rect 100 74 112 86
rect 140 74 152 86
rect 180 74 192 86
rect 220 74 232 86
<< metal1 >>
rect -6 246 286 248
rect -6 232 286 234
rect 7 226 19 232
rect 47 226 59 232
rect 87 226 99 232
rect 127 226 139 232
rect 167 226 179 232
rect 207 226 219 232
rect 247 226 259 232
rect 26 140 38 146
rect 66 140 78 146
rect 107 140 119 146
rect 146 140 158 146
rect 187 140 199 146
rect 226 140 238 146
rect 26 132 53 140
rect 66 132 92 140
rect 107 132 132 140
rect 146 132 174 140
rect 187 132 208 140
rect 226 132 248 140
rect 45 86 53 132
rect 84 86 92 132
rect 124 86 132 132
rect 166 86 174 132
rect 200 86 208 132
rect 240 103 248 132
rect 240 89 243 103
rect 45 74 60 86
rect 84 74 100 86
rect 124 74 140 86
rect 166 74 180 86
rect 200 74 220 86
rect 45 68 53 74
rect 84 68 92 74
rect 124 68 132 74
rect 166 68 174 74
rect 200 68 208 74
rect 240 68 248 89
rect 27 60 53 68
rect 67 60 92 68
rect 107 60 132 68
rect 146 60 174 68
rect 187 60 208 68
rect 227 60 248 68
rect 27 54 39 60
rect 67 54 79 60
rect 107 54 119 60
rect 146 54 158 60
rect 187 54 199 60
rect 227 54 239 60
rect 7 8 19 14
rect 47 8 59 14
rect 87 8 99 14
rect 127 8 139 14
rect 167 8 179 14
rect 207 8 219 14
rect 247 8 259 14
rect -6 6 286 8
rect -6 -8 286 -6
<< m2contact >>
rect 23 89 37 103
rect 243 89 257 103
<< metal2 >>
rect 23 103 37 117
rect 243 103 257 117
<< m1p >>
rect -6 232 286 248
rect -6 -8 286 8
<< m2p >>
rect 23 103 37 117
rect 243 103 257 117
<< labels >>
rlabel metal1 -6 -8 286 8 0 gnd
port 3 nsew ground bidirectional abutment
rlabel metal1 -6 232 286 248 0 vdd
port 2 nsew power bidirectional abutment
rlabel metal2 23 103 37 117 0 A
port 0 nsew signal input
rlabel metal2 243 103 257 117 0 Y
port 1 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 280 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
