magic
tech scmos
magscale 1 3
timestamp 1555589239
<< checkpaint >>
rect -60 -90 619 480
<< metal1 >>
rect 68 204 285 220
rect 108 176 468 192
<< metal2 >>
rect 0 220 20 420
rect 149 396 168 420
rect 149 376 391 396
rect 149 276 168 376
rect 149 256 180 276
rect 371 256 391 376
rect 0 200 54 220
rect 238 -30 258 46
rect 511 -24 531 46
use INV  INV_0
timestamp 1555589239
transform 1 0 15 0 1 47
box -1 -21 93 307
use NAND2  NAND2_0
timestamp 1555589239
transform 1 0 392 0 1 47
box -1 -21 167 307
use NOR2  NOR2_0
timestamp 1555589239
transform 1 0 149 0 1 47
box -32 -21 212 323
use via1_CDNS_704676826054  via1_CDNS_704676826054_0
timestamp 1555589239
transform 1 0 245 0 1 200
box 0 0 20 20
use via1_CDNS_704676826054  via1_CDNS_704676826054_1
timestamp 1555589239
transform 1 0 108 0 1 176
box 0 0 20 20
use via1_CDNS_704676826054  via1_CDNS_704676826054_2
timestamp 1555589239
transform 1 0 48 0 1 200
box 0 0 20 20
use via1_CDNS_704676826054  via1_CDNS_704676826054_3
timestamp 1555589239
transform 1 0 478 0 1 176
box 0 0 20 20
use via1_CDNS_704676826054  via1_CDNS_704676826054_4
timestamp 1555589239
transform 1 0 265 0 1 200
box 0 0 20 20
use via1_CDNS_704676826054  via1_CDNS_704676826054_5
timestamp 1555589239
transform 1 0 28 0 1 200
box 0 0 20 20
use via1_CDNS_704676826054  via1_CDNS_704676826054_6
timestamp 1555589239
transform 1 0 88 0 1 176
box 0 0 20 20
use via1_CDNS_704676826054  via1_CDNS_704676826054_7
timestamp 1555589239
transform 1 0 458 0 1 176
box 0 0 20 20
<< labels >>
flabel m2p s 520 -17 520 -17 0 FreeSans 19 0 0 0 ND
flabel m2p s 247 -17 247 -17 0 FreeSans 19 0 0 0 PD
flabel m2p s 158 417 158 417 0 FreeSans 19 0 0 0 A
flabel m2p s 7 420 7 420 0 FreeSans 19 0 0 0 OE
<< end >>
