magic
tech scmos
magscale 1 2
timestamp 1702310787
<< nwell >>
rect -13 154 93 272
<< ntransistor >>
rect 18 14 22 74
rect 28 14 32 74
rect 42 14 46 74
<< ptransistor >>
rect 18 206 22 246
rect 38 206 42 246
rect 58 206 62 246
<< ndiffusion >>
rect 16 14 18 74
rect 22 14 28 74
rect 32 14 42 74
rect 46 73 60 74
rect 46 14 48 73
<< pdiffusion >>
rect 16 206 18 246
rect 22 206 24 246
rect 36 206 38 246
rect 42 210 44 246
rect 56 210 58 246
rect 42 206 58 210
rect 62 206 64 246
<< ndcontact >>
rect 4 14 16 74
rect 48 14 60 73
<< pdcontact >>
rect 4 206 16 246
rect 24 206 36 246
rect 44 210 56 246
rect 64 206 76 246
<< psubstratepcontact >>
rect -6 -6 86 6
<< nsubstratencontact >>
rect -6 254 86 266
<< polysilicon >>
rect 18 246 22 250
rect 38 246 42 250
rect 58 246 62 250
rect 18 198 22 206
rect 38 198 42 206
rect 13 193 22 198
rect 28 193 42 198
rect 13 117 18 193
rect 17 105 22 117
rect 18 74 22 105
rect 28 100 32 193
rect 58 120 62 206
rect 57 108 62 120
rect 28 88 30 100
rect 28 74 32 88
rect 58 80 62 108
rect 42 76 62 80
rect 42 74 46 76
rect 18 10 22 14
rect 28 10 32 14
rect 42 10 46 14
<< polycontact >>
rect 5 105 17 117
rect 45 108 57 120
rect 30 88 42 100
<< metal1 >>
rect -6 266 86 268
rect -6 252 86 254
rect 4 246 16 252
rect 44 246 56 252
rect 26 204 36 206
rect 64 204 74 206
rect 26 198 74 204
rect 3 123 17 137
rect 43 123 57 137
rect 5 117 17 123
rect 45 120 57 123
rect 23 103 37 117
rect 66 117 74 198
rect 63 103 77 117
rect 26 100 37 103
rect 26 88 30 100
rect 66 76 74 103
rect 48 73 74 76
rect 60 70 74 73
rect 4 8 16 14
rect -6 6 86 8
rect -6 -8 86 -6
<< m1p >>
rect -6 252 86 268
rect 3 123 17 137
rect 43 123 57 137
rect 23 103 37 117
rect 63 103 77 117
rect -6 -8 86 8
<< labels >>
rlabel nsubstratencontact 40 260 40 260 0 vdd
port 5 nsew power bidirectional abutment
rlabel psubstratepcontact 40 0 40 0 0 gnd
port 6 nsew ground bidirectional abutment
rlabel metal1 10 131 10 131 0 A
port 1 nsew signal input
rlabel metal1 30 110 30 110 0 B
port 2 nsew signal input
rlabel metal1 50 131 50 131 0 C
port 3 nsew signal input
rlabel metal1 70 111 70 111 0 Y
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 80 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
