magic
tech scmos
magscale 1 2
timestamp 1727907586
<< nwell >>
rect -13 134 112 252
<< ntransistor >>
rect 20 14 24 54
rect 28 14 32 54
rect 50 14 54 34
<< ptransistor >>
rect 20 186 24 226
rect 40 186 44 226
rect 60 186 64 226
<< ndiffusion >>
rect 18 14 20 54
rect 24 14 28 54
rect 32 14 34 54
rect 46 14 50 34
rect 54 14 56 34
<< pdiffusion >>
rect 18 186 20 226
rect 24 186 26 226
rect 38 186 40 226
rect 44 186 46 226
rect 58 186 60 226
rect 64 186 66 226
<< ndcontact >>
rect 6 14 18 54
rect 34 14 46 54
rect 56 14 68 34
<< pdcontact >>
rect 6 186 18 226
rect 26 186 38 226
rect 46 186 58 226
rect 66 186 78 226
<< psubstratepcontact >>
rect -6 -6 106 6
<< nsubstratencontact >>
rect -6 234 106 246
<< polysilicon >>
rect 20 226 24 230
rect 40 226 44 230
rect 60 226 64 230
rect 20 103 24 186
rect 16 91 24 103
rect 20 54 24 91
rect 40 87 44 186
rect 60 182 64 186
rect 60 178 68 182
rect 28 80 44 87
rect 28 54 32 80
rect 64 72 68 178
rect 56 60 68 72
rect 50 34 54 60
rect 20 10 24 14
rect 28 10 32 14
rect 50 10 54 14
<< polycontact >>
rect 4 91 16 103
rect 44 137 56 149
rect 44 60 56 72
<< metal1 >>
rect -6 246 106 248
rect -6 232 106 234
rect 6 226 18 232
rect 46 226 58 232
rect 3 103 17 117
rect 26 72 34 186
rect 43 123 57 137
rect 66 97 74 186
rect 63 83 77 97
rect 10 64 44 72
rect 10 54 18 64
rect 63 42 71 83
rect 56 34 71 42
rect 34 8 46 14
rect -6 6 106 8
rect -6 -8 106 -6
<< m1p >>
rect 43 123 57 137
rect 3 103 17 117
rect 63 83 77 97
<< labels >>
rlabel metal1 -6 -8 106 8 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 -6 232 106 248 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 43 123 57 137 0 B
port 1 nsew signal input
rlabel metal1 3 103 17 117 0 A
port 0 nsew signal input
rlabel metal1 63 83 77 97 0 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 100 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
