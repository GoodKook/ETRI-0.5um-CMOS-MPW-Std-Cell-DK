magic
tech scmos
magscale 1 3
timestamp 1569139307
<< checkpaint >>
rect -70 -108 70 108
<< metal1 >>
rect -10 44 10 48
rect -10 36 -4 44
rect 4 36 10 44
rect -10 28 10 36
rect -10 20 -4 28
rect 4 20 10 28
rect -10 12 10 20
rect -10 4 -4 12
rect 4 4 10 12
rect -10 -4 10 4
rect -10 -12 -4 -4
rect 4 -12 10 -4
rect -10 -20 10 -12
rect -10 -28 -4 -20
rect 4 -28 10 -20
rect -10 -36 10 -28
rect -10 -44 -4 -36
rect 4 -44 10 -36
rect -10 -48 10 -44
<< m2contact >>
rect -4 36 4 44
rect -4 20 4 28
rect -4 4 4 12
rect -4 -12 4 -4
rect -4 -28 4 -20
rect -4 -44 4 -36
<< metal2 >>
rect -10 44 10 48
rect -10 36 -4 44
rect 4 36 10 44
rect -10 28 10 36
rect -10 20 -4 28
rect 4 20 10 28
rect -10 12 10 20
rect -10 4 -4 12
rect 4 4 10 12
rect -10 -4 10 4
rect -10 -12 -4 -4
rect 4 -12 10 -4
rect -10 -20 10 -12
rect -10 -28 -4 -20
rect 4 -28 10 -20
rect -10 -36 10 -28
rect -10 -44 -4 -36
rect 4 -44 10 -36
rect -10 -48 10 -44
<< end >>
