magic
tech scmos
magscale 1 2
timestamp 1728305106
<< nwell >>
rect -12 134 92 252
<< ntransistor >>
rect 21 14 25 34
rect 41 14 45 34
<< ptransistor >>
rect 21 146 25 226
rect 29 146 33 226
<< ndiffusion >>
rect 19 14 21 34
rect 25 14 27 34
rect 39 14 41 34
rect 45 14 47 34
<< pdiffusion >>
rect 19 146 21 226
rect 25 146 29 226
rect 33 146 35 226
<< ndcontact >>
rect 7 14 19 34
rect 27 14 39 34
rect 47 14 59 34
<< pdcontact >>
rect 7 146 19 226
rect 35 146 47 226
<< psubstratepcontact >>
rect -6 -6 86 6
<< nsubstratencontact >>
rect -6 234 86 246
<< polysilicon >>
rect 21 226 25 230
rect 29 226 33 230
rect 21 123 25 146
rect 16 111 25 123
rect 29 123 33 146
rect 29 111 44 123
rect 21 34 25 111
rect 41 34 45 111
rect 21 10 25 14
rect 41 10 45 14
<< polycontact >>
rect 4 111 16 123
rect 44 111 56 123
<< metal1 >>
rect -6 246 86 248
rect -6 232 86 234
rect 7 226 19 232
rect 30 139 47 146
rect 30 91 37 139
rect 30 34 37 77
rect 7 8 19 14
rect 47 8 59 14
rect -6 6 86 8
rect -6 -8 86 -6
<< m2contact >>
rect 3 97 17 111
rect 43 97 57 111
rect 23 77 37 91
<< metal2 >>
rect 3 83 17 97
rect 43 83 57 97
rect 23 63 37 77
<< m1p >>
rect -6 232 86 248
rect -6 -8 86 8
<< m2p >>
rect 3 83 17 97
rect 43 83 57 97
rect 23 63 37 77
<< labels >>
rlabel metal1 -6 -8 86 8 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 -6 232 86 248 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal2 43 83 57 97 0 B
port 1 nsew signal input
rlabel metal2 3 83 17 97 0 A
port 0 nsew signal input
rlabel metal2 23 63 37 77 0 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 80 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
