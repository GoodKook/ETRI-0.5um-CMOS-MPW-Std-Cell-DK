VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fir_pe
  CLASS BLOCK ;
  FOREIGN fir_pe ;
  ORIGIN 6.000 6.000 ;
  SIZE 909.000 BY 912.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 897.300 906.450 899.700 ;
        RECT 16.800 893.400 18.600 897.300 ;
        RECT 29.700 890.400 31.500 897.300 ;
        RECT 44.850 893.400 46.650 897.300 ;
        RECT 53.850 893.400 55.650 897.300 ;
        RECT 60.750 893.400 62.550 897.300 ;
        RECT 70.050 893.400 71.850 897.300 ;
        RECT 80.850 893.400 82.650 897.300 ;
        RECT 89.850 893.400 91.650 897.300 ;
        RECT 96.750 893.400 98.550 897.300 ;
        RECT 106.050 893.400 107.850 897.300 ;
        RECT 122.400 890.400 124.200 897.300 ;
        RECT 128.400 890.400 130.200 897.300 ;
        RECT 134.400 890.400 136.200 897.300 ;
        RECT 140.400 890.400 142.200 897.300 ;
        RECT 146.400 890.400 148.200 897.300 ;
        RECT 164.400 891.300 166.200 897.300 ;
        RECT 173.100 891.300 174.900 897.300 ;
        RECT 199.500 890.400 201.300 897.300 ;
        RECT 220.500 890.400 222.300 897.300 ;
        RECT 238.500 890.400 240.300 897.300 ;
        RECT 247.500 890.400 249.300 897.300 ;
        RECT 271.800 887.400 273.600 897.300 ;
        RECT 289.800 893.400 291.600 897.300 ;
        RECT 313.800 887.400 315.600 897.300 ;
        RECT 331.800 893.400 333.600 897.300 ;
        RECT 347.400 893.400 349.200 897.300 ;
        RECT 353.400 893.400 355.200 897.300 ;
        RECT 371.400 892.200 373.200 897.300 ;
        RECT 403.800 887.400 405.600 897.300 ;
        RECT 416.400 893.400 418.200 897.300 ;
        RECT 448.800 887.400 450.600 897.300 ;
        RECT 462.000 890.400 463.800 897.300 ;
        RECT 469.500 893.400 471.300 897.300 ;
        RECT 488.400 892.200 490.200 897.300 ;
        RECT 509.400 893.400 511.200 897.300 ;
        RECT 528.000 890.400 529.800 897.300 ;
        RECT 535.500 893.400 537.300 897.300 ;
        RECT 557.100 891.300 558.900 897.300 ;
        RECT 565.800 891.300 567.600 897.300 ;
        RECT 584.400 892.200 586.200 897.300 ;
        RECT 616.800 887.400 618.600 897.300 ;
        RECT 637.800 892.200 639.600 897.300 ;
        RECT 664.800 887.400 666.600 897.300 ;
        RECT 677.700 890.400 679.500 897.300 ;
        RECT 701.700 893.400 703.500 897.300 ;
        RECT 709.200 890.400 711.000 897.300 ;
        RECT 733.800 887.400 735.600 897.300 ;
        RECT 757.800 887.400 759.600 897.300 ;
        RECT 771.000 890.400 772.800 897.300 ;
        RECT 778.500 893.400 780.300 897.300 ;
        RECT 799.800 893.400 801.600 897.300 ;
        RECT 812.400 893.400 814.200 897.300 ;
        RECT 831.000 890.400 832.800 897.300 ;
        RECT 838.500 893.400 840.300 897.300 ;
        RECT 857.400 892.200 859.200 897.300 ;
        RECT 878.400 887.400 880.200 897.300 ;
        RECT 15.900 821.700 17.700 828.600 ;
        RECT 35.400 821.700 37.200 825.600 ;
        RECT 47.850 821.700 49.650 825.600 ;
        RECT 56.850 821.700 58.650 825.600 ;
        RECT 63.750 821.700 65.550 825.600 ;
        RECT 73.050 821.700 74.850 825.600 ;
        RECT 92.400 821.700 94.200 827.100 ;
        RECT 119.400 821.700 121.200 827.100 ;
        RECT 143.700 821.700 145.500 828.600 ;
        RECT 167.700 821.700 169.500 828.600 ;
        RECT 191.700 821.700 193.500 825.600 ;
        RECT 199.200 821.700 201.000 828.600 ;
        RECT 212.400 821.700 214.200 831.600 ;
        RECT 237.000 821.700 238.800 828.600 ;
        RECT 244.500 821.700 246.300 825.600 ;
        RECT 268.800 821.700 270.600 826.800 ;
        RECT 287.700 821.700 289.500 825.600 ;
        RECT 295.200 821.700 297.000 828.600 ;
        RECT 309.000 821.700 310.800 828.600 ;
        RECT 316.500 821.700 318.300 825.600 ;
        RECT 340.800 821.700 342.600 826.800 ;
        RECT 359.700 821.700 361.500 825.600 ;
        RECT 367.200 821.700 369.000 828.600 ;
        RECT 380.400 821.700 382.200 831.600 ;
        RECT 407.400 821.700 409.200 826.800 ;
        RECT 439.800 821.700 441.600 831.600 ;
        RECT 463.800 821.700 465.600 831.600 ;
        RECT 484.800 821.700 486.600 826.800 ;
        RECT 503.400 821.700 505.200 826.800 ;
        RECT 527.700 821.700 529.500 825.600 ;
        RECT 535.200 821.700 537.000 828.600 ;
        RECT 559.800 821.700 561.600 831.600 ;
        RECT 577.800 821.700 579.600 827.700 ;
        RECT 586.800 821.700 588.600 827.700 ;
        RECT 602.400 821.700 604.200 831.600 ;
        RECT 629.400 821.700 631.200 826.800 ;
        RECT 658.500 821.700 660.300 828.600 ;
        RECT 679.500 821.700 681.300 828.600 ;
        RECT 692.700 821.700 694.500 828.600 ;
        RECT 720.300 821.700 722.100 828.600 ;
        RECT 748.800 821.700 750.600 831.600 ;
        RECT 762.000 821.700 763.800 828.600 ;
        RECT 769.500 821.700 771.300 825.600 ;
        RECT 788.400 821.700 790.200 826.800 ;
        RECT 809.400 821.700 811.200 831.600 ;
        RECT 841.800 821.700 843.600 826.800 ;
        RECT 863.700 821.700 865.500 825.600 ;
        RECT 871.200 821.700 873.000 828.600 ;
        RECT 897.450 821.700 906.450 897.300 ;
        RECT 0.600 819.300 906.450 821.700 ;
        RECT 11.700 812.400 13.500 819.300 ;
        RECT 32.400 815.400 34.200 819.300 ;
        RECT 58.800 814.200 60.600 819.300 ;
        RECT 69.150 815.400 70.950 819.300 ;
        RECT 78.450 815.400 80.250 819.300 ;
        RECT 85.350 815.400 87.150 819.300 ;
        RECT 94.350 815.400 96.150 819.300 ;
        RECT 110.400 815.400 112.200 819.300 ;
        RECT 131.400 814.200 133.200 819.300 ;
        RECT 157.800 815.400 159.600 819.300 ;
        RECT 178.500 812.400 180.300 819.300 ;
        RECT 196.800 815.400 198.600 819.300 ;
        RECT 223.800 809.400 225.600 819.300 ;
        RECT 241.800 815.400 243.600 819.300 ;
        RECT 257.400 814.200 259.200 819.300 ;
        RECT 289.800 809.400 291.600 819.300 ;
        RECT 303.000 812.400 304.800 819.300 ;
        RECT 310.500 815.400 312.300 819.300 ;
        RECT 337.800 809.400 339.600 819.300 ;
        RECT 355.800 815.400 357.600 819.300 ;
        RECT 379.800 809.400 381.600 819.300 ;
        RECT 400.800 814.200 402.600 819.300 ;
        RECT 424.500 812.400 426.300 819.300 ;
        RECT 448.800 809.400 450.600 819.300 ;
        RECT 464.700 815.400 466.500 819.300 ;
        RECT 472.200 812.400 474.000 819.300 ;
        RECT 492.300 812.400 494.100 819.300 ;
        RECT 517.500 812.400 519.300 819.300 ;
        RECT 538.800 815.400 540.600 819.300 ;
        RECT 552.000 812.400 553.800 819.300 ;
        RECT 559.500 815.400 561.300 819.300 ;
        RECT 583.800 814.200 585.600 819.300 ;
        RECT 602.400 814.200 604.200 819.300 ;
        RECT 637.800 809.400 639.600 819.300 ;
        RECT 661.800 809.400 663.600 819.300 ;
        RECT 675.000 812.400 676.800 819.300 ;
        RECT 682.500 815.400 684.300 819.300 ;
        RECT 701.400 814.200 703.200 819.300 ;
        RECT 730.800 814.200 732.600 819.300 ;
        RECT 746.400 809.400 748.200 819.300 ;
        RECT 778.800 814.200 780.600 819.300 ;
        RECT 805.800 809.400 807.600 819.300 ;
        RECT 819.000 812.400 820.800 819.300 ;
        RECT 826.500 815.400 828.300 819.300 ;
        RECT 845.700 815.400 847.500 819.300 ;
        RECT 853.200 812.400 855.000 819.300 ;
        RECT 877.800 809.400 879.600 819.300 ;
        RECT 16.800 743.700 18.600 747.600 ;
        RECT 29.700 743.700 31.500 750.600 ;
        RECT 53.400 743.700 55.200 748.800 ;
        RECT 74.700 743.700 76.500 750.600 ;
        RECT 95.400 743.700 97.200 747.600 ;
        RECT 101.400 743.700 103.200 747.600 ;
        RECT 116.400 743.700 118.200 747.600 ;
        RECT 122.400 743.700 124.200 747.600 ;
        RECT 137.400 743.700 139.200 747.600 ;
        RECT 143.400 743.700 145.200 747.600 ;
        RECT 158.400 743.700 160.200 747.600 ;
        RECT 179.400 743.700 181.200 749.100 ;
        RECT 214.800 743.700 216.600 753.600 ;
        RECT 238.800 743.700 240.600 753.600 ;
        RECT 265.800 743.700 267.600 753.600 ;
        RECT 281.700 743.700 283.500 747.600 ;
        RECT 289.200 743.700 291.000 750.600 ;
        RECT 302.400 743.700 304.200 753.600 ;
        RECT 326.700 743.700 328.500 750.600 ;
        RECT 352.800 743.700 354.600 747.600 ;
        RECT 373.800 743.700 375.600 748.800 ;
        RECT 397.800 743.700 399.600 747.600 ;
        RECT 410.700 743.700 412.500 750.600 ;
        RECT 442.800 743.700 444.600 749.100 ;
        RECT 458.400 743.700 460.200 747.600 ;
        RECT 464.400 743.700 466.200 747.600 ;
        RECT 482.400 743.700 484.200 748.800 ;
        RECT 506.400 743.700 508.200 753.600 ;
        RECT 535.800 743.700 537.600 747.600 ;
        RECT 548.400 743.700 550.200 753.600 ;
        RECT 580.800 743.700 582.600 748.800 ;
        RECT 596.700 743.700 598.500 750.600 ;
        RECT 617.400 743.700 619.200 753.600 ;
        RECT 646.800 743.700 648.600 747.600 ;
        RECT 664.800 743.700 666.600 747.600 ;
        RECT 677.400 743.700 679.200 753.600 ;
        RECT 712.800 743.700 714.600 753.600 ;
        RECT 726.000 743.700 727.800 750.600 ;
        RECT 733.500 743.700 735.300 747.600 ;
        RECT 749.700 743.700 751.500 750.600 ;
        RECT 778.500 743.700 780.300 750.600 ;
        RECT 795.900 743.700 797.700 750.600 ;
        RECT 816.000 743.700 817.800 750.600 ;
        RECT 823.500 743.700 825.300 747.600 ;
        RECT 847.800 743.700 849.600 747.600 ;
        RECT 860.400 743.700 862.200 753.600 ;
        RECT 897.450 743.700 906.450 819.300 ;
        RECT 0.600 741.300 906.450 743.700 ;
        RECT 11.700 734.400 13.500 741.300 ;
        RECT 32.400 737.400 34.200 741.300 ;
        RECT 55.800 737.400 57.600 741.300 ;
        RECT 76.800 736.200 78.600 741.300 ;
        RECT 97.800 737.400 99.600 741.300 ;
        RECT 104.850 737.400 106.650 741.300 ;
        RECT 113.850 737.400 115.650 741.300 ;
        RECT 120.750 737.400 122.550 741.300 ;
        RECT 130.050 737.400 131.850 741.300 ;
        RECT 154.800 736.200 156.600 741.300 ;
        RECT 164.850 737.400 166.650 741.300 ;
        RECT 173.850 737.400 175.650 741.300 ;
        RECT 180.750 737.400 182.550 741.300 ;
        RECT 190.050 737.400 191.850 741.300 ;
        RECT 209.700 737.400 211.500 741.300 ;
        RECT 217.200 734.400 219.000 741.300 ;
        RECT 238.800 736.200 240.600 741.300 ;
        RECT 257.400 736.200 259.200 741.300 ;
        RECT 281.700 737.400 283.500 741.300 ;
        RECT 289.200 734.400 291.000 741.300 ;
        RECT 313.800 731.400 315.600 741.300 ;
        RECT 326.400 737.400 328.200 741.300 ;
        RECT 345.000 734.400 346.800 741.300 ;
        RECT 352.500 737.400 354.300 741.300 ;
        RECT 371.400 736.200 373.200 741.300 ;
        RECT 392.400 737.400 394.200 741.300 ;
        RECT 398.400 737.400 400.200 741.300 ;
        RECT 413.700 734.400 415.500 741.300 ;
        RECT 439.800 737.400 441.600 741.300 ;
        RECT 463.800 736.200 465.600 741.300 ;
        RECT 484.800 737.400 486.600 741.300 ;
        RECT 505.500 734.400 507.300 741.300 ;
        RECT 518.700 734.400 520.500 741.300 ;
        RECT 539.700 734.400 541.500 741.300 ;
        RECT 560.700 734.400 562.500 741.300 ;
        RECT 588.300 734.400 590.100 741.300 ;
        RECT 608.400 736.200 610.200 741.300 ;
        RECT 636.300 734.400 638.100 741.300 ;
        RECT 653.700 734.400 655.500 741.300 ;
        RECT 677.700 737.400 679.500 741.300 ;
        RECT 685.200 734.400 687.000 741.300 ;
        RECT 698.400 731.400 700.200 741.300 ;
        RECT 730.800 736.200 732.600 741.300 ;
        RECT 746.700 734.400 748.500 741.300 ;
        RECT 767.400 737.400 769.200 741.300 ;
        RECT 796.800 731.400 798.600 741.300 ;
        RECT 810.000 734.400 811.800 741.300 ;
        RECT 817.500 737.400 819.300 741.300 ;
        RECT 836.400 731.400 838.200 741.300 ;
        RECT 863.400 736.200 865.200 741.300 ;
        RECT 19.800 665.700 21.600 670.800 ;
        RECT 38.400 665.700 40.200 670.800 ;
        RECT 66.300 665.700 68.100 672.600 ;
        RECT 91.800 665.700 93.600 669.600 ;
        RECT 97.800 666.600 99.600 669.600 ;
        RECT 98.400 665.700 99.600 666.600 ;
        RECT 110.700 665.700 112.500 672.600 ;
        RECT 131.700 665.700 133.500 672.600 ;
        RECT 157.800 665.700 159.600 669.600 ;
        RECT 178.800 665.700 180.600 669.600 ;
        RECT 202.800 665.700 204.600 675.600 ;
        RECT 216.000 665.700 217.800 672.600 ;
        RECT 223.500 665.700 225.300 669.600 ;
        RECT 247.800 665.700 249.600 670.800 ;
        RECT 266.700 665.700 268.500 669.600 ;
        RECT 274.200 665.700 276.000 672.600 ;
        RECT 295.500 665.700 297.300 672.600 ;
        RECT 316.500 665.700 318.300 672.600 ;
        RECT 336.300 665.700 338.100 672.600 ;
        RECT 358.500 665.700 360.300 672.600 ;
        RECT 367.500 665.700 369.300 672.600 ;
        RECT 388.500 665.700 390.300 672.600 ;
        RECT 409.800 665.700 411.600 670.800 ;
        RECT 430.500 665.700 432.300 672.600 ;
        RECT 439.500 665.700 441.300 672.600 ;
        RECT 458.400 665.700 460.200 670.800 ;
        RECT 482.400 665.700 484.200 670.800 ;
        RECT 510.300 665.700 512.100 672.600 ;
        RECT 530.400 665.700 532.200 670.800 ;
        RECT 551.700 665.700 553.500 672.600 ;
        RECT 575.400 665.700 577.200 670.800 ;
        RECT 599.400 665.700 601.200 670.800 ;
        RECT 627.300 665.700 629.100 672.600 ;
        RECT 644.400 665.700 646.200 669.600 ;
        RECT 650.400 665.700 652.200 669.600 ;
        RECT 671.700 665.700 673.500 669.600 ;
        RECT 679.200 665.700 681.000 672.600 ;
        RECT 703.800 665.700 705.600 675.600 ;
        RECT 724.800 665.700 726.600 670.800 ;
        RECT 743.400 665.700 745.200 670.800 ;
        RECT 775.800 665.700 777.600 675.600 ;
        RECT 789.000 665.700 790.800 672.600 ;
        RECT 796.500 665.700 798.300 669.600 ;
        RECT 815.400 665.700 817.200 670.800 ;
        RECT 839.700 665.700 841.500 669.600 ;
        RECT 847.200 665.700 849.000 672.600 ;
        RECT 860.400 665.700 862.200 675.600 ;
        RECT 887.400 665.700 889.200 669.600 ;
        RECT 897.450 665.700 906.450 741.300 ;
        RECT 0.600 663.300 906.450 665.700 ;
        RECT 13.800 659.400 15.600 663.300 ;
        RECT 19.800 659.400 21.600 663.300 ;
        RECT 32.400 659.400 34.200 663.300 ;
        RECT 53.400 658.200 55.200 663.300 ;
        RECT 76.800 659.400 78.600 663.300 ;
        RECT 82.800 659.400 84.600 663.300 ;
        RECT 98.400 653.400 100.200 663.300 ;
        RECT 127.800 659.400 129.600 663.300 ;
        RECT 134.850 659.400 136.650 663.300 ;
        RECT 143.850 659.400 145.650 663.300 ;
        RECT 150.750 659.400 152.550 663.300 ;
        RECT 160.050 659.400 161.850 663.300 ;
        RECT 179.400 658.200 181.200 663.300 ;
        RECT 205.800 659.400 207.600 663.300 ;
        RECT 226.800 658.200 228.600 663.300 ;
        RECT 245.700 659.400 247.500 663.300 ;
        RECT 253.200 656.400 255.000 663.300 ;
        RECT 266.400 653.400 268.200 663.300 ;
        RECT 301.800 658.200 303.600 663.300 ;
        RECT 317.400 659.400 319.200 663.300 ;
        RECT 323.400 659.400 325.200 663.300 ;
        RECT 338.700 656.400 340.500 663.300 ;
        RECT 366.300 656.400 368.100 663.300 ;
        RECT 391.800 658.200 393.600 663.300 ;
        RECT 407.700 656.400 409.500 663.300 ;
        RECT 428.700 656.400 430.500 663.300 ;
        RECT 457.800 658.200 459.600 663.300 ;
        RECT 481.500 656.400 483.300 663.300 ;
        RECT 498.900 656.400 500.700 663.300 ;
        RECT 518.700 656.400 520.500 663.300 ;
        RECT 539.400 656.400 541.200 663.300 ;
        RECT 562.800 656.400 564.600 663.300 ;
        RECT 583.800 658.200 585.600 663.300 ;
        RECT 604.800 659.400 606.600 663.300 ;
        RECT 631.800 653.400 633.600 663.300 ;
        RECT 652.500 656.400 654.300 663.300 ;
        RECT 665.700 656.400 667.500 663.300 ;
        RECT 691.500 656.400 693.300 663.300 ;
        RECT 700.500 656.400 702.300 663.300 ;
        RECT 713.700 656.400 715.500 663.300 ;
        RECT 722.700 656.400 724.500 663.300 ;
        RECT 743.700 659.400 745.500 663.300 ;
        RECT 751.200 656.400 753.000 663.300 ;
        RECT 764.400 653.400 766.200 663.300 ;
        RECT 788.400 653.400 790.200 663.300 ;
        RECT 815.400 659.400 817.200 663.300 ;
        RECT 834.000 656.400 835.800 663.300 ;
        RECT 841.500 659.400 843.300 663.300 ;
        RECT 868.800 653.400 870.600 663.300 ;
        RECT 882.000 656.400 883.800 663.300 ;
        RECT 889.500 659.400 891.300 663.300 ;
        RECT 18.300 587.700 20.100 594.600 ;
        RECT 41.100 587.700 42.900 593.700 ;
        RECT 49.800 587.700 51.600 593.700 ;
        RECT 70.800 587.700 72.600 593.700 ;
        RECT 79.800 587.700 81.600 593.700 ;
        RECT 96.000 587.700 97.800 594.600 ;
        RECT 103.500 587.700 105.300 591.600 ;
        RECT 119.700 587.700 121.500 594.600 ;
        RECT 142.800 587.700 144.600 591.600 ;
        RECT 148.800 587.700 150.600 591.600 ;
        RECT 166.800 587.700 168.600 591.600 ;
        RECT 184.800 587.700 186.600 591.600 ;
        RECT 190.800 587.700 192.600 591.600 ;
        RECT 198.150 587.700 199.950 591.600 ;
        RECT 207.450 587.700 209.250 591.600 ;
        RECT 214.350 587.700 216.150 591.600 ;
        RECT 223.350 587.700 225.150 591.600 ;
        RECT 247.800 587.700 249.600 592.800 ;
        RECT 266.400 587.700 268.200 593.700 ;
        RECT 275.100 587.700 276.900 593.700 ;
        RECT 293.400 587.700 295.200 591.600 ;
        RECT 299.400 587.700 301.200 591.600 ;
        RECT 322.500 587.700 324.300 594.600 ;
        RECT 342.300 587.700 344.100 594.600 ;
        RECT 359.700 587.700 361.500 594.600 ;
        RECT 380.700 587.700 382.500 594.600 ;
        RECT 389.700 587.700 391.500 594.600 ;
        RECT 412.800 587.700 414.600 591.600 ;
        RECT 433.800 587.700 435.600 591.600 ;
        RECT 454.800 587.700 456.600 591.600 ;
        RECT 478.800 587.700 480.600 592.800 ;
        RECT 489.150 587.700 490.950 591.600 ;
        RECT 498.450 587.700 500.250 591.600 ;
        RECT 505.350 587.700 507.150 591.600 ;
        RECT 514.350 587.700 516.150 591.600 ;
        RECT 541.800 587.700 543.600 592.800 ;
        RECT 552.150 587.700 553.950 591.600 ;
        RECT 561.450 587.700 563.250 591.600 ;
        RECT 568.350 587.700 570.150 591.600 ;
        RECT 577.350 587.700 579.150 591.600 ;
        RECT 601.500 587.700 603.300 594.600 ;
        RECT 622.800 587.700 624.600 592.800 ;
        RECT 646.500 587.700 648.300 594.600 ;
        RECT 662.400 587.700 664.200 592.800 ;
        RECT 686.400 587.700 688.200 591.600 ;
        RECT 707.400 587.700 709.200 591.600 ;
        RECT 725.700 587.700 727.500 594.600 ;
        RECT 746.400 587.700 748.200 597.600 ;
        RECT 770.700 587.700 772.500 594.600 ;
        RECT 779.700 587.700 781.500 594.600 ;
        RECT 797.400 587.700 799.200 591.600 ;
        RECT 823.800 587.700 825.600 592.800 ;
        RECT 839.400 587.700 841.200 597.600 ;
        RECT 866.700 587.700 868.500 591.600 ;
        RECT 874.200 587.700 876.000 594.600 ;
        RECT 892.800 587.700 894.600 591.600 ;
        RECT 897.450 587.700 906.450 663.300 ;
        RECT 0.600 585.300 906.450 587.700 ;
        RECT 13.800 581.400 15.600 585.300 ;
        RECT 19.800 581.400 21.600 585.300 ;
        RECT 40.500 578.400 42.300 585.300 ;
        RECT 64.800 580.200 66.600 585.300 ;
        RECT 83.400 580.200 85.200 585.300 ;
        RECT 107.400 581.400 109.200 585.300 ;
        RECT 125.700 578.400 127.500 585.300 ;
        RECT 149.400 580.200 151.200 585.300 ;
        RECT 175.800 581.400 177.600 585.300 ;
        RECT 188.700 578.400 190.500 585.300 ;
        RECT 203.850 581.400 205.650 585.300 ;
        RECT 212.850 581.400 214.650 585.300 ;
        RECT 219.750 581.400 221.550 585.300 ;
        RECT 229.050 581.400 230.850 585.300 ;
        RECT 245.700 578.400 247.500 585.300 ;
        RECT 266.700 578.400 268.500 585.300 ;
        RECT 287.400 578.400 289.200 585.300 ;
        RECT 293.400 578.400 295.200 585.300 ;
        RECT 299.400 578.400 301.200 585.300 ;
        RECT 305.400 578.400 307.200 585.300 ;
        RECT 311.400 578.400 313.200 585.300 ;
        RECT 326.400 575.400 328.200 585.300 ;
        RECT 350.400 578.400 352.200 585.300 ;
        RECT 356.400 578.400 358.200 585.300 ;
        RECT 362.400 578.400 364.200 585.300 ;
        RECT 368.400 578.400 370.200 585.300 ;
        RECT 374.400 578.400 376.200 585.300 ;
        RECT 394.800 581.400 396.600 585.300 ;
        RECT 412.800 581.400 414.600 585.300 ;
        RECT 433.800 581.400 435.600 585.300 ;
        RECT 446.700 578.400 448.500 585.300 ;
        RECT 475.500 578.400 477.300 585.300 ;
        RECT 496.500 578.400 498.300 585.300 ;
        RECT 509.700 578.400 511.500 585.300 ;
        RECT 538.800 580.200 540.600 585.300 ;
        RECT 549.150 581.400 550.950 585.300 ;
        RECT 558.450 581.400 560.250 585.300 ;
        RECT 565.350 581.400 567.150 585.300 ;
        RECT 574.350 581.400 576.150 585.300 ;
        RECT 590.400 581.400 592.200 585.300 ;
        RECT 608.400 578.400 610.200 585.300 ;
        RECT 634.500 578.400 636.300 585.300 ;
        RECT 650.400 581.400 652.200 585.300 ;
        RECT 675.300 578.400 677.100 585.300 ;
        RECT 700.500 578.400 702.300 585.300 ;
        RECT 716.400 580.200 718.200 585.300 ;
        RECT 745.500 578.400 747.300 585.300 ;
        RECT 758.400 575.400 760.200 585.300 ;
        RECT 785.700 578.400 787.500 585.300 ;
        RECT 794.700 578.400 796.500 585.300 ;
        RECT 820.800 580.200 822.600 585.300 ;
        RECT 839.400 580.200 841.200 585.300 ;
        RECT 860.400 575.400 862.200 585.300 ;
        RECT 14.400 509.700 16.200 514.800 ;
        RECT 43.500 509.700 45.300 516.600 ;
        RECT 61.800 509.700 63.600 515.700 ;
        RECT 70.800 509.700 72.600 515.700 ;
        RECT 80.850 509.700 82.650 513.600 ;
        RECT 89.850 509.700 91.650 513.600 ;
        RECT 96.750 509.700 98.550 513.600 ;
        RECT 106.050 509.700 107.850 513.600 ;
        RECT 125.400 509.700 127.200 514.800 ;
        RECT 146.700 509.700 148.500 516.600 ;
        RECT 161.850 509.700 163.650 513.600 ;
        RECT 170.850 509.700 172.650 513.600 ;
        RECT 177.750 509.700 179.550 513.600 ;
        RECT 187.050 509.700 188.850 513.600 ;
        RECT 203.400 509.700 205.200 513.600 ;
        RECT 224.400 509.700 226.200 514.800 ;
        RECT 251.400 509.700 253.200 513.600 ;
        RECT 269.700 509.700 271.500 516.600 ;
        RECT 290.400 509.700 292.200 513.600 ;
        RECT 310.800 509.700 312.600 513.600 ;
        RECT 316.800 509.700 318.600 513.600 ;
        RECT 323.850 509.700 325.650 513.600 ;
        RECT 332.850 509.700 334.650 513.600 ;
        RECT 339.750 509.700 341.550 513.600 ;
        RECT 349.050 509.700 350.850 513.600 ;
        RECT 373.500 509.700 375.300 516.600 ;
        RECT 391.800 509.700 393.600 516.600 ;
        RECT 412.800 509.700 414.600 514.800 ;
        RECT 423.150 509.700 424.950 513.600 ;
        RECT 432.450 509.700 434.250 513.600 ;
        RECT 439.350 509.700 441.150 513.600 ;
        RECT 448.350 509.700 450.150 513.600 ;
        RECT 464.700 509.700 466.500 516.600 ;
        RECT 493.500 509.700 495.300 516.600 ;
        RECT 514.800 509.700 516.600 514.800 ;
        RECT 525.150 509.700 526.950 513.600 ;
        RECT 534.450 509.700 536.250 513.600 ;
        RECT 541.350 509.700 543.150 513.600 ;
        RECT 550.350 509.700 552.150 513.600 ;
        RECT 569.400 509.700 571.200 514.800 ;
        RECT 597.300 509.700 599.100 516.600 ;
        RECT 625.800 509.700 627.600 519.600 ;
        RECT 638.400 509.700 640.200 513.600 ;
        RECT 664.500 509.700 666.300 516.600 ;
        RECT 680.400 509.700 682.200 514.800 ;
        RECT 704.400 509.700 706.200 513.600 ;
        RECT 725.400 509.700 727.200 514.800 ;
        RECT 750.900 509.700 752.700 516.600 ;
        RECT 778.500 509.700 780.300 516.600 ;
        RECT 799.500 509.700 801.300 516.600 ;
        RECT 816.900 509.700 818.700 516.600 ;
        RECT 839.700 509.700 841.500 513.600 ;
        RECT 847.200 509.700 849.000 516.600 ;
        RECT 863.400 509.700 865.200 514.800 ;
        RECT 897.450 509.700 906.450 585.300 ;
        RECT 0.600 507.300 906.450 509.700 ;
        RECT 6.150 503.400 7.950 507.300 ;
        RECT 15.450 503.400 17.250 507.300 ;
        RECT 22.350 503.400 24.150 507.300 ;
        RECT 31.350 503.400 33.150 507.300 ;
        RECT 47.700 500.400 49.500 507.300 ;
        RECT 76.500 500.400 78.300 507.300 ;
        RECT 83.850 503.400 85.650 507.300 ;
        RECT 92.850 503.400 94.650 507.300 ;
        RECT 99.750 503.400 101.550 507.300 ;
        RECT 109.050 503.400 110.850 507.300 ;
        RECT 128.700 503.400 130.500 507.300 ;
        RECT 136.200 500.400 138.000 507.300 ;
        RECT 149.400 503.400 151.200 507.300 ;
        RECT 155.400 503.400 157.200 507.300 ;
        RECT 170.400 503.400 172.200 507.300 ;
        RECT 191.700 500.400 193.500 507.300 ;
        RECT 219.300 500.400 221.100 507.300 ;
        RECT 236.700 500.400 238.500 507.300 ;
        RECT 265.800 502.200 267.600 507.300 ;
        RECT 275.850 503.400 277.650 507.300 ;
        RECT 284.850 503.400 286.650 507.300 ;
        RECT 291.750 503.400 293.550 507.300 ;
        RECT 301.050 503.400 302.850 507.300 ;
        RECT 320.400 502.200 322.200 507.300 ;
        RECT 349.800 502.200 351.600 507.300 ;
        RECT 359.850 503.400 361.650 507.300 ;
        RECT 368.850 503.400 370.650 507.300 ;
        RECT 375.750 503.400 377.550 507.300 ;
        RECT 385.050 503.400 386.850 507.300 ;
        RECT 409.500 500.400 411.300 507.300 ;
        RECT 430.800 502.200 432.600 507.300 ;
        RECT 454.800 502.200 456.600 507.300 ;
        RECT 465.150 503.400 466.950 507.300 ;
        RECT 474.450 503.400 476.250 507.300 ;
        RECT 481.350 503.400 483.150 507.300 ;
        RECT 490.350 503.400 492.150 507.300 ;
        RECT 509.400 502.200 511.200 507.300 ;
        RECT 530.400 500.400 532.200 507.300 ;
        RECT 551.400 503.400 553.200 507.300 ;
        RECT 577.500 500.400 579.300 507.300 ;
        RECT 598.800 502.200 600.600 507.300 ;
        RECT 617.400 502.200 619.200 507.300 ;
        RECT 638.700 500.400 640.500 507.300 ;
        RECT 659.400 497.400 661.200 507.300 ;
        RECT 683.700 500.400 685.500 507.300 ;
        RECT 710.400 502.200 712.200 507.300 ;
        RECT 732.000 500.400 733.800 507.300 ;
        RECT 739.500 503.400 741.300 507.300 ;
        RECT 762.300 500.400 764.100 507.300 ;
        RECT 779.700 500.400 781.500 507.300 ;
        RECT 788.700 500.400 790.500 507.300 ;
        RECT 806.400 503.400 808.200 507.300 ;
        RECT 812.400 503.400 814.200 507.300 ;
        RECT 827.700 500.400 829.500 507.300 ;
        RECT 856.800 502.200 858.600 507.300 ;
        RECT 872.400 497.400 874.200 507.300 ;
        RECT 6.150 431.700 7.950 435.600 ;
        RECT 15.450 431.700 17.250 435.600 ;
        RECT 22.350 431.700 24.150 435.600 ;
        RECT 31.350 431.700 33.150 435.600 ;
        RECT 55.800 431.700 57.600 436.800 ;
        RECT 76.800 431.700 78.600 435.600 ;
        RECT 95.400 431.700 97.200 437.700 ;
        RECT 104.100 431.700 105.900 437.700 ;
        RECT 127.800 431.700 129.600 437.700 ;
        RECT 136.800 431.700 138.600 437.700 ;
        RECT 157.800 431.700 159.600 435.600 ;
        RECT 173.400 431.700 175.200 435.600 ;
        RECT 199.800 431.700 201.600 436.800 ;
        RECT 215.700 431.700 217.500 438.600 ;
        RECT 230.850 431.700 232.650 435.600 ;
        RECT 239.850 431.700 241.650 435.600 ;
        RECT 246.750 431.700 248.550 435.600 ;
        RECT 256.050 431.700 257.850 435.600 ;
        RECT 272.700 431.700 274.500 438.600 ;
        RECT 287.850 431.700 289.650 435.600 ;
        RECT 296.850 431.700 298.650 435.600 ;
        RECT 303.750 431.700 305.550 435.600 ;
        RECT 313.050 431.700 314.850 435.600 ;
        RECT 337.800 431.700 339.600 436.800 ;
        RECT 361.800 431.700 363.600 436.800 ;
        RECT 379.800 431.700 381.600 435.600 ;
        RECT 385.800 431.700 387.600 435.600 ;
        RECT 392.850 431.700 394.650 435.600 ;
        RECT 401.850 431.700 403.650 435.600 ;
        RECT 408.750 431.700 410.550 435.600 ;
        RECT 418.050 431.700 419.850 435.600 ;
        RECT 439.800 431.700 441.600 435.600 ;
        RECT 449.850 431.700 451.650 435.600 ;
        RECT 458.850 431.700 460.650 435.600 ;
        RECT 465.750 431.700 467.550 435.600 ;
        RECT 475.050 431.700 476.850 435.600 ;
        RECT 494.400 431.700 496.200 435.600 ;
        RECT 512.400 431.700 514.200 438.600 ;
        RECT 538.500 431.700 540.300 438.600 ;
        RECT 559.800 431.700 561.600 438.600 ;
        RECT 577.800 431.700 579.600 438.600 ;
        RECT 590.700 431.700 592.500 438.600 ;
        RECT 613.800 431.700 615.600 435.600 ;
        RECT 619.800 431.700 621.600 435.600 ;
        RECT 636.900 431.700 638.700 438.600 ;
        RECT 661.500 431.700 663.300 438.600 ;
        RECT 670.500 431.700 672.300 438.600 ;
        RECT 691.500 431.700 693.300 438.600 ;
        RECT 707.400 431.700 709.200 436.800 ;
        RECT 728.700 431.700 730.500 438.600 ;
        RECT 757.500 431.700 759.300 438.600 ;
        RECT 778.500 431.700 780.300 438.600 ;
        RECT 796.800 431.700 798.600 437.700 ;
        RECT 805.800 431.700 807.600 437.700 ;
        RECT 824.400 431.700 826.200 436.800 ;
        RECT 850.800 431.700 852.600 435.600 ;
        RECT 863.400 431.700 865.200 435.600 ;
        RECT 882.000 431.700 883.800 438.600 ;
        RECT 889.500 431.700 891.300 435.600 ;
        RECT 897.450 431.700 906.450 507.300 ;
        RECT 0.600 429.300 906.450 431.700 ;
        RECT 6.150 425.400 7.950 429.300 ;
        RECT 15.450 425.400 17.250 429.300 ;
        RECT 22.350 425.400 24.150 429.300 ;
        RECT 31.350 425.400 33.150 429.300 ;
        RECT 47.700 422.400 49.500 429.300 ;
        RECT 71.400 424.200 73.200 429.300 ;
        RECT 100.800 424.200 102.600 429.300 ;
        RECT 119.700 422.400 121.500 429.300 ;
        RECT 135.150 425.400 136.950 429.300 ;
        RECT 144.450 425.400 146.250 429.300 ;
        RECT 151.350 425.400 153.150 429.300 ;
        RECT 160.350 425.400 162.150 429.300 ;
        RECT 184.800 424.200 186.600 429.300 ;
        RECT 202.800 425.400 204.600 429.300 ;
        RECT 208.800 425.400 210.600 429.300 ;
        RECT 226.800 425.400 228.600 429.300 ;
        RECT 244.800 425.400 246.600 429.300 ;
        RECT 251.850 425.400 253.650 429.300 ;
        RECT 260.850 425.400 262.650 429.300 ;
        RECT 267.750 425.400 269.550 429.300 ;
        RECT 277.050 425.400 278.850 429.300 ;
        RECT 293.700 422.400 295.500 429.300 ;
        RECT 317.400 424.200 319.200 429.300 ;
        RECT 349.800 424.200 351.600 429.300 ;
        RECT 368.400 424.200 370.200 429.300 ;
        RECT 390.000 422.400 391.800 429.300 ;
        RECT 397.500 425.400 399.300 429.300 ;
        RECT 421.800 424.200 423.600 429.300 ;
        RECT 432.150 425.400 433.950 429.300 ;
        RECT 441.450 425.400 443.250 429.300 ;
        RECT 448.350 425.400 450.150 429.300 ;
        RECT 457.350 425.400 459.150 429.300 ;
        RECT 478.800 425.400 480.600 429.300 ;
        RECT 494.700 422.400 496.500 429.300 ;
        RECT 523.800 424.200 525.600 429.300 ;
        RECT 542.400 424.200 544.200 429.300 ;
        RECT 563.400 425.400 565.200 429.300 ;
        RECT 569.400 425.400 571.200 429.300 ;
        RECT 592.800 424.200 594.600 429.300 ;
        RECT 608.700 422.400 610.500 429.300 ;
        RECT 629.400 425.400 631.200 429.300 ;
        RECT 635.400 425.400 637.200 429.300 ;
        RECT 650.700 422.400 652.500 429.300 ;
        RECT 672.000 422.400 673.800 429.300 ;
        RECT 679.500 425.400 681.300 429.300 ;
        RECT 695.700 422.400 697.500 429.300 ;
        RECT 704.700 422.400 706.500 429.300 ;
        RECT 729.300 422.400 731.100 429.300 ;
        RECT 754.800 424.200 756.600 429.300 ;
        RECT 770.700 422.400 772.500 429.300 ;
        RECT 791.400 428.400 792.600 429.300 ;
        RECT 791.400 425.400 793.200 428.400 ;
        RECT 797.400 425.400 799.200 429.300 ;
        RECT 823.800 424.200 825.600 429.300 ;
        RECT 839.400 425.400 841.200 429.300 ;
        RECT 845.400 425.400 847.200 429.300 ;
        RECT 863.400 424.200 865.200 429.300 ;
        RECT 884.700 422.400 886.500 429.300 ;
        RECT 6.150 353.700 7.950 357.600 ;
        RECT 15.450 353.700 17.250 357.600 ;
        RECT 22.350 353.700 24.150 357.600 ;
        RECT 31.350 353.700 33.150 357.600 ;
        RECT 55.800 353.700 57.600 358.800 ;
        RECT 79.500 353.700 81.300 360.600 ;
        RECT 86.850 353.700 88.650 357.600 ;
        RECT 95.850 353.700 97.650 357.600 ;
        RECT 102.750 353.700 104.550 357.600 ;
        RECT 112.050 353.700 113.850 357.600 ;
        RECT 133.800 353.700 135.600 357.600 ;
        RECT 151.800 353.700 153.600 357.600 ;
        RECT 157.800 353.700 159.600 357.600 ;
        RECT 173.400 353.700 175.200 358.800 ;
        RECT 196.800 353.700 198.600 357.600 ;
        RECT 202.800 353.700 204.600 357.600 ;
        RECT 209.850 353.700 211.650 357.600 ;
        RECT 218.850 353.700 220.650 357.600 ;
        RECT 225.750 353.700 227.550 357.600 ;
        RECT 235.050 353.700 236.850 357.600 ;
        RECT 254.400 353.700 256.200 358.800 ;
        RECT 278.700 353.700 280.500 360.600 ;
        RECT 299.400 353.700 301.200 360.600 ;
        RECT 325.800 353.700 327.600 357.600 ;
        RECT 341.400 353.700 343.200 358.800 ;
        RECT 356.850 353.700 358.650 357.600 ;
        RECT 365.850 353.700 367.650 357.600 ;
        RECT 372.750 353.700 374.550 357.600 ;
        RECT 382.050 353.700 383.850 357.600 ;
        RECT 392.850 353.700 394.650 357.600 ;
        RECT 401.850 353.700 403.650 357.600 ;
        RECT 408.750 353.700 410.550 357.600 ;
        RECT 418.050 353.700 419.850 357.600 ;
        RECT 429.150 353.700 430.950 357.600 ;
        RECT 438.450 353.700 440.250 357.600 ;
        RECT 445.350 353.700 447.150 357.600 ;
        RECT 454.350 353.700 456.150 357.600 ;
        RECT 470.400 353.700 472.200 357.600 ;
        RECT 476.400 353.700 478.200 357.600 ;
        RECT 495.000 353.700 496.800 360.600 ;
        RECT 502.500 353.700 504.300 357.600 ;
        RECT 526.800 353.700 528.600 357.600 ;
        RECT 532.800 354.600 534.600 357.600 ;
        RECT 533.400 353.700 534.600 354.600 ;
        RECT 551.400 353.700 553.200 358.800 ;
        RECT 575.400 353.700 577.200 358.800 ;
        RECT 599.400 353.700 601.200 359.100 ;
        RECT 623.400 353.700 625.200 357.600 ;
        RECT 649.800 353.700 651.600 358.800 ;
        RECT 665.700 353.700 667.500 360.600 ;
        RECT 692.400 353.700 694.200 359.700 ;
        RECT 701.100 353.700 702.900 359.700 ;
        RECT 727.800 353.700 729.600 358.800 ;
        RECT 743.400 353.700 745.200 357.600 ;
        RECT 749.400 353.700 751.200 357.600 ;
        RECT 767.400 353.700 769.200 359.700 ;
        RECT 776.400 353.700 778.200 359.700 ;
        RECT 802.800 353.700 804.600 358.800 ;
        RECT 818.700 353.700 820.500 360.600 ;
        RECT 842.400 353.700 844.200 358.800 ;
        RECT 864.000 353.700 865.800 360.600 ;
        RECT 871.500 353.700 873.300 357.600 ;
        RECT 897.450 353.700 906.450 429.300 ;
        RECT 0.600 351.300 906.450 353.700 ;
        RECT 6.150 347.400 7.950 351.300 ;
        RECT 15.450 347.400 17.250 351.300 ;
        RECT 22.350 347.400 24.150 351.300 ;
        RECT 31.350 347.400 33.150 351.300 ;
        RECT 47.700 344.400 49.500 351.300 ;
        RECT 76.500 344.400 78.300 351.300 ;
        RECT 85.500 344.400 87.300 351.300 ;
        RECT 101.700 344.400 103.500 351.300 ;
        RECT 130.800 346.200 132.600 351.300 ;
        RECT 154.500 344.400 156.300 351.300 ;
        RECT 175.500 344.400 177.300 351.300 ;
        RECT 188.400 347.400 190.200 351.300 ;
        RECT 209.400 347.400 211.200 351.300 ;
        RECT 229.800 347.400 231.600 351.300 ;
        RECT 235.800 347.400 237.600 351.300 ;
        RECT 249.000 344.400 250.800 351.300 ;
        RECT 256.500 347.400 258.300 351.300 ;
        RECT 272.400 347.400 274.200 351.300 ;
        RECT 278.400 347.400 280.200 351.300 ;
        RECT 288.150 347.400 289.950 351.300 ;
        RECT 297.450 347.400 299.250 351.300 ;
        RECT 304.350 347.400 306.150 351.300 ;
        RECT 313.350 347.400 315.150 351.300 ;
        RECT 329.400 347.400 331.200 351.300 ;
        RECT 347.400 344.400 349.200 351.300 ;
        RECT 353.400 344.400 355.200 351.300 ;
        RECT 359.400 344.400 361.200 351.300 ;
        RECT 365.400 344.400 367.200 351.300 ;
        RECT 371.400 344.400 373.200 351.300 ;
        RECT 388.800 347.400 390.600 351.300 ;
        RECT 394.800 347.400 396.600 351.300 ;
        RECT 410.700 347.400 412.500 351.300 ;
        RECT 418.200 344.400 420.000 351.300 ;
        RECT 436.800 347.400 438.600 351.300 ;
        RECT 455.400 347.400 457.200 351.300 ;
        RECT 475.800 347.400 477.600 351.300 ;
        RECT 481.800 347.400 483.600 351.300 ;
        RECT 494.400 341.400 496.200 351.300 ;
        RECT 521.400 346.200 523.200 351.300 ;
        RECT 545.400 346.200 547.200 351.300 ;
        RECT 574.500 344.400 576.300 351.300 ;
        RECT 593.400 345.300 595.200 351.300 ;
        RECT 602.400 345.300 604.200 351.300 ;
        RECT 628.800 346.200 630.600 351.300 ;
        RECT 655.800 341.400 657.600 351.300 ;
        RECT 669.000 344.400 670.800 351.300 ;
        RECT 676.500 347.400 678.300 351.300 ;
        RECT 703.800 341.400 705.600 351.300 ;
        RECT 716.400 341.400 718.200 351.300 ;
        RECT 743.700 347.400 745.500 351.300 ;
        RECT 751.200 344.400 753.000 351.300 ;
        RECT 767.400 341.400 769.200 351.300 ;
        RECT 792.000 344.400 793.800 351.300 ;
        RECT 799.500 347.400 801.300 351.300 ;
        RECT 823.800 346.200 825.600 351.300 ;
        RECT 842.400 346.200 844.200 351.300 ;
        RECT 863.400 341.400 865.200 351.300 ;
        RECT 13.800 275.700 15.600 282.600 ;
        RECT 19.800 275.700 21.600 282.600 ;
        RECT 25.800 275.700 27.600 282.600 ;
        RECT 31.800 275.700 33.600 282.600 ;
        RECT 37.800 275.700 39.600 282.600 ;
        RECT 55.500 275.700 57.300 282.600 ;
        RECT 64.500 275.700 66.300 282.600 ;
        RECT 82.500 275.700 84.300 282.600 ;
        RECT 91.500 275.700 93.300 282.600 ;
        RECT 98.850 275.700 100.650 279.600 ;
        RECT 107.850 275.700 109.650 279.600 ;
        RECT 114.750 275.700 116.550 279.600 ;
        RECT 124.050 275.700 125.850 279.600 ;
        RECT 135.150 275.700 136.950 279.600 ;
        RECT 144.450 275.700 146.250 279.600 ;
        RECT 151.350 275.700 153.150 279.600 ;
        RECT 160.350 275.700 162.150 279.600 ;
        RECT 171.150 275.700 172.950 279.600 ;
        RECT 180.450 275.700 182.250 279.600 ;
        RECT 187.350 275.700 189.150 279.600 ;
        RECT 196.350 275.700 198.150 279.600 ;
        RECT 220.500 275.700 222.300 282.600 ;
        RECT 241.500 275.700 243.300 282.600 ;
        RECT 248.850 275.700 250.650 279.600 ;
        RECT 257.850 275.700 259.650 279.600 ;
        RECT 264.750 275.700 266.550 279.600 ;
        RECT 274.050 275.700 275.850 279.600 ;
        RECT 293.400 275.700 295.200 280.800 ;
        RECT 322.500 275.700 324.300 282.600 ;
        RECT 337.800 275.700 339.600 279.600 ;
        RECT 343.800 275.700 345.600 279.600 ;
        RECT 350.850 275.700 352.650 279.600 ;
        RECT 359.850 275.700 361.650 279.600 ;
        RECT 366.750 275.700 368.550 279.600 ;
        RECT 376.050 275.700 377.850 279.600 ;
        RECT 395.700 275.700 397.500 279.600 ;
        RECT 403.200 275.700 405.000 282.600 ;
        RECT 419.400 275.700 421.200 279.600 ;
        RECT 437.700 275.700 439.500 282.600 ;
        RECT 460.800 275.700 462.600 279.600 ;
        RECT 466.800 275.700 468.600 279.600 ;
        RECT 480.000 275.700 481.800 282.600 ;
        RECT 487.500 275.700 489.300 279.600 ;
        RECT 498.150 275.700 499.950 279.600 ;
        RECT 507.450 275.700 509.250 279.600 ;
        RECT 514.350 275.700 516.150 279.600 ;
        RECT 523.350 275.700 525.150 279.600 ;
        RECT 546.300 275.700 548.100 282.600 ;
        RECT 568.800 275.700 570.600 279.600 ;
        RECT 581.400 276.600 583.200 279.600 ;
        RECT 581.400 275.700 582.600 276.600 ;
        RECT 587.400 275.700 589.200 279.600 ;
        RECT 605.400 275.700 607.200 279.600 ;
        RECT 627.000 275.700 628.800 282.600 ;
        RECT 634.500 275.700 636.300 279.600 ;
        RECT 655.800 275.700 657.600 279.600 ;
        RECT 668.400 275.700 670.200 279.600 ;
        RECT 686.400 275.700 688.200 285.600 ;
        RECT 716.400 275.700 718.200 280.800 ;
        RECT 740.400 275.700 742.200 280.800 ;
        RECT 761.400 275.700 763.200 285.600 ;
        RECT 785.400 275.700 787.200 285.600 ;
        RECT 812.400 275.700 814.200 279.600 ;
        RECT 831.000 275.700 832.800 282.600 ;
        RECT 838.500 275.700 840.300 279.600 ;
        RECT 865.800 275.700 867.600 285.600 ;
        RECT 879.000 275.700 880.800 282.600 ;
        RECT 886.500 275.700 888.300 279.600 ;
        RECT 897.450 275.700 906.450 351.300 ;
        RECT 0.600 273.300 906.450 275.700 ;
        RECT 13.800 266.400 15.600 273.300 ;
        RECT 19.800 266.400 21.600 273.300 ;
        RECT 25.800 266.400 27.600 273.300 ;
        RECT 31.800 266.400 33.600 273.300 ;
        RECT 37.800 266.400 39.600 273.300 ;
        RECT 58.800 268.200 60.600 273.300 ;
        RECT 82.800 269.400 84.600 273.300 ;
        RECT 103.800 266.400 105.600 273.300 ;
        RECT 121.500 266.400 123.300 273.300 ;
        RECT 130.500 266.400 132.300 273.300 ;
        RECT 151.500 266.400 153.300 273.300 ;
        RECT 158.850 269.400 160.650 273.300 ;
        RECT 167.850 269.400 169.650 273.300 ;
        RECT 174.750 269.400 176.550 273.300 ;
        RECT 184.050 269.400 185.850 273.300 ;
        RECT 208.800 268.200 210.600 273.300 ;
        RECT 224.400 263.400 226.200 273.300 ;
        RECT 250.800 269.400 252.600 273.300 ;
        RECT 256.800 269.400 258.600 273.300 ;
        RECT 263.850 269.400 265.650 273.300 ;
        RECT 272.850 269.400 274.650 273.300 ;
        RECT 279.750 269.400 281.550 273.300 ;
        RECT 289.050 269.400 290.850 273.300 ;
        RECT 305.400 266.400 307.200 273.300 ;
        RECT 311.400 266.400 313.200 273.300 ;
        RECT 317.400 266.400 319.200 273.300 ;
        RECT 332.400 269.400 334.200 273.300 ;
        RECT 353.400 269.400 355.200 273.300 ;
        RECT 366.150 269.400 367.950 273.300 ;
        RECT 375.450 269.400 377.250 273.300 ;
        RECT 382.350 269.400 384.150 273.300 ;
        RECT 391.350 269.400 393.150 273.300 ;
        RECT 407.400 269.400 409.200 273.300 ;
        RECT 428.400 268.200 430.200 273.300 ;
        RECT 452.400 269.400 454.200 273.300 ;
        RECT 465.150 269.400 466.950 273.300 ;
        RECT 474.450 269.400 476.250 273.300 ;
        RECT 481.350 269.400 483.150 273.300 ;
        RECT 490.350 269.400 492.150 273.300 ;
        RECT 509.400 268.200 511.200 273.300 ;
        RECT 530.700 266.400 532.500 273.300 ;
        RECT 559.500 266.400 561.300 273.300 ;
        RECT 577.800 269.400 579.600 273.300 ;
        RECT 584.400 272.400 585.600 273.300 ;
        RECT 583.800 269.400 585.600 272.400 ;
        RECT 604.500 266.400 606.300 273.300 ;
        RECT 620.400 268.200 622.200 273.300 ;
        RECT 650.100 267.300 651.900 273.300 ;
        RECT 658.800 267.300 660.600 273.300 ;
        RECT 682.500 266.400 684.300 273.300 ;
        RECT 698.700 269.400 700.500 273.300 ;
        RECT 706.200 266.400 708.000 273.300 ;
        RECT 719.400 263.400 721.200 273.300 ;
        RECT 754.800 263.400 756.600 273.300 ;
        RECT 775.500 266.400 777.300 273.300 ;
        RECT 788.400 263.400 790.200 273.300 ;
        RECT 820.800 268.200 822.600 273.300 ;
        RECT 836.400 263.400 838.200 273.300 ;
        RECT 863.700 269.400 865.500 273.300 ;
        RECT 871.200 266.400 873.000 273.300 ;
        RECT 6.150 197.700 7.950 201.600 ;
        RECT 15.450 197.700 17.250 201.600 ;
        RECT 22.350 197.700 24.150 201.600 ;
        RECT 31.350 197.700 33.150 201.600 ;
        RECT 55.800 197.700 57.600 202.800 ;
        RECT 71.400 197.700 73.200 201.600 ;
        RECT 97.800 197.700 99.600 202.800 ;
        RECT 113.400 197.700 115.200 201.600 ;
        RECT 119.400 197.700 121.200 201.600 ;
        RECT 136.800 197.700 138.600 201.600 ;
        RECT 142.800 197.700 144.600 201.600 ;
        RECT 163.800 197.700 165.600 202.800 ;
        RECT 179.400 197.700 181.200 201.600 ;
        RECT 185.400 197.700 187.200 201.600 ;
        RECT 211.800 197.700 213.600 202.800 ;
        RECT 221.850 197.700 223.650 201.600 ;
        RECT 230.850 197.700 232.650 201.600 ;
        RECT 237.750 197.700 239.550 201.600 ;
        RECT 247.050 197.700 248.850 201.600 ;
        RECT 263.700 197.700 265.500 204.600 ;
        RECT 292.800 197.700 294.600 202.800 ;
        RECT 316.800 197.700 318.600 202.800 ;
        RECT 334.800 197.700 336.600 201.600 ;
        RECT 340.800 197.700 342.600 201.600 ;
        RECT 358.800 197.700 360.600 201.600 ;
        RECT 378.300 197.700 380.100 204.600 ;
        RECT 400.800 197.700 402.600 201.600 ;
        RECT 406.800 198.600 408.600 201.600 ;
        RECT 407.400 197.700 408.600 198.600 ;
        RECT 419.700 197.700 421.500 204.600 ;
        RECT 435.150 197.700 436.950 201.600 ;
        RECT 444.450 197.700 446.250 201.600 ;
        RECT 451.350 197.700 453.150 201.600 ;
        RECT 460.350 197.700 462.150 201.600 ;
        RECT 476.400 197.700 478.200 201.600 ;
        RECT 497.400 197.700 499.200 202.800 ;
        RECT 518.700 197.700 520.500 204.600 ;
        RECT 533.850 197.700 535.650 201.600 ;
        RECT 542.850 197.700 544.650 201.600 ;
        RECT 549.750 197.700 551.550 201.600 ;
        RECT 559.050 197.700 560.850 201.600 ;
        RECT 578.700 197.700 580.500 204.600 ;
        RECT 607.800 197.700 609.600 202.800 ;
        RECT 627.900 197.700 629.700 204.600 ;
        RECT 651.900 197.700 653.700 204.600 ;
        RECT 674.700 197.700 676.500 201.600 ;
        RECT 682.200 197.700 684.000 204.600 ;
        RECT 698.400 197.700 700.200 203.700 ;
        RECT 707.400 197.700 709.200 203.700 ;
        RECT 730.800 197.700 732.600 203.700 ;
        RECT 739.800 197.700 741.600 203.700 ;
        RECT 758.700 197.700 760.500 201.600 ;
        RECT 766.200 197.700 768.000 204.600 ;
        RECT 784.800 197.700 786.600 201.600 ;
        RECT 797.700 197.700 799.500 204.600 ;
        RECT 825.300 197.700 827.100 204.600 ;
        RECT 842.400 197.700 844.200 207.600 ;
        RECT 874.800 197.700 876.600 202.800 ;
        RECT 897.450 197.700 906.450 273.300 ;
        RECT 0.600 195.300 906.450 197.700 ;
        RECT 19.800 190.200 21.600 195.300 ;
        RECT 35.700 188.400 37.500 195.300 ;
        RECT 64.800 190.200 66.600 195.300 ;
        RECT 83.400 190.200 85.200 195.300 ;
        RECT 98.850 191.400 100.650 195.300 ;
        RECT 107.850 191.400 109.650 195.300 ;
        RECT 114.750 191.400 116.550 195.300 ;
        RECT 124.050 191.400 125.850 195.300 ;
        RECT 140.700 188.400 142.500 195.300 ;
        RECT 169.800 190.200 171.600 195.300 ;
        RECT 185.700 188.400 187.500 195.300 ;
        RECT 214.500 188.400 216.300 195.300 ;
        RECT 221.850 191.400 223.650 195.300 ;
        RECT 230.850 191.400 232.650 195.300 ;
        RECT 237.750 191.400 239.550 195.300 ;
        RECT 247.050 191.400 248.850 195.300 ;
        RECT 271.800 190.200 273.600 195.300 ;
        RECT 290.700 191.400 292.500 195.300 ;
        RECT 298.200 188.400 300.000 195.300 ;
        RECT 313.800 191.400 315.600 195.300 ;
        RECT 319.800 191.400 321.600 195.300 ;
        RECT 337.800 189.300 339.600 195.300 ;
        RECT 346.800 189.300 348.600 195.300 ;
        RECT 365.400 190.200 367.200 195.300 ;
        RECT 391.800 191.400 393.600 195.300 ;
        RECT 412.800 190.200 414.600 195.300 ;
        RECT 431.400 191.400 433.200 195.300 ;
        RECT 437.400 191.400 439.200 195.300 ;
        RECT 452.400 191.400 454.200 195.300 ;
        RECT 475.800 191.400 477.600 195.300 ;
        RECT 482.850 191.400 484.650 195.300 ;
        RECT 491.850 191.400 493.650 195.300 ;
        RECT 498.750 191.400 500.550 195.300 ;
        RECT 508.050 191.400 509.850 195.300 ;
        RECT 524.400 191.400 526.200 195.300 ;
        RECT 530.400 191.400 532.200 195.300 ;
        RECT 545.700 188.400 547.500 195.300 ;
        RECT 561.150 191.400 562.950 195.300 ;
        RECT 570.450 191.400 572.250 195.300 ;
        RECT 577.350 191.400 579.150 195.300 ;
        RECT 586.350 191.400 588.150 195.300 ;
        RECT 610.800 190.200 612.600 195.300 ;
        RECT 626.700 188.400 628.500 195.300 ;
        RECT 655.800 190.200 657.600 195.300 ;
        RECT 674.700 188.400 676.500 195.300 ;
        RECT 683.700 188.400 685.500 195.300 ;
        RECT 701.400 191.400 703.200 195.300 ;
        RECT 707.400 191.400 709.200 195.300 ;
        RECT 722.400 191.400 724.200 195.300 ;
        RECT 743.400 190.200 745.200 195.300 ;
        RECT 764.400 191.400 766.200 195.300 ;
        RECT 783.000 188.400 784.800 195.300 ;
        RECT 790.500 191.400 792.300 195.300 ;
        RECT 808.800 191.400 810.600 195.300 ;
        RECT 814.800 191.400 816.600 195.300 ;
        RECT 827.700 188.400 829.500 195.300 ;
        RECT 848.700 188.400 850.500 195.300 ;
        RECT 869.700 188.400 871.500 195.300 ;
        RECT 16.800 119.700 18.600 123.600 ;
        RECT 32.400 119.700 34.200 126.600 ;
        RECT 38.400 119.700 40.200 126.600 ;
        RECT 44.400 119.700 46.200 126.600 ;
        RECT 50.400 119.700 52.200 126.600 ;
        RECT 56.400 119.700 58.200 126.600 ;
        RECT 79.500 119.700 81.300 126.600 ;
        RECT 96.900 119.700 98.700 126.600 ;
        RECT 127.800 119.700 129.600 124.800 ;
        RECT 146.400 119.700 148.200 124.800 ;
        RECT 172.800 119.700 174.600 123.600 ;
        RECT 193.800 119.700 195.600 123.600 ;
        RECT 200.850 119.700 202.650 123.600 ;
        RECT 209.850 119.700 211.650 123.600 ;
        RECT 216.750 119.700 218.550 123.600 ;
        RECT 226.050 119.700 227.850 123.600 ;
        RECT 245.400 119.700 247.200 124.800 ;
        RECT 274.500 119.700 276.300 126.600 ;
        RECT 295.800 119.700 297.600 124.800 ;
        RECT 305.850 119.700 307.650 123.600 ;
        RECT 314.850 119.700 316.650 123.600 ;
        RECT 321.750 119.700 323.550 123.600 ;
        RECT 331.050 119.700 332.850 123.600 ;
        RECT 352.800 119.700 354.600 123.600 ;
        RECT 368.700 119.700 370.500 126.600 ;
        RECT 389.400 119.700 391.200 126.600 ;
        RECT 395.400 119.700 397.200 126.600 ;
        RECT 401.400 119.700 403.200 126.600 ;
        RECT 407.400 119.700 409.200 126.600 ;
        RECT 413.400 119.700 415.200 126.600 ;
        RECT 436.500 119.700 438.300 126.600 ;
        RECT 457.800 119.700 459.600 124.800 ;
        RECT 467.850 119.700 469.650 123.600 ;
        RECT 476.850 119.700 478.650 123.600 ;
        RECT 483.750 119.700 485.550 123.600 ;
        RECT 493.050 119.700 494.850 123.600 ;
        RECT 509.700 119.700 511.500 126.600 ;
        RECT 518.700 119.700 520.500 126.600 ;
        RECT 541.800 119.700 543.600 123.600 ;
        RECT 547.800 120.600 549.600 123.600 ;
        RECT 548.400 119.700 549.600 120.600 ;
        RECT 564.000 119.700 565.800 126.600 ;
        RECT 571.500 119.700 573.300 123.600 ;
        RECT 587.400 119.700 589.200 123.600 ;
        RECT 610.800 119.700 612.600 123.600 ;
        RECT 617.850 119.700 619.650 123.600 ;
        RECT 626.850 119.700 628.650 123.600 ;
        RECT 633.750 119.700 635.550 123.600 ;
        RECT 643.050 119.700 644.850 123.600 ;
        RECT 664.800 119.700 666.600 123.600 ;
        RECT 671.850 119.700 673.650 123.600 ;
        RECT 680.850 119.700 682.650 123.600 ;
        RECT 687.750 119.700 689.550 123.600 ;
        RECT 697.050 119.700 698.850 123.600 ;
        RECT 716.400 119.700 718.200 125.100 ;
        RECT 743.400 119.700 745.200 124.800 ;
        RECT 767.700 119.700 769.500 123.600 ;
        RECT 775.200 119.700 777.000 126.600 ;
        RECT 791.400 119.700 793.200 124.800 ;
        RECT 817.800 119.700 819.600 123.600 ;
        RECT 838.800 119.700 840.600 124.800 ;
        RECT 859.800 119.700 861.600 123.600 ;
        RECT 872.400 119.700 874.200 129.600 ;
        RECT 897.450 119.700 906.450 195.300 ;
        RECT 0.600 117.300 906.450 119.700 ;
        RECT 16.800 111.300 18.600 117.300 ;
        RECT 25.800 111.300 27.600 117.300 ;
        RECT 43.800 113.400 45.600 117.300 ;
        RECT 49.800 113.400 51.600 117.300 ;
        RECT 70.500 110.400 72.300 117.300 ;
        RECT 85.800 113.400 87.600 117.300 ;
        RECT 91.800 113.400 93.600 117.300 ;
        RECT 104.400 113.400 106.200 117.300 ;
        RECT 124.800 113.400 126.600 117.300 ;
        RECT 130.800 113.400 132.600 117.300 ;
        RECT 146.400 113.400 148.200 117.300 ;
        RECT 166.800 113.400 168.600 117.300 ;
        RECT 172.800 113.400 174.600 117.300 ;
        RECT 187.800 113.400 189.600 117.300 ;
        RECT 193.800 113.400 195.600 117.300 ;
        RECT 214.800 113.400 216.600 117.300 ;
        RECT 221.850 113.400 223.650 117.300 ;
        RECT 230.850 113.400 232.650 117.300 ;
        RECT 237.750 113.400 239.550 117.300 ;
        RECT 247.050 113.400 248.850 117.300 ;
        RECT 266.400 112.200 268.200 117.300 ;
        RECT 292.800 113.400 294.600 117.300 ;
        RECT 299.850 113.400 301.650 117.300 ;
        RECT 308.850 113.400 310.650 117.300 ;
        RECT 315.750 113.400 317.550 117.300 ;
        RECT 325.050 113.400 326.850 117.300 ;
        RECT 344.400 111.900 346.200 117.300 ;
        RECT 370.800 113.400 372.600 117.300 ;
        RECT 376.800 113.400 378.600 117.300 ;
        RECT 383.850 113.400 385.650 117.300 ;
        RECT 392.850 113.400 394.650 117.300 ;
        RECT 399.750 113.400 401.550 117.300 ;
        RECT 409.050 113.400 410.850 117.300 ;
        RECT 428.700 113.400 430.500 117.300 ;
        RECT 436.200 110.400 438.000 117.300 ;
        RECT 451.800 113.400 453.600 117.300 ;
        RECT 457.800 113.400 459.600 117.300 ;
        RECT 478.800 112.200 480.600 117.300 ;
        RECT 494.400 113.400 496.200 117.300 ;
        RECT 514.800 113.400 516.600 117.300 ;
        RECT 520.800 113.400 522.600 117.300 ;
        RECT 536.400 112.200 538.200 117.300 ;
        RECT 562.800 113.400 564.600 117.300 ;
        RECT 579.900 110.400 581.700 117.300 ;
        RECT 607.500 110.400 609.300 117.300 ;
        RECT 623.400 113.400 625.200 117.300 ;
        RECT 629.400 113.400 631.200 117.300 ;
        RECT 649.800 113.400 651.600 117.300 ;
        RECT 656.850 113.400 658.650 117.300 ;
        RECT 665.850 113.400 667.650 117.300 ;
        RECT 672.750 113.400 674.550 117.300 ;
        RECT 682.050 113.400 683.850 117.300 ;
        RECT 709.800 107.400 711.600 117.300 ;
        RECT 722.700 110.400 724.500 117.300 ;
        RECT 746.400 111.300 748.200 117.300 ;
        RECT 755.400 111.300 757.200 117.300 ;
        RECT 774.000 110.400 775.800 117.300 ;
        RECT 781.500 113.400 783.300 117.300 ;
        RECT 798.000 110.400 799.800 117.300 ;
        RECT 805.500 113.400 807.300 117.300 ;
        RECT 823.800 113.400 825.600 117.300 ;
        RECT 829.800 113.400 831.600 117.300 ;
        RECT 842.400 113.400 844.200 117.300 ;
        RECT 848.400 113.400 850.200 117.300 ;
        RECT 863.400 113.400 865.200 117.300 ;
        RECT 869.400 113.400 871.200 117.300 ;
        RECT 884.400 113.400 886.200 117.300 ;
        RECT 13.800 41.700 15.600 45.600 ;
        RECT 19.800 41.700 21.600 45.600 ;
        RECT 32.400 41.700 34.200 45.600 ;
        RECT 38.400 41.700 40.200 45.600 ;
        RECT 54.000 41.700 55.800 48.600 ;
        RECT 61.500 41.700 63.300 45.600 ;
        RECT 85.800 41.700 87.600 46.800 ;
        RECT 101.700 41.700 103.500 48.600 ;
        RECT 122.700 41.700 124.500 48.600 ;
        RECT 137.850 41.700 139.650 45.600 ;
        RECT 146.850 41.700 148.650 45.600 ;
        RECT 153.750 41.700 155.550 45.600 ;
        RECT 163.050 41.700 164.850 45.600 ;
        RECT 179.400 41.700 181.200 45.600 ;
        RECT 185.400 41.700 187.200 45.600 ;
        RECT 203.700 41.700 205.500 45.600 ;
        RECT 211.200 41.700 213.000 48.600 ;
        RECT 227.400 41.700 229.200 46.800 ;
        RECT 242.850 41.700 244.650 45.600 ;
        RECT 251.850 41.700 253.650 45.600 ;
        RECT 258.750 41.700 260.550 45.600 ;
        RECT 268.050 41.700 269.850 45.600 ;
        RECT 284.400 41.700 286.200 45.600 ;
        RECT 310.500 41.700 312.300 48.600 ;
        RECT 334.800 41.700 336.600 51.600 ;
        RECT 347.400 41.700 349.200 45.600 ;
        RECT 353.400 41.700 355.200 45.600 ;
        RECT 376.800 41.700 378.600 46.800 ;
        RECT 397.800 41.700 399.600 45.600 ;
        RECT 413.400 41.700 415.200 46.800 ;
        RECT 434.400 41.700 436.200 45.600 ;
        RECT 455.400 41.700 457.200 46.800 ;
        RECT 481.800 41.700 483.600 45.600 ;
        RECT 497.700 41.700 499.500 45.600 ;
        RECT 505.200 41.700 507.000 48.600 ;
        RECT 526.800 41.700 528.600 45.600 ;
        RECT 544.800 41.700 546.600 45.600 ;
        RECT 560.700 41.700 562.500 45.600 ;
        RECT 568.200 41.700 570.000 48.600 ;
        RECT 583.800 41.700 585.600 45.600 ;
        RECT 589.800 41.700 591.600 45.600 ;
        RECT 604.800 41.700 606.600 45.600 ;
        RECT 610.800 41.700 612.600 45.600 ;
        RECT 628.800 41.700 630.600 45.600 ;
        RECT 641.400 41.700 643.200 45.600 ;
        RECT 647.400 41.700 649.200 45.600 ;
        RECT 673.800 41.700 675.600 51.600 ;
        RECT 697.800 41.700 699.600 51.600 ;
        RECT 710.400 41.700 712.200 45.600 ;
        RECT 728.400 41.700 730.200 51.600 ;
        RECT 760.500 41.700 762.300 48.600 ;
        RECT 773.400 41.700 775.200 51.600 ;
        RECT 797.400 41.700 799.200 45.600 ;
        RECT 815.400 41.700 817.200 45.600 ;
        RECT 836.400 41.700 838.200 45.600 ;
        RECT 854.400 41.700 856.200 51.600 ;
        RECT 878.400 41.700 880.200 45.600 ;
        RECT 897.450 41.700 906.450 117.300 ;
        RECT 0.600 39.300 906.450 41.700 ;
        RECT 16.800 35.400 18.600 39.300 ;
        RECT 29.700 32.400 31.500 39.300 ;
        RECT 55.800 35.400 57.600 39.300 ;
        RECT 76.800 35.400 78.600 39.300 ;
        RECT 86.850 35.400 88.650 39.300 ;
        RECT 95.850 35.400 97.650 39.300 ;
        RECT 102.750 35.400 104.550 39.300 ;
        RECT 112.050 35.400 113.850 39.300 ;
        RECT 131.400 35.400 133.200 39.300 ;
        RECT 152.400 34.200 154.200 39.300 ;
        RECT 173.700 32.400 175.500 39.300 ;
        RECT 188.850 35.400 190.650 39.300 ;
        RECT 197.850 35.400 199.650 39.300 ;
        RECT 204.750 35.400 206.550 39.300 ;
        RECT 214.050 35.400 215.850 39.300 ;
        RECT 238.500 32.400 240.300 39.300 ;
        RECT 259.500 32.400 261.300 39.300 ;
        RECT 280.800 34.200 282.600 39.300 ;
        RECT 291.150 35.400 292.950 39.300 ;
        RECT 300.450 35.400 302.250 39.300 ;
        RECT 307.350 35.400 309.150 39.300 ;
        RECT 316.350 35.400 318.150 39.300 ;
        RECT 332.400 35.400 334.200 39.300 ;
        RECT 355.800 35.400 357.600 39.300 ;
        RECT 362.850 35.400 364.650 39.300 ;
        RECT 371.850 35.400 373.650 39.300 ;
        RECT 378.750 35.400 380.550 39.300 ;
        RECT 388.050 35.400 389.850 39.300 ;
        RECT 407.400 34.200 409.200 39.300 ;
        RECT 428.700 32.400 430.500 39.300 ;
        RECT 449.700 32.400 451.500 39.300 ;
        RECT 464.850 35.400 466.650 39.300 ;
        RECT 473.850 35.400 475.650 39.300 ;
        RECT 480.750 35.400 482.550 39.300 ;
        RECT 490.050 35.400 491.850 39.300 ;
        RECT 506.400 35.400 508.200 39.300 ;
        RECT 527.400 34.200 529.200 39.300 ;
        RECT 556.500 32.400 558.300 39.300 ;
        RECT 564.150 35.400 565.950 39.300 ;
        RECT 573.450 35.400 575.250 39.300 ;
        RECT 580.350 35.400 582.150 39.300 ;
        RECT 589.350 35.400 591.150 39.300 ;
        RECT 613.500 32.400 615.300 39.300 ;
        RECT 629.400 34.200 631.200 39.300 ;
        RECT 644.850 35.400 646.650 39.300 ;
        RECT 653.850 35.400 655.650 39.300 ;
        RECT 660.750 35.400 662.550 39.300 ;
        RECT 670.050 35.400 671.850 39.300 ;
        RECT 694.500 32.400 696.300 39.300 ;
        RECT 715.800 34.200 717.600 39.300 ;
        RECT 731.700 32.400 733.500 39.300 ;
        RECT 757.800 35.400 759.600 39.300 ;
        RECT 764.400 38.400 765.600 39.300 ;
        RECT 763.800 35.400 765.600 38.400 ;
        RECT 783.300 32.400 785.100 39.300 ;
        RECT 803.400 34.200 805.200 39.300 ;
        RECT 824.400 35.400 826.200 39.300 ;
        RECT 843.000 32.400 844.800 39.300 ;
        RECT 850.500 35.400 852.300 39.300 ;
        RECT 874.800 34.200 876.600 39.300 ;
        RECT 897.450 0.300 906.450 39.300 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -9.450 860.700 -0.450 899.700 ;
        RECT 16.800 860.700 18.600 867.600 ;
        RECT 29.400 860.700 31.200 867.600 ;
        RECT 35.400 860.700 37.200 867.600 ;
        RECT 44.550 860.700 46.350 864.600 ;
        RECT 53.250 860.700 55.050 867.600 ;
        RECT 59.850 860.700 61.650 867.600 ;
        RECT 70.050 860.700 71.850 867.600 ;
        RECT 80.550 860.700 82.350 864.600 ;
        RECT 89.250 860.700 91.050 867.600 ;
        RECT 95.850 860.700 97.650 867.600 ;
        RECT 106.050 860.700 107.850 867.600 ;
        RECT 122.400 860.700 124.200 873.600 ;
        RECT 128.400 860.700 130.200 873.600 ;
        RECT 134.400 860.700 136.200 873.600 ;
        RECT 140.400 860.700 142.200 873.600 ;
        RECT 146.400 860.700 148.200 873.600 ;
        RECT 164.400 860.700 166.200 871.500 ;
        RECT 173.100 860.700 175.200 871.500 ;
        RECT 193.800 860.700 195.600 867.600 ;
        RECT 199.800 860.700 201.600 867.600 ;
        RECT 214.800 860.700 216.600 867.600 ;
        RECT 220.800 860.700 222.600 867.600 ;
        RECT 244.800 860.700 246.600 871.500 ;
        RECT 265.800 860.700 267.600 867.000 ;
        RECT 271.800 860.700 273.600 867.600 ;
        RECT 289.800 860.700 291.600 867.600 ;
        RECT 307.800 860.700 309.600 867.000 ;
        RECT 313.800 860.700 315.600 867.600 ;
        RECT 331.800 860.700 333.600 867.600 ;
        RECT 347.400 860.700 349.200 873.600 ;
        RECT 368.700 860.700 370.500 873.600 ;
        RECT 376.800 860.700 378.600 867.600 ;
        RECT 397.800 860.700 399.600 867.000 ;
        RECT 403.800 860.700 405.600 867.600 ;
        RECT 416.400 860.700 418.200 867.600 ;
        RECT 442.800 860.700 444.600 867.000 ;
        RECT 448.800 860.700 450.600 867.600 ;
        RECT 464.400 860.700 466.200 871.800 ;
        RECT 485.700 860.700 487.500 873.600 ;
        RECT 493.800 860.700 495.600 867.600 ;
        RECT 509.400 860.700 511.200 867.600 ;
        RECT 530.400 860.700 532.200 871.800 ;
        RECT 556.800 860.700 558.900 871.500 ;
        RECT 565.800 860.700 567.600 871.500 ;
        RECT 581.700 860.700 583.500 873.600 ;
        RECT 589.800 860.700 591.600 867.600 ;
        RECT 610.800 860.700 612.600 867.000 ;
        RECT 616.800 860.700 618.600 867.600 ;
        RECT 632.400 860.700 634.200 867.600 ;
        RECT 640.500 860.700 642.300 873.600 ;
        RECT 658.800 860.700 660.600 867.000 ;
        RECT 664.800 860.700 666.600 867.600 ;
        RECT 677.400 860.700 679.200 867.600 ;
        RECT 683.400 860.700 685.200 867.600 ;
        RECT 706.800 860.700 708.600 871.800 ;
        RECT 727.800 860.700 729.600 867.000 ;
        RECT 733.800 860.700 735.600 867.600 ;
        RECT 751.800 860.700 753.600 867.000 ;
        RECT 757.800 860.700 759.600 867.600 ;
        RECT 773.400 860.700 775.200 871.800 ;
        RECT 799.800 860.700 801.600 867.600 ;
        RECT 812.400 860.700 814.200 867.600 ;
        RECT 833.400 860.700 835.200 871.800 ;
        RECT 854.700 860.700 856.500 873.600 ;
        RECT 862.800 860.700 864.600 867.600 ;
        RECT 878.400 860.700 880.200 867.600 ;
        RECT 884.400 860.700 886.200 867.000 ;
        RECT -9.450 858.300 896.400 860.700 ;
        RECT -9.450 782.700 -0.450 858.300 ;
        RECT 11.400 851.400 13.200 858.300 ;
        RECT 17.400 851.400 19.200 858.300 ;
        RECT 35.400 851.400 37.200 858.300 ;
        RECT 47.550 854.400 49.350 858.300 ;
        RECT 56.250 851.400 58.050 858.300 ;
        RECT 62.850 851.400 64.650 858.300 ;
        RECT 73.050 851.400 74.850 858.300 ;
        RECT 89.400 845.400 91.200 858.300 ;
        RECT 99.900 845.400 101.700 858.300 ;
        RECT 116.400 845.400 118.200 858.300 ;
        RECT 126.900 845.400 128.700 858.300 ;
        RECT 143.400 851.400 145.200 858.300 ;
        RECT 149.400 851.400 151.200 858.300 ;
        RECT 167.400 851.400 169.200 858.300 ;
        RECT 173.400 851.400 175.200 858.300 ;
        RECT 196.800 847.200 198.600 858.300 ;
        RECT 212.400 851.400 214.200 858.300 ;
        RECT 218.400 852.000 220.200 858.300 ;
        RECT 239.400 847.200 241.200 858.300 ;
        RECT 263.400 851.400 265.200 858.300 ;
        RECT 271.500 845.400 273.300 858.300 ;
        RECT 292.800 847.200 294.600 858.300 ;
        RECT 311.400 847.200 313.200 858.300 ;
        RECT 335.400 851.400 337.200 858.300 ;
        RECT 343.500 845.400 345.300 858.300 ;
        RECT 364.800 847.200 366.600 858.300 ;
        RECT 380.400 851.400 382.200 858.300 ;
        RECT 386.400 852.000 388.200 858.300 ;
        RECT 404.700 845.400 406.500 858.300 ;
        RECT 412.800 851.400 414.600 858.300 ;
        RECT 433.800 852.000 435.600 858.300 ;
        RECT 439.800 851.400 441.600 858.300 ;
        RECT 457.800 852.000 459.600 858.300 ;
        RECT 463.800 851.400 465.600 858.300 ;
        RECT 479.400 851.400 481.200 858.300 ;
        RECT 487.500 845.400 489.300 858.300 ;
        RECT 500.700 845.400 502.500 858.300 ;
        RECT 508.800 851.400 510.600 858.300 ;
        RECT 532.800 847.200 534.600 858.300 ;
        RECT 553.800 852.000 555.600 858.300 ;
        RECT 559.800 851.400 561.600 858.300 ;
        RECT 577.800 847.500 579.600 858.300 ;
        RECT 586.800 847.500 588.600 858.300 ;
        RECT 602.400 851.400 604.200 858.300 ;
        RECT 608.400 852.000 610.200 858.300 ;
        RECT 626.700 845.400 628.500 858.300 ;
        RECT 634.800 851.400 636.600 858.300 ;
        RECT 652.800 851.400 654.600 858.300 ;
        RECT 658.800 851.400 660.600 858.300 ;
        RECT 673.800 851.400 675.600 858.300 ;
        RECT 679.800 851.400 681.600 858.300 ;
        RECT 692.400 851.400 694.200 858.300 ;
        RECT 698.400 851.400 700.200 858.300 ;
        RECT 718.800 851.400 720.600 858.300 ;
        RECT 724.800 851.400 726.600 858.300 ;
        RECT 742.800 852.000 744.600 858.300 ;
        RECT 748.800 851.400 750.600 858.300 ;
        RECT 764.400 847.200 766.200 858.300 ;
        RECT 785.700 845.400 787.500 858.300 ;
        RECT 793.800 851.400 795.600 858.300 ;
        RECT 809.400 851.400 811.200 858.300 ;
        RECT 815.400 852.000 817.200 858.300 ;
        RECT 836.400 851.400 838.200 858.300 ;
        RECT 844.500 845.400 846.300 858.300 ;
        RECT 868.800 847.200 870.600 858.300 ;
        RECT 11.400 782.700 13.200 789.600 ;
        RECT 17.400 782.700 19.200 789.600 ;
        RECT 32.400 782.700 34.200 789.600 ;
        RECT 53.400 782.700 55.200 789.600 ;
        RECT 61.500 782.700 63.300 795.600 ;
        RECT 69.150 782.700 70.950 789.600 ;
        RECT 79.350 782.700 81.150 789.600 ;
        RECT 85.950 782.700 87.750 789.600 ;
        RECT 94.650 782.700 96.450 786.600 ;
        RECT 110.400 782.700 112.200 789.600 ;
        RECT 128.700 782.700 130.500 795.600 ;
        RECT 136.800 782.700 138.600 789.600 ;
        RECT 157.800 782.700 159.600 789.600 ;
        RECT 172.800 782.700 174.600 789.600 ;
        RECT 178.800 782.700 180.600 789.600 ;
        RECT 196.800 782.700 198.600 789.600 ;
        RECT 217.800 782.700 219.600 789.000 ;
        RECT 223.800 782.700 225.600 789.600 ;
        RECT 241.800 782.700 243.600 789.600 ;
        RECT 254.700 782.700 256.500 795.600 ;
        RECT 262.800 782.700 264.600 789.600 ;
        RECT 283.800 782.700 285.600 789.000 ;
        RECT 289.800 782.700 291.600 789.600 ;
        RECT 305.400 782.700 307.200 793.800 ;
        RECT 331.800 782.700 333.600 789.000 ;
        RECT 337.800 782.700 339.600 789.600 ;
        RECT 355.800 782.700 357.600 789.600 ;
        RECT 373.800 782.700 375.600 789.000 ;
        RECT 379.800 782.700 381.600 789.600 ;
        RECT 395.400 782.700 397.200 789.600 ;
        RECT 403.500 782.700 405.300 795.600 ;
        RECT 418.800 782.700 420.600 789.600 ;
        RECT 424.800 782.700 426.600 789.600 ;
        RECT 442.800 782.700 444.600 789.000 ;
        RECT 448.800 782.700 450.600 789.600 ;
        RECT 469.800 782.700 471.600 793.800 ;
        RECT 490.800 782.700 492.600 789.600 ;
        RECT 496.800 782.700 498.600 789.600 ;
        RECT 511.800 782.700 513.600 789.600 ;
        RECT 517.800 782.700 519.600 789.600 ;
        RECT 538.800 782.700 540.600 789.600 ;
        RECT 554.400 782.700 556.200 793.800 ;
        RECT 578.400 782.700 580.200 789.600 ;
        RECT 586.500 782.700 588.300 795.600 ;
        RECT 599.700 782.700 601.500 795.600 ;
        RECT 607.800 782.700 609.600 789.600 ;
        RECT 631.800 782.700 633.600 789.000 ;
        RECT 637.800 782.700 639.600 789.600 ;
        RECT 655.800 782.700 657.600 789.000 ;
        RECT 661.800 782.700 663.600 789.600 ;
        RECT 677.400 782.700 679.200 793.800 ;
        RECT 698.700 782.700 700.500 795.600 ;
        RECT 706.800 782.700 708.600 789.600 ;
        RECT 725.400 782.700 727.200 789.600 ;
        RECT 733.500 782.700 735.300 795.600 ;
        RECT 746.400 782.700 748.200 789.600 ;
        RECT 752.400 782.700 754.200 789.000 ;
        RECT 773.400 782.700 775.200 789.600 ;
        RECT 781.500 782.700 783.300 795.600 ;
        RECT 799.800 782.700 801.600 789.000 ;
        RECT 805.800 782.700 807.600 789.600 ;
        RECT 821.400 782.700 823.200 793.800 ;
        RECT 850.800 782.700 852.600 793.800 ;
        RECT 871.800 782.700 873.600 789.000 ;
        RECT 877.800 782.700 879.600 789.600 ;
        RECT -9.450 780.300 896.400 782.700 ;
        RECT -9.450 704.700 -0.450 780.300 ;
        RECT 16.800 773.400 18.600 780.300 ;
        RECT 29.400 773.400 31.200 780.300 ;
        RECT 35.400 773.400 37.200 780.300 ;
        RECT 50.700 767.400 52.500 780.300 ;
        RECT 58.800 773.400 60.600 780.300 ;
        RECT 74.400 773.400 76.200 780.300 ;
        RECT 80.400 773.400 82.200 780.300 ;
        RECT 95.400 767.400 97.200 780.300 ;
        RECT 116.400 767.400 118.200 780.300 ;
        RECT 137.400 767.400 139.200 780.300 ;
        RECT 158.400 773.400 160.200 780.300 ;
        RECT 176.400 767.400 178.200 780.300 ;
        RECT 186.900 767.400 188.700 780.300 ;
        RECT 208.800 774.000 210.600 780.300 ;
        RECT 214.800 773.400 216.600 780.300 ;
        RECT 232.800 774.000 234.600 780.300 ;
        RECT 238.800 773.400 240.600 780.300 ;
        RECT 259.800 774.000 261.600 780.300 ;
        RECT 265.800 773.400 267.600 780.300 ;
        RECT 286.800 769.200 288.600 780.300 ;
        RECT 302.400 773.400 304.200 780.300 ;
        RECT 308.400 774.000 310.200 780.300 ;
        RECT 326.400 773.400 328.200 780.300 ;
        RECT 332.400 773.400 334.200 780.300 ;
        RECT 352.800 773.400 354.600 780.300 ;
        RECT 368.400 773.400 370.200 780.300 ;
        RECT 376.500 767.400 378.300 780.300 ;
        RECT 397.800 773.400 399.600 780.300 ;
        RECT 410.400 773.400 412.200 780.300 ;
        RECT 416.400 773.400 418.200 780.300 ;
        RECT 435.300 767.400 437.100 780.300 ;
        RECT 445.800 767.400 447.600 780.300 ;
        RECT 458.400 767.400 460.200 780.300 ;
        RECT 479.700 767.400 481.500 780.300 ;
        RECT 487.800 773.400 489.600 780.300 ;
        RECT 506.400 773.400 508.200 780.300 ;
        RECT 512.400 774.000 514.200 780.300 ;
        RECT 535.800 773.400 537.600 780.300 ;
        RECT 548.400 773.400 550.200 780.300 ;
        RECT 554.400 774.000 556.200 780.300 ;
        RECT 575.400 773.400 577.200 780.300 ;
        RECT 583.500 767.400 585.300 780.300 ;
        RECT 596.400 773.400 598.200 780.300 ;
        RECT 602.400 773.400 604.200 780.300 ;
        RECT 617.400 773.400 619.200 780.300 ;
        RECT 623.400 774.000 625.200 780.300 ;
        RECT 646.800 773.400 648.600 780.300 ;
        RECT 664.800 773.400 666.600 780.300 ;
        RECT 677.400 773.400 679.200 780.300 ;
        RECT 683.400 774.000 685.200 780.300 ;
        RECT 706.800 774.000 708.600 780.300 ;
        RECT 712.800 773.400 714.600 780.300 ;
        RECT 728.400 769.200 730.200 780.300 ;
        RECT 749.400 773.400 751.200 780.300 ;
        RECT 755.400 773.400 757.200 780.300 ;
        RECT 772.800 773.400 774.600 780.300 ;
        RECT 778.800 773.400 780.600 780.300 ;
        RECT 791.400 773.400 793.200 780.300 ;
        RECT 797.400 773.400 799.200 780.300 ;
        RECT 818.400 769.200 820.200 780.300 ;
        RECT 847.800 773.400 849.600 780.300 ;
        RECT 860.400 773.400 862.200 780.300 ;
        RECT 866.400 774.000 868.200 780.300 ;
        RECT 11.400 704.700 13.200 711.600 ;
        RECT 17.400 704.700 19.200 711.600 ;
        RECT 32.400 704.700 34.200 711.600 ;
        RECT 55.800 704.700 57.600 711.600 ;
        RECT 71.400 704.700 73.200 711.600 ;
        RECT 79.500 704.700 81.300 717.600 ;
        RECT 97.800 704.700 99.600 711.600 ;
        RECT 104.550 704.700 106.350 708.600 ;
        RECT 113.250 704.700 115.050 711.600 ;
        RECT 119.850 704.700 121.650 711.600 ;
        RECT 130.050 704.700 131.850 711.600 ;
        RECT 149.400 704.700 151.200 711.600 ;
        RECT 157.500 704.700 159.300 717.600 ;
        RECT 164.550 704.700 166.350 708.600 ;
        RECT 173.250 704.700 175.050 711.600 ;
        RECT 179.850 704.700 181.650 711.600 ;
        RECT 190.050 704.700 191.850 711.600 ;
        RECT 214.800 704.700 216.600 715.800 ;
        RECT 233.400 704.700 235.200 711.600 ;
        RECT 241.500 704.700 243.300 717.600 ;
        RECT 254.700 704.700 256.500 717.600 ;
        RECT 262.800 704.700 264.600 711.600 ;
        RECT 286.800 704.700 288.600 715.800 ;
        RECT 307.800 704.700 309.600 711.000 ;
        RECT 313.800 704.700 315.600 711.600 ;
        RECT 326.400 704.700 328.200 711.600 ;
        RECT 347.400 704.700 349.200 715.800 ;
        RECT 368.700 704.700 370.500 717.600 ;
        RECT 376.800 704.700 378.600 711.600 ;
        RECT 392.400 704.700 394.200 717.600 ;
        RECT 413.400 704.700 415.200 711.600 ;
        RECT 419.400 704.700 421.200 711.600 ;
        RECT 439.800 704.700 441.600 711.600 ;
        RECT 458.400 704.700 460.200 711.600 ;
        RECT 466.500 704.700 468.300 717.600 ;
        RECT 484.800 704.700 486.600 711.600 ;
        RECT 499.800 704.700 501.600 711.600 ;
        RECT 505.800 704.700 507.600 711.600 ;
        RECT 518.400 704.700 520.200 711.600 ;
        RECT 524.400 704.700 526.200 711.600 ;
        RECT 539.400 704.700 541.200 711.600 ;
        RECT 545.400 704.700 547.200 711.600 ;
        RECT 560.400 704.700 562.200 711.600 ;
        RECT 566.400 704.700 568.200 711.600 ;
        RECT 586.800 704.700 588.600 711.600 ;
        RECT 592.800 704.700 594.600 711.600 ;
        RECT 605.700 704.700 607.500 717.600 ;
        RECT 613.800 704.700 615.600 711.600 ;
        RECT 634.800 704.700 636.600 711.600 ;
        RECT 640.800 704.700 642.600 711.600 ;
        RECT 653.400 704.700 655.200 711.600 ;
        RECT 659.400 704.700 661.200 711.600 ;
        RECT 682.800 704.700 684.600 715.800 ;
        RECT 698.400 704.700 700.200 711.600 ;
        RECT 704.400 704.700 706.200 711.000 ;
        RECT 725.400 704.700 727.200 711.600 ;
        RECT 733.500 704.700 735.300 717.600 ;
        RECT 746.400 704.700 748.200 711.600 ;
        RECT 752.400 704.700 754.200 711.600 ;
        RECT 767.400 704.700 769.200 711.600 ;
        RECT 790.800 704.700 792.600 711.000 ;
        RECT 796.800 704.700 798.600 711.600 ;
        RECT 812.400 704.700 814.200 715.800 ;
        RECT 836.400 704.700 838.200 711.600 ;
        RECT 842.400 704.700 844.200 711.000 ;
        RECT 860.700 704.700 862.500 717.600 ;
        RECT 868.800 704.700 870.600 711.600 ;
        RECT -9.450 702.300 896.400 704.700 ;
        RECT -9.450 626.700 -0.450 702.300 ;
        RECT 14.400 695.400 16.200 702.300 ;
        RECT 22.500 689.400 24.300 702.300 ;
        RECT 35.700 689.400 37.500 702.300 ;
        RECT 43.800 695.400 45.600 702.300 ;
        RECT 64.800 695.400 66.600 702.300 ;
        RECT 70.800 695.400 72.600 702.300 ;
        RECT 93.300 689.400 95.100 702.300 ;
        RECT 110.400 695.400 112.200 702.300 ;
        RECT 116.400 695.400 118.200 702.300 ;
        RECT 131.400 695.400 133.200 702.300 ;
        RECT 137.400 695.400 139.200 702.300 ;
        RECT 157.800 695.400 159.600 702.300 ;
        RECT 178.800 695.400 180.600 702.300 ;
        RECT 196.800 696.000 198.600 702.300 ;
        RECT 202.800 695.400 204.600 702.300 ;
        RECT 218.400 691.200 220.200 702.300 ;
        RECT 242.400 695.400 244.200 702.300 ;
        RECT 250.500 689.400 252.300 702.300 ;
        RECT 271.800 691.200 273.600 702.300 ;
        RECT 289.800 695.400 291.600 702.300 ;
        RECT 295.800 695.400 297.600 702.300 ;
        RECT 310.800 695.400 312.600 702.300 ;
        RECT 316.800 695.400 318.600 702.300 ;
        RECT 334.800 695.400 336.600 702.300 ;
        RECT 340.800 695.400 342.600 702.300 ;
        RECT 364.800 691.500 366.600 702.300 ;
        RECT 382.800 695.400 384.600 702.300 ;
        RECT 388.800 695.400 390.600 702.300 ;
        RECT 404.400 695.400 406.200 702.300 ;
        RECT 412.500 689.400 414.300 702.300 ;
        RECT 436.800 691.500 438.600 702.300 ;
        RECT 455.700 689.400 457.500 702.300 ;
        RECT 463.800 695.400 465.600 702.300 ;
        RECT 479.700 689.400 481.500 702.300 ;
        RECT 487.800 695.400 489.600 702.300 ;
        RECT 508.800 695.400 510.600 702.300 ;
        RECT 514.800 695.400 516.600 702.300 ;
        RECT 527.700 689.400 529.500 702.300 ;
        RECT 535.800 695.400 537.600 702.300 ;
        RECT 551.400 695.400 553.200 702.300 ;
        RECT 557.400 695.400 559.200 702.300 ;
        RECT 572.700 689.400 574.500 702.300 ;
        RECT 580.800 695.400 582.600 702.300 ;
        RECT 596.700 689.400 598.500 702.300 ;
        RECT 604.800 695.400 606.600 702.300 ;
        RECT 625.800 695.400 627.600 702.300 ;
        RECT 631.800 695.400 633.600 702.300 ;
        RECT 644.400 689.400 646.200 702.300 ;
        RECT 676.800 691.200 678.600 702.300 ;
        RECT 697.800 696.000 699.600 702.300 ;
        RECT 703.800 695.400 705.600 702.300 ;
        RECT 719.400 695.400 721.200 702.300 ;
        RECT 727.500 689.400 729.300 702.300 ;
        RECT 740.700 689.400 742.500 702.300 ;
        RECT 748.800 695.400 750.600 702.300 ;
        RECT 769.800 696.000 771.600 702.300 ;
        RECT 775.800 695.400 777.600 702.300 ;
        RECT 791.400 691.200 793.200 702.300 ;
        RECT 812.700 689.400 814.500 702.300 ;
        RECT 820.800 695.400 822.600 702.300 ;
        RECT 844.800 691.200 846.600 702.300 ;
        RECT 860.400 695.400 862.200 702.300 ;
        RECT 866.400 696.000 868.200 702.300 ;
        RECT 887.400 695.400 889.200 702.300 ;
        RECT 19.800 626.700 21.600 639.600 ;
        RECT 32.400 626.700 34.200 633.600 ;
        RECT 50.700 626.700 52.500 639.600 ;
        RECT 58.800 626.700 60.600 633.600 ;
        RECT 82.800 626.700 84.600 639.600 ;
        RECT 98.400 626.700 100.200 633.600 ;
        RECT 104.400 626.700 106.200 633.000 ;
        RECT 127.800 626.700 129.600 633.600 ;
        RECT 134.550 626.700 136.350 630.600 ;
        RECT 143.250 626.700 145.050 633.600 ;
        RECT 149.850 626.700 151.650 633.600 ;
        RECT 160.050 626.700 161.850 633.600 ;
        RECT 176.700 626.700 178.500 639.600 ;
        RECT 184.800 626.700 186.600 633.600 ;
        RECT 205.800 626.700 207.600 633.600 ;
        RECT 221.400 626.700 223.200 633.600 ;
        RECT 229.500 626.700 231.300 639.600 ;
        RECT 250.800 626.700 252.600 637.800 ;
        RECT 266.400 626.700 268.200 633.600 ;
        RECT 272.400 626.700 274.200 633.000 ;
        RECT 296.400 626.700 298.200 633.600 ;
        RECT 304.500 626.700 306.300 639.600 ;
        RECT 317.400 626.700 319.200 639.600 ;
        RECT 338.400 626.700 340.200 633.600 ;
        RECT 344.400 626.700 346.200 633.600 ;
        RECT 364.800 626.700 366.600 633.600 ;
        RECT 370.800 626.700 372.600 633.600 ;
        RECT 386.400 626.700 388.200 633.600 ;
        RECT 394.500 626.700 396.300 639.600 ;
        RECT 407.400 626.700 409.200 633.600 ;
        RECT 413.400 626.700 415.200 633.600 ;
        RECT 428.400 626.700 430.200 633.600 ;
        RECT 434.400 626.700 436.200 633.600 ;
        RECT 452.400 626.700 454.200 633.600 ;
        RECT 460.500 626.700 462.300 639.600 ;
        RECT 475.800 626.700 477.600 633.600 ;
        RECT 481.800 626.700 483.600 633.600 ;
        RECT 494.400 626.700 496.200 633.600 ;
        RECT 500.400 626.700 502.200 633.600 ;
        RECT 518.400 626.700 520.200 633.600 ;
        RECT 524.400 626.700 526.200 633.600 ;
        RECT 539.400 626.700 541.200 639.600 ;
        RECT 562.800 626.700 564.600 639.600 ;
        RECT 578.400 626.700 580.200 633.600 ;
        RECT 586.500 626.700 588.300 639.600 ;
        RECT 604.800 626.700 606.600 633.600 ;
        RECT 625.800 626.700 627.600 633.000 ;
        RECT 631.800 626.700 633.600 633.600 ;
        RECT 646.800 626.700 648.600 633.600 ;
        RECT 652.800 626.700 654.600 633.600 ;
        RECT 665.400 626.700 667.200 633.600 ;
        RECT 671.400 626.700 673.200 633.600 ;
        RECT 697.800 626.700 699.600 637.500 ;
        RECT 716.400 626.700 718.200 637.500 ;
        RECT 748.800 626.700 750.600 637.800 ;
        RECT 764.400 626.700 766.200 633.600 ;
        RECT 770.400 626.700 772.200 633.000 ;
        RECT 788.400 626.700 790.200 633.600 ;
        RECT 794.400 626.700 796.200 633.000 ;
        RECT 815.400 626.700 817.200 633.600 ;
        RECT 836.400 626.700 838.200 637.800 ;
        RECT 862.800 626.700 864.600 633.000 ;
        RECT 868.800 626.700 870.600 633.600 ;
        RECT 884.400 626.700 886.200 637.800 ;
        RECT -9.450 624.300 896.400 626.700 ;
        RECT -9.450 548.700 -0.450 624.300 ;
        RECT 16.800 617.400 18.600 624.300 ;
        RECT 22.800 617.400 24.600 624.300 ;
        RECT 40.800 613.500 42.900 624.300 ;
        RECT 49.800 613.500 51.600 624.300 ;
        RECT 70.800 613.500 72.600 624.300 ;
        RECT 79.800 613.500 81.600 624.300 ;
        RECT 98.400 613.200 100.200 624.300 ;
        RECT 119.400 617.400 121.200 624.300 ;
        RECT 125.400 617.400 127.200 624.300 ;
        RECT 148.800 611.400 150.600 624.300 ;
        RECT 166.800 617.400 168.600 624.300 ;
        RECT 190.800 611.400 192.600 624.300 ;
        RECT 198.150 617.400 199.950 624.300 ;
        RECT 208.350 617.400 210.150 624.300 ;
        RECT 214.950 617.400 216.750 624.300 ;
        RECT 223.650 620.400 225.450 624.300 ;
        RECT 242.400 617.400 244.200 624.300 ;
        RECT 250.500 611.400 252.300 624.300 ;
        RECT 266.400 613.500 268.200 624.300 ;
        RECT 275.100 613.500 277.200 624.300 ;
        RECT 293.400 611.400 295.200 624.300 ;
        RECT 316.800 617.400 318.600 624.300 ;
        RECT 322.800 617.400 324.600 624.300 ;
        RECT 340.800 617.400 342.600 624.300 ;
        RECT 346.800 617.400 348.600 624.300 ;
        RECT 359.400 617.400 361.200 624.300 ;
        RECT 365.400 617.400 367.200 624.300 ;
        RECT 383.400 613.500 385.200 624.300 ;
        RECT 412.800 617.400 414.600 624.300 ;
        RECT 433.800 617.400 435.600 624.300 ;
        RECT 454.800 617.400 456.600 624.300 ;
        RECT 473.400 617.400 475.200 624.300 ;
        RECT 481.500 611.400 483.300 624.300 ;
        RECT 489.150 617.400 490.950 624.300 ;
        RECT 499.350 617.400 501.150 624.300 ;
        RECT 505.950 617.400 507.750 624.300 ;
        RECT 514.650 620.400 516.450 624.300 ;
        RECT 536.400 617.400 538.200 624.300 ;
        RECT 544.500 611.400 546.300 624.300 ;
        RECT 552.150 617.400 553.950 624.300 ;
        RECT 562.350 617.400 564.150 624.300 ;
        RECT 568.950 617.400 570.750 624.300 ;
        RECT 577.650 620.400 579.450 624.300 ;
        RECT 595.800 617.400 597.600 624.300 ;
        RECT 601.800 617.400 603.600 624.300 ;
        RECT 617.400 617.400 619.200 624.300 ;
        RECT 625.500 611.400 627.300 624.300 ;
        RECT 640.800 617.400 642.600 624.300 ;
        RECT 646.800 617.400 648.600 624.300 ;
        RECT 659.700 611.400 661.500 624.300 ;
        RECT 667.800 617.400 669.600 624.300 ;
        RECT 686.400 617.400 688.200 624.300 ;
        RECT 707.400 617.400 709.200 624.300 ;
        RECT 725.400 617.400 727.200 624.300 ;
        RECT 731.400 617.400 733.200 624.300 ;
        RECT 746.400 617.400 748.200 624.300 ;
        RECT 752.400 618.000 754.200 624.300 ;
        RECT 773.400 613.500 775.200 624.300 ;
        RECT 797.400 617.400 799.200 624.300 ;
        RECT 818.400 617.400 820.200 624.300 ;
        RECT 826.500 611.400 828.300 624.300 ;
        RECT 839.400 617.400 841.200 624.300 ;
        RECT 845.400 618.000 847.200 624.300 ;
        RECT 871.800 613.200 873.600 624.300 ;
        RECT 892.800 617.400 894.600 624.300 ;
        RECT 19.800 548.700 21.600 561.600 ;
        RECT 34.800 548.700 36.600 555.600 ;
        RECT 40.800 548.700 42.600 555.600 ;
        RECT 59.400 548.700 61.200 555.600 ;
        RECT 67.500 548.700 69.300 561.600 ;
        RECT 80.700 548.700 82.500 561.600 ;
        RECT 88.800 548.700 90.600 555.600 ;
        RECT 107.400 548.700 109.200 555.600 ;
        RECT 125.400 548.700 127.200 555.600 ;
        RECT 131.400 548.700 133.200 555.600 ;
        RECT 146.700 548.700 148.500 561.600 ;
        RECT 154.800 548.700 156.600 555.600 ;
        RECT 175.800 548.700 177.600 555.600 ;
        RECT 188.400 548.700 190.200 555.600 ;
        RECT 194.400 548.700 196.200 555.600 ;
        RECT 203.550 548.700 205.350 552.600 ;
        RECT 212.250 548.700 214.050 555.600 ;
        RECT 218.850 548.700 220.650 555.600 ;
        RECT 229.050 548.700 230.850 555.600 ;
        RECT 245.400 548.700 247.200 555.600 ;
        RECT 251.400 548.700 253.200 555.600 ;
        RECT 266.400 548.700 268.200 555.600 ;
        RECT 272.400 548.700 274.200 555.600 ;
        RECT 287.400 548.700 289.200 561.600 ;
        RECT 293.400 548.700 295.200 561.600 ;
        RECT 299.400 548.700 301.200 561.600 ;
        RECT 305.400 548.700 307.200 561.600 ;
        RECT 311.400 548.700 313.200 561.600 ;
        RECT 326.400 548.700 328.200 555.600 ;
        RECT 332.400 548.700 334.200 555.000 ;
        RECT 350.400 548.700 352.200 561.600 ;
        RECT 356.400 548.700 358.200 561.600 ;
        RECT 362.400 548.700 364.200 561.600 ;
        RECT 368.400 548.700 370.200 561.600 ;
        RECT 374.400 548.700 376.200 561.600 ;
        RECT 394.800 548.700 396.600 555.600 ;
        RECT 412.800 548.700 414.600 555.600 ;
        RECT 433.800 548.700 435.600 555.600 ;
        RECT 446.400 548.700 448.200 555.600 ;
        RECT 452.400 548.700 454.200 555.600 ;
        RECT 469.800 548.700 471.600 555.600 ;
        RECT 475.800 548.700 477.600 555.600 ;
        RECT 490.800 548.700 492.600 555.600 ;
        RECT 496.800 548.700 498.600 555.600 ;
        RECT 509.400 548.700 511.200 555.600 ;
        RECT 515.400 548.700 517.200 555.600 ;
        RECT 533.400 548.700 535.200 555.600 ;
        RECT 541.500 548.700 543.300 561.600 ;
        RECT 549.150 548.700 550.950 555.600 ;
        RECT 559.350 548.700 561.150 555.600 ;
        RECT 565.950 548.700 567.750 555.600 ;
        RECT 574.650 548.700 576.450 552.600 ;
        RECT 590.400 548.700 592.200 555.600 ;
        RECT 608.400 548.700 610.200 561.600 ;
        RECT 628.800 548.700 630.600 555.600 ;
        RECT 634.800 548.700 636.600 555.600 ;
        RECT 650.400 548.700 652.200 555.600 ;
        RECT 673.800 548.700 675.600 555.600 ;
        RECT 679.800 548.700 681.600 555.600 ;
        RECT 694.800 548.700 696.600 555.600 ;
        RECT 700.800 548.700 702.600 555.600 ;
        RECT 713.700 548.700 715.500 561.600 ;
        RECT 721.800 548.700 723.600 555.600 ;
        RECT 739.800 548.700 741.600 555.600 ;
        RECT 745.800 548.700 747.600 555.600 ;
        RECT 758.400 548.700 760.200 555.600 ;
        RECT 764.400 548.700 766.200 555.000 ;
        RECT 788.400 548.700 790.200 559.500 ;
        RECT 815.400 548.700 817.200 555.600 ;
        RECT 823.500 548.700 825.300 561.600 ;
        RECT 836.700 548.700 838.500 561.600 ;
        RECT 844.800 548.700 846.600 555.600 ;
        RECT 860.400 548.700 862.200 555.600 ;
        RECT 866.400 548.700 868.200 555.000 ;
        RECT -9.450 546.300 896.400 548.700 ;
        RECT -9.450 470.700 -0.450 546.300 ;
        RECT 11.700 533.400 13.500 546.300 ;
        RECT 19.800 539.400 21.600 546.300 ;
        RECT 37.800 539.400 39.600 546.300 ;
        RECT 43.800 539.400 45.600 546.300 ;
        RECT 61.800 535.500 63.600 546.300 ;
        RECT 70.800 535.500 72.600 546.300 ;
        RECT 80.550 542.400 82.350 546.300 ;
        RECT 89.250 539.400 91.050 546.300 ;
        RECT 95.850 539.400 97.650 546.300 ;
        RECT 106.050 539.400 107.850 546.300 ;
        RECT 122.700 533.400 124.500 546.300 ;
        RECT 130.800 539.400 132.600 546.300 ;
        RECT 146.400 539.400 148.200 546.300 ;
        RECT 152.400 539.400 154.200 546.300 ;
        RECT 161.550 542.400 163.350 546.300 ;
        RECT 170.250 539.400 172.050 546.300 ;
        RECT 176.850 539.400 178.650 546.300 ;
        RECT 187.050 539.400 188.850 546.300 ;
        RECT 203.400 539.400 205.200 546.300 ;
        RECT 221.700 533.400 223.500 546.300 ;
        RECT 229.800 539.400 231.600 546.300 ;
        RECT 251.400 539.400 253.200 546.300 ;
        RECT 269.400 539.400 271.200 546.300 ;
        RECT 275.400 539.400 277.200 546.300 ;
        RECT 290.400 539.400 292.200 546.300 ;
        RECT 316.800 533.400 318.600 546.300 ;
        RECT 323.550 542.400 325.350 546.300 ;
        RECT 332.250 539.400 334.050 546.300 ;
        RECT 338.850 539.400 340.650 546.300 ;
        RECT 349.050 539.400 350.850 546.300 ;
        RECT 367.800 539.400 369.600 546.300 ;
        RECT 373.800 539.400 375.600 546.300 ;
        RECT 391.800 533.400 393.600 546.300 ;
        RECT 407.400 539.400 409.200 546.300 ;
        RECT 415.500 533.400 417.300 546.300 ;
        RECT 423.150 539.400 424.950 546.300 ;
        RECT 433.350 539.400 435.150 546.300 ;
        RECT 439.950 539.400 441.750 546.300 ;
        RECT 448.650 542.400 450.450 546.300 ;
        RECT 464.400 539.400 466.200 546.300 ;
        RECT 470.400 539.400 472.200 546.300 ;
        RECT 487.800 539.400 489.600 546.300 ;
        RECT 493.800 539.400 495.600 546.300 ;
        RECT 509.400 539.400 511.200 546.300 ;
        RECT 517.500 533.400 519.300 546.300 ;
        RECT 525.150 539.400 526.950 546.300 ;
        RECT 535.350 539.400 537.150 546.300 ;
        RECT 541.950 539.400 543.750 546.300 ;
        RECT 550.650 542.400 552.450 546.300 ;
        RECT 566.700 533.400 568.500 546.300 ;
        RECT 574.800 539.400 576.600 546.300 ;
        RECT 595.800 539.400 597.600 546.300 ;
        RECT 601.800 539.400 603.600 546.300 ;
        RECT 619.800 540.000 621.600 546.300 ;
        RECT 625.800 539.400 627.600 546.300 ;
        RECT 638.400 539.400 640.200 546.300 ;
        RECT 658.800 539.400 660.600 546.300 ;
        RECT 664.800 539.400 666.600 546.300 ;
        RECT 677.700 533.400 679.500 546.300 ;
        RECT 685.800 539.400 687.600 546.300 ;
        RECT 704.400 539.400 706.200 546.300 ;
        RECT 722.700 533.400 724.500 546.300 ;
        RECT 730.800 539.400 732.600 546.300 ;
        RECT 746.400 539.400 748.200 546.300 ;
        RECT 752.400 539.400 754.200 546.300 ;
        RECT 772.800 539.400 774.600 546.300 ;
        RECT 778.800 539.400 780.600 546.300 ;
        RECT 793.800 539.400 795.600 546.300 ;
        RECT 799.800 539.400 801.600 546.300 ;
        RECT 812.400 539.400 814.200 546.300 ;
        RECT 818.400 539.400 820.200 546.300 ;
        RECT 844.800 535.200 846.600 546.300 ;
        RECT 860.700 533.400 862.500 546.300 ;
        RECT 868.800 539.400 870.600 546.300 ;
        RECT 6.150 470.700 7.950 477.600 ;
        RECT 16.350 470.700 18.150 477.600 ;
        RECT 22.950 470.700 24.750 477.600 ;
        RECT 31.650 470.700 33.450 474.600 ;
        RECT 47.400 470.700 49.200 477.600 ;
        RECT 53.400 470.700 55.200 477.600 ;
        RECT 70.800 470.700 72.600 477.600 ;
        RECT 76.800 470.700 78.600 477.600 ;
        RECT 83.550 470.700 85.350 474.600 ;
        RECT 92.250 470.700 94.050 477.600 ;
        RECT 98.850 470.700 100.650 477.600 ;
        RECT 109.050 470.700 110.850 477.600 ;
        RECT 133.800 470.700 135.600 481.800 ;
        RECT 149.400 470.700 151.200 483.600 ;
        RECT 170.400 470.700 172.200 477.600 ;
        RECT 191.400 470.700 193.200 477.600 ;
        RECT 197.400 470.700 199.200 477.600 ;
        RECT 217.800 470.700 219.600 477.600 ;
        RECT 223.800 470.700 225.600 477.600 ;
        RECT 236.400 470.700 238.200 477.600 ;
        RECT 242.400 470.700 244.200 477.600 ;
        RECT 260.400 470.700 262.200 477.600 ;
        RECT 268.500 470.700 270.300 483.600 ;
        RECT 275.550 470.700 277.350 474.600 ;
        RECT 284.250 470.700 286.050 477.600 ;
        RECT 290.850 470.700 292.650 477.600 ;
        RECT 301.050 470.700 302.850 477.600 ;
        RECT 317.700 470.700 319.500 483.600 ;
        RECT 325.800 470.700 327.600 477.600 ;
        RECT 344.400 470.700 346.200 477.600 ;
        RECT 352.500 470.700 354.300 483.600 ;
        RECT 359.550 470.700 361.350 474.600 ;
        RECT 368.250 470.700 370.050 477.600 ;
        RECT 374.850 470.700 376.650 477.600 ;
        RECT 385.050 470.700 386.850 477.600 ;
        RECT 403.800 470.700 405.600 477.600 ;
        RECT 409.800 470.700 411.600 477.600 ;
        RECT 425.400 470.700 427.200 477.600 ;
        RECT 433.500 470.700 435.300 483.600 ;
        RECT 449.400 470.700 451.200 477.600 ;
        RECT 457.500 470.700 459.300 483.600 ;
        RECT 465.150 470.700 466.950 477.600 ;
        RECT 475.350 470.700 477.150 477.600 ;
        RECT 481.950 470.700 483.750 477.600 ;
        RECT 490.650 470.700 492.450 474.600 ;
        RECT 506.700 470.700 508.500 483.600 ;
        RECT 514.800 470.700 516.600 477.600 ;
        RECT 530.400 470.700 532.200 483.600 ;
        RECT 551.400 470.700 553.200 477.600 ;
        RECT 571.800 470.700 573.600 477.600 ;
        RECT 577.800 470.700 579.600 477.600 ;
        RECT 593.400 470.700 595.200 477.600 ;
        RECT 601.500 470.700 603.300 483.600 ;
        RECT 614.700 470.700 616.500 483.600 ;
        RECT 622.800 470.700 624.600 477.600 ;
        RECT 638.400 470.700 640.200 477.600 ;
        RECT 644.400 470.700 646.200 477.600 ;
        RECT 659.400 470.700 661.200 477.600 ;
        RECT 665.400 470.700 667.200 477.000 ;
        RECT 683.400 470.700 685.200 477.600 ;
        RECT 689.400 470.700 691.200 477.600 ;
        RECT 707.700 470.700 709.500 483.600 ;
        RECT 715.800 470.700 717.600 477.600 ;
        RECT 734.400 470.700 736.200 481.800 ;
        RECT 760.800 470.700 762.600 477.600 ;
        RECT 766.800 470.700 768.600 477.600 ;
        RECT 782.400 470.700 784.200 481.500 ;
        RECT 806.400 470.700 808.200 483.600 ;
        RECT 827.400 470.700 829.200 477.600 ;
        RECT 833.400 470.700 835.200 477.600 ;
        RECT 851.400 470.700 853.200 477.600 ;
        RECT 859.500 470.700 861.300 483.600 ;
        RECT 872.400 470.700 874.200 477.600 ;
        RECT 878.400 470.700 880.200 477.000 ;
        RECT -9.450 468.300 896.400 470.700 ;
        RECT -9.450 392.700 -0.450 468.300 ;
        RECT 6.150 461.400 7.950 468.300 ;
        RECT 16.350 461.400 18.150 468.300 ;
        RECT 22.950 461.400 24.750 468.300 ;
        RECT 31.650 464.400 33.450 468.300 ;
        RECT 50.400 461.400 52.200 468.300 ;
        RECT 58.500 455.400 60.300 468.300 ;
        RECT 76.800 461.400 78.600 468.300 ;
        RECT 95.400 457.500 97.200 468.300 ;
        RECT 104.100 457.500 106.200 468.300 ;
        RECT 127.800 457.500 129.600 468.300 ;
        RECT 136.800 457.500 138.600 468.300 ;
        RECT 157.800 461.400 159.600 468.300 ;
        RECT 173.400 461.400 175.200 468.300 ;
        RECT 194.400 461.400 196.200 468.300 ;
        RECT 202.500 455.400 204.300 468.300 ;
        RECT 215.400 461.400 217.200 468.300 ;
        RECT 221.400 461.400 223.200 468.300 ;
        RECT 230.550 464.400 232.350 468.300 ;
        RECT 239.250 461.400 241.050 468.300 ;
        RECT 245.850 461.400 247.650 468.300 ;
        RECT 256.050 461.400 257.850 468.300 ;
        RECT 272.400 461.400 274.200 468.300 ;
        RECT 278.400 461.400 280.200 468.300 ;
        RECT 287.550 464.400 289.350 468.300 ;
        RECT 296.250 461.400 298.050 468.300 ;
        RECT 302.850 461.400 304.650 468.300 ;
        RECT 313.050 461.400 314.850 468.300 ;
        RECT 332.400 461.400 334.200 468.300 ;
        RECT 340.500 455.400 342.300 468.300 ;
        RECT 356.400 461.400 358.200 468.300 ;
        RECT 364.500 455.400 366.300 468.300 ;
        RECT 385.800 455.400 387.600 468.300 ;
        RECT 392.550 464.400 394.350 468.300 ;
        RECT 401.250 461.400 403.050 468.300 ;
        RECT 407.850 461.400 409.650 468.300 ;
        RECT 418.050 461.400 419.850 468.300 ;
        RECT 439.800 461.400 441.600 468.300 ;
        RECT 449.550 464.400 451.350 468.300 ;
        RECT 458.250 461.400 460.050 468.300 ;
        RECT 464.850 461.400 466.650 468.300 ;
        RECT 475.050 461.400 476.850 468.300 ;
        RECT 494.400 461.400 496.200 468.300 ;
        RECT 512.400 455.400 514.200 468.300 ;
        RECT 532.800 461.400 534.600 468.300 ;
        RECT 538.800 461.400 540.600 468.300 ;
        RECT 559.800 455.400 561.600 468.300 ;
        RECT 577.800 455.400 579.600 468.300 ;
        RECT 590.400 461.400 592.200 468.300 ;
        RECT 596.400 461.400 598.200 468.300 ;
        RECT 619.800 455.400 621.600 468.300 ;
        RECT 632.400 461.400 634.200 468.300 ;
        RECT 638.400 461.400 640.200 468.300 ;
        RECT 667.800 457.500 669.600 468.300 ;
        RECT 685.800 461.400 687.600 468.300 ;
        RECT 691.800 461.400 693.600 468.300 ;
        RECT 704.700 455.400 706.500 468.300 ;
        RECT 712.800 461.400 714.600 468.300 ;
        RECT 728.400 461.400 730.200 468.300 ;
        RECT 734.400 461.400 736.200 468.300 ;
        RECT 751.800 461.400 753.600 468.300 ;
        RECT 757.800 461.400 759.600 468.300 ;
        RECT 772.800 461.400 774.600 468.300 ;
        RECT 778.800 461.400 780.600 468.300 ;
        RECT 796.800 457.500 798.600 468.300 ;
        RECT 805.800 457.500 807.600 468.300 ;
        RECT 821.700 455.400 823.500 468.300 ;
        RECT 829.800 461.400 831.600 468.300 ;
        RECT 850.800 461.400 852.600 468.300 ;
        RECT 863.400 461.400 865.200 468.300 ;
        RECT 884.400 457.200 886.200 468.300 ;
        RECT 6.150 392.700 7.950 399.600 ;
        RECT 16.350 392.700 18.150 399.600 ;
        RECT 22.950 392.700 24.750 399.600 ;
        RECT 31.650 392.700 33.450 396.600 ;
        RECT 47.400 392.700 49.200 399.600 ;
        RECT 53.400 392.700 55.200 399.600 ;
        RECT 68.700 392.700 70.500 405.600 ;
        RECT 76.800 392.700 78.600 399.600 ;
        RECT 95.400 392.700 97.200 399.600 ;
        RECT 103.500 392.700 105.300 405.600 ;
        RECT 119.400 392.700 121.200 399.600 ;
        RECT 125.400 392.700 127.200 399.600 ;
        RECT 135.150 392.700 136.950 399.600 ;
        RECT 145.350 392.700 147.150 399.600 ;
        RECT 151.950 392.700 153.750 399.600 ;
        RECT 160.650 392.700 162.450 396.600 ;
        RECT 179.400 392.700 181.200 399.600 ;
        RECT 187.500 392.700 189.300 405.600 ;
        RECT 208.800 392.700 210.600 405.600 ;
        RECT 226.800 392.700 228.600 399.600 ;
        RECT 244.800 392.700 246.600 399.600 ;
        RECT 251.550 392.700 253.350 396.600 ;
        RECT 260.250 392.700 262.050 399.600 ;
        RECT 266.850 392.700 268.650 399.600 ;
        RECT 277.050 392.700 278.850 399.600 ;
        RECT 293.400 392.700 295.200 399.600 ;
        RECT 299.400 392.700 301.200 399.600 ;
        RECT 314.700 392.700 316.500 405.600 ;
        RECT 322.800 392.700 324.600 399.600 ;
        RECT 344.400 392.700 346.200 399.600 ;
        RECT 352.500 392.700 354.300 405.600 ;
        RECT 365.700 392.700 367.500 405.600 ;
        RECT 373.800 392.700 375.600 399.600 ;
        RECT 392.400 392.700 394.200 403.800 ;
        RECT 416.400 392.700 418.200 399.600 ;
        RECT 424.500 392.700 426.300 405.600 ;
        RECT 432.150 392.700 433.950 399.600 ;
        RECT 442.350 392.700 444.150 399.600 ;
        RECT 448.950 392.700 450.750 399.600 ;
        RECT 457.650 392.700 459.450 396.600 ;
        RECT 478.800 392.700 480.600 399.600 ;
        RECT 494.400 392.700 496.200 399.600 ;
        RECT 500.400 392.700 502.200 399.600 ;
        RECT 518.400 392.700 520.200 399.600 ;
        RECT 526.500 392.700 528.300 405.600 ;
        RECT 539.700 392.700 541.500 405.600 ;
        RECT 547.800 392.700 549.600 399.600 ;
        RECT 563.400 392.700 565.200 405.600 ;
        RECT 587.400 392.700 589.200 399.600 ;
        RECT 595.500 392.700 597.300 405.600 ;
        RECT 608.400 392.700 610.200 399.600 ;
        RECT 614.400 392.700 616.200 399.600 ;
        RECT 629.400 392.700 631.200 405.600 ;
        RECT 650.400 392.700 652.200 399.600 ;
        RECT 656.400 392.700 658.200 399.600 ;
        RECT 674.400 392.700 676.200 403.800 ;
        RECT 698.400 392.700 700.200 403.500 ;
        RECT 727.800 392.700 729.600 399.600 ;
        RECT 733.800 392.700 735.600 399.600 ;
        RECT 749.400 392.700 751.200 399.600 ;
        RECT 757.500 392.700 759.300 405.600 ;
        RECT 770.400 392.700 772.200 399.600 ;
        RECT 776.400 392.700 778.200 399.600 ;
        RECT 795.900 392.700 797.700 405.600 ;
        RECT 818.400 392.700 820.200 399.600 ;
        RECT 826.500 392.700 828.300 405.600 ;
        RECT 839.400 392.700 841.200 405.600 ;
        RECT 860.700 392.700 862.500 405.600 ;
        RECT 868.800 392.700 870.600 399.600 ;
        RECT 884.400 392.700 886.200 399.600 ;
        RECT 890.400 392.700 892.200 399.600 ;
        RECT -9.450 390.300 896.400 392.700 ;
        RECT -9.450 314.700 -0.450 390.300 ;
        RECT 6.150 383.400 7.950 390.300 ;
        RECT 16.350 383.400 18.150 390.300 ;
        RECT 22.950 383.400 24.750 390.300 ;
        RECT 31.650 386.400 33.450 390.300 ;
        RECT 50.400 383.400 52.200 390.300 ;
        RECT 58.500 377.400 60.300 390.300 ;
        RECT 73.800 383.400 75.600 390.300 ;
        RECT 79.800 383.400 81.600 390.300 ;
        RECT 86.550 386.400 88.350 390.300 ;
        RECT 95.250 383.400 97.050 390.300 ;
        RECT 101.850 383.400 103.650 390.300 ;
        RECT 112.050 383.400 113.850 390.300 ;
        RECT 133.800 383.400 135.600 390.300 ;
        RECT 157.800 377.400 159.600 390.300 ;
        RECT 170.700 377.400 172.500 390.300 ;
        RECT 178.800 383.400 180.600 390.300 ;
        RECT 202.800 377.400 204.600 390.300 ;
        RECT 209.550 386.400 211.350 390.300 ;
        RECT 218.250 383.400 220.050 390.300 ;
        RECT 224.850 383.400 226.650 390.300 ;
        RECT 235.050 383.400 236.850 390.300 ;
        RECT 251.700 377.400 253.500 390.300 ;
        RECT 259.800 383.400 261.600 390.300 ;
        RECT 278.400 383.400 280.200 390.300 ;
        RECT 284.400 383.400 286.200 390.300 ;
        RECT 299.400 377.400 301.200 390.300 ;
        RECT 325.800 383.400 327.600 390.300 ;
        RECT 338.700 377.400 340.500 390.300 ;
        RECT 346.800 383.400 348.600 390.300 ;
        RECT 356.550 386.400 358.350 390.300 ;
        RECT 365.250 383.400 367.050 390.300 ;
        RECT 371.850 383.400 373.650 390.300 ;
        RECT 382.050 383.400 383.850 390.300 ;
        RECT 392.550 386.400 394.350 390.300 ;
        RECT 401.250 383.400 403.050 390.300 ;
        RECT 407.850 383.400 409.650 390.300 ;
        RECT 418.050 383.400 419.850 390.300 ;
        RECT 429.150 383.400 430.950 390.300 ;
        RECT 439.350 383.400 441.150 390.300 ;
        RECT 445.950 383.400 447.750 390.300 ;
        RECT 454.650 386.400 456.450 390.300 ;
        RECT 470.400 377.400 472.200 390.300 ;
        RECT 497.400 379.200 499.200 390.300 ;
        RECT 528.300 377.400 530.100 390.300 ;
        RECT 548.700 377.400 550.500 390.300 ;
        RECT 556.800 383.400 558.600 390.300 ;
        RECT 572.700 377.400 574.500 390.300 ;
        RECT 580.800 383.400 582.600 390.300 ;
        RECT 596.400 377.400 598.200 390.300 ;
        RECT 606.900 377.400 608.700 390.300 ;
        RECT 623.400 383.400 625.200 390.300 ;
        RECT 644.400 383.400 646.200 390.300 ;
        RECT 652.500 377.400 654.300 390.300 ;
        RECT 665.400 383.400 667.200 390.300 ;
        RECT 671.400 383.400 673.200 390.300 ;
        RECT 692.400 379.500 694.200 390.300 ;
        RECT 701.100 379.500 703.200 390.300 ;
        RECT 722.400 383.400 724.200 390.300 ;
        RECT 730.500 377.400 732.300 390.300 ;
        RECT 743.400 377.400 745.200 390.300 ;
        RECT 767.400 379.500 769.200 390.300 ;
        RECT 776.400 379.500 778.200 390.300 ;
        RECT 797.400 383.400 799.200 390.300 ;
        RECT 805.500 377.400 807.300 390.300 ;
        RECT 818.400 383.400 820.200 390.300 ;
        RECT 824.400 383.400 826.200 390.300 ;
        RECT 839.700 377.400 841.500 390.300 ;
        RECT 847.800 383.400 849.600 390.300 ;
        RECT 866.400 379.200 868.200 390.300 ;
        RECT 6.150 314.700 7.950 321.600 ;
        RECT 16.350 314.700 18.150 321.600 ;
        RECT 22.950 314.700 24.750 321.600 ;
        RECT 31.650 314.700 33.450 318.600 ;
        RECT 47.400 314.700 49.200 321.600 ;
        RECT 53.400 314.700 55.200 321.600 ;
        RECT 82.800 314.700 84.600 325.500 ;
        RECT 101.400 314.700 103.200 321.600 ;
        RECT 107.400 314.700 109.200 321.600 ;
        RECT 125.400 314.700 127.200 321.600 ;
        RECT 133.500 314.700 135.300 327.600 ;
        RECT 148.800 314.700 150.600 321.600 ;
        RECT 154.800 314.700 156.600 321.600 ;
        RECT 169.800 314.700 171.600 321.600 ;
        RECT 175.800 314.700 177.600 321.600 ;
        RECT 188.400 314.700 190.200 321.600 ;
        RECT 209.400 314.700 211.200 321.600 ;
        RECT 235.800 314.700 237.600 327.600 ;
        RECT 251.400 314.700 253.200 325.800 ;
        RECT 272.400 314.700 274.200 327.600 ;
        RECT 288.150 314.700 289.950 321.600 ;
        RECT 298.350 314.700 300.150 321.600 ;
        RECT 304.950 314.700 306.750 321.600 ;
        RECT 313.650 314.700 315.450 318.600 ;
        RECT 329.400 314.700 331.200 321.600 ;
        RECT 347.400 314.700 349.200 327.600 ;
        RECT 353.400 314.700 355.200 327.600 ;
        RECT 359.400 314.700 361.200 327.600 ;
        RECT 365.400 314.700 367.200 327.600 ;
        RECT 371.400 314.700 373.200 327.600 ;
        RECT 394.800 314.700 396.600 327.600 ;
        RECT 415.800 314.700 417.600 325.800 ;
        RECT 436.800 314.700 438.600 321.600 ;
        RECT 455.400 314.700 457.200 321.600 ;
        RECT 481.800 314.700 483.600 327.600 ;
        RECT 494.400 314.700 496.200 321.600 ;
        RECT 500.400 314.700 502.200 321.000 ;
        RECT 518.700 314.700 520.500 327.600 ;
        RECT 526.800 314.700 528.600 321.600 ;
        RECT 542.700 314.700 544.500 327.600 ;
        RECT 550.800 314.700 552.600 321.600 ;
        RECT 568.800 314.700 570.600 321.600 ;
        RECT 574.800 314.700 576.600 321.600 ;
        RECT 593.400 314.700 595.200 325.500 ;
        RECT 602.400 314.700 604.200 325.500 ;
        RECT 623.400 314.700 625.200 321.600 ;
        RECT 631.500 314.700 633.300 327.600 ;
        RECT 649.800 314.700 651.600 321.000 ;
        RECT 655.800 314.700 657.600 321.600 ;
        RECT 671.400 314.700 673.200 325.800 ;
        RECT 697.800 314.700 699.600 321.000 ;
        RECT 703.800 314.700 705.600 321.600 ;
        RECT 716.400 314.700 718.200 321.600 ;
        RECT 722.400 314.700 724.200 321.000 ;
        RECT 748.800 314.700 750.600 325.800 ;
        RECT 767.400 314.700 769.200 321.600 ;
        RECT 773.400 314.700 775.200 321.000 ;
        RECT 794.400 314.700 796.200 325.800 ;
        RECT 818.400 314.700 820.200 321.600 ;
        RECT 826.500 314.700 828.300 327.600 ;
        RECT 839.700 314.700 841.500 327.600 ;
        RECT 847.800 314.700 849.600 321.600 ;
        RECT 863.400 314.700 865.200 321.600 ;
        RECT 869.400 314.700 871.200 321.000 ;
        RECT -9.450 312.300 896.400 314.700 ;
        RECT -9.450 236.700 -0.450 312.300 ;
        RECT 13.800 299.400 15.600 312.300 ;
        RECT 19.800 299.400 21.600 312.300 ;
        RECT 25.800 299.400 27.600 312.300 ;
        RECT 31.800 299.400 33.600 312.300 ;
        RECT 37.800 299.400 39.600 312.300 ;
        RECT 61.800 301.500 63.600 312.300 ;
        RECT 88.800 301.500 90.600 312.300 ;
        RECT 98.550 308.400 100.350 312.300 ;
        RECT 107.250 305.400 109.050 312.300 ;
        RECT 113.850 305.400 115.650 312.300 ;
        RECT 124.050 305.400 125.850 312.300 ;
        RECT 135.150 305.400 136.950 312.300 ;
        RECT 145.350 305.400 147.150 312.300 ;
        RECT 151.950 305.400 153.750 312.300 ;
        RECT 160.650 308.400 162.450 312.300 ;
        RECT 171.150 305.400 172.950 312.300 ;
        RECT 181.350 305.400 183.150 312.300 ;
        RECT 187.950 305.400 189.750 312.300 ;
        RECT 196.650 308.400 198.450 312.300 ;
        RECT 214.800 305.400 216.600 312.300 ;
        RECT 220.800 305.400 222.600 312.300 ;
        RECT 235.800 305.400 237.600 312.300 ;
        RECT 241.800 305.400 243.600 312.300 ;
        RECT 248.550 308.400 250.350 312.300 ;
        RECT 257.250 305.400 259.050 312.300 ;
        RECT 263.850 305.400 265.650 312.300 ;
        RECT 274.050 305.400 275.850 312.300 ;
        RECT 290.700 299.400 292.500 312.300 ;
        RECT 298.800 305.400 300.600 312.300 ;
        RECT 316.800 305.400 318.600 312.300 ;
        RECT 322.800 305.400 324.600 312.300 ;
        RECT 343.800 299.400 345.600 312.300 ;
        RECT 350.550 308.400 352.350 312.300 ;
        RECT 359.250 305.400 361.050 312.300 ;
        RECT 365.850 305.400 367.650 312.300 ;
        RECT 376.050 305.400 377.850 312.300 ;
        RECT 400.800 301.200 402.600 312.300 ;
        RECT 419.400 305.400 421.200 312.300 ;
        RECT 437.400 305.400 439.200 312.300 ;
        RECT 443.400 305.400 445.200 312.300 ;
        RECT 466.800 299.400 468.600 312.300 ;
        RECT 482.400 301.200 484.200 312.300 ;
        RECT 498.150 305.400 499.950 312.300 ;
        RECT 508.350 305.400 510.150 312.300 ;
        RECT 514.950 305.400 516.750 312.300 ;
        RECT 523.650 308.400 525.450 312.300 ;
        RECT 544.800 305.400 546.600 312.300 ;
        RECT 550.800 305.400 552.600 312.300 ;
        RECT 568.800 305.400 570.600 312.300 ;
        RECT 585.900 299.400 587.700 312.300 ;
        RECT 605.400 305.400 607.200 312.300 ;
        RECT 629.400 301.200 631.200 312.300 ;
        RECT 655.800 305.400 657.600 312.300 ;
        RECT 668.400 305.400 670.200 312.300 ;
        RECT 686.400 305.400 688.200 312.300 ;
        RECT 692.400 306.000 694.200 312.300 ;
        RECT 713.700 299.400 715.500 312.300 ;
        RECT 721.800 305.400 723.600 312.300 ;
        RECT 737.700 299.400 739.500 312.300 ;
        RECT 745.800 305.400 747.600 312.300 ;
        RECT 761.400 305.400 763.200 312.300 ;
        RECT 767.400 306.000 769.200 312.300 ;
        RECT 785.400 305.400 787.200 312.300 ;
        RECT 791.400 306.000 793.200 312.300 ;
        RECT 812.400 305.400 814.200 312.300 ;
        RECT 833.400 301.200 835.200 312.300 ;
        RECT 859.800 306.000 861.600 312.300 ;
        RECT 865.800 305.400 867.600 312.300 ;
        RECT 881.400 301.200 883.200 312.300 ;
        RECT 13.800 236.700 15.600 249.600 ;
        RECT 19.800 236.700 21.600 249.600 ;
        RECT 25.800 236.700 27.600 249.600 ;
        RECT 31.800 236.700 33.600 249.600 ;
        RECT 37.800 236.700 39.600 249.600 ;
        RECT 53.400 236.700 55.200 243.600 ;
        RECT 61.500 236.700 63.300 249.600 ;
        RECT 82.800 236.700 84.600 243.600 ;
        RECT 103.800 236.700 105.600 249.600 ;
        RECT 127.800 236.700 129.600 247.500 ;
        RECT 145.800 236.700 147.600 243.600 ;
        RECT 151.800 236.700 153.600 243.600 ;
        RECT 158.550 236.700 160.350 240.600 ;
        RECT 167.250 236.700 169.050 243.600 ;
        RECT 173.850 236.700 175.650 243.600 ;
        RECT 184.050 236.700 185.850 243.600 ;
        RECT 203.400 236.700 205.200 243.600 ;
        RECT 211.500 236.700 213.300 249.600 ;
        RECT 224.400 236.700 226.200 243.600 ;
        RECT 230.400 236.700 232.200 243.000 ;
        RECT 256.800 236.700 258.600 249.600 ;
        RECT 263.550 236.700 265.350 240.600 ;
        RECT 272.250 236.700 274.050 243.600 ;
        RECT 278.850 236.700 280.650 243.600 ;
        RECT 289.050 236.700 290.850 243.600 ;
        RECT 305.400 236.700 307.200 249.600 ;
        RECT 311.400 236.700 313.200 249.600 ;
        RECT 317.400 236.700 319.200 249.600 ;
        RECT 332.400 236.700 334.200 243.600 ;
        RECT 353.400 236.700 355.200 243.600 ;
        RECT 366.150 236.700 367.950 243.600 ;
        RECT 376.350 236.700 378.150 243.600 ;
        RECT 382.950 236.700 384.750 243.600 ;
        RECT 391.650 236.700 393.450 240.600 ;
        RECT 407.400 236.700 409.200 243.600 ;
        RECT 425.700 236.700 427.500 249.600 ;
        RECT 433.800 236.700 435.600 243.600 ;
        RECT 452.400 236.700 454.200 243.600 ;
        RECT 465.150 236.700 466.950 243.600 ;
        RECT 475.350 236.700 477.150 243.600 ;
        RECT 481.950 236.700 483.750 243.600 ;
        RECT 490.650 236.700 492.450 240.600 ;
        RECT 506.700 236.700 508.500 249.600 ;
        RECT 514.800 236.700 516.600 243.600 ;
        RECT 530.400 236.700 532.200 243.600 ;
        RECT 536.400 236.700 538.200 243.600 ;
        RECT 553.800 236.700 555.600 243.600 ;
        RECT 559.800 236.700 561.600 243.600 ;
        RECT 579.300 236.700 581.100 249.600 ;
        RECT 598.800 236.700 600.600 243.600 ;
        RECT 604.800 236.700 606.600 243.600 ;
        RECT 617.700 236.700 619.500 249.600 ;
        RECT 625.800 236.700 627.600 243.600 ;
        RECT 649.800 236.700 651.900 247.500 ;
        RECT 658.800 236.700 660.600 247.500 ;
        RECT 676.800 236.700 678.600 243.600 ;
        RECT 682.800 236.700 684.600 243.600 ;
        RECT 703.800 236.700 705.600 247.800 ;
        RECT 719.400 236.700 721.200 243.600 ;
        RECT 725.400 236.700 727.200 243.000 ;
        RECT 748.800 236.700 750.600 243.000 ;
        RECT 754.800 236.700 756.600 243.600 ;
        RECT 769.800 236.700 771.600 243.600 ;
        RECT 775.800 236.700 777.600 243.600 ;
        RECT 788.400 236.700 790.200 243.600 ;
        RECT 794.400 236.700 796.200 243.000 ;
        RECT 815.400 236.700 817.200 243.600 ;
        RECT 823.500 236.700 825.300 249.600 ;
        RECT 836.400 236.700 838.200 243.600 ;
        RECT 842.400 236.700 844.200 243.000 ;
        RECT 868.800 236.700 870.600 247.800 ;
        RECT -9.450 234.300 896.400 236.700 ;
        RECT -9.450 158.700 -0.450 234.300 ;
        RECT 6.150 227.400 7.950 234.300 ;
        RECT 16.350 227.400 18.150 234.300 ;
        RECT 22.950 227.400 24.750 234.300 ;
        RECT 31.650 230.400 33.450 234.300 ;
        RECT 50.400 227.400 52.200 234.300 ;
        RECT 58.500 221.400 60.300 234.300 ;
        RECT 71.400 227.400 73.200 234.300 ;
        RECT 92.400 227.400 94.200 234.300 ;
        RECT 100.500 221.400 102.300 234.300 ;
        RECT 113.400 221.400 115.200 234.300 ;
        RECT 142.800 221.400 144.600 234.300 ;
        RECT 158.400 227.400 160.200 234.300 ;
        RECT 166.500 221.400 168.300 234.300 ;
        RECT 179.400 221.400 181.200 234.300 ;
        RECT 206.400 227.400 208.200 234.300 ;
        RECT 214.500 221.400 216.300 234.300 ;
        RECT 221.550 230.400 223.350 234.300 ;
        RECT 230.250 227.400 232.050 234.300 ;
        RECT 236.850 227.400 238.650 234.300 ;
        RECT 247.050 227.400 248.850 234.300 ;
        RECT 263.400 227.400 265.200 234.300 ;
        RECT 269.400 227.400 271.200 234.300 ;
        RECT 287.400 227.400 289.200 234.300 ;
        RECT 295.500 221.400 297.300 234.300 ;
        RECT 311.400 227.400 313.200 234.300 ;
        RECT 319.500 221.400 321.300 234.300 ;
        RECT 340.800 221.400 342.600 234.300 ;
        RECT 358.800 227.400 360.600 234.300 ;
        RECT 376.800 227.400 378.600 234.300 ;
        RECT 382.800 227.400 384.600 234.300 ;
        RECT 402.300 221.400 404.100 234.300 ;
        RECT 419.400 227.400 421.200 234.300 ;
        RECT 425.400 227.400 427.200 234.300 ;
        RECT 435.150 227.400 436.950 234.300 ;
        RECT 445.350 227.400 447.150 234.300 ;
        RECT 451.950 227.400 453.750 234.300 ;
        RECT 460.650 230.400 462.450 234.300 ;
        RECT 476.400 227.400 478.200 234.300 ;
        RECT 494.700 221.400 496.500 234.300 ;
        RECT 502.800 227.400 504.600 234.300 ;
        RECT 518.400 227.400 520.200 234.300 ;
        RECT 524.400 227.400 526.200 234.300 ;
        RECT 533.550 230.400 535.350 234.300 ;
        RECT 542.250 227.400 544.050 234.300 ;
        RECT 548.850 227.400 550.650 234.300 ;
        RECT 559.050 227.400 560.850 234.300 ;
        RECT 578.400 227.400 580.200 234.300 ;
        RECT 584.400 227.400 586.200 234.300 ;
        RECT 602.400 227.400 604.200 234.300 ;
        RECT 610.500 221.400 612.300 234.300 ;
        RECT 623.400 227.400 625.200 234.300 ;
        RECT 629.400 227.400 631.200 234.300 ;
        RECT 647.400 227.400 649.200 234.300 ;
        RECT 653.400 227.400 655.200 234.300 ;
        RECT 679.800 223.200 681.600 234.300 ;
        RECT 698.400 223.500 700.200 234.300 ;
        RECT 707.400 223.500 709.200 234.300 ;
        RECT 730.800 223.500 732.600 234.300 ;
        RECT 739.800 223.500 741.600 234.300 ;
        RECT 763.800 223.200 765.600 234.300 ;
        RECT 784.800 227.400 786.600 234.300 ;
        RECT 797.400 227.400 799.200 234.300 ;
        RECT 803.400 227.400 805.200 234.300 ;
        RECT 823.800 227.400 825.600 234.300 ;
        RECT 829.800 227.400 831.600 234.300 ;
        RECT 842.400 227.400 844.200 234.300 ;
        RECT 848.400 228.000 850.200 234.300 ;
        RECT 869.400 227.400 871.200 234.300 ;
        RECT 877.500 221.400 879.300 234.300 ;
        RECT 14.400 158.700 16.200 165.600 ;
        RECT 22.500 158.700 24.300 171.600 ;
        RECT 35.400 158.700 37.200 165.600 ;
        RECT 41.400 158.700 43.200 165.600 ;
        RECT 59.400 158.700 61.200 165.600 ;
        RECT 67.500 158.700 69.300 171.600 ;
        RECT 80.700 158.700 82.500 171.600 ;
        RECT 88.800 158.700 90.600 165.600 ;
        RECT 98.550 158.700 100.350 162.600 ;
        RECT 107.250 158.700 109.050 165.600 ;
        RECT 113.850 158.700 115.650 165.600 ;
        RECT 124.050 158.700 125.850 165.600 ;
        RECT 140.400 158.700 142.200 165.600 ;
        RECT 146.400 158.700 148.200 165.600 ;
        RECT 164.400 158.700 166.200 165.600 ;
        RECT 172.500 158.700 174.300 171.600 ;
        RECT 185.400 158.700 187.200 165.600 ;
        RECT 191.400 158.700 193.200 165.600 ;
        RECT 208.800 158.700 210.600 165.600 ;
        RECT 214.800 158.700 216.600 165.600 ;
        RECT 221.550 158.700 223.350 162.600 ;
        RECT 230.250 158.700 232.050 165.600 ;
        RECT 236.850 158.700 238.650 165.600 ;
        RECT 247.050 158.700 248.850 165.600 ;
        RECT 266.400 158.700 268.200 165.600 ;
        RECT 274.500 158.700 276.300 171.600 ;
        RECT 295.800 158.700 297.600 169.800 ;
        RECT 319.800 158.700 321.600 171.600 ;
        RECT 337.800 158.700 339.600 169.500 ;
        RECT 346.800 158.700 348.600 169.500 ;
        RECT 362.700 158.700 364.500 171.600 ;
        RECT 370.800 158.700 372.600 165.600 ;
        RECT 391.800 158.700 393.600 165.600 ;
        RECT 407.400 158.700 409.200 165.600 ;
        RECT 415.500 158.700 417.300 171.600 ;
        RECT 431.400 158.700 433.200 171.600 ;
        RECT 452.400 158.700 454.200 165.600 ;
        RECT 475.800 158.700 477.600 165.600 ;
        RECT 482.550 158.700 484.350 162.600 ;
        RECT 491.250 158.700 493.050 165.600 ;
        RECT 497.850 158.700 499.650 165.600 ;
        RECT 508.050 158.700 509.850 165.600 ;
        RECT 524.400 158.700 526.200 171.600 ;
        RECT 545.400 158.700 547.200 165.600 ;
        RECT 551.400 158.700 553.200 165.600 ;
        RECT 561.150 158.700 562.950 165.600 ;
        RECT 571.350 158.700 573.150 165.600 ;
        RECT 577.950 158.700 579.750 165.600 ;
        RECT 586.650 158.700 588.450 162.600 ;
        RECT 605.400 158.700 607.200 165.600 ;
        RECT 613.500 158.700 615.300 171.600 ;
        RECT 626.400 158.700 628.200 165.600 ;
        RECT 632.400 158.700 634.200 165.600 ;
        RECT 650.400 158.700 652.200 165.600 ;
        RECT 658.500 158.700 660.300 171.600 ;
        RECT 677.400 158.700 679.200 169.500 ;
        RECT 701.400 158.700 703.200 171.600 ;
        RECT 722.400 158.700 724.200 165.600 ;
        RECT 740.700 158.700 742.500 171.600 ;
        RECT 748.800 158.700 750.600 165.600 ;
        RECT 764.400 158.700 766.200 165.600 ;
        RECT 785.400 158.700 787.200 169.800 ;
        RECT 814.800 158.700 816.600 171.600 ;
        RECT 827.400 158.700 829.200 165.600 ;
        RECT 833.400 158.700 835.200 165.600 ;
        RECT 848.400 158.700 850.200 165.600 ;
        RECT 854.400 158.700 856.200 165.600 ;
        RECT 869.400 158.700 871.200 165.600 ;
        RECT 875.400 158.700 877.200 165.600 ;
        RECT -9.450 156.300 896.400 158.700 ;
        RECT -9.450 80.700 -0.450 156.300 ;
        RECT 16.800 149.400 18.600 156.300 ;
        RECT 32.400 143.400 34.200 156.300 ;
        RECT 38.400 143.400 40.200 156.300 ;
        RECT 44.400 143.400 46.200 156.300 ;
        RECT 50.400 143.400 52.200 156.300 ;
        RECT 56.400 143.400 58.200 156.300 ;
        RECT 73.800 149.400 75.600 156.300 ;
        RECT 79.800 149.400 81.600 156.300 ;
        RECT 92.400 149.400 94.200 156.300 ;
        RECT 98.400 149.400 100.200 156.300 ;
        RECT 122.400 149.400 124.200 156.300 ;
        RECT 130.500 143.400 132.300 156.300 ;
        RECT 143.700 143.400 145.500 156.300 ;
        RECT 151.800 149.400 153.600 156.300 ;
        RECT 172.800 149.400 174.600 156.300 ;
        RECT 193.800 149.400 195.600 156.300 ;
        RECT 200.550 152.400 202.350 156.300 ;
        RECT 209.250 149.400 211.050 156.300 ;
        RECT 215.850 149.400 217.650 156.300 ;
        RECT 226.050 149.400 227.850 156.300 ;
        RECT 242.700 143.400 244.500 156.300 ;
        RECT 250.800 149.400 252.600 156.300 ;
        RECT 268.800 149.400 270.600 156.300 ;
        RECT 274.800 149.400 276.600 156.300 ;
        RECT 290.400 149.400 292.200 156.300 ;
        RECT 298.500 143.400 300.300 156.300 ;
        RECT 305.550 152.400 307.350 156.300 ;
        RECT 314.250 149.400 316.050 156.300 ;
        RECT 320.850 149.400 322.650 156.300 ;
        RECT 331.050 149.400 332.850 156.300 ;
        RECT 352.800 149.400 354.600 156.300 ;
        RECT 368.400 149.400 370.200 156.300 ;
        RECT 374.400 149.400 376.200 156.300 ;
        RECT 389.400 143.400 391.200 156.300 ;
        RECT 395.400 143.400 397.200 156.300 ;
        RECT 401.400 143.400 403.200 156.300 ;
        RECT 407.400 143.400 409.200 156.300 ;
        RECT 413.400 143.400 415.200 156.300 ;
        RECT 430.800 149.400 432.600 156.300 ;
        RECT 436.800 149.400 438.600 156.300 ;
        RECT 452.400 149.400 454.200 156.300 ;
        RECT 460.500 143.400 462.300 156.300 ;
        RECT 467.550 152.400 469.350 156.300 ;
        RECT 476.250 149.400 478.050 156.300 ;
        RECT 482.850 149.400 484.650 156.300 ;
        RECT 493.050 149.400 494.850 156.300 ;
        RECT 512.400 145.500 514.200 156.300 ;
        RECT 543.300 143.400 545.100 156.300 ;
        RECT 566.400 145.200 568.200 156.300 ;
        RECT 587.400 149.400 589.200 156.300 ;
        RECT 610.800 149.400 612.600 156.300 ;
        RECT 617.550 152.400 619.350 156.300 ;
        RECT 626.250 149.400 628.050 156.300 ;
        RECT 632.850 149.400 634.650 156.300 ;
        RECT 643.050 149.400 644.850 156.300 ;
        RECT 664.800 149.400 666.600 156.300 ;
        RECT 671.550 152.400 673.350 156.300 ;
        RECT 680.250 149.400 682.050 156.300 ;
        RECT 686.850 149.400 688.650 156.300 ;
        RECT 697.050 149.400 698.850 156.300 ;
        RECT 713.400 143.400 715.200 156.300 ;
        RECT 723.900 143.400 725.700 156.300 ;
        RECT 740.700 143.400 742.500 156.300 ;
        RECT 748.800 149.400 750.600 156.300 ;
        RECT 772.800 145.200 774.600 156.300 ;
        RECT 788.700 143.400 790.500 156.300 ;
        RECT 796.800 149.400 798.600 156.300 ;
        RECT 817.800 149.400 819.600 156.300 ;
        RECT 833.400 149.400 835.200 156.300 ;
        RECT 841.500 143.400 843.300 156.300 ;
        RECT 859.800 149.400 861.600 156.300 ;
        RECT 872.400 149.400 874.200 156.300 ;
        RECT 878.400 150.000 880.200 156.300 ;
        RECT 16.800 80.700 18.600 91.500 ;
        RECT 25.800 80.700 27.600 91.500 ;
        RECT 49.800 80.700 51.600 93.600 ;
        RECT 64.800 80.700 66.600 87.600 ;
        RECT 70.800 80.700 72.600 87.600 ;
        RECT 91.800 80.700 93.600 93.600 ;
        RECT 104.400 80.700 106.200 87.600 ;
        RECT 130.800 80.700 132.600 93.600 ;
        RECT 146.400 80.700 148.200 87.600 ;
        RECT 172.800 80.700 174.600 93.600 ;
        RECT 193.800 80.700 195.600 93.600 ;
        RECT 214.800 80.700 216.600 87.600 ;
        RECT 221.550 80.700 223.350 84.600 ;
        RECT 230.250 80.700 232.050 87.600 ;
        RECT 236.850 80.700 238.650 87.600 ;
        RECT 247.050 80.700 248.850 87.600 ;
        RECT 263.700 80.700 265.500 93.600 ;
        RECT 271.800 80.700 273.600 87.600 ;
        RECT 292.800 80.700 294.600 87.600 ;
        RECT 299.550 80.700 301.350 84.600 ;
        RECT 308.250 80.700 310.050 87.600 ;
        RECT 314.850 80.700 316.650 87.600 ;
        RECT 325.050 80.700 326.850 87.600 ;
        RECT 341.400 80.700 343.200 93.600 ;
        RECT 351.900 80.700 353.700 93.600 ;
        RECT 376.800 80.700 378.600 93.600 ;
        RECT 383.550 80.700 385.350 84.600 ;
        RECT 392.250 80.700 394.050 87.600 ;
        RECT 398.850 80.700 400.650 87.600 ;
        RECT 409.050 80.700 410.850 87.600 ;
        RECT 433.800 80.700 435.600 91.800 ;
        RECT 457.800 80.700 459.600 93.600 ;
        RECT 473.400 80.700 475.200 87.600 ;
        RECT 481.500 80.700 483.300 93.600 ;
        RECT 494.400 80.700 496.200 87.600 ;
        RECT 520.800 80.700 522.600 93.600 ;
        RECT 533.700 80.700 535.500 93.600 ;
        RECT 541.800 80.700 543.600 87.600 ;
        RECT 562.800 80.700 564.600 87.600 ;
        RECT 575.400 80.700 577.200 87.600 ;
        RECT 581.400 80.700 583.200 87.600 ;
        RECT 601.800 80.700 603.600 87.600 ;
        RECT 607.800 80.700 609.600 87.600 ;
        RECT 623.400 80.700 625.200 93.600 ;
        RECT 649.800 80.700 651.600 87.600 ;
        RECT 656.550 80.700 658.350 84.600 ;
        RECT 665.250 80.700 667.050 87.600 ;
        RECT 671.850 80.700 673.650 87.600 ;
        RECT 682.050 80.700 683.850 87.600 ;
        RECT 703.800 80.700 705.600 87.000 ;
        RECT 709.800 80.700 711.600 87.600 ;
        RECT 722.400 80.700 724.200 87.600 ;
        RECT 728.400 80.700 730.200 87.600 ;
        RECT 746.400 80.700 748.200 91.500 ;
        RECT 755.400 80.700 757.200 91.500 ;
        RECT 776.400 80.700 778.200 91.800 ;
        RECT 800.400 80.700 802.200 91.800 ;
        RECT 829.800 80.700 831.600 93.600 ;
        RECT 842.400 80.700 844.200 93.600 ;
        RECT 863.400 80.700 865.200 93.600 ;
        RECT 884.400 80.700 886.200 87.600 ;
        RECT -9.450 78.300 896.400 80.700 ;
        RECT -9.450 2.700 -0.450 78.300 ;
        RECT 19.800 65.400 21.600 78.300 ;
        RECT 32.400 65.400 34.200 78.300 ;
        RECT 56.400 67.200 58.200 78.300 ;
        RECT 80.400 71.400 82.200 78.300 ;
        RECT 88.500 65.400 90.300 78.300 ;
        RECT 101.400 71.400 103.200 78.300 ;
        RECT 107.400 71.400 109.200 78.300 ;
        RECT 122.400 71.400 124.200 78.300 ;
        RECT 128.400 71.400 130.200 78.300 ;
        RECT 137.550 74.400 139.350 78.300 ;
        RECT 146.250 71.400 148.050 78.300 ;
        RECT 152.850 71.400 154.650 78.300 ;
        RECT 163.050 71.400 164.850 78.300 ;
        RECT 179.400 65.400 181.200 78.300 ;
        RECT 208.800 67.200 210.600 78.300 ;
        RECT 224.700 65.400 226.500 78.300 ;
        RECT 232.800 71.400 234.600 78.300 ;
        RECT 242.550 74.400 244.350 78.300 ;
        RECT 251.250 71.400 253.050 78.300 ;
        RECT 257.850 71.400 259.650 78.300 ;
        RECT 268.050 71.400 269.850 78.300 ;
        RECT 284.400 71.400 286.200 78.300 ;
        RECT 304.800 71.400 306.600 78.300 ;
        RECT 310.800 71.400 312.600 78.300 ;
        RECT 328.800 72.000 330.600 78.300 ;
        RECT 334.800 71.400 336.600 78.300 ;
        RECT 347.400 65.400 349.200 78.300 ;
        RECT 371.400 71.400 373.200 78.300 ;
        RECT 379.500 65.400 381.300 78.300 ;
        RECT 397.800 71.400 399.600 78.300 ;
        RECT 410.700 65.400 412.500 78.300 ;
        RECT 418.800 71.400 420.600 78.300 ;
        RECT 434.400 71.400 436.200 78.300 ;
        RECT 452.700 65.400 454.500 78.300 ;
        RECT 460.800 71.400 462.600 78.300 ;
        RECT 481.800 71.400 483.600 78.300 ;
        RECT 502.800 67.200 504.600 78.300 ;
        RECT 526.800 71.400 528.600 78.300 ;
        RECT 544.800 71.400 546.600 78.300 ;
        RECT 565.800 67.200 567.600 78.300 ;
        RECT 589.800 65.400 591.600 78.300 ;
        RECT 610.800 65.400 612.600 78.300 ;
        RECT 628.800 71.400 630.600 78.300 ;
        RECT 641.400 65.400 643.200 78.300 ;
        RECT 667.800 72.000 669.600 78.300 ;
        RECT 673.800 71.400 675.600 78.300 ;
        RECT 691.800 72.000 693.600 78.300 ;
        RECT 697.800 71.400 699.600 78.300 ;
        RECT 710.400 71.400 712.200 78.300 ;
        RECT 728.400 71.400 730.200 78.300 ;
        RECT 734.400 72.000 736.200 78.300 ;
        RECT 754.800 71.400 756.600 78.300 ;
        RECT 760.800 71.400 762.600 78.300 ;
        RECT 773.400 71.400 775.200 78.300 ;
        RECT 779.400 72.000 781.200 78.300 ;
        RECT 797.400 71.400 799.200 78.300 ;
        RECT 815.400 71.400 817.200 78.300 ;
        RECT 836.400 71.400 838.200 78.300 ;
        RECT 854.400 71.400 856.200 78.300 ;
        RECT 860.400 72.000 862.200 78.300 ;
        RECT 878.400 71.400 880.200 78.300 ;
        RECT 16.800 2.700 18.600 9.600 ;
        RECT 29.400 2.700 31.200 9.600 ;
        RECT 35.400 2.700 37.200 9.600 ;
        RECT 55.800 2.700 57.600 9.600 ;
        RECT 76.800 2.700 78.600 9.600 ;
        RECT 86.550 2.700 88.350 6.600 ;
        RECT 95.250 2.700 97.050 9.600 ;
        RECT 101.850 2.700 103.650 9.600 ;
        RECT 112.050 2.700 113.850 9.600 ;
        RECT 131.400 2.700 133.200 9.600 ;
        RECT 149.700 2.700 151.500 15.600 ;
        RECT 157.800 2.700 159.600 9.600 ;
        RECT 173.400 2.700 175.200 9.600 ;
        RECT 179.400 2.700 181.200 9.600 ;
        RECT 188.550 2.700 190.350 6.600 ;
        RECT 197.250 2.700 199.050 9.600 ;
        RECT 203.850 2.700 205.650 9.600 ;
        RECT 214.050 2.700 215.850 9.600 ;
        RECT 232.800 2.700 234.600 9.600 ;
        RECT 238.800 2.700 240.600 9.600 ;
        RECT 253.800 2.700 255.600 9.600 ;
        RECT 259.800 2.700 261.600 9.600 ;
        RECT 275.400 2.700 277.200 9.600 ;
        RECT 283.500 2.700 285.300 15.600 ;
        RECT 291.150 2.700 292.950 9.600 ;
        RECT 301.350 2.700 303.150 9.600 ;
        RECT 307.950 2.700 309.750 9.600 ;
        RECT 316.650 2.700 318.450 6.600 ;
        RECT 332.400 2.700 334.200 9.600 ;
        RECT 355.800 2.700 357.600 9.600 ;
        RECT 362.550 2.700 364.350 6.600 ;
        RECT 371.250 2.700 373.050 9.600 ;
        RECT 377.850 2.700 379.650 9.600 ;
        RECT 388.050 2.700 389.850 9.600 ;
        RECT 404.700 2.700 406.500 15.600 ;
        RECT 412.800 2.700 414.600 9.600 ;
        RECT 428.400 2.700 430.200 9.600 ;
        RECT 434.400 2.700 436.200 9.600 ;
        RECT 449.400 2.700 451.200 9.600 ;
        RECT 455.400 2.700 457.200 9.600 ;
        RECT 464.550 2.700 466.350 6.600 ;
        RECT 473.250 2.700 475.050 9.600 ;
        RECT 479.850 2.700 481.650 9.600 ;
        RECT 490.050 2.700 491.850 9.600 ;
        RECT 506.400 2.700 508.200 9.600 ;
        RECT 524.700 2.700 526.500 15.600 ;
        RECT 532.800 2.700 534.600 9.600 ;
        RECT 550.800 2.700 552.600 9.600 ;
        RECT 556.800 2.700 558.600 9.600 ;
        RECT 564.150 2.700 565.950 9.600 ;
        RECT 574.350 2.700 576.150 9.600 ;
        RECT 580.950 2.700 582.750 9.600 ;
        RECT 589.650 2.700 591.450 6.600 ;
        RECT 607.800 2.700 609.600 9.600 ;
        RECT 613.800 2.700 615.600 9.600 ;
        RECT 626.700 2.700 628.500 15.600 ;
        RECT 634.800 2.700 636.600 9.600 ;
        RECT 644.550 2.700 646.350 6.600 ;
        RECT 653.250 2.700 655.050 9.600 ;
        RECT 659.850 2.700 661.650 9.600 ;
        RECT 670.050 2.700 671.850 9.600 ;
        RECT 688.800 2.700 690.600 9.600 ;
        RECT 694.800 2.700 696.600 9.600 ;
        RECT 710.400 2.700 712.200 9.600 ;
        RECT 718.500 2.700 720.300 15.600 ;
        RECT 731.400 2.700 733.200 9.600 ;
        RECT 737.400 2.700 739.200 9.600 ;
        RECT 759.300 2.700 761.100 15.600 ;
        RECT 781.800 2.700 783.600 9.600 ;
        RECT 787.800 2.700 789.600 9.600 ;
        RECT 800.700 2.700 802.500 15.600 ;
        RECT 808.800 2.700 810.600 9.600 ;
        RECT 824.400 2.700 826.200 9.600 ;
        RECT 845.400 2.700 847.200 13.800 ;
        RECT 869.400 2.700 871.200 9.600 ;
        RECT 877.500 2.700 879.300 15.600 ;
        RECT -9.450 0.300 896.400 2.700 ;
    END
  END vdd
  PIN Cin[5]
    PORT
      LAYER metal1 ;
        RECT 706.950 876.450 709.050 877.050 ;
        RECT 718.950 876.450 721.050 877.050 ;
        RECT 706.950 875.550 721.050 876.450 ;
        RECT 706.950 874.950 709.050 875.550 ;
        RECT 718.950 874.950 721.050 875.550 ;
        RECT 604.950 762.450 609.000 763.050 ;
        RECT 604.950 760.950 609.450 762.450 ;
        RECT 608.550 757.050 609.450 760.950 ;
        RECT 604.950 755.550 609.450 757.050 ;
        RECT 604.950 754.950 609.000 755.550 ;
        RECT 580.950 567.450 583.050 568.050 ;
        RECT 586.950 567.450 589.050 568.050 ;
        RECT 580.950 566.550 589.050 567.450 ;
        RECT 580.950 565.950 583.050 566.550 ;
        RECT 586.950 565.950 589.050 566.550 ;
      LAYER metal2 ;
        RECT 731.400 898.050 732.600 906.600 ;
        RECT 718.950 895.950 721.050 898.050 ;
        RECT 730.950 895.950 733.050 898.050 ;
        RECT 719.400 877.050 720.600 895.950 ;
        RECT 706.950 874.950 709.050 877.050 ;
        RECT 718.950 874.950 721.050 877.050 ;
        RECT 707.400 859.050 708.600 874.950 ;
        RECT 619.950 856.950 622.050 859.050 ;
        RECT 706.950 856.950 709.050 859.050 ;
        RECT 620.400 793.050 621.600 856.950 ;
        RECT 604.950 790.950 607.050 793.050 ;
        RECT 619.800 790.950 621.900 793.050 ;
        RECT 605.400 763.050 606.600 790.950 ;
        RECT 603.000 762.600 607.050 763.050 ;
        RECT 602.400 760.950 607.050 762.600 ;
        RECT 602.400 760.050 603.600 760.950 ;
        RECT 601.950 757.950 604.050 760.050 ;
        RECT 604.950 754.950 607.050 757.050 ;
        RECT 605.400 745.050 606.600 754.950 ;
        RECT 577.950 742.950 580.050 745.050 ;
        RECT 604.950 742.950 607.050 745.050 ;
        RECT 565.950 724.950 568.050 727.050 ;
        RECT 566.400 723.900 567.600 724.950 ;
        RECT 578.400 724.050 579.600 742.950 ;
        RECT 565.950 721.800 568.050 723.900 ;
        RECT 577.950 721.950 580.050 724.050 ;
        RECT 601.950 721.800 604.050 723.900 ;
        RECT 602.400 706.050 603.600 721.800 ;
        RECT 601.950 703.950 604.050 706.050 ;
        RECT 613.950 703.950 616.050 706.050 ;
        RECT 614.400 625.050 615.600 703.950 ;
        RECT 583.950 622.950 586.050 625.050 ;
        RECT 613.950 622.950 616.050 625.050 ;
        RECT 584.400 600.600 585.600 622.950 ;
        RECT 581.400 599.400 585.600 600.600 ;
        RECT 581.400 568.050 582.600 599.400 ;
        RECT 628.950 568.950 631.050 571.050 ;
        RECT 580.950 565.950 583.050 568.050 ;
        RECT 586.950 565.950 589.050 568.050 ;
        RECT 587.400 541.050 588.600 565.950 ;
        RECT 629.400 541.050 630.600 568.950 ;
        RECT 586.950 538.950 589.050 541.050 ;
        RECT 628.950 538.950 631.050 541.050 ;
        RECT 587.400 502.050 588.600 538.950 ;
        RECT 565.950 499.950 568.050 502.050 ;
        RECT 586.950 499.950 589.050 502.050 ;
        RECT 566.400 460.050 567.600 499.950 ;
        RECT 565.950 457.950 568.050 460.050 ;
        RECT 577.950 457.950 580.050 460.050 ;
        RECT 578.400 448.050 579.600 457.950 ;
        RECT 577.950 445.950 580.050 448.050 ;
      LAYER metal3 ;
        RECT 718.950 897.600 721.050 898.050 ;
        RECT 730.950 897.600 733.050 898.050 ;
        RECT 718.950 896.400 733.050 897.600 ;
        RECT 718.950 895.950 721.050 896.400 ;
        RECT 730.950 895.950 733.050 896.400 ;
        RECT 619.950 858.600 622.050 859.050 ;
        RECT 706.950 858.600 709.050 859.050 ;
        RECT 619.950 857.400 709.050 858.600 ;
        RECT 619.950 856.950 622.050 857.400 ;
        RECT 706.950 856.950 709.050 857.400 ;
        RECT 604.950 792.600 607.050 793.050 ;
        RECT 619.800 792.600 621.900 793.050 ;
        RECT 604.950 791.400 621.900 792.600 ;
        RECT 604.950 790.950 607.050 791.400 ;
        RECT 619.800 790.950 621.900 791.400 ;
        RECT 577.950 744.600 580.050 745.050 ;
        RECT 604.950 744.600 607.050 745.050 ;
        RECT 577.950 743.400 607.050 744.600 ;
        RECT 577.950 742.950 580.050 743.400 ;
        RECT 604.950 742.950 607.050 743.400 ;
        RECT 565.950 723.450 568.050 723.900 ;
        RECT 577.950 723.450 580.050 724.050 ;
        RECT 601.950 723.450 604.050 723.900 ;
        RECT 565.950 722.250 604.050 723.450 ;
        RECT 565.950 721.800 568.050 722.250 ;
        RECT 577.950 721.950 580.050 722.250 ;
        RECT 601.950 721.800 604.050 722.250 ;
        RECT 601.950 705.600 604.050 706.050 ;
        RECT 613.950 705.600 616.050 706.050 ;
        RECT 601.950 704.400 616.050 705.600 ;
        RECT 601.950 703.950 604.050 704.400 ;
        RECT 613.950 703.950 616.050 704.400 ;
        RECT 583.950 624.600 586.050 625.050 ;
        RECT 613.950 624.600 616.050 625.050 ;
        RECT 583.950 623.400 616.050 624.600 ;
        RECT 583.950 622.950 586.050 623.400 ;
        RECT 613.950 622.950 616.050 623.400 ;
        RECT 586.950 540.600 589.050 541.050 ;
        RECT 628.950 540.600 631.050 541.050 ;
        RECT 586.950 539.400 631.050 540.600 ;
        RECT 586.950 538.950 589.050 539.400 ;
        RECT 628.950 538.950 631.050 539.400 ;
        RECT 565.950 501.600 568.050 502.050 ;
        RECT 586.950 501.600 589.050 502.050 ;
        RECT 565.950 500.400 589.050 501.600 ;
        RECT 565.950 499.950 568.050 500.400 ;
        RECT 586.950 499.950 589.050 500.400 ;
        RECT 565.950 459.600 568.050 460.050 ;
        RECT 577.950 459.600 580.050 460.050 ;
        RECT 565.950 458.400 580.050 459.600 ;
        RECT 565.950 457.950 568.050 458.400 ;
        RECT 577.950 457.950 580.050 458.400 ;
    END
  END Cin[5]
  PIN Cin[4]
    PORT
      LAYER metal1 ;
        RECT 652.950 607.950 655.050 610.050 ;
        RECT 653.550 601.050 654.450 607.950 ;
        RECT 649.950 599.550 654.450 601.050 ;
        RECT 649.950 598.950 654.000 599.550 ;
      LAYER metal2 ;
        RECT 725.400 892.050 726.600 906.600 ;
        RECT 691.950 889.950 694.050 892.050 ;
        RECT 724.950 889.950 727.050 892.050 ;
        RECT 692.400 853.050 693.600 889.950 ;
        RECT 646.950 850.950 649.050 853.050 ;
        RECT 691.800 850.950 693.900 853.050 ;
        RECT 647.400 778.050 648.600 850.950 ;
        RECT 634.950 775.950 637.050 778.050 ;
        RECT 646.950 775.950 649.050 778.050 ;
        RECT 586.950 733.950 589.050 736.050 ;
        RECT 595.950 733.950 598.050 736.050 ;
        RECT 587.400 727.050 588.600 733.950 ;
        RECT 596.400 730.050 597.600 733.950 ;
        RECT 635.400 730.200 636.600 775.950 ;
        RECT 595.950 727.950 598.050 730.050 ;
        RECT 634.950 728.100 637.050 730.200 ;
        RECT 664.950 728.100 667.050 730.200 ;
        RECT 635.400 727.050 636.600 728.100 ;
        RECT 544.950 724.950 547.050 727.050 ;
        RECT 586.950 724.950 589.050 727.050 ;
        RECT 634.950 724.950 637.050 727.050 ;
        RECT 545.400 723.900 546.600 724.950 ;
        RECT 544.950 721.800 547.050 723.900 ;
        RECT 556.950 721.950 559.050 724.050 ;
        RECT 557.400 682.050 558.600 721.950 ;
        RECT 665.400 699.600 666.600 728.100 ;
        RECT 662.400 698.400 666.600 699.600 ;
        RECT 556.950 679.950 559.050 682.050 ;
        RECT 662.400 670.050 663.600 698.400 ;
        RECT 640.950 667.950 643.050 670.050 ;
        RECT 661.950 667.950 664.050 670.050 ;
        RECT 641.400 631.050 642.600 667.950 ;
        RECT 640.950 628.950 643.050 631.050 ;
        RECT 652.950 628.950 655.050 631.050 ;
        RECT 653.400 610.050 654.600 628.950 ;
        RECT 652.950 607.950 655.050 610.050 ;
        RECT 649.950 598.950 652.050 601.050 ;
        RECT 650.400 574.050 651.600 598.950 ;
        RECT 649.950 571.950 652.050 574.050 ;
        RECT 649.950 565.950 652.050 568.050 ;
        RECT 595.950 523.950 598.050 526.050 ;
        RECT 596.400 511.050 597.600 523.950 ;
        RECT 650.400 514.050 651.600 565.950 ;
        RECT 649.950 511.950 652.050 514.050 ;
        RECT 595.950 508.950 598.050 511.050 ;
        RECT 625.950 508.950 628.050 511.050 ;
        RECT 626.400 496.050 627.600 508.950 ;
        RECT 625.950 493.950 628.050 496.050 ;
        RECT 625.950 487.950 628.050 490.050 ;
        RECT 626.400 466.050 627.600 487.950 ;
        RECT 598.950 463.950 601.050 466.050 ;
        RECT 625.950 463.950 628.050 466.050 ;
        RECT 646.950 463.950 649.050 466.050 ;
        RECT 511.950 449.100 514.050 451.200 ;
        RECT 532.950 449.100 535.050 451.200 ;
        RECT 595.950 450.600 598.050 451.050 ;
        RECT 599.400 450.600 600.600 463.950 ;
        RECT 595.950 449.400 600.600 450.600 ;
        RECT 512.400 448.050 513.600 449.100 ;
        RECT 533.400 448.050 534.600 449.100 ;
        RECT 595.950 448.950 598.050 449.400 ;
        RECT 596.400 448.050 597.600 448.950 ;
        RECT 511.950 445.950 514.050 448.050 ;
        RECT 532.950 445.950 535.050 448.050 ;
        RECT 595.950 445.950 598.050 448.050 ;
        RECT 647.400 442.050 648.600 463.950 ;
        RECT 667.950 445.950 670.050 448.050 ;
        RECT 668.400 444.000 669.600 445.950 ;
        RECT 646.950 439.950 649.050 442.050 ;
        RECT 667.950 441.600 670.050 444.000 ;
        RECT 665.400 440.400 670.050 441.600 ;
        RECT 665.400 421.050 666.600 440.400 ;
        RECT 667.950 439.950 670.050 440.400 ;
        RECT 664.950 418.950 667.050 421.050 ;
        RECT 727.800 420.000 729.900 421.050 ;
        RECT 727.800 418.950 730.050 420.000 ;
        RECT 655.950 412.950 658.050 415.050 ;
        RECT 656.400 411.900 657.600 412.950 ;
        RECT 665.400 411.900 666.600 418.950 ;
        RECT 727.950 417.000 730.050 418.950 ;
        RECT 728.400 415.050 729.600 417.000 ;
        RECT 727.950 412.950 730.050 415.050 ;
        RECT 655.950 409.800 658.050 411.900 ;
        RECT 664.950 409.800 667.050 411.900 ;
      LAYER metal3 ;
        RECT 691.950 891.600 694.050 892.050 ;
        RECT 724.950 891.600 727.050 892.050 ;
        RECT 691.950 890.400 727.050 891.600 ;
        RECT 691.950 889.950 694.050 890.400 ;
        RECT 724.950 889.950 727.050 890.400 ;
        RECT 646.950 852.600 649.050 853.050 ;
        RECT 691.800 852.600 693.900 853.050 ;
        RECT 646.950 851.400 693.900 852.600 ;
        RECT 646.950 850.950 649.050 851.400 ;
        RECT 691.800 850.950 693.900 851.400 ;
        RECT 634.950 777.600 637.050 778.050 ;
        RECT 646.950 777.600 649.050 778.050 ;
        RECT 634.950 776.400 649.050 777.600 ;
        RECT 634.950 775.950 637.050 776.400 ;
        RECT 646.950 775.950 649.050 776.400 ;
        RECT 586.950 735.600 589.050 736.050 ;
        RECT 595.950 735.600 598.050 736.050 ;
        RECT 586.950 734.400 598.050 735.600 ;
        RECT 586.950 733.950 589.050 734.400 ;
        RECT 595.950 733.950 598.050 734.400 ;
        RECT 595.950 729.600 598.050 730.050 ;
        RECT 634.950 729.750 637.050 730.200 ;
        RECT 664.950 729.750 667.050 730.200 ;
        RECT 634.950 729.600 667.050 729.750 ;
        RECT 593.400 728.550 667.050 729.600 ;
        RECT 593.400 728.400 637.050 728.550 ;
        RECT 593.400 726.600 594.600 728.400 ;
        RECT 595.950 727.950 598.050 728.400 ;
        RECT 634.950 728.100 637.050 728.400 ;
        RECT 664.950 728.100 667.050 728.550 ;
        RECT 551.400 725.400 594.600 726.600 ;
        RECT 544.950 723.600 547.050 723.900 ;
        RECT 551.400 723.600 552.600 725.400 ;
        RECT 556.950 723.600 559.050 724.050 ;
        RECT 544.950 722.400 559.050 723.600 ;
        RECT 544.950 721.800 547.050 722.400 ;
        RECT 556.950 721.950 559.050 722.400 ;
        RECT 640.950 669.600 643.050 670.050 ;
        RECT 661.950 669.600 664.050 670.050 ;
        RECT 640.950 668.400 664.050 669.600 ;
        RECT 640.950 667.950 643.050 668.400 ;
        RECT 661.950 667.950 664.050 668.400 ;
        RECT 640.950 630.600 643.050 631.050 ;
        RECT 652.950 630.600 655.050 631.050 ;
        RECT 640.950 629.400 655.050 630.600 ;
        RECT 640.950 628.950 643.050 629.400 ;
        RECT 652.950 628.950 655.050 629.400 ;
        RECT 649.950 571.950 652.050 574.050 ;
        RECT 650.400 568.050 651.600 571.950 ;
        RECT 649.950 565.950 652.050 568.050 ;
        RECT 649.950 513.600 652.050 514.050 ;
        RECT 626.400 512.400 652.050 513.600 ;
        RECT 626.400 511.050 627.600 512.400 ;
        RECT 649.950 511.950 652.050 512.400 ;
        RECT 595.950 510.600 598.050 511.050 ;
        RECT 625.950 510.600 628.050 511.050 ;
        RECT 595.950 509.400 628.050 510.600 ;
        RECT 595.950 508.950 598.050 509.400 ;
        RECT 625.950 508.950 628.050 509.400 ;
        RECT 625.950 493.950 628.050 496.050 ;
        RECT 626.400 490.050 627.600 493.950 ;
        RECT 625.950 487.950 628.050 490.050 ;
        RECT 598.950 465.600 601.050 466.050 ;
        RECT 625.950 465.600 628.050 466.050 ;
        RECT 646.950 465.600 649.050 466.050 ;
        RECT 598.950 464.400 649.050 465.600 ;
        RECT 598.950 463.950 601.050 464.400 ;
        RECT 625.950 463.950 628.050 464.400 ;
        RECT 646.950 463.950 649.050 464.400 ;
        RECT 511.950 450.600 514.050 451.200 ;
        RECT 532.950 450.600 535.050 451.200 ;
        RECT 595.950 450.600 598.050 451.050 ;
        RECT 511.950 449.400 535.050 450.600 ;
        RECT 511.950 449.100 514.050 449.400 ;
        RECT 532.950 449.100 535.050 449.400 ;
        RECT 593.400 449.400 598.050 450.600 ;
        RECT 533.400 447.600 534.600 449.100 ;
        RECT 593.400 447.600 594.600 449.400 ;
        RECT 595.950 448.950 598.050 449.400 ;
        RECT 533.400 446.400 594.600 447.600 ;
        RECT 646.950 441.600 649.050 442.050 ;
        RECT 667.950 441.600 670.050 442.050 ;
        RECT 646.950 440.400 670.050 441.600 ;
        RECT 646.950 439.950 649.050 440.400 ;
        RECT 667.950 439.950 670.050 440.400 ;
        RECT 664.950 420.600 667.050 421.050 ;
        RECT 727.800 420.600 729.900 421.050 ;
        RECT 664.950 419.400 729.900 420.600 ;
        RECT 664.950 418.950 667.050 419.400 ;
        RECT 727.800 418.950 729.900 419.400 ;
        RECT 655.950 411.450 658.050 411.900 ;
        RECT 664.950 411.450 667.050 411.900 ;
        RECT 655.950 410.250 667.050 411.450 ;
        RECT 655.950 409.800 658.050 410.250 ;
        RECT 664.950 409.800 667.050 410.250 ;
    END
  END Cin[4]
  PIN Cin[3]
    PORT
      LAYER metal1 ;
        RECT 573.000 651.450 577.050 652.050 ;
        RECT 572.550 649.950 577.050 651.450 ;
        RECT 572.550 646.050 573.450 649.950 ;
        RECT 572.550 644.550 577.050 646.050 ;
        RECT 573.000 643.950 577.050 644.550 ;
      LAYER metal2 ;
        RECT 707.400 905.400 711.600 906.600 ;
        RECT 694.950 895.950 697.050 898.050 ;
        RECT 700.950 897.600 703.050 898.050 ;
        RECT 707.400 897.600 708.600 905.400 ;
        RECT 700.950 896.400 708.600 897.600 ;
        RECT 700.950 895.950 703.050 896.400 ;
        RECT 695.400 853.050 696.600 895.950 ;
        RECT 694.950 850.950 697.050 853.050 ;
        RECT 706.950 850.950 709.050 853.050 ;
        RECT 707.400 835.050 708.600 850.950 ;
        RECT 700.950 832.950 703.050 835.050 ;
        RECT 706.950 832.950 709.050 835.050 ;
        RECT 701.400 817.050 702.600 832.950 ;
        RECT 691.950 814.950 694.050 817.050 ;
        RECT 700.950 814.950 703.050 817.050 ;
        RECT 692.400 739.050 693.600 814.950 ;
        RECT 667.950 736.950 670.050 739.050 ;
        RECT 691.950 736.950 694.050 739.050 ;
        RECT 523.950 724.950 526.050 727.050 ;
        RECT 524.400 685.050 525.600 724.950 ;
        RECT 668.400 718.050 669.600 736.950 ;
        RECT 637.950 715.950 640.050 718.050 ;
        RECT 667.950 715.950 670.050 718.050 ;
        RECT 523.950 682.950 526.050 685.050 ;
        RECT 508.950 679.950 511.050 682.050 ;
        RECT 625.950 679.950 628.050 682.050 ;
        RECT 509.400 678.600 510.600 679.950 ;
        RECT 511.950 678.600 514.050 679.050 ;
        RECT 509.400 677.400 514.050 678.600 ;
        RECT 626.400 678.000 627.600 679.950 ;
        RECT 511.950 676.950 514.050 677.400 ;
        RECT 512.400 673.050 513.600 676.950 ;
        RECT 604.950 673.950 607.050 676.050 ;
        RECT 625.950 673.950 628.050 678.000 ;
        RECT 638.400 676.050 639.600 715.950 ;
        RECT 637.950 673.950 640.050 676.050 ;
        RECT 511.950 670.950 514.050 673.050 ;
        RECT 532.950 670.950 535.050 673.050 ;
        RECT 523.950 646.950 526.050 649.050 ;
        RECT 524.400 645.900 525.600 646.950 ;
        RECT 533.400 646.050 534.600 670.950 ;
        RECT 605.400 658.050 606.600 673.950 ;
        RECT 574.950 655.950 577.050 658.050 ;
        RECT 604.950 655.950 607.050 658.050 ;
        RECT 575.400 652.050 576.600 655.950 ;
        RECT 574.950 649.950 577.050 652.050 ;
        RECT 538.950 646.950 541.050 649.050 ;
        RECT 523.950 643.800 526.050 645.900 ;
        RECT 532.950 643.950 535.050 646.050 ;
        RECT 539.400 645.900 540.600 646.950 ;
        RECT 538.950 643.800 541.050 645.900 ;
        RECT 574.950 643.950 577.050 646.050 ;
        RECT 524.400 553.050 525.600 643.800 ;
        RECT 539.400 631.050 540.600 643.800 ;
        RECT 575.400 631.050 576.600 643.950 ;
        RECT 538.950 628.950 541.050 631.050 ;
        RECT 574.950 628.950 577.050 631.050 ;
        RECT 523.950 550.950 526.050 553.050 ;
        RECT 541.950 550.950 544.050 553.050 ;
        RECT 542.400 484.050 543.600 550.950 ;
        RECT 571.950 490.950 574.050 493.050 ;
        RECT 572.400 484.050 573.600 490.950 ;
        RECT 541.950 481.950 544.050 484.050 ;
        RECT 571.950 481.950 574.050 484.050 ;
        RECT 572.400 469.050 573.600 481.950 ;
        RECT 571.950 466.950 574.050 469.050 ;
        RECT 583.950 466.950 586.050 469.050 ;
        RECT 584.400 436.050 585.600 466.950 ;
        RECT 637.950 445.950 640.050 448.050 ;
        RECT 661.950 445.950 664.050 448.050 ;
        RECT 638.400 444.900 639.600 445.950 ;
        RECT 637.950 442.800 640.050 444.900 ;
        RECT 643.950 442.950 646.050 445.050 ;
        RECT 662.400 444.900 663.600 445.950 ;
        RECT 644.400 436.050 645.600 442.950 ;
        RECT 661.950 442.800 664.050 444.900 ;
        RECT 583.950 433.950 586.050 436.050 ;
        RECT 643.950 433.950 646.050 436.050 ;
        RECT 613.950 412.950 616.050 415.050 ;
        RECT 614.400 411.900 615.600 412.950 ;
        RECT 644.400 411.900 645.600 433.950 ;
        RECT 613.950 409.800 616.050 411.900 ;
        RECT 643.950 411.600 646.050 411.900 ;
        RECT 643.950 410.400 648.600 411.600 ;
        RECT 643.950 409.800 646.050 410.400 ;
        RECT 647.400 376.050 648.600 410.400 ;
        RECT 646.950 373.950 649.050 376.050 ;
        RECT 670.950 372.000 673.050 376.050 ;
        RECT 671.400 370.050 672.600 372.000 ;
        RECT 670.950 367.950 673.050 370.050 ;
      LAYER metal3 ;
        RECT 694.950 897.600 697.050 898.050 ;
        RECT 700.950 897.600 703.050 898.050 ;
        RECT 694.950 896.400 703.050 897.600 ;
        RECT 694.950 895.950 697.050 896.400 ;
        RECT 700.950 895.950 703.050 896.400 ;
        RECT 694.950 852.600 697.050 853.050 ;
        RECT 706.950 852.600 709.050 853.050 ;
        RECT 694.950 851.400 709.050 852.600 ;
        RECT 694.950 850.950 697.050 851.400 ;
        RECT 706.950 850.950 709.050 851.400 ;
        RECT 700.950 834.600 703.050 835.050 ;
        RECT 706.950 834.600 709.050 835.050 ;
        RECT 700.950 833.400 709.050 834.600 ;
        RECT 700.950 832.950 703.050 833.400 ;
        RECT 706.950 832.950 709.050 833.400 ;
        RECT 691.950 816.600 694.050 817.050 ;
        RECT 700.950 816.600 703.050 817.050 ;
        RECT 691.950 815.400 703.050 816.600 ;
        RECT 691.950 814.950 694.050 815.400 ;
        RECT 700.950 814.950 703.050 815.400 ;
        RECT 667.950 738.600 670.050 739.050 ;
        RECT 691.950 738.600 694.050 739.050 ;
        RECT 667.950 737.400 694.050 738.600 ;
        RECT 667.950 736.950 670.050 737.400 ;
        RECT 691.950 736.950 694.050 737.400 ;
        RECT 637.950 717.600 640.050 718.050 ;
        RECT 667.950 717.600 670.050 718.050 ;
        RECT 637.950 716.400 670.050 717.600 ;
        RECT 637.950 715.950 640.050 716.400 ;
        RECT 667.950 715.950 670.050 716.400 ;
        RECT 523.950 682.950 526.050 685.050 ;
        RECT 511.950 678.600 514.050 679.050 ;
        RECT 524.400 678.600 525.600 682.950 ;
        RECT 511.950 677.400 525.600 678.600 ;
        RECT 511.950 676.950 514.050 677.400 ;
        RECT 604.950 675.600 607.050 676.050 ;
        RECT 625.950 675.600 628.050 676.050 ;
        RECT 637.950 675.600 640.050 676.050 ;
        RECT 604.950 674.400 640.050 675.600 ;
        RECT 604.950 673.950 607.050 674.400 ;
        RECT 625.950 673.950 628.050 674.400 ;
        RECT 637.950 673.950 640.050 674.400 ;
        RECT 511.950 672.600 514.050 673.050 ;
        RECT 532.950 672.600 535.050 673.050 ;
        RECT 511.950 671.400 535.050 672.600 ;
        RECT 511.950 670.950 514.050 671.400 ;
        RECT 532.950 670.950 535.050 671.400 ;
        RECT 574.950 657.600 577.050 658.050 ;
        RECT 604.950 657.600 607.050 658.050 ;
        RECT 574.950 656.400 607.050 657.600 ;
        RECT 574.950 655.950 577.050 656.400 ;
        RECT 604.950 655.950 607.050 656.400 ;
        RECT 523.950 645.600 526.050 645.900 ;
        RECT 532.950 645.600 535.050 646.050 ;
        RECT 538.950 645.600 541.050 645.900 ;
        RECT 523.950 644.400 541.050 645.600 ;
        RECT 523.950 643.800 526.050 644.400 ;
        RECT 532.950 643.950 535.050 644.400 ;
        RECT 538.950 643.800 541.050 644.400 ;
        RECT 538.950 630.600 541.050 631.050 ;
        RECT 574.950 630.600 577.050 631.050 ;
        RECT 538.950 629.400 577.050 630.600 ;
        RECT 538.950 628.950 541.050 629.400 ;
        RECT 574.950 628.950 577.050 629.400 ;
        RECT 523.950 552.600 526.050 553.050 ;
        RECT 541.950 552.600 544.050 553.050 ;
        RECT 523.950 551.400 544.050 552.600 ;
        RECT 523.950 550.950 526.050 551.400 ;
        RECT 541.950 550.950 544.050 551.400 ;
        RECT 541.950 483.600 544.050 484.050 ;
        RECT 571.950 483.600 574.050 484.050 ;
        RECT 541.950 482.400 574.050 483.600 ;
        RECT 541.950 481.950 544.050 482.400 ;
        RECT 571.950 481.950 574.050 482.400 ;
        RECT 571.950 468.600 574.050 469.050 ;
        RECT 583.950 468.600 586.050 469.050 ;
        RECT 571.950 467.400 586.050 468.600 ;
        RECT 571.950 466.950 574.050 467.400 ;
        RECT 583.950 466.950 586.050 467.400 ;
        RECT 637.950 444.600 640.050 444.900 ;
        RECT 643.950 444.600 646.050 445.050 ;
        RECT 661.950 444.600 664.050 444.900 ;
        RECT 637.950 443.400 664.050 444.600 ;
        RECT 637.950 442.800 640.050 443.400 ;
        RECT 643.950 442.950 646.050 443.400 ;
        RECT 661.950 442.800 664.050 443.400 ;
        RECT 583.950 435.600 586.050 436.050 ;
        RECT 643.950 435.600 646.050 436.050 ;
        RECT 583.950 434.400 646.050 435.600 ;
        RECT 583.950 433.950 586.050 434.400 ;
        RECT 643.950 433.950 646.050 434.400 ;
        RECT 613.950 411.450 616.050 411.900 ;
        RECT 643.950 411.450 646.050 411.900 ;
        RECT 613.950 410.250 646.050 411.450 ;
        RECT 613.950 409.800 616.050 410.250 ;
        RECT 643.950 409.800 646.050 410.250 ;
        RECT 646.950 375.600 649.050 376.050 ;
        RECT 670.950 375.600 673.050 376.050 ;
        RECT 646.950 374.400 673.050 375.600 ;
        RECT 646.950 373.950 649.050 374.400 ;
        RECT 670.950 373.950 673.050 374.400 ;
    END
  END Cin[3]
  PIN Cin[2]
    PORT
      LAYER metal1 ;
        RECT 331.950 765.450 334.050 766.050 ;
        RECT 340.950 765.450 343.050 766.050 ;
        RECT 331.950 764.550 343.050 765.450 ;
        RECT 331.950 763.950 334.050 764.550 ;
        RECT 340.950 763.950 343.050 764.550 ;
        RECT 415.950 765.450 418.050 766.050 ;
        RECT 433.950 765.450 436.050 766.050 ;
        RECT 415.950 764.550 436.050 765.450 ;
        RECT 415.950 763.950 418.050 764.550 ;
        RECT 433.950 763.950 436.050 764.550 ;
        RECT 757.950 762.450 762.000 763.050 ;
        RECT 757.950 760.950 762.450 762.450 ;
        RECT 761.550 756.450 762.450 760.950 ;
        RECT 769.950 756.450 772.050 757.050 ;
        RECT 761.550 755.550 772.050 756.450 ;
        RECT 769.950 754.950 772.050 755.550 ;
        RECT 730.950 630.450 733.050 631.050 ;
        RECT 736.950 630.450 739.050 631.050 ;
        RECT 730.950 629.550 739.050 630.450 ;
        RECT 730.950 628.950 733.050 629.550 ;
        RECT 736.950 628.950 739.050 629.550 ;
        RECT 768.000 528.450 772.050 529.050 ;
        RECT 767.550 526.950 772.050 528.450 ;
        RECT 767.550 525.450 768.450 526.950 ;
        RECT 764.550 524.550 768.450 525.450 ;
        RECT 757.950 522.450 760.050 523.050 ;
        RECT 764.550 522.450 765.450 524.550 ;
        RECT 757.950 521.550 765.450 522.450 ;
        RECT 757.950 520.950 760.050 521.550 ;
        RECT 733.950 453.450 736.050 454.050 ;
        RECT 751.950 453.450 754.050 454.050 ;
        RECT 733.950 452.550 754.050 453.450 ;
        RECT 733.950 451.950 736.050 452.550 ;
        RECT 751.950 451.950 754.050 452.550 ;
      LAYER metal2 ;
        RECT 704.400 901.050 705.600 906.600 ;
        RECT 703.950 898.950 706.050 901.050 ;
        RECT 715.950 898.950 718.050 901.050 ;
        RECT 716.400 862.050 717.600 898.950 ;
        RECT 709.950 859.950 712.050 862.050 ;
        RECT 715.950 859.950 718.050 862.050 ;
        RECT 710.400 829.050 711.600 859.950 ;
        RECT 688.950 826.950 691.050 829.050 ;
        RECT 709.950 826.950 712.050 829.050 ;
        RECT 715.950 826.950 718.050 829.050 ;
        RECT 689.400 820.050 690.600 826.950 ;
        RECT 616.950 817.950 619.050 820.050 ;
        RECT 688.950 817.950 691.050 820.050 ;
        RECT 617.400 796.050 618.600 817.950 ;
        RECT 553.950 793.950 556.050 796.050 ;
        RECT 616.950 793.950 619.050 796.050 ;
        RECT 340.950 781.950 343.050 784.050 ;
        RECT 415.950 781.950 418.050 784.050 ;
        RECT 433.950 781.950 436.050 784.050 ;
        RECT 466.950 781.950 469.050 784.050 ;
        RECT 341.400 766.050 342.600 781.950 ;
        RECT 416.400 766.050 417.600 781.950 ;
        RECT 434.400 766.050 435.600 781.950 ;
        RECT 467.400 775.050 468.600 781.950 ;
        RECT 554.400 775.050 555.600 793.950 ;
        RECT 716.400 793.050 717.600 826.950 ;
        RECT 715.950 790.950 718.050 793.050 ;
        RECT 757.950 790.950 760.050 793.050 ;
        RECT 466.950 772.950 469.050 775.050 ;
        RECT 553.950 772.950 556.050 775.050 ;
        RECT 331.950 762.000 334.050 766.050 ;
        RECT 340.950 765.600 343.050 766.050 ;
        RECT 338.400 764.400 343.050 765.600 ;
        RECT 332.400 760.050 333.600 762.000 ;
        RECT 331.950 757.950 334.050 760.050 ;
        RECT 338.400 709.050 339.600 764.400 ;
        RECT 340.950 763.950 343.050 764.400 ;
        RECT 415.950 762.000 418.050 766.050 ;
        RECT 433.950 763.950 436.050 766.050 ;
        RECT 758.400 763.050 759.600 790.950 ;
        RECT 416.400 760.050 417.600 762.000 ;
        RECT 757.950 760.950 760.050 763.050 ;
        RECT 415.950 757.950 418.050 760.050 ;
        RECT 769.950 754.950 772.050 757.050 ;
        RECT 770.400 748.050 771.600 754.950 ;
        RECT 769.950 745.950 772.050 748.050 ;
        RECT 778.950 745.950 781.050 748.050 ;
        RECT 751.950 724.950 754.050 727.050 ;
        RECT 752.400 721.050 753.600 724.950 ;
        RECT 779.400 721.050 780.600 745.950 ;
        RECT 751.950 718.950 754.050 721.050 ;
        RECT 778.950 718.950 781.050 721.050 ;
        RECT 289.950 706.950 292.050 709.050 ;
        RECT 337.950 706.950 340.050 709.050 ;
        RECT 290.400 682.050 291.600 706.950 ;
        RECT 752.400 699.600 753.600 718.950 ;
        RECT 752.400 698.400 756.600 699.600 ;
        RECT 289.950 679.950 292.050 682.050 ;
        RECT 755.400 658.050 756.600 698.400 ;
        RECT 715.950 655.950 718.050 658.050 ;
        RECT 736.950 655.950 739.050 658.050 ;
        RECT 754.950 655.950 757.050 658.050 ;
        RECT 716.400 649.050 717.600 655.950 ;
        RECT 715.950 646.950 718.050 649.050 ;
        RECT 737.400 631.050 738.600 655.950 ;
        RECT 730.950 628.950 733.050 631.050 ;
        RECT 736.950 628.950 739.050 631.050 ;
        RECT 731.400 607.200 732.600 628.950 ;
        RECT 730.950 605.100 733.050 607.200 ;
        RECT 731.400 604.050 732.600 605.100 ;
        RECT 763.800 604.950 765.900 607.050 ;
        RECT 730.950 601.950 733.050 604.050 ;
        RECT 764.400 586.050 765.600 604.950 ;
        RECT 763.950 583.950 766.050 586.050 ;
        RECT 778.950 583.950 781.050 586.050 ;
        RECT 779.400 556.050 780.600 583.950 ;
        RECT 769.950 553.950 772.050 556.050 ;
        RECT 778.950 553.950 781.050 556.050 ;
        RECT 770.400 529.050 771.600 553.950 ;
        RECT 769.950 526.950 772.050 529.050 ;
        RECT 757.950 520.950 760.050 523.050 ;
        RECT 758.400 499.050 759.600 520.950 ;
        RECT 751.950 496.950 754.050 499.050 ;
        RECT 757.950 496.950 760.050 499.050 ;
        RECT 685.950 454.950 688.050 457.050 ;
        RECT 686.400 448.050 687.600 454.950 ;
        RECT 733.950 450.000 736.050 457.050 ;
        RECT 752.400 454.050 753.600 496.950 ;
        RECT 751.950 451.950 754.050 454.050 ;
        RECT 734.400 448.050 735.600 450.000 ;
        RECT 752.400 448.050 753.600 451.950 ;
        RECT 685.950 445.950 688.050 448.050 ;
        RECT 733.950 445.950 736.050 448.050 ;
        RECT 751.950 445.950 754.050 448.050 ;
      LAYER metal3 ;
        RECT 703.950 900.600 706.050 901.050 ;
        RECT 715.950 900.600 718.050 901.050 ;
        RECT 703.950 899.400 718.050 900.600 ;
        RECT 703.950 898.950 706.050 899.400 ;
        RECT 715.950 898.950 718.050 899.400 ;
        RECT 709.950 861.600 712.050 862.050 ;
        RECT 715.950 861.600 718.050 862.050 ;
        RECT 709.950 860.400 718.050 861.600 ;
        RECT 709.950 859.950 712.050 860.400 ;
        RECT 715.950 859.950 718.050 860.400 ;
        RECT 688.950 828.600 691.050 829.050 ;
        RECT 709.950 828.600 712.050 829.050 ;
        RECT 715.950 828.600 718.050 829.050 ;
        RECT 688.950 827.400 718.050 828.600 ;
        RECT 688.950 826.950 691.050 827.400 ;
        RECT 709.950 826.950 712.050 827.400 ;
        RECT 715.950 826.950 718.050 827.400 ;
        RECT 616.950 819.600 619.050 820.050 ;
        RECT 688.950 819.600 691.050 820.050 ;
        RECT 616.950 818.400 691.050 819.600 ;
        RECT 616.950 817.950 619.050 818.400 ;
        RECT 688.950 817.950 691.050 818.400 ;
        RECT 553.950 795.600 556.050 796.050 ;
        RECT 616.950 795.600 619.050 796.050 ;
        RECT 553.950 794.400 619.050 795.600 ;
        RECT 553.950 793.950 556.050 794.400 ;
        RECT 616.950 793.950 619.050 794.400 ;
        RECT 715.950 792.600 718.050 793.050 ;
        RECT 757.950 792.600 760.050 793.050 ;
        RECT 715.950 791.400 760.050 792.600 ;
        RECT 715.950 790.950 718.050 791.400 ;
        RECT 757.950 790.950 760.050 791.400 ;
        RECT 340.950 783.600 343.050 784.050 ;
        RECT 415.950 783.600 418.050 784.050 ;
        RECT 340.950 782.400 418.050 783.600 ;
        RECT 340.950 781.950 343.050 782.400 ;
        RECT 415.950 781.950 418.050 782.400 ;
        RECT 433.950 783.600 436.050 784.050 ;
        RECT 466.950 783.600 469.050 784.050 ;
        RECT 433.950 782.400 469.050 783.600 ;
        RECT 433.950 781.950 436.050 782.400 ;
        RECT 466.950 781.950 469.050 782.400 ;
        RECT 466.950 774.600 469.050 775.050 ;
        RECT 553.950 774.600 556.050 775.050 ;
        RECT 466.950 773.400 556.050 774.600 ;
        RECT 466.950 772.950 469.050 773.400 ;
        RECT 553.950 772.950 556.050 773.400 ;
        RECT 769.950 747.600 772.050 748.050 ;
        RECT 778.950 747.600 781.050 748.050 ;
        RECT 769.950 746.400 781.050 747.600 ;
        RECT 769.950 745.950 772.050 746.400 ;
        RECT 778.950 745.950 781.050 746.400 ;
        RECT 751.950 720.600 754.050 721.050 ;
        RECT 778.950 720.600 781.050 721.050 ;
        RECT 751.950 719.400 781.050 720.600 ;
        RECT 751.950 718.950 754.050 719.400 ;
        RECT 778.950 718.950 781.050 719.400 ;
        RECT 289.950 708.600 292.050 709.050 ;
        RECT 337.950 708.600 340.050 709.050 ;
        RECT 289.950 707.400 340.050 708.600 ;
        RECT 289.950 706.950 292.050 707.400 ;
        RECT 337.950 706.950 340.050 707.400 ;
        RECT 715.950 657.600 718.050 658.050 ;
        RECT 736.950 657.600 739.050 658.050 ;
        RECT 754.950 657.600 757.050 658.050 ;
        RECT 715.950 656.400 757.050 657.600 ;
        RECT 715.950 655.950 718.050 656.400 ;
        RECT 736.950 655.950 739.050 656.400 ;
        RECT 754.950 655.950 757.050 656.400 ;
        RECT 730.950 606.600 733.050 607.200 ;
        RECT 763.800 606.600 765.900 607.050 ;
        RECT 730.950 605.400 765.900 606.600 ;
        RECT 730.950 605.100 733.050 605.400 ;
        RECT 763.800 604.950 765.900 605.400 ;
        RECT 763.950 585.600 766.050 586.050 ;
        RECT 778.950 585.600 781.050 586.050 ;
        RECT 763.950 584.400 781.050 585.600 ;
        RECT 763.950 583.950 766.050 584.400 ;
        RECT 778.950 583.950 781.050 584.400 ;
        RECT 769.950 555.600 772.050 556.050 ;
        RECT 778.950 555.600 781.050 556.050 ;
        RECT 769.950 554.400 781.050 555.600 ;
        RECT 769.950 553.950 772.050 554.400 ;
        RECT 778.950 553.950 781.050 554.400 ;
        RECT 751.950 498.600 754.050 499.050 ;
        RECT 757.950 498.600 760.050 499.050 ;
        RECT 751.950 497.400 760.050 498.600 ;
        RECT 751.950 496.950 754.050 497.400 ;
        RECT 757.950 496.950 760.050 497.400 ;
        RECT 685.950 456.600 688.050 457.050 ;
        RECT 733.950 456.600 736.050 457.050 ;
        RECT 685.950 455.400 736.050 456.600 ;
        RECT 685.950 454.950 688.050 455.400 ;
        RECT 733.950 454.950 736.050 455.400 ;
    END
  END Cin[2]
  PIN Cin[1]
    PORT
      LAYER metal1 ;
        RECT 568.950 729.450 573.000 730.050 ;
        RECT 568.950 727.950 573.450 729.450 ;
        RECT 572.550 724.050 573.450 727.950 ;
        RECT 568.950 722.550 573.450 724.050 ;
        RECT 568.950 721.950 573.000 722.550 ;
        RECT 567.000 684.450 571.050 685.050 ;
        RECT 566.550 682.950 571.050 684.450 ;
        RECT 566.550 679.050 567.450 682.950 ;
        RECT 566.550 677.550 571.050 679.050 ;
        RECT 567.000 676.950 571.050 677.550 ;
      LAYER metal2 ;
        RECT 530.400 901.050 531.600 906.600 ;
        RECT 529.950 898.950 532.050 901.050 ;
        RECT 571.950 898.950 574.050 901.050 ;
        RECT 572.400 876.600 573.600 898.950 ;
        RECT 569.400 875.400 573.600 876.600 ;
        RECT 569.400 730.050 570.600 875.400 ;
        RECT 568.950 727.950 571.050 730.050 ;
        RECT 568.950 721.950 571.050 724.050 ;
        RECT 569.400 685.050 570.600 721.950 ;
        RECT 568.950 682.950 571.050 685.050 ;
        RECT 568.950 676.950 571.050 679.050 ;
        RECT 569.400 616.050 570.600 676.950 ;
        RECT 445.950 613.950 448.050 616.050 ;
        RECT 568.950 613.950 571.050 616.050 ;
        RECT 697.950 613.950 700.050 616.050 ;
        RECT 436.950 601.950 439.050 604.050 ;
        RECT 437.400 600.000 438.600 601.950 ;
        RECT 436.950 595.950 439.050 600.000 ;
        RECT 446.400 598.050 447.600 613.950 ;
        RECT 457.950 601.950 460.050 604.050 ;
        RECT 458.400 600.000 459.600 601.950 ;
        RECT 698.400 600.900 699.600 613.950 ;
        RECT 703.950 601.950 706.050 604.050 ;
        RECT 704.400 600.900 705.600 601.950 ;
        RECT 445.950 595.950 448.050 598.050 ;
        RECT 457.950 595.950 460.050 600.000 ;
        RECT 697.950 598.800 700.050 600.900 ;
        RECT 703.800 598.800 705.900 600.900 ;
        RECT 698.400 583.050 699.600 598.800 ;
        RECT 688.950 580.950 691.050 583.050 ;
        RECT 697.950 580.950 700.050 583.050 ;
        RECT 689.400 535.050 690.600 580.950 ;
        RECT 688.950 532.950 691.050 535.050 ;
        RECT 694.950 532.950 697.050 535.050 ;
        RECT 695.400 522.900 696.600 532.950 ;
        RECT 700.950 523.950 703.050 526.050 ;
        RECT 701.400 522.900 702.600 523.950 ;
        RECT 694.950 520.800 697.050 522.900 ;
        RECT 700.950 520.800 703.050 522.900 ;
      LAYER metal3 ;
        RECT 529.950 900.600 532.050 901.050 ;
        RECT 571.950 900.600 574.050 901.050 ;
        RECT 529.950 899.400 574.050 900.600 ;
        RECT 529.950 898.950 532.050 899.400 ;
        RECT 571.950 898.950 574.050 899.400 ;
        RECT 445.950 615.600 448.050 616.050 ;
        RECT 568.950 615.600 571.050 616.050 ;
        RECT 697.950 615.600 700.050 616.050 ;
        RECT 445.950 614.400 700.050 615.600 ;
        RECT 445.950 613.950 448.050 614.400 ;
        RECT 568.950 613.950 571.050 614.400 ;
        RECT 697.950 613.950 700.050 614.400 ;
        RECT 697.950 600.450 700.050 600.900 ;
        RECT 703.800 600.450 705.900 600.900 ;
        RECT 697.950 599.250 705.900 600.450 ;
        RECT 697.950 598.800 700.050 599.250 ;
        RECT 703.800 598.800 705.900 599.250 ;
        RECT 436.950 597.600 439.050 598.050 ;
        RECT 445.950 597.600 448.050 598.050 ;
        RECT 457.950 597.600 460.050 598.050 ;
        RECT 436.950 596.400 460.050 597.600 ;
        RECT 436.950 595.950 439.050 596.400 ;
        RECT 445.950 595.950 448.050 596.400 ;
        RECT 457.950 595.950 460.050 596.400 ;
        RECT 688.950 582.600 691.050 583.050 ;
        RECT 697.950 582.600 700.050 583.050 ;
        RECT 688.950 581.400 700.050 582.600 ;
        RECT 688.950 580.950 691.050 581.400 ;
        RECT 697.950 580.950 700.050 581.400 ;
        RECT 688.950 534.600 691.050 535.050 ;
        RECT 694.950 534.600 697.050 535.050 ;
        RECT 688.950 533.400 697.050 534.600 ;
        RECT 688.950 532.950 691.050 533.400 ;
        RECT 694.950 532.950 697.050 533.400 ;
        RECT 694.950 522.450 697.050 522.900 ;
        RECT 700.950 522.450 703.050 522.900 ;
        RECT 694.950 521.250 703.050 522.450 ;
        RECT 694.950 520.800 697.050 521.250 ;
        RECT 700.950 520.800 703.050 521.250 ;
    END
  END Cin[1]
  PIN Cin[0]
    PORT
      LAYER metal1 ;
        RECT 423.000 684.450 427.050 685.050 ;
        RECT 422.550 682.950 427.050 684.450 ;
        RECT 422.550 679.050 423.450 682.950 ;
        RECT 422.550 677.550 427.050 679.050 ;
        RECT 423.000 676.950 427.050 677.550 ;
        RECT 418.950 672.450 421.050 672.900 ;
        RECT 424.950 672.450 427.050 673.050 ;
        RECT 418.950 671.550 427.050 672.450 ;
        RECT 418.950 670.800 421.050 671.550 ;
        RECT 424.950 670.950 427.050 671.550 ;
        RECT 595.950 609.450 598.050 610.050 ;
        RECT 584.550 608.550 598.050 609.450 ;
        RECT 584.550 598.050 585.450 608.550 ;
        RECT 595.950 607.950 598.050 608.550 ;
        RECT 583.950 595.950 586.050 598.050 ;
        RECT 496.950 576.450 499.050 577.050 ;
        RECT 508.950 576.450 511.050 577.050 ;
        RECT 496.950 575.550 511.050 576.450 ;
        RECT 496.950 574.950 499.050 575.550 ;
        RECT 508.950 574.950 511.050 575.550 ;
      LAYER metal2 ;
        RECT 440.400 901.050 441.600 906.600 ;
        RECT 433.950 898.950 436.050 901.050 ;
        RECT 439.950 898.950 442.050 901.050 ;
        RECT 434.400 877.050 435.600 898.950 ;
        RECT 418.950 874.950 421.050 877.050 ;
        RECT 433.950 874.950 436.050 877.050 ;
        RECT 419.400 820.050 420.600 874.950 ;
        RECT 412.950 817.950 415.050 820.050 ;
        RECT 418.950 817.950 421.050 820.050 ;
        RECT 413.400 793.050 414.600 817.950 ;
        RECT 412.950 790.950 415.050 793.050 ;
        RECT 421.950 790.950 424.050 793.050 ;
        RECT 422.400 730.050 423.600 790.950 ;
        RECT 421.950 727.950 424.050 730.050 ;
        RECT 427.950 728.100 430.050 730.200 ;
        RECT 442.950 728.100 445.050 730.200 ;
        RECT 428.400 717.600 429.600 728.100 ;
        RECT 443.400 727.050 444.600 728.100 ;
        RECT 442.950 724.950 445.050 727.050 ;
        RECT 425.400 716.400 429.600 717.600 ;
        RECT 425.400 685.050 426.600 716.400 ;
        RECT 424.950 682.950 427.050 685.050 ;
        RECT 424.950 676.950 427.050 679.050 ;
        RECT 425.400 673.050 426.600 676.950 ;
        RECT 418.950 670.800 421.050 672.900 ;
        RECT 424.950 670.950 427.050 673.050 ;
        RECT 415.950 579.600 418.050 580.050 ;
        RECT 419.400 579.600 420.600 670.800 ;
        RECT 604.950 651.600 609.000 652.050 ;
        RECT 604.950 649.950 609.600 651.600 ;
        RECT 608.400 649.050 609.600 649.950 ;
        RECT 607.950 646.950 610.050 649.050 ;
        RECT 604.950 643.950 607.050 646.050 ;
        RECT 605.400 613.050 606.600 643.950 ;
        RECT 595.950 607.950 598.050 613.050 ;
        RECT 604.950 610.950 607.050 613.050 ;
        RECT 637.800 610.950 639.900 613.050 ;
        RECT 638.400 606.600 639.600 610.950 ;
        RECT 635.400 605.400 639.600 606.600 ;
        RECT 635.400 600.600 636.600 605.400 ;
        RECT 635.400 600.000 639.600 600.600 ;
        RECT 635.400 599.400 640.050 600.000 ;
        RECT 583.950 595.950 586.050 598.050 ;
        RECT 637.950 595.950 640.050 599.400 ;
        RECT 646.950 595.950 649.050 598.050 ;
        RECT 584.400 583.050 585.600 595.950 ;
        RECT 508.950 580.950 511.050 583.050 ;
        RECT 583.950 580.950 586.050 583.050 ;
        RECT 415.950 578.400 420.600 579.600 ;
        RECT 415.950 577.950 418.050 578.400 ;
        RECT 416.400 571.050 417.600 577.950 ;
        RECT 496.950 574.950 499.050 580.050 ;
        RECT 509.400 577.050 510.600 580.950 ;
        RECT 508.950 574.950 511.050 577.050 ;
        RECT 647.400 571.050 648.600 595.950 ;
        RECT 415.950 568.950 418.050 571.050 ;
        RECT 646.950 568.950 649.050 571.050 ;
      LAYER metal3 ;
        RECT 433.950 900.600 436.050 901.050 ;
        RECT 439.950 900.600 442.050 901.050 ;
        RECT 433.950 899.400 442.050 900.600 ;
        RECT 433.950 898.950 436.050 899.400 ;
        RECT 439.950 898.950 442.050 899.400 ;
        RECT 418.950 876.600 421.050 877.050 ;
        RECT 433.950 876.600 436.050 877.050 ;
        RECT 418.950 875.400 436.050 876.600 ;
        RECT 418.950 874.950 421.050 875.400 ;
        RECT 433.950 874.950 436.050 875.400 ;
        RECT 412.950 819.600 415.050 820.050 ;
        RECT 418.950 819.600 421.050 820.050 ;
        RECT 412.950 818.400 421.050 819.600 ;
        RECT 412.950 817.950 415.050 818.400 ;
        RECT 418.950 817.950 421.050 818.400 ;
        RECT 412.950 792.600 415.050 793.050 ;
        RECT 421.950 792.600 424.050 793.050 ;
        RECT 412.950 791.400 424.050 792.600 ;
        RECT 412.950 790.950 415.050 791.400 ;
        RECT 421.950 790.950 424.050 791.400 ;
        RECT 421.950 729.600 424.050 730.050 ;
        RECT 427.950 729.750 430.050 730.200 ;
        RECT 442.950 729.750 445.050 730.200 ;
        RECT 427.950 729.600 445.050 729.750 ;
        RECT 421.950 728.550 445.050 729.600 ;
        RECT 421.950 728.400 430.050 728.550 ;
        RECT 421.950 727.950 424.050 728.400 ;
        RECT 427.950 728.100 430.050 728.400 ;
        RECT 442.950 728.100 445.050 728.550 ;
        RECT 604.950 649.950 607.050 652.050 ;
        RECT 605.400 646.050 606.600 649.950 ;
        RECT 604.950 643.950 607.050 646.050 ;
        RECT 595.950 612.600 598.050 613.050 ;
        RECT 604.950 612.600 607.050 613.050 ;
        RECT 637.800 612.600 639.900 613.050 ;
        RECT 595.950 611.400 639.900 612.600 ;
        RECT 595.950 610.950 598.050 611.400 ;
        RECT 604.950 610.950 607.050 611.400 ;
        RECT 637.800 610.950 639.900 611.400 ;
        RECT 637.950 597.600 640.050 598.050 ;
        RECT 646.950 597.600 649.050 598.050 ;
        RECT 637.950 596.400 649.050 597.600 ;
        RECT 637.950 595.950 640.050 596.400 ;
        RECT 646.950 595.950 649.050 596.400 ;
        RECT 508.950 582.600 511.050 583.050 ;
        RECT 583.950 582.600 586.050 583.050 ;
        RECT 508.950 581.400 586.050 582.600 ;
        RECT 508.950 580.950 511.050 581.400 ;
        RECT 583.950 580.950 586.050 581.400 ;
        RECT 415.950 579.600 418.050 580.050 ;
        RECT 496.950 579.600 499.050 580.050 ;
        RECT 415.950 578.400 499.050 579.600 ;
        RECT 415.950 577.950 418.050 578.400 ;
        RECT 496.950 577.950 499.050 578.400 ;
    END
  END Cin[0]
  PIN Rdy
    PORT
      LAYER metal2 ;
        RECT 13.950 334.950 16.050 337.050 ;
        RECT 14.400 328.050 15.600 334.950 ;
        RECT 13.950 325.950 16.050 328.050 ;
      LAYER metal3 ;
        RECT -3.600 330.600 -2.400 333.600 ;
        RECT -3.600 329.400 0.600 330.600 ;
        RECT -0.600 327.600 0.600 329.400 ;
        RECT 13.950 327.600 16.050 328.050 ;
        RECT -0.600 326.400 16.050 327.600 ;
        RECT 13.950 325.950 16.050 326.400 ;
    END
  END Rdy
  PIN Vld
    PORT
      LAYER metal2 ;
        RECT 835.950 67.950 838.050 70.050 ;
        RECT 895.950 67.950 898.050 70.050 ;
        RECT 836.400 63.600 837.600 67.950 ;
        RECT 836.400 62.400 840.600 63.600 ;
        RECT 839.400 58.050 840.600 62.400 ;
        RECT 896.400 61.050 897.600 67.950 ;
        RECT 895.950 58.950 898.050 61.050 ;
        RECT 838.950 55.950 841.050 58.050 ;
      LAYER metal3 ;
        RECT 835.950 69.600 838.050 70.050 ;
        RECT 895.950 69.600 898.050 70.050 ;
        RECT 835.950 68.400 898.050 69.600 ;
        RECT 835.950 67.950 838.050 68.400 ;
        RECT 895.950 67.950 898.050 68.400 ;
        RECT 895.950 60.600 898.050 61.050 ;
        RECT 895.950 59.400 903.600 60.600 ;
        RECT 895.950 58.950 898.050 59.400 ;
    END
  END Vld
  PIN Xin[3]
    PORT
      LAYER metal1 ;
        RECT 22.950 573.450 27.000 574.050 ;
        RECT 22.950 571.950 27.450 573.450 ;
        RECT 26.550 567.450 27.450 571.950 ;
        RECT 31.950 567.450 34.050 568.050 ;
        RECT 26.550 566.550 34.050 567.450 ;
        RECT 31.950 565.950 34.050 566.550 ;
        RECT 454.950 534.450 457.050 535.050 ;
        RECT 463.950 534.450 466.050 535.050 ;
        RECT 454.950 533.550 466.050 534.450 ;
        RECT 454.950 532.950 457.050 533.550 ;
        RECT 463.950 532.950 466.050 533.550 ;
      LAYER metal2 ;
        RECT 22.950 577.950 25.050 580.050 ;
        RECT 23.400 574.050 24.600 577.950 ;
        RECT 22.950 571.950 25.050 574.050 ;
        RECT 31.950 565.950 34.050 568.050 ;
        RECT 32.400 547.050 33.600 565.950 ;
        RECT 31.950 544.950 34.050 547.050 ;
        RECT 367.950 544.950 370.050 547.050 ;
        RECT 454.950 544.950 457.050 547.050 ;
        RECT 368.400 526.050 369.600 544.950 ;
        RECT 455.400 535.050 456.600 544.950 ;
        RECT 454.950 532.950 457.050 535.050 ;
        RECT 463.950 532.950 466.050 535.050 ;
        RECT 464.400 526.050 465.600 532.950 ;
        RECT 367.950 523.950 370.050 526.050 ;
        RECT 463.950 523.950 466.050 526.050 ;
      LAYER metal3 ;
        RECT 22.950 579.600 25.050 580.050 ;
        RECT -3.600 578.400 25.050 579.600 ;
        RECT 22.950 577.950 25.050 578.400 ;
        RECT 31.950 546.600 34.050 547.050 ;
        RECT 367.950 546.600 370.050 547.050 ;
        RECT 454.950 546.600 457.050 547.050 ;
        RECT 31.950 545.400 457.050 546.600 ;
        RECT 31.950 544.950 34.050 545.400 ;
        RECT 367.950 544.950 370.050 545.400 ;
        RECT 454.950 544.950 457.050 545.400 ;
    END
  END Xin[3]
  PIN Xin[2]
    PORT
      LAYER metal2 ;
        RECT 1.950 625.800 4.050 627.900 ;
        RECT 127.950 625.950 130.050 628.050 ;
        RECT 2.400 574.050 3.600 625.800 ;
        RECT 128.400 616.050 129.600 625.950 ;
        RECT 127.950 613.950 130.050 616.050 ;
        RECT 283.950 613.950 286.050 616.050 ;
        RECT 284.400 580.050 285.600 613.950 ;
        RECT 283.950 577.950 286.050 580.050 ;
        RECT 403.950 577.950 406.050 580.050 ;
        RECT 1.950 571.950 4.050 574.050 ;
        RECT 404.400 559.050 405.600 577.950 ;
        RECT 445.950 568.950 448.050 571.050 ;
        RECT 490.950 568.950 493.050 571.050 ;
        RECT 446.400 559.050 447.600 568.950 ;
        RECT 403.950 556.950 406.050 559.050 ;
        RECT 445.950 556.950 448.050 559.050 ;
        RECT 446.400 553.050 447.600 556.950 ;
        RECT 491.400 553.050 492.600 568.950 ;
        RECT 445.950 550.950 448.050 553.050 ;
        RECT 490.950 550.950 493.050 553.050 ;
      LAYER metal3 ;
        RECT 1.950 627.600 4.050 627.900 ;
        RECT 127.950 627.600 130.050 628.050 ;
        RECT 1.950 626.400 130.050 627.600 ;
        RECT 1.950 625.800 4.050 626.400 ;
        RECT 127.950 625.950 130.050 626.400 ;
        RECT 127.950 615.600 130.050 616.050 ;
        RECT 283.950 615.600 286.050 616.050 ;
        RECT 127.950 614.400 286.050 615.600 ;
        RECT 127.950 613.950 130.050 614.400 ;
        RECT 283.950 613.950 286.050 614.400 ;
        RECT 283.950 579.600 286.050 580.050 ;
        RECT 403.950 579.600 406.050 580.050 ;
        RECT 283.950 578.400 406.050 579.600 ;
        RECT 283.950 577.950 286.050 578.400 ;
        RECT 403.950 577.950 406.050 578.400 ;
        RECT 1.950 573.600 4.050 574.050 ;
        RECT -3.600 572.400 4.050 573.600 ;
        RECT 1.950 571.950 4.050 572.400 ;
        RECT 403.950 558.600 406.050 559.050 ;
        RECT 445.950 558.600 448.050 559.050 ;
        RECT 403.950 557.400 448.050 558.600 ;
        RECT 403.950 556.950 406.050 557.400 ;
        RECT 445.950 556.950 448.050 557.400 ;
        RECT 445.950 552.600 448.050 553.050 ;
        RECT 490.950 552.600 493.050 553.050 ;
        RECT 445.950 551.400 493.050 552.600 ;
        RECT 445.950 550.950 448.050 551.400 ;
        RECT 490.950 550.950 493.050 551.400 ;
    END
  END Xin[2]
  PIN Xin[1]
    PORT
      LAYER metal2 ;
        RECT 469.950 568.950 472.050 571.050 ;
        RECT 508.950 568.950 511.050 571.050 ;
        RECT 1.950 565.950 4.050 568.050 ;
        RECT 2.400 559.050 3.600 565.950 ;
        RECT 470.400 562.050 471.600 568.950 ;
        RECT 509.400 562.050 510.600 568.950 ;
        RECT 400.950 559.950 403.050 562.050 ;
        RECT 469.950 559.950 472.050 562.050 ;
        RECT 508.950 559.950 511.050 562.050 ;
        RECT 1.950 556.950 4.050 559.050 ;
        RECT 55.950 556.800 58.050 558.900 ;
        RECT 56.400 553.050 57.600 556.800 ;
        RECT 401.400 553.050 402.600 559.950 ;
        RECT 55.950 550.950 58.050 553.050 ;
        RECT 400.950 550.950 403.050 553.050 ;
      LAYER metal3 ;
        RECT 1.950 567.600 4.050 568.050 ;
        RECT -3.600 566.400 4.050 567.600 ;
        RECT 1.950 565.950 4.050 566.400 ;
        RECT 400.950 561.600 403.050 562.050 ;
        RECT 469.950 561.600 474.000 562.050 ;
        RECT 508.950 561.600 511.050 562.050 ;
        RECT 400.950 560.400 474.600 561.600 ;
        RECT 400.950 559.950 403.050 560.400 ;
        RECT 469.950 559.950 474.600 560.400 ;
        RECT 1.950 558.600 4.050 559.050 ;
        RECT 55.950 558.600 58.050 558.900 ;
        RECT 1.950 557.400 58.050 558.600 ;
        RECT 473.400 558.600 474.600 559.950 ;
        RECT 500.400 560.400 511.050 561.600 ;
        RECT 500.400 558.600 501.600 560.400 ;
        RECT 508.950 559.950 511.050 560.400 ;
        RECT 473.400 557.400 501.600 558.600 ;
        RECT 1.950 556.950 4.050 557.400 ;
        RECT 55.950 556.800 58.050 557.400 ;
        RECT 55.950 552.600 58.050 553.050 ;
        RECT 400.950 552.600 403.050 553.050 ;
        RECT 55.950 551.400 403.050 552.600 ;
        RECT 55.950 550.950 58.050 551.400 ;
        RECT 400.950 550.950 403.050 551.400 ;
    END
  END Xin[1]
  PIN Xin[0]
    PORT
      LAYER metal2 ;
        RECT 403.950 490.950 406.050 493.050 ;
        RECT 268.950 484.950 271.050 487.050 ;
        RECT 269.400 481.050 270.600 484.950 ;
        RECT 404.400 484.050 405.600 490.950 ;
        RECT 367.950 481.950 370.050 484.050 ;
        RECT 403.950 481.950 406.050 484.050 ;
        RECT 430.950 481.950 433.050 484.050 ;
        RECT 13.950 478.950 16.050 481.050 ;
        RECT 268.950 478.950 271.050 481.050 ;
        RECT 14.400 453.600 15.600 478.950 ;
        RECT 368.400 469.050 369.600 481.950 ;
        RECT 404.400 469.050 405.600 481.950 ;
        RECT 367.950 466.950 370.050 469.050 ;
        RECT 403.950 466.950 406.050 469.050 ;
        RECT 11.400 453.000 15.600 453.600 ;
        RECT 10.950 452.400 15.600 453.000 ;
        RECT 10.950 451.050 13.050 452.400 ;
        RECT 10.800 450.000 13.050 451.050 ;
        RECT 10.800 448.950 12.900 450.000 ;
        RECT 431.400 436.050 432.600 481.950 ;
        RECT 430.950 433.950 433.050 436.050 ;
        RECT 484.950 433.950 487.050 436.050 ;
        RECT 485.400 418.050 486.600 433.950 ;
        RECT 484.950 415.950 487.050 418.050 ;
        RECT 493.950 412.950 496.050 415.050 ;
        RECT 494.400 411.900 495.600 412.950 ;
        RECT 493.950 409.800 496.050 411.900 ;
      LAYER metal3 ;
        RECT 268.950 486.600 271.050 487.050 ;
        RECT 268.950 485.400 309.600 486.600 ;
        RECT 268.950 484.950 271.050 485.400 ;
        RECT 308.400 483.600 309.600 485.400 ;
        RECT 367.950 483.600 370.050 484.050 ;
        RECT 308.400 482.400 370.050 483.600 ;
        RECT 367.950 481.950 370.050 482.400 ;
        RECT 403.950 483.600 406.050 484.050 ;
        RECT 430.950 483.600 433.050 484.050 ;
        RECT 403.950 482.400 433.050 483.600 ;
        RECT 403.950 481.950 406.050 482.400 ;
        RECT 430.950 481.950 433.050 482.400 ;
        RECT 13.950 480.600 16.050 481.050 ;
        RECT 268.950 480.600 271.050 481.050 ;
        RECT 13.950 479.400 271.050 480.600 ;
        RECT 13.950 478.950 16.050 479.400 ;
        RECT 268.950 478.950 271.050 479.400 ;
        RECT 367.950 468.600 370.050 469.050 ;
        RECT 403.950 468.600 406.050 469.050 ;
        RECT 367.950 467.400 406.050 468.600 ;
        RECT 367.950 466.950 370.050 467.400 ;
        RECT 403.950 466.950 406.050 467.400 ;
        RECT 10.800 450.600 12.900 451.050 ;
        RECT -3.600 449.400 12.900 450.600 ;
        RECT 10.800 448.950 12.900 449.400 ;
        RECT 430.950 435.600 433.050 436.050 ;
        RECT 484.950 435.600 487.050 436.050 ;
        RECT 430.950 434.400 487.050 435.600 ;
        RECT 430.950 433.950 433.050 434.400 ;
        RECT 484.950 433.950 487.050 434.400 ;
        RECT 484.950 417.600 487.050 418.050 ;
        RECT 484.950 416.400 492.600 417.600 ;
        RECT 484.950 415.950 487.050 416.400 ;
        RECT 491.400 414.600 492.600 416.400 ;
        RECT 491.400 413.400 495.600 414.600 ;
        RECT 494.400 411.900 495.600 413.400 ;
        RECT 493.950 409.800 496.050 411.900 ;
    END
  END Xin[0]
  PIN Xout[3]
    PORT
      LAYER metal2 ;
        RECT 889.950 683.100 892.050 685.200 ;
        RECT 890.400 682.050 891.600 683.100 ;
        RECT 889.950 679.950 892.050 682.050 ;
      LAYER metal3 ;
        RECT 889.950 684.600 892.050 685.200 ;
        RECT 889.950 683.400 903.600 684.600 ;
        RECT 889.950 683.100 892.050 683.400 ;
    END
  END Xout[3]
  PIN Xout[2]
    PORT
      LAYER metal2 ;
        RECT 826.950 658.950 829.050 661.050 ;
        RECT 817.950 646.950 820.050 649.050 ;
        RECT 818.400 645.900 819.600 646.950 ;
        RECT 827.400 646.050 828.600 658.950 ;
        RECT 895.950 655.950 898.050 658.050 ;
        RECT 896.400 649.050 897.600 655.950 ;
        RECT 895.950 646.950 898.050 649.050 ;
        RECT 817.950 643.800 820.050 645.900 ;
        RECT 826.950 643.950 829.050 646.050 ;
      LAYER metal3 ;
        RECT 826.950 660.600 829.050 661.050 ;
        RECT 826.950 659.400 861.600 660.600 ;
        RECT 826.950 658.950 829.050 659.400 ;
        RECT 860.400 657.600 861.600 659.400 ;
        RECT 895.950 657.600 898.050 658.050 ;
        RECT 860.400 656.400 898.050 657.600 ;
        RECT 895.950 655.950 898.050 656.400 ;
        RECT 895.950 648.600 898.050 649.050 ;
        RECT 895.950 647.400 903.600 648.600 ;
        RECT 895.950 646.950 898.050 647.400 ;
        RECT 817.950 645.600 820.050 645.900 ;
        RECT 826.950 645.600 829.050 646.050 ;
        RECT 817.950 644.400 829.050 645.600 ;
        RECT 902.400 644.400 903.600 647.400 ;
        RECT 817.950 643.800 820.050 644.400 ;
        RECT 826.950 643.950 829.050 644.400 ;
    END
  END Xout[2]
  PIN Xout[1]
    PORT
      LAYER metal2 ;
        RECT 745.950 622.800 748.050 624.900 ;
        RECT 895.950 622.950 898.050 625.050 ;
        RECT 746.400 613.050 747.600 622.800 ;
        RECT 688.950 610.950 691.050 613.050 ;
        RECT 745.950 610.950 748.050 613.050 ;
        RECT 689.400 604.050 690.600 610.950 ;
        RECT 896.400 607.050 897.600 622.950 ;
        RECT 895.950 604.950 898.050 607.050 ;
        RECT 688.950 601.950 691.050 604.050 ;
      LAYER metal3 ;
        RECT 745.950 624.600 748.050 624.900 ;
        RECT 895.950 624.600 898.050 625.050 ;
        RECT 745.950 623.400 898.050 624.600 ;
        RECT 745.950 622.800 748.050 623.400 ;
        RECT 895.950 622.950 898.050 623.400 ;
        RECT 688.950 612.600 691.050 613.050 ;
        RECT 745.950 612.600 748.050 613.050 ;
        RECT 688.950 611.400 748.050 612.600 ;
        RECT 688.950 610.950 691.050 611.400 ;
        RECT 745.950 610.950 748.050 611.400 ;
        RECT 895.950 606.600 898.050 607.050 ;
        RECT 895.950 605.400 903.600 606.600 ;
        RECT 895.950 604.950 898.050 605.400 ;
    END
  END Xout[1]
  PIN Xout[0]
    PORT
      LAYER metal2 ;
        RECT 553.950 490.950 556.050 493.050 ;
        RECT 554.400 475.050 555.600 490.950 ;
        RECT 895.950 487.950 898.050 490.050 ;
        RECT 896.400 481.050 897.600 487.950 ;
        RECT 832.950 478.800 835.050 480.900 ;
        RECT 895.950 478.950 898.050 481.050 ;
        RECT 553.950 472.950 556.050 475.050 ;
        RECT 833.400 472.050 834.600 478.800 ;
        RECT 832.950 469.950 835.050 472.050 ;
      LAYER metal3 ;
        RECT 895.950 489.600 898.050 490.050 ;
        RECT 895.950 488.400 903.600 489.600 ;
        RECT 895.950 487.950 898.050 488.400 ;
        RECT 832.950 480.600 835.050 480.900 ;
        RECT 895.950 480.600 898.050 481.050 ;
        RECT 832.950 479.400 898.050 480.600 ;
        RECT 832.950 478.800 835.050 479.400 ;
        RECT 895.950 478.950 898.050 479.400 ;
        RECT 553.950 474.600 556.050 475.050 ;
        RECT 553.950 473.400 753.600 474.600 ;
        RECT 553.950 472.950 556.050 473.400 ;
        RECT 752.400 471.600 753.600 473.400 ;
        RECT 832.950 471.600 835.050 472.050 ;
        RECT 752.400 470.400 835.050 471.600 ;
        RECT 832.950 469.950 835.050 470.400 ;
    END
  END Xout[0]
  PIN Yin[3]
    PORT
      LAYER metal1 ;
        RECT 274.950 51.450 277.050 52.050 ;
        RECT 283.950 51.450 286.050 52.050 ;
        RECT 274.950 50.550 286.050 51.450 ;
        RECT 274.950 49.950 277.050 50.550 ;
        RECT 283.950 49.950 286.050 50.550 ;
      LAYER metal2 ;
        RECT 283.950 55.950 286.050 58.050 ;
        RECT 284.400 54.000 285.600 55.950 ;
        RECT 274.950 49.950 277.050 52.050 ;
        RECT 283.950 49.950 286.050 54.000 ;
        RECT 275.400 31.050 276.600 49.950 ;
        RECT 274.950 28.950 277.050 31.050 ;
        RECT 283.950 16.950 286.050 19.050 ;
        RECT 284.400 -2.400 285.600 16.950 ;
        RECT 284.400 -3.600 288.600 -2.400 ;
      LAYER metal3 ;
        RECT 274.950 28.950 277.050 31.050 ;
        RECT 275.400 24.600 276.600 28.950 ;
        RECT 275.400 23.400 279.600 24.600 ;
        RECT 278.400 18.600 279.600 23.400 ;
        RECT 283.950 18.600 286.050 19.050 ;
        RECT 278.400 17.400 286.050 18.600 ;
        RECT 283.950 16.950 286.050 17.400 ;
    END
  END Yin[3]
  PIN Yin[2]
    PORT
      LAYER metal2 ;
        RECT 433.950 55.950 436.050 58.050 ;
        RECT 434.400 31.050 435.600 55.950 ;
        RECT 433.950 28.950 436.050 31.050 ;
        RECT 439.950 28.950 442.050 31.050 ;
        RECT 440.400 -2.400 441.600 28.950 ;
        RECT 437.400 -3.600 441.600 -2.400 ;
      LAYER metal3 ;
        RECT 433.950 30.600 436.050 31.050 ;
        RECT 439.950 30.600 442.050 31.050 ;
        RECT 433.950 29.400 442.050 30.600 ;
        RECT 433.950 28.950 436.050 29.400 ;
        RECT 439.950 28.950 442.050 29.400 ;
    END
  END Yin[2]
  PIN Yin[1]
    PORT
      LAYER metal2 ;
        RECT 505.950 26.100 508.050 28.200 ;
        RECT 506.400 25.050 507.600 26.100 ;
        RECT 505.950 22.950 508.050 25.050 ;
        RECT 502.950 19.950 505.050 22.050 ;
        RECT 503.400 4.050 504.600 19.950 ;
        RECT 502.950 1.950 505.050 4.050 ;
        RECT 508.950 1.950 511.050 4.050 ;
        RECT 509.400 -3.600 510.600 1.950 ;
      LAYER metal3 ;
        RECT 505.950 27.600 508.050 28.200 ;
        RECT 503.400 26.400 508.050 27.600 ;
        RECT 503.400 22.050 504.600 26.400 ;
        RECT 505.950 26.100 508.050 26.400 ;
        RECT 502.950 19.950 505.050 22.050 ;
        RECT 502.950 3.600 505.050 4.050 ;
        RECT 508.950 3.600 511.050 4.050 ;
        RECT 502.950 2.400 511.050 3.600 ;
        RECT 502.950 1.950 505.050 2.400 ;
        RECT 508.950 1.950 511.050 2.400 ;
    END
  END Yin[1]
  PIN Yin[0]
    PORT
      LAYER metal2 ;
        RECT 526.950 55.950 529.050 58.050 ;
        RECT 527.400 34.050 528.600 55.950 ;
        RECT 517.950 31.950 520.050 34.050 ;
        RECT 526.950 31.950 529.050 34.050 ;
        RECT 518.400 4.050 519.600 31.950 ;
        RECT 517.950 1.950 520.050 4.050 ;
        RECT 523.950 1.950 526.050 4.050 ;
        RECT 524.400 -3.600 525.600 1.950 ;
      LAYER metal3 ;
        RECT 517.950 33.600 520.050 34.050 ;
        RECT 526.950 33.600 529.050 34.050 ;
        RECT 517.950 32.400 529.050 33.600 ;
        RECT 517.950 31.950 520.050 32.400 ;
        RECT 526.950 31.950 529.050 32.400 ;
        RECT 517.950 3.600 520.050 4.050 ;
        RECT 523.950 3.600 526.050 4.050 ;
        RECT 517.950 2.400 526.050 3.600 ;
        RECT 517.950 1.950 520.050 2.400 ;
        RECT 523.950 1.950 526.050 2.400 ;
    END
  END Yin[0]
  PIN Yout[3]
    PORT
      LAYER metal2 ;
        RECT 7.950 136.950 10.050 139.050 ;
        RECT 13.950 137.100 16.050 139.200 ;
        RECT 8.400 4.050 9.600 136.950 ;
        RECT 14.400 136.050 15.600 137.100 ;
        RECT 13.950 133.950 16.050 136.050 ;
        RECT 7.950 1.950 10.050 4.050 ;
        RECT 13.950 1.950 16.050 4.050 ;
        RECT 14.400 -3.600 15.600 1.950 ;
      LAYER metal3 ;
        RECT 7.950 138.600 10.050 139.050 ;
        RECT 13.950 138.600 16.050 139.200 ;
        RECT 7.950 137.400 16.050 138.600 ;
        RECT 7.950 136.950 10.050 137.400 ;
        RECT 13.950 137.100 16.050 137.400 ;
        RECT 7.950 3.600 10.050 4.050 ;
        RECT 13.950 3.600 16.050 4.050 ;
        RECT 7.950 2.400 16.050 3.600 ;
        RECT 7.950 1.950 10.050 2.400 ;
        RECT 13.950 1.950 16.050 2.400 ;
    END
  END Yout[3]
  PIN Yout[2]
    PORT
      LAYER metal2 ;
        RECT 52.950 22.950 55.050 25.050 ;
        RECT 53.400 -3.600 54.600 22.950 ;
    END
  END Yout[2]
  PIN Yout[1]
    PORT
      LAYER metal2 ;
        RECT 73.950 22.950 76.050 25.050 ;
        RECT 74.400 -3.600 75.600 22.950 ;
    END
  END Yout[1]
  PIN Yout[0]
    PORT
      LAYER metal2 ;
        RECT 148.950 100.950 151.050 103.050 ;
        RECT 149.400 70.050 150.600 100.950 ;
        RECT 148.950 67.950 151.050 70.050 ;
        RECT 154.950 67.950 157.050 70.050 ;
        RECT 155.400 64.050 156.600 67.950 ;
        RECT 154.950 61.950 157.050 64.050 ;
        RECT 157.950 51.600 160.050 55.050 ;
        RECT 155.400 51.000 160.050 51.600 ;
        RECT 155.400 50.400 159.600 51.000 ;
        RECT 155.400 43.050 156.600 50.400 ;
        RECT 142.950 40.950 145.050 43.050 ;
        RECT 154.950 40.950 157.050 43.050 ;
        RECT 143.400 -2.400 144.600 40.950 ;
        RECT 143.400 -3.600 147.600 -2.400 ;
      LAYER metal3 ;
        RECT 148.950 69.600 151.050 70.050 ;
        RECT 154.950 69.600 157.050 70.050 ;
        RECT 148.950 68.400 157.050 69.600 ;
        RECT 148.950 67.950 151.050 68.400 ;
        RECT 154.950 67.950 157.050 68.400 ;
        RECT 154.950 63.600 159.000 64.050 ;
        RECT 154.950 61.950 159.600 63.600 ;
        RECT 158.400 55.050 159.600 61.950 ;
        RECT 157.950 52.950 160.050 55.050 ;
        RECT 142.950 42.600 145.050 43.050 ;
        RECT 154.950 42.600 157.050 43.050 ;
        RECT 142.950 41.400 157.050 42.600 ;
        RECT 142.950 40.950 145.050 41.400 ;
        RECT 154.950 40.950 157.050 41.400 ;
    END
  END Yout[0]
  PIN clk
    PORT
      LAYER metal2 ;
        RECT 122.400 901.050 123.600 906.600 ;
        RECT 121.950 898.950 124.050 901.050 ;
        RECT 136.950 898.950 139.050 901.050 ;
        RECT 124.950 880.950 127.050 883.050 ;
        RECT 125.400 879.000 126.600 880.950 ;
        RECT 124.950 874.950 127.050 879.000 ;
        RECT 137.400 877.050 138.600 898.950 ;
        RECT 136.950 874.950 139.050 877.050 ;
        RECT 137.400 820.050 138.600 874.950 ;
        RECT 136.950 817.950 139.050 820.050 ;
        RECT 145.950 817.950 148.050 820.050 ;
        RECT 146.400 796.050 147.600 817.950 ;
        RECT 145.950 793.950 148.050 796.050 ;
        RECT 169.950 793.950 172.050 796.050 ;
        RECT 170.400 756.600 171.600 793.950 ;
        RECT 170.400 755.400 174.600 756.600 ;
        RECT 173.400 708.600 174.600 755.400 ;
        RECT 170.400 707.400 174.600 708.600 ;
        RECT 170.400 628.050 171.600 707.400 ;
        RECT 169.950 625.950 172.050 628.050 ;
        RECT 259.950 625.950 262.050 628.050 ;
        RECT 260.400 556.050 261.600 625.950 ;
        RECT 289.950 568.950 292.050 571.050 ;
        RECT 352.950 568.950 355.050 571.050 ;
        RECT 290.400 556.050 291.600 568.950 ;
        RECT 353.400 559.050 354.600 568.950 ;
        RECT 352.950 556.950 355.050 559.050 ;
        RECT 361.950 556.950 364.050 559.050 ;
        RECT 259.950 553.950 262.050 556.050 ;
        RECT 289.950 553.950 292.050 556.050 ;
        RECT 362.400 523.050 363.600 556.950 ;
        RECT 361.950 520.950 364.050 523.050 ;
        RECT 394.950 520.950 397.050 523.050 ;
        RECT 395.400 466.050 396.600 520.950 ;
        RECT 394.950 463.950 397.050 466.050 ;
        RECT 403.950 463.800 406.050 465.900 ;
        RECT 404.400 352.050 405.600 463.800 ;
        RECT 382.950 349.950 385.050 352.050 ;
        RECT 403.950 349.950 406.050 352.050 ;
        RECT 349.950 334.950 352.050 337.050 ;
        RECT 350.400 333.900 351.600 334.950 ;
        RECT 383.400 333.900 384.600 349.950 ;
        RECT 349.950 331.800 352.050 333.900 ;
        RECT 382.950 331.800 385.050 333.900 ;
        RECT 350.400 322.050 351.600 331.800 ;
        RECT 349.950 319.950 352.050 322.050 ;
        RECT 82.950 316.950 85.050 319.050 ;
        RECT 124.950 316.950 127.050 319.050 ;
        RECT 184.950 316.950 187.050 319.050 ;
        RECT 83.400 307.050 84.600 316.950 ;
        RECT 125.400 310.050 126.600 316.950 ;
        RECT 185.400 310.050 186.600 316.950 ;
        RECT 124.950 307.950 127.050 310.050 ;
        RECT 184.950 307.950 187.050 310.050 ;
        RECT 28.950 304.950 31.050 307.050 ;
        RECT 34.950 304.950 37.050 307.050 ;
        RECT 82.950 304.950 85.050 307.050 ;
        RECT 19.950 253.950 22.050 256.050 ;
        RECT 29.400 255.900 30.600 304.950 ;
        RECT 35.400 292.050 36.600 304.950 ;
        RECT 34.950 289.950 37.050 292.050 ;
        RECT 34.950 256.950 37.050 259.050 ;
        RECT 35.400 255.900 36.600 256.950 ;
        RECT 20.400 199.050 21.600 253.950 ;
        RECT 28.950 253.800 31.050 255.900 ;
        RECT 34.950 253.800 37.050 255.900 ;
        RECT 383.400 238.050 384.600 331.800 ;
        RECT 382.950 235.950 385.050 238.050 ;
        RECT 388.950 235.950 391.050 238.050 ;
        RECT 389.400 208.050 390.600 235.950 ;
        RECT 382.950 205.950 385.050 208.050 ;
        RECT 388.950 205.950 391.050 208.050 ;
        RECT 7.950 196.950 10.050 199.050 ;
        RECT 19.950 196.950 22.050 199.050 ;
        RECT 8.400 145.050 9.600 196.950 ;
        RECT 383.400 160.050 384.600 205.950 ;
        RECT 382.950 157.950 385.050 160.050 ;
        RECT 391.950 157.950 394.050 160.050 ;
        RECT 7.950 142.950 10.050 145.050 ;
        RECT 34.950 142.950 37.050 145.050 ;
        RECT 35.400 136.050 36.600 142.950 ;
        RECT 392.400 136.050 393.600 157.950 ;
        RECT 34.950 133.950 37.050 136.050 ;
        RECT 391.950 133.950 394.050 136.050 ;
      LAYER metal3 ;
        RECT 121.950 900.600 124.050 901.050 ;
        RECT 136.950 900.600 139.050 901.050 ;
        RECT 121.950 899.400 139.050 900.600 ;
        RECT 121.950 898.950 124.050 899.400 ;
        RECT 136.950 898.950 139.050 899.400 ;
        RECT 124.950 876.600 127.050 877.050 ;
        RECT 136.950 876.600 139.050 877.050 ;
        RECT 124.950 875.400 139.050 876.600 ;
        RECT 124.950 874.950 127.050 875.400 ;
        RECT 136.950 874.950 139.050 875.400 ;
        RECT 136.950 819.600 139.050 820.050 ;
        RECT 145.950 819.600 148.050 820.050 ;
        RECT 136.950 818.400 148.050 819.600 ;
        RECT 136.950 817.950 139.050 818.400 ;
        RECT 145.950 817.950 148.050 818.400 ;
        RECT 145.950 795.600 148.050 796.050 ;
        RECT 169.950 795.600 172.050 796.050 ;
        RECT 145.950 794.400 172.050 795.600 ;
        RECT 145.950 793.950 148.050 794.400 ;
        RECT 169.950 793.950 172.050 794.400 ;
        RECT 169.950 627.600 172.050 628.050 ;
        RECT 259.950 627.600 262.050 628.050 ;
        RECT 169.950 626.400 262.050 627.600 ;
        RECT 169.950 625.950 172.050 626.400 ;
        RECT 259.950 625.950 262.050 626.400 ;
        RECT 352.950 558.600 355.050 559.050 ;
        RECT 361.950 558.600 364.050 559.050 ;
        RECT 352.950 557.400 364.050 558.600 ;
        RECT 352.950 556.950 355.050 557.400 ;
        RECT 361.950 556.950 364.050 557.400 ;
        RECT 259.950 555.600 262.050 556.050 ;
        RECT 289.950 555.600 292.050 556.050 ;
        RECT 353.400 555.600 354.600 556.950 ;
        RECT 259.950 554.400 354.600 555.600 ;
        RECT 259.950 553.950 262.050 554.400 ;
        RECT 289.950 553.950 292.050 554.400 ;
        RECT 361.950 522.600 364.050 523.050 ;
        RECT 394.950 522.600 397.050 523.050 ;
        RECT 361.950 521.400 397.050 522.600 ;
        RECT 361.950 520.950 364.050 521.400 ;
        RECT 394.950 520.950 397.050 521.400 ;
        RECT 394.950 465.600 397.050 466.050 ;
        RECT 403.950 465.600 406.050 465.900 ;
        RECT 394.950 464.400 406.050 465.600 ;
        RECT 394.950 463.950 397.050 464.400 ;
        RECT 403.950 463.800 406.050 464.400 ;
        RECT 382.950 351.600 385.050 352.050 ;
        RECT 403.950 351.600 406.050 352.050 ;
        RECT 382.950 350.400 406.050 351.600 ;
        RECT 382.950 349.950 385.050 350.400 ;
        RECT 403.950 349.950 406.050 350.400 ;
        RECT 349.950 333.450 352.050 333.900 ;
        RECT 382.950 333.450 385.050 333.900 ;
        RECT 349.950 332.250 385.050 333.450 ;
        RECT 349.950 331.800 352.050 332.250 ;
        RECT 382.950 331.800 385.050 332.250 ;
        RECT 349.950 321.600 352.050 322.050 ;
        RECT 278.400 320.400 352.050 321.600 ;
        RECT 82.950 318.600 85.050 319.050 ;
        RECT 124.950 318.600 127.050 319.050 ;
        RECT 82.950 317.400 127.050 318.600 ;
        RECT 82.950 316.950 85.050 317.400 ;
        RECT 124.950 316.950 127.050 317.400 ;
        RECT 184.950 318.600 187.050 319.050 ;
        RECT 278.400 318.600 279.600 320.400 ;
        RECT 349.950 319.950 352.050 320.400 ;
        RECT 184.950 317.400 279.600 318.600 ;
        RECT 184.950 316.950 187.050 317.400 ;
        RECT 124.950 309.600 127.050 310.050 ;
        RECT 184.950 309.600 187.050 310.050 ;
        RECT 124.950 308.400 187.050 309.600 ;
        RECT 124.950 307.950 127.050 308.400 ;
        RECT 184.950 307.950 187.050 308.400 ;
        RECT 28.950 306.600 31.050 307.050 ;
        RECT 34.950 306.600 37.050 307.050 ;
        RECT 82.950 306.600 85.050 307.050 ;
        RECT 28.950 305.400 85.050 306.600 ;
        RECT 28.950 304.950 31.050 305.400 ;
        RECT 34.950 304.950 37.050 305.400 ;
        RECT 82.950 304.950 85.050 305.400 ;
        RECT 19.950 255.600 22.050 256.050 ;
        RECT 28.950 255.600 31.050 255.900 ;
        RECT 19.950 255.450 31.050 255.600 ;
        RECT 34.950 255.450 37.050 255.900 ;
        RECT 19.950 254.400 37.050 255.450 ;
        RECT 19.950 253.950 22.050 254.400 ;
        RECT 28.950 254.250 37.050 254.400 ;
        RECT 28.950 253.800 31.050 254.250 ;
        RECT 34.950 253.800 37.050 254.250 ;
        RECT 382.950 237.600 385.050 238.050 ;
        RECT 388.950 237.600 391.050 238.050 ;
        RECT 382.950 236.400 391.050 237.600 ;
        RECT 382.950 235.950 385.050 236.400 ;
        RECT 388.950 235.950 391.050 236.400 ;
        RECT 382.950 207.600 385.050 208.050 ;
        RECT 388.950 207.600 391.050 208.050 ;
        RECT 382.950 206.400 391.050 207.600 ;
        RECT 382.950 205.950 385.050 206.400 ;
        RECT 388.950 205.950 391.050 206.400 ;
        RECT 7.950 198.600 10.050 199.050 ;
        RECT 19.950 198.600 22.050 199.050 ;
        RECT 7.950 197.400 22.050 198.600 ;
        RECT 7.950 196.950 10.050 197.400 ;
        RECT 19.950 196.950 22.050 197.400 ;
        RECT 382.950 159.600 385.050 160.050 ;
        RECT 391.950 159.600 394.050 160.050 ;
        RECT 382.950 158.400 394.050 159.600 ;
        RECT 382.950 157.950 385.050 158.400 ;
        RECT 391.950 157.950 394.050 158.400 ;
        RECT 7.950 144.600 10.050 145.050 ;
        RECT 34.950 144.600 37.050 145.050 ;
        RECT 7.950 143.400 37.050 144.600 ;
        RECT 7.950 142.950 10.050 143.400 ;
        RECT 34.950 142.950 37.050 143.400 ;
    END
  END clk
  OBS
      LAYER metal1 ;
        RECT 13.800 893.400 15.600 896.400 ;
        RECT 14.400 883.050 15.600 893.400 ;
        RECT 34.800 889.200 36.600 896.400 ;
        RECT 32.400 888.300 36.600 889.200 ;
        RECT 41.550 890.400 43.350 896.400 ;
        RECT 49.650 893.400 51.450 896.400 ;
        RECT 57.450 893.400 59.250 896.400 ;
        RECT 65.250 894.300 67.050 896.400 ;
        RECT 65.250 893.400 69.000 894.300 ;
        RECT 49.650 892.500 50.700 893.400 ;
        RECT 46.950 891.300 50.700 892.500 ;
        RECT 58.200 892.500 59.250 893.400 ;
        RECT 67.950 892.500 69.000 893.400 ;
        RECT 58.200 891.450 63.150 892.500 ;
        RECT 46.950 890.400 49.050 891.300 ;
        RECT 61.350 890.700 63.150 891.450 ;
        RECT 29.100 883.050 30.900 884.850 ;
        RECT 32.400 883.050 33.600 888.300 ;
        RECT 35.100 883.050 36.900 884.850 ;
        RECT 41.550 883.050 42.750 890.400 ;
        RECT 64.650 889.800 66.450 891.600 ;
        RECT 67.950 890.400 70.050 892.500 ;
        RECT 73.050 890.400 74.850 896.400 ;
        RECT 54.150 888.000 55.950 888.600 ;
        RECT 65.100 888.000 66.150 889.800 ;
        RECT 54.150 886.800 66.150 888.000 ;
        RECT 13.950 880.950 16.050 883.050 ;
        RECT 16.950 880.950 19.050 883.050 ;
        RECT 28.950 880.950 31.050 883.050 ;
        RECT 31.950 880.950 34.050 883.050 ;
        RECT 34.950 880.950 37.050 883.050 ;
        RECT 41.550 881.250 47.850 883.050 ;
        RECT 41.550 880.950 46.050 881.250 ;
        RECT 14.400 867.600 15.600 880.950 ;
        RECT 17.100 879.150 18.900 880.950 ;
        RECT 13.800 861.600 15.600 867.600 ;
        RECT 32.400 867.600 33.600 880.950 ;
        RECT 41.550 873.600 42.750 880.950 ;
        RECT 43.950 875.400 45.750 877.200 ;
        RECT 44.850 874.200 49.050 875.400 ;
        RECT 54.150 874.200 55.050 886.800 ;
        RECT 65.100 885.600 72.000 886.800 ;
        RECT 65.100 885.000 66.900 885.600 ;
        RECT 71.100 884.850 72.000 885.600 ;
        RECT 68.100 883.800 69.900 884.400 ;
        RECT 61.950 882.600 69.900 883.800 ;
        RECT 71.100 883.050 72.900 884.850 ;
        RECT 61.950 880.950 64.050 882.600 ;
        RECT 70.950 880.950 73.050 883.050 ;
        RECT 63.750 875.700 65.550 876.000 ;
        RECT 73.950 875.700 74.850 890.400 ;
        RECT 63.750 875.100 74.850 875.700 ;
        RECT 32.400 861.600 34.200 867.600 ;
        RECT 41.550 861.600 43.350 873.600 ;
        RECT 46.950 873.300 49.050 874.200 ;
        RECT 49.950 873.300 55.050 874.200 ;
        RECT 57.150 874.500 74.850 875.100 ;
        RECT 57.150 874.200 65.550 874.500 ;
        RECT 49.950 872.400 50.850 873.300 ;
        RECT 48.150 870.600 50.850 872.400 ;
        RECT 51.750 872.100 53.550 872.400 ;
        RECT 57.150 872.100 58.050 874.200 ;
        RECT 73.950 873.600 74.850 874.500 ;
        RECT 51.750 871.200 58.050 872.100 ;
        RECT 58.950 872.700 60.750 873.300 ;
        RECT 58.950 871.500 66.450 872.700 ;
        RECT 51.750 870.600 53.550 871.200 ;
        RECT 65.250 870.600 66.450 871.500 ;
        RECT 46.950 867.600 50.850 869.700 ;
        RECT 55.950 869.550 57.750 870.300 ;
        RECT 60.750 869.550 62.550 870.300 ;
        RECT 55.950 868.500 62.550 869.550 ;
        RECT 65.250 868.500 70.050 870.600 ;
        RECT 49.050 861.600 50.850 867.600 ;
        RECT 56.850 861.600 58.650 868.500 ;
        RECT 65.250 867.600 66.450 868.500 ;
        RECT 64.650 861.600 66.450 867.600 ;
        RECT 73.050 861.600 74.850 873.600 ;
        RECT 77.550 890.400 79.350 896.400 ;
        RECT 85.650 893.400 87.450 896.400 ;
        RECT 93.450 893.400 95.250 896.400 ;
        RECT 101.250 894.300 103.050 896.400 ;
        RECT 101.250 893.400 105.000 894.300 ;
        RECT 85.650 892.500 86.700 893.400 ;
        RECT 82.950 891.300 86.700 892.500 ;
        RECT 94.200 892.500 95.250 893.400 ;
        RECT 103.950 892.500 105.000 893.400 ;
        RECT 94.200 891.450 99.150 892.500 ;
        RECT 82.950 890.400 85.050 891.300 ;
        RECT 97.350 890.700 99.150 891.450 ;
        RECT 77.550 883.050 78.750 890.400 ;
        RECT 100.650 889.800 102.450 891.600 ;
        RECT 103.950 890.400 106.050 892.500 ;
        RECT 109.050 890.400 110.850 896.400 ;
        RECT 90.150 888.000 91.950 888.600 ;
        RECT 101.100 888.000 102.150 889.800 ;
        RECT 90.150 886.800 102.150 888.000 ;
        RECT 77.550 881.250 83.850 883.050 ;
        RECT 77.550 880.950 82.050 881.250 ;
        RECT 77.550 873.600 78.750 880.950 ;
        RECT 79.950 875.400 81.750 877.200 ;
        RECT 80.850 874.200 85.050 875.400 ;
        RECT 90.150 874.200 91.050 886.800 ;
        RECT 101.100 885.600 108.000 886.800 ;
        RECT 101.100 885.000 102.900 885.600 ;
        RECT 107.100 884.850 108.000 885.600 ;
        RECT 104.100 883.800 105.900 884.400 ;
        RECT 97.950 882.600 105.900 883.800 ;
        RECT 107.100 883.050 108.900 884.850 ;
        RECT 97.950 880.950 100.050 882.600 ;
        RECT 106.950 880.950 109.050 883.050 ;
        RECT 99.750 875.700 101.550 876.000 ;
        RECT 109.950 875.700 110.850 890.400 ;
        RECT 125.400 889.500 127.200 896.400 ;
        RECT 131.400 889.500 133.200 896.400 ;
        RECT 137.400 889.500 139.200 896.400 ;
        RECT 143.400 889.500 145.200 896.400 ;
        RECT 161.400 890.400 163.200 896.400 ;
        RECT 168.600 891.000 170.400 896.400 ;
        RECT 161.400 889.500 162.900 890.400 ;
        RECT 125.400 888.300 129.300 889.500 ;
        RECT 131.400 888.300 135.300 889.500 ;
        RECT 137.400 888.300 141.300 889.500 ;
        RECT 143.400 888.300 146.100 889.500 ;
        RECT 128.100 887.400 129.300 888.300 ;
        RECT 134.100 887.400 135.300 888.300 ;
        RECT 140.100 887.400 141.300 888.300 ;
        RECT 128.100 886.200 132.300 887.400 ;
        RECT 125.100 883.050 126.900 884.850 ;
        RECT 124.950 880.950 127.050 883.050 ;
        RECT 128.100 875.700 129.300 886.200 ;
        RECT 130.500 885.600 132.300 886.200 ;
        RECT 134.100 886.200 138.300 887.400 ;
        RECT 134.100 875.700 135.300 886.200 ;
        RECT 136.500 885.600 138.300 886.200 ;
        RECT 140.100 886.200 144.300 887.400 ;
        RECT 140.100 875.700 141.300 886.200 ;
        RECT 142.500 885.600 144.300 886.200 ;
        RECT 145.200 883.050 146.100 888.300 ;
        RECT 161.400 888.000 165.750 889.500 ;
        RECT 163.650 887.400 165.750 888.000 ;
        RECT 169.350 888.900 170.400 891.000 ;
        RECT 176.400 890.400 178.200 896.400 ;
        RECT 173.700 889.200 178.200 890.400 ;
        RECT 194.400 889.200 196.200 896.400 ;
        RECT 215.400 889.200 217.200 896.400 ;
        RECT 243.000 890.400 244.800 896.400 ;
        RECT 166.650 885.900 168.450 887.700 ;
        RECT 169.350 886.800 172.500 888.900 ;
        RECT 173.700 887.100 175.800 889.200 ;
        RECT 194.400 888.300 198.600 889.200 ;
        RECT 215.400 888.300 219.600 889.200 ;
        RECT 166.200 885.000 168.300 885.900 ;
        RECT 161.700 883.800 168.300 885.000 ;
        RECT 161.700 883.200 163.500 883.800 ;
        RECT 145.200 880.950 148.050 883.050 ;
        RECT 161.400 881.100 163.500 883.200 ;
        RECT 145.200 875.700 146.100 880.950 ;
        RECT 166.200 880.800 168.300 882.900 ;
        RECT 166.200 879.000 168.000 880.800 ;
        RECT 169.350 880.200 170.250 886.800 ;
        RECT 171.150 882.900 173.250 885.000 ;
        RECT 171.300 881.100 173.100 882.900 ;
        RECT 175.950 881.100 178.050 883.200 ;
        RECT 194.100 883.050 195.900 884.850 ;
        RECT 197.400 883.050 198.600 888.300 ;
        RECT 200.100 883.050 201.900 884.850 ;
        RECT 215.100 883.050 216.900 884.850 ;
        RECT 218.400 883.050 219.600 888.300 ;
        RECT 221.100 883.050 222.900 884.850 ;
        RECT 236.100 883.050 237.900 884.850 ;
        RECT 243.000 883.050 244.050 890.400 ;
        RECT 265.200 888.000 267.000 896.400 ;
        RECT 286.800 893.400 288.600 896.400 ;
        RECT 263.700 886.800 267.000 888.000 ;
        RECT 248.100 883.050 249.900 884.850 ;
        RECT 263.700 883.050 264.600 886.800 ;
        RECT 266.100 883.050 267.900 884.850 ;
        RECT 272.100 883.050 273.900 884.850 ;
        RECT 287.400 883.050 288.600 893.400 ;
        RECT 307.200 888.000 309.000 896.400 ;
        RECT 328.800 893.400 330.600 896.400 ;
        RECT 350.400 893.400 352.200 896.400 ;
        RECT 305.700 886.800 309.000 888.000 ;
        RECT 305.700 883.050 306.600 886.800 ;
        RECT 308.100 883.050 309.900 884.850 ;
        RECT 314.100 883.050 315.900 884.850 ;
        RECT 329.400 883.050 330.600 893.400 ;
        RECT 350.700 883.050 351.600 893.400 ;
        RECT 368.400 891.300 370.200 896.400 ;
        RECT 374.400 891.300 376.200 896.400 ;
        RECT 368.400 889.950 376.200 891.300 ;
        RECT 377.400 890.400 379.200 896.400 ;
        RECT 377.400 888.300 378.600 890.400 ;
        RECT 374.850 887.250 378.600 888.300 ;
        RECT 397.200 888.000 399.000 896.400 ;
        RECT 371.100 883.050 372.900 884.850 ;
        RECT 374.850 883.050 376.050 887.250 ;
        RECT 395.700 886.800 399.000 888.000 ;
        RECT 419.400 893.400 421.200 896.400 ;
        RECT 377.100 883.050 378.900 884.850 ;
        RECT 395.700 883.050 396.600 886.800 ;
        RECT 398.100 883.050 399.900 884.850 ;
        RECT 404.100 883.050 405.900 884.850 ;
        RECT 419.400 883.050 420.600 893.400 ;
        RECT 442.200 888.000 444.000 896.400 ;
        RECT 466.500 891.600 468.300 896.400 ;
        RECT 466.500 890.400 471.600 891.600 ;
        RECT 440.700 886.800 444.000 888.000 ;
        RECT 440.700 883.050 441.600 886.800 ;
        RECT 443.100 883.050 444.900 884.850 ;
        RECT 449.100 883.050 450.900 884.850 ;
        RECT 461.100 883.050 462.900 884.850 ;
        RECT 467.100 883.050 468.900 884.850 ;
        RECT 470.700 883.050 471.600 890.400 ;
        RECT 485.400 891.300 487.200 896.400 ;
        RECT 491.400 891.300 493.200 896.400 ;
        RECT 485.400 889.950 493.200 891.300 ;
        RECT 494.400 890.400 496.200 896.400 ;
        RECT 512.400 893.400 514.200 896.400 ;
        RECT 494.400 888.300 495.600 890.400 ;
        RECT 491.850 887.250 495.600 888.300 ;
        RECT 488.100 883.050 489.900 884.850 ;
        RECT 491.850 883.050 493.050 887.250 ;
        RECT 494.100 883.050 495.900 884.850 ;
        RECT 512.400 883.050 513.600 893.400 ;
        RECT 532.500 891.600 534.300 896.400 ;
        RECT 532.500 890.400 537.600 891.600 ;
        RECT 527.100 883.050 528.900 884.850 ;
        RECT 533.100 883.050 534.900 884.850 ;
        RECT 536.700 883.050 537.600 890.400 ;
        RECT 553.800 890.400 555.600 896.400 ;
        RECT 561.600 891.000 563.400 896.400 ;
        RECT 553.800 889.200 558.300 890.400 ;
        RECT 556.200 887.100 558.300 889.200 ;
        RECT 561.600 888.900 562.650 891.000 ;
        RECT 568.800 890.400 570.600 896.400 ;
        RECT 569.100 889.500 570.600 890.400 ;
        RECT 581.400 891.300 583.200 896.400 ;
        RECT 587.400 891.300 589.200 896.400 ;
        RECT 581.400 889.950 589.200 891.300 ;
        RECT 590.400 890.400 592.200 896.400 ;
        RECT 559.500 886.800 562.650 888.900 ;
        RECT 566.250 888.000 570.600 889.500 ;
        RECT 590.400 888.300 591.600 890.400 ;
        RECT 169.350 878.700 172.500 880.200 ;
        RECT 176.100 879.450 177.900 881.100 ;
        RECT 193.950 880.950 196.050 883.050 ;
        RECT 196.950 880.950 199.050 883.050 ;
        RECT 199.950 880.950 202.050 883.050 ;
        RECT 214.950 880.950 217.050 883.050 ;
        RECT 217.950 880.950 220.050 883.050 ;
        RECT 220.950 880.950 223.050 883.050 ;
        RECT 235.950 880.950 238.050 883.050 ;
        RECT 238.950 880.950 241.050 883.050 ;
        RECT 241.950 880.950 244.050 883.050 ;
        RECT 244.950 880.950 247.050 883.050 ;
        RECT 247.950 880.950 250.050 883.050 ;
        RECT 262.950 880.950 265.050 883.050 ;
        RECT 265.950 880.950 268.050 883.050 ;
        RECT 268.950 880.950 271.050 883.050 ;
        RECT 271.950 880.950 274.050 883.050 ;
        RECT 286.950 880.950 289.050 883.050 ;
        RECT 289.950 880.950 292.050 883.050 ;
        RECT 304.950 880.950 307.050 883.050 ;
        RECT 307.950 880.950 310.050 883.050 ;
        RECT 310.950 880.950 313.050 883.050 ;
        RECT 313.950 880.950 316.050 883.050 ;
        RECT 328.950 880.950 331.050 883.050 ;
        RECT 331.950 880.950 334.050 883.050 ;
        RECT 346.950 880.950 349.050 883.050 ;
        RECT 349.950 880.950 352.050 883.050 ;
        RECT 352.950 880.950 355.050 883.050 ;
        RECT 367.950 880.950 370.050 883.050 ;
        RECT 370.950 880.950 373.050 883.050 ;
        RECT 373.950 880.950 376.050 883.050 ;
        RECT 376.950 880.950 379.050 883.050 ;
        RECT 394.950 880.950 397.050 883.050 ;
        RECT 397.950 880.950 400.050 883.050 ;
        RECT 400.950 880.950 403.050 883.050 ;
        RECT 403.950 880.950 406.050 883.050 ;
        RECT 415.950 880.950 418.050 883.050 ;
        RECT 418.950 880.950 421.050 883.050 ;
        RECT 439.950 880.950 442.050 883.050 ;
        RECT 442.950 880.950 445.050 883.050 ;
        RECT 445.950 880.950 448.050 883.050 ;
        RECT 448.950 880.950 451.050 883.050 ;
        RECT 460.950 880.950 463.050 883.050 ;
        RECT 463.950 880.950 466.050 883.050 ;
        RECT 466.950 880.950 469.050 883.050 ;
        RECT 469.950 880.950 472.050 883.050 ;
        RECT 484.950 880.950 487.050 883.050 ;
        RECT 487.950 880.950 490.050 883.050 ;
        RECT 490.950 880.950 493.050 883.050 ;
        RECT 493.950 880.950 496.050 883.050 ;
        RECT 508.950 880.950 511.050 883.050 ;
        RECT 511.950 880.950 514.050 883.050 ;
        RECT 526.950 880.950 529.050 883.050 ;
        RECT 529.950 880.950 532.050 883.050 ;
        RECT 532.950 880.950 535.050 883.050 ;
        RECT 535.950 880.950 538.050 883.050 ;
        RECT 541.950 882.450 544.050 883.050 ;
        RECT 553.950 882.450 556.050 883.200 ;
        RECT 558.750 882.900 560.850 885.000 ;
        RECT 541.950 881.550 556.050 882.450 ;
        RECT 541.950 880.950 544.050 881.550 ;
        RECT 553.950 881.100 556.050 881.550 ;
        RECT 558.900 881.100 560.700 882.900 ;
        RECT 181.950 879.450 184.050 880.050 ;
        RECT 176.100 879.300 184.050 879.450 ;
        RECT 170.400 878.100 172.500 878.700 ;
        RECT 176.550 878.550 184.050 879.300 ;
        RECT 167.700 875.700 169.500 877.800 ;
        RECT 99.750 875.100 110.850 875.700 ;
        RECT 77.550 861.600 79.350 873.600 ;
        RECT 82.950 873.300 85.050 874.200 ;
        RECT 85.950 873.300 91.050 874.200 ;
        RECT 93.150 874.500 110.850 875.100 ;
        RECT 93.150 874.200 101.550 874.500 ;
        RECT 85.950 872.400 86.850 873.300 ;
        RECT 84.150 870.600 86.850 872.400 ;
        RECT 87.750 872.100 89.550 872.400 ;
        RECT 93.150 872.100 94.050 874.200 ;
        RECT 109.950 873.600 110.850 874.500 ;
        RECT 87.750 871.200 94.050 872.100 ;
        RECT 94.950 872.700 96.750 873.300 ;
        RECT 94.950 871.500 102.450 872.700 ;
        RECT 87.750 870.600 89.550 871.200 ;
        RECT 101.250 870.600 102.450 871.500 ;
        RECT 82.950 867.600 86.850 869.700 ;
        RECT 91.950 869.550 93.750 870.300 ;
        RECT 96.750 869.550 98.550 870.300 ;
        RECT 91.950 868.500 98.550 869.550 ;
        RECT 101.250 868.500 106.050 870.600 ;
        RECT 85.050 861.600 86.850 867.600 ;
        RECT 92.850 861.600 94.650 868.500 ;
        RECT 101.250 867.600 102.450 868.500 ;
        RECT 100.650 861.600 102.450 867.600 ;
        RECT 109.050 861.600 110.850 873.600 ;
        RECT 125.400 874.500 129.300 875.700 ;
        RECT 131.400 874.500 135.300 875.700 ;
        RECT 137.400 874.500 141.300 875.700 ;
        RECT 143.400 874.500 146.100 875.700 ;
        RECT 164.100 874.800 169.500 875.700 ;
        RECT 125.400 861.600 127.200 874.500 ;
        RECT 131.400 861.600 133.200 874.500 ;
        RECT 137.400 861.600 139.200 874.500 ;
        RECT 143.400 861.600 145.200 874.500 ;
        RECT 164.100 873.900 166.200 874.800 ;
        RECT 161.400 872.700 166.200 873.900 ;
        RECT 171.000 873.600 172.200 878.100 ;
        RECT 181.950 877.950 184.050 878.550 ;
        RECT 168.900 872.700 172.200 873.600 ;
        RECT 173.100 873.600 175.200 874.500 ;
        RECT 161.400 861.600 163.200 872.700 ;
        RECT 168.900 861.600 170.700 872.700 ;
        RECT 173.100 872.400 178.200 873.600 ;
        RECT 176.400 861.600 178.200 872.400 ;
        RECT 197.400 867.600 198.600 880.950 ;
        RECT 218.400 867.600 219.600 880.950 ;
        RECT 239.100 879.150 240.900 880.950 ;
        RECT 243.000 875.400 243.900 880.950 ;
        RECT 245.100 879.150 246.900 880.950 ;
        RECT 238.800 874.500 243.900 875.400 ;
        RECT 196.800 861.600 198.600 867.600 ;
        RECT 217.800 861.600 219.600 867.600 ;
        RECT 235.800 862.500 237.600 873.600 ;
        RECT 238.800 863.400 240.600 874.500 ;
        RECT 241.800 872.400 249.600 873.300 ;
        RECT 241.800 862.500 243.600 872.400 ;
        RECT 235.800 861.600 243.600 862.500 ;
        RECT 247.800 861.600 249.600 872.400 ;
        RECT 263.700 868.800 264.600 880.950 ;
        RECT 269.100 879.150 270.900 880.950 ;
        RECT 263.700 867.900 270.300 868.800 ;
        RECT 263.700 867.600 264.600 867.900 ;
        RECT 262.800 861.600 264.600 867.600 ;
        RECT 268.800 867.600 270.300 867.900 ;
        RECT 287.400 867.600 288.600 880.950 ;
        RECT 290.100 879.150 291.900 880.950 ;
        RECT 305.700 868.800 306.600 880.950 ;
        RECT 311.100 879.150 312.900 880.950 ;
        RECT 305.700 867.900 312.300 868.800 ;
        RECT 305.700 867.600 306.600 867.900 ;
        RECT 268.800 861.600 270.600 867.600 ;
        RECT 286.800 861.600 288.600 867.600 ;
        RECT 304.800 861.600 306.600 867.600 ;
        RECT 310.800 867.600 312.300 867.900 ;
        RECT 329.400 867.600 330.600 880.950 ;
        RECT 332.100 879.150 333.900 880.950 ;
        RECT 347.100 879.150 348.900 880.950 ;
        RECT 350.700 873.600 351.600 880.950 ;
        RECT 353.100 879.150 354.900 880.950 ;
        RECT 368.100 879.150 369.900 880.950 ;
        RECT 350.700 872.400 354.300 873.600 ;
        RECT 310.800 861.600 312.600 867.600 ;
        RECT 328.800 861.600 330.600 867.600 ;
        RECT 352.500 861.600 354.300 872.400 ;
        RECT 373.950 867.600 375.150 880.950 ;
        RECT 395.700 868.800 396.600 880.950 ;
        RECT 401.100 879.150 402.900 880.950 ;
        RECT 416.100 879.150 417.900 880.950 ;
        RECT 395.700 867.900 402.300 868.800 ;
        RECT 395.700 867.600 396.600 867.900 ;
        RECT 373.800 861.600 375.600 867.600 ;
        RECT 394.800 861.600 396.600 867.600 ;
        RECT 400.800 867.600 402.300 867.900 ;
        RECT 419.400 867.600 420.600 880.950 ;
        RECT 421.950 879.450 424.050 880.050 ;
        RECT 430.950 879.450 433.050 880.050 ;
        RECT 421.950 878.550 433.050 879.450 ;
        RECT 421.950 877.950 424.050 878.550 ;
        RECT 430.950 877.950 433.050 878.550 ;
        RECT 440.700 868.800 441.600 880.950 ;
        RECT 446.100 879.150 447.900 880.950 ;
        RECT 464.100 879.150 465.900 880.950 ;
        RECT 442.950 876.450 445.050 877.050 ;
        RECT 466.950 876.450 469.050 877.050 ;
        RECT 442.950 875.550 469.050 876.450 ;
        RECT 442.950 874.950 445.050 875.550 ;
        RECT 466.950 874.950 469.050 875.550 ;
        RECT 448.950 873.450 451.050 874.050 ;
        RECT 454.950 873.450 457.050 874.050 ;
        RECT 470.700 873.600 471.600 880.950 ;
        RECT 485.100 879.150 486.900 880.950 ;
        RECT 448.950 872.550 457.050 873.450 ;
        RECT 448.950 871.950 451.050 872.550 ;
        RECT 454.950 871.950 457.050 872.550 ;
        RECT 461.400 872.700 469.200 873.600 ;
        RECT 440.700 867.900 447.300 868.800 ;
        RECT 440.700 867.600 441.600 867.900 ;
        RECT 400.800 861.600 402.600 867.600 ;
        RECT 419.400 861.600 421.200 867.600 ;
        RECT 439.800 861.600 441.600 867.600 ;
        RECT 445.800 867.600 447.300 867.900 ;
        RECT 445.800 861.600 447.600 867.600 ;
        RECT 461.400 861.600 463.200 872.700 ;
        RECT 467.400 861.600 469.200 872.700 ;
        RECT 470.400 861.600 472.200 873.600 ;
        RECT 490.950 867.600 492.150 880.950 ;
        RECT 509.100 879.150 510.900 880.950 ;
        RECT 512.400 867.600 513.600 880.950 ;
        RECT 530.100 879.150 531.900 880.950 ;
        RECT 536.700 873.600 537.600 880.950 ;
        RECT 554.100 879.300 555.900 881.100 ;
        RECT 561.750 880.200 562.650 886.800 ;
        RECT 563.550 885.900 565.350 887.700 ;
        RECT 566.250 887.400 568.350 888.000 ;
        RECT 587.850 887.250 591.600 888.300 ;
        RECT 610.200 888.000 612.000 896.400 ;
        RECT 631.800 890.400 633.600 896.400 ;
        RECT 563.700 885.000 565.800 885.900 ;
        RECT 563.700 883.800 570.300 885.000 ;
        RECT 568.500 883.200 570.300 883.800 ;
        RECT 563.700 880.800 565.800 882.900 ;
        RECT 568.500 881.100 570.600 883.200 ;
        RECT 584.100 883.050 585.900 884.850 ;
        RECT 587.850 883.050 589.050 887.250 ;
        RECT 608.700 886.800 612.000 888.000 ;
        RECT 632.400 888.300 633.600 890.400 ;
        RECT 634.800 891.300 636.600 896.400 ;
        RECT 640.800 891.300 642.600 896.400 ;
        RECT 634.800 889.950 642.600 891.300 ;
        RECT 632.400 887.250 636.150 888.300 ;
        RECT 658.200 888.000 660.000 896.400 ;
        RECT 682.800 889.200 684.600 896.400 ;
        RECT 704.700 891.600 706.500 896.400 ;
        RECT 592.950 885.450 597.000 886.050 ;
        RECT 590.100 883.050 591.900 884.850 ;
        RECT 592.950 883.950 597.450 885.450 ;
        RECT 580.950 880.950 583.050 883.050 ;
        RECT 583.950 880.950 586.050 883.050 ;
        RECT 586.950 880.950 589.050 883.050 ;
        RECT 589.950 880.950 592.050 883.050 ;
        RECT 559.500 878.700 562.650 880.200 ;
        RECT 564.000 879.000 565.800 880.800 ;
        RECT 581.100 879.150 582.900 880.950 ;
        RECT 559.500 878.100 561.600 878.700 ;
        RECT 556.800 873.600 558.900 874.500 ;
        RECT 527.400 872.700 535.200 873.600 ;
        RECT 490.800 861.600 492.600 867.600 ;
        RECT 512.400 861.600 514.200 867.600 ;
        RECT 527.400 861.600 529.200 872.700 ;
        RECT 533.400 861.600 535.200 872.700 ;
        RECT 536.400 861.600 538.200 873.600 ;
        RECT 553.800 872.400 558.900 873.600 ;
        RECT 559.800 873.600 561.000 878.100 ;
        RECT 562.500 875.700 564.300 877.800 ;
        RECT 562.500 874.800 567.900 875.700 ;
        RECT 565.800 873.900 567.900 874.800 ;
        RECT 559.800 872.700 563.100 873.600 ;
        RECT 565.800 872.700 570.600 873.900 ;
        RECT 553.800 861.600 555.600 872.400 ;
        RECT 561.300 861.600 563.100 872.700 ;
        RECT 568.800 861.600 570.600 872.700 ;
        RECT 586.950 867.600 588.150 880.950 ;
        RECT 596.550 880.050 597.450 883.950 ;
        RECT 608.700 883.050 609.600 886.800 ;
        RECT 611.100 883.050 612.900 884.850 ;
        RECT 617.100 883.050 618.900 884.850 ;
        RECT 632.100 883.050 633.900 884.850 ;
        RECT 634.950 883.050 636.150 887.250 ;
        RECT 656.700 886.800 660.000 888.000 ;
        RECT 680.400 888.300 684.600 889.200 ;
        RECT 701.400 890.400 706.500 891.600 ;
        RECT 638.100 883.050 639.900 884.850 ;
        RECT 656.700 883.050 657.600 886.800 ;
        RECT 659.100 883.050 660.900 884.850 ;
        RECT 665.100 883.050 666.900 884.850 ;
        RECT 677.100 883.050 678.900 884.850 ;
        RECT 680.400 883.050 681.600 888.300 ;
        RECT 683.100 883.050 684.900 884.850 ;
        RECT 701.400 883.050 702.300 890.400 ;
        RECT 706.950 888.450 709.050 889.200 ;
        RECT 721.950 888.450 724.050 889.050 ;
        RECT 706.950 887.550 724.050 888.450 ;
        RECT 727.200 888.000 729.000 896.400 ;
        RECT 751.200 888.000 753.000 896.400 ;
        RECT 775.500 891.600 777.300 896.400 ;
        RECT 796.800 893.400 798.600 896.400 ;
        RECT 775.500 890.400 780.600 891.600 ;
        RECT 706.950 887.100 709.050 887.550 ;
        RECT 721.950 886.950 724.050 887.550 ;
        RECT 725.700 886.800 729.000 888.000 ;
        RECT 749.700 886.800 753.000 888.000 ;
        RECT 704.100 883.050 705.900 884.850 ;
        RECT 710.100 883.050 711.900 884.850 ;
        RECT 725.700 883.050 726.600 886.800 ;
        RECT 728.100 883.050 729.900 884.850 ;
        RECT 734.100 883.050 735.900 884.850 ;
        RECT 749.700 883.050 750.600 886.800 ;
        RECT 752.100 883.050 753.900 884.850 ;
        RECT 758.100 883.050 759.900 884.850 ;
        RECT 770.100 883.050 771.900 884.850 ;
        RECT 776.100 883.050 777.900 884.850 ;
        RECT 779.700 883.050 780.600 890.400 ;
        RECT 797.400 883.050 798.600 893.400 ;
        RECT 815.400 893.400 817.200 896.400 ;
        RECT 815.400 883.050 816.600 893.400 ;
        RECT 835.500 891.600 837.300 896.400 ;
        RECT 835.500 890.400 840.600 891.600 ;
        RECT 830.100 883.050 831.900 884.850 ;
        RECT 836.100 883.050 837.900 884.850 ;
        RECT 839.700 883.050 840.600 890.400 ;
        RECT 854.400 891.300 856.200 896.400 ;
        RECT 860.400 891.300 862.200 896.400 ;
        RECT 854.400 889.950 862.200 891.300 ;
        RECT 863.400 890.400 865.200 896.400 ;
        RECT 863.400 888.300 864.600 890.400 ;
        RECT 860.850 887.250 864.600 888.300 ;
        RECT 885.000 888.000 886.800 896.400 ;
        RECT 857.100 883.050 858.900 884.850 ;
        RECT 860.850 883.050 862.050 887.250 ;
        RECT 885.000 886.800 888.300 888.000 ;
        RECT 863.100 883.050 864.900 884.850 ;
        RECT 878.100 883.050 879.900 884.850 ;
        RECT 884.100 883.050 885.900 884.850 ;
        RECT 887.400 883.050 888.300 886.800 ;
        RECT 607.950 880.950 610.050 883.050 ;
        RECT 610.950 880.950 613.050 883.050 ;
        RECT 613.950 880.950 616.050 883.050 ;
        RECT 616.950 880.950 619.050 883.050 ;
        RECT 631.950 880.950 634.050 883.050 ;
        RECT 634.950 880.950 637.050 883.050 ;
        RECT 637.950 880.950 640.050 883.050 ;
        RECT 640.950 880.950 643.050 883.050 ;
        RECT 655.950 880.950 658.050 883.050 ;
        RECT 658.950 880.950 661.050 883.050 ;
        RECT 661.950 880.950 664.050 883.050 ;
        RECT 664.950 880.950 667.050 883.050 ;
        RECT 676.950 880.950 679.050 883.050 ;
        RECT 679.950 880.950 682.050 883.050 ;
        RECT 682.950 880.950 685.050 883.050 ;
        RECT 700.950 880.950 703.050 883.050 ;
        RECT 703.950 880.950 706.050 883.050 ;
        RECT 706.950 880.950 709.050 883.050 ;
        RECT 709.950 880.950 712.050 883.050 ;
        RECT 724.950 880.950 727.050 883.050 ;
        RECT 727.950 880.950 730.050 883.050 ;
        RECT 730.950 880.950 733.050 883.050 ;
        RECT 733.950 880.950 736.050 883.050 ;
        RECT 748.950 880.950 751.050 883.050 ;
        RECT 751.950 880.950 754.050 883.050 ;
        RECT 754.950 880.950 757.050 883.050 ;
        RECT 757.950 880.950 760.050 883.050 ;
        RECT 769.950 880.950 772.050 883.050 ;
        RECT 772.950 880.950 775.050 883.050 ;
        RECT 775.950 880.950 778.050 883.050 ;
        RECT 778.950 880.950 781.050 883.050 ;
        RECT 796.950 880.950 799.050 883.050 ;
        RECT 799.950 880.950 802.050 883.050 ;
        RECT 811.950 880.950 814.050 883.050 ;
        RECT 814.950 880.950 817.050 883.050 ;
        RECT 829.950 880.950 832.050 883.050 ;
        RECT 832.950 880.950 835.050 883.050 ;
        RECT 835.950 880.950 838.050 883.050 ;
        RECT 838.950 880.950 841.050 883.050 ;
        RECT 853.950 880.950 856.050 883.050 ;
        RECT 856.950 880.950 859.050 883.050 ;
        RECT 859.950 880.950 862.050 883.050 ;
        RECT 862.950 880.950 865.050 883.050 ;
        RECT 877.950 880.950 880.050 883.050 ;
        RECT 880.950 880.950 883.050 883.050 ;
        RECT 883.950 880.950 886.050 883.050 ;
        RECT 886.950 880.950 889.050 883.050 ;
        RECT 592.950 878.550 597.450 880.050 ;
        RECT 592.950 877.950 597.000 878.550 ;
        RECT 608.700 868.800 609.600 880.950 ;
        RECT 614.100 879.150 615.900 880.950 ;
        RECT 610.950 876.450 613.050 877.050 ;
        RECT 622.950 876.450 625.050 877.050 ;
        RECT 610.950 875.550 625.050 876.450 ;
        RECT 610.950 874.950 613.050 875.550 ;
        RECT 622.950 874.950 625.050 875.550 ;
        RECT 608.700 867.900 615.300 868.800 ;
        RECT 608.700 867.600 609.600 867.900 ;
        RECT 586.800 861.600 588.600 867.600 ;
        RECT 607.800 861.600 609.600 867.600 ;
        RECT 613.800 867.600 615.300 867.900 ;
        RECT 635.850 867.600 637.050 880.950 ;
        RECT 641.100 879.150 642.900 880.950 ;
        RECT 656.700 868.800 657.600 880.950 ;
        RECT 662.100 879.150 663.900 880.950 ;
        RECT 656.700 867.900 663.300 868.800 ;
        RECT 656.700 867.600 657.600 867.900 ;
        RECT 613.800 861.600 615.600 867.600 ;
        RECT 635.400 861.600 637.200 867.600 ;
        RECT 655.800 861.600 657.600 867.600 ;
        RECT 661.800 867.600 663.300 867.900 ;
        RECT 680.400 867.600 681.600 880.950 ;
        RECT 701.400 873.600 702.300 880.950 ;
        RECT 707.100 879.150 708.900 880.950 ;
        RECT 661.800 861.600 663.600 867.600 ;
        RECT 680.400 861.600 682.200 867.600 ;
        RECT 700.800 861.600 702.600 873.600 ;
        RECT 703.800 872.700 711.600 873.600 ;
        RECT 703.800 861.600 705.600 872.700 ;
        RECT 709.800 861.600 711.600 872.700 ;
        RECT 725.700 868.800 726.600 880.950 ;
        RECT 731.100 879.150 732.900 880.950 ;
        RECT 730.950 873.450 733.050 877.050 ;
        RECT 739.950 873.450 742.050 874.050 ;
        RECT 730.950 873.000 742.050 873.450 ;
        RECT 731.550 872.550 742.050 873.000 ;
        RECT 739.950 871.950 742.050 872.550 ;
        RECT 749.700 868.800 750.600 880.950 ;
        RECT 755.100 879.150 756.900 880.950 ;
        RECT 773.100 879.150 774.900 880.950 ;
        RECT 757.950 876.450 760.050 877.050 ;
        RECT 775.950 876.450 778.050 877.050 ;
        RECT 757.950 875.550 778.050 876.450 ;
        RECT 757.950 874.950 760.050 875.550 ;
        RECT 775.950 874.950 778.050 875.550 ;
        RECT 779.700 873.600 780.600 880.950 ;
        RECT 770.400 872.700 778.200 873.600 ;
        RECT 725.700 867.900 732.300 868.800 ;
        RECT 725.700 867.600 726.600 867.900 ;
        RECT 724.800 861.600 726.600 867.600 ;
        RECT 730.800 867.600 732.300 867.900 ;
        RECT 749.700 867.900 756.300 868.800 ;
        RECT 749.700 867.600 750.600 867.900 ;
        RECT 730.800 861.600 732.600 867.600 ;
        RECT 748.800 861.600 750.600 867.600 ;
        RECT 754.800 867.600 756.300 867.900 ;
        RECT 754.800 861.600 756.600 867.600 ;
        RECT 770.400 861.600 772.200 872.700 ;
        RECT 776.400 861.600 778.200 872.700 ;
        RECT 779.400 861.600 781.200 873.600 ;
        RECT 797.400 867.600 798.600 880.950 ;
        RECT 800.100 879.150 801.900 880.950 ;
        RECT 812.100 879.150 813.900 880.950 ;
        RECT 796.800 861.600 798.600 867.600 ;
        RECT 815.400 867.600 816.600 880.950 ;
        RECT 833.100 879.150 834.900 880.950 ;
        RECT 839.700 873.600 840.600 880.950 ;
        RECT 854.100 879.150 855.900 880.950 ;
        RECT 830.400 872.700 838.200 873.600 ;
        RECT 815.400 861.600 817.200 867.600 ;
        RECT 830.400 861.600 832.200 872.700 ;
        RECT 836.400 861.600 838.200 872.700 ;
        RECT 839.400 861.600 841.200 873.600 ;
        RECT 859.950 867.600 861.150 880.950 ;
        RECT 881.100 879.150 882.900 880.950 ;
        RECT 887.400 868.800 888.300 880.950 ;
        RECT 881.700 867.900 888.300 868.800 ;
        RECT 881.700 867.600 883.200 867.900 ;
        RECT 859.800 861.600 861.600 867.600 ;
        RECT 881.400 861.600 883.200 867.600 ;
        RECT 887.400 867.600 888.300 867.900 ;
        RECT 887.400 861.600 889.200 867.600 ;
        RECT 14.400 851.400 16.200 857.400 ;
        RECT 10.950 835.950 13.050 838.050 ;
        RECT 11.100 834.150 12.900 835.950 ;
        RECT 14.400 831.300 15.300 851.400 ;
        RECT 20.400 845.400 22.200 857.400 ;
        RECT 38.400 851.400 40.200 857.400 ;
        RECT 17.100 838.050 18.900 839.850 ;
        RECT 20.700 838.050 21.600 845.400 ;
        RECT 35.100 838.050 36.900 839.850 ;
        RECT 38.400 838.050 39.600 851.400 ;
        RECT 44.550 845.400 46.350 857.400 ;
        RECT 52.050 851.400 53.850 857.400 ;
        RECT 49.950 849.300 53.850 851.400 ;
        RECT 59.850 850.500 61.650 857.400 ;
        RECT 67.650 851.400 69.450 857.400 ;
        RECT 68.250 850.500 69.450 851.400 ;
        RECT 58.950 849.450 65.550 850.500 ;
        RECT 58.950 848.700 60.750 849.450 ;
        RECT 63.750 848.700 65.550 849.450 ;
        RECT 68.250 848.400 73.050 850.500 ;
        RECT 51.150 846.600 53.850 848.400 ;
        RECT 54.750 847.800 56.550 848.400 ;
        RECT 54.750 846.900 61.050 847.800 ;
        RECT 68.250 847.500 69.450 848.400 ;
        RECT 54.750 846.600 56.550 846.900 ;
        RECT 52.950 845.700 53.850 846.600 ;
        RECT 44.550 838.050 45.750 845.400 ;
        RECT 49.950 844.800 52.050 845.700 ;
        RECT 52.950 844.800 58.050 845.700 ;
        RECT 47.850 843.600 52.050 844.800 ;
        RECT 46.950 841.800 48.750 843.600 ;
        RECT 16.950 835.950 19.050 838.050 ;
        RECT 19.950 835.950 22.050 838.050 ;
        RECT 34.950 835.950 37.050 838.050 ;
        RECT 37.950 835.950 40.050 838.050 ;
        RECT 44.550 837.750 49.050 838.050 ;
        RECT 44.550 835.950 50.850 837.750 ;
        RECT 11.400 830.400 18.900 831.300 ;
        RECT 11.400 822.600 13.200 830.400 ;
        RECT 17.100 829.500 18.900 830.400 ;
        RECT 20.700 828.600 21.600 835.950 ;
        RECT 18.900 826.800 21.600 828.600 ;
        RECT 18.900 822.600 20.700 826.800 ;
        RECT 38.400 825.600 39.600 835.950 ;
        RECT 44.550 828.600 45.750 835.950 ;
        RECT 57.150 832.200 58.050 844.800 ;
        RECT 60.150 844.800 61.050 846.900 ;
        RECT 61.950 846.300 69.450 847.500 ;
        RECT 61.950 845.700 63.750 846.300 ;
        RECT 76.050 845.400 77.850 857.400 ;
        RECT 93.900 845.400 97.200 857.400 ;
        RECT 120.900 845.400 124.200 857.400 ;
        RECT 146.400 851.400 148.200 857.400 ;
        RECT 170.400 851.400 172.200 857.400 ;
        RECT 60.150 844.500 68.550 844.800 ;
        RECT 76.950 844.500 77.850 845.400 ;
        RECT 60.150 843.900 77.850 844.500 ;
        RECT 66.750 843.300 77.850 843.900 ;
        RECT 66.750 843.000 68.550 843.300 ;
        RECT 64.950 836.400 67.050 838.050 ;
        RECT 64.950 835.200 72.900 836.400 ;
        RECT 73.950 835.950 76.050 838.050 ;
        RECT 71.100 834.600 72.900 835.200 ;
        RECT 74.100 834.150 75.900 835.950 ;
        RECT 68.100 833.400 69.900 834.000 ;
        RECT 74.100 833.400 75.000 834.150 ;
        RECT 68.100 832.200 75.000 833.400 ;
        RECT 57.150 831.000 69.150 832.200 ;
        RECT 57.150 830.400 58.950 831.000 ;
        RECT 68.100 829.200 69.150 831.000 ;
        RECT 38.400 822.600 40.200 825.600 ;
        RECT 44.550 822.600 46.350 828.600 ;
        RECT 49.950 827.700 52.050 828.600 ;
        RECT 49.950 826.500 53.700 827.700 ;
        RECT 64.350 827.550 66.150 828.300 ;
        RECT 52.650 825.600 53.700 826.500 ;
        RECT 61.200 826.500 66.150 827.550 ;
        RECT 67.650 827.400 69.450 829.200 ;
        RECT 76.950 828.600 77.850 843.300 ;
        RECT 89.100 838.050 90.900 839.850 ;
        RECT 95.100 838.050 96.300 845.400 ;
        RECT 101.100 838.050 102.900 839.850 ;
        RECT 116.100 838.050 117.900 839.850 ;
        RECT 122.100 838.050 123.300 845.400 ;
        RECT 128.100 838.050 129.900 839.850 ;
        RECT 146.400 838.050 147.600 851.400 ;
        RECT 170.400 838.050 171.600 851.400 ;
        RECT 190.800 845.400 192.600 857.400 ;
        RECT 193.800 846.300 195.600 857.400 ;
        RECT 199.800 846.300 201.600 857.400 ;
        RECT 215.400 851.400 217.200 857.400 ;
        RECT 215.700 851.100 217.200 851.400 ;
        RECT 221.400 851.400 223.200 857.400 ;
        RECT 221.400 851.100 222.300 851.400 ;
        RECT 215.700 850.200 222.300 851.100 ;
        RECT 193.800 845.400 201.600 846.300 ;
        RECT 191.400 838.050 192.300 845.400 ;
        RECT 197.100 838.050 198.900 839.850 ;
        RECT 215.100 838.050 216.900 839.850 ;
        RECT 221.400 838.050 222.300 850.200 ;
        RECT 236.400 846.300 238.200 857.400 ;
        RECT 242.400 846.300 244.200 857.400 ;
        RECT 236.400 845.400 244.200 846.300 ;
        RECT 245.400 845.400 247.200 857.400 ;
        RECT 266.400 851.400 268.200 857.400 ;
        RECT 239.100 838.050 240.900 839.850 ;
        RECT 245.700 838.050 246.600 845.400 ;
        RECT 253.950 843.450 256.050 844.050 ;
        RECT 262.950 843.450 265.050 844.050 ;
        RECT 253.950 842.550 265.050 843.450 ;
        RECT 253.950 841.950 256.050 842.550 ;
        RECT 262.950 841.950 265.050 842.550 ;
        RECT 266.850 838.050 268.050 851.400 ;
        RECT 286.800 845.400 288.600 857.400 ;
        RECT 289.800 846.300 291.600 857.400 ;
        RECT 295.800 846.300 297.600 857.400 ;
        RECT 289.800 845.400 297.600 846.300 ;
        RECT 308.400 846.300 310.200 857.400 ;
        RECT 314.400 846.300 316.200 857.400 ;
        RECT 308.400 845.400 316.200 846.300 ;
        RECT 317.400 845.400 319.200 857.400 ;
        RECT 338.400 851.400 340.200 857.400 ;
        RECT 272.100 838.050 273.900 839.850 ;
        RECT 287.400 838.050 288.300 845.400 ;
        RECT 293.100 838.050 294.900 839.850 ;
        RECT 311.100 838.050 312.900 839.850 ;
        RECT 317.700 838.050 318.600 845.400 ;
        RECT 338.850 838.050 340.050 851.400 ;
        RECT 358.800 845.400 360.600 857.400 ;
        RECT 361.800 846.300 363.600 857.400 ;
        RECT 367.800 846.300 369.600 857.400 ;
        RECT 383.400 851.400 385.200 857.400 ;
        RECT 383.700 851.100 385.200 851.400 ;
        RECT 389.400 851.400 391.200 857.400 ;
        RECT 409.800 851.400 411.600 857.400 ;
        RECT 430.800 851.400 432.600 857.400 ;
        RECT 389.400 851.100 390.300 851.400 ;
        RECT 383.700 850.200 390.300 851.100 ;
        RECT 361.800 845.400 369.600 846.300 ;
        RECT 344.100 838.050 345.900 839.850 ;
        RECT 359.400 838.050 360.300 845.400 ;
        RECT 361.950 843.450 364.050 844.050 ;
        RECT 373.950 843.450 376.050 844.050 ;
        RECT 379.950 843.450 382.050 844.050 ;
        RECT 361.950 842.550 382.050 843.450 ;
        RECT 361.950 841.950 364.050 842.550 ;
        RECT 373.950 841.950 376.050 842.550 ;
        RECT 379.950 841.950 382.050 842.550 ;
        RECT 365.100 838.050 366.900 839.850 ;
        RECT 383.100 838.050 384.900 839.850 ;
        RECT 389.400 838.050 390.300 850.200 ;
        RECT 404.100 838.050 405.900 839.850 ;
        RECT 409.950 838.050 411.150 851.400 ;
        RECT 431.700 851.100 432.600 851.400 ;
        RECT 436.800 851.400 438.600 857.400 ;
        RECT 454.800 851.400 456.600 857.400 ;
        RECT 436.800 851.100 438.300 851.400 ;
        RECT 431.700 850.200 438.300 851.100 ;
        RECT 455.700 851.100 456.600 851.400 ;
        RECT 460.800 851.400 462.600 857.400 ;
        RECT 482.400 851.400 484.200 857.400 ;
        RECT 505.800 851.400 507.600 857.400 ;
        RECT 460.800 851.100 462.300 851.400 ;
        RECT 455.700 850.200 462.300 851.100 ;
        RECT 431.700 838.050 432.600 850.200 ;
        RECT 437.100 838.050 438.900 839.850 ;
        RECT 455.700 838.050 456.600 850.200 ;
        RECT 461.100 838.050 462.900 839.850 ;
        RECT 482.850 838.050 484.050 851.400 ;
        RECT 488.100 838.050 489.900 839.850 ;
        RECT 500.100 838.050 501.900 839.850 ;
        RECT 505.950 838.050 507.150 851.400 ;
        RECT 526.800 845.400 528.600 857.400 ;
        RECT 529.800 846.300 531.600 857.400 ;
        RECT 535.800 846.300 537.600 857.400 ;
        RECT 550.800 851.400 552.600 857.400 ;
        RECT 529.800 845.400 537.600 846.300 ;
        RECT 551.700 851.100 552.600 851.400 ;
        RECT 556.800 851.400 558.600 857.400 ;
        RECT 556.800 851.100 558.300 851.400 ;
        RECT 551.700 850.200 558.300 851.100 ;
        RECT 527.400 838.050 528.300 845.400 ;
        RECT 533.100 838.050 534.900 839.850 ;
        RECT 551.700 838.050 552.600 850.200 ;
        RECT 574.800 846.600 576.600 857.400 ;
        RECT 574.800 845.400 579.600 846.600 ;
        RECT 577.500 844.500 579.600 845.400 ;
        RECT 582.300 845.400 584.100 857.400 ;
        RECT 589.800 846.300 591.600 857.400 ;
        RECT 605.400 851.400 607.200 857.400 ;
        RECT 605.700 851.100 607.200 851.400 ;
        RECT 611.400 851.400 613.200 857.400 ;
        RECT 631.800 851.400 633.600 857.400 ;
        RECT 655.800 851.400 657.600 857.400 ;
        RECT 676.800 851.400 678.600 857.400 ;
        RECT 611.400 851.100 612.300 851.400 ;
        RECT 605.700 850.200 612.300 851.100 ;
        RECT 587.100 845.400 591.600 846.300 ;
        RECT 582.300 843.900 583.500 845.400 ;
        RECT 582.000 843.000 583.500 843.900 ;
        RECT 587.100 843.300 589.200 845.400 ;
        RECT 582.000 840.900 582.900 843.000 ;
        RECT 557.100 838.050 558.900 839.850 ;
        RECT 575.100 838.050 576.900 839.850 ;
        RECT 580.800 838.800 582.900 840.900 ;
        RECT 583.800 841.500 585.900 841.800 ;
        RECT 583.800 839.700 587.700 841.500 ;
        RECT 88.950 835.950 91.050 838.050 ;
        RECT 91.950 835.950 94.050 838.050 ;
        RECT 94.950 835.950 97.050 838.050 ;
        RECT 97.950 835.950 100.050 838.050 ;
        RECT 100.950 835.950 103.050 838.050 ;
        RECT 115.950 835.950 118.050 838.050 ;
        RECT 118.950 835.950 121.050 838.050 ;
        RECT 121.950 835.950 124.050 838.050 ;
        RECT 124.950 835.950 127.050 838.050 ;
        RECT 127.950 835.950 130.050 838.050 ;
        RECT 142.950 835.950 145.050 838.050 ;
        RECT 145.950 835.950 148.050 838.050 ;
        RECT 148.950 835.950 151.050 838.050 ;
        RECT 166.950 835.950 169.050 838.050 ;
        RECT 169.950 835.950 172.050 838.050 ;
        RECT 172.950 835.950 175.050 838.050 ;
        RECT 190.950 835.950 193.050 838.050 ;
        RECT 193.950 835.950 196.050 838.050 ;
        RECT 196.950 835.950 199.050 838.050 ;
        RECT 199.950 835.950 202.050 838.050 ;
        RECT 211.950 835.950 214.050 838.050 ;
        RECT 214.950 835.950 217.050 838.050 ;
        RECT 217.950 835.950 220.050 838.050 ;
        RECT 220.950 835.950 223.050 838.050 ;
        RECT 235.950 835.950 238.050 838.050 ;
        RECT 238.950 835.950 241.050 838.050 ;
        RECT 241.950 835.950 244.050 838.050 ;
        RECT 244.950 835.950 247.050 838.050 ;
        RECT 262.950 835.950 265.050 838.050 ;
        RECT 265.950 835.950 268.050 838.050 ;
        RECT 268.950 835.950 271.050 838.050 ;
        RECT 271.950 835.950 274.050 838.050 ;
        RECT 286.950 835.950 289.050 838.050 ;
        RECT 289.950 835.950 292.050 838.050 ;
        RECT 292.950 835.950 295.050 838.050 ;
        RECT 295.950 835.950 298.050 838.050 ;
        RECT 307.950 835.950 310.050 838.050 ;
        RECT 310.950 835.950 313.050 838.050 ;
        RECT 313.950 835.950 316.050 838.050 ;
        RECT 316.950 835.950 319.050 838.050 ;
        RECT 334.950 835.950 337.050 838.050 ;
        RECT 337.950 835.950 340.050 838.050 ;
        RECT 340.950 835.950 343.050 838.050 ;
        RECT 343.950 835.950 346.050 838.050 ;
        RECT 358.950 835.950 361.050 838.050 ;
        RECT 361.950 835.950 364.050 838.050 ;
        RECT 364.950 835.950 367.050 838.050 ;
        RECT 367.950 835.950 370.050 838.050 ;
        RECT 379.950 835.950 382.050 838.050 ;
        RECT 382.950 835.950 385.050 838.050 ;
        RECT 385.950 835.950 388.050 838.050 ;
        RECT 388.950 835.950 391.050 838.050 ;
        RECT 403.950 835.950 406.050 838.050 ;
        RECT 406.950 835.950 409.050 838.050 ;
        RECT 409.950 835.950 412.050 838.050 ;
        RECT 412.950 835.950 415.050 838.050 ;
        RECT 430.950 835.950 433.050 838.050 ;
        RECT 433.950 835.950 436.050 838.050 ;
        RECT 436.950 835.950 439.050 838.050 ;
        RECT 439.950 835.950 442.050 838.050 ;
        RECT 454.950 835.950 457.050 838.050 ;
        RECT 457.950 835.950 460.050 838.050 ;
        RECT 460.950 835.950 463.050 838.050 ;
        RECT 463.950 835.950 466.050 838.050 ;
        RECT 478.950 835.950 481.050 838.050 ;
        RECT 481.950 835.950 484.050 838.050 ;
        RECT 484.950 835.950 487.050 838.050 ;
        RECT 487.950 835.950 490.050 838.050 ;
        RECT 499.950 835.950 502.050 838.050 ;
        RECT 502.950 835.950 505.050 838.050 ;
        RECT 505.950 835.950 508.050 838.050 ;
        RECT 508.950 835.950 511.050 838.050 ;
        RECT 526.950 835.950 529.050 838.050 ;
        RECT 529.950 835.950 532.050 838.050 ;
        RECT 532.950 835.950 535.050 838.050 ;
        RECT 535.950 835.950 538.050 838.050 ;
        RECT 550.950 835.950 553.050 838.050 ;
        RECT 553.950 835.950 556.050 838.050 ;
        RECT 556.950 835.950 559.050 838.050 ;
        RECT 559.950 835.950 562.050 838.050 ;
        RECT 565.950 837.450 568.050 838.050 ;
        RECT 574.950 837.450 577.050 838.050 ;
        RECT 581.400 837.900 583.800 838.800 ;
        RECT 565.950 836.550 577.050 837.450 ;
        RECT 565.950 835.950 568.050 836.550 ;
        RECT 574.950 835.950 577.050 836.550 ;
        RECT 92.100 834.150 93.900 835.950 ;
        RECT 94.950 831.300 96.300 835.950 ;
        RECT 98.100 834.150 99.900 835.950 ;
        RECT 119.100 834.150 120.900 835.950 ;
        RECT 121.950 831.300 123.300 835.950 ;
        RECT 125.100 834.150 126.900 835.950 ;
        RECT 143.100 834.150 144.900 835.950 ;
        RECT 94.950 830.100 99.600 831.300 ;
        RECT 121.950 830.100 126.600 831.300 ;
        RECT 70.950 826.500 73.050 828.600 ;
        RECT 61.200 825.600 62.250 826.500 ;
        RECT 70.950 825.600 72.000 826.500 ;
        RECT 52.650 822.600 54.450 825.600 ;
        RECT 60.450 822.600 62.250 825.600 ;
        RECT 68.250 824.700 72.000 825.600 ;
        RECT 68.250 822.600 70.050 824.700 ;
        RECT 76.050 822.600 77.850 828.600 ;
        RECT 89.400 828.000 97.200 828.900 ;
        RECT 98.700 828.600 99.600 830.100 ;
        RECT 89.400 822.600 91.200 828.000 ;
        RECT 95.400 823.500 97.200 828.000 ;
        RECT 98.400 824.400 100.200 828.600 ;
        RECT 101.400 823.500 103.200 828.600 ;
        RECT 95.400 822.600 103.200 823.500 ;
        RECT 116.400 828.000 124.200 828.900 ;
        RECT 125.700 828.600 126.600 830.100 ;
        RECT 146.400 830.700 147.600 835.950 ;
        RECT 149.100 834.150 150.900 835.950 ;
        RECT 167.100 834.150 168.900 835.950 ;
        RECT 170.400 830.700 171.600 835.950 ;
        RECT 173.100 834.150 174.900 835.950 ;
        RECT 146.400 829.800 150.600 830.700 ;
        RECT 170.400 829.800 174.600 830.700 ;
        RECT 116.400 822.600 118.200 828.000 ;
        RECT 122.400 823.500 124.200 828.000 ;
        RECT 125.400 824.400 127.200 828.600 ;
        RECT 128.400 823.500 130.200 828.600 ;
        RECT 122.400 822.600 130.200 823.500 ;
        RECT 148.800 822.600 150.600 829.800 ;
        RECT 172.800 822.600 174.600 829.800 ;
        RECT 191.400 828.600 192.300 835.950 ;
        RECT 194.100 834.150 195.900 835.950 ;
        RECT 200.100 834.150 201.900 835.950 ;
        RECT 212.100 834.150 213.900 835.950 ;
        RECT 218.100 834.150 219.900 835.950 ;
        RECT 221.400 832.200 222.300 835.950 ;
        RECT 236.100 834.150 237.900 835.950 ;
        RECT 242.100 834.150 243.900 835.950 ;
        RECT 219.000 831.000 222.300 832.200 ;
        RECT 191.400 827.400 196.500 828.600 ;
        RECT 194.700 822.600 196.500 827.400 ;
        RECT 219.000 822.600 220.800 831.000 ;
        RECT 245.700 828.600 246.600 835.950 ;
        RECT 263.100 834.150 264.900 835.950 ;
        RECT 265.950 831.750 267.150 835.950 ;
        RECT 269.100 834.150 270.900 835.950 ;
        RECT 263.400 830.700 267.150 831.750 ;
        RECT 263.400 828.600 264.600 830.700 ;
        RECT 241.500 827.400 246.600 828.600 ;
        RECT 241.500 822.600 243.300 827.400 ;
        RECT 262.800 822.600 264.600 828.600 ;
        RECT 265.800 827.700 273.600 829.050 ;
        RECT 265.800 822.600 267.600 827.700 ;
        RECT 271.800 822.600 273.600 827.700 ;
        RECT 287.400 828.600 288.300 835.950 ;
        RECT 290.100 834.150 291.900 835.950 ;
        RECT 296.100 834.150 297.900 835.950 ;
        RECT 308.100 834.150 309.900 835.950 ;
        RECT 314.100 834.150 315.900 835.950 ;
        RECT 317.700 828.600 318.600 835.950 ;
        RECT 335.100 834.150 336.900 835.950 ;
        RECT 337.950 831.750 339.150 835.950 ;
        RECT 341.100 834.150 342.900 835.950 ;
        RECT 335.400 830.700 339.150 831.750 ;
        RECT 335.400 828.600 336.600 830.700 ;
        RECT 287.400 827.400 292.500 828.600 ;
        RECT 290.700 822.600 292.500 827.400 ;
        RECT 313.500 827.400 318.600 828.600 ;
        RECT 313.500 822.600 315.300 827.400 ;
        RECT 334.800 822.600 336.600 828.600 ;
        RECT 337.800 827.700 345.600 829.050 ;
        RECT 337.800 822.600 339.600 827.700 ;
        RECT 343.800 822.600 345.600 827.700 ;
        RECT 359.400 828.600 360.300 835.950 ;
        RECT 362.100 834.150 363.900 835.950 ;
        RECT 368.100 834.150 369.900 835.950 ;
        RECT 380.100 834.150 381.900 835.950 ;
        RECT 386.100 834.150 387.900 835.950 ;
        RECT 389.400 832.200 390.300 835.950 ;
        RECT 407.100 834.150 408.900 835.950 ;
        RECT 364.950 831.450 367.050 832.050 ;
        RECT 370.950 831.450 373.050 832.050 ;
        RECT 364.950 830.550 373.050 831.450 ;
        RECT 364.950 829.950 367.050 830.550 ;
        RECT 370.950 829.950 373.050 830.550 ;
        RECT 387.000 831.000 390.300 832.200 ;
        RECT 410.850 831.750 412.050 835.950 ;
        RECT 413.100 834.150 414.900 835.950 ;
        RECT 431.700 832.200 432.600 835.950 ;
        RECT 434.100 834.150 435.900 835.950 ;
        RECT 440.100 834.150 441.900 835.950 ;
        RECT 451.950 834.450 454.050 835.050 ;
        RECT 443.550 834.000 454.050 834.450 ;
        RECT 442.950 833.550 454.050 834.000 ;
        RECT 359.400 827.400 364.500 828.600 ;
        RECT 362.700 822.600 364.500 827.400 ;
        RECT 387.000 822.600 388.800 831.000 ;
        RECT 410.850 830.700 414.600 831.750 ;
        RECT 431.700 831.000 435.000 832.200 ;
        RECT 404.400 827.700 412.200 829.050 ;
        RECT 404.400 822.600 406.200 827.700 ;
        RECT 410.400 822.600 412.200 827.700 ;
        RECT 413.400 828.600 414.600 830.700 ;
        RECT 413.400 822.600 415.200 828.600 ;
        RECT 433.200 822.600 435.000 831.000 ;
        RECT 442.950 829.950 445.050 833.550 ;
        RECT 451.950 832.950 454.050 833.550 ;
        RECT 455.700 832.200 456.600 835.950 ;
        RECT 458.100 834.150 459.900 835.950 ;
        RECT 464.100 834.150 465.900 835.950 ;
        RECT 479.100 834.150 480.900 835.950 ;
        RECT 455.700 831.000 459.000 832.200 ;
        RECT 481.950 831.750 483.150 835.950 ;
        RECT 485.100 834.150 486.900 835.950 ;
        RECT 503.100 834.150 504.900 835.950 ;
        RECT 457.200 822.600 459.000 831.000 ;
        RECT 479.400 830.700 483.150 831.750 ;
        RECT 506.850 831.750 508.050 835.950 ;
        RECT 509.100 834.150 510.900 835.950 ;
        RECT 506.850 830.700 510.600 831.750 ;
        RECT 511.950 831.450 514.050 835.050 ;
        RECT 520.950 831.450 523.050 832.050 ;
        RECT 511.950 831.000 523.050 831.450 ;
        RECT 479.400 828.600 480.600 830.700 ;
        RECT 478.800 822.600 480.600 828.600 ;
        RECT 481.800 827.700 489.600 829.050 ;
        RECT 481.800 822.600 483.600 827.700 ;
        RECT 487.800 822.600 489.600 827.700 ;
        RECT 500.400 827.700 508.200 829.050 ;
        RECT 500.400 822.600 502.200 827.700 ;
        RECT 506.400 822.600 508.200 827.700 ;
        RECT 509.400 828.600 510.600 830.700 ;
        RECT 512.550 830.550 523.050 831.000 ;
        RECT 520.950 829.950 523.050 830.550 ;
        RECT 527.400 828.600 528.300 835.950 ;
        RECT 530.100 834.150 531.900 835.950 ;
        RECT 536.100 834.150 537.900 835.950 ;
        RECT 551.700 832.200 552.600 835.950 ;
        RECT 554.100 834.150 555.900 835.950 ;
        RECT 560.100 834.150 561.900 835.950 ;
        RECT 579.600 835.200 581.400 837.000 ;
        RECT 579.750 833.100 581.850 835.200 ;
        RECT 582.750 832.200 583.800 837.900 ;
        RECT 584.700 837.900 586.500 838.500 ;
        RECT 605.100 838.050 606.900 839.850 ;
        RECT 611.400 838.050 612.300 850.200 ;
        RECT 626.100 838.050 627.900 839.850 ;
        RECT 631.950 838.050 633.150 851.400 ;
        RECT 656.400 838.050 657.600 851.400 ;
        RECT 664.950 843.450 667.050 844.050 ;
        RECT 673.950 843.450 676.050 844.050 ;
        RECT 664.950 842.550 676.050 843.450 ;
        RECT 664.950 841.950 667.050 842.550 ;
        RECT 673.950 841.950 676.050 842.550 ;
        RECT 677.400 838.050 678.600 851.400 ;
        RECT 695.400 851.400 697.200 857.400 ;
        RECT 695.400 838.050 696.600 851.400 ;
        RECT 715.800 845.400 717.600 857.400 ;
        RECT 721.800 851.400 723.600 857.400 ;
        RECT 739.800 851.400 741.600 857.400 ;
        RECT 716.400 838.050 717.300 845.400 ;
        RECT 719.100 838.050 720.900 839.850 ;
        RECT 589.500 837.900 595.050 838.050 ;
        RECT 584.700 836.700 595.050 837.900 ;
        RECT 589.500 835.950 595.050 836.700 ;
        RECT 601.950 835.950 604.050 838.050 ;
        RECT 604.950 835.950 607.050 838.050 ;
        RECT 607.950 835.950 610.050 838.050 ;
        RECT 610.950 835.950 613.050 838.050 ;
        RECT 625.950 835.950 628.050 838.050 ;
        RECT 628.950 835.950 631.050 838.050 ;
        RECT 631.950 835.950 634.050 838.050 ;
        RECT 634.950 835.950 637.050 838.050 ;
        RECT 652.950 835.950 655.050 838.050 ;
        RECT 655.950 835.950 658.050 838.050 ;
        RECT 658.950 835.950 661.050 838.050 ;
        RECT 673.950 835.950 676.050 838.050 ;
        RECT 676.950 835.950 679.050 838.050 ;
        RECT 679.950 835.950 682.050 838.050 ;
        RECT 691.950 835.950 694.050 838.050 ;
        RECT 694.950 835.950 697.050 838.050 ;
        RECT 697.950 835.950 700.050 838.050 ;
        RECT 715.950 835.950 718.050 838.050 ;
        RECT 718.950 835.950 721.050 838.050 ;
        RECT 551.700 831.000 555.000 832.200 ;
        RECT 509.400 822.600 511.200 828.600 ;
        RECT 527.400 827.400 532.500 828.600 ;
        RECT 530.700 822.600 532.500 827.400 ;
        RECT 553.200 822.600 555.000 831.000 ;
        RECT 577.500 829.500 579.600 830.700 ;
        RECT 580.800 830.100 583.800 832.200 ;
        RECT 584.700 833.400 586.500 835.200 ;
        RECT 589.800 834.150 591.600 835.950 ;
        RECT 602.100 834.150 603.900 835.950 ;
        RECT 608.100 834.150 609.900 835.950 ;
        RECT 584.700 831.300 586.800 833.400 ;
        RECT 611.400 832.200 612.300 835.950 ;
        RECT 629.100 834.150 630.900 835.950 ;
        RECT 584.700 830.400 591.000 831.300 ;
        RECT 574.800 828.600 579.600 829.500 ;
        RECT 582.600 828.600 583.800 830.100 ;
        RECT 589.800 828.600 591.000 830.400 ;
        RECT 609.000 831.000 612.300 832.200 ;
        RECT 632.850 831.750 634.050 835.950 ;
        RECT 635.100 834.150 636.900 835.950 ;
        RECT 653.100 834.150 654.900 835.950 ;
        RECT 574.800 822.600 576.600 828.600 ;
        RECT 582.300 822.600 584.100 828.600 ;
        RECT 589.800 822.600 591.600 828.600 ;
        RECT 609.000 822.600 610.800 831.000 ;
        RECT 632.850 830.700 636.600 831.750 ;
        RECT 656.400 830.700 657.600 835.950 ;
        RECT 659.100 834.150 660.900 835.950 ;
        RECT 674.100 834.150 675.900 835.950 ;
        RECT 677.400 830.700 678.600 835.950 ;
        RECT 680.100 834.150 681.900 835.950 ;
        RECT 692.100 834.150 693.900 835.950 ;
        RECT 626.400 827.700 634.200 829.050 ;
        RECT 626.400 822.600 628.200 827.700 ;
        RECT 632.400 822.600 634.200 827.700 ;
        RECT 635.400 828.600 636.600 830.700 ;
        RECT 653.400 829.800 657.600 830.700 ;
        RECT 674.400 829.800 678.600 830.700 ;
        RECT 695.400 830.700 696.600 835.950 ;
        RECT 698.100 834.150 699.900 835.950 ;
        RECT 695.400 829.800 699.600 830.700 ;
        RECT 635.400 822.600 637.200 828.600 ;
        RECT 653.400 822.600 655.200 829.800 ;
        RECT 674.400 822.600 676.200 829.800 ;
        RECT 697.800 822.600 699.600 829.800 ;
        RECT 716.400 828.600 717.300 835.950 ;
        RECT 722.700 831.300 723.600 851.400 ;
        RECT 740.700 851.100 741.600 851.400 ;
        RECT 745.800 851.400 747.600 857.400 ;
        RECT 745.800 851.100 747.300 851.400 ;
        RECT 740.700 850.200 747.300 851.100 ;
        RECT 740.700 838.050 741.600 850.200 ;
        RECT 761.400 846.300 763.200 857.400 ;
        RECT 767.400 846.300 769.200 857.400 ;
        RECT 761.400 845.400 769.200 846.300 ;
        RECT 770.400 845.400 772.200 857.400 ;
        RECT 790.800 851.400 792.600 857.400 ;
        RECT 812.400 851.400 814.200 857.400 ;
        RECT 742.950 843.450 745.050 844.050 ;
        RECT 754.950 843.450 757.050 844.050 ;
        RECT 742.950 842.550 757.050 843.450 ;
        RECT 742.950 841.950 745.050 842.550 ;
        RECT 754.950 841.950 757.050 842.550 ;
        RECT 751.950 840.450 756.000 841.050 ;
        RECT 746.100 838.050 747.900 839.850 ;
        RECT 751.950 838.950 756.450 840.450 ;
        RECT 724.950 835.950 727.050 838.050 ;
        RECT 739.950 835.950 742.050 838.050 ;
        RECT 742.950 835.950 745.050 838.050 ;
        RECT 745.950 835.950 748.050 838.050 ;
        RECT 748.950 835.950 751.050 838.050 ;
        RECT 725.100 834.150 726.900 835.950 ;
        RECT 740.700 832.200 741.600 835.950 ;
        RECT 743.100 834.150 744.900 835.950 ;
        RECT 749.100 834.150 750.900 835.950 ;
        RECT 755.550 835.050 756.450 838.950 ;
        RECT 764.100 838.050 765.900 839.850 ;
        RECT 770.700 838.050 771.600 845.400 ;
        RECT 772.950 840.450 777.000 841.050 ;
        RECT 772.950 838.950 777.450 840.450 ;
        RECT 760.950 835.950 763.050 838.050 ;
        RECT 763.950 835.950 766.050 838.050 ;
        RECT 766.950 835.950 769.050 838.050 ;
        RECT 769.950 835.950 772.050 838.050 ;
        RECT 751.950 833.550 756.450 835.050 ;
        RECT 761.100 834.150 762.900 835.950 ;
        RECT 767.100 834.150 768.900 835.950 ;
        RECT 751.950 832.950 756.000 833.550 ;
        RECT 719.100 830.400 726.600 831.300 ;
        RECT 740.700 831.000 744.000 832.200 ;
        RECT 719.100 829.500 720.900 830.400 ;
        RECT 716.400 826.800 719.100 828.600 ;
        RECT 717.300 822.600 719.100 826.800 ;
        RECT 724.800 822.600 726.600 830.400 ;
        RECT 742.200 822.600 744.000 831.000 ;
        RECT 770.700 828.600 771.600 835.950 ;
        RECT 776.550 831.900 777.450 838.950 ;
        RECT 785.100 838.050 786.900 839.850 ;
        RECT 790.950 838.050 792.150 851.400 ;
        RECT 812.700 851.100 814.200 851.400 ;
        RECT 818.400 851.400 820.200 857.400 ;
        RECT 839.400 851.400 841.200 857.400 ;
        RECT 818.400 851.100 819.300 851.400 ;
        RECT 812.700 850.200 819.300 851.100 ;
        RECT 812.100 838.050 813.900 839.850 ;
        RECT 818.400 838.050 819.300 850.200 ;
        RECT 839.850 838.050 841.050 851.400 ;
        RECT 862.800 845.400 864.600 857.400 ;
        RECT 865.800 846.300 867.600 857.400 ;
        RECT 871.800 846.300 873.600 857.400 ;
        RECT 865.800 845.400 873.600 846.300 ;
        RECT 845.100 838.050 846.900 839.850 ;
        RECT 863.400 838.050 864.300 845.400 ;
        RECT 865.950 843.450 868.050 844.050 ;
        RECT 877.950 843.450 880.050 844.050 ;
        RECT 886.950 843.450 889.050 844.050 ;
        RECT 865.950 842.550 889.050 843.450 ;
        RECT 865.950 841.950 868.050 842.550 ;
        RECT 877.950 841.950 880.050 842.550 ;
        RECT 886.950 841.950 889.050 842.550 ;
        RECT 869.100 838.050 870.900 839.850 ;
        RECT 784.950 835.950 787.050 838.050 ;
        RECT 787.950 835.950 790.050 838.050 ;
        RECT 790.950 835.950 793.050 838.050 ;
        RECT 793.950 835.950 796.050 838.050 ;
        RECT 808.950 835.950 811.050 838.050 ;
        RECT 811.950 835.950 814.050 838.050 ;
        RECT 814.950 835.950 817.050 838.050 ;
        RECT 817.950 835.950 820.050 838.050 ;
        RECT 835.950 835.950 838.050 838.050 ;
        RECT 838.950 835.950 841.050 838.050 ;
        RECT 841.950 835.950 844.050 838.050 ;
        RECT 844.950 835.950 847.050 838.050 ;
        RECT 862.950 835.950 865.050 838.050 ;
        RECT 865.950 835.950 868.050 838.050 ;
        RECT 868.950 835.950 871.050 838.050 ;
        RECT 871.950 835.950 874.050 838.050 ;
        RECT 788.100 834.150 789.900 835.950 ;
        RECT 775.950 829.800 778.050 831.900 ;
        RECT 791.850 831.750 793.050 835.950 ;
        RECT 794.100 834.150 795.900 835.950 ;
        RECT 809.100 834.150 810.900 835.950 ;
        RECT 815.100 834.150 816.900 835.950 ;
        RECT 818.400 832.200 819.300 835.950 ;
        RECT 836.100 834.150 837.900 835.950 ;
        RECT 791.850 830.700 795.600 831.750 ;
        RECT 766.500 827.400 771.600 828.600 ;
        RECT 785.400 827.700 793.200 829.050 ;
        RECT 766.500 822.600 768.300 827.400 ;
        RECT 785.400 822.600 787.200 827.700 ;
        RECT 791.400 822.600 793.200 827.700 ;
        RECT 794.400 828.600 795.600 830.700 ;
        RECT 816.000 831.000 819.300 832.200 ;
        RECT 838.950 831.750 840.150 835.950 ;
        RECT 842.100 834.150 843.900 835.950 ;
        RECT 794.400 822.600 796.200 828.600 ;
        RECT 816.000 822.600 817.800 831.000 ;
        RECT 836.400 830.700 840.150 831.750 ;
        RECT 836.400 828.600 837.600 830.700 ;
        RECT 835.800 822.600 837.600 828.600 ;
        RECT 838.800 827.700 846.600 829.050 ;
        RECT 838.800 822.600 840.600 827.700 ;
        RECT 844.800 822.600 846.600 827.700 ;
        RECT 863.400 828.600 864.300 835.950 ;
        RECT 866.100 834.150 867.900 835.950 ;
        RECT 872.100 834.150 873.900 835.950 ;
        RECT 863.400 827.400 868.500 828.600 ;
        RECT 866.700 822.600 868.500 827.400 ;
        RECT 16.800 811.200 18.600 818.400 ;
        RECT 14.400 810.300 18.600 811.200 ;
        RECT 35.400 815.400 37.200 818.400 ;
        RECT 11.100 805.050 12.900 806.850 ;
        RECT 14.400 805.050 15.600 810.300 ;
        RECT 19.950 807.450 22.050 808.050 ;
        RECT 17.100 805.050 18.900 806.850 ;
        RECT 19.950 806.550 27.450 807.450 ;
        RECT 19.950 805.950 22.050 806.550 ;
        RECT 10.950 802.950 13.050 805.050 ;
        RECT 13.950 802.950 16.050 805.050 ;
        RECT 16.950 802.950 19.050 805.050 ;
        RECT 14.400 789.600 15.600 802.950 ;
        RECT 26.550 802.050 27.450 806.550 ;
        RECT 35.400 805.050 36.600 815.400 ;
        RECT 52.800 812.400 54.600 818.400 ;
        RECT 53.400 810.300 54.600 812.400 ;
        RECT 55.800 813.300 57.600 818.400 ;
        RECT 61.800 813.300 63.600 818.400 ;
        RECT 55.800 811.950 63.600 813.300 ;
        RECT 66.150 812.400 67.950 818.400 ;
        RECT 73.950 816.300 75.750 818.400 ;
        RECT 72.000 815.400 75.750 816.300 ;
        RECT 81.750 815.400 83.550 818.400 ;
        RECT 89.550 815.400 91.350 818.400 ;
        RECT 72.000 814.500 73.050 815.400 ;
        RECT 81.750 814.500 82.800 815.400 ;
        RECT 70.950 812.400 73.050 814.500 ;
        RECT 53.400 809.250 57.150 810.300 ;
        RECT 53.100 805.050 54.900 806.850 ;
        RECT 55.950 805.050 57.150 809.250 ;
        RECT 59.100 805.050 60.900 806.850 ;
        RECT 31.950 802.950 34.050 805.050 ;
        RECT 34.950 802.950 37.050 805.050 ;
        RECT 52.950 802.950 55.050 805.050 ;
        RECT 55.950 802.950 58.050 805.050 ;
        RECT 58.950 802.950 61.050 805.050 ;
        RECT 61.950 802.950 64.050 805.050 ;
        RECT 26.550 800.550 31.050 802.050 ;
        RECT 32.100 801.150 33.900 802.950 ;
        RECT 27.000 799.950 31.050 800.550 ;
        RECT 35.400 789.600 36.600 802.950 ;
        RECT 40.950 798.450 43.050 798.900 ;
        RECT 52.950 798.450 55.050 799.050 ;
        RECT 40.950 797.550 55.050 798.450 ;
        RECT 40.950 796.800 43.050 797.550 ;
        RECT 52.950 796.950 55.050 797.550 ;
        RECT 56.850 789.600 58.050 802.950 ;
        RECT 62.100 801.150 63.900 802.950 ;
        RECT 66.150 797.700 67.050 812.400 ;
        RECT 74.550 811.800 76.350 813.600 ;
        RECT 77.850 813.450 82.800 814.500 ;
        RECT 90.300 814.500 91.350 815.400 ;
        RECT 77.850 812.700 79.650 813.450 ;
        RECT 90.300 813.300 94.050 814.500 ;
        RECT 91.950 812.400 94.050 813.300 ;
        RECT 97.650 812.400 99.450 818.400 ;
        RECT 74.850 810.000 75.900 811.800 ;
        RECT 85.050 810.000 86.850 810.600 ;
        RECT 74.850 808.800 86.850 810.000 ;
        RECT 69.000 807.600 75.900 808.800 ;
        RECT 69.000 806.850 69.900 807.600 ;
        RECT 74.100 807.000 75.900 807.600 ;
        RECT 68.100 805.050 69.900 806.850 ;
        RECT 71.100 805.800 72.900 806.400 ;
        RECT 67.950 802.950 70.050 805.050 ;
        RECT 71.100 804.600 79.050 805.800 ;
        RECT 76.950 802.950 79.050 804.600 ;
        RECT 75.450 797.700 77.250 798.000 ;
        RECT 66.150 797.100 77.250 797.700 ;
        RECT 66.150 796.500 83.850 797.100 ;
        RECT 66.150 795.600 67.050 796.500 ;
        RECT 75.450 796.200 83.850 796.500 ;
        RECT 14.400 783.600 16.200 789.600 ;
        RECT 35.400 783.600 37.200 789.600 ;
        RECT 56.400 783.600 58.200 789.600 ;
        RECT 66.150 783.600 67.950 795.600 ;
        RECT 80.250 794.700 82.050 795.300 ;
        RECT 74.550 793.500 82.050 794.700 ;
        RECT 82.950 794.100 83.850 796.200 ;
        RECT 85.950 796.200 86.850 808.800 ;
        RECT 98.250 805.050 99.450 812.400 ;
        RECT 113.400 815.400 115.200 818.400 ;
        RECT 113.400 805.050 114.600 815.400 ;
        RECT 128.400 813.300 130.200 818.400 ;
        RECT 134.400 813.300 136.200 818.400 ;
        RECT 128.400 811.950 136.200 813.300 ;
        RECT 137.400 812.400 139.200 818.400 ;
        RECT 154.800 815.400 156.600 818.400 ;
        RECT 137.400 810.300 138.600 812.400 ;
        RECT 134.850 809.250 138.600 810.300 ;
        RECT 131.100 805.050 132.900 806.850 ;
        RECT 134.850 805.050 136.050 809.250 ;
        RECT 137.100 805.050 138.900 806.850 ;
        RECT 155.400 805.050 156.600 815.400 ;
        RECT 173.400 811.200 175.200 818.400 ;
        RECT 193.800 815.400 195.600 818.400 ;
        RECT 173.400 810.300 177.600 811.200 ;
        RECT 173.100 805.050 174.900 806.850 ;
        RECT 176.400 805.050 177.600 810.300 ;
        RECT 179.100 805.050 180.900 806.850 ;
        RECT 194.400 805.050 195.600 815.400 ;
        RECT 217.200 810.000 219.000 818.400 ;
        RECT 238.800 815.400 240.600 818.400 ;
        RECT 215.700 808.800 219.000 810.000 ;
        RECT 215.700 805.050 216.600 808.800 ;
        RECT 218.100 805.050 219.900 806.850 ;
        RECT 224.100 805.050 225.900 806.850 ;
        RECT 239.400 805.050 240.600 815.400 ;
        RECT 254.400 813.300 256.200 818.400 ;
        RECT 260.400 813.300 262.200 818.400 ;
        RECT 254.400 811.950 262.200 813.300 ;
        RECT 263.400 812.400 265.200 818.400 ;
        RECT 263.400 810.300 264.600 812.400 ;
        RECT 260.850 809.250 264.600 810.300 ;
        RECT 283.200 810.000 285.000 818.400 ;
        RECT 307.500 813.600 309.300 818.400 ;
        RECT 307.500 812.400 312.600 813.600 ;
        RECT 257.100 805.050 258.900 806.850 ;
        RECT 260.850 805.050 262.050 809.250 ;
        RECT 281.700 808.800 285.000 810.000 ;
        RECT 263.100 805.050 264.900 806.850 ;
        RECT 281.700 805.050 282.600 808.800 ;
        RECT 284.100 805.050 285.900 806.850 ;
        RECT 290.100 805.050 291.900 806.850 ;
        RECT 302.100 805.050 303.900 806.850 ;
        RECT 308.100 805.050 309.900 806.850 ;
        RECT 311.700 805.050 312.600 812.400 ;
        RECT 331.200 810.000 333.000 818.400 ;
        RECT 352.800 815.400 354.600 818.400 ;
        RECT 329.700 808.800 333.000 810.000 ;
        RECT 329.700 805.050 330.600 808.800 ;
        RECT 332.100 805.050 333.900 806.850 ;
        RECT 338.100 805.050 339.900 806.850 ;
        RECT 353.400 805.050 354.600 815.400 ;
        RECT 373.200 810.000 375.000 818.400 ;
        RECT 394.800 812.400 396.600 818.400 ;
        RECT 371.700 808.800 375.000 810.000 ;
        RECT 395.400 810.300 396.600 812.400 ;
        RECT 397.800 813.300 399.600 818.400 ;
        RECT 403.800 813.300 405.600 818.400 ;
        RECT 397.800 811.950 405.600 813.300 ;
        RECT 419.400 811.200 421.200 818.400 ;
        RECT 419.400 810.300 423.600 811.200 ;
        RECT 395.400 809.250 399.150 810.300 ;
        RECT 371.700 805.050 372.600 808.800 ;
        RECT 374.100 805.050 375.900 806.850 ;
        RECT 380.100 805.050 381.900 806.850 ;
        RECT 395.100 805.050 396.900 806.850 ;
        RECT 397.950 805.050 399.150 809.250 ;
        RECT 401.100 805.050 402.900 806.850 ;
        RECT 419.100 805.050 420.900 806.850 ;
        RECT 422.400 805.050 423.600 810.300 ;
        RECT 442.200 810.000 444.000 818.400 ;
        RECT 467.700 813.600 469.500 818.400 ;
        RECT 489.300 814.200 491.100 818.400 ;
        RECT 440.700 808.800 444.000 810.000 ;
        RECT 464.400 812.400 469.500 813.600 ;
        RECT 488.400 812.400 491.100 814.200 ;
        RECT 425.100 805.050 426.900 806.850 ;
        RECT 440.700 805.050 441.600 808.800 ;
        RECT 443.100 805.050 444.900 806.850 ;
        RECT 449.100 805.050 450.900 806.850 ;
        RECT 464.400 805.050 465.300 812.400 ;
        RECT 467.100 805.050 468.900 806.850 ;
        RECT 473.100 805.050 474.900 806.850 ;
        RECT 488.400 805.050 489.300 812.400 ;
        RECT 491.100 810.600 492.900 811.500 ;
        RECT 496.800 810.600 498.600 818.400 ;
        RECT 491.100 809.700 498.600 810.600 ;
        RECT 512.400 811.200 514.200 818.400 ;
        RECT 535.800 815.400 537.600 818.400 ;
        RECT 512.400 810.300 516.600 811.200 ;
        RECT 93.150 803.250 99.450 805.050 ;
        RECT 94.950 802.950 99.450 803.250 ;
        RECT 109.950 802.950 112.050 805.050 ;
        RECT 112.950 802.950 115.050 805.050 ;
        RECT 127.950 802.950 130.050 805.050 ;
        RECT 130.950 802.950 133.050 805.050 ;
        RECT 133.950 802.950 136.050 805.050 ;
        RECT 136.950 802.950 139.050 805.050 ;
        RECT 154.950 802.950 157.050 805.050 ;
        RECT 157.950 802.950 160.050 805.050 ;
        RECT 172.950 802.950 175.050 805.050 ;
        RECT 175.950 802.950 178.050 805.050 ;
        RECT 178.950 802.950 181.050 805.050 ;
        RECT 193.950 802.950 196.050 805.050 ;
        RECT 196.950 802.950 199.050 805.050 ;
        RECT 214.950 802.950 217.050 805.050 ;
        RECT 217.950 802.950 220.050 805.050 ;
        RECT 220.950 802.950 223.050 805.050 ;
        RECT 223.950 802.950 226.050 805.050 ;
        RECT 238.950 802.950 241.050 805.050 ;
        RECT 241.950 802.950 244.050 805.050 ;
        RECT 253.950 802.950 256.050 805.050 ;
        RECT 256.950 802.950 259.050 805.050 ;
        RECT 259.950 802.950 262.050 805.050 ;
        RECT 262.950 802.950 265.050 805.050 ;
        RECT 280.950 802.950 283.050 805.050 ;
        RECT 283.950 802.950 286.050 805.050 ;
        RECT 286.950 802.950 289.050 805.050 ;
        RECT 289.950 802.950 292.050 805.050 ;
        RECT 301.950 802.950 304.050 805.050 ;
        RECT 304.950 802.950 307.050 805.050 ;
        RECT 307.950 802.950 310.050 805.050 ;
        RECT 310.950 802.950 313.050 805.050 ;
        RECT 328.950 802.950 331.050 805.050 ;
        RECT 331.950 802.950 334.050 805.050 ;
        RECT 334.950 802.950 337.050 805.050 ;
        RECT 337.950 802.950 340.050 805.050 ;
        RECT 352.950 802.950 355.050 805.050 ;
        RECT 355.950 802.950 358.050 805.050 ;
        RECT 370.950 802.950 373.050 805.050 ;
        RECT 373.950 802.950 376.050 805.050 ;
        RECT 376.950 802.950 379.050 805.050 ;
        RECT 379.950 802.950 382.050 805.050 ;
        RECT 394.950 802.950 397.050 805.050 ;
        RECT 397.950 802.950 400.050 805.050 ;
        RECT 400.950 802.950 403.050 805.050 ;
        RECT 403.950 802.950 406.050 805.050 ;
        RECT 418.950 802.950 421.050 805.050 ;
        RECT 421.950 802.950 424.050 805.050 ;
        RECT 424.950 802.950 427.050 805.050 ;
        RECT 439.950 802.950 442.050 805.050 ;
        RECT 442.950 802.950 445.050 805.050 ;
        RECT 445.950 802.950 448.050 805.050 ;
        RECT 448.950 802.950 451.050 805.050 ;
        RECT 463.950 802.950 466.050 805.050 ;
        RECT 466.950 802.950 469.050 805.050 ;
        RECT 469.950 802.950 472.050 805.050 ;
        RECT 472.950 802.950 475.050 805.050 ;
        RECT 487.950 802.950 490.050 805.050 ;
        RECT 490.950 802.950 493.050 805.050 ;
        RECT 95.250 797.400 97.050 799.200 ;
        RECT 91.950 796.200 96.150 797.400 ;
        RECT 85.950 795.300 91.050 796.200 ;
        RECT 91.950 795.300 94.050 796.200 ;
        RECT 98.250 795.600 99.450 802.950 ;
        RECT 110.100 801.150 111.900 802.950 ;
        RECT 90.150 794.400 91.050 795.300 ;
        RECT 87.450 794.100 89.250 794.400 ;
        RECT 74.550 792.600 75.750 793.500 ;
        RECT 82.950 793.200 89.250 794.100 ;
        RECT 87.450 792.600 89.250 793.200 ;
        RECT 90.150 792.600 92.850 794.400 ;
        RECT 70.950 790.500 75.750 792.600 ;
        RECT 78.450 791.550 80.250 792.300 ;
        RECT 83.250 791.550 85.050 792.300 ;
        RECT 78.450 790.500 85.050 791.550 ;
        RECT 74.550 789.600 75.750 790.500 ;
        RECT 74.550 783.600 76.350 789.600 ;
        RECT 82.350 783.600 84.150 790.500 ;
        RECT 90.150 789.600 94.050 791.700 ;
        RECT 90.150 783.600 91.950 789.600 ;
        RECT 97.650 783.600 99.450 795.600 ;
        RECT 113.400 789.600 114.600 802.950 ;
        RECT 128.100 801.150 129.900 802.950 ;
        RECT 133.950 789.600 135.150 802.950 ;
        RECT 155.400 789.600 156.600 802.950 ;
        RECT 158.100 801.150 159.900 802.950 ;
        RECT 176.400 789.600 177.600 802.950 ;
        RECT 194.400 789.600 195.600 802.950 ;
        RECT 197.100 801.150 198.900 802.950 ;
        RECT 215.700 790.800 216.600 802.950 ;
        RECT 221.100 801.150 222.900 802.950 ;
        RECT 226.950 801.450 229.050 802.050 ;
        RECT 235.950 801.450 238.050 802.050 ;
        RECT 226.950 800.550 238.050 801.450 ;
        RECT 226.950 799.950 229.050 800.550 ;
        RECT 235.950 799.950 238.050 800.550 ;
        RECT 217.950 798.450 220.050 799.050 ;
        RECT 229.950 798.450 232.050 799.050 ;
        RECT 217.950 797.550 232.050 798.450 ;
        RECT 217.950 796.950 220.050 797.550 ;
        RECT 229.950 796.950 232.050 797.550 ;
        RECT 215.700 789.900 222.300 790.800 ;
        RECT 215.700 789.600 216.600 789.900 ;
        RECT 113.400 783.600 115.200 789.600 ;
        RECT 133.800 783.600 135.600 789.600 ;
        RECT 154.800 783.600 156.600 789.600 ;
        RECT 175.800 783.600 177.600 789.600 ;
        RECT 193.800 783.600 195.600 789.600 ;
        RECT 214.800 783.600 216.600 789.600 ;
        RECT 220.800 789.600 222.300 789.900 ;
        RECT 239.400 789.600 240.600 802.950 ;
        RECT 242.100 801.150 243.900 802.950 ;
        RECT 254.100 801.150 255.900 802.950 ;
        RECT 259.950 789.600 261.150 802.950 ;
        RECT 281.700 790.800 282.600 802.950 ;
        RECT 287.100 801.150 288.900 802.950 ;
        RECT 305.100 801.150 306.900 802.950 ;
        RECT 283.950 798.450 286.050 799.050 ;
        RECT 307.950 798.450 310.050 799.050 ;
        RECT 283.950 797.550 310.050 798.450 ;
        RECT 283.950 796.950 286.050 797.550 ;
        RECT 307.950 796.950 310.050 797.550 ;
        RECT 311.700 795.600 312.600 802.950 ;
        RECT 302.400 794.700 310.200 795.600 ;
        RECT 281.700 789.900 288.300 790.800 ;
        RECT 281.700 789.600 282.600 789.900 ;
        RECT 220.800 783.600 222.600 789.600 ;
        RECT 238.800 783.600 240.600 789.600 ;
        RECT 259.800 783.600 261.600 789.600 ;
        RECT 280.800 783.600 282.600 789.600 ;
        RECT 286.800 789.600 288.300 789.900 ;
        RECT 286.800 783.600 288.600 789.600 ;
        RECT 302.400 783.600 304.200 794.700 ;
        RECT 308.400 783.600 310.200 794.700 ;
        RECT 311.400 783.600 313.200 795.600 ;
        RECT 329.700 790.800 330.600 802.950 ;
        RECT 335.100 801.150 336.900 802.950 ;
        RECT 329.700 789.900 336.300 790.800 ;
        RECT 329.700 789.600 330.600 789.900 ;
        RECT 328.800 783.600 330.600 789.600 ;
        RECT 334.800 789.600 336.300 789.900 ;
        RECT 353.400 789.600 354.600 802.950 ;
        RECT 356.100 801.150 357.900 802.950 ;
        RECT 371.700 790.800 372.600 802.950 ;
        RECT 377.100 801.150 378.900 802.950 ;
        RECT 379.950 798.450 382.050 799.050 ;
        RECT 394.950 798.450 397.050 799.050 ;
        RECT 379.950 797.550 397.050 798.450 ;
        RECT 379.950 796.950 382.050 797.550 ;
        RECT 394.950 796.950 397.050 797.550 ;
        RECT 371.700 789.900 378.300 790.800 ;
        RECT 371.700 789.600 372.600 789.900 ;
        RECT 334.800 783.600 336.600 789.600 ;
        RECT 352.800 783.600 354.600 789.600 ;
        RECT 370.800 783.600 372.600 789.600 ;
        RECT 376.800 789.600 378.300 789.900 ;
        RECT 398.850 789.600 400.050 802.950 ;
        RECT 404.100 801.150 405.900 802.950 ;
        RECT 422.400 789.600 423.600 802.950 ;
        RECT 440.700 790.800 441.600 802.950 ;
        RECT 446.100 801.150 447.900 802.950 ;
        RECT 464.400 795.600 465.300 802.950 ;
        RECT 470.100 801.150 471.900 802.950 ;
        RECT 488.400 795.600 489.300 802.950 ;
        RECT 491.100 801.150 492.900 802.950 ;
        RECT 440.700 789.900 447.300 790.800 ;
        RECT 440.700 789.600 441.600 789.900 ;
        RECT 376.800 783.600 378.600 789.600 ;
        RECT 398.400 783.600 400.200 789.600 ;
        RECT 421.800 783.600 423.600 789.600 ;
        RECT 439.800 783.600 441.600 789.600 ;
        RECT 445.800 789.600 447.300 789.900 ;
        RECT 445.800 783.600 447.600 789.600 ;
        RECT 463.800 783.600 465.600 795.600 ;
        RECT 466.800 794.700 474.600 795.600 ;
        RECT 466.800 783.600 468.600 794.700 ;
        RECT 472.800 783.600 474.600 794.700 ;
        RECT 487.800 783.600 489.600 795.600 ;
        RECT 494.700 789.600 495.600 809.700 ;
        RECT 497.100 805.050 498.900 806.850 ;
        RECT 512.100 805.050 513.900 806.850 ;
        RECT 515.400 805.050 516.600 810.300 ;
        RECT 518.100 805.050 519.900 806.850 ;
        RECT 536.400 805.050 537.600 815.400 ;
        RECT 556.500 813.600 558.300 818.400 ;
        RECT 556.500 812.400 561.600 813.600 ;
        RECT 577.800 812.400 579.600 818.400 ;
        RECT 551.100 805.050 552.900 806.850 ;
        RECT 557.100 805.050 558.900 806.850 ;
        RECT 560.700 805.050 561.600 812.400 ;
        RECT 578.400 810.300 579.600 812.400 ;
        RECT 580.800 813.300 582.600 818.400 ;
        RECT 586.800 813.300 588.600 818.400 ;
        RECT 580.800 811.950 588.600 813.300 ;
        RECT 599.400 813.300 601.200 818.400 ;
        RECT 605.400 813.300 607.200 818.400 ;
        RECT 599.400 811.950 607.200 813.300 ;
        RECT 608.400 812.400 610.200 818.400 ;
        RECT 608.400 810.300 609.600 812.400 ;
        RECT 578.400 809.250 582.150 810.300 ;
        RECT 578.100 805.050 579.900 806.850 ;
        RECT 580.950 805.050 582.150 809.250 ;
        RECT 605.850 809.250 609.600 810.300 ;
        RECT 631.200 810.000 633.000 818.400 ;
        RECT 655.200 810.000 657.000 818.400 ;
        RECT 679.500 813.600 681.300 818.400 ;
        RECT 679.500 812.400 684.600 813.600 ;
        RECT 584.100 805.050 585.900 806.850 ;
        RECT 602.100 805.050 603.900 806.850 ;
        RECT 605.850 805.050 607.050 809.250 ;
        RECT 629.700 808.800 633.000 810.000 ;
        RECT 653.700 808.800 657.000 810.000 ;
        RECT 608.100 805.050 609.900 806.850 ;
        RECT 629.700 805.050 630.600 808.800 ;
        RECT 640.950 807.450 643.050 808.050 ;
        RECT 632.100 805.050 633.900 806.850 ;
        RECT 638.100 805.050 639.900 806.850 ;
        RECT 640.950 806.550 648.450 807.450 ;
        RECT 640.950 805.950 643.050 806.550 ;
        RECT 496.950 802.950 499.050 805.050 ;
        RECT 511.950 802.950 514.050 805.050 ;
        RECT 514.950 802.950 517.050 805.050 ;
        RECT 517.950 802.950 520.050 805.050 ;
        RECT 535.950 802.950 538.050 805.050 ;
        RECT 538.950 802.950 541.050 805.050 ;
        RECT 550.950 802.950 553.050 805.050 ;
        RECT 553.950 802.950 556.050 805.050 ;
        RECT 556.950 802.950 559.050 805.050 ;
        RECT 559.950 802.950 562.050 805.050 ;
        RECT 577.950 802.950 580.050 805.050 ;
        RECT 580.950 802.950 583.050 805.050 ;
        RECT 583.950 802.950 586.050 805.050 ;
        RECT 586.950 802.950 589.050 805.050 ;
        RECT 598.950 802.950 601.050 805.050 ;
        RECT 601.950 802.950 604.050 805.050 ;
        RECT 604.950 802.950 607.050 805.050 ;
        RECT 607.950 802.950 610.050 805.050 ;
        RECT 628.950 802.950 631.050 805.050 ;
        RECT 631.950 802.950 634.050 805.050 ;
        RECT 634.950 802.950 637.050 805.050 ;
        RECT 637.950 802.950 640.050 805.050 ;
        RECT 515.400 789.600 516.600 802.950 ;
        RECT 536.400 789.600 537.600 802.950 ;
        RECT 539.100 801.150 540.900 802.950 ;
        RECT 554.100 801.150 555.900 802.950 ;
        RECT 560.700 795.600 561.600 802.950 ;
        RECT 493.800 783.600 495.600 789.600 ;
        RECT 514.800 783.600 516.600 789.600 ;
        RECT 535.800 783.600 537.600 789.600 ;
        RECT 551.400 794.700 559.200 795.600 ;
        RECT 551.400 783.600 553.200 794.700 ;
        RECT 557.400 783.600 559.200 794.700 ;
        RECT 560.400 783.600 562.200 795.600 ;
        RECT 581.850 789.600 583.050 802.950 ;
        RECT 587.100 801.150 588.900 802.950 ;
        RECT 599.100 801.150 600.900 802.950 ;
        RECT 604.950 789.600 606.150 802.950 ;
        RECT 629.700 790.800 630.600 802.950 ;
        RECT 635.100 801.150 636.900 802.950 ;
        RECT 647.550 802.050 648.450 806.550 ;
        RECT 653.700 805.050 654.600 808.800 ;
        RECT 656.100 805.050 657.900 806.850 ;
        RECT 662.100 805.050 663.900 806.850 ;
        RECT 674.100 805.050 675.900 806.850 ;
        RECT 680.100 805.050 681.900 806.850 ;
        RECT 683.700 805.050 684.600 812.400 ;
        RECT 698.400 813.300 700.200 818.400 ;
        RECT 704.400 813.300 706.200 818.400 ;
        RECT 698.400 811.950 706.200 813.300 ;
        RECT 707.400 812.400 709.200 818.400 ;
        RECT 724.800 812.400 726.600 818.400 ;
        RECT 707.400 810.300 708.600 812.400 ;
        RECT 704.850 809.250 708.600 810.300 ;
        RECT 725.400 810.300 726.600 812.400 ;
        RECT 727.800 813.300 729.600 818.400 ;
        RECT 733.800 813.300 735.600 818.400 ;
        RECT 727.800 811.950 735.600 813.300 ;
        RECT 725.400 809.250 729.150 810.300 ;
        RECT 701.100 805.050 702.900 806.850 ;
        RECT 704.850 805.050 706.050 809.250 ;
        RECT 707.100 805.050 708.900 806.850 ;
        RECT 725.100 805.050 726.900 806.850 ;
        RECT 727.950 805.050 729.150 809.250 ;
        RECT 753.000 810.000 754.800 818.400 ;
        RECT 772.800 812.400 774.600 818.400 ;
        RECT 773.400 810.300 774.600 812.400 ;
        RECT 775.800 813.300 777.600 818.400 ;
        RECT 781.800 813.300 783.600 818.400 ;
        RECT 775.800 811.950 783.600 813.300 ;
        RECT 753.000 808.800 756.300 810.000 ;
        RECT 773.400 809.250 777.150 810.300 ;
        RECT 799.200 810.000 801.000 818.400 ;
        RECT 823.500 813.600 825.300 818.400 ;
        RECT 848.700 813.600 850.500 818.400 ;
        RECT 823.500 812.400 828.600 813.600 ;
        RECT 731.100 805.050 732.900 806.850 ;
        RECT 746.100 805.050 747.900 806.850 ;
        RECT 752.100 805.050 753.900 806.850 ;
        RECT 755.400 805.050 756.300 808.800 ;
        RECT 773.100 805.050 774.900 806.850 ;
        RECT 775.950 805.050 777.150 809.250 ;
        RECT 797.700 808.800 801.000 810.000 ;
        RECT 779.100 805.050 780.900 806.850 ;
        RECT 797.700 805.050 798.600 808.800 ;
        RECT 800.100 805.050 801.900 806.850 ;
        RECT 806.100 805.050 807.900 806.850 ;
        RECT 818.100 805.050 819.900 806.850 ;
        RECT 824.100 805.050 825.900 806.850 ;
        RECT 827.700 805.050 828.600 812.400 ;
        RECT 845.400 812.400 850.500 813.600 ;
        RECT 845.400 805.050 846.300 812.400 ;
        RECT 871.200 810.000 873.000 818.400 ;
        RECT 869.700 808.800 873.000 810.000 ;
        RECT 848.100 805.050 849.900 806.850 ;
        RECT 854.100 805.050 855.900 806.850 ;
        RECT 869.700 805.050 870.600 808.800 ;
        RECT 872.100 805.050 873.900 806.850 ;
        RECT 878.100 805.050 879.900 806.850 ;
        RECT 652.950 802.950 655.050 805.050 ;
        RECT 655.950 802.950 658.050 805.050 ;
        RECT 658.950 802.950 661.050 805.050 ;
        RECT 661.950 802.950 664.050 805.050 ;
        RECT 673.950 802.950 676.050 805.050 ;
        RECT 676.950 802.950 679.050 805.050 ;
        RECT 679.950 802.950 682.050 805.050 ;
        RECT 682.950 802.950 685.050 805.050 ;
        RECT 697.950 802.950 700.050 805.050 ;
        RECT 700.950 802.950 703.050 805.050 ;
        RECT 703.950 802.950 706.050 805.050 ;
        RECT 706.950 802.950 709.050 805.050 ;
        RECT 724.950 802.950 727.050 805.050 ;
        RECT 727.950 802.950 730.050 805.050 ;
        RECT 730.950 802.950 733.050 805.050 ;
        RECT 733.950 802.950 736.050 805.050 ;
        RECT 745.950 802.950 748.050 805.050 ;
        RECT 748.950 802.950 751.050 805.050 ;
        RECT 751.950 802.950 754.050 805.050 ;
        RECT 754.950 802.950 757.050 805.050 ;
        RECT 772.950 802.950 775.050 805.050 ;
        RECT 775.950 802.950 778.050 805.050 ;
        RECT 778.950 802.950 781.050 805.050 ;
        RECT 781.950 802.950 784.050 805.050 ;
        RECT 796.950 802.950 799.050 805.050 ;
        RECT 799.950 802.950 802.050 805.050 ;
        RECT 802.950 802.950 805.050 805.050 ;
        RECT 805.950 802.950 808.050 805.050 ;
        RECT 817.950 802.950 820.050 805.050 ;
        RECT 820.950 802.950 823.050 805.050 ;
        RECT 823.950 802.950 826.050 805.050 ;
        RECT 826.950 802.950 829.050 805.050 ;
        RECT 844.950 802.950 847.050 805.050 ;
        RECT 847.950 802.950 850.050 805.050 ;
        RECT 850.950 802.950 853.050 805.050 ;
        RECT 853.950 802.950 856.050 805.050 ;
        RECT 868.950 802.950 871.050 805.050 ;
        RECT 871.950 802.950 874.050 805.050 ;
        RECT 874.950 802.950 877.050 805.050 ;
        RECT 877.950 802.950 880.050 805.050 ;
        RECT 647.550 800.550 652.050 802.050 ;
        RECT 648.000 799.950 652.050 800.550 ;
        RECT 631.950 798.450 634.050 799.050 ;
        RECT 643.950 798.450 646.050 798.900 ;
        RECT 631.950 797.550 646.050 798.450 ;
        RECT 631.950 796.950 634.050 797.550 ;
        RECT 643.950 796.800 646.050 797.550 ;
        RECT 653.700 790.800 654.600 802.950 ;
        RECT 659.100 801.150 660.900 802.950 ;
        RECT 677.100 801.150 678.900 802.950 ;
        RECT 655.950 798.450 658.050 799.050 ;
        RECT 673.950 798.450 676.050 799.050 ;
        RECT 655.950 797.550 676.050 798.450 ;
        RECT 655.950 796.950 658.050 797.550 ;
        RECT 673.950 796.950 676.050 797.550 ;
        RECT 683.700 795.600 684.600 802.950 ;
        RECT 698.100 801.150 699.900 802.950 ;
        RECT 674.400 794.700 682.200 795.600 ;
        RECT 629.700 789.900 636.300 790.800 ;
        RECT 629.700 789.600 630.600 789.900 ;
        RECT 581.400 783.600 583.200 789.600 ;
        RECT 604.800 783.600 606.600 789.600 ;
        RECT 628.800 783.600 630.600 789.600 ;
        RECT 634.800 789.600 636.300 789.900 ;
        RECT 653.700 789.900 660.300 790.800 ;
        RECT 653.700 789.600 654.600 789.900 ;
        RECT 634.800 783.600 636.600 789.600 ;
        RECT 652.800 783.600 654.600 789.600 ;
        RECT 658.800 789.600 660.300 789.900 ;
        RECT 658.800 783.600 660.600 789.600 ;
        RECT 674.400 783.600 676.200 794.700 ;
        RECT 680.400 783.600 682.200 794.700 ;
        RECT 683.400 783.600 685.200 795.600 ;
        RECT 703.950 789.600 705.150 802.950 ;
        RECT 728.850 789.600 730.050 802.950 ;
        RECT 734.100 801.150 735.900 802.950 ;
        RECT 749.100 801.150 750.900 802.950 ;
        RECT 755.400 790.800 756.300 802.950 ;
        RECT 749.700 789.900 756.300 790.800 ;
        RECT 749.700 789.600 751.200 789.900 ;
        RECT 703.800 783.600 705.600 789.600 ;
        RECT 728.400 783.600 730.200 789.600 ;
        RECT 749.400 783.600 751.200 789.600 ;
        RECT 755.400 789.600 756.300 789.900 ;
        RECT 776.850 789.600 778.050 802.950 ;
        RECT 782.100 801.150 783.900 802.950 ;
        RECT 797.700 790.800 798.600 802.950 ;
        RECT 803.100 801.150 804.900 802.950 ;
        RECT 821.100 801.150 822.900 802.950 ;
        RECT 808.950 798.450 811.050 799.050 ;
        RECT 817.950 798.450 820.050 799.050 ;
        RECT 808.950 797.550 820.050 798.450 ;
        RECT 808.950 796.950 811.050 797.550 ;
        RECT 817.950 796.950 820.050 797.550 ;
        RECT 827.700 795.600 828.600 802.950 ;
        RECT 845.400 795.600 846.300 802.950 ;
        RECT 851.100 801.150 852.900 802.950 ;
        RECT 818.400 794.700 826.200 795.600 ;
        RECT 797.700 789.900 804.300 790.800 ;
        RECT 797.700 789.600 798.600 789.900 ;
        RECT 755.400 783.600 757.200 789.600 ;
        RECT 776.400 783.600 778.200 789.600 ;
        RECT 796.800 783.600 798.600 789.600 ;
        RECT 802.800 789.600 804.300 789.900 ;
        RECT 802.800 783.600 804.600 789.600 ;
        RECT 818.400 783.600 820.200 794.700 ;
        RECT 824.400 783.600 826.200 794.700 ;
        RECT 827.400 783.600 829.200 795.600 ;
        RECT 844.800 783.600 846.600 795.600 ;
        RECT 847.800 794.700 855.600 795.600 ;
        RECT 847.800 783.600 849.600 794.700 ;
        RECT 853.800 783.600 855.600 794.700 ;
        RECT 869.700 790.800 870.600 802.950 ;
        RECT 875.100 801.150 876.900 802.950 ;
        RECT 871.950 798.450 874.050 799.050 ;
        RECT 880.950 798.450 883.050 799.050 ;
        RECT 871.950 797.550 883.050 798.450 ;
        RECT 871.950 796.950 874.050 797.550 ;
        RECT 880.950 796.950 883.050 797.550 ;
        RECT 869.700 789.900 876.300 790.800 ;
        RECT 869.700 789.600 870.600 789.900 ;
        RECT 868.800 783.600 870.600 789.600 ;
        RECT 874.800 789.600 876.300 789.900 ;
        RECT 874.800 783.600 876.600 789.600 ;
        RECT 13.800 773.400 15.600 779.400 ;
        RECT 14.400 760.050 15.600 773.400 ;
        RECT 32.400 773.400 34.200 779.400 ;
        RECT 55.800 773.400 57.600 779.400 ;
        RECT 77.400 773.400 79.200 779.400 ;
        RECT 17.100 760.050 18.900 761.850 ;
        RECT 32.400 760.050 33.600 773.400 ;
        RECT 45.000 762.450 49.050 763.050 ;
        RECT 44.550 760.950 49.050 762.450 ;
        RECT 13.950 757.950 16.050 760.050 ;
        RECT 16.950 757.950 19.050 760.050 ;
        RECT 28.950 757.950 31.050 760.050 ;
        RECT 31.950 757.950 34.050 760.050 ;
        RECT 34.950 757.950 37.050 760.050 ;
        RECT 14.400 747.600 15.600 757.950 ;
        RECT 29.100 756.150 30.900 757.950 ;
        RECT 32.400 752.700 33.600 757.950 ;
        RECT 35.100 756.150 36.900 757.950 ;
        RECT 44.550 757.050 45.450 760.950 ;
        RECT 50.100 760.050 51.900 761.850 ;
        RECT 55.950 760.050 57.150 773.400 ;
        RECT 77.400 760.050 78.600 773.400 ;
        RECT 100.500 768.600 102.300 779.400 ;
        RECT 121.500 768.600 123.300 779.400 ;
        RECT 142.500 768.600 144.300 779.400 ;
        RECT 98.700 767.400 102.300 768.600 ;
        RECT 119.700 767.400 123.300 768.600 ;
        RECT 140.700 767.400 144.300 768.600 ;
        RECT 161.400 773.400 163.200 779.400 ;
        RECT 95.100 760.050 96.900 761.850 ;
        RECT 98.700 760.050 99.600 767.400 ;
        RECT 101.100 760.050 102.900 761.850 ;
        RECT 116.100 760.050 117.900 761.850 ;
        RECT 119.700 760.050 120.600 767.400 ;
        RECT 122.100 760.050 123.900 761.850 ;
        RECT 137.100 760.050 138.900 761.850 ;
        RECT 140.700 760.050 141.600 767.400 ;
        RECT 143.100 760.050 144.900 761.850 ;
        RECT 158.100 760.050 159.900 761.850 ;
        RECT 161.400 760.050 162.600 773.400 ;
        RECT 180.900 767.400 184.200 779.400 ;
        RECT 205.800 773.400 207.600 779.400 ;
        RECT 206.700 773.100 207.600 773.400 ;
        RECT 211.800 773.400 213.600 779.400 ;
        RECT 229.800 773.400 231.600 779.400 ;
        RECT 211.800 773.100 213.300 773.400 ;
        RECT 206.700 772.200 213.300 773.100 ;
        RECT 230.700 773.100 231.600 773.400 ;
        RECT 235.800 773.400 237.600 779.400 ;
        RECT 256.800 773.400 258.600 779.400 ;
        RECT 235.800 773.100 237.300 773.400 ;
        RECT 230.700 772.200 237.300 773.100 ;
        RECT 257.700 773.100 258.600 773.400 ;
        RECT 262.800 773.400 264.600 779.400 ;
        RECT 262.800 773.100 264.300 773.400 ;
        RECT 257.700 772.200 264.300 773.100 ;
        RECT 176.100 760.050 177.900 761.850 ;
        RECT 182.100 760.050 183.300 767.400 ;
        RECT 188.100 760.050 189.900 761.850 ;
        RECT 206.700 760.050 207.600 772.200 ;
        RECT 212.100 760.050 213.900 761.850 ;
        RECT 230.700 760.050 231.600 772.200 ;
        RECT 236.100 760.050 237.900 761.850 ;
        RECT 257.700 760.050 258.600 772.200 ;
        RECT 280.800 767.400 282.600 779.400 ;
        RECT 283.800 768.300 285.600 779.400 ;
        RECT 289.800 768.300 291.600 779.400 ;
        RECT 305.400 773.400 307.200 779.400 ;
        RECT 305.700 773.100 307.200 773.400 ;
        RECT 311.400 773.400 313.200 779.400 ;
        RECT 329.400 773.400 331.200 779.400 ;
        RECT 349.800 773.400 351.600 779.400 ;
        RECT 371.400 773.400 373.200 779.400 ;
        RECT 394.800 773.400 396.600 779.400 ;
        RECT 311.400 773.100 312.300 773.400 ;
        RECT 305.700 772.200 312.300 773.100 ;
        RECT 283.800 767.400 291.600 768.300 ;
        RECT 263.100 760.050 264.900 761.850 ;
        RECT 281.400 760.050 282.300 767.400 ;
        RECT 283.950 765.450 286.050 766.050 ;
        RECT 301.950 765.450 304.050 766.050 ;
        RECT 283.950 764.550 304.050 765.450 ;
        RECT 283.950 763.950 286.050 764.550 ;
        RECT 301.950 763.950 304.050 764.550 ;
        RECT 287.100 760.050 288.900 761.850 ;
        RECT 305.100 760.050 306.900 761.850 ;
        RECT 311.400 760.050 312.300 772.200 ;
        RECT 329.400 760.050 330.600 773.400 ;
        RECT 350.400 760.050 351.600 773.400 ;
        RECT 353.100 760.050 354.900 761.850 ;
        RECT 371.850 760.050 373.050 773.400 ;
        RECT 377.100 760.050 378.900 761.850 ;
        RECT 395.400 760.050 396.600 773.400 ;
        RECT 413.400 773.400 415.200 779.400 ;
        RECT 405.000 762.450 409.050 763.050 ;
        RECT 398.100 760.050 399.900 761.850 ;
        RECT 404.550 760.950 409.050 762.450 ;
        RECT 49.950 757.950 52.050 760.050 ;
        RECT 52.950 757.950 55.050 760.050 ;
        RECT 55.950 757.950 58.050 760.050 ;
        RECT 58.950 757.950 61.050 760.050 ;
        RECT 73.950 757.950 76.050 760.050 ;
        RECT 76.950 757.950 79.050 760.050 ;
        RECT 79.950 757.950 82.050 760.050 ;
        RECT 94.950 757.950 97.050 760.050 ;
        RECT 97.950 757.950 100.050 760.050 ;
        RECT 100.950 757.950 103.050 760.050 ;
        RECT 115.950 757.950 118.050 760.050 ;
        RECT 118.950 757.950 121.050 760.050 ;
        RECT 121.950 757.950 124.050 760.050 ;
        RECT 136.950 757.950 139.050 760.050 ;
        RECT 139.950 757.950 142.050 760.050 ;
        RECT 142.950 757.950 145.050 760.050 ;
        RECT 157.950 757.950 160.050 760.050 ;
        RECT 160.950 757.950 163.050 760.050 ;
        RECT 175.950 757.950 178.050 760.050 ;
        RECT 178.950 757.950 181.050 760.050 ;
        RECT 181.950 757.950 184.050 760.050 ;
        RECT 184.950 757.950 187.050 760.050 ;
        RECT 187.950 757.950 190.050 760.050 ;
        RECT 205.950 757.950 208.050 760.050 ;
        RECT 208.950 757.950 211.050 760.050 ;
        RECT 211.950 757.950 214.050 760.050 ;
        RECT 214.950 757.950 217.050 760.050 ;
        RECT 229.950 757.950 232.050 760.050 ;
        RECT 232.950 757.950 235.050 760.050 ;
        RECT 235.950 757.950 238.050 760.050 ;
        RECT 238.950 757.950 241.050 760.050 ;
        RECT 256.950 757.950 259.050 760.050 ;
        RECT 259.950 757.950 262.050 760.050 ;
        RECT 262.950 757.950 265.050 760.050 ;
        RECT 265.950 757.950 268.050 760.050 ;
        RECT 280.950 757.950 283.050 760.050 ;
        RECT 283.950 757.950 286.050 760.050 ;
        RECT 286.950 757.950 289.050 760.050 ;
        RECT 289.950 757.950 292.050 760.050 ;
        RECT 301.950 757.950 304.050 760.050 ;
        RECT 304.950 757.950 307.050 760.050 ;
        RECT 307.950 757.950 310.050 760.050 ;
        RECT 310.950 757.950 313.050 760.050 ;
        RECT 325.950 757.950 328.050 760.050 ;
        RECT 328.950 757.950 331.050 760.050 ;
        RECT 331.950 757.950 334.050 760.050 ;
        RECT 349.950 757.950 352.050 760.050 ;
        RECT 352.950 757.950 355.050 760.050 ;
        RECT 367.950 757.950 370.050 760.050 ;
        RECT 370.950 757.950 373.050 760.050 ;
        RECT 373.950 757.950 376.050 760.050 ;
        RECT 376.950 757.950 379.050 760.050 ;
        RECT 394.950 757.950 397.050 760.050 ;
        RECT 397.950 757.950 400.050 760.050 ;
        RECT 44.550 755.550 49.050 757.050 ;
        RECT 53.100 756.150 54.900 757.950 ;
        RECT 45.000 754.950 49.050 755.550 ;
        RECT 56.850 753.750 58.050 757.950 ;
        RECT 59.100 756.150 60.900 757.950 ;
        RECT 74.100 756.150 75.900 757.950 ;
        RECT 56.850 752.700 60.600 753.750 ;
        RECT 32.400 751.800 36.600 752.700 ;
        RECT 13.800 744.600 15.600 747.600 ;
        RECT 34.800 744.600 36.600 751.800 ;
        RECT 50.400 749.700 58.200 751.050 ;
        RECT 50.400 744.600 52.200 749.700 ;
        RECT 56.400 744.600 58.200 749.700 ;
        RECT 59.400 750.600 60.600 752.700 ;
        RECT 77.400 752.700 78.600 757.950 ;
        RECT 80.100 756.150 81.900 757.950 ;
        RECT 77.400 751.800 81.600 752.700 ;
        RECT 59.400 744.600 61.200 750.600 ;
        RECT 79.800 744.600 81.600 751.800 ;
        RECT 98.700 747.600 99.600 757.950 ;
        RECT 119.700 747.600 120.600 757.950 ;
        RECT 140.700 747.600 141.600 757.950 ;
        RECT 161.400 747.600 162.600 757.950 ;
        RECT 179.100 756.150 180.900 757.950 ;
        RECT 181.950 753.300 183.300 757.950 ;
        RECT 185.100 756.150 186.900 757.950 ;
        RECT 206.700 754.200 207.600 757.950 ;
        RECT 209.100 756.150 210.900 757.950 ;
        RECT 215.100 756.150 216.900 757.950 ;
        RECT 230.700 754.200 231.600 757.950 ;
        RECT 233.100 756.150 234.900 757.950 ;
        RECT 239.100 756.150 240.900 757.950 ;
        RECT 257.700 754.200 258.600 757.950 ;
        RECT 260.100 756.150 261.900 757.950 ;
        RECT 266.100 756.150 267.900 757.950 ;
        RECT 181.950 752.100 186.600 753.300 ;
        RECT 206.700 753.000 210.000 754.200 ;
        RECT 230.700 753.000 234.000 754.200 ;
        RECT 257.700 753.000 261.000 754.200 ;
        RECT 176.400 750.000 184.200 750.900 ;
        RECT 185.700 750.600 186.600 752.100 ;
        RECT 98.400 744.600 100.200 747.600 ;
        RECT 119.400 744.600 121.200 747.600 ;
        RECT 140.400 744.600 142.200 747.600 ;
        RECT 161.400 744.600 163.200 747.600 ;
        RECT 176.400 744.600 178.200 750.000 ;
        RECT 182.400 745.500 184.200 750.000 ;
        RECT 185.400 746.400 187.200 750.600 ;
        RECT 188.400 745.500 190.200 750.600 ;
        RECT 182.400 744.600 190.200 745.500 ;
        RECT 208.200 744.600 210.000 753.000 ;
        RECT 232.200 744.600 234.000 753.000 ;
        RECT 259.200 744.600 261.000 753.000 ;
        RECT 281.400 750.600 282.300 757.950 ;
        RECT 284.100 756.150 285.900 757.950 ;
        RECT 290.100 756.150 291.900 757.950 ;
        RECT 302.100 756.150 303.900 757.950 ;
        RECT 308.100 756.150 309.900 757.950 ;
        RECT 311.400 754.200 312.300 757.950 ;
        RECT 326.100 756.150 327.900 757.950 ;
        RECT 309.000 753.000 312.300 754.200 ;
        RECT 281.400 749.400 286.500 750.600 ;
        RECT 284.700 744.600 286.500 749.400 ;
        RECT 309.000 744.600 310.800 753.000 ;
        RECT 329.400 752.700 330.600 757.950 ;
        RECT 332.100 756.150 333.900 757.950 ;
        RECT 329.400 751.800 333.600 752.700 ;
        RECT 331.800 744.600 333.600 751.800 ;
        RECT 350.400 747.600 351.600 757.950 ;
        RECT 368.100 756.150 369.900 757.950 ;
        RECT 370.950 753.750 372.150 757.950 ;
        RECT 374.100 756.150 375.900 757.950 ;
        RECT 368.400 752.700 372.150 753.750 ;
        RECT 368.400 750.600 369.600 752.700 ;
        RECT 349.800 744.600 351.600 747.600 ;
        RECT 367.800 744.600 369.600 750.600 ;
        RECT 370.800 749.700 378.600 751.050 ;
        RECT 370.800 744.600 372.600 749.700 ;
        RECT 376.800 744.600 378.600 749.700 ;
        RECT 395.400 747.600 396.600 757.950 ;
        RECT 404.550 757.050 405.450 760.950 ;
        RECT 413.400 760.050 414.600 773.400 ;
        RECT 439.800 767.400 443.100 779.400 ;
        RECT 463.500 768.600 465.300 779.400 ;
        RECT 484.800 773.400 486.600 779.400 ;
        RECT 509.400 773.400 511.200 779.400 ;
        RECT 461.700 767.400 465.300 768.600 ;
        RECT 434.100 760.050 435.900 761.850 ;
        RECT 440.700 760.050 441.900 767.400 ;
        RECT 446.100 760.050 447.900 761.850 ;
        RECT 458.100 760.050 459.900 761.850 ;
        RECT 461.700 760.050 462.600 767.400 ;
        RECT 464.100 760.050 465.900 761.850 ;
        RECT 479.100 760.050 480.900 761.850 ;
        RECT 484.950 760.050 486.150 773.400 ;
        RECT 509.700 773.100 511.200 773.400 ;
        RECT 515.400 773.400 517.200 779.400 ;
        RECT 532.800 773.400 534.600 779.400 ;
        RECT 551.400 773.400 553.200 779.400 ;
        RECT 515.400 773.100 516.300 773.400 ;
        RECT 509.700 772.200 516.300 773.100 ;
        RECT 493.950 768.450 496.050 769.050 ;
        RECT 505.950 768.450 508.050 769.050 ;
        RECT 493.950 767.550 508.050 768.450 ;
        RECT 493.950 766.950 496.050 767.550 ;
        RECT 505.950 766.950 508.050 767.550 ;
        RECT 499.950 765.450 502.050 766.050 ;
        RECT 511.950 765.450 514.050 766.050 ;
        RECT 499.950 764.550 514.050 765.450 ;
        RECT 499.950 763.950 502.050 764.550 ;
        RECT 511.950 763.950 514.050 764.550 ;
        RECT 509.100 760.050 510.900 761.850 ;
        RECT 515.400 760.050 516.300 772.200 ;
        RECT 533.400 760.050 534.600 773.400 ;
        RECT 551.700 773.100 553.200 773.400 ;
        RECT 557.400 773.400 559.200 779.400 ;
        RECT 578.400 773.400 580.200 779.400 ;
        RECT 599.400 773.400 601.200 779.400 ;
        RECT 620.400 773.400 622.200 779.400 ;
        RECT 557.400 773.100 558.300 773.400 ;
        RECT 551.700 772.200 558.300 773.100 ;
        RECT 536.100 760.050 537.900 761.850 ;
        RECT 551.100 760.050 552.900 761.850 ;
        RECT 557.400 760.050 558.300 772.200 ;
        RECT 570.000 762.450 574.050 763.050 ;
        RECT 569.550 760.950 574.050 762.450 ;
        RECT 409.950 757.950 412.050 760.050 ;
        RECT 412.950 757.950 415.050 760.050 ;
        RECT 415.950 757.950 418.050 760.050 ;
        RECT 433.950 757.950 436.050 760.050 ;
        RECT 436.950 757.950 439.050 760.050 ;
        RECT 439.950 757.950 442.050 760.050 ;
        RECT 442.950 757.950 445.050 760.050 ;
        RECT 445.950 757.950 448.050 760.050 ;
        RECT 457.950 757.950 460.050 760.050 ;
        RECT 460.950 757.950 463.050 760.050 ;
        RECT 463.950 757.950 466.050 760.050 ;
        RECT 478.950 757.950 481.050 760.050 ;
        RECT 481.950 757.950 484.050 760.050 ;
        RECT 484.950 757.950 487.050 760.050 ;
        RECT 487.950 757.950 490.050 760.050 ;
        RECT 505.950 757.950 508.050 760.050 ;
        RECT 508.950 757.950 511.050 760.050 ;
        RECT 511.950 757.950 514.050 760.050 ;
        RECT 514.950 757.950 517.050 760.050 ;
        RECT 532.950 757.950 535.050 760.050 ;
        RECT 535.950 757.950 538.050 760.050 ;
        RECT 547.950 757.950 550.050 760.050 ;
        RECT 550.950 757.950 553.050 760.050 ;
        RECT 553.950 757.950 556.050 760.050 ;
        RECT 556.950 757.950 559.050 760.050 ;
        RECT 404.550 755.550 409.050 757.050 ;
        RECT 410.100 756.150 411.900 757.950 ;
        RECT 405.000 754.950 409.050 755.550 ;
        RECT 413.400 752.700 414.600 757.950 ;
        RECT 416.100 756.150 417.900 757.950 ;
        RECT 437.100 756.150 438.900 757.950 ;
        RECT 440.700 753.300 442.050 757.950 ;
        RECT 443.100 756.150 444.900 757.950 ;
        RECT 413.400 751.800 417.600 752.700 ;
        RECT 394.800 744.600 396.600 747.600 ;
        RECT 415.800 744.600 417.600 751.800 ;
        RECT 437.400 752.100 442.050 753.300 ;
        RECT 437.400 750.600 438.300 752.100 ;
        RECT 433.800 745.500 435.600 750.600 ;
        RECT 436.800 746.400 438.600 750.600 ;
        RECT 439.800 750.000 447.600 750.900 ;
        RECT 439.800 745.500 441.600 750.000 ;
        RECT 433.800 744.600 441.600 745.500 ;
        RECT 445.800 744.600 447.600 750.000 ;
        RECT 461.700 747.600 462.600 757.950 ;
        RECT 482.100 756.150 483.900 757.950 ;
        RECT 485.850 753.750 487.050 757.950 ;
        RECT 488.100 756.150 489.900 757.950 ;
        RECT 506.100 756.150 507.900 757.950 ;
        RECT 512.100 756.150 513.900 757.950 ;
        RECT 515.400 754.200 516.300 757.950 ;
        RECT 485.850 752.700 489.600 753.750 ;
        RECT 479.400 749.700 487.200 751.050 ;
        RECT 461.400 744.600 463.200 747.600 ;
        RECT 479.400 744.600 481.200 749.700 ;
        RECT 485.400 744.600 487.200 749.700 ;
        RECT 488.400 750.600 489.600 752.700 ;
        RECT 513.000 753.000 516.300 754.200 ;
        RECT 488.400 744.600 490.200 750.600 ;
        RECT 513.000 744.600 514.800 753.000 ;
        RECT 533.400 747.600 534.600 757.950 ;
        RECT 548.100 756.150 549.900 757.950 ;
        RECT 554.100 756.150 555.900 757.950 ;
        RECT 557.400 754.200 558.300 757.950 ;
        RECT 559.950 756.450 562.050 757.050 ;
        RECT 569.550 756.450 570.450 760.950 ;
        RECT 578.850 760.050 580.050 773.400 ;
        RECT 584.100 760.050 585.900 761.850 ;
        RECT 599.400 760.050 600.600 773.400 ;
        RECT 620.700 773.100 622.200 773.400 ;
        RECT 626.400 773.400 628.200 779.400 ;
        RECT 643.800 773.400 645.600 779.400 ;
        RECT 661.800 773.400 663.600 779.400 ;
        RECT 680.400 773.400 682.200 779.400 ;
        RECT 626.400 773.100 627.300 773.400 ;
        RECT 620.700 772.200 627.300 773.100 ;
        RECT 620.100 760.050 621.900 761.850 ;
        RECT 626.400 760.050 627.300 772.200 ;
        RECT 644.400 760.050 645.600 773.400 ;
        RECT 647.100 760.050 648.900 761.850 ;
        RECT 662.400 760.050 663.600 773.400 ;
        RECT 680.700 773.100 682.200 773.400 ;
        RECT 686.400 773.400 688.200 779.400 ;
        RECT 703.800 773.400 705.600 779.400 ;
        RECT 686.400 773.100 687.300 773.400 ;
        RECT 680.700 772.200 687.300 773.100 ;
        RECT 667.950 762.450 672.000 763.050 ;
        RECT 665.100 760.050 666.900 761.850 ;
        RECT 667.950 760.950 672.450 762.450 ;
        RECT 574.950 757.950 577.050 760.050 ;
        RECT 577.950 757.950 580.050 760.050 ;
        RECT 580.950 757.950 583.050 760.050 ;
        RECT 583.950 757.950 586.050 760.050 ;
        RECT 595.950 757.950 598.050 760.050 ;
        RECT 598.950 757.950 601.050 760.050 ;
        RECT 601.950 757.950 604.050 760.050 ;
        RECT 616.950 757.950 619.050 760.050 ;
        RECT 619.950 757.950 622.050 760.050 ;
        RECT 622.950 757.950 625.050 760.050 ;
        RECT 625.950 757.950 628.050 760.050 ;
        RECT 643.950 757.950 646.050 760.050 ;
        RECT 646.950 757.950 649.050 760.050 ;
        RECT 661.950 757.950 664.050 760.050 ;
        RECT 664.950 757.950 667.050 760.050 ;
        RECT 559.950 755.550 570.450 756.450 ;
        RECT 575.100 756.150 576.900 757.950 ;
        RECT 559.950 754.950 562.050 755.550 ;
        RECT 532.800 744.600 534.600 747.600 ;
        RECT 555.000 753.000 558.300 754.200 ;
        RECT 577.950 753.750 579.150 757.950 ;
        RECT 581.100 756.150 582.900 757.950 ;
        RECT 596.100 756.150 597.900 757.950 ;
        RECT 555.000 744.600 556.800 753.000 ;
        RECT 575.400 752.700 579.150 753.750 ;
        RECT 599.400 752.700 600.600 757.950 ;
        RECT 602.100 756.150 603.900 757.950 ;
        RECT 617.100 756.150 618.900 757.950 ;
        RECT 623.100 756.150 624.900 757.950 ;
        RECT 626.400 754.200 627.300 757.950 ;
        RECT 624.000 753.000 627.300 754.200 ;
        RECT 575.400 750.600 576.600 752.700 ;
        RECT 599.400 751.800 603.600 752.700 ;
        RECT 574.800 744.600 576.600 750.600 ;
        RECT 577.800 749.700 585.600 751.050 ;
        RECT 577.800 744.600 579.600 749.700 ;
        RECT 583.800 744.600 585.600 749.700 ;
        RECT 601.800 744.600 603.600 751.800 ;
        RECT 624.000 744.600 625.800 753.000 ;
        RECT 644.400 747.600 645.600 757.950 ;
        RECT 662.400 747.600 663.600 757.950 ;
        RECT 671.550 757.050 672.450 760.950 ;
        RECT 680.100 760.050 681.900 761.850 ;
        RECT 686.400 760.050 687.300 772.200 ;
        RECT 704.700 773.100 705.600 773.400 ;
        RECT 709.800 773.400 711.600 779.400 ;
        RECT 709.800 773.100 711.300 773.400 ;
        RECT 704.700 772.200 711.300 773.100 ;
        RECT 704.700 760.050 705.600 772.200 ;
        RECT 709.950 768.450 712.050 769.050 ;
        RECT 715.950 768.450 718.050 769.050 ;
        RECT 709.950 767.550 718.050 768.450 ;
        RECT 709.950 766.950 712.050 767.550 ;
        RECT 715.950 766.950 718.050 767.550 ;
        RECT 725.400 768.300 727.200 779.400 ;
        RECT 731.400 768.300 733.200 779.400 ;
        RECT 725.400 767.400 733.200 768.300 ;
        RECT 734.400 767.400 736.200 779.400 ;
        RECT 752.400 773.400 754.200 779.400 ;
        RECT 775.800 773.400 777.600 779.400 ;
        RECT 710.100 760.050 711.900 761.850 ;
        RECT 728.100 760.050 729.900 761.850 ;
        RECT 734.700 760.050 735.600 767.400 ;
        RECT 752.400 760.050 753.600 773.400 ;
        RECT 776.400 760.050 777.600 773.400 ;
        RECT 794.400 773.400 796.200 779.400 ;
        RECT 676.950 757.950 679.050 760.050 ;
        RECT 679.950 757.950 682.050 760.050 ;
        RECT 682.950 757.950 685.050 760.050 ;
        RECT 685.950 757.950 688.050 760.050 ;
        RECT 703.950 757.950 706.050 760.050 ;
        RECT 706.950 757.950 709.050 760.050 ;
        RECT 709.950 757.950 712.050 760.050 ;
        RECT 712.950 757.950 715.050 760.050 ;
        RECT 724.950 757.950 727.050 760.050 ;
        RECT 727.950 757.950 730.050 760.050 ;
        RECT 730.950 757.950 733.050 760.050 ;
        RECT 733.950 757.950 736.050 760.050 ;
        RECT 748.950 757.950 751.050 760.050 ;
        RECT 751.950 757.950 754.050 760.050 ;
        RECT 754.950 757.950 757.050 760.050 ;
        RECT 772.950 757.950 775.050 760.050 ;
        RECT 775.950 757.950 778.050 760.050 ;
        RECT 778.950 757.950 781.050 760.050 ;
        RECT 790.950 757.950 793.050 760.050 ;
        RECT 671.550 755.550 676.050 757.050 ;
        RECT 677.100 756.150 678.900 757.950 ;
        RECT 683.100 756.150 684.900 757.950 ;
        RECT 672.000 754.950 676.050 755.550 ;
        RECT 686.400 754.200 687.300 757.950 ;
        RECT 643.800 744.600 645.600 747.600 ;
        RECT 661.800 744.600 663.600 747.600 ;
        RECT 684.000 753.000 687.300 754.200 ;
        RECT 704.700 754.200 705.600 757.950 ;
        RECT 707.100 756.150 708.900 757.950 ;
        RECT 713.100 756.150 714.900 757.950 ;
        RECT 725.100 756.150 726.900 757.950 ;
        RECT 731.100 756.150 732.900 757.950 ;
        RECT 704.700 753.000 708.000 754.200 ;
        RECT 684.000 744.600 685.800 753.000 ;
        RECT 706.200 744.600 708.000 753.000 ;
        RECT 718.950 753.450 721.050 754.050 ;
        RECT 730.950 753.450 733.050 754.050 ;
        RECT 718.950 752.550 733.050 753.450 ;
        RECT 718.950 751.950 721.050 752.550 ;
        RECT 730.950 751.950 733.050 752.550 ;
        RECT 734.700 750.600 735.600 757.950 ;
        RECT 749.100 756.150 750.900 757.950 ;
        RECT 752.400 752.700 753.600 757.950 ;
        RECT 755.100 756.150 756.900 757.950 ;
        RECT 773.100 756.150 774.900 757.950 ;
        RECT 776.400 752.700 777.600 757.950 ;
        RECT 779.100 756.150 780.900 757.950 ;
        RECT 791.100 756.150 792.900 757.950 ;
        RECT 794.400 753.300 795.300 773.400 ;
        RECT 800.400 767.400 802.200 779.400 ;
        RECT 815.400 768.300 817.200 779.400 ;
        RECT 821.400 768.300 823.200 779.400 ;
        RECT 815.400 767.400 823.200 768.300 ;
        RECT 824.400 767.400 826.200 779.400 ;
        RECT 844.800 773.400 846.600 779.400 ;
        RECT 863.400 773.400 865.200 779.400 ;
        RECT 797.100 760.050 798.900 761.850 ;
        RECT 800.700 760.050 801.600 767.400 ;
        RECT 818.100 760.050 819.900 761.850 ;
        RECT 824.700 760.050 825.600 767.400 ;
        RECT 829.950 762.450 832.050 763.050 ;
        RECT 841.950 762.450 844.050 763.050 ;
        RECT 829.950 761.550 844.050 762.450 ;
        RECT 829.950 760.950 832.050 761.550 ;
        RECT 841.950 760.950 844.050 761.550 ;
        RECT 845.400 760.050 846.600 773.400 ;
        RECT 863.700 773.100 865.200 773.400 ;
        RECT 869.400 773.400 871.200 779.400 ;
        RECT 869.400 773.100 870.300 773.400 ;
        RECT 863.700 772.200 870.300 773.100 ;
        RECT 850.950 765.450 853.050 766.050 ;
        RECT 865.950 765.450 868.050 766.050 ;
        RECT 850.950 764.550 868.050 765.450 ;
        RECT 850.950 763.950 853.050 764.550 ;
        RECT 865.950 763.950 868.050 764.550 ;
        RECT 855.000 762.450 859.050 763.050 ;
        RECT 848.100 760.050 849.900 761.850 ;
        RECT 854.550 760.950 859.050 762.450 ;
        RECT 796.950 757.950 799.050 760.050 ;
        RECT 799.950 757.950 802.050 760.050 ;
        RECT 814.950 757.950 817.050 760.050 ;
        RECT 817.950 757.950 820.050 760.050 ;
        RECT 820.950 757.950 823.050 760.050 ;
        RECT 823.950 757.950 826.050 760.050 ;
        RECT 844.950 757.950 847.050 760.050 ;
        RECT 847.950 757.950 850.050 760.050 ;
        RECT 752.400 751.800 756.600 752.700 ;
        RECT 730.500 749.400 735.600 750.600 ;
        RECT 730.500 744.600 732.300 749.400 ;
        RECT 754.800 744.600 756.600 751.800 ;
        RECT 773.400 751.800 777.600 752.700 ;
        RECT 791.400 752.400 798.900 753.300 ;
        RECT 773.400 744.600 775.200 751.800 ;
        RECT 791.400 744.600 793.200 752.400 ;
        RECT 797.100 751.500 798.900 752.400 ;
        RECT 800.700 750.600 801.600 757.950 ;
        RECT 815.100 756.150 816.900 757.950 ;
        RECT 821.100 756.150 822.900 757.950 ;
        RECT 824.700 750.600 825.600 757.950 ;
        RECT 798.900 748.800 801.600 750.600 ;
        RECT 820.500 749.400 825.600 750.600 ;
        RECT 798.900 744.600 800.700 748.800 ;
        RECT 820.500 744.600 822.300 749.400 ;
        RECT 845.400 747.600 846.600 757.950 ;
        RECT 854.550 757.050 855.450 760.950 ;
        RECT 863.100 760.050 864.900 761.850 ;
        RECT 869.400 760.050 870.300 772.200 ;
        RECT 859.950 757.950 862.050 760.050 ;
        RECT 862.950 757.950 865.050 760.050 ;
        RECT 865.950 757.950 868.050 760.050 ;
        RECT 868.950 757.950 871.050 760.050 ;
        RECT 850.950 755.550 855.450 757.050 ;
        RECT 860.100 756.150 861.900 757.950 ;
        RECT 866.100 756.150 867.900 757.950 ;
        RECT 850.950 754.950 855.000 755.550 ;
        RECT 869.400 754.200 870.300 757.950 ;
        RECT 844.800 744.600 846.600 747.600 ;
        RECT 867.000 753.000 870.300 754.200 ;
        RECT 867.000 744.600 868.800 753.000 ;
        RECT 16.800 733.200 18.600 740.400 ;
        RECT 14.400 732.300 18.600 733.200 ;
        RECT 35.400 737.400 37.200 740.400 ;
        RECT 52.800 737.400 54.600 740.400 ;
        RECT 11.100 727.050 12.900 728.850 ;
        RECT 14.400 727.050 15.600 732.300 ;
        RECT 17.100 727.050 18.900 728.850 ;
        RECT 35.400 727.050 36.600 737.400 ;
        RECT 53.400 727.050 54.600 737.400 ;
        RECT 70.800 734.400 72.600 740.400 ;
        RECT 71.400 732.300 72.600 734.400 ;
        RECT 73.800 735.300 75.600 740.400 ;
        RECT 79.800 735.300 81.600 740.400 ;
        RECT 94.800 737.400 96.600 740.400 ;
        RECT 73.800 733.950 81.600 735.300 ;
        RECT 71.400 731.250 75.150 732.300 ;
        RECT 71.100 727.050 72.900 728.850 ;
        RECT 73.950 727.050 75.150 731.250 ;
        RECT 77.100 727.050 78.900 728.850 ;
        RECT 95.400 727.050 96.600 737.400 ;
        RECT 101.550 734.400 103.350 740.400 ;
        RECT 109.650 737.400 111.450 740.400 ;
        RECT 117.450 737.400 119.250 740.400 ;
        RECT 125.250 738.300 127.050 740.400 ;
        RECT 125.250 737.400 129.000 738.300 ;
        RECT 109.650 736.500 110.700 737.400 ;
        RECT 106.950 735.300 110.700 736.500 ;
        RECT 118.200 736.500 119.250 737.400 ;
        RECT 127.950 736.500 129.000 737.400 ;
        RECT 118.200 735.450 123.150 736.500 ;
        RECT 106.950 734.400 109.050 735.300 ;
        RECT 121.350 734.700 123.150 735.450 ;
        RECT 101.550 727.050 102.750 734.400 ;
        RECT 124.650 733.800 126.450 735.600 ;
        RECT 127.950 734.400 130.050 736.500 ;
        RECT 133.050 734.400 134.850 740.400 ;
        RECT 148.800 734.400 150.600 740.400 ;
        RECT 114.150 732.000 115.950 732.600 ;
        RECT 125.100 732.000 126.150 733.800 ;
        RECT 114.150 730.800 126.150 732.000 ;
        RECT 10.950 724.950 13.050 727.050 ;
        RECT 13.950 724.950 16.050 727.050 ;
        RECT 16.950 724.950 19.050 727.050 ;
        RECT 31.950 724.950 34.050 727.050 ;
        RECT 34.950 724.950 37.050 727.050 ;
        RECT 52.950 724.950 55.050 727.050 ;
        RECT 55.950 724.950 58.050 727.050 ;
        RECT 70.950 724.950 73.050 727.050 ;
        RECT 73.950 724.950 76.050 727.050 ;
        RECT 76.950 724.950 79.050 727.050 ;
        RECT 79.950 724.950 82.050 727.050 ;
        RECT 94.950 724.950 97.050 727.050 ;
        RECT 97.950 724.950 100.050 727.050 ;
        RECT 101.550 725.250 107.850 727.050 ;
        RECT 101.550 724.950 106.050 725.250 ;
        RECT 14.400 711.600 15.600 724.950 ;
        RECT 32.100 723.150 33.900 724.950 ;
        RECT 35.400 711.600 36.600 724.950 ;
        RECT 40.950 723.450 43.050 724.050 ;
        RECT 49.950 723.450 52.050 724.050 ;
        RECT 40.950 722.550 52.050 723.450 ;
        RECT 40.950 721.950 43.050 722.550 ;
        RECT 49.950 721.950 52.050 722.550 ;
        RECT 53.400 711.600 54.600 724.950 ;
        RECT 56.100 723.150 57.900 724.950 ;
        RECT 74.850 711.600 76.050 724.950 ;
        RECT 80.100 723.150 81.900 724.950 ;
        RECT 95.400 711.600 96.600 724.950 ;
        RECT 98.100 723.150 99.900 724.950 ;
        RECT 14.400 705.600 16.200 711.600 ;
        RECT 35.400 705.600 37.200 711.600 ;
        RECT 52.800 705.600 54.600 711.600 ;
        RECT 74.400 705.600 76.200 711.600 ;
        RECT 94.800 705.600 96.600 711.600 ;
        RECT 101.550 717.600 102.750 724.950 ;
        RECT 103.950 719.400 105.750 721.200 ;
        RECT 104.850 718.200 109.050 719.400 ;
        RECT 114.150 718.200 115.050 730.800 ;
        RECT 125.100 729.600 132.000 730.800 ;
        RECT 125.100 729.000 126.900 729.600 ;
        RECT 131.100 728.850 132.000 729.600 ;
        RECT 128.100 727.800 129.900 728.400 ;
        RECT 121.950 726.600 129.900 727.800 ;
        RECT 131.100 727.050 132.900 728.850 ;
        RECT 121.950 724.950 124.050 726.600 ;
        RECT 130.950 724.950 133.050 727.050 ;
        RECT 123.750 719.700 125.550 720.000 ;
        RECT 133.950 719.700 134.850 734.400 ;
        RECT 149.400 732.300 150.600 734.400 ;
        RECT 151.800 735.300 153.600 740.400 ;
        RECT 157.800 735.300 159.600 740.400 ;
        RECT 151.800 733.950 159.600 735.300 ;
        RECT 161.550 734.400 163.350 740.400 ;
        RECT 169.650 737.400 171.450 740.400 ;
        RECT 177.450 737.400 179.250 740.400 ;
        RECT 185.250 738.300 187.050 740.400 ;
        RECT 185.250 737.400 189.000 738.300 ;
        RECT 169.650 736.500 170.700 737.400 ;
        RECT 166.950 735.300 170.700 736.500 ;
        RECT 178.200 736.500 179.250 737.400 ;
        RECT 187.950 736.500 189.000 737.400 ;
        RECT 178.200 735.450 183.150 736.500 ;
        RECT 166.950 734.400 169.050 735.300 ;
        RECT 181.350 734.700 183.150 735.450 ;
        RECT 149.400 731.250 153.150 732.300 ;
        RECT 149.100 727.050 150.900 728.850 ;
        RECT 151.950 727.050 153.150 731.250 ;
        RECT 155.100 727.050 156.900 728.850 ;
        RECT 161.550 727.050 162.750 734.400 ;
        RECT 184.650 733.800 186.450 735.600 ;
        RECT 187.950 734.400 190.050 736.500 ;
        RECT 193.050 734.400 194.850 740.400 ;
        RECT 212.700 735.600 214.500 740.400 ;
        RECT 174.150 732.000 175.950 732.600 ;
        RECT 185.100 732.000 186.150 733.800 ;
        RECT 174.150 730.800 186.150 732.000 ;
        RECT 148.950 724.950 151.050 727.050 ;
        RECT 151.950 724.950 154.050 727.050 ;
        RECT 154.950 724.950 157.050 727.050 ;
        RECT 157.950 724.950 160.050 727.050 ;
        RECT 161.550 725.250 167.850 727.050 ;
        RECT 161.550 724.950 166.050 725.250 ;
        RECT 123.750 719.100 134.850 719.700 ;
        RECT 101.550 705.600 103.350 717.600 ;
        RECT 106.950 717.300 109.050 718.200 ;
        RECT 109.950 717.300 115.050 718.200 ;
        RECT 117.150 718.500 134.850 719.100 ;
        RECT 117.150 718.200 125.550 718.500 ;
        RECT 109.950 716.400 110.850 717.300 ;
        RECT 108.150 714.600 110.850 716.400 ;
        RECT 111.750 716.100 113.550 716.400 ;
        RECT 117.150 716.100 118.050 718.200 ;
        RECT 133.950 717.600 134.850 718.500 ;
        RECT 111.750 715.200 118.050 716.100 ;
        RECT 118.950 716.700 120.750 717.300 ;
        RECT 118.950 715.500 126.450 716.700 ;
        RECT 111.750 714.600 113.550 715.200 ;
        RECT 125.250 714.600 126.450 715.500 ;
        RECT 106.950 711.600 110.850 713.700 ;
        RECT 115.950 713.550 117.750 714.300 ;
        RECT 120.750 713.550 122.550 714.300 ;
        RECT 115.950 712.500 122.550 713.550 ;
        RECT 125.250 712.500 130.050 714.600 ;
        RECT 109.050 705.600 110.850 711.600 ;
        RECT 116.850 705.600 118.650 712.500 ;
        RECT 125.250 711.600 126.450 712.500 ;
        RECT 124.650 705.600 126.450 711.600 ;
        RECT 133.050 705.600 134.850 717.600 ;
        RECT 152.850 711.600 154.050 724.950 ;
        RECT 158.100 723.150 159.900 724.950 ;
        RECT 161.550 717.600 162.750 724.950 ;
        RECT 163.950 719.400 165.750 721.200 ;
        RECT 164.850 718.200 169.050 719.400 ;
        RECT 174.150 718.200 175.050 730.800 ;
        RECT 185.100 729.600 192.000 730.800 ;
        RECT 185.100 729.000 186.900 729.600 ;
        RECT 191.100 728.850 192.000 729.600 ;
        RECT 188.100 727.800 189.900 728.400 ;
        RECT 181.950 726.600 189.900 727.800 ;
        RECT 191.100 727.050 192.900 728.850 ;
        RECT 181.950 724.950 184.050 726.600 ;
        RECT 190.950 724.950 193.050 727.050 ;
        RECT 183.750 719.700 185.550 720.000 ;
        RECT 193.950 719.700 194.850 734.400 ;
        RECT 209.400 734.400 214.500 735.600 ;
        RECT 232.800 734.400 234.600 740.400 ;
        RECT 209.400 727.050 210.300 734.400 ;
        RECT 233.400 732.300 234.600 734.400 ;
        RECT 235.800 735.300 237.600 740.400 ;
        RECT 241.800 735.300 243.600 740.400 ;
        RECT 235.800 733.950 243.600 735.300 ;
        RECT 254.400 735.300 256.200 740.400 ;
        RECT 260.400 735.300 262.200 740.400 ;
        RECT 254.400 733.950 262.200 735.300 ;
        RECT 263.400 734.400 265.200 740.400 ;
        RECT 284.700 735.600 286.500 740.400 ;
        RECT 281.400 734.400 286.500 735.600 ;
        RECT 263.400 732.300 264.600 734.400 ;
        RECT 233.400 731.250 237.150 732.300 ;
        RECT 212.100 727.050 213.900 728.850 ;
        RECT 218.100 727.050 219.900 728.850 ;
        RECT 233.100 727.050 234.900 728.850 ;
        RECT 235.950 727.050 237.150 731.250 ;
        RECT 260.850 731.250 264.600 732.300 ;
        RECT 239.100 727.050 240.900 728.850 ;
        RECT 257.100 727.050 258.900 728.850 ;
        RECT 260.850 727.050 262.050 731.250 ;
        RECT 263.100 727.050 264.900 728.850 ;
        RECT 281.400 727.050 282.300 734.400 ;
        RECT 307.200 732.000 309.000 740.400 ;
        RECT 305.700 730.800 309.000 732.000 ;
        RECT 329.400 737.400 331.200 740.400 ;
        RECT 284.100 727.050 285.900 728.850 ;
        RECT 290.100 727.050 291.900 728.850 ;
        RECT 305.700 727.050 306.600 730.800 ;
        RECT 308.100 727.050 309.900 728.850 ;
        RECT 314.100 727.050 315.900 728.850 ;
        RECT 329.400 727.050 330.600 737.400 ;
        RECT 349.500 735.600 351.300 740.400 ;
        RECT 349.500 734.400 354.600 735.600 ;
        RECT 344.100 727.050 345.900 728.850 ;
        RECT 350.100 727.050 351.900 728.850 ;
        RECT 353.700 727.050 354.600 734.400 ;
        RECT 368.400 735.300 370.200 740.400 ;
        RECT 374.400 735.300 376.200 740.400 ;
        RECT 368.400 733.950 376.200 735.300 ;
        RECT 377.400 734.400 379.200 740.400 ;
        RECT 395.400 737.400 397.200 740.400 ;
        RECT 377.400 732.300 378.600 734.400 ;
        RECT 374.850 731.250 378.600 732.300 ;
        RECT 371.100 727.050 372.900 728.850 ;
        RECT 374.850 727.050 376.050 731.250 ;
        RECT 377.100 727.050 378.900 728.850 ;
        RECT 395.700 727.050 396.600 737.400 ;
        RECT 418.800 733.200 420.600 740.400 ;
        RECT 416.400 732.300 420.600 733.200 ;
        RECT 436.800 734.400 438.600 740.400 ;
        RECT 442.800 737.400 444.600 740.400 ;
        RECT 413.100 727.050 414.900 728.850 ;
        RECT 416.400 727.050 417.600 732.300 ;
        RECT 419.100 727.050 420.900 728.850 ;
        RECT 436.800 727.050 438.000 734.400 ;
        RECT 443.400 733.500 444.600 737.400 ;
        RECT 457.800 734.400 459.600 740.400 ;
        RECT 438.900 732.600 444.600 733.500 ;
        RECT 438.900 731.700 440.850 732.600 ;
        RECT 208.950 724.950 211.050 727.050 ;
        RECT 211.950 724.950 214.050 727.050 ;
        RECT 214.950 724.950 217.050 727.050 ;
        RECT 217.950 724.950 220.050 727.050 ;
        RECT 232.950 724.950 235.050 727.050 ;
        RECT 235.950 724.950 238.050 727.050 ;
        RECT 238.950 724.950 241.050 727.050 ;
        RECT 241.950 724.950 244.050 727.050 ;
        RECT 253.950 724.950 256.050 727.050 ;
        RECT 256.950 724.950 259.050 727.050 ;
        RECT 259.950 724.950 262.050 727.050 ;
        RECT 262.950 724.950 265.050 727.050 ;
        RECT 280.950 724.950 283.050 727.050 ;
        RECT 283.950 724.950 286.050 727.050 ;
        RECT 286.950 724.950 289.050 727.050 ;
        RECT 289.950 724.950 292.050 727.050 ;
        RECT 304.950 724.950 307.050 727.050 ;
        RECT 307.950 724.950 310.050 727.050 ;
        RECT 310.950 724.950 313.050 727.050 ;
        RECT 313.950 724.950 316.050 727.050 ;
        RECT 325.950 724.950 328.050 727.050 ;
        RECT 328.950 724.950 331.050 727.050 ;
        RECT 343.950 724.950 346.050 727.050 ;
        RECT 346.950 724.950 349.050 727.050 ;
        RECT 349.950 724.950 352.050 727.050 ;
        RECT 352.950 724.950 355.050 727.050 ;
        RECT 367.950 724.950 370.050 727.050 ;
        RECT 370.950 724.950 373.050 727.050 ;
        RECT 373.950 724.950 376.050 727.050 ;
        RECT 376.950 724.950 379.050 727.050 ;
        RECT 391.950 724.950 394.050 727.050 ;
        RECT 394.950 724.950 397.050 727.050 ;
        RECT 397.950 724.950 400.050 727.050 ;
        RECT 412.950 724.950 415.050 727.050 ;
        RECT 415.950 724.950 418.050 727.050 ;
        RECT 418.950 724.950 421.050 727.050 ;
        RECT 436.800 724.950 439.050 727.050 ;
        RECT 183.750 719.100 194.850 719.700 ;
        RECT 152.400 705.600 154.200 711.600 ;
        RECT 161.550 705.600 163.350 717.600 ;
        RECT 166.950 717.300 169.050 718.200 ;
        RECT 169.950 717.300 175.050 718.200 ;
        RECT 177.150 718.500 194.850 719.100 ;
        RECT 177.150 718.200 185.550 718.500 ;
        RECT 169.950 716.400 170.850 717.300 ;
        RECT 168.150 714.600 170.850 716.400 ;
        RECT 171.750 716.100 173.550 716.400 ;
        RECT 177.150 716.100 178.050 718.200 ;
        RECT 193.950 717.600 194.850 718.500 ;
        RECT 209.400 717.600 210.300 724.950 ;
        RECT 215.100 723.150 216.900 724.950 ;
        RECT 171.750 715.200 178.050 716.100 ;
        RECT 178.950 716.700 180.750 717.300 ;
        RECT 178.950 715.500 186.450 716.700 ;
        RECT 171.750 714.600 173.550 715.200 ;
        RECT 185.250 714.600 186.450 715.500 ;
        RECT 166.950 711.600 170.850 713.700 ;
        RECT 175.950 713.550 177.750 714.300 ;
        RECT 180.750 713.550 182.550 714.300 ;
        RECT 175.950 712.500 182.550 713.550 ;
        RECT 185.250 712.500 190.050 714.600 ;
        RECT 169.050 705.600 170.850 711.600 ;
        RECT 176.850 705.600 178.650 712.500 ;
        RECT 185.250 711.600 186.450 712.500 ;
        RECT 184.650 705.600 186.450 711.600 ;
        RECT 193.050 705.600 194.850 717.600 ;
        RECT 208.800 705.600 210.600 717.600 ;
        RECT 211.800 716.700 219.600 717.600 ;
        RECT 211.800 705.600 213.600 716.700 ;
        RECT 217.800 705.600 219.600 716.700 ;
        RECT 236.850 711.600 238.050 724.950 ;
        RECT 242.100 723.150 243.900 724.950 ;
        RECT 254.100 723.150 255.900 724.950 ;
        RECT 259.950 711.600 261.150 724.950 ;
        RECT 281.400 717.600 282.300 724.950 ;
        RECT 287.100 723.150 288.900 724.950 ;
        RECT 236.400 705.600 238.200 711.600 ;
        RECT 259.800 705.600 261.600 711.600 ;
        RECT 280.800 705.600 282.600 717.600 ;
        RECT 283.800 716.700 291.600 717.600 ;
        RECT 283.800 705.600 285.600 716.700 ;
        RECT 289.800 705.600 291.600 716.700 ;
        RECT 305.700 712.800 306.600 724.950 ;
        RECT 311.100 723.150 312.900 724.950 ;
        RECT 326.100 723.150 327.900 724.950 ;
        RECT 307.950 720.450 310.050 721.050 ;
        RECT 319.950 720.450 322.050 721.050 ;
        RECT 307.950 719.550 322.050 720.450 ;
        RECT 307.950 718.950 310.050 719.550 ;
        RECT 319.950 718.950 322.050 719.550 ;
        RECT 305.700 711.900 312.300 712.800 ;
        RECT 305.700 711.600 306.600 711.900 ;
        RECT 304.800 705.600 306.600 711.600 ;
        RECT 310.800 711.600 312.300 711.900 ;
        RECT 329.400 711.600 330.600 724.950 ;
        RECT 347.100 723.150 348.900 724.950 ;
        RECT 353.700 717.600 354.600 724.950 ;
        RECT 368.100 723.150 369.900 724.950 ;
        RECT 344.400 716.700 352.200 717.600 ;
        RECT 310.800 705.600 312.600 711.600 ;
        RECT 329.400 705.600 331.200 711.600 ;
        RECT 344.400 705.600 346.200 716.700 ;
        RECT 350.400 705.600 352.200 716.700 ;
        RECT 353.400 705.600 355.200 717.600 ;
        RECT 373.950 711.600 375.150 724.950 ;
        RECT 392.100 723.150 393.900 724.950 ;
        RECT 395.700 717.600 396.600 724.950 ;
        RECT 398.100 723.150 399.900 724.950 ;
        RECT 395.700 716.400 399.300 717.600 ;
        RECT 373.800 705.600 375.600 711.600 ;
        RECT 397.500 705.600 399.300 716.400 ;
        RECT 416.400 711.600 417.600 724.950 ;
        RECT 436.800 717.600 438.000 724.950 ;
        RECT 439.950 720.300 440.850 731.700 ;
        RECT 458.400 732.300 459.600 734.400 ;
        RECT 460.800 735.300 462.600 740.400 ;
        RECT 466.800 735.300 468.600 740.400 ;
        RECT 481.800 737.400 483.600 740.400 ;
        RECT 460.800 733.950 468.600 735.300 ;
        RECT 458.400 731.250 462.150 732.300 ;
        RECT 458.100 727.050 459.900 728.850 ;
        RECT 460.950 727.050 462.150 731.250 ;
        RECT 464.100 727.050 465.900 728.850 ;
        RECT 482.400 727.050 483.600 737.400 ;
        RECT 500.400 733.200 502.200 740.400 ;
        RECT 523.800 733.200 525.600 740.400 ;
        RECT 544.800 733.200 546.600 740.400 ;
        RECT 565.800 733.200 567.600 740.400 ;
        RECT 585.300 736.200 587.100 740.400 ;
        RECT 500.400 732.300 504.600 733.200 ;
        RECT 500.100 727.050 501.900 728.850 ;
        RECT 503.400 727.050 504.600 732.300 ;
        RECT 521.400 732.300 525.600 733.200 ;
        RECT 542.400 732.300 546.600 733.200 ;
        RECT 563.400 732.300 567.600 733.200 ;
        RECT 584.400 734.400 587.100 736.200 ;
        RECT 506.100 727.050 507.900 728.850 ;
        RECT 518.100 727.050 519.900 728.850 ;
        RECT 521.400 727.050 522.600 732.300 ;
        RECT 524.100 727.050 525.900 728.850 ;
        RECT 539.100 727.050 540.900 728.850 ;
        RECT 542.400 727.050 543.600 732.300 ;
        RECT 545.100 727.050 546.900 728.850 ;
        RECT 560.100 727.050 561.900 728.850 ;
        RECT 563.400 727.050 564.600 732.300 ;
        RECT 566.100 727.050 567.900 728.850 ;
        RECT 584.400 727.050 585.300 734.400 ;
        RECT 587.100 732.600 588.900 733.500 ;
        RECT 592.800 732.600 594.600 740.400 ;
        RECT 605.400 735.300 607.200 740.400 ;
        RECT 611.400 735.300 613.200 740.400 ;
        RECT 605.400 733.950 613.200 735.300 ;
        RECT 614.400 734.400 616.200 740.400 ;
        RECT 633.300 736.200 635.100 740.400 ;
        RECT 632.400 734.400 635.100 736.200 ;
        RECT 587.100 731.700 594.600 732.600 ;
        RECT 614.400 732.300 615.600 734.400 ;
        RECT 442.950 724.950 445.050 727.050 ;
        RECT 457.950 724.950 460.050 727.050 ;
        RECT 460.950 724.950 463.050 727.050 ;
        RECT 463.950 724.950 466.050 727.050 ;
        RECT 466.950 724.950 469.050 727.050 ;
        RECT 481.950 724.950 484.050 727.050 ;
        RECT 484.950 724.950 487.050 727.050 ;
        RECT 499.950 724.950 502.050 727.050 ;
        RECT 502.950 724.950 505.050 727.050 ;
        RECT 505.950 724.950 508.050 727.050 ;
        RECT 517.950 724.950 520.050 727.050 ;
        RECT 520.950 724.950 523.050 727.050 ;
        RECT 523.950 724.950 526.050 727.050 ;
        RECT 538.950 724.950 541.050 727.050 ;
        RECT 541.950 724.950 544.050 727.050 ;
        RECT 544.950 724.950 547.050 727.050 ;
        RECT 559.950 724.950 562.050 727.050 ;
        RECT 562.950 724.950 565.050 727.050 ;
        RECT 565.950 724.950 568.050 727.050 ;
        RECT 583.950 724.950 586.050 727.050 ;
        RECT 586.950 724.950 589.050 727.050 ;
        RECT 443.100 723.150 444.900 724.950 ;
        RECT 438.900 719.400 440.850 720.300 ;
        RECT 438.900 718.500 444.600 719.400 ;
        RECT 416.400 705.600 418.200 711.600 ;
        RECT 436.800 705.600 438.600 717.600 ;
        RECT 443.400 711.600 444.600 718.500 ;
        RECT 461.850 711.600 463.050 724.950 ;
        RECT 467.100 723.150 468.900 724.950 ;
        RECT 482.400 711.600 483.600 724.950 ;
        RECT 485.100 723.150 486.900 724.950 ;
        RECT 503.400 711.600 504.600 724.950 ;
        RECT 442.800 705.600 444.600 711.600 ;
        RECT 461.400 705.600 463.200 711.600 ;
        RECT 481.800 705.600 483.600 711.600 ;
        RECT 502.800 705.600 504.600 711.600 ;
        RECT 521.400 711.600 522.600 724.950 ;
        RECT 542.400 711.600 543.600 724.950 ;
        RECT 563.400 711.600 564.600 724.950 ;
        RECT 584.400 717.600 585.300 724.950 ;
        RECT 587.100 723.150 588.900 724.950 ;
        RECT 521.400 705.600 523.200 711.600 ;
        RECT 542.400 705.600 544.200 711.600 ;
        RECT 563.400 705.600 565.200 711.600 ;
        RECT 583.800 705.600 585.600 717.600 ;
        RECT 590.700 711.600 591.600 731.700 ;
        RECT 611.850 731.250 615.600 732.300 ;
        RECT 593.100 727.050 594.900 728.850 ;
        RECT 608.100 727.050 609.900 728.850 ;
        RECT 611.850 727.050 613.050 731.250 ;
        RECT 614.100 727.050 615.900 728.850 ;
        RECT 632.400 727.050 633.300 734.400 ;
        RECT 635.100 732.600 636.900 733.500 ;
        RECT 640.800 732.600 642.600 740.400 ;
        RECT 658.800 733.200 660.600 740.400 ;
        RECT 680.700 735.600 682.500 740.400 ;
        RECT 635.100 731.700 642.600 732.600 ;
        RECT 656.400 732.300 660.600 733.200 ;
        RECT 677.400 734.400 682.500 735.600 ;
        RECT 592.950 724.950 595.050 727.050 ;
        RECT 604.950 724.950 607.050 727.050 ;
        RECT 607.950 724.950 610.050 727.050 ;
        RECT 610.950 724.950 613.050 727.050 ;
        RECT 613.950 724.950 616.050 727.050 ;
        RECT 631.950 724.950 634.050 727.050 ;
        RECT 634.950 724.950 637.050 727.050 ;
        RECT 605.100 723.150 606.900 724.950 ;
        RECT 610.950 711.600 612.150 724.950 ;
        RECT 632.400 717.600 633.300 724.950 ;
        RECT 635.100 723.150 636.900 724.950 ;
        RECT 589.800 705.600 591.600 711.600 ;
        RECT 610.800 705.600 612.600 711.600 ;
        RECT 631.800 705.600 633.600 717.600 ;
        RECT 638.700 711.600 639.600 731.700 ;
        RECT 641.100 727.050 642.900 728.850 ;
        RECT 653.100 727.050 654.900 728.850 ;
        RECT 656.400 727.050 657.600 732.300 ;
        RECT 659.100 727.050 660.900 728.850 ;
        RECT 677.400 727.050 678.300 734.400 ;
        RECT 705.000 732.000 706.800 740.400 ;
        RECT 724.800 734.400 726.600 740.400 ;
        RECT 725.400 732.300 726.600 734.400 ;
        RECT 727.800 735.300 729.600 740.400 ;
        RECT 733.800 735.300 735.600 740.400 ;
        RECT 727.800 733.950 735.600 735.300 ;
        RECT 751.800 733.200 753.600 740.400 ;
        RECT 749.400 732.300 753.600 733.200 ;
        RECT 770.400 737.400 772.200 740.400 ;
        RECT 705.000 730.800 708.300 732.000 ;
        RECT 725.400 731.250 729.150 732.300 ;
        RECT 680.100 727.050 681.900 728.850 ;
        RECT 686.100 727.050 687.900 728.850 ;
        RECT 698.100 727.050 699.900 728.850 ;
        RECT 704.100 727.050 705.900 728.850 ;
        RECT 707.400 727.050 708.300 730.800 ;
        RECT 725.100 727.050 726.900 728.850 ;
        RECT 727.950 727.050 729.150 731.250 ;
        RECT 731.100 727.050 732.900 728.850 ;
        RECT 746.100 727.050 747.900 728.850 ;
        RECT 749.400 727.050 750.600 732.300 ;
        RECT 752.100 727.050 753.900 728.850 ;
        RECT 770.400 727.050 771.600 737.400 ;
        RECT 790.200 732.000 792.000 740.400 ;
        RECT 814.500 735.600 816.300 740.400 ;
        RECT 814.500 734.400 819.600 735.600 ;
        RECT 788.700 730.800 792.000 732.000 ;
        RECT 788.700 727.050 789.600 730.800 ;
        RECT 791.100 727.050 792.900 728.850 ;
        RECT 797.100 727.050 798.900 728.850 ;
        RECT 809.100 727.050 810.900 728.850 ;
        RECT 815.100 727.050 816.900 728.850 ;
        RECT 818.700 727.050 819.600 734.400 ;
        RECT 843.000 732.000 844.800 740.400 ;
        RECT 860.400 735.300 862.200 740.400 ;
        RECT 866.400 735.300 868.200 740.400 ;
        RECT 860.400 733.950 868.200 735.300 ;
        RECT 869.400 734.400 871.200 740.400 ;
        RECT 869.400 732.300 870.600 734.400 ;
        RECT 843.000 730.800 846.300 732.000 ;
        RECT 836.100 727.050 837.900 728.850 ;
        RECT 842.100 727.050 843.900 728.850 ;
        RECT 845.400 727.050 846.300 730.800 ;
        RECT 866.850 731.250 870.600 732.300 ;
        RECT 847.950 729.450 852.000 730.050 ;
        RECT 855.000 729.450 859.050 730.050 ;
        RECT 847.950 727.950 852.450 729.450 ;
        RECT 640.950 724.950 643.050 727.050 ;
        RECT 652.950 724.950 655.050 727.050 ;
        RECT 655.950 724.950 658.050 727.050 ;
        RECT 658.950 724.950 661.050 727.050 ;
        RECT 676.950 724.950 679.050 727.050 ;
        RECT 679.950 724.950 682.050 727.050 ;
        RECT 682.950 724.950 685.050 727.050 ;
        RECT 685.950 724.950 688.050 727.050 ;
        RECT 697.950 724.950 700.050 727.050 ;
        RECT 700.950 724.950 703.050 727.050 ;
        RECT 703.950 724.950 706.050 727.050 ;
        RECT 706.950 724.950 709.050 727.050 ;
        RECT 724.950 724.950 727.050 727.050 ;
        RECT 727.950 724.950 730.050 727.050 ;
        RECT 730.950 724.950 733.050 727.050 ;
        RECT 733.950 724.950 736.050 727.050 ;
        RECT 745.950 724.950 748.050 727.050 ;
        RECT 748.950 724.950 751.050 727.050 ;
        RECT 751.950 724.950 754.050 727.050 ;
        RECT 766.950 724.950 769.050 727.050 ;
        RECT 769.950 724.950 772.050 727.050 ;
        RECT 787.950 724.950 790.050 727.050 ;
        RECT 790.950 724.950 793.050 727.050 ;
        RECT 793.950 724.950 796.050 727.050 ;
        RECT 796.950 724.950 799.050 727.050 ;
        RECT 808.950 724.950 811.050 727.050 ;
        RECT 811.950 724.950 814.050 727.050 ;
        RECT 814.950 724.950 817.050 727.050 ;
        RECT 817.950 724.950 820.050 727.050 ;
        RECT 835.950 724.950 838.050 727.050 ;
        RECT 838.950 724.950 841.050 727.050 ;
        RECT 841.950 724.950 844.050 727.050 ;
        RECT 844.950 724.950 847.050 727.050 ;
        RECT 640.950 717.450 643.050 718.050 ;
        RECT 652.950 717.450 655.050 718.050 ;
        RECT 640.950 716.550 655.050 717.450 ;
        RECT 640.950 715.950 643.050 716.550 ;
        RECT 652.950 715.950 655.050 716.550 ;
        RECT 637.800 705.600 639.600 711.600 ;
        RECT 656.400 711.600 657.600 724.950 ;
        RECT 677.400 717.600 678.300 724.950 ;
        RECT 683.100 723.150 684.900 724.950 ;
        RECT 701.100 723.150 702.900 724.950 ;
        RECT 656.400 705.600 658.200 711.600 ;
        RECT 676.800 705.600 678.600 717.600 ;
        RECT 679.800 716.700 687.600 717.600 ;
        RECT 679.800 705.600 681.600 716.700 ;
        RECT 685.800 705.600 687.600 716.700 ;
        RECT 707.400 712.800 708.300 724.950 ;
        RECT 701.700 711.900 708.300 712.800 ;
        RECT 701.700 711.600 703.200 711.900 ;
        RECT 701.400 705.600 703.200 711.600 ;
        RECT 707.400 711.600 708.300 711.900 ;
        RECT 728.850 711.600 730.050 724.950 ;
        RECT 734.100 723.150 735.900 724.950 ;
        RECT 749.400 711.600 750.600 724.950 ;
        RECT 767.100 723.150 768.900 724.950 ;
        RECT 770.400 711.600 771.600 724.950 ;
        RECT 788.700 712.800 789.600 724.950 ;
        RECT 794.100 723.150 795.900 724.950 ;
        RECT 812.100 723.150 813.900 724.950 ;
        RECT 796.950 720.450 799.050 721.050 ;
        RECT 814.950 720.450 817.050 721.050 ;
        RECT 796.950 719.550 817.050 720.450 ;
        RECT 796.950 718.950 799.050 719.550 ;
        RECT 814.950 718.950 817.050 719.550 ;
        RECT 818.700 717.600 819.600 724.950 ;
        RECT 839.100 723.150 840.900 724.950 ;
        RECT 809.400 716.700 817.200 717.600 ;
        RECT 788.700 711.900 795.300 712.800 ;
        RECT 788.700 711.600 789.600 711.900 ;
        RECT 707.400 705.600 709.200 711.600 ;
        RECT 728.400 705.600 730.200 711.600 ;
        RECT 749.400 705.600 751.200 711.600 ;
        RECT 770.400 705.600 772.200 711.600 ;
        RECT 787.800 705.600 789.600 711.600 ;
        RECT 793.800 711.600 795.300 711.900 ;
        RECT 793.800 705.600 795.600 711.600 ;
        RECT 809.400 705.600 811.200 716.700 ;
        RECT 815.400 705.600 817.200 716.700 ;
        RECT 818.400 705.600 820.200 717.600 ;
        RECT 845.400 712.800 846.300 724.950 ;
        RECT 851.550 720.450 852.450 727.950 ;
        RECT 854.550 727.950 859.050 729.450 ;
        RECT 854.550 724.050 855.450 727.950 ;
        RECT 863.100 727.050 864.900 728.850 ;
        RECT 866.850 727.050 868.050 731.250 ;
        RECT 869.100 727.050 870.900 728.850 ;
        RECT 859.950 724.950 862.050 727.050 ;
        RECT 862.950 724.950 865.050 727.050 ;
        RECT 865.950 724.950 868.050 727.050 ;
        RECT 868.950 724.950 871.050 727.050 ;
        RECT 854.550 722.550 859.050 724.050 ;
        RECT 860.100 723.150 861.900 724.950 ;
        RECT 855.000 721.950 859.050 722.550 ;
        RECT 859.950 720.450 862.050 721.050 ;
        RECT 851.550 719.550 862.050 720.450 ;
        RECT 859.950 718.950 862.050 719.550 ;
        RECT 839.700 711.900 846.300 712.800 ;
        RECT 839.700 711.600 841.200 711.900 ;
        RECT 839.400 705.600 841.200 711.600 ;
        RECT 845.400 711.600 846.300 711.900 ;
        RECT 865.950 711.600 867.150 724.950 ;
        RECT 871.950 723.450 874.050 724.050 ;
        RECT 889.950 723.450 892.050 724.050 ;
        RECT 871.950 722.550 892.050 723.450 ;
        RECT 871.950 721.950 874.050 722.550 ;
        RECT 889.950 721.950 892.050 722.550 ;
        RECT 845.400 705.600 847.200 711.600 ;
        RECT 865.800 705.600 867.600 711.600 ;
        RECT 17.400 695.400 19.200 701.400 ;
        RECT 40.800 695.400 42.600 701.400 ;
        RECT 17.850 682.050 19.050 695.400 ;
        RECT 22.950 687.450 25.050 688.050 ;
        RECT 22.950 686.550 30.450 687.450 ;
        RECT 22.950 685.950 25.050 686.550 ;
        RECT 23.100 682.050 24.900 683.850 ;
        RECT 13.950 679.950 16.050 682.050 ;
        RECT 16.950 679.950 19.050 682.050 ;
        RECT 19.950 679.950 22.050 682.050 ;
        RECT 22.950 679.950 25.050 682.050 ;
        RECT 14.100 678.150 15.900 679.950 ;
        RECT 16.950 675.750 18.150 679.950 ;
        RECT 20.100 678.150 21.900 679.950 ;
        RECT 29.550 679.050 30.450 686.550 ;
        RECT 35.100 682.050 36.900 683.850 ;
        RECT 40.950 682.050 42.150 695.400 ;
        RECT 61.800 689.400 63.600 701.400 ;
        RECT 67.800 695.400 69.600 701.400 ;
        RECT 46.950 684.450 49.050 685.050 ;
        RECT 55.950 684.450 58.050 685.050 ;
        RECT 46.950 683.550 58.050 684.450 ;
        RECT 46.950 682.950 49.050 683.550 ;
        RECT 55.950 682.950 58.050 683.550 ;
        RECT 62.400 682.050 63.300 689.400 ;
        RECT 65.100 682.050 66.900 683.850 ;
        RECT 34.950 679.950 37.050 682.050 ;
        RECT 37.950 679.950 40.050 682.050 ;
        RECT 40.950 679.950 43.050 682.050 ;
        RECT 43.950 679.950 46.050 682.050 ;
        RECT 61.950 679.950 64.050 682.050 ;
        RECT 64.950 679.950 67.050 682.050 ;
        RECT 29.550 677.550 34.050 679.050 ;
        RECT 38.100 678.150 39.900 679.950 ;
        RECT 30.000 676.950 34.050 677.550 ;
        RECT 14.400 674.700 18.150 675.750 ;
        RECT 41.850 675.750 43.050 679.950 ;
        RECT 44.100 678.150 45.900 679.950 ;
        RECT 41.850 674.700 45.600 675.750 ;
        RECT 14.400 672.600 15.600 674.700 ;
        RECT 13.800 666.600 15.600 672.600 ;
        RECT 16.800 671.700 24.600 673.050 ;
        RECT 16.800 666.600 18.600 671.700 ;
        RECT 22.800 666.600 24.600 671.700 ;
        RECT 35.400 671.700 43.200 673.050 ;
        RECT 35.400 666.600 37.200 671.700 ;
        RECT 41.400 666.600 43.200 671.700 ;
        RECT 44.400 672.600 45.600 674.700 ;
        RECT 62.400 672.600 63.300 679.950 ;
        RECT 68.700 675.300 69.600 695.400 ;
        RECT 90.300 690.900 92.100 701.400 ;
        RECT 89.700 689.400 92.100 690.900 ;
        RECT 97.800 689.400 99.600 701.400 ;
        RECT 89.700 682.050 91.050 689.400 ;
        RECT 98.400 687.900 99.600 689.400 ;
        RECT 70.950 679.950 73.050 682.050 ;
        RECT 88.950 679.950 91.050 682.050 ;
        RECT 92.400 686.700 99.600 687.900 ;
        RECT 113.400 695.400 115.200 701.400 ;
        RECT 134.400 695.400 136.200 701.400 ;
        RECT 92.400 686.100 94.200 686.700 ;
        RECT 71.100 678.150 72.900 679.950 ;
        RECT 65.100 674.400 72.600 675.300 ;
        RECT 65.100 673.500 66.900 674.400 ;
        RECT 44.400 666.600 46.200 672.600 ;
        RECT 62.400 670.800 65.100 672.600 ;
        RECT 63.300 666.600 65.100 670.800 ;
        RECT 70.800 666.600 72.600 674.400 ;
        RECT 88.950 672.600 90.000 679.950 ;
        RECT 92.400 675.600 93.300 686.100 ;
        RECT 95.100 682.050 96.900 683.850 ;
        RECT 113.400 682.050 114.600 695.400 ;
        RECT 134.400 682.050 135.600 695.400 ;
        RECT 154.800 689.400 156.600 701.400 ;
        RECT 160.800 695.400 162.600 701.400 ;
        RECT 175.800 695.400 177.600 701.400 ;
        RECT 193.800 695.400 195.600 701.400 ;
        RECT 154.800 682.050 156.000 689.400 ;
        RECT 161.400 688.500 162.600 695.400 ;
        RECT 156.900 687.600 162.600 688.500 ;
        RECT 156.900 686.700 158.850 687.600 ;
        RECT 94.950 679.950 97.050 682.050 ;
        RECT 97.950 679.950 100.050 682.050 ;
        RECT 109.950 679.950 112.050 682.050 ;
        RECT 112.950 679.950 115.050 682.050 ;
        RECT 115.950 679.950 118.050 682.050 ;
        RECT 130.950 679.950 133.050 682.050 ;
        RECT 133.950 679.950 136.050 682.050 ;
        RECT 136.950 679.950 139.050 682.050 ;
        RECT 154.800 679.950 157.050 682.050 ;
        RECT 98.100 678.150 99.900 679.950 ;
        RECT 110.100 678.150 111.900 679.950 ;
        RECT 92.400 674.700 94.200 675.600 ;
        RECT 113.400 674.700 114.600 679.950 ;
        RECT 116.100 678.150 117.900 679.950 ;
        RECT 131.100 678.150 132.900 679.950 ;
        RECT 134.400 674.700 135.600 679.950 ;
        RECT 137.100 678.150 138.900 679.950 ;
        RECT 92.400 673.800 95.700 674.700 ;
        RECT 113.400 673.800 117.600 674.700 ;
        RECT 134.400 673.800 138.600 674.700 ;
        RECT 88.800 666.600 90.600 672.600 ;
        RECT 94.800 669.600 95.700 673.800 ;
        RECT 94.800 666.600 96.600 669.600 ;
        RECT 115.800 666.600 117.600 673.800 ;
        RECT 118.950 669.450 121.050 670.050 ;
        RECT 127.950 669.450 130.050 670.050 ;
        RECT 118.950 668.550 130.050 669.450 ;
        RECT 118.950 667.950 121.050 668.550 ;
        RECT 127.950 667.950 130.050 668.550 ;
        RECT 136.800 666.600 138.600 673.800 ;
        RECT 154.800 672.600 156.000 679.950 ;
        RECT 157.950 675.300 158.850 686.700 ;
        RECT 161.100 682.050 162.900 683.850 ;
        RECT 176.400 682.050 177.600 695.400 ;
        RECT 194.700 695.100 195.600 695.400 ;
        RECT 199.800 695.400 201.600 701.400 ;
        RECT 199.800 695.100 201.300 695.400 ;
        RECT 194.700 694.200 201.300 695.100 ;
        RECT 179.100 682.050 180.900 683.850 ;
        RECT 194.700 682.050 195.600 694.200 ;
        RECT 215.400 690.300 217.200 701.400 ;
        RECT 221.400 690.300 223.200 701.400 ;
        RECT 215.400 689.400 223.200 690.300 ;
        RECT 224.400 689.400 226.200 701.400 ;
        RECT 245.400 695.400 247.200 701.400 ;
        RECT 196.950 687.450 199.050 688.050 ;
        RECT 196.950 686.550 207.450 687.450 ;
        RECT 196.950 685.950 199.050 686.550 ;
        RECT 206.550 684.450 207.450 686.550 ;
        RECT 200.100 682.050 201.900 683.850 ;
        RECT 206.550 683.550 210.450 684.450 ;
        RECT 160.950 679.950 163.050 682.050 ;
        RECT 175.950 679.950 178.050 682.050 ;
        RECT 178.950 679.950 181.050 682.050 ;
        RECT 193.950 679.950 196.050 682.050 ;
        RECT 196.950 679.950 199.050 682.050 ;
        RECT 199.950 679.950 202.050 682.050 ;
        RECT 202.950 679.950 205.050 682.050 ;
        RECT 156.900 674.400 158.850 675.300 ;
        RECT 156.900 673.500 162.600 674.400 ;
        RECT 154.800 666.600 156.600 672.600 ;
        RECT 161.400 669.600 162.600 673.500 ;
        RECT 176.400 669.600 177.600 679.950 ;
        RECT 194.700 676.200 195.600 679.950 ;
        RECT 197.100 678.150 198.900 679.950 ;
        RECT 203.100 678.150 204.900 679.950 ;
        RECT 209.550 679.050 210.450 683.550 ;
        RECT 218.100 682.050 219.900 683.850 ;
        RECT 224.700 682.050 225.600 689.400 ;
        RECT 245.850 682.050 247.050 695.400 ;
        RECT 265.800 689.400 267.600 701.400 ;
        RECT 268.800 690.300 270.600 701.400 ;
        RECT 274.800 690.300 276.600 701.400 ;
        RECT 292.800 695.400 294.600 701.400 ;
        RECT 313.800 695.400 315.600 701.400 ;
        RECT 268.800 689.400 276.600 690.300 ;
        RECT 251.100 682.050 252.900 683.850 ;
        RECT 266.400 682.050 267.300 689.400 ;
        RECT 272.100 682.050 273.900 683.850 ;
        RECT 293.400 682.050 294.600 695.400 ;
        RECT 314.400 682.050 315.600 695.400 ;
        RECT 331.800 689.400 333.600 701.400 ;
        RECT 337.800 695.400 339.600 701.400 ;
        RECT 332.400 682.050 333.300 689.400 ;
        RECT 335.100 682.050 336.900 683.850 ;
        RECT 214.950 679.950 217.050 682.050 ;
        RECT 217.950 679.950 220.050 682.050 ;
        RECT 220.950 679.950 223.050 682.050 ;
        RECT 223.950 679.950 226.050 682.050 ;
        RECT 241.950 679.950 244.050 682.050 ;
        RECT 244.950 679.950 247.050 682.050 ;
        RECT 247.950 679.950 250.050 682.050 ;
        RECT 250.950 679.950 253.050 682.050 ;
        RECT 265.950 679.950 268.050 682.050 ;
        RECT 268.950 679.950 271.050 682.050 ;
        RECT 271.950 679.950 274.050 682.050 ;
        RECT 274.950 679.950 277.050 682.050 ;
        RECT 289.950 679.950 292.050 682.050 ;
        RECT 292.950 679.950 295.050 682.050 ;
        RECT 295.950 679.950 298.050 682.050 ;
        RECT 310.950 679.950 313.050 682.050 ;
        RECT 313.950 679.950 316.050 682.050 ;
        RECT 316.950 679.950 319.050 682.050 ;
        RECT 331.950 679.950 334.050 682.050 ;
        RECT 334.950 679.950 337.050 682.050 ;
        RECT 205.950 677.550 210.450 679.050 ;
        RECT 215.100 678.150 216.900 679.950 ;
        RECT 221.100 678.150 222.900 679.950 ;
        RECT 205.950 676.950 210.000 677.550 ;
        RECT 194.700 675.000 198.000 676.200 ;
        RECT 160.800 666.600 162.600 669.600 ;
        RECT 175.800 666.600 177.600 669.600 ;
        RECT 196.200 666.600 198.000 675.000 ;
        RECT 224.700 672.600 225.600 679.950 ;
        RECT 242.100 678.150 243.900 679.950 ;
        RECT 244.950 675.750 246.150 679.950 ;
        RECT 248.100 678.150 249.900 679.950 ;
        RECT 242.400 674.700 246.150 675.750 ;
        RECT 242.400 672.600 243.600 674.700 ;
        RECT 220.500 671.400 225.600 672.600 ;
        RECT 220.500 666.600 222.300 671.400 ;
        RECT 241.800 666.600 243.600 672.600 ;
        RECT 244.800 671.700 252.600 673.050 ;
        RECT 244.800 666.600 246.600 671.700 ;
        RECT 250.800 666.600 252.600 671.700 ;
        RECT 266.400 672.600 267.300 679.950 ;
        RECT 269.100 678.150 270.900 679.950 ;
        RECT 275.100 678.150 276.900 679.950 ;
        RECT 290.100 678.150 291.900 679.950 ;
        RECT 293.400 674.700 294.600 679.950 ;
        RECT 296.100 678.150 297.900 679.950 ;
        RECT 311.100 678.150 312.900 679.950 ;
        RECT 314.400 674.700 315.600 679.950 ;
        RECT 317.100 678.150 318.900 679.950 ;
        RECT 290.400 673.800 294.600 674.700 ;
        RECT 311.400 673.800 315.600 674.700 ;
        RECT 266.400 671.400 271.500 672.600 ;
        RECT 269.700 666.600 271.500 671.400 ;
        RECT 290.400 666.600 292.200 673.800 ;
        RECT 311.400 666.600 313.200 673.800 ;
        RECT 332.400 672.600 333.300 679.950 ;
        RECT 338.700 675.300 339.600 695.400 ;
        RECT 355.800 700.500 363.600 701.400 ;
        RECT 355.800 689.400 357.600 700.500 ;
        RECT 358.800 688.500 360.600 699.600 ;
        RECT 361.800 690.600 363.600 700.500 ;
        RECT 367.800 690.600 369.600 701.400 ;
        RECT 385.800 695.400 387.600 701.400 ;
        RECT 407.400 695.400 409.200 701.400 ;
        RECT 427.800 700.500 435.600 701.400 ;
        RECT 415.950 696.450 418.050 697.050 ;
        RECT 421.950 696.450 424.050 697.050 ;
        RECT 415.950 695.550 424.050 696.450 ;
        RECT 361.800 689.700 369.600 690.600 ;
        RECT 358.800 687.600 363.900 688.500 ;
        RECT 359.100 682.050 360.900 683.850 ;
        RECT 363.000 682.050 363.900 687.600 ;
        RECT 365.100 682.050 366.900 683.850 ;
        RECT 386.400 682.050 387.600 695.400 ;
        RECT 407.850 682.050 409.050 695.400 ;
        RECT 415.950 694.950 418.050 695.550 ;
        RECT 421.950 694.950 424.050 695.550 ;
        RECT 427.800 689.400 429.600 700.500 ;
        RECT 430.800 688.500 432.600 699.600 ;
        RECT 433.800 690.600 435.600 700.500 ;
        RECT 439.800 690.600 441.600 701.400 ;
        RECT 460.800 695.400 462.600 701.400 ;
        RECT 484.800 695.400 486.600 701.400 ;
        RECT 433.800 689.700 441.600 690.600 ;
        RECT 430.800 687.600 435.900 688.500 ;
        RECT 413.100 682.050 414.900 683.850 ;
        RECT 431.100 682.050 432.900 683.850 ;
        RECT 435.000 682.050 435.900 687.600 ;
        RECT 437.100 682.050 438.900 683.850 ;
        RECT 455.100 682.050 456.900 683.850 ;
        RECT 460.950 682.050 462.150 695.400 ;
        RECT 479.100 682.050 480.900 683.850 ;
        RECT 484.950 682.050 486.150 695.400 ;
        RECT 505.800 689.400 507.600 701.400 ;
        RECT 511.800 695.400 513.600 701.400 ;
        RECT 532.800 695.400 534.600 701.400 ;
        RECT 538.950 699.450 541.050 700.050 ;
        RECT 544.950 699.450 547.050 700.050 ;
        RECT 538.950 698.550 547.050 699.450 ;
        RECT 538.950 697.950 541.050 698.550 ;
        RECT 544.950 697.950 547.050 698.550 ;
        RECT 554.400 695.400 556.200 701.400 ;
        RECT 577.800 695.400 579.600 701.400 ;
        RECT 601.800 695.400 603.600 701.400 ;
        RECT 490.950 684.450 495.000 685.050 ;
        RECT 490.950 682.950 495.450 684.450 ;
        RECT 340.950 679.950 343.050 682.050 ;
        RECT 355.950 679.950 358.050 682.050 ;
        RECT 358.950 679.950 361.050 682.050 ;
        RECT 361.950 679.950 364.050 682.050 ;
        RECT 364.950 679.950 367.050 682.050 ;
        RECT 367.950 679.950 370.050 682.050 ;
        RECT 382.950 679.950 385.050 682.050 ;
        RECT 385.950 679.950 388.050 682.050 ;
        RECT 388.950 679.950 391.050 682.050 ;
        RECT 403.950 679.950 406.050 682.050 ;
        RECT 406.950 679.950 409.050 682.050 ;
        RECT 409.950 679.950 412.050 682.050 ;
        RECT 412.950 679.950 415.050 682.050 ;
        RECT 427.950 679.950 430.050 682.050 ;
        RECT 430.950 679.950 433.050 682.050 ;
        RECT 433.950 679.950 436.050 682.050 ;
        RECT 436.950 679.950 439.050 682.050 ;
        RECT 439.950 679.950 442.050 682.050 ;
        RECT 454.950 679.950 457.050 682.050 ;
        RECT 457.950 679.950 460.050 682.050 ;
        RECT 460.950 679.950 463.050 682.050 ;
        RECT 463.950 679.950 466.050 682.050 ;
        RECT 478.950 679.950 481.050 682.050 ;
        RECT 481.950 679.950 484.050 682.050 ;
        RECT 484.950 679.950 487.050 682.050 ;
        RECT 487.950 679.950 490.050 682.050 ;
        RECT 494.550 681.450 495.450 682.950 ;
        RECT 506.400 682.050 507.300 689.400 ;
        RECT 509.100 682.050 510.900 683.850 ;
        RECT 499.950 681.450 502.050 681.900 ;
        RECT 494.550 680.550 502.050 681.450 ;
        RECT 341.100 678.150 342.900 679.950 ;
        RECT 356.100 678.150 357.900 679.950 ;
        RECT 335.100 674.400 342.600 675.300 ;
        RECT 335.100 673.500 336.900 674.400 ;
        RECT 332.400 670.800 335.100 672.600 ;
        RECT 333.300 666.600 335.100 670.800 ;
        RECT 340.800 666.600 342.600 674.400 ;
        RECT 363.000 672.600 364.050 679.950 ;
        RECT 368.100 678.150 369.900 679.950 ;
        RECT 383.100 678.150 384.900 679.950 ;
        RECT 386.400 674.700 387.600 679.950 ;
        RECT 389.100 678.150 390.900 679.950 ;
        RECT 404.100 678.150 405.900 679.950 ;
        RECT 406.950 675.750 408.150 679.950 ;
        RECT 410.100 678.150 411.900 679.950 ;
        RECT 428.100 678.150 429.900 679.950 ;
        RECT 383.400 673.800 387.600 674.700 ;
        RECT 404.400 674.700 408.150 675.750 ;
        RECT 346.950 669.450 349.050 670.050 ;
        RECT 352.950 669.450 355.050 670.050 ;
        RECT 346.950 668.550 355.050 669.450 ;
        RECT 346.950 667.950 349.050 668.550 ;
        RECT 352.950 667.950 355.050 668.550 ;
        RECT 363.000 666.600 364.800 672.600 ;
        RECT 383.400 666.600 385.200 673.800 ;
        RECT 404.400 672.600 405.600 674.700 ;
        RECT 403.800 666.600 405.600 672.600 ;
        RECT 406.800 671.700 414.600 673.050 ;
        RECT 406.800 666.600 408.600 671.700 ;
        RECT 412.800 666.600 414.600 671.700 ;
        RECT 435.000 672.600 436.050 679.950 ;
        RECT 440.100 678.150 441.900 679.950 ;
        RECT 458.100 678.150 459.900 679.950 ;
        RECT 461.850 675.750 463.050 679.950 ;
        RECT 464.100 678.150 465.900 679.950 ;
        RECT 466.950 678.450 469.050 679.050 ;
        RECT 475.950 678.450 478.050 679.050 ;
        RECT 466.950 677.550 478.050 678.450 ;
        RECT 482.100 678.150 483.900 679.950 ;
        RECT 466.950 676.950 469.050 677.550 ;
        RECT 475.950 676.950 478.050 677.550 ;
        RECT 485.850 675.750 487.050 679.950 ;
        RECT 488.100 678.150 489.900 679.950 ;
        RECT 499.950 679.800 502.050 680.550 ;
        RECT 505.950 679.950 508.050 682.050 ;
        RECT 508.950 679.950 511.050 682.050 ;
        RECT 461.850 674.700 465.600 675.750 ;
        RECT 485.850 674.700 489.600 675.750 ;
        RECT 435.000 666.600 436.800 672.600 ;
        RECT 455.400 671.700 463.200 673.050 ;
        RECT 455.400 666.600 457.200 671.700 ;
        RECT 461.400 666.600 463.200 671.700 ;
        RECT 464.400 672.600 465.600 674.700 ;
        RECT 464.400 666.600 466.200 672.600 ;
        RECT 479.400 671.700 487.200 673.050 ;
        RECT 479.400 666.600 481.200 671.700 ;
        RECT 485.400 666.600 487.200 671.700 ;
        RECT 488.400 672.600 489.600 674.700 ;
        RECT 506.400 672.600 507.300 679.950 ;
        RECT 512.700 675.300 513.600 695.400 ;
        RECT 527.100 682.050 528.900 683.850 ;
        RECT 532.950 682.050 534.150 695.400 ;
        RECT 554.400 682.050 555.600 695.400 ;
        RECT 572.100 682.050 573.900 683.850 ;
        RECT 577.950 682.050 579.150 695.400 ;
        RECT 583.950 684.450 588.000 685.050 ;
        RECT 583.950 682.950 588.450 684.450 ;
        RECT 514.950 679.950 517.050 682.050 ;
        RECT 526.950 679.950 529.050 682.050 ;
        RECT 529.950 679.950 532.050 682.050 ;
        RECT 532.950 679.950 535.050 682.050 ;
        RECT 535.950 679.950 538.050 682.050 ;
        RECT 550.950 679.950 553.050 682.050 ;
        RECT 553.950 679.950 556.050 682.050 ;
        RECT 556.950 679.950 559.050 682.050 ;
        RECT 571.950 679.950 574.050 682.050 ;
        RECT 574.950 679.950 577.050 682.050 ;
        RECT 577.950 679.950 580.050 682.050 ;
        RECT 580.950 679.950 583.050 682.050 ;
        RECT 515.100 678.150 516.900 679.950 ;
        RECT 530.100 678.150 531.900 679.950 ;
        RECT 533.850 675.750 535.050 679.950 ;
        RECT 536.100 678.150 537.900 679.950 ;
        RECT 551.100 678.150 552.900 679.950 ;
        RECT 509.100 674.400 516.600 675.300 ;
        RECT 533.850 674.700 537.600 675.750 ;
        RECT 509.100 673.500 510.900 674.400 ;
        RECT 488.400 666.600 490.200 672.600 ;
        RECT 506.400 670.800 509.100 672.600 ;
        RECT 507.300 666.600 509.100 670.800 ;
        RECT 514.800 666.600 516.600 674.400 ;
        RECT 527.400 671.700 535.200 673.050 ;
        RECT 527.400 666.600 529.200 671.700 ;
        RECT 533.400 666.600 535.200 671.700 ;
        RECT 536.400 672.600 537.600 674.700 ;
        RECT 554.400 674.700 555.600 679.950 ;
        RECT 557.100 678.150 558.900 679.950 ;
        RECT 575.100 678.150 576.900 679.950 ;
        RECT 578.850 675.750 580.050 679.950 ;
        RECT 581.100 678.150 582.900 679.950 ;
        RECT 587.550 679.050 588.450 682.950 ;
        RECT 596.100 682.050 597.900 683.850 ;
        RECT 601.950 682.050 603.150 695.400 ;
        RECT 622.800 689.400 624.600 701.400 ;
        RECT 628.800 695.400 630.600 701.400 ;
        RECT 623.400 682.050 624.300 689.400 ;
        RECT 626.100 682.050 627.900 683.850 ;
        RECT 595.950 679.950 598.050 682.050 ;
        RECT 598.950 679.950 601.050 682.050 ;
        RECT 601.950 679.950 604.050 682.050 ;
        RECT 604.950 679.950 607.050 682.050 ;
        RECT 622.950 679.950 625.050 682.050 ;
        RECT 625.950 679.950 628.050 682.050 ;
        RECT 583.950 677.550 588.450 679.050 ;
        RECT 599.100 678.150 600.900 679.950 ;
        RECT 583.950 676.950 588.000 677.550 ;
        RECT 602.850 675.750 604.050 679.950 ;
        RECT 605.100 678.150 606.900 679.950 ;
        RECT 578.850 674.700 582.600 675.750 ;
        RECT 602.850 674.700 606.600 675.750 ;
        RECT 554.400 673.800 558.600 674.700 ;
        RECT 536.400 666.600 538.200 672.600 ;
        RECT 556.800 666.600 558.600 673.800 ;
        RECT 572.400 671.700 580.200 673.050 ;
        RECT 572.400 666.600 574.200 671.700 ;
        RECT 578.400 666.600 580.200 671.700 ;
        RECT 581.400 672.600 582.600 674.700 ;
        RECT 581.400 666.600 583.200 672.600 ;
        RECT 596.400 671.700 604.200 673.050 ;
        RECT 596.400 666.600 598.200 671.700 ;
        RECT 602.400 666.600 604.200 671.700 ;
        RECT 605.400 672.600 606.600 674.700 ;
        RECT 623.400 672.600 624.300 679.950 ;
        RECT 629.700 675.300 630.600 695.400 ;
        RECT 649.500 690.600 651.300 701.400 ;
        RECT 647.700 689.400 651.300 690.600 ;
        RECT 670.800 689.400 672.600 701.400 ;
        RECT 673.800 690.300 675.600 701.400 ;
        RECT 679.800 690.300 681.600 701.400 ;
        RECT 694.800 695.400 696.600 701.400 ;
        RECT 673.800 689.400 681.600 690.300 ;
        RECT 695.700 695.100 696.600 695.400 ;
        RECT 700.800 695.400 702.600 701.400 ;
        RECT 722.400 695.400 724.200 701.400 ;
        RECT 745.800 695.400 747.600 701.400 ;
        RECT 766.800 695.400 768.600 701.400 ;
        RECT 700.800 695.100 702.300 695.400 ;
        RECT 695.700 694.200 702.300 695.100 ;
        RECT 644.100 682.050 645.900 683.850 ;
        RECT 647.700 682.050 648.600 689.400 ;
        RECT 649.950 687.450 652.050 688.050 ;
        RECT 667.950 687.450 670.050 688.050 ;
        RECT 649.950 686.550 670.050 687.450 ;
        RECT 649.950 685.950 652.050 686.550 ;
        RECT 667.950 685.950 670.050 686.550 ;
        RECT 650.100 682.050 651.900 683.850 ;
        RECT 671.400 682.050 672.300 689.400 ;
        RECT 690.000 684.450 694.050 685.050 ;
        RECT 677.100 682.050 678.900 683.850 ;
        RECT 689.550 682.950 694.050 684.450 ;
        RECT 631.950 679.950 634.050 682.050 ;
        RECT 643.950 679.950 646.050 682.050 ;
        RECT 646.950 679.950 649.050 682.050 ;
        RECT 649.950 679.950 652.050 682.050 ;
        RECT 670.950 679.950 673.050 682.050 ;
        RECT 673.950 679.950 676.050 682.050 ;
        RECT 676.950 679.950 679.050 682.050 ;
        RECT 679.950 679.950 682.050 682.050 ;
        RECT 632.100 678.150 633.900 679.950 ;
        RECT 626.100 674.400 633.600 675.300 ;
        RECT 626.100 673.500 627.900 674.400 ;
        RECT 605.400 666.600 607.200 672.600 ;
        RECT 623.400 670.800 626.100 672.600 ;
        RECT 624.300 666.600 626.100 670.800 ;
        RECT 631.800 666.600 633.600 674.400 ;
        RECT 647.700 669.600 648.600 679.950 ;
        RECT 671.400 672.600 672.300 679.950 ;
        RECT 674.100 678.150 675.900 679.950 ;
        RECT 680.100 678.150 681.900 679.950 ;
        RECT 682.950 678.450 685.050 679.050 ;
        RECT 689.550 678.450 690.450 682.950 ;
        RECT 695.700 682.050 696.600 694.200 ;
        RECT 701.100 682.050 702.900 683.850 ;
        RECT 722.850 682.050 724.050 695.400 ;
        RECT 728.100 682.050 729.900 683.850 ;
        RECT 740.100 682.050 741.900 683.850 ;
        RECT 745.950 682.050 747.150 695.400 ;
        RECT 767.700 695.100 768.600 695.400 ;
        RECT 772.800 695.400 774.600 701.400 ;
        RECT 772.800 695.100 774.300 695.400 ;
        RECT 767.700 694.200 774.300 695.100 ;
        RECT 767.700 682.050 768.600 694.200 ;
        RECT 788.400 690.300 790.200 701.400 ;
        RECT 794.400 690.300 796.200 701.400 ;
        RECT 788.400 689.400 796.200 690.300 ;
        RECT 797.400 689.400 799.200 701.400 ;
        RECT 817.800 695.400 819.600 701.400 ;
        RECT 773.100 682.050 774.900 683.850 ;
        RECT 791.100 682.050 792.900 683.850 ;
        RECT 797.700 682.050 798.600 689.400 ;
        RECT 812.100 682.050 813.900 683.850 ;
        RECT 817.950 682.050 819.150 695.400 ;
        RECT 838.800 689.400 840.600 701.400 ;
        RECT 841.800 690.300 843.600 701.400 ;
        RECT 847.800 690.300 849.600 701.400 ;
        RECT 863.400 695.400 865.200 701.400 ;
        RECT 863.700 695.100 865.200 695.400 ;
        RECT 869.400 695.400 871.200 701.400 ;
        RECT 884.400 695.400 886.200 701.400 ;
        RECT 869.400 695.100 870.300 695.400 ;
        RECT 863.700 694.200 870.300 695.100 ;
        RECT 841.800 689.400 849.600 690.300 ;
        RECT 839.400 682.050 840.300 689.400 ;
        RECT 847.950 687.450 850.050 688.050 ;
        RECT 856.950 687.450 859.050 688.050 ;
        RECT 865.950 687.450 868.050 688.050 ;
        RECT 847.950 686.550 868.050 687.450 ;
        RECT 847.950 685.950 850.050 686.550 ;
        RECT 856.950 685.950 859.050 686.550 ;
        RECT 865.950 685.950 868.050 686.550 ;
        RECT 845.100 682.050 846.900 683.850 ;
        RECT 863.100 682.050 864.900 683.850 ;
        RECT 869.400 682.050 870.300 694.200 ;
        RECT 884.400 688.500 885.600 695.400 ;
        RECT 890.400 689.400 892.200 701.400 ;
        RECT 884.400 687.600 890.100 688.500 ;
        RECT 888.150 686.700 890.100 687.600 ;
        RECT 871.950 684.450 876.000 685.050 ;
        RECT 871.950 682.950 876.450 684.450 ;
        RECT 694.950 679.950 697.050 682.050 ;
        RECT 697.950 679.950 700.050 682.050 ;
        RECT 700.950 679.950 703.050 682.050 ;
        RECT 703.950 679.950 706.050 682.050 ;
        RECT 718.950 679.950 721.050 682.050 ;
        RECT 721.950 679.950 724.050 682.050 ;
        RECT 724.950 679.950 727.050 682.050 ;
        RECT 727.950 679.950 730.050 682.050 ;
        RECT 739.950 679.950 742.050 682.050 ;
        RECT 742.950 679.950 745.050 682.050 ;
        RECT 745.950 679.950 748.050 682.050 ;
        RECT 748.950 679.950 751.050 682.050 ;
        RECT 766.950 679.950 769.050 682.050 ;
        RECT 769.950 679.950 772.050 682.050 ;
        RECT 772.950 679.950 775.050 682.050 ;
        RECT 775.950 679.950 778.050 682.050 ;
        RECT 787.950 679.950 790.050 682.050 ;
        RECT 790.950 679.950 793.050 682.050 ;
        RECT 793.950 679.950 796.050 682.050 ;
        RECT 796.950 679.950 799.050 682.050 ;
        RECT 811.950 679.950 814.050 682.050 ;
        RECT 814.950 679.950 817.050 682.050 ;
        RECT 817.950 679.950 820.050 682.050 ;
        RECT 820.950 679.950 823.050 682.050 ;
        RECT 838.950 679.950 841.050 682.050 ;
        RECT 841.950 679.950 844.050 682.050 ;
        RECT 844.950 679.950 847.050 682.050 ;
        RECT 847.950 679.950 850.050 682.050 ;
        RECT 859.950 679.950 862.050 682.050 ;
        RECT 862.950 679.950 865.050 682.050 ;
        RECT 865.950 679.950 868.050 682.050 ;
        RECT 868.950 679.950 871.050 682.050 ;
        RECT 682.950 677.550 690.450 678.450 ;
        RECT 682.950 676.950 685.050 677.550 ;
        RECT 695.700 676.200 696.600 679.950 ;
        RECT 698.100 678.150 699.900 679.950 ;
        RECT 704.100 678.150 705.900 679.950 ;
        RECT 719.100 678.150 720.900 679.950 ;
        RECT 695.700 675.000 699.000 676.200 ;
        RECT 721.950 675.750 723.150 679.950 ;
        RECT 725.100 678.150 726.900 679.950 ;
        RECT 743.100 678.150 744.900 679.950 ;
        RECT 671.400 671.400 676.500 672.600 ;
        RECT 647.400 666.600 649.200 669.600 ;
        RECT 674.700 666.600 676.500 671.400 ;
        RECT 697.200 666.600 699.000 675.000 ;
        RECT 719.400 674.700 723.150 675.750 ;
        RECT 746.850 675.750 748.050 679.950 ;
        RECT 749.100 678.150 750.900 679.950 ;
        RECT 767.700 676.200 768.600 679.950 ;
        RECT 770.100 678.150 771.900 679.950 ;
        RECT 776.100 678.150 777.900 679.950 ;
        RECT 788.100 678.150 789.900 679.950 ;
        RECT 794.100 678.150 795.900 679.950 ;
        RECT 746.850 674.700 750.600 675.750 ;
        RECT 767.700 675.000 771.000 676.200 ;
        RECT 719.400 672.600 720.600 674.700 ;
        RECT 718.800 666.600 720.600 672.600 ;
        RECT 721.800 671.700 729.600 673.050 ;
        RECT 721.800 666.600 723.600 671.700 ;
        RECT 727.800 666.600 729.600 671.700 ;
        RECT 740.400 671.700 748.200 673.050 ;
        RECT 740.400 666.600 742.200 671.700 ;
        RECT 746.400 666.600 748.200 671.700 ;
        RECT 749.400 672.600 750.600 674.700 ;
        RECT 749.400 666.600 751.200 672.600 ;
        RECT 769.200 666.600 771.000 675.000 ;
        RECT 797.700 672.600 798.600 679.950 ;
        RECT 799.950 678.450 802.050 679.050 ;
        RECT 805.950 678.450 808.050 679.050 ;
        RECT 799.950 677.550 808.050 678.450 ;
        RECT 815.100 678.150 816.900 679.950 ;
        RECT 799.950 676.950 802.050 677.550 ;
        RECT 805.950 676.950 808.050 677.550 ;
        RECT 818.850 675.750 820.050 679.950 ;
        RECT 821.100 678.150 822.900 679.950 ;
        RECT 818.850 674.700 822.600 675.750 ;
        RECT 793.500 671.400 798.600 672.600 ;
        RECT 812.400 671.700 820.200 673.050 ;
        RECT 793.500 666.600 795.300 671.400 ;
        RECT 812.400 666.600 814.200 671.700 ;
        RECT 818.400 666.600 820.200 671.700 ;
        RECT 821.400 672.600 822.600 674.700 ;
        RECT 839.400 672.600 840.300 679.950 ;
        RECT 842.100 678.150 843.900 679.950 ;
        RECT 848.100 678.150 849.900 679.950 ;
        RECT 860.100 678.150 861.900 679.950 ;
        RECT 866.100 678.150 867.900 679.950 ;
        RECT 869.400 676.200 870.300 679.950 ;
        RECT 875.550 679.050 876.450 682.950 ;
        RECT 884.100 682.050 885.900 683.850 ;
        RECT 883.950 679.950 886.050 682.050 ;
        RECT 871.950 678.450 876.450 679.050 ;
        RECT 880.950 678.450 883.050 679.050 ;
        RECT 871.950 677.550 883.050 678.450 ;
        RECT 871.950 676.950 876.000 677.550 ;
        RECT 880.950 676.950 883.050 677.550 ;
        RECT 867.000 675.000 870.300 676.200 ;
        RECT 888.150 675.300 889.050 686.700 ;
        RECT 891.000 682.050 892.200 689.400 ;
        RECT 889.950 679.950 892.200 682.050 ;
        RECT 821.400 666.600 823.200 672.600 ;
        RECT 839.400 671.400 844.500 672.600 ;
        RECT 842.700 666.600 844.500 671.400 ;
        RECT 867.000 666.600 868.800 675.000 ;
        RECT 888.150 674.400 890.100 675.300 ;
        RECT 884.400 673.500 890.100 674.400 ;
        RECT 884.400 669.600 885.600 673.500 ;
        RECT 891.000 672.600 892.200 679.950 ;
        RECT 884.400 666.600 886.200 669.600 ;
        RECT 890.400 666.600 892.200 672.600 ;
        RECT 16.800 659.400 18.600 662.400 ;
        RECT 35.400 659.400 37.200 662.400 ;
        RECT 7.950 657.450 10.050 658.050 ;
        RECT 13.950 657.450 16.050 658.050 ;
        RECT 7.950 656.550 16.050 657.450 ;
        RECT 7.950 655.950 10.050 656.550 ;
        RECT 13.950 655.950 16.050 656.550 ;
        RECT 17.400 649.050 18.300 659.400 ;
        RECT 27.000 651.450 31.050 652.050 ;
        RECT 26.550 649.950 31.050 651.450 ;
        RECT 13.950 646.950 16.050 649.050 ;
        RECT 16.950 646.950 19.050 649.050 ;
        RECT 19.950 646.950 22.050 649.050 ;
        RECT 14.100 645.150 15.900 646.950 ;
        RECT 17.400 639.600 18.300 646.950 ;
        RECT 20.100 645.150 21.900 646.950 ;
        RECT 26.550 646.050 27.450 649.950 ;
        RECT 35.400 649.050 36.600 659.400 ;
        RECT 50.400 657.300 52.200 662.400 ;
        RECT 56.400 657.300 58.200 662.400 ;
        RECT 50.400 655.950 58.200 657.300 ;
        RECT 59.400 656.400 61.200 662.400 ;
        RECT 79.800 659.400 81.600 662.400 ;
        RECT 64.950 657.450 67.050 658.050 ;
        RECT 76.950 657.450 79.050 658.050 ;
        RECT 64.950 656.550 79.050 657.450 ;
        RECT 59.400 654.300 60.600 656.400 ;
        RECT 64.950 655.950 67.050 656.550 ;
        RECT 76.950 655.950 79.050 656.550 ;
        RECT 56.850 653.250 60.600 654.300 ;
        RECT 53.100 649.050 54.900 650.850 ;
        RECT 56.850 649.050 58.050 653.250 ;
        RECT 59.100 649.050 60.900 650.850 ;
        RECT 80.400 649.050 81.300 659.400 ;
        RECT 82.950 654.450 85.050 655.200 ;
        RECT 88.950 654.450 91.050 655.050 ;
        RECT 82.950 653.550 91.050 654.450 ;
        RECT 82.950 653.100 85.050 653.550 ;
        RECT 88.950 652.950 91.050 653.550 ;
        RECT 105.000 654.000 106.800 662.400 ;
        RECT 124.800 659.400 126.600 662.400 ;
        RECT 105.000 652.800 108.300 654.000 ;
        RECT 98.100 649.050 99.900 650.850 ;
        RECT 104.100 649.050 105.900 650.850 ;
        RECT 107.400 649.050 108.300 652.800 ;
        RECT 125.400 649.050 126.600 659.400 ;
        RECT 131.550 656.400 133.350 662.400 ;
        RECT 139.650 659.400 141.450 662.400 ;
        RECT 147.450 659.400 149.250 662.400 ;
        RECT 155.250 660.300 157.050 662.400 ;
        RECT 155.250 659.400 159.000 660.300 ;
        RECT 139.650 658.500 140.700 659.400 ;
        RECT 136.950 657.300 140.700 658.500 ;
        RECT 148.200 658.500 149.250 659.400 ;
        RECT 157.950 658.500 159.000 659.400 ;
        RECT 148.200 657.450 153.150 658.500 ;
        RECT 136.950 656.400 139.050 657.300 ;
        RECT 151.350 656.700 153.150 657.450 ;
        RECT 131.550 649.050 132.750 656.400 ;
        RECT 154.650 655.800 156.450 657.600 ;
        RECT 157.950 656.400 160.050 658.500 ;
        RECT 163.050 656.400 164.850 662.400 ;
        RECT 144.150 654.000 145.950 654.600 ;
        RECT 155.100 654.000 156.150 655.800 ;
        RECT 144.150 652.800 156.150 654.000 ;
        RECT 31.950 646.950 34.050 649.050 ;
        RECT 34.950 646.950 37.050 649.050 ;
        RECT 49.950 646.950 52.050 649.050 ;
        RECT 52.950 646.950 55.050 649.050 ;
        RECT 55.950 646.950 58.050 649.050 ;
        RECT 58.950 646.950 61.050 649.050 ;
        RECT 76.950 646.950 79.050 649.050 ;
        RECT 79.950 646.950 82.050 649.050 ;
        RECT 82.950 646.950 85.050 649.050 ;
        RECT 97.950 646.950 100.050 649.050 ;
        RECT 100.950 646.950 103.050 649.050 ;
        RECT 103.950 646.950 106.050 649.050 ;
        RECT 106.950 646.950 109.050 649.050 ;
        RECT 124.950 646.950 127.050 649.050 ;
        RECT 127.950 646.950 130.050 649.050 ;
        RECT 131.550 647.250 137.850 649.050 ;
        RECT 131.550 646.950 136.050 647.250 ;
        RECT 26.550 644.550 31.050 646.050 ;
        RECT 32.100 645.150 33.900 646.950 ;
        RECT 27.000 643.950 31.050 644.550 ;
        RECT 14.700 638.400 18.300 639.600 ;
        RECT 1.950 630.450 4.050 631.050 ;
        RECT 7.950 630.450 10.050 631.050 ;
        RECT 1.950 629.550 10.050 630.450 ;
        RECT 1.950 628.950 4.050 629.550 ;
        RECT 7.950 628.950 10.050 629.550 ;
        RECT 14.700 627.600 16.500 638.400 ;
        RECT 35.400 633.600 36.600 646.950 ;
        RECT 50.100 645.150 51.900 646.950 ;
        RECT 55.950 633.600 57.150 646.950 ;
        RECT 77.100 645.150 78.900 646.950 ;
        RECT 80.400 639.600 81.300 646.950 ;
        RECT 83.100 645.150 84.900 646.950 ;
        RECT 101.100 645.150 102.900 646.950 ;
        RECT 77.700 638.400 81.300 639.600 ;
        RECT 35.400 627.600 37.200 633.600 ;
        RECT 55.800 627.600 57.600 633.600 ;
        RECT 77.700 627.600 79.500 638.400 ;
        RECT 107.400 634.800 108.300 646.950 ;
        RECT 101.700 633.900 108.300 634.800 ;
        RECT 101.700 633.600 103.200 633.900 ;
        RECT 101.400 627.600 103.200 633.600 ;
        RECT 107.400 633.600 108.300 633.900 ;
        RECT 125.400 633.600 126.600 646.950 ;
        RECT 128.100 645.150 129.900 646.950 ;
        RECT 107.400 627.600 109.200 633.600 ;
        RECT 124.800 627.600 126.600 633.600 ;
        RECT 131.550 639.600 132.750 646.950 ;
        RECT 133.950 641.400 135.750 643.200 ;
        RECT 134.850 640.200 139.050 641.400 ;
        RECT 144.150 640.200 145.050 652.800 ;
        RECT 155.100 651.600 162.000 652.800 ;
        RECT 155.100 651.000 156.900 651.600 ;
        RECT 161.100 650.850 162.000 651.600 ;
        RECT 158.100 649.800 159.900 650.400 ;
        RECT 151.950 648.600 159.900 649.800 ;
        RECT 161.100 649.050 162.900 650.850 ;
        RECT 151.950 646.950 154.050 648.600 ;
        RECT 160.950 646.950 163.050 649.050 ;
        RECT 153.750 641.700 155.550 642.000 ;
        RECT 163.950 641.700 164.850 656.400 ;
        RECT 176.400 657.300 178.200 662.400 ;
        RECT 182.400 657.300 184.200 662.400 ;
        RECT 176.400 655.950 184.200 657.300 ;
        RECT 185.400 656.400 187.200 662.400 ;
        RECT 202.800 659.400 204.600 662.400 ;
        RECT 185.400 654.300 186.600 656.400 ;
        RECT 182.850 653.250 186.600 654.300 ;
        RECT 179.100 649.050 180.900 650.850 ;
        RECT 182.850 649.050 184.050 653.250 ;
        RECT 185.100 649.050 186.900 650.850 ;
        RECT 203.400 649.050 204.600 659.400 ;
        RECT 220.800 656.400 222.600 662.400 ;
        RECT 205.950 654.450 208.050 655.050 ;
        RECT 214.950 654.450 217.050 655.050 ;
        RECT 205.950 653.550 217.050 654.450 ;
        RECT 205.950 652.950 208.050 653.550 ;
        RECT 214.950 652.950 217.050 653.550 ;
        RECT 221.400 654.300 222.600 656.400 ;
        RECT 223.800 657.300 225.600 662.400 ;
        RECT 229.800 657.300 231.600 662.400 ;
        RECT 248.700 657.600 250.500 662.400 ;
        RECT 223.800 655.950 231.600 657.300 ;
        RECT 245.400 656.400 250.500 657.600 ;
        RECT 221.400 653.250 225.150 654.300 ;
        RECT 221.100 649.050 222.900 650.850 ;
        RECT 223.950 649.050 225.150 653.250 ;
        RECT 227.100 649.050 228.900 650.850 ;
        RECT 245.400 649.050 246.300 656.400 ;
        RECT 273.000 654.000 274.800 662.400 ;
        RECT 295.800 656.400 297.600 662.400 ;
        RECT 296.400 654.300 297.600 656.400 ;
        RECT 298.800 657.300 300.600 662.400 ;
        RECT 304.800 657.300 306.600 662.400 ;
        RECT 320.400 659.400 322.200 662.400 ;
        RECT 298.800 655.950 306.600 657.300 ;
        RECT 307.950 657.450 310.050 658.050 ;
        RECT 316.950 657.450 319.050 658.050 ;
        RECT 307.950 656.550 319.050 657.450 ;
        RECT 307.950 655.950 310.050 656.550 ;
        RECT 316.950 655.950 319.050 656.550 ;
        RECT 273.000 652.800 276.300 654.000 ;
        RECT 296.400 653.250 300.150 654.300 ;
        RECT 248.100 649.050 249.900 650.850 ;
        RECT 254.100 649.050 255.900 650.850 ;
        RECT 266.100 649.050 267.900 650.850 ;
        RECT 272.100 649.050 273.900 650.850 ;
        RECT 275.400 649.050 276.300 652.800 ;
        RECT 296.100 649.050 297.900 650.850 ;
        RECT 298.950 649.050 300.150 653.250 ;
        RECT 302.100 649.050 303.900 650.850 ;
        RECT 320.700 649.050 321.600 659.400 ;
        RECT 343.800 655.200 345.600 662.400 ;
        RECT 363.300 658.200 365.100 662.400 ;
        RECT 341.400 654.300 345.600 655.200 ;
        RECT 362.400 656.400 365.100 658.200 ;
        RECT 338.100 649.050 339.900 650.850 ;
        RECT 341.400 649.050 342.600 654.300 ;
        RECT 344.100 649.050 345.900 650.850 ;
        RECT 362.400 649.050 363.300 656.400 ;
        RECT 365.100 654.600 366.900 655.500 ;
        RECT 370.800 654.600 372.600 662.400 ;
        RECT 385.800 656.400 387.600 662.400 ;
        RECT 365.100 653.700 372.600 654.600 ;
        RECT 386.400 654.300 387.600 656.400 ;
        RECT 388.800 657.300 390.600 662.400 ;
        RECT 394.800 657.300 396.600 662.400 ;
        RECT 388.800 655.950 396.600 657.300 ;
        RECT 412.800 655.200 414.600 662.400 ;
        RECT 433.800 655.200 435.600 662.400 ;
        RECT 451.800 656.400 453.600 662.400 ;
        RECT 410.400 654.300 414.600 655.200 ;
        RECT 431.400 654.300 435.600 655.200 ;
        RECT 452.400 654.300 453.600 656.400 ;
        RECT 454.800 657.300 456.600 662.400 ;
        RECT 460.800 657.300 462.600 662.400 ;
        RECT 454.800 655.950 462.600 657.300 ;
        RECT 476.400 655.200 478.200 662.400 ;
        RECT 476.400 654.300 480.600 655.200 ;
        RECT 175.950 646.950 178.050 649.050 ;
        RECT 178.950 646.950 181.050 649.050 ;
        RECT 181.950 646.950 184.050 649.050 ;
        RECT 184.950 646.950 187.050 649.050 ;
        RECT 202.950 646.950 205.050 649.050 ;
        RECT 205.950 646.950 208.050 649.050 ;
        RECT 220.950 646.950 223.050 649.050 ;
        RECT 223.950 646.950 226.050 649.050 ;
        RECT 226.950 646.950 229.050 649.050 ;
        RECT 229.950 646.950 232.050 649.050 ;
        RECT 244.950 646.950 247.050 649.050 ;
        RECT 247.950 646.950 250.050 649.050 ;
        RECT 250.950 646.950 253.050 649.050 ;
        RECT 253.950 646.950 256.050 649.050 ;
        RECT 265.950 646.950 268.050 649.050 ;
        RECT 268.950 646.950 271.050 649.050 ;
        RECT 271.950 646.950 274.050 649.050 ;
        RECT 274.950 646.950 277.050 649.050 ;
        RECT 295.950 646.950 298.050 649.050 ;
        RECT 298.950 646.950 301.050 649.050 ;
        RECT 301.950 646.950 304.050 649.050 ;
        RECT 304.950 646.950 307.050 649.050 ;
        RECT 316.950 646.950 319.050 649.050 ;
        RECT 319.950 646.950 322.050 649.050 ;
        RECT 322.950 646.950 325.050 649.050 ;
        RECT 337.950 646.950 340.050 649.050 ;
        RECT 340.950 646.950 343.050 649.050 ;
        RECT 343.950 646.950 346.050 649.050 ;
        RECT 361.950 646.950 364.050 649.050 ;
        RECT 364.950 646.950 367.050 649.050 ;
        RECT 176.100 645.150 177.900 646.950 ;
        RECT 153.750 641.100 164.850 641.700 ;
        RECT 131.550 627.600 133.350 639.600 ;
        RECT 136.950 639.300 139.050 640.200 ;
        RECT 139.950 639.300 145.050 640.200 ;
        RECT 147.150 640.500 164.850 641.100 ;
        RECT 147.150 640.200 155.550 640.500 ;
        RECT 139.950 638.400 140.850 639.300 ;
        RECT 138.150 636.600 140.850 638.400 ;
        RECT 141.750 638.100 143.550 638.400 ;
        RECT 147.150 638.100 148.050 640.200 ;
        RECT 163.950 639.600 164.850 640.500 ;
        RECT 141.750 637.200 148.050 638.100 ;
        RECT 148.950 638.700 150.750 639.300 ;
        RECT 148.950 637.500 156.450 638.700 ;
        RECT 141.750 636.600 143.550 637.200 ;
        RECT 155.250 636.600 156.450 637.500 ;
        RECT 136.950 633.600 140.850 635.700 ;
        RECT 145.950 635.550 147.750 636.300 ;
        RECT 150.750 635.550 152.550 636.300 ;
        RECT 145.950 634.500 152.550 635.550 ;
        RECT 155.250 634.500 160.050 636.600 ;
        RECT 139.050 627.600 140.850 633.600 ;
        RECT 146.850 627.600 148.650 634.500 ;
        RECT 155.250 633.600 156.450 634.500 ;
        RECT 154.650 627.600 156.450 633.600 ;
        RECT 163.050 627.600 164.850 639.600 ;
        RECT 181.950 633.600 183.150 646.950 ;
        RECT 203.400 633.600 204.600 646.950 ;
        RECT 206.100 645.150 207.900 646.950 ;
        RECT 224.850 633.600 226.050 646.950 ;
        RECT 230.100 645.150 231.900 646.950 ;
        RECT 245.400 639.600 246.300 646.950 ;
        RECT 251.100 645.150 252.900 646.950 ;
        RECT 269.100 645.150 270.900 646.950 ;
        RECT 181.800 627.600 183.600 633.600 ;
        RECT 202.800 627.600 204.600 633.600 ;
        RECT 224.400 627.600 226.200 633.600 ;
        RECT 244.800 627.600 246.600 639.600 ;
        RECT 247.800 638.700 255.600 639.600 ;
        RECT 247.800 627.600 249.600 638.700 ;
        RECT 253.800 627.600 255.600 638.700 ;
        RECT 275.400 634.800 276.300 646.950 ;
        RECT 269.700 633.900 276.300 634.800 ;
        RECT 269.700 633.600 271.200 633.900 ;
        RECT 269.400 627.600 271.200 633.600 ;
        RECT 275.400 633.600 276.300 633.900 ;
        RECT 299.850 633.600 301.050 646.950 ;
        RECT 305.100 645.150 306.900 646.950 ;
        RECT 317.100 645.150 318.900 646.950 ;
        RECT 320.700 639.600 321.600 646.950 ;
        RECT 323.100 645.150 324.900 646.950 ;
        RECT 320.700 638.400 324.300 639.600 ;
        RECT 275.400 627.600 277.200 633.600 ;
        RECT 299.400 627.600 301.200 633.600 ;
        RECT 322.500 627.600 324.300 638.400 ;
        RECT 341.400 633.600 342.600 646.950 ;
        RECT 362.400 639.600 363.300 646.950 ;
        RECT 365.100 645.150 366.900 646.950 ;
        RECT 341.400 627.600 343.200 633.600 ;
        RECT 361.800 627.600 363.600 639.600 ;
        RECT 368.700 633.600 369.600 653.700 ;
        RECT 386.400 653.250 390.150 654.300 ;
        RECT 371.100 649.050 372.900 650.850 ;
        RECT 386.100 649.050 387.900 650.850 ;
        RECT 388.950 649.050 390.150 653.250 ;
        RECT 392.100 649.050 393.900 650.850 ;
        RECT 407.100 649.050 408.900 650.850 ;
        RECT 410.400 649.050 411.600 654.300 ;
        RECT 415.950 651.450 420.000 652.050 ;
        RECT 413.100 649.050 414.900 650.850 ;
        RECT 415.950 649.950 420.450 651.450 ;
        RECT 370.950 646.950 373.050 649.050 ;
        RECT 385.950 646.950 388.050 649.050 ;
        RECT 388.950 646.950 391.050 649.050 ;
        RECT 391.950 646.950 394.050 649.050 ;
        RECT 394.950 646.950 397.050 649.050 ;
        RECT 406.950 646.950 409.050 649.050 ;
        RECT 409.950 646.950 412.050 649.050 ;
        RECT 412.950 646.950 415.050 649.050 ;
        RECT 389.850 633.600 391.050 646.950 ;
        RECT 395.100 645.150 396.900 646.950 ;
        RECT 410.400 633.600 411.600 646.950 ;
        RECT 419.550 646.050 420.450 649.950 ;
        RECT 428.100 649.050 429.900 650.850 ;
        RECT 431.400 649.050 432.600 654.300 ;
        RECT 452.400 653.250 456.150 654.300 ;
        RECT 434.100 649.050 435.900 650.850 ;
        RECT 452.100 649.050 453.900 650.850 ;
        RECT 454.950 649.050 456.150 653.250 ;
        RECT 458.100 649.050 459.900 650.850 ;
        RECT 476.100 649.050 477.900 650.850 ;
        RECT 479.400 649.050 480.600 654.300 ;
        RECT 494.400 654.600 496.200 662.400 ;
        RECT 501.900 658.200 503.700 662.400 ;
        RECT 501.900 656.400 504.600 658.200 ;
        RECT 500.100 654.600 501.900 655.500 ;
        RECT 494.400 653.700 501.900 654.600 ;
        RECT 482.100 649.050 483.900 650.850 ;
        RECT 494.100 649.050 495.900 650.850 ;
        RECT 427.950 646.950 430.050 649.050 ;
        RECT 430.950 646.950 433.050 649.050 ;
        RECT 433.950 646.950 436.050 649.050 ;
        RECT 451.950 646.950 454.050 649.050 ;
        RECT 454.950 646.950 457.050 649.050 ;
        RECT 457.950 646.950 460.050 649.050 ;
        RECT 460.950 646.950 463.050 649.050 ;
        RECT 475.950 646.950 478.050 649.050 ;
        RECT 478.950 646.950 481.050 649.050 ;
        RECT 481.950 646.950 484.050 649.050 ;
        RECT 493.950 646.950 496.050 649.050 ;
        RECT 415.950 644.550 420.450 646.050 ;
        RECT 415.950 643.950 420.000 644.550 ;
        RECT 412.950 636.450 415.050 637.050 ;
        RECT 427.950 636.450 430.050 637.050 ;
        RECT 412.950 635.550 430.050 636.450 ;
        RECT 412.950 634.950 415.050 635.550 ;
        RECT 427.950 634.950 430.050 635.550 ;
        RECT 431.400 633.600 432.600 646.950 ;
        RECT 433.950 642.450 436.050 643.050 ;
        RECT 445.950 642.450 448.050 643.050 ;
        RECT 433.950 641.550 448.050 642.450 ;
        RECT 433.950 640.950 436.050 641.550 ;
        RECT 445.950 640.950 448.050 641.550 ;
        RECT 455.850 633.600 457.050 646.950 ;
        RECT 461.100 645.150 462.900 646.950 ;
        RECT 479.400 633.600 480.600 646.950 ;
        RECT 367.800 627.600 369.600 633.600 ;
        RECT 389.400 627.600 391.200 633.600 ;
        RECT 410.400 627.600 412.200 633.600 ;
        RECT 431.400 627.600 433.200 633.600 ;
        RECT 455.400 627.600 457.200 633.600 ;
        RECT 478.800 627.600 480.600 633.600 ;
        RECT 497.400 633.600 498.300 653.700 ;
        RECT 503.700 649.050 504.600 656.400 ;
        RECT 523.800 655.200 525.600 662.400 ;
        RECT 521.400 654.300 525.600 655.200 ;
        RECT 542.400 656.400 544.200 662.400 ;
        RECT 559.800 656.400 561.600 662.400 ;
        RECT 577.800 656.400 579.600 662.400 ;
        RECT 518.100 649.050 519.900 650.850 ;
        RECT 521.400 649.050 522.600 654.300 ;
        RECT 524.100 649.050 525.900 650.850 ;
        RECT 539.100 649.050 540.900 650.850 ;
        RECT 542.400 649.050 543.600 656.400 ;
        RECT 544.950 654.450 547.050 655.050 ;
        RECT 556.950 654.450 559.050 655.050 ;
        RECT 544.950 653.550 559.050 654.450 ;
        RECT 544.950 652.950 547.050 653.550 ;
        RECT 556.950 652.950 559.050 653.550 ;
        RECT 560.400 649.050 561.600 656.400 ;
        RECT 578.400 654.300 579.600 656.400 ;
        RECT 580.800 657.300 582.600 662.400 ;
        RECT 586.800 657.300 588.600 662.400 ;
        RECT 580.800 655.950 588.600 657.300 ;
        RECT 601.800 656.400 603.600 662.400 ;
        RECT 607.800 659.400 609.600 662.400 ;
        RECT 578.400 653.250 582.150 654.300 ;
        RECT 563.100 649.050 564.900 650.850 ;
        RECT 578.100 649.050 579.900 650.850 ;
        RECT 580.950 649.050 582.150 653.250 ;
        RECT 584.100 649.050 585.900 650.850 ;
        RECT 601.800 649.050 603.000 656.400 ;
        RECT 608.400 655.500 609.600 659.400 ;
        RECT 603.900 654.600 609.600 655.500 ;
        RECT 603.900 653.700 605.850 654.600 ;
        RECT 625.200 654.000 627.000 662.400 ;
        RECT 647.400 655.200 649.200 662.400 ;
        RECT 670.800 655.200 672.600 662.400 ;
        RECT 696.000 656.400 697.800 662.400 ;
        RECT 718.200 656.400 720.000 662.400 ;
        RECT 746.700 657.600 748.500 662.400 ;
        RECT 647.400 654.300 651.600 655.200 ;
        RECT 499.950 646.950 502.050 649.050 ;
        RECT 502.950 646.950 505.050 649.050 ;
        RECT 517.950 646.950 520.050 649.050 ;
        RECT 520.950 646.950 523.050 649.050 ;
        RECT 523.950 646.950 526.050 649.050 ;
        RECT 538.950 646.950 541.050 649.050 ;
        RECT 541.950 646.950 544.050 649.050 ;
        RECT 559.950 646.950 562.050 649.050 ;
        RECT 562.950 646.950 565.050 649.050 ;
        RECT 577.950 646.950 580.050 649.050 ;
        RECT 580.950 646.950 583.050 649.050 ;
        RECT 583.950 646.950 586.050 649.050 ;
        RECT 586.950 646.950 589.050 649.050 ;
        RECT 601.800 646.950 604.050 649.050 ;
        RECT 500.100 645.150 501.900 646.950 ;
        RECT 503.700 639.600 504.600 646.950 ;
        RECT 497.400 627.600 499.200 633.600 ;
        RECT 503.400 627.600 505.200 639.600 ;
        RECT 521.400 633.600 522.600 646.950 ;
        RECT 542.400 639.600 543.600 646.950 ;
        RECT 560.400 639.600 561.600 646.950 ;
        RECT 521.400 627.600 523.200 633.600 ;
        RECT 542.400 627.600 544.200 639.600 ;
        RECT 559.800 627.600 561.600 639.600 ;
        RECT 581.850 633.600 583.050 646.950 ;
        RECT 587.100 645.150 588.900 646.950 ;
        RECT 601.800 639.600 603.000 646.950 ;
        RECT 604.950 642.300 605.850 653.700 ;
        RECT 623.700 652.800 627.000 654.000 ;
        RECT 623.700 649.050 624.600 652.800 ;
        RECT 626.100 649.050 627.900 650.850 ;
        RECT 632.100 649.050 633.900 650.850 ;
        RECT 647.100 649.050 648.900 650.850 ;
        RECT 650.400 649.050 651.600 654.300 ;
        RECT 668.400 654.300 672.600 655.200 ;
        RECT 679.950 654.450 682.050 655.050 ;
        RECT 691.950 654.450 694.050 655.200 ;
        RECT 655.950 651.450 660.000 652.050 ;
        RECT 653.100 649.050 654.900 650.850 ;
        RECT 655.950 649.950 660.450 651.450 ;
        RECT 607.950 646.950 610.050 649.050 ;
        RECT 622.950 646.950 625.050 649.050 ;
        RECT 625.950 646.950 628.050 649.050 ;
        RECT 628.950 646.950 631.050 649.050 ;
        RECT 631.950 646.950 634.050 649.050 ;
        RECT 646.950 646.950 649.050 649.050 ;
        RECT 649.950 646.950 652.050 649.050 ;
        RECT 652.950 646.950 655.050 649.050 ;
        RECT 608.100 645.150 609.900 646.950 ;
        RECT 603.900 641.400 605.850 642.300 ;
        RECT 603.900 640.500 609.600 641.400 ;
        RECT 581.400 627.600 583.200 633.600 ;
        RECT 601.800 627.600 603.600 639.600 ;
        RECT 608.400 633.600 609.600 640.500 ;
        RECT 623.700 634.800 624.600 646.950 ;
        RECT 629.100 645.150 630.900 646.950 ;
        RECT 631.950 642.450 634.050 643.050 ;
        RECT 643.950 642.450 646.050 643.050 ;
        RECT 631.950 641.550 646.050 642.450 ;
        RECT 631.950 640.950 634.050 641.550 ;
        RECT 643.950 640.950 646.050 641.550 ;
        RECT 623.700 633.900 630.300 634.800 ;
        RECT 623.700 633.600 624.600 633.900 ;
        RECT 607.800 627.600 609.600 633.600 ;
        RECT 622.800 627.600 624.600 633.600 ;
        RECT 628.800 633.600 630.300 633.900 ;
        RECT 650.400 633.600 651.600 646.950 ;
        RECT 659.550 646.050 660.450 649.950 ;
        RECT 665.100 649.050 666.900 650.850 ;
        RECT 668.400 649.050 669.600 654.300 ;
        RECT 679.950 653.550 694.050 654.450 ;
        RECT 679.950 652.950 682.050 653.550 ;
        RECT 691.950 653.100 694.050 653.550 ;
        RECT 671.100 649.050 672.900 650.850 ;
        RECT 689.100 649.050 690.900 650.850 ;
        RECT 696.000 649.050 697.050 656.400 ;
        RECT 703.950 651.450 706.050 655.050 ;
        RECT 703.950 651.000 708.450 651.450 ;
        RECT 701.100 649.050 702.900 650.850 ;
        RECT 704.550 650.550 708.450 651.000 ;
        RECT 664.950 646.950 667.050 649.050 ;
        RECT 667.950 646.950 670.050 649.050 ;
        RECT 670.950 646.950 673.050 649.050 ;
        RECT 655.950 644.550 660.450 646.050 ;
        RECT 655.950 643.950 660.000 644.550 ;
        RECT 628.800 627.600 630.600 633.600 ;
        RECT 649.800 627.600 651.600 633.600 ;
        RECT 668.400 633.600 669.600 646.950 ;
        RECT 676.950 646.050 679.050 649.050 ;
        RECT 688.950 646.950 691.050 649.050 ;
        RECT 691.950 646.950 694.050 649.050 ;
        RECT 694.950 646.950 697.050 649.050 ;
        RECT 697.950 646.950 700.050 649.050 ;
        RECT 700.950 646.950 703.050 649.050 ;
        RECT 673.950 645.000 679.050 646.050 ;
        RECT 692.100 645.150 693.900 646.950 ;
        RECT 673.950 644.550 678.450 645.000 ;
        RECT 673.950 643.950 678.000 644.550 ;
        RECT 670.950 642.450 673.050 643.050 ;
        RECT 676.950 642.450 679.050 643.050 ;
        RECT 670.950 641.550 679.050 642.450 ;
        RECT 670.950 640.950 673.050 641.550 ;
        RECT 676.950 640.950 679.050 641.550 ;
        RECT 696.000 641.400 696.900 646.950 ;
        RECT 698.100 645.150 699.900 646.950 ;
        RECT 707.550 646.050 708.450 650.550 ;
        RECT 713.100 649.050 714.900 650.850 ;
        RECT 718.950 649.050 720.000 656.400 ;
        RECT 743.400 656.400 748.500 657.600 ;
        RECT 727.950 651.450 732.000 652.050 ;
        RECT 725.100 649.050 726.900 650.850 ;
        RECT 727.950 649.950 732.450 651.450 ;
        RECT 712.950 646.950 715.050 649.050 ;
        RECT 715.950 646.950 718.050 649.050 ;
        RECT 718.950 646.950 721.050 649.050 ;
        RECT 721.950 646.950 724.050 649.050 ;
        RECT 724.950 646.950 727.050 649.050 ;
        RECT 707.550 644.550 712.050 646.050 ;
        RECT 716.100 645.150 717.900 646.950 ;
        RECT 708.000 643.950 712.050 644.550 ;
        RECT 691.800 640.500 696.900 641.400 ;
        RECT 719.100 641.400 720.000 646.950 ;
        RECT 722.100 645.150 723.900 646.950 ;
        RECT 731.550 646.050 732.450 649.950 ;
        RECT 743.400 649.050 744.300 656.400 ;
        RECT 748.950 654.450 751.050 655.200 ;
        RECT 760.950 654.450 763.050 655.050 ;
        RECT 748.950 653.550 763.050 654.450 ;
        RECT 748.950 653.100 751.050 653.550 ;
        RECT 760.950 652.950 763.050 653.550 ;
        RECT 771.000 654.000 772.800 662.400 ;
        RECT 795.000 654.000 796.800 662.400 ;
        RECT 812.400 659.400 814.200 662.400 ;
        RECT 812.400 655.500 813.600 659.400 ;
        RECT 818.400 656.400 820.200 662.400 ;
        RECT 838.500 657.600 840.300 662.400 ;
        RECT 844.950 660.450 847.050 661.050 ;
        RECT 850.950 660.450 853.050 661.050 ;
        RECT 844.950 659.550 853.050 660.450 ;
        RECT 844.950 658.950 847.050 659.550 ;
        RECT 850.950 658.950 853.050 659.550 ;
        RECT 838.500 656.400 843.600 657.600 ;
        RECT 812.400 654.600 818.100 655.500 ;
        RECT 771.000 652.800 774.300 654.000 ;
        RECT 795.000 652.800 798.300 654.000 ;
        RECT 746.100 649.050 747.900 650.850 ;
        RECT 752.100 649.050 753.900 650.850 ;
        RECT 764.100 649.050 765.900 650.850 ;
        RECT 770.100 649.050 771.900 650.850 ;
        RECT 773.400 649.050 774.300 652.800 ;
        RECT 788.100 649.050 789.900 650.850 ;
        RECT 794.100 649.050 795.900 650.850 ;
        RECT 797.400 649.050 798.300 652.800 ;
        RECT 816.150 653.700 818.100 654.600 ;
        RECT 742.950 646.950 745.050 649.050 ;
        RECT 745.950 646.950 748.050 649.050 ;
        RECT 748.950 646.950 751.050 649.050 ;
        RECT 751.950 646.950 754.050 649.050 ;
        RECT 763.950 646.950 766.050 649.050 ;
        RECT 766.950 646.950 769.050 649.050 ;
        RECT 769.950 646.950 772.050 649.050 ;
        RECT 772.950 646.950 775.050 649.050 ;
        RECT 787.950 646.950 790.050 649.050 ;
        RECT 790.950 646.950 793.050 649.050 ;
        RECT 793.950 646.950 796.050 649.050 ;
        RECT 796.950 646.950 799.050 649.050 ;
        RECT 811.950 646.950 814.050 649.050 ;
        RECT 727.950 644.550 732.450 646.050 ;
        RECT 727.950 643.950 732.000 644.550 ;
        RECT 719.100 640.500 724.200 641.400 ;
        RECT 668.400 627.600 670.200 633.600 ;
        RECT 688.800 628.500 690.600 639.600 ;
        RECT 691.800 629.400 693.600 640.500 ;
        RECT 694.800 638.400 702.600 639.300 ;
        RECT 694.800 628.500 696.600 638.400 ;
        RECT 688.800 627.600 696.600 628.500 ;
        RECT 700.800 627.600 702.600 638.400 ;
        RECT 713.400 638.400 721.200 639.300 ;
        RECT 713.400 627.600 715.200 638.400 ;
        RECT 719.400 628.500 721.200 638.400 ;
        RECT 722.400 629.400 724.200 640.500 ;
        RECT 743.400 639.600 744.300 646.950 ;
        RECT 749.100 645.150 750.900 646.950 ;
        RECT 767.100 645.150 768.900 646.950 ;
        RECT 745.950 642.450 748.050 643.050 ;
        RECT 763.950 642.450 766.050 643.050 ;
        RECT 745.950 641.550 766.050 642.450 ;
        RECT 745.950 640.950 748.050 641.550 ;
        RECT 763.950 640.950 766.050 641.550 ;
        RECT 725.400 628.500 727.200 639.600 ;
        RECT 719.400 627.600 727.200 628.500 ;
        RECT 742.800 627.600 744.600 639.600 ;
        RECT 745.800 638.700 753.600 639.600 ;
        RECT 745.800 627.600 747.600 638.700 ;
        RECT 751.800 627.600 753.600 638.700 ;
        RECT 754.950 639.450 757.050 640.050 ;
        RECT 766.950 639.450 769.050 640.050 ;
        RECT 754.950 638.550 769.050 639.450 ;
        RECT 754.950 637.950 757.050 638.550 ;
        RECT 766.950 637.950 769.050 638.550 ;
        RECT 773.400 634.800 774.300 646.950 ;
        RECT 791.100 645.150 792.900 646.950 ;
        RECT 797.400 634.800 798.300 646.950 ;
        RECT 812.100 645.150 813.900 646.950 ;
        RECT 816.150 642.300 817.050 653.700 ;
        RECT 819.000 649.050 820.200 656.400 ;
        RECT 828.000 651.450 832.050 652.050 ;
        RECT 817.950 646.950 820.200 649.050 ;
        RECT 816.150 641.400 818.100 642.300 ;
        RECT 767.700 633.900 774.300 634.800 ;
        RECT 767.700 633.600 769.200 633.900 ;
        RECT 767.400 627.600 769.200 633.600 ;
        RECT 773.400 633.600 774.300 633.900 ;
        RECT 791.700 633.900 798.300 634.800 ;
        RECT 791.700 633.600 793.200 633.900 ;
        RECT 773.400 627.600 775.200 633.600 ;
        RECT 791.400 627.600 793.200 633.600 ;
        RECT 797.400 633.600 798.300 633.900 ;
        RECT 812.400 640.500 818.100 641.400 ;
        RECT 812.400 633.600 813.600 640.500 ;
        RECT 819.000 639.600 820.200 646.950 ;
        RECT 827.550 649.950 832.050 651.450 ;
        RECT 827.550 646.050 828.450 649.950 ;
        RECT 833.100 649.050 834.900 650.850 ;
        RECT 839.100 649.050 840.900 650.850 ;
        RECT 842.700 649.050 843.600 656.400 ;
        RECT 862.200 654.000 864.000 662.400 ;
        RECT 886.500 657.600 888.300 662.400 ;
        RECT 886.500 656.400 891.600 657.600 ;
        RECT 860.700 652.800 864.000 654.000 ;
        RECT 860.700 649.050 861.600 652.800 ;
        RECT 871.950 651.450 876.000 652.050 ;
        RECT 863.100 649.050 864.900 650.850 ;
        RECT 869.100 649.050 870.900 650.850 ;
        RECT 871.950 649.950 876.450 651.450 ;
        RECT 832.950 646.950 835.050 649.050 ;
        RECT 835.950 646.950 838.050 649.050 ;
        RECT 838.950 646.950 841.050 649.050 ;
        RECT 841.950 646.950 844.050 649.050 ;
        RECT 859.950 646.950 862.050 649.050 ;
        RECT 862.950 646.950 865.050 649.050 ;
        RECT 865.950 646.950 868.050 649.050 ;
        RECT 868.950 646.950 871.050 649.050 ;
        RECT 827.550 644.550 832.050 646.050 ;
        RECT 836.100 645.150 837.900 646.950 ;
        RECT 828.000 643.950 832.050 644.550 ;
        RECT 842.700 639.600 843.600 646.950 ;
        RECT 797.400 627.600 799.200 633.600 ;
        RECT 812.400 627.600 814.200 633.600 ;
        RECT 818.400 627.600 820.200 639.600 ;
        RECT 833.400 638.700 841.200 639.600 ;
        RECT 833.400 627.600 835.200 638.700 ;
        RECT 839.400 627.600 841.200 638.700 ;
        RECT 842.400 627.600 844.200 639.600 ;
        RECT 860.700 634.800 861.600 646.950 ;
        RECT 866.100 645.150 867.900 646.950 ;
        RECT 875.550 646.050 876.450 649.950 ;
        RECT 881.100 649.050 882.900 650.850 ;
        RECT 887.100 649.050 888.900 650.850 ;
        RECT 890.700 649.050 891.600 656.400 ;
        RECT 880.950 646.950 883.050 649.050 ;
        RECT 883.950 646.950 886.050 649.050 ;
        RECT 886.950 646.950 889.050 649.050 ;
        RECT 889.950 646.950 892.050 649.050 ;
        RECT 871.950 644.550 876.450 646.050 ;
        RECT 884.100 645.150 885.900 646.950 ;
        RECT 871.950 643.950 876.000 644.550 ;
        RECT 862.950 642.450 865.050 643.050 ;
        RECT 880.950 642.450 883.050 643.050 ;
        RECT 862.950 641.550 883.050 642.450 ;
        RECT 862.950 640.950 865.050 641.550 ;
        RECT 880.950 640.950 883.050 641.550 ;
        RECT 890.700 639.600 891.600 646.950 ;
        RECT 881.400 638.700 889.200 639.600 ;
        RECT 860.700 633.900 867.300 634.800 ;
        RECT 860.700 633.600 861.600 633.900 ;
        RECT 859.800 627.600 861.600 633.600 ;
        RECT 865.800 633.600 867.300 633.900 ;
        RECT 865.800 627.600 867.600 633.600 ;
        RECT 881.400 627.600 883.200 638.700 ;
        RECT 887.400 627.600 889.200 638.700 ;
        RECT 890.400 627.600 892.200 639.600 ;
        RECT 13.800 611.400 15.600 623.400 ;
        RECT 19.800 617.400 21.600 623.400 ;
        RECT 14.400 604.050 15.300 611.400 ;
        RECT 17.100 604.050 18.900 605.850 ;
        RECT 13.950 601.950 16.050 604.050 ;
        RECT 16.950 601.950 19.050 604.050 ;
        RECT 14.400 594.600 15.300 601.950 ;
        RECT 20.700 597.300 21.600 617.400 ;
        RECT 37.800 612.600 39.600 623.400 ;
        RECT 37.800 611.400 42.900 612.600 ;
        RECT 45.300 612.300 47.100 623.400 ;
        RECT 52.800 612.300 54.600 623.400 ;
        RECT 40.800 610.500 42.900 611.400 ;
        RECT 43.800 611.400 47.100 612.300 ;
        RECT 22.950 609.450 25.050 610.050 ;
        RECT 22.950 608.550 36.450 609.450 ;
        RECT 22.950 607.950 25.050 608.550 ;
        RECT 35.550 606.450 36.450 608.550 ;
        RECT 43.800 606.900 45.000 611.400 ;
        RECT 49.800 611.100 54.600 612.300 ;
        RECT 67.800 612.600 69.600 623.400 ;
        RECT 67.800 611.400 72.600 612.600 ;
        RECT 49.800 610.200 51.900 611.100 ;
        RECT 70.500 610.500 72.600 611.400 ;
        RECT 75.300 611.400 77.100 623.400 ;
        RECT 82.800 612.300 84.600 623.400 ;
        RECT 85.950 618.450 88.050 619.050 ;
        RECT 85.950 617.550 93.450 618.450 ;
        RECT 85.950 616.950 88.050 617.550 ;
        RECT 80.100 611.400 84.600 612.300 ;
        RECT 46.500 609.300 51.900 610.200 ;
        RECT 75.300 609.900 76.500 611.400 ;
        RECT 46.500 607.200 48.300 609.300 ;
        RECT 75.000 609.000 76.500 609.900 ;
        RECT 80.100 609.300 82.200 611.400 ;
        RECT 92.550 610.050 93.450 617.550 ;
        RECT 95.400 612.300 97.200 623.400 ;
        RECT 101.400 612.300 103.200 623.400 ;
        RECT 95.400 611.400 103.200 612.300 ;
        RECT 104.400 611.400 106.200 623.400 ;
        RECT 122.400 617.400 124.200 623.400 ;
        RECT 75.000 606.900 75.900 609.000 ;
        RECT 92.550 608.550 97.050 610.050 ;
        RECT 93.000 607.950 97.050 608.550 ;
        RECT 35.550 605.700 39.450 606.450 ;
        RECT 43.500 606.300 45.600 606.900 ;
        RECT 35.550 605.550 39.900 605.700 ;
        RECT 22.950 601.950 25.050 604.050 ;
        RECT 38.100 603.900 39.900 605.550 ;
        RECT 43.500 604.800 46.650 606.300 ;
        RECT 23.100 600.150 24.900 601.950 ;
        RECT 37.950 601.800 40.050 603.900 ;
        RECT 42.900 602.100 44.700 603.900 ;
        RECT 42.750 600.000 44.850 602.100 ;
        RECT 45.750 598.200 46.650 604.800 ;
        RECT 48.000 604.200 49.800 606.000 ;
        RECT 47.700 602.100 49.800 604.200 ;
        RECT 68.100 604.050 69.900 605.850 ;
        RECT 73.800 604.800 75.900 606.900 ;
        RECT 76.800 607.500 78.900 607.800 ;
        RECT 76.800 605.700 80.700 607.500 ;
        RECT 52.500 601.800 54.600 603.900 ;
        RECT 55.950 603.450 58.050 604.050 ;
        RECT 67.950 603.450 70.050 604.050 ;
        RECT 74.400 603.900 76.800 604.800 ;
        RECT 55.950 602.550 70.050 603.450 ;
        RECT 55.950 601.950 58.050 602.550 ;
        RECT 67.950 601.950 70.050 602.550 ;
        RECT 52.500 601.200 54.300 601.800 ;
        RECT 72.600 601.200 74.400 603.000 ;
        RECT 47.700 600.000 54.300 601.200 ;
        RECT 47.700 599.100 49.800 600.000 ;
        RECT 72.750 599.100 74.850 601.200 ;
        RECT 17.100 596.400 24.600 597.300 ;
        RECT 17.100 595.500 18.900 596.400 ;
        RECT 14.400 592.800 17.100 594.600 ;
        RECT 15.300 588.600 17.100 592.800 ;
        RECT 22.800 588.600 24.600 596.400 ;
        RECT 40.200 595.800 42.300 597.900 ;
        RECT 43.500 596.100 46.650 598.200 ;
        RECT 47.550 597.300 49.350 599.100 ;
        RECT 75.750 598.200 76.800 603.900 ;
        RECT 77.700 603.900 79.500 604.500 ;
        RECT 98.100 604.050 99.900 605.850 ;
        RECT 104.700 604.050 105.600 611.400 ;
        RECT 122.400 604.050 123.600 617.400 ;
        RECT 143.700 612.600 145.500 623.400 ;
        RECT 143.700 611.400 147.300 612.600 ;
        RECT 143.100 604.050 144.900 605.850 ;
        RECT 146.400 604.050 147.300 611.400 ;
        RECT 163.800 611.400 165.600 623.400 ;
        RECT 169.800 617.400 171.600 623.400 ;
        RECT 149.100 604.050 150.900 605.850 ;
        RECT 163.800 604.050 165.000 611.400 ;
        RECT 170.400 610.500 171.600 617.400 ;
        RECT 185.700 612.600 187.500 623.400 ;
        RECT 185.700 611.400 189.300 612.600 ;
        RECT 165.900 609.600 171.600 610.500 ;
        RECT 165.900 608.700 167.850 609.600 ;
        RECT 82.500 603.900 84.600 604.050 ;
        RECT 77.700 602.700 84.600 603.900 ;
        RECT 82.500 601.950 84.600 602.700 ;
        RECT 94.950 601.950 97.050 604.050 ;
        RECT 97.950 601.950 100.050 604.050 ;
        RECT 100.950 601.950 103.050 604.050 ;
        RECT 103.950 601.950 106.050 604.050 ;
        RECT 118.950 601.950 121.050 604.050 ;
        RECT 121.950 601.950 124.050 604.050 ;
        RECT 124.950 601.950 127.050 604.050 ;
        RECT 142.950 601.950 145.050 604.050 ;
        RECT 145.950 601.950 148.050 604.050 ;
        RECT 148.950 601.950 151.050 604.050 ;
        RECT 163.800 601.950 166.050 604.050 ;
        RECT 37.800 594.600 42.300 595.800 ;
        RECT 37.800 588.600 39.600 594.600 ;
        RECT 45.600 594.000 46.650 596.100 ;
        RECT 50.250 597.000 52.350 597.600 ;
        RECT 50.250 595.500 54.600 597.000 ;
        RECT 70.500 595.500 72.600 596.700 ;
        RECT 73.800 596.100 76.800 598.200 ;
        RECT 77.700 599.400 79.500 601.200 ;
        RECT 82.800 600.150 84.600 601.950 ;
        RECT 95.100 600.150 96.900 601.950 ;
        RECT 101.100 600.150 102.900 601.950 ;
        RECT 77.700 597.300 79.800 599.400 ;
        RECT 77.700 596.400 84.000 597.300 ;
        RECT 53.100 594.600 54.600 595.500 ;
        RECT 45.600 588.600 47.400 594.000 ;
        RECT 52.800 588.600 54.600 594.600 ;
        RECT 67.800 594.600 72.600 595.500 ;
        RECT 75.600 594.600 76.800 596.100 ;
        RECT 82.800 594.600 84.000 596.400 ;
        RECT 104.700 594.600 105.600 601.950 ;
        RECT 119.100 600.150 120.900 601.950 ;
        RECT 122.400 596.700 123.600 601.950 ;
        RECT 125.100 600.150 126.900 601.950 ;
        RECT 122.400 595.800 126.600 596.700 ;
        RECT 67.800 588.600 69.600 594.600 ;
        RECT 75.300 588.600 77.100 594.600 ;
        RECT 82.800 588.600 84.600 594.600 ;
        RECT 100.500 593.400 105.600 594.600 ;
        RECT 100.500 588.600 102.300 593.400 ;
        RECT 124.800 588.600 126.600 595.800 ;
        RECT 146.400 591.600 147.300 601.950 ;
        RECT 163.800 594.600 165.000 601.950 ;
        RECT 166.950 597.300 167.850 608.700 ;
        RECT 170.100 604.050 171.900 605.850 ;
        RECT 185.100 604.050 186.900 605.850 ;
        RECT 188.400 604.050 189.300 611.400 ;
        RECT 195.150 611.400 196.950 623.400 ;
        RECT 203.550 617.400 205.350 623.400 ;
        RECT 203.550 616.500 204.750 617.400 ;
        RECT 211.350 616.500 213.150 623.400 ;
        RECT 219.150 617.400 220.950 623.400 ;
        RECT 199.950 614.400 204.750 616.500 ;
        RECT 207.450 615.450 214.050 616.500 ;
        RECT 207.450 614.700 209.250 615.450 ;
        RECT 212.250 614.700 214.050 615.450 ;
        RECT 219.150 615.300 223.050 617.400 ;
        RECT 203.550 613.500 204.750 614.400 ;
        RECT 216.450 613.800 218.250 614.400 ;
        RECT 203.550 612.300 211.050 613.500 ;
        RECT 209.250 611.700 211.050 612.300 ;
        RECT 211.950 612.900 218.250 613.800 ;
        RECT 195.150 610.500 196.050 611.400 ;
        RECT 211.950 610.800 212.850 612.900 ;
        RECT 216.450 612.600 218.250 612.900 ;
        RECT 219.150 612.600 221.850 614.400 ;
        RECT 219.150 611.700 220.050 612.600 ;
        RECT 204.450 610.500 212.850 610.800 ;
        RECT 195.150 609.900 212.850 610.500 ;
        RECT 214.950 610.800 220.050 611.700 ;
        RECT 220.950 610.800 223.050 611.700 ;
        RECT 226.650 611.400 228.450 623.400 ;
        RECT 245.400 617.400 247.200 623.400 ;
        RECT 195.150 609.300 206.250 609.900 ;
        RECT 191.100 604.050 192.900 605.850 ;
        RECT 169.950 601.950 172.050 604.050 ;
        RECT 184.950 601.950 187.050 604.050 ;
        RECT 187.950 601.950 190.050 604.050 ;
        RECT 190.950 601.950 193.050 604.050 ;
        RECT 165.900 596.400 167.850 597.300 ;
        RECT 165.900 595.500 171.600 596.400 ;
        RECT 145.800 588.600 147.600 591.600 ;
        RECT 163.800 588.600 165.600 594.600 ;
        RECT 170.400 591.600 171.600 595.500 ;
        RECT 188.400 591.600 189.300 601.950 ;
        RECT 195.150 594.600 196.050 609.300 ;
        RECT 204.450 609.000 206.250 609.300 ;
        RECT 196.950 601.950 199.050 604.050 ;
        RECT 205.950 602.400 208.050 604.050 ;
        RECT 197.100 600.150 198.900 601.950 ;
        RECT 200.100 601.200 208.050 602.400 ;
        RECT 200.100 600.600 201.900 601.200 ;
        RECT 198.000 599.400 198.900 600.150 ;
        RECT 203.100 599.400 204.900 600.000 ;
        RECT 198.000 598.200 204.900 599.400 ;
        RECT 214.950 598.200 215.850 610.800 ;
        RECT 220.950 609.600 225.150 610.800 ;
        RECT 224.250 607.800 226.050 609.600 ;
        RECT 227.250 604.050 228.450 611.400 ;
        RECT 245.850 604.050 247.050 617.400 ;
        RECT 263.400 612.300 265.200 623.400 ;
        RECT 270.900 612.300 272.700 623.400 ;
        RECT 278.400 612.600 280.200 623.400 ;
        RECT 298.500 612.600 300.300 623.400 ;
        RECT 319.800 617.400 321.600 623.400 ;
        RECT 263.400 611.100 268.200 612.300 ;
        RECT 270.900 611.400 274.200 612.300 ;
        RECT 266.100 610.200 268.200 611.100 ;
        RECT 266.100 609.300 271.500 610.200 ;
        RECT 269.700 607.200 271.500 609.300 ;
        RECT 273.000 606.900 274.200 611.400 ;
        RECT 275.100 611.400 280.200 612.600 ;
        RECT 296.700 611.400 300.300 612.600 ;
        RECT 275.100 610.500 277.200 611.400 ;
        RECT 272.400 606.300 274.500 606.900 ;
        RECT 286.950 606.450 289.050 607.050 ;
        RECT 251.100 604.050 252.900 605.850 ;
        RECT 268.200 604.200 270.000 606.000 ;
        RECT 271.350 604.800 274.500 606.300 ;
        RECT 278.550 605.700 289.050 606.450 ;
        RECT 278.100 605.550 289.050 605.700 ;
        RECT 223.950 603.750 228.450 604.050 ;
        RECT 222.150 601.950 228.450 603.750 ;
        RECT 241.950 601.950 244.050 604.050 ;
        RECT 244.950 601.950 247.050 604.050 ;
        RECT 247.950 601.950 250.050 604.050 ;
        RECT 250.950 601.950 253.050 604.050 ;
        RECT 203.850 597.000 215.850 598.200 ;
        RECT 203.850 595.200 204.900 597.000 ;
        RECT 214.050 596.400 215.850 597.000 ;
        RECT 169.800 588.600 171.600 591.600 ;
        RECT 187.800 588.600 189.600 591.600 ;
        RECT 195.150 588.600 196.950 594.600 ;
        RECT 199.950 592.500 202.050 594.600 ;
        RECT 203.550 593.400 205.350 595.200 ;
        RECT 227.250 594.600 228.450 601.950 ;
        RECT 242.100 600.150 243.900 601.950 ;
        RECT 244.950 597.750 246.150 601.950 ;
        RECT 248.100 600.150 249.900 601.950 ;
        RECT 263.400 601.800 265.500 603.900 ;
        RECT 268.200 602.100 270.300 604.200 ;
        RECT 263.700 601.200 265.500 601.800 ;
        RECT 263.700 600.000 270.300 601.200 ;
        RECT 268.200 599.100 270.300 600.000 ;
        RECT 242.400 596.700 246.150 597.750 ;
        RECT 265.650 597.000 267.750 597.600 ;
        RECT 268.650 597.300 270.450 599.100 ;
        RECT 271.350 598.200 272.250 604.800 ;
        RECT 278.100 603.900 279.900 605.550 ;
        RECT 286.950 604.950 289.050 605.550 ;
        RECT 293.100 604.050 294.900 605.850 ;
        RECT 296.700 604.050 297.600 611.400 ;
        RECT 299.100 604.050 300.900 605.850 ;
        RECT 320.400 604.050 321.600 617.400 ;
        RECT 337.800 611.400 339.600 623.400 ;
        RECT 343.800 617.400 345.600 623.400 ;
        RECT 338.400 604.050 339.300 611.400 ;
        RECT 341.100 604.050 342.900 605.850 ;
        RECT 273.300 602.100 275.100 603.900 ;
        RECT 273.150 600.000 275.250 602.100 ;
        RECT 277.950 601.800 280.050 603.900 ;
        RECT 292.950 601.950 295.050 604.050 ;
        RECT 295.950 601.950 298.050 604.050 ;
        RECT 298.950 601.950 301.050 604.050 ;
        RECT 316.950 601.950 319.050 604.050 ;
        RECT 319.950 601.950 322.050 604.050 ;
        RECT 322.950 601.950 325.050 604.050 ;
        RECT 337.950 601.950 340.050 604.050 ;
        RECT 340.950 601.950 343.050 604.050 ;
        RECT 242.400 594.600 243.600 596.700 ;
        RECT 263.400 595.500 267.750 597.000 ;
        RECT 271.350 596.100 274.500 598.200 ;
        RECT 206.850 593.550 208.650 594.300 ;
        RECT 220.950 593.700 223.050 594.600 ;
        RECT 206.850 592.500 211.800 593.550 ;
        RECT 201.000 591.600 202.050 592.500 ;
        RECT 210.750 591.600 211.800 592.500 ;
        RECT 219.300 592.500 223.050 593.700 ;
        RECT 219.300 591.600 220.350 592.500 ;
        RECT 201.000 590.700 204.750 591.600 ;
        RECT 202.950 588.600 204.750 590.700 ;
        RECT 210.750 588.600 212.550 591.600 ;
        RECT 218.550 588.600 220.350 591.600 ;
        RECT 226.650 588.600 228.450 594.600 ;
        RECT 241.800 588.600 243.600 594.600 ;
        RECT 244.800 593.700 252.600 595.050 ;
        RECT 244.800 588.600 246.600 593.700 ;
        RECT 250.800 588.600 252.600 593.700 ;
        RECT 263.400 594.600 264.900 595.500 ;
        RECT 263.400 588.600 265.200 594.600 ;
        RECT 271.350 594.000 272.400 596.100 ;
        RECT 275.700 595.800 277.800 597.900 ;
        RECT 275.700 594.600 280.200 595.800 ;
        RECT 270.600 588.600 272.400 594.000 ;
        RECT 278.400 588.600 280.200 594.600 ;
        RECT 296.700 591.600 297.600 601.950 ;
        RECT 317.100 600.150 318.900 601.950 ;
        RECT 320.400 596.700 321.600 601.950 ;
        RECT 323.100 600.150 324.900 601.950 ;
        RECT 317.400 595.800 321.600 596.700 ;
        RECT 322.950 597.450 325.050 598.050 ;
        RECT 328.950 597.450 331.050 598.050 ;
        RECT 322.950 596.550 331.050 597.450 ;
        RECT 322.950 595.950 325.050 596.550 ;
        RECT 328.950 595.950 331.050 596.550 ;
        RECT 296.400 588.600 298.200 591.600 ;
        RECT 317.400 588.600 319.200 595.800 ;
        RECT 338.400 594.600 339.300 601.950 ;
        RECT 344.700 597.300 345.600 617.400 ;
        RECT 362.400 617.400 364.200 623.400 ;
        RECT 362.400 604.050 363.600 617.400 ;
        RECT 380.400 612.600 382.200 623.400 ;
        RECT 386.400 622.500 394.200 623.400 ;
        RECT 386.400 612.600 388.200 622.500 ;
        RECT 380.400 611.700 388.200 612.600 ;
        RECT 389.400 610.500 391.200 621.600 ;
        RECT 392.400 611.400 394.200 622.500 ;
        RECT 409.800 617.400 411.600 623.400 ;
        RECT 364.950 609.450 367.050 610.050 ;
        RECT 373.950 609.450 376.050 610.050 ;
        RECT 382.950 609.450 385.050 610.050 ;
        RECT 364.950 608.550 385.050 609.450 ;
        RECT 364.950 607.950 367.050 608.550 ;
        RECT 373.950 607.950 376.050 608.550 ;
        RECT 382.950 607.950 385.050 608.550 ;
        RECT 386.100 609.600 391.200 610.500 ;
        RECT 383.100 604.050 384.900 605.850 ;
        RECT 386.100 604.050 387.000 609.600 ;
        RECT 389.100 604.050 390.900 605.850 ;
        RECT 410.400 604.050 411.600 617.400 ;
        RECT 430.800 611.400 432.600 623.400 ;
        RECT 436.800 617.400 438.600 623.400 ;
        RECT 413.100 604.050 414.900 605.850 ;
        RECT 430.800 604.050 432.000 611.400 ;
        RECT 437.400 610.500 438.600 617.400 ;
        RECT 432.900 609.600 438.600 610.500 ;
        RECT 451.800 611.400 453.600 623.400 ;
        RECT 457.800 617.400 459.600 623.400 ;
        RECT 476.400 617.400 478.200 623.400 ;
        RECT 432.900 608.700 434.850 609.600 ;
        RECT 346.950 601.950 349.050 604.050 ;
        RECT 358.950 601.950 361.050 604.050 ;
        RECT 361.950 601.950 364.050 604.050 ;
        RECT 364.950 601.950 367.050 604.050 ;
        RECT 379.950 601.950 382.050 604.050 ;
        RECT 382.950 601.950 385.050 604.050 ;
        RECT 385.950 601.950 388.050 604.050 ;
        RECT 388.950 601.950 391.050 604.050 ;
        RECT 391.950 601.950 394.050 604.050 ;
        RECT 409.950 601.950 412.050 604.050 ;
        RECT 412.950 601.950 415.050 604.050 ;
        RECT 430.800 601.950 433.050 604.050 ;
        RECT 347.100 600.150 348.900 601.950 ;
        RECT 359.100 600.150 360.900 601.950 ;
        RECT 341.100 596.400 348.600 597.300 ;
        RECT 341.100 595.500 342.900 596.400 ;
        RECT 338.400 592.800 341.100 594.600 ;
        RECT 339.300 588.600 341.100 592.800 ;
        RECT 346.800 588.600 348.600 596.400 ;
        RECT 362.400 596.700 363.600 601.950 ;
        RECT 365.100 600.150 366.900 601.950 ;
        RECT 380.100 600.150 381.900 601.950 ;
        RECT 362.400 595.800 366.600 596.700 ;
        RECT 364.800 588.600 366.600 595.800 ;
        RECT 385.950 594.600 387.000 601.950 ;
        RECT 392.100 600.150 393.900 601.950 ;
        RECT 385.200 588.600 387.000 594.600 ;
        RECT 410.400 591.600 411.600 601.950 ;
        RECT 409.800 588.600 411.600 591.600 ;
        RECT 430.800 594.600 432.000 601.950 ;
        RECT 433.950 597.300 434.850 608.700 ;
        RECT 437.100 604.050 438.900 605.850 ;
        RECT 451.800 604.050 453.000 611.400 ;
        RECT 458.400 610.500 459.600 617.400 ;
        RECT 453.900 609.600 459.600 610.500 ;
        RECT 453.900 608.700 455.850 609.600 ;
        RECT 436.950 601.950 439.050 604.050 ;
        RECT 451.800 601.950 454.050 604.050 ;
        RECT 432.900 596.400 434.850 597.300 ;
        RECT 432.900 595.500 438.600 596.400 ;
        RECT 430.800 588.600 432.600 594.600 ;
        RECT 437.400 591.600 438.600 595.500 ;
        RECT 436.800 588.600 438.600 591.600 ;
        RECT 451.800 594.600 453.000 601.950 ;
        RECT 454.950 597.300 455.850 608.700 ;
        RECT 458.100 604.050 459.900 605.850 ;
        RECT 476.850 604.050 478.050 617.400 ;
        RECT 486.150 611.400 487.950 623.400 ;
        RECT 494.550 617.400 496.350 623.400 ;
        RECT 494.550 616.500 495.750 617.400 ;
        RECT 502.350 616.500 504.150 623.400 ;
        RECT 510.150 617.400 511.950 623.400 ;
        RECT 490.950 614.400 495.750 616.500 ;
        RECT 498.450 615.450 505.050 616.500 ;
        RECT 498.450 614.700 500.250 615.450 ;
        RECT 503.250 614.700 505.050 615.450 ;
        RECT 510.150 615.300 514.050 617.400 ;
        RECT 494.550 613.500 495.750 614.400 ;
        RECT 507.450 613.800 509.250 614.400 ;
        RECT 494.550 612.300 502.050 613.500 ;
        RECT 500.250 611.700 502.050 612.300 ;
        RECT 502.950 612.900 509.250 613.800 ;
        RECT 486.150 610.500 487.050 611.400 ;
        RECT 502.950 610.800 503.850 612.900 ;
        RECT 507.450 612.600 509.250 612.900 ;
        RECT 510.150 612.600 512.850 614.400 ;
        RECT 510.150 611.700 511.050 612.600 ;
        RECT 495.450 610.500 503.850 610.800 ;
        RECT 486.150 609.900 503.850 610.500 ;
        RECT 505.950 610.800 511.050 611.700 ;
        RECT 511.950 610.800 514.050 611.700 ;
        RECT 517.650 611.400 519.450 623.400 ;
        RECT 539.400 617.400 541.200 623.400 ;
        RECT 486.150 609.300 497.250 609.900 ;
        RECT 482.100 604.050 483.900 605.850 ;
        RECT 457.950 601.950 460.050 604.050 ;
        RECT 472.950 601.950 475.050 604.050 ;
        RECT 475.950 601.950 478.050 604.050 ;
        RECT 478.950 601.950 481.050 604.050 ;
        RECT 481.950 601.950 484.050 604.050 ;
        RECT 473.100 600.150 474.900 601.950 ;
        RECT 475.950 597.750 477.150 601.950 ;
        RECT 479.100 600.150 480.900 601.950 ;
        RECT 453.900 596.400 455.850 597.300 ;
        RECT 473.400 596.700 477.150 597.750 ;
        RECT 453.900 595.500 459.600 596.400 ;
        RECT 451.800 588.600 453.600 594.600 ;
        RECT 458.400 591.600 459.600 595.500 ;
        RECT 473.400 594.600 474.600 596.700 ;
        RECT 457.800 588.600 459.600 591.600 ;
        RECT 472.800 588.600 474.600 594.600 ;
        RECT 475.800 593.700 483.600 595.050 ;
        RECT 475.800 588.600 477.600 593.700 ;
        RECT 481.800 588.600 483.600 593.700 ;
        RECT 486.150 594.600 487.050 609.300 ;
        RECT 495.450 609.000 497.250 609.300 ;
        RECT 487.950 601.950 490.050 604.050 ;
        RECT 496.950 602.400 499.050 604.050 ;
        RECT 488.100 600.150 489.900 601.950 ;
        RECT 491.100 601.200 499.050 602.400 ;
        RECT 491.100 600.600 492.900 601.200 ;
        RECT 489.000 599.400 489.900 600.150 ;
        RECT 494.100 599.400 495.900 600.000 ;
        RECT 489.000 598.200 495.900 599.400 ;
        RECT 505.950 598.200 506.850 610.800 ;
        RECT 511.950 609.600 516.150 610.800 ;
        RECT 515.250 607.800 517.050 609.600 ;
        RECT 518.250 604.050 519.450 611.400 ;
        RECT 539.850 604.050 541.050 617.400 ;
        RECT 549.150 611.400 550.950 623.400 ;
        RECT 557.550 617.400 559.350 623.400 ;
        RECT 557.550 616.500 558.750 617.400 ;
        RECT 565.350 616.500 567.150 623.400 ;
        RECT 573.150 617.400 574.950 623.400 ;
        RECT 553.950 614.400 558.750 616.500 ;
        RECT 561.450 615.450 568.050 616.500 ;
        RECT 561.450 614.700 563.250 615.450 ;
        RECT 566.250 614.700 568.050 615.450 ;
        RECT 573.150 615.300 577.050 617.400 ;
        RECT 557.550 613.500 558.750 614.400 ;
        RECT 570.450 613.800 572.250 614.400 ;
        RECT 557.550 612.300 565.050 613.500 ;
        RECT 563.250 611.700 565.050 612.300 ;
        RECT 565.950 612.900 572.250 613.800 ;
        RECT 549.150 610.500 550.050 611.400 ;
        RECT 565.950 610.800 566.850 612.900 ;
        RECT 570.450 612.600 572.250 612.900 ;
        RECT 573.150 612.600 575.850 614.400 ;
        RECT 573.150 611.700 574.050 612.600 ;
        RECT 558.450 610.500 566.850 610.800 ;
        RECT 549.150 609.900 566.850 610.500 ;
        RECT 568.950 610.800 574.050 611.700 ;
        RECT 574.950 610.800 577.050 611.700 ;
        RECT 580.650 611.400 582.450 623.400 ;
        RECT 598.800 617.400 600.600 623.400 ;
        RECT 620.400 617.400 622.200 623.400 ;
        RECT 643.800 617.400 645.600 623.400 ;
        RECT 664.800 617.400 666.600 623.400 ;
        RECT 683.400 617.400 685.200 623.400 ;
        RECT 549.150 609.300 560.250 609.900 ;
        RECT 545.100 604.050 546.900 605.850 ;
        RECT 514.950 603.750 519.450 604.050 ;
        RECT 513.150 601.950 519.450 603.750 ;
        RECT 535.950 601.950 538.050 604.050 ;
        RECT 538.950 601.950 541.050 604.050 ;
        RECT 541.950 601.950 544.050 604.050 ;
        RECT 544.950 601.950 547.050 604.050 ;
        RECT 494.850 597.000 506.850 598.200 ;
        RECT 494.850 595.200 495.900 597.000 ;
        RECT 505.050 596.400 506.850 597.000 ;
        RECT 486.150 588.600 487.950 594.600 ;
        RECT 490.950 592.500 493.050 594.600 ;
        RECT 494.550 593.400 496.350 595.200 ;
        RECT 518.250 594.600 519.450 601.950 ;
        RECT 520.950 600.450 523.050 601.050 ;
        RECT 532.950 600.450 535.050 601.050 ;
        RECT 520.950 599.550 535.050 600.450 ;
        RECT 536.100 600.150 537.900 601.950 ;
        RECT 520.950 598.950 523.050 599.550 ;
        RECT 532.950 598.950 535.050 599.550 ;
        RECT 538.950 597.750 540.150 601.950 ;
        RECT 542.100 600.150 543.900 601.950 ;
        RECT 536.400 596.700 540.150 597.750 ;
        RECT 536.400 594.600 537.600 596.700 ;
        RECT 497.850 593.550 499.650 594.300 ;
        RECT 511.950 593.700 514.050 594.600 ;
        RECT 497.850 592.500 502.800 593.550 ;
        RECT 492.000 591.600 493.050 592.500 ;
        RECT 501.750 591.600 502.800 592.500 ;
        RECT 510.300 592.500 514.050 593.700 ;
        RECT 510.300 591.600 511.350 592.500 ;
        RECT 492.000 590.700 495.750 591.600 ;
        RECT 493.950 588.600 495.750 590.700 ;
        RECT 501.750 588.600 503.550 591.600 ;
        RECT 509.550 588.600 511.350 591.600 ;
        RECT 517.650 588.600 519.450 594.600 ;
        RECT 535.800 588.600 537.600 594.600 ;
        RECT 538.800 593.700 546.600 595.050 ;
        RECT 538.800 588.600 540.600 593.700 ;
        RECT 544.800 588.600 546.600 593.700 ;
        RECT 549.150 594.600 550.050 609.300 ;
        RECT 558.450 609.000 560.250 609.300 ;
        RECT 550.950 601.950 553.050 604.050 ;
        RECT 559.950 602.400 562.050 604.050 ;
        RECT 551.100 600.150 552.900 601.950 ;
        RECT 554.100 601.200 562.050 602.400 ;
        RECT 554.100 600.600 555.900 601.200 ;
        RECT 552.000 599.400 552.900 600.150 ;
        RECT 557.100 599.400 558.900 600.000 ;
        RECT 552.000 598.200 558.900 599.400 ;
        RECT 568.950 598.200 569.850 610.800 ;
        RECT 574.950 609.600 579.150 610.800 ;
        RECT 578.250 607.800 580.050 609.600 ;
        RECT 581.250 604.050 582.450 611.400 ;
        RECT 599.400 604.050 600.600 617.400 ;
        RECT 610.950 609.450 613.050 610.050 ;
        RECT 616.950 609.450 619.050 610.050 ;
        RECT 610.950 608.550 619.050 609.450 ;
        RECT 610.950 607.950 613.050 608.550 ;
        RECT 616.950 607.950 619.050 608.550 ;
        RECT 613.950 606.450 616.050 607.050 ;
        RECT 608.550 605.550 616.050 606.450 ;
        RECT 577.950 603.750 582.450 604.050 ;
        RECT 576.150 601.950 582.450 603.750 ;
        RECT 595.950 601.950 598.050 604.050 ;
        RECT 598.950 601.950 601.050 604.050 ;
        RECT 601.950 601.950 604.050 604.050 ;
        RECT 557.850 597.000 569.850 598.200 ;
        RECT 557.850 595.200 558.900 597.000 ;
        RECT 568.050 596.400 569.850 597.000 ;
        RECT 549.150 588.600 550.950 594.600 ;
        RECT 553.950 592.500 556.050 594.600 ;
        RECT 557.550 593.400 559.350 595.200 ;
        RECT 581.250 594.600 582.450 601.950 ;
        RECT 596.100 600.150 597.900 601.950 ;
        RECT 599.400 596.700 600.600 601.950 ;
        RECT 602.100 600.150 603.900 601.950 ;
        RECT 608.550 601.050 609.450 605.550 ;
        RECT 613.950 604.950 616.050 605.550 ;
        RECT 620.850 604.050 622.050 617.400 ;
        RECT 628.950 606.450 631.050 610.050 ;
        RECT 634.950 607.950 637.050 610.050 ;
        RECT 628.950 606.000 633.450 606.450 ;
        RECT 626.100 604.050 627.900 605.850 ;
        RECT 629.550 605.550 633.450 606.000 ;
        RECT 616.950 601.950 619.050 604.050 ;
        RECT 619.950 601.950 622.050 604.050 ;
        RECT 622.950 601.950 625.050 604.050 ;
        RECT 625.950 601.950 628.050 604.050 ;
        RECT 604.950 599.550 609.450 601.050 ;
        RECT 617.100 600.150 618.900 601.950 ;
        RECT 604.950 598.950 609.000 599.550 ;
        RECT 619.950 597.750 621.150 601.950 ;
        RECT 623.100 600.150 624.900 601.950 ;
        RECT 632.550 601.050 633.450 605.550 ;
        RECT 628.950 599.550 633.450 601.050 ;
        RECT 628.950 598.950 633.000 599.550 ;
        RECT 635.550 598.050 636.450 607.950 ;
        RECT 644.400 604.050 645.600 617.400 ;
        RECT 659.100 604.050 660.900 605.850 ;
        RECT 664.950 604.050 666.150 617.400 ;
        RECT 683.400 610.500 684.600 617.400 ;
        RECT 689.400 611.400 691.200 623.400 ;
        RECT 683.400 609.600 689.100 610.500 ;
        RECT 687.150 608.700 689.100 609.600 ;
        RECT 683.100 604.050 684.900 605.850 ;
        RECT 640.950 601.950 643.050 604.050 ;
        RECT 643.950 601.950 646.050 604.050 ;
        RECT 646.950 601.950 649.050 604.050 ;
        RECT 658.950 601.950 661.050 604.050 ;
        RECT 661.950 601.950 664.050 604.050 ;
        RECT 664.950 601.950 667.050 604.050 ;
        RECT 667.950 601.950 670.050 604.050 ;
        RECT 682.950 601.950 685.050 604.050 ;
        RECT 641.100 600.150 642.900 601.950 ;
        RECT 560.850 593.550 562.650 594.300 ;
        RECT 574.950 593.700 577.050 594.600 ;
        RECT 560.850 592.500 565.800 593.550 ;
        RECT 555.000 591.600 556.050 592.500 ;
        RECT 564.750 591.600 565.800 592.500 ;
        RECT 573.300 592.500 577.050 593.700 ;
        RECT 573.300 591.600 574.350 592.500 ;
        RECT 555.000 590.700 558.750 591.600 ;
        RECT 556.950 588.600 558.750 590.700 ;
        RECT 564.750 588.600 566.550 591.600 ;
        RECT 572.550 588.600 574.350 591.600 ;
        RECT 580.650 588.600 582.450 594.600 ;
        RECT 596.400 595.800 600.600 596.700 ;
        RECT 617.400 596.700 621.150 597.750 ;
        RECT 596.400 588.600 598.200 595.800 ;
        RECT 617.400 594.600 618.600 596.700 ;
        RECT 634.950 595.950 637.050 598.050 ;
        RECT 644.400 596.700 645.600 601.950 ;
        RECT 647.100 600.150 648.900 601.950 ;
        RECT 662.100 600.150 663.900 601.950 ;
        RECT 665.850 597.750 667.050 601.950 ;
        RECT 668.100 600.150 669.900 601.950 ;
        RECT 665.850 596.700 669.600 597.750 ;
        RECT 641.400 595.800 645.600 596.700 ;
        RECT 616.800 588.600 618.600 594.600 ;
        RECT 619.800 593.700 627.600 595.050 ;
        RECT 619.800 588.600 621.600 593.700 ;
        RECT 625.800 588.600 627.600 593.700 ;
        RECT 641.400 588.600 643.200 595.800 ;
        RECT 659.400 593.700 667.200 595.050 ;
        RECT 659.400 588.600 661.200 593.700 ;
        RECT 665.400 588.600 667.200 593.700 ;
        RECT 668.400 594.600 669.600 596.700 ;
        RECT 687.150 597.300 688.050 608.700 ;
        RECT 690.000 604.050 691.200 611.400 ;
        RECT 704.400 617.400 706.200 623.400 ;
        RECT 704.400 610.500 705.600 617.400 ;
        RECT 710.400 611.400 712.200 623.400 ;
        RECT 704.400 609.600 710.100 610.500 ;
        RECT 708.150 608.700 710.100 609.600 ;
        RECT 699.000 606.450 703.050 607.050 ;
        RECT 688.950 601.950 691.200 604.050 ;
        RECT 687.150 596.400 689.100 597.300 ;
        RECT 683.400 595.500 689.100 596.400 ;
        RECT 668.400 588.600 670.200 594.600 ;
        RECT 683.400 591.600 684.600 595.500 ;
        RECT 690.000 594.600 691.200 601.950 ;
        RECT 698.550 604.950 703.050 606.450 ;
        RECT 698.550 601.050 699.450 604.950 ;
        RECT 704.100 604.050 705.900 605.850 ;
        RECT 703.950 601.950 706.050 604.050 ;
        RECT 698.550 599.550 703.050 601.050 ;
        RECT 699.000 598.950 703.050 599.550 ;
        RECT 708.150 597.300 709.050 608.700 ;
        RECT 711.000 604.050 712.200 611.400 ;
        RECT 728.400 617.400 730.200 623.400 ;
        RECT 749.400 617.400 751.200 623.400 ;
        RECT 718.950 609.450 721.050 610.050 ;
        RECT 724.950 609.450 727.050 610.050 ;
        RECT 718.950 608.550 727.050 609.450 ;
        RECT 718.950 607.950 721.050 608.550 ;
        RECT 724.950 607.950 727.050 608.550 ;
        RECT 728.400 604.050 729.600 617.400 ;
        RECT 749.700 617.100 751.200 617.400 ;
        RECT 755.400 617.400 757.200 623.400 ;
        RECT 760.950 618.450 763.050 619.050 ;
        RECT 766.950 618.450 769.050 619.050 ;
        RECT 760.950 617.550 769.050 618.450 ;
        RECT 755.400 617.100 756.300 617.400 ;
        RECT 749.700 616.200 756.300 617.100 ;
        RECT 760.950 616.950 763.050 617.550 ;
        RECT 766.950 616.950 769.050 617.550 ;
        RECT 739.950 609.450 742.050 610.050 ;
        RECT 751.950 609.450 754.050 610.050 ;
        RECT 739.950 608.550 754.050 609.450 ;
        RECT 739.950 607.950 742.050 608.550 ;
        RECT 751.950 607.950 754.050 608.550 ;
        RECT 733.950 606.450 738.000 607.050 ;
        RECT 741.000 606.450 745.050 607.050 ;
        RECT 733.950 604.950 738.450 606.450 ;
        RECT 709.950 601.950 712.200 604.050 ;
        RECT 724.950 601.950 727.050 604.050 ;
        RECT 727.950 601.950 730.050 604.050 ;
        RECT 730.950 601.950 733.050 604.050 ;
        RECT 708.150 596.400 710.100 597.300 ;
        RECT 683.400 588.600 685.200 591.600 ;
        RECT 689.400 588.600 691.200 594.600 ;
        RECT 704.400 595.500 710.100 596.400 ;
        RECT 704.400 591.600 705.600 595.500 ;
        RECT 711.000 594.600 712.200 601.950 ;
        RECT 725.100 600.150 726.900 601.950 ;
        RECT 728.400 596.700 729.600 601.950 ;
        RECT 731.100 600.150 732.900 601.950 ;
        RECT 737.550 600.450 738.450 604.950 ;
        RECT 734.550 600.000 738.450 600.450 ;
        RECT 733.950 599.550 738.450 600.000 ;
        RECT 740.550 604.950 745.050 606.450 ;
        RECT 740.550 601.050 741.450 604.950 ;
        RECT 749.100 604.050 750.900 605.850 ;
        RECT 755.400 604.050 756.300 616.200 ;
        RECT 770.400 612.600 772.200 623.400 ;
        RECT 776.400 622.500 784.200 623.400 ;
        RECT 776.400 612.600 778.200 622.500 ;
        RECT 770.400 611.700 778.200 612.600 ;
        RECT 779.400 610.500 781.200 621.600 ;
        RECT 782.400 611.400 784.200 622.500 ;
        RECT 800.400 617.400 802.200 623.400 ;
        RECT 821.400 617.400 823.200 623.400 ;
        RECT 842.400 617.400 844.200 623.400 ;
        RECT 776.100 609.600 781.200 610.500 ;
        RECT 757.950 606.450 760.050 607.050 ;
        RECT 757.950 605.550 765.450 606.450 ;
        RECT 757.950 604.950 760.050 605.550 ;
        RECT 745.950 601.950 748.050 604.050 ;
        RECT 748.950 601.950 751.050 604.050 ;
        RECT 751.950 601.950 754.050 604.050 ;
        RECT 754.950 601.950 757.050 604.050 ;
        RECT 740.550 599.550 745.050 601.050 ;
        RECT 746.100 600.150 747.900 601.950 ;
        RECT 752.100 600.150 753.900 601.950 ;
        RECT 728.400 595.800 732.600 596.700 ;
        RECT 733.950 595.950 736.050 599.550 ;
        RECT 741.000 598.950 745.050 599.550 ;
        RECT 755.400 598.200 756.300 601.950 ;
        RECT 764.550 601.050 765.450 605.550 ;
        RECT 773.100 604.050 774.900 605.850 ;
        RECT 776.100 604.050 777.000 609.600 ;
        RECT 790.950 609.450 793.050 610.050 ;
        RECT 796.950 609.450 799.050 613.050 ;
        RECT 790.950 609.000 799.050 609.450 ;
        RECT 790.950 608.550 798.450 609.000 ;
        RECT 790.950 607.950 793.050 608.550 ;
        RECT 784.950 606.450 787.050 607.050 ;
        RECT 790.950 606.450 793.050 606.900 ;
        RECT 779.100 604.050 780.900 605.850 ;
        RECT 784.950 605.550 793.050 606.450 ;
        RECT 784.950 604.950 787.050 605.550 ;
        RECT 790.950 604.800 793.050 605.550 ;
        RECT 797.100 604.050 798.900 605.850 ;
        RECT 800.400 604.050 801.600 617.400 ;
        RECT 821.850 604.050 823.050 617.400 ;
        RECT 842.700 617.100 844.200 617.400 ;
        RECT 848.400 617.400 850.200 623.400 ;
        RECT 848.400 617.100 849.300 617.400 ;
        RECT 842.700 616.200 849.300 617.100 ;
        RECT 834.000 606.450 838.050 607.050 ;
        RECT 827.100 604.050 828.900 605.850 ;
        RECT 833.550 604.950 838.050 606.450 ;
        RECT 769.950 601.950 772.050 604.050 ;
        RECT 772.950 601.950 775.050 604.050 ;
        RECT 775.950 601.950 778.050 604.050 ;
        RECT 778.950 601.950 781.050 604.050 ;
        RECT 781.950 601.950 784.050 604.050 ;
        RECT 796.950 601.950 799.050 604.050 ;
        RECT 799.950 601.950 802.050 604.050 ;
        RECT 817.950 601.950 820.050 604.050 ;
        RECT 820.950 601.950 823.050 604.050 ;
        RECT 823.950 601.950 826.050 604.050 ;
        RECT 826.950 601.950 829.050 604.050 ;
        RECT 764.550 599.550 769.050 601.050 ;
        RECT 770.100 600.150 771.900 601.950 ;
        RECT 765.000 598.950 769.050 599.550 ;
        RECT 753.000 597.000 756.300 598.200 ;
        RECT 704.400 588.600 706.200 591.600 ;
        RECT 710.400 588.600 712.200 594.600 ;
        RECT 730.800 588.600 732.600 595.800 ;
        RECT 753.000 588.600 754.800 597.000 ;
        RECT 775.950 594.600 777.000 601.950 ;
        RECT 782.100 600.150 783.900 601.950 ;
        RECT 775.200 588.600 777.000 594.600 ;
        RECT 784.950 594.450 787.050 595.050 ;
        RECT 796.950 594.450 799.050 595.050 ;
        RECT 784.950 593.550 799.050 594.450 ;
        RECT 784.950 592.950 787.050 593.550 ;
        RECT 796.950 592.950 799.050 593.550 ;
        RECT 800.400 591.600 801.600 601.950 ;
        RECT 818.100 600.150 819.900 601.950 ;
        RECT 820.950 597.750 822.150 601.950 ;
        RECT 824.100 600.150 825.900 601.950 ;
        RECT 833.550 601.050 834.450 604.950 ;
        RECT 842.100 604.050 843.900 605.850 ;
        RECT 848.400 604.050 849.300 616.200 ;
        RECT 865.800 611.400 867.600 623.400 ;
        RECT 868.800 612.300 870.600 623.400 ;
        RECT 874.800 612.300 876.600 623.400 ;
        RECT 889.800 617.400 891.600 623.400 ;
        RECT 868.800 611.400 876.600 612.300 ;
        RECT 866.400 604.050 867.300 611.400 ;
        RECT 868.950 609.450 871.050 610.050 ;
        RECT 886.950 609.450 889.050 610.050 ;
        RECT 868.950 608.550 889.050 609.450 ;
        RECT 868.950 607.950 871.050 608.550 ;
        RECT 886.950 607.950 889.050 608.550 ;
        RECT 872.100 604.050 873.900 605.850 ;
        RECT 890.400 604.050 891.600 617.400 ;
        RECT 893.100 604.050 894.900 605.850 ;
        RECT 838.950 601.950 841.050 604.050 ;
        RECT 841.950 601.950 844.050 604.050 ;
        RECT 844.950 601.950 847.050 604.050 ;
        RECT 847.950 601.950 850.050 604.050 ;
        RECT 865.950 601.950 868.050 604.050 ;
        RECT 868.950 601.950 871.050 604.050 ;
        RECT 871.950 601.950 874.050 604.050 ;
        RECT 874.950 601.950 877.050 604.050 ;
        RECT 889.950 601.950 892.050 604.050 ;
        RECT 892.950 601.950 895.050 604.050 ;
        RECT 829.950 599.550 834.450 601.050 ;
        RECT 839.100 600.150 840.900 601.950 ;
        RECT 845.100 600.150 846.900 601.950 ;
        RECT 829.950 598.950 834.000 599.550 ;
        RECT 848.400 598.200 849.300 601.950 ;
        RECT 818.400 596.700 822.150 597.750 ;
        RECT 846.000 597.000 849.300 598.200 ;
        RECT 853.950 597.450 856.050 597.900 ;
        RECT 859.950 597.450 862.050 598.050 ;
        RECT 818.400 594.600 819.600 596.700 ;
        RECT 800.400 588.600 802.200 591.600 ;
        RECT 817.800 588.600 819.600 594.600 ;
        RECT 820.800 593.700 828.600 595.050 ;
        RECT 820.800 588.600 822.600 593.700 ;
        RECT 826.800 588.600 828.600 593.700 ;
        RECT 846.000 588.600 847.800 597.000 ;
        RECT 853.950 596.550 862.050 597.450 ;
        RECT 853.950 595.800 856.050 596.550 ;
        RECT 859.950 595.950 862.050 596.550 ;
        RECT 866.400 594.600 867.300 601.950 ;
        RECT 869.100 600.150 870.900 601.950 ;
        RECT 875.100 600.150 876.900 601.950 ;
        RECT 866.400 593.400 871.500 594.600 ;
        RECT 869.700 588.600 871.500 593.400 ;
        RECT 890.400 591.600 891.600 601.950 ;
        RECT 889.800 588.600 891.600 591.600 ;
        RECT 16.800 581.400 18.600 584.400 ;
        RECT 17.400 571.050 18.300 581.400 ;
        RECT 35.400 577.200 37.200 584.400 ;
        RECT 58.800 578.400 60.600 584.400 ;
        RECT 35.400 576.300 39.600 577.200 ;
        RECT 35.100 571.050 36.900 572.850 ;
        RECT 38.400 571.050 39.600 576.300 ;
        RECT 59.400 576.300 60.600 578.400 ;
        RECT 61.800 579.300 63.600 584.400 ;
        RECT 67.800 579.300 69.600 584.400 ;
        RECT 61.800 577.950 69.600 579.300 ;
        RECT 80.400 579.300 82.200 584.400 ;
        RECT 86.400 579.300 88.200 584.400 ;
        RECT 80.400 577.950 88.200 579.300 ;
        RECT 89.400 578.400 91.200 584.400 ;
        RECT 110.400 581.400 112.200 584.400 ;
        RECT 89.400 576.300 90.600 578.400 ;
        RECT 59.400 575.250 63.150 576.300 ;
        RECT 41.100 571.050 42.900 572.850 ;
        RECT 59.100 571.050 60.900 572.850 ;
        RECT 61.950 571.050 63.150 575.250 ;
        RECT 86.850 575.250 90.600 576.300 ;
        RECT 65.100 571.050 66.900 572.850 ;
        RECT 83.100 571.050 84.900 572.850 ;
        RECT 86.850 571.050 88.050 575.250 ;
        RECT 89.100 571.050 90.900 572.850 ;
        RECT 110.400 571.050 111.600 581.400 ;
        RECT 130.800 577.200 132.600 584.400 ;
        RECT 146.400 579.300 148.200 584.400 ;
        RECT 152.400 579.300 154.200 584.400 ;
        RECT 146.400 577.950 154.200 579.300 ;
        RECT 155.400 578.400 157.200 584.400 ;
        RECT 172.800 581.400 174.600 584.400 ;
        RECT 128.400 576.300 132.600 577.200 ;
        RECT 155.400 576.300 156.600 578.400 ;
        RECT 125.100 571.050 126.900 572.850 ;
        RECT 128.400 571.050 129.600 576.300 ;
        RECT 152.850 575.250 156.600 576.300 ;
        RECT 131.100 571.050 132.900 572.850 ;
        RECT 149.100 571.050 150.900 572.850 ;
        RECT 152.850 571.050 154.050 575.250 ;
        RECT 155.100 571.050 156.900 572.850 ;
        RECT 173.400 571.050 174.600 581.400 ;
        RECT 193.800 577.200 195.600 584.400 ;
        RECT 191.400 576.300 195.600 577.200 ;
        RECT 200.550 578.400 202.350 584.400 ;
        RECT 208.650 581.400 210.450 584.400 ;
        RECT 216.450 581.400 218.250 584.400 ;
        RECT 224.250 582.300 226.050 584.400 ;
        RECT 224.250 581.400 228.000 582.300 ;
        RECT 208.650 580.500 209.700 581.400 ;
        RECT 205.950 579.300 209.700 580.500 ;
        RECT 217.200 580.500 218.250 581.400 ;
        RECT 226.950 580.500 228.000 581.400 ;
        RECT 217.200 579.450 222.150 580.500 ;
        RECT 205.950 578.400 208.050 579.300 ;
        RECT 220.350 578.700 222.150 579.450 ;
        RECT 188.100 571.050 189.900 572.850 ;
        RECT 191.400 571.050 192.600 576.300 ;
        RECT 194.100 571.050 195.900 572.850 ;
        RECT 200.550 571.050 201.750 578.400 ;
        RECT 223.650 577.800 225.450 579.600 ;
        RECT 226.950 578.400 229.050 580.500 ;
        RECT 232.050 578.400 233.850 584.400 ;
        RECT 213.150 576.000 214.950 576.600 ;
        RECT 224.100 576.000 225.150 577.800 ;
        RECT 213.150 574.800 225.150 576.000 ;
        RECT 13.950 568.950 16.050 571.050 ;
        RECT 16.950 568.950 19.050 571.050 ;
        RECT 19.950 568.950 22.050 571.050 ;
        RECT 34.950 568.950 37.050 571.050 ;
        RECT 37.950 568.950 40.050 571.050 ;
        RECT 40.950 568.950 43.050 571.050 ;
        RECT 58.950 568.950 61.050 571.050 ;
        RECT 61.950 568.950 64.050 571.050 ;
        RECT 64.950 568.950 67.050 571.050 ;
        RECT 67.950 568.950 70.050 571.050 ;
        RECT 79.950 568.950 82.050 571.050 ;
        RECT 82.950 568.950 85.050 571.050 ;
        RECT 85.950 568.950 88.050 571.050 ;
        RECT 88.950 568.950 91.050 571.050 ;
        RECT 106.950 568.950 109.050 571.050 ;
        RECT 109.950 568.950 112.050 571.050 ;
        RECT 124.950 568.950 127.050 571.050 ;
        RECT 127.950 568.950 130.050 571.050 ;
        RECT 130.950 568.950 133.050 571.050 ;
        RECT 145.950 568.950 148.050 571.050 ;
        RECT 148.950 568.950 151.050 571.050 ;
        RECT 151.950 568.950 154.050 571.050 ;
        RECT 154.950 568.950 157.050 571.050 ;
        RECT 172.950 568.950 175.050 571.050 ;
        RECT 175.950 568.950 178.050 571.050 ;
        RECT 187.950 568.950 190.050 571.050 ;
        RECT 190.950 568.950 193.050 571.050 ;
        RECT 193.950 568.950 196.050 571.050 ;
        RECT 200.550 569.250 206.850 571.050 ;
        RECT 200.550 568.950 205.050 569.250 ;
        RECT 14.100 567.150 15.900 568.950 ;
        RECT 17.400 561.600 18.300 568.950 ;
        RECT 20.100 567.150 21.900 568.950 ;
        RECT 14.700 560.400 18.300 561.600 ;
        RECT 14.700 549.600 16.500 560.400 ;
        RECT 38.400 555.600 39.600 568.950 ;
        RECT 46.950 564.450 49.050 565.050 ;
        RECT 58.950 564.450 61.050 565.050 ;
        RECT 46.950 563.550 61.050 564.450 ;
        RECT 46.950 562.950 49.050 563.550 ;
        RECT 58.950 562.950 61.050 563.550 ;
        RECT 62.850 555.600 64.050 568.950 ;
        RECT 68.100 567.150 69.900 568.950 ;
        RECT 80.100 567.150 81.900 568.950 ;
        RECT 85.950 555.600 87.150 568.950 ;
        RECT 107.100 567.150 108.900 568.950 ;
        RECT 110.400 555.600 111.600 568.950 ;
        RECT 128.400 555.600 129.600 568.950 ;
        RECT 146.100 567.150 147.900 568.950 ;
        RECT 151.950 555.600 153.150 568.950 ;
        RECT 154.950 564.450 157.050 565.050 ;
        RECT 166.950 564.450 169.050 565.050 ;
        RECT 154.950 563.550 169.050 564.450 ;
        RECT 154.950 562.950 157.050 563.550 ;
        RECT 166.950 562.950 169.050 563.550 ;
        RECT 173.400 555.600 174.600 568.950 ;
        RECT 176.100 567.150 177.900 568.950 ;
        RECT 181.950 564.450 184.050 565.050 ;
        RECT 187.950 564.450 190.050 565.050 ;
        RECT 181.950 563.550 190.050 564.450 ;
        RECT 181.950 562.950 184.050 563.550 ;
        RECT 187.950 562.950 190.050 563.550 ;
        RECT 37.800 549.600 39.600 555.600 ;
        RECT 43.950 552.450 46.050 553.050 ;
        RECT 52.950 552.450 55.050 553.050 ;
        RECT 43.950 551.550 55.050 552.450 ;
        RECT 43.950 550.950 46.050 551.550 ;
        RECT 52.950 550.950 55.050 551.550 ;
        RECT 62.400 549.600 64.200 555.600 ;
        RECT 85.800 549.600 87.600 555.600 ;
        RECT 110.400 549.600 112.200 555.600 ;
        RECT 128.400 549.600 130.200 555.600 ;
        RECT 151.800 549.600 153.600 555.600 ;
        RECT 172.800 549.600 174.600 555.600 ;
        RECT 191.400 555.600 192.600 568.950 ;
        RECT 200.550 561.600 201.750 568.950 ;
        RECT 202.950 563.400 204.750 565.200 ;
        RECT 203.850 562.200 208.050 563.400 ;
        RECT 213.150 562.200 214.050 574.800 ;
        RECT 224.100 573.600 231.000 574.800 ;
        RECT 224.100 573.000 225.900 573.600 ;
        RECT 230.100 572.850 231.000 573.600 ;
        RECT 227.100 571.800 228.900 572.400 ;
        RECT 220.950 570.600 228.900 571.800 ;
        RECT 230.100 571.050 231.900 572.850 ;
        RECT 220.950 568.950 223.050 570.600 ;
        RECT 229.950 568.950 232.050 571.050 ;
        RECT 222.750 563.700 224.550 564.000 ;
        RECT 232.950 563.700 233.850 578.400 ;
        RECT 250.800 577.200 252.600 584.400 ;
        RECT 271.800 577.200 273.600 584.400 ;
        RECT 248.400 576.300 252.600 577.200 ;
        RECT 269.400 576.300 273.600 577.200 ;
        RECT 290.400 577.500 292.200 584.400 ;
        RECT 296.400 577.500 298.200 584.400 ;
        RECT 302.400 577.500 304.200 584.400 ;
        RECT 308.400 577.500 310.200 584.400 ;
        RECT 290.400 576.300 294.300 577.500 ;
        RECT 296.400 576.300 300.300 577.500 ;
        RECT 302.400 576.300 306.300 577.500 ;
        RECT 308.400 576.300 311.100 577.500 ;
        RECT 245.100 571.050 246.900 572.850 ;
        RECT 248.400 571.050 249.600 576.300 ;
        RECT 251.100 571.050 252.900 572.850 ;
        RECT 266.100 571.050 267.900 572.850 ;
        RECT 269.400 571.050 270.600 576.300 ;
        RECT 293.100 575.400 294.300 576.300 ;
        RECT 299.100 575.400 300.300 576.300 ;
        RECT 305.100 575.400 306.300 576.300 ;
        RECT 293.100 574.200 297.300 575.400 ;
        RECT 272.100 571.050 273.900 572.850 ;
        RECT 290.100 571.050 291.900 572.850 ;
        RECT 244.950 568.950 247.050 571.050 ;
        RECT 247.950 568.950 250.050 571.050 ;
        RECT 250.950 568.950 253.050 571.050 ;
        RECT 265.950 568.950 268.050 571.050 ;
        RECT 268.950 568.950 271.050 571.050 ;
        RECT 271.950 568.950 274.050 571.050 ;
        RECT 289.950 568.950 292.050 571.050 ;
        RECT 222.750 563.100 233.850 563.700 ;
        RECT 191.400 549.600 193.200 555.600 ;
        RECT 200.550 549.600 202.350 561.600 ;
        RECT 205.950 561.300 208.050 562.200 ;
        RECT 208.950 561.300 214.050 562.200 ;
        RECT 216.150 562.500 233.850 563.100 ;
        RECT 216.150 562.200 224.550 562.500 ;
        RECT 208.950 560.400 209.850 561.300 ;
        RECT 207.150 558.600 209.850 560.400 ;
        RECT 210.750 560.100 212.550 560.400 ;
        RECT 216.150 560.100 217.050 562.200 ;
        RECT 232.950 561.600 233.850 562.500 ;
        RECT 210.750 559.200 217.050 560.100 ;
        RECT 217.950 560.700 219.750 561.300 ;
        RECT 217.950 559.500 225.450 560.700 ;
        RECT 210.750 558.600 212.550 559.200 ;
        RECT 224.250 558.600 225.450 559.500 ;
        RECT 205.950 555.600 209.850 557.700 ;
        RECT 214.950 557.550 216.750 558.300 ;
        RECT 219.750 557.550 221.550 558.300 ;
        RECT 214.950 556.500 221.550 557.550 ;
        RECT 224.250 556.500 229.050 558.600 ;
        RECT 208.050 549.600 209.850 555.600 ;
        RECT 215.850 549.600 217.650 556.500 ;
        RECT 224.250 555.600 225.450 556.500 ;
        RECT 223.650 549.600 225.450 555.600 ;
        RECT 232.050 549.600 233.850 561.600 ;
        RECT 248.400 555.600 249.600 568.950 ;
        RECT 269.400 555.600 270.600 568.950 ;
        RECT 293.100 563.700 294.300 574.200 ;
        RECT 295.500 573.600 297.300 574.200 ;
        RECT 299.100 574.200 303.300 575.400 ;
        RECT 299.100 563.700 300.300 574.200 ;
        RECT 301.500 573.600 303.300 574.200 ;
        RECT 305.100 574.200 309.300 575.400 ;
        RECT 305.100 563.700 306.300 574.200 ;
        RECT 307.500 573.600 309.300 574.200 ;
        RECT 310.200 571.050 311.100 576.300 ;
        RECT 333.000 576.000 334.800 584.400 ;
        RECT 353.400 577.500 355.200 584.400 ;
        RECT 359.400 577.500 361.200 584.400 ;
        RECT 365.400 577.500 367.200 584.400 ;
        RECT 371.400 577.500 373.200 584.400 ;
        RECT 391.800 581.400 393.600 584.400 ;
        RECT 353.400 576.300 357.300 577.500 ;
        RECT 359.400 576.300 363.300 577.500 ;
        RECT 365.400 576.300 369.300 577.500 ;
        RECT 371.400 576.300 374.100 577.500 ;
        RECT 333.000 574.800 336.300 576.000 ;
        RECT 326.100 571.050 327.900 572.850 ;
        RECT 332.100 571.050 333.900 572.850 ;
        RECT 335.400 571.050 336.300 574.800 ;
        RECT 356.100 575.400 357.300 576.300 ;
        RECT 362.100 575.400 363.300 576.300 ;
        RECT 368.100 575.400 369.300 576.300 ;
        RECT 356.100 574.200 360.300 575.400 ;
        RECT 353.100 571.050 354.900 572.850 ;
        RECT 310.200 568.950 313.050 571.050 ;
        RECT 325.950 568.950 328.050 571.050 ;
        RECT 328.950 568.950 331.050 571.050 ;
        RECT 331.950 568.950 334.050 571.050 ;
        RECT 334.950 568.950 337.050 571.050 ;
        RECT 352.950 568.950 355.050 571.050 ;
        RECT 310.200 563.700 311.100 568.950 ;
        RECT 329.100 567.150 330.900 568.950 ;
        RECT 290.400 562.500 294.300 563.700 ;
        RECT 296.400 562.500 300.300 563.700 ;
        RECT 302.400 562.500 306.300 563.700 ;
        RECT 308.400 562.500 311.100 563.700 ;
        RECT 248.400 549.600 250.200 555.600 ;
        RECT 269.400 549.600 271.200 555.600 ;
        RECT 290.400 549.600 292.200 562.500 ;
        RECT 296.400 549.600 298.200 562.500 ;
        RECT 302.400 549.600 304.200 562.500 ;
        RECT 308.400 549.600 310.200 562.500 ;
        RECT 335.400 556.800 336.300 568.950 ;
        RECT 356.100 563.700 357.300 574.200 ;
        RECT 358.500 573.600 360.300 574.200 ;
        RECT 362.100 574.200 366.300 575.400 ;
        RECT 362.100 563.700 363.300 574.200 ;
        RECT 364.500 573.600 366.300 574.200 ;
        RECT 368.100 574.200 372.300 575.400 ;
        RECT 368.100 563.700 369.300 574.200 ;
        RECT 370.500 573.600 372.300 574.200 ;
        RECT 373.200 571.050 374.100 576.300 ;
        RECT 392.400 571.050 393.600 581.400 ;
        RECT 409.800 578.400 411.600 584.400 ;
        RECT 415.800 581.400 417.600 584.400 ;
        RECT 430.800 581.400 432.600 584.400 ;
        RECT 409.800 571.050 411.000 578.400 ;
        RECT 416.400 577.500 417.600 581.400 ;
        RECT 411.900 576.600 417.600 577.500 ;
        RECT 411.900 575.700 413.850 576.600 ;
        RECT 373.200 568.950 376.050 571.050 ;
        RECT 391.950 568.950 394.050 571.050 ;
        RECT 394.950 568.950 397.050 571.050 ;
        RECT 409.800 568.950 412.050 571.050 ;
        RECT 373.200 563.700 374.100 568.950 ;
        RECT 329.700 555.900 336.300 556.800 ;
        RECT 329.700 555.600 331.200 555.900 ;
        RECT 329.400 549.600 331.200 555.600 ;
        RECT 335.400 555.600 336.300 555.900 ;
        RECT 353.400 562.500 357.300 563.700 ;
        RECT 359.400 562.500 363.300 563.700 ;
        RECT 365.400 562.500 369.300 563.700 ;
        RECT 371.400 562.500 374.100 563.700 ;
        RECT 335.400 549.600 337.200 555.600 ;
        RECT 353.400 549.600 355.200 562.500 ;
        RECT 359.400 549.600 361.200 562.500 ;
        RECT 365.400 549.600 367.200 562.500 ;
        RECT 371.400 549.600 373.200 562.500 ;
        RECT 392.400 555.600 393.600 568.950 ;
        RECT 395.100 567.150 396.900 568.950 ;
        RECT 391.800 549.600 393.600 555.600 ;
        RECT 409.800 561.600 411.000 568.950 ;
        RECT 412.950 564.300 413.850 575.700 ;
        RECT 431.400 571.050 432.600 581.400 ;
        RECT 451.800 577.200 453.600 584.400 ;
        RECT 449.400 576.300 453.600 577.200 ;
        RECT 470.400 577.200 472.200 584.400 ;
        RECT 491.400 577.200 493.200 584.400 ;
        RECT 514.800 577.200 516.600 584.400 ;
        RECT 532.800 578.400 534.600 584.400 ;
        RECT 470.400 576.300 474.600 577.200 ;
        RECT 491.400 576.300 495.600 577.200 ;
        RECT 446.100 571.050 447.900 572.850 ;
        RECT 449.400 571.050 450.600 576.300 ;
        RECT 452.100 571.050 453.900 572.850 ;
        RECT 470.100 571.050 471.900 572.850 ;
        RECT 473.400 571.050 474.600 576.300 ;
        RECT 476.100 571.050 477.900 572.850 ;
        RECT 491.100 571.050 492.900 572.850 ;
        RECT 494.400 571.050 495.600 576.300 ;
        RECT 512.400 576.300 516.600 577.200 ;
        RECT 533.400 576.300 534.600 578.400 ;
        RECT 535.800 579.300 537.600 584.400 ;
        RECT 541.800 579.300 543.600 584.400 ;
        RECT 535.800 577.950 543.600 579.300 ;
        RECT 546.150 578.400 547.950 584.400 ;
        RECT 553.950 582.300 555.750 584.400 ;
        RECT 552.000 581.400 555.750 582.300 ;
        RECT 561.750 581.400 563.550 584.400 ;
        RECT 569.550 581.400 571.350 584.400 ;
        RECT 552.000 580.500 553.050 581.400 ;
        RECT 561.750 580.500 562.800 581.400 ;
        RECT 550.950 578.400 553.050 580.500 ;
        RECT 497.100 571.050 498.900 572.850 ;
        RECT 509.100 571.050 510.900 572.850 ;
        RECT 512.400 571.050 513.600 576.300 ;
        RECT 533.400 575.250 537.150 576.300 ;
        RECT 515.100 571.050 516.900 572.850 ;
        RECT 533.100 571.050 534.900 572.850 ;
        RECT 535.950 571.050 537.150 575.250 ;
        RECT 539.100 571.050 540.900 572.850 ;
        RECT 415.950 568.950 418.050 571.050 ;
        RECT 430.950 568.950 433.050 571.050 ;
        RECT 433.950 568.950 436.050 571.050 ;
        RECT 445.950 568.950 448.050 571.050 ;
        RECT 448.950 568.950 451.050 571.050 ;
        RECT 451.950 568.950 454.050 571.050 ;
        RECT 469.950 568.950 472.050 571.050 ;
        RECT 472.950 568.950 475.050 571.050 ;
        RECT 475.950 568.950 478.050 571.050 ;
        RECT 490.950 568.950 493.050 571.050 ;
        RECT 493.950 568.950 496.050 571.050 ;
        RECT 496.950 568.950 499.050 571.050 ;
        RECT 508.950 568.950 511.050 571.050 ;
        RECT 511.950 568.950 514.050 571.050 ;
        RECT 514.950 568.950 517.050 571.050 ;
        RECT 532.950 568.950 535.050 571.050 ;
        RECT 535.950 568.950 538.050 571.050 ;
        RECT 538.950 568.950 541.050 571.050 ;
        RECT 541.950 568.950 544.050 571.050 ;
        RECT 416.100 567.150 417.900 568.950 ;
        RECT 411.900 563.400 413.850 564.300 ;
        RECT 411.900 562.500 417.600 563.400 ;
        RECT 409.800 549.600 411.600 561.600 ;
        RECT 416.400 555.600 417.600 562.500 ;
        RECT 431.400 555.600 432.600 568.950 ;
        RECT 434.100 567.150 435.900 568.950 ;
        RECT 415.800 549.600 417.600 555.600 ;
        RECT 430.800 549.600 432.600 555.600 ;
        RECT 449.400 555.600 450.600 568.950 ;
        RECT 473.400 555.600 474.600 568.950 ;
        RECT 494.400 555.600 495.600 568.950 ;
        RECT 449.400 549.600 451.200 555.600 ;
        RECT 472.800 549.600 474.600 555.600 ;
        RECT 493.800 549.600 495.600 555.600 ;
        RECT 512.400 555.600 513.600 568.950 ;
        RECT 536.850 555.600 538.050 568.950 ;
        RECT 542.100 567.150 543.900 568.950 ;
        RECT 546.150 563.700 547.050 578.400 ;
        RECT 554.550 577.800 556.350 579.600 ;
        RECT 557.850 579.450 562.800 580.500 ;
        RECT 570.300 580.500 571.350 581.400 ;
        RECT 557.850 578.700 559.650 579.450 ;
        RECT 570.300 579.300 574.050 580.500 ;
        RECT 571.950 578.400 574.050 579.300 ;
        RECT 577.650 578.400 579.450 584.400 ;
        RECT 554.850 576.000 555.900 577.800 ;
        RECT 565.050 576.000 566.850 576.600 ;
        RECT 554.850 574.800 566.850 576.000 ;
        RECT 549.000 573.600 555.900 574.800 ;
        RECT 549.000 572.850 549.900 573.600 ;
        RECT 554.100 573.000 555.900 573.600 ;
        RECT 548.100 571.050 549.900 572.850 ;
        RECT 551.100 571.800 552.900 572.400 ;
        RECT 547.950 568.950 550.050 571.050 ;
        RECT 551.100 570.600 559.050 571.800 ;
        RECT 556.950 568.950 559.050 570.600 ;
        RECT 555.450 563.700 557.250 564.000 ;
        RECT 546.150 563.100 557.250 563.700 ;
        RECT 546.150 562.500 563.850 563.100 ;
        RECT 546.150 561.600 547.050 562.500 ;
        RECT 555.450 562.200 563.850 562.500 ;
        RECT 512.400 549.600 514.200 555.600 ;
        RECT 536.400 549.600 538.200 555.600 ;
        RECT 546.150 549.600 547.950 561.600 ;
        RECT 560.250 560.700 562.050 561.300 ;
        RECT 554.550 559.500 562.050 560.700 ;
        RECT 562.950 560.100 563.850 562.200 ;
        RECT 565.950 562.200 566.850 574.800 ;
        RECT 578.250 571.050 579.450 578.400 ;
        RECT 593.400 581.400 595.200 584.400 ;
        RECT 593.400 571.050 594.600 581.400 ;
        RECT 611.400 578.400 613.200 584.400 ;
        RECT 608.100 571.050 609.900 572.850 ;
        RECT 611.400 571.050 612.600 578.400 ;
        RECT 629.400 577.200 631.200 584.400 ;
        RECT 647.400 581.400 649.200 584.400 ;
        RECT 647.400 577.500 648.600 581.400 ;
        RECT 653.400 578.400 655.200 584.400 ;
        RECT 672.300 580.200 674.100 584.400 ;
        RECT 629.400 576.300 633.600 577.200 ;
        RECT 647.400 576.600 653.100 577.500 ;
        RECT 629.100 571.050 630.900 572.850 ;
        RECT 632.400 571.050 633.600 576.300 ;
        RECT 651.150 575.700 653.100 576.600 ;
        RECT 635.100 571.050 636.900 572.850 ;
        RECT 573.150 569.250 579.450 571.050 ;
        RECT 574.950 568.950 579.450 569.250 ;
        RECT 589.950 568.950 592.050 571.050 ;
        RECT 592.950 568.950 595.050 571.050 ;
        RECT 607.950 568.950 610.050 571.050 ;
        RECT 610.950 568.950 613.050 571.050 ;
        RECT 628.950 568.950 631.050 571.050 ;
        RECT 631.950 568.950 634.050 571.050 ;
        RECT 634.950 568.950 637.050 571.050 ;
        RECT 646.950 568.950 649.050 571.050 ;
        RECT 575.250 563.400 577.050 565.200 ;
        RECT 571.950 562.200 576.150 563.400 ;
        RECT 565.950 561.300 571.050 562.200 ;
        RECT 571.950 561.300 574.050 562.200 ;
        RECT 578.250 561.600 579.450 568.950 ;
        RECT 590.100 567.150 591.900 568.950 ;
        RECT 570.150 560.400 571.050 561.300 ;
        RECT 567.450 560.100 569.250 560.400 ;
        RECT 554.550 558.600 555.750 559.500 ;
        RECT 562.950 559.200 569.250 560.100 ;
        RECT 567.450 558.600 569.250 559.200 ;
        RECT 570.150 558.600 572.850 560.400 ;
        RECT 550.950 556.500 555.750 558.600 ;
        RECT 558.450 557.550 560.250 558.300 ;
        RECT 563.250 557.550 565.050 558.300 ;
        RECT 558.450 556.500 565.050 557.550 ;
        RECT 554.550 555.600 555.750 556.500 ;
        RECT 554.550 549.600 556.350 555.600 ;
        RECT 562.350 549.600 564.150 556.500 ;
        RECT 570.150 555.600 574.050 557.700 ;
        RECT 570.150 549.600 571.950 555.600 ;
        RECT 577.650 549.600 579.450 561.600 ;
        RECT 593.400 555.600 594.600 568.950 ;
        RECT 611.400 561.600 612.600 568.950 ;
        RECT 593.400 549.600 595.200 555.600 ;
        RECT 611.400 549.600 613.200 561.600 ;
        RECT 632.400 555.600 633.600 568.950 ;
        RECT 647.100 567.150 648.900 568.950 ;
        RECT 651.150 564.300 652.050 575.700 ;
        RECT 654.000 571.050 655.200 578.400 ;
        RECT 671.400 578.400 674.100 580.200 ;
        RECT 666.000 573.450 670.050 574.050 ;
        RECT 652.950 568.950 655.200 571.050 ;
        RECT 651.150 563.400 653.100 564.300 ;
        RECT 631.800 549.600 633.600 555.600 ;
        RECT 647.400 562.500 653.100 563.400 ;
        RECT 647.400 555.600 648.600 562.500 ;
        RECT 654.000 561.600 655.200 568.950 ;
        RECT 665.550 571.950 670.050 573.450 ;
        RECT 665.550 568.050 666.450 571.950 ;
        RECT 671.400 571.050 672.300 578.400 ;
        RECT 674.100 576.600 675.900 577.500 ;
        RECT 679.800 576.600 681.600 584.400 ;
        RECT 674.100 575.700 681.600 576.600 ;
        RECT 695.400 577.200 697.200 584.400 ;
        RECT 713.400 579.300 715.200 584.400 ;
        RECT 719.400 579.300 721.200 584.400 ;
        RECT 713.400 577.950 721.200 579.300 ;
        RECT 722.400 578.400 724.200 584.400 ;
        RECT 695.400 576.300 699.600 577.200 ;
        RECT 722.400 576.300 723.600 578.400 ;
        RECT 670.950 568.950 673.050 571.050 ;
        RECT 673.950 568.950 676.050 571.050 ;
        RECT 665.550 566.550 670.050 568.050 ;
        RECT 666.000 565.950 670.050 566.550 ;
        RECT 671.400 561.600 672.300 568.950 ;
        RECT 674.100 567.150 675.900 568.950 ;
        RECT 647.400 549.600 649.200 555.600 ;
        RECT 653.400 549.600 655.200 561.600 ;
        RECT 670.800 549.600 672.600 561.600 ;
        RECT 677.700 555.600 678.600 575.700 ;
        RECT 691.950 573.450 694.050 574.050 ;
        RECT 680.100 571.050 681.900 572.850 ;
        RECT 686.550 572.550 694.050 573.450 ;
        RECT 679.950 568.950 682.050 571.050 ;
        RECT 686.550 568.050 687.450 572.550 ;
        RECT 691.950 571.950 694.050 572.550 ;
        RECT 695.100 571.050 696.900 572.850 ;
        RECT 698.400 571.050 699.600 576.300 ;
        RECT 719.850 575.250 723.600 576.300 ;
        RECT 724.950 576.450 727.050 577.050 ;
        RECT 736.950 576.450 739.050 580.050 ;
        RECT 724.950 576.000 739.050 576.450 ;
        RECT 740.400 577.200 742.200 584.400 ;
        RECT 740.400 576.300 744.600 577.200 ;
        RECT 724.950 575.550 738.450 576.000 ;
        RECT 701.100 571.050 702.900 572.850 ;
        RECT 706.950 571.950 709.050 574.050 ;
        RECT 694.950 568.950 697.050 571.050 ;
        RECT 697.950 568.950 700.050 571.050 ;
        RECT 700.950 568.950 703.050 571.050 ;
        RECT 682.950 566.550 687.450 568.050 ;
        RECT 682.950 565.950 687.000 566.550 ;
        RECT 698.400 555.600 699.600 568.950 ;
        RECT 707.550 568.050 708.450 571.950 ;
        RECT 716.100 571.050 717.900 572.850 ;
        RECT 719.850 571.050 721.050 575.250 ;
        RECT 724.950 574.950 727.050 575.550 ;
        RECT 722.100 571.050 723.900 572.850 ;
        RECT 740.100 571.050 741.900 572.850 ;
        RECT 743.400 571.050 744.600 576.300 ;
        RECT 765.000 576.000 766.800 584.400 ;
        RECT 790.200 578.400 792.000 584.400 ;
        RECT 814.800 578.400 816.600 584.400 ;
        RECT 765.000 574.800 768.300 576.000 ;
        RECT 753.000 573.450 757.050 574.050 ;
        RECT 746.100 571.050 747.900 572.850 ;
        RECT 752.550 571.950 757.050 573.450 ;
        RECT 712.950 568.950 715.050 571.050 ;
        RECT 715.950 568.950 718.050 571.050 ;
        RECT 718.950 568.950 721.050 571.050 ;
        RECT 721.950 568.950 724.050 571.050 ;
        RECT 739.950 568.950 742.050 571.050 ;
        RECT 742.950 568.950 745.050 571.050 ;
        RECT 745.950 568.950 748.050 571.050 ;
        RECT 706.950 565.950 709.050 568.050 ;
        RECT 713.100 567.150 714.900 568.950 ;
        RECT 718.950 555.600 720.150 568.950 ;
        RECT 743.400 555.600 744.600 568.950 ;
        RECT 752.550 568.050 753.450 571.950 ;
        RECT 758.100 571.050 759.900 572.850 ;
        RECT 764.100 571.050 765.900 572.850 ;
        RECT 767.400 571.050 768.300 574.800 ;
        RECT 780.000 573.450 784.050 574.050 ;
        RECT 779.550 571.950 784.050 573.450 ;
        RECT 757.950 568.950 760.050 571.050 ;
        RECT 760.950 568.950 763.050 571.050 ;
        RECT 763.950 568.950 766.050 571.050 ;
        RECT 766.950 568.950 769.050 571.050 ;
        RECT 748.950 566.550 753.450 568.050 ;
        RECT 761.100 567.150 762.900 568.950 ;
        RECT 748.950 565.950 753.000 566.550 ;
        RECT 767.400 556.800 768.300 568.950 ;
        RECT 779.550 568.050 780.450 571.950 ;
        RECT 785.100 571.050 786.900 572.850 ;
        RECT 790.950 571.050 792.000 578.400 ;
        RECT 802.950 576.450 807.000 577.050 ;
        RECT 802.950 574.950 807.450 576.450 ;
        RECT 815.400 576.300 816.600 578.400 ;
        RECT 817.800 579.300 819.600 584.400 ;
        RECT 823.800 579.300 825.600 584.400 ;
        RECT 829.950 580.950 832.050 583.050 ;
        RECT 817.800 577.950 825.600 579.300 ;
        RECT 815.400 575.250 819.150 576.300 ;
        RECT 799.950 573.450 804.000 574.050 ;
        RECT 797.100 571.050 798.900 572.850 ;
        RECT 799.950 571.950 804.450 573.450 ;
        RECT 784.950 568.950 787.050 571.050 ;
        RECT 787.950 568.950 790.050 571.050 ;
        RECT 790.950 568.950 793.050 571.050 ;
        RECT 793.950 568.950 796.050 571.050 ;
        RECT 796.950 568.950 799.050 571.050 ;
        RECT 779.550 566.550 784.050 568.050 ;
        RECT 788.100 567.150 789.900 568.950 ;
        RECT 780.000 565.950 784.050 566.550 ;
        RECT 769.950 564.450 772.050 565.050 ;
        RECT 787.950 564.450 790.050 565.050 ;
        RECT 769.950 563.550 790.050 564.450 ;
        RECT 769.950 562.950 772.050 563.550 ;
        RECT 787.950 562.950 790.050 563.550 ;
        RECT 791.100 563.400 792.000 568.950 ;
        RECT 794.100 567.150 795.900 568.950 ;
        RECT 803.550 568.050 804.450 571.950 ;
        RECT 806.550 571.050 807.450 574.950 ;
        RECT 815.100 571.050 816.900 572.850 ;
        RECT 817.950 571.050 819.150 575.250 ;
        RECT 821.100 571.050 822.900 572.850 ;
        RECT 806.550 570.900 810.000 571.050 ;
        RECT 806.550 569.550 811.050 570.900 ;
        RECT 807.000 568.950 811.050 569.550 ;
        RECT 814.950 568.950 817.050 571.050 ;
        RECT 817.950 568.950 820.050 571.050 ;
        RECT 820.950 568.950 823.050 571.050 ;
        RECT 823.950 568.950 826.050 571.050 ;
        RECT 808.950 568.800 811.050 568.950 ;
        RECT 799.950 566.550 804.450 568.050 ;
        RECT 799.950 565.950 804.000 566.550 ;
        RECT 791.100 562.500 796.200 563.400 ;
        RECT 761.700 555.900 768.300 556.800 ;
        RECT 761.700 555.600 763.200 555.900 ;
        RECT 676.800 549.600 678.600 555.600 ;
        RECT 697.800 549.600 699.600 555.600 ;
        RECT 718.800 549.600 720.600 555.600 ;
        RECT 742.800 549.600 744.600 555.600 ;
        RECT 761.400 549.600 763.200 555.600 ;
        RECT 767.400 555.600 768.300 555.900 ;
        RECT 785.400 560.400 793.200 561.300 ;
        RECT 767.400 549.600 769.200 555.600 ;
        RECT 785.400 549.600 787.200 560.400 ;
        RECT 791.400 550.500 793.200 560.400 ;
        RECT 794.400 551.400 796.200 562.500 ;
        RECT 797.400 550.500 799.200 561.600 ;
        RECT 818.850 555.600 820.050 568.950 ;
        RECT 824.100 567.150 825.900 568.950 ;
        RECT 830.550 567.450 831.450 580.950 ;
        RECT 836.400 579.300 838.200 584.400 ;
        RECT 842.400 579.300 844.200 584.400 ;
        RECT 836.400 577.950 844.200 579.300 ;
        RECT 845.400 578.400 847.200 584.400 ;
        RECT 845.400 576.300 846.600 578.400 ;
        RECT 842.850 575.250 846.600 576.300 ;
        RECT 867.000 576.000 868.800 584.400 ;
        RECT 839.100 571.050 840.900 572.850 ;
        RECT 842.850 571.050 844.050 575.250 ;
        RECT 867.000 574.800 870.300 576.000 ;
        RECT 845.100 571.050 846.900 572.850 ;
        RECT 860.100 571.050 861.900 572.850 ;
        RECT 866.100 571.050 867.900 572.850 ;
        RECT 869.400 571.050 870.300 574.800 ;
        RECT 835.950 568.950 838.050 571.050 ;
        RECT 838.950 568.950 841.050 571.050 ;
        RECT 841.950 568.950 844.050 571.050 ;
        RECT 844.950 568.950 847.050 571.050 ;
        RECT 859.950 568.950 862.050 571.050 ;
        RECT 862.950 568.950 865.050 571.050 ;
        RECT 865.950 568.950 868.050 571.050 ;
        RECT 868.950 568.950 871.050 571.050 ;
        RECT 830.550 566.550 834.450 567.450 ;
        RECT 836.100 567.150 837.900 568.950 ;
        RECT 833.550 565.050 834.450 566.550 ;
        RECT 833.550 563.550 838.050 565.050 ;
        RECT 834.000 562.950 838.050 563.550 ;
        RECT 841.950 555.600 843.150 568.950 ;
        RECT 863.100 567.150 864.900 568.950 ;
        RECT 869.400 556.800 870.300 568.950 ;
        RECT 863.700 555.900 870.300 556.800 ;
        RECT 863.700 555.600 865.200 555.900 ;
        RECT 791.400 549.600 799.200 550.500 ;
        RECT 818.400 549.600 820.200 555.600 ;
        RECT 841.800 549.600 843.600 555.600 ;
        RECT 863.400 549.600 865.200 555.600 ;
        RECT 869.400 555.600 870.300 555.900 ;
        RECT 869.400 549.600 871.200 555.600 ;
        RECT 16.800 539.400 18.600 545.400 ;
        RECT 40.800 539.400 42.600 545.400 ;
        RECT 11.100 526.050 12.900 527.850 ;
        RECT 16.950 526.050 18.150 539.400 ;
        RECT 41.400 526.050 42.600 539.400 ;
        RECT 58.800 534.600 60.600 545.400 ;
        RECT 58.800 533.400 63.600 534.600 ;
        RECT 61.500 532.500 63.600 533.400 ;
        RECT 66.300 533.400 68.100 545.400 ;
        RECT 73.800 534.300 75.600 545.400 ;
        RECT 71.100 533.400 75.600 534.300 ;
        RECT 77.550 533.400 79.350 545.400 ;
        RECT 85.050 539.400 86.850 545.400 ;
        RECT 82.950 537.300 86.850 539.400 ;
        RECT 92.850 538.500 94.650 545.400 ;
        RECT 100.650 539.400 102.450 545.400 ;
        RECT 101.250 538.500 102.450 539.400 ;
        RECT 91.950 537.450 98.550 538.500 ;
        RECT 91.950 536.700 93.750 537.450 ;
        RECT 96.750 536.700 98.550 537.450 ;
        RECT 101.250 536.400 106.050 538.500 ;
        RECT 84.150 534.600 86.850 536.400 ;
        RECT 87.750 535.800 89.550 536.400 ;
        RECT 87.750 534.900 94.050 535.800 ;
        RECT 101.250 535.500 102.450 536.400 ;
        RECT 87.750 534.600 89.550 534.900 ;
        RECT 85.950 533.700 86.850 534.600 ;
        RECT 66.300 531.900 67.500 533.400 ;
        RECT 66.000 531.000 67.500 531.900 ;
        RECT 71.100 531.300 73.200 533.400 ;
        RECT 66.000 528.900 66.900 531.000 ;
        RECT 59.100 526.050 60.900 527.850 ;
        RECT 64.800 526.800 66.900 528.900 ;
        RECT 67.800 529.500 69.900 529.800 ;
        RECT 67.800 527.700 71.700 529.500 ;
        RECT 10.950 523.950 13.050 526.050 ;
        RECT 13.950 523.950 16.050 526.050 ;
        RECT 16.950 523.950 19.050 526.050 ;
        RECT 19.950 523.950 22.050 526.050 ;
        RECT 37.950 523.950 40.050 526.050 ;
        RECT 40.950 523.950 43.050 526.050 ;
        RECT 43.950 523.950 46.050 526.050 ;
        RECT 52.950 525.450 57.000 526.050 ;
        RECT 58.950 525.450 61.050 526.050 ;
        RECT 65.400 525.900 67.800 526.800 ;
        RECT 52.950 524.550 61.050 525.450 ;
        RECT 52.950 523.950 57.000 524.550 ;
        RECT 58.950 523.950 61.050 524.550 ;
        RECT 14.100 522.150 15.900 523.950 ;
        RECT 17.850 519.750 19.050 523.950 ;
        RECT 20.100 522.150 21.900 523.950 ;
        RECT 38.100 522.150 39.900 523.950 ;
        RECT 17.850 518.700 21.600 519.750 ;
        RECT 41.400 518.700 42.600 523.950 ;
        RECT 44.100 522.150 45.900 523.950 ;
        RECT 63.600 523.200 65.400 525.000 ;
        RECT 63.750 521.100 65.850 523.200 ;
        RECT 66.750 520.200 67.800 525.900 ;
        RECT 68.700 525.900 70.500 526.500 ;
        RECT 77.550 526.050 78.750 533.400 ;
        RECT 82.950 532.800 85.050 533.700 ;
        RECT 85.950 532.800 91.050 533.700 ;
        RECT 80.850 531.600 85.050 532.800 ;
        RECT 79.950 529.800 81.750 531.600 ;
        RECT 73.500 525.900 75.600 526.050 ;
        RECT 68.700 524.700 75.600 525.900 ;
        RECT 73.500 523.950 75.600 524.700 ;
        RECT 11.400 515.700 19.200 517.050 ;
        RECT 11.400 510.600 13.200 515.700 ;
        RECT 17.400 510.600 19.200 515.700 ;
        RECT 20.400 516.600 21.600 518.700 ;
        RECT 38.400 517.800 42.600 518.700 ;
        RECT 20.400 510.600 22.200 516.600 ;
        RECT 38.400 510.600 40.200 517.800 ;
        RECT 61.500 517.500 63.600 518.700 ;
        RECT 64.800 518.100 67.800 520.200 ;
        RECT 68.700 521.400 70.500 523.200 ;
        RECT 73.800 522.150 75.600 523.950 ;
        RECT 77.550 525.750 82.050 526.050 ;
        RECT 77.550 523.950 83.850 525.750 ;
        RECT 68.700 519.300 70.800 521.400 ;
        RECT 68.700 518.400 75.000 519.300 ;
        RECT 58.800 516.600 63.600 517.500 ;
        RECT 66.600 516.600 67.800 518.100 ;
        RECT 73.800 516.600 75.000 518.400 ;
        RECT 77.550 516.600 78.750 523.950 ;
        RECT 90.150 520.200 91.050 532.800 ;
        RECT 93.150 532.800 94.050 534.900 ;
        RECT 94.950 534.300 102.450 535.500 ;
        RECT 94.950 533.700 96.750 534.300 ;
        RECT 109.050 533.400 110.850 545.400 ;
        RECT 127.800 539.400 129.600 545.400 ;
        RECT 149.400 539.400 151.200 545.400 ;
        RECT 93.150 532.500 101.550 532.800 ;
        RECT 109.950 532.500 110.850 533.400 ;
        RECT 93.150 531.900 110.850 532.500 ;
        RECT 99.750 531.300 110.850 531.900 ;
        RECT 99.750 531.000 101.550 531.300 ;
        RECT 97.950 524.400 100.050 526.050 ;
        RECT 97.950 523.200 105.900 524.400 ;
        RECT 106.950 523.950 109.050 526.050 ;
        RECT 104.100 522.600 105.900 523.200 ;
        RECT 107.100 522.150 108.900 523.950 ;
        RECT 101.100 521.400 102.900 522.000 ;
        RECT 107.100 521.400 108.000 522.150 ;
        RECT 101.100 520.200 108.000 521.400 ;
        RECT 90.150 519.000 102.150 520.200 ;
        RECT 90.150 518.400 91.950 519.000 ;
        RECT 101.100 517.200 102.150 519.000 ;
        RECT 58.800 510.600 60.600 516.600 ;
        RECT 66.300 510.600 68.100 516.600 ;
        RECT 73.800 510.600 75.600 516.600 ;
        RECT 77.550 510.600 79.350 516.600 ;
        RECT 82.950 515.700 85.050 516.600 ;
        RECT 82.950 514.500 86.700 515.700 ;
        RECT 97.350 515.550 99.150 516.300 ;
        RECT 85.650 513.600 86.700 514.500 ;
        RECT 94.200 514.500 99.150 515.550 ;
        RECT 100.650 515.400 102.450 517.200 ;
        RECT 109.950 516.600 110.850 531.300 ;
        RECT 122.100 526.050 123.900 527.850 ;
        RECT 127.950 526.050 129.150 539.400 ;
        RECT 130.950 531.450 133.050 532.050 ;
        RECT 136.950 531.450 139.050 532.050 ;
        RECT 130.950 530.550 139.050 531.450 ;
        RECT 130.950 529.950 133.050 530.550 ;
        RECT 136.950 529.950 139.050 530.550 ;
        RECT 149.400 526.050 150.600 539.400 ;
        RECT 158.550 533.400 160.350 545.400 ;
        RECT 166.050 539.400 167.850 545.400 ;
        RECT 163.950 537.300 167.850 539.400 ;
        RECT 173.850 538.500 175.650 545.400 ;
        RECT 181.650 539.400 183.450 545.400 ;
        RECT 182.250 538.500 183.450 539.400 ;
        RECT 172.950 537.450 179.550 538.500 ;
        RECT 172.950 536.700 174.750 537.450 ;
        RECT 177.750 536.700 179.550 537.450 ;
        RECT 182.250 536.400 187.050 538.500 ;
        RECT 165.150 534.600 167.850 536.400 ;
        RECT 168.750 535.800 170.550 536.400 ;
        RECT 168.750 534.900 175.050 535.800 ;
        RECT 182.250 535.500 183.450 536.400 ;
        RECT 168.750 534.600 170.550 534.900 ;
        RECT 166.950 533.700 167.850 534.600 ;
        RECT 158.550 526.050 159.750 533.400 ;
        RECT 163.950 532.800 166.050 533.700 ;
        RECT 166.950 532.800 172.050 533.700 ;
        RECT 161.850 531.600 166.050 532.800 ;
        RECT 160.950 529.800 162.750 531.600 ;
        RECT 121.950 523.950 124.050 526.050 ;
        RECT 124.950 523.950 127.050 526.050 ;
        RECT 127.950 523.950 130.050 526.050 ;
        RECT 130.950 523.950 133.050 526.050 ;
        RECT 145.950 523.950 148.050 526.050 ;
        RECT 148.950 523.950 151.050 526.050 ;
        RECT 151.950 523.950 154.050 526.050 ;
        RECT 158.550 525.750 163.050 526.050 ;
        RECT 158.550 523.950 164.850 525.750 ;
        RECT 125.100 522.150 126.900 523.950 ;
        RECT 128.850 519.750 130.050 523.950 ;
        RECT 131.100 522.150 132.900 523.950 ;
        RECT 146.100 522.150 147.900 523.950 ;
        RECT 128.850 518.700 132.600 519.750 ;
        RECT 103.950 514.500 106.050 516.600 ;
        RECT 94.200 513.600 95.250 514.500 ;
        RECT 103.950 513.600 105.000 514.500 ;
        RECT 85.650 510.600 87.450 513.600 ;
        RECT 93.450 510.600 95.250 513.600 ;
        RECT 101.250 512.700 105.000 513.600 ;
        RECT 101.250 510.600 103.050 512.700 ;
        RECT 109.050 510.600 110.850 516.600 ;
        RECT 122.400 515.700 130.200 517.050 ;
        RECT 122.400 510.600 124.200 515.700 ;
        RECT 128.400 510.600 130.200 515.700 ;
        RECT 131.400 516.600 132.600 518.700 ;
        RECT 149.400 518.700 150.600 523.950 ;
        RECT 152.100 522.150 153.900 523.950 ;
        RECT 149.400 517.800 153.600 518.700 ;
        RECT 131.400 510.600 133.200 516.600 ;
        RECT 151.800 510.600 153.600 517.800 ;
        RECT 158.550 516.600 159.750 523.950 ;
        RECT 171.150 520.200 172.050 532.800 ;
        RECT 174.150 532.800 175.050 534.900 ;
        RECT 175.950 534.300 183.450 535.500 ;
        RECT 175.950 533.700 177.750 534.300 ;
        RECT 190.050 533.400 191.850 545.400 ;
        RECT 174.150 532.500 182.550 532.800 ;
        RECT 190.950 532.500 191.850 533.400 ;
        RECT 174.150 531.900 191.850 532.500 ;
        RECT 180.750 531.300 191.850 531.900 ;
        RECT 180.750 531.000 182.550 531.300 ;
        RECT 178.950 524.400 181.050 526.050 ;
        RECT 178.950 523.200 186.900 524.400 ;
        RECT 187.950 523.950 190.050 526.050 ;
        RECT 185.100 522.600 186.900 523.200 ;
        RECT 188.100 522.150 189.900 523.950 ;
        RECT 182.100 521.400 183.900 522.000 ;
        RECT 188.100 521.400 189.000 522.150 ;
        RECT 182.100 520.200 189.000 521.400 ;
        RECT 171.150 519.000 183.150 520.200 ;
        RECT 171.150 518.400 172.950 519.000 ;
        RECT 182.100 517.200 183.150 519.000 ;
        RECT 158.550 510.600 160.350 516.600 ;
        RECT 163.950 515.700 166.050 516.600 ;
        RECT 163.950 514.500 167.700 515.700 ;
        RECT 178.350 515.550 180.150 516.300 ;
        RECT 166.650 513.600 167.700 514.500 ;
        RECT 175.200 514.500 180.150 515.550 ;
        RECT 181.650 515.400 183.450 517.200 ;
        RECT 190.950 516.600 191.850 531.300 ;
        RECT 206.400 539.400 208.200 545.400 ;
        RECT 226.800 539.400 228.600 545.400 ;
        RECT 248.400 539.400 250.200 545.400 ;
        RECT 203.100 526.050 204.900 527.850 ;
        RECT 206.400 526.050 207.600 539.400 ;
        RECT 221.100 526.050 222.900 527.850 ;
        RECT 226.950 526.050 228.150 539.400 ;
        RECT 248.400 532.500 249.600 539.400 ;
        RECT 254.400 533.400 256.200 545.400 ;
        RECT 248.400 531.600 254.100 532.500 ;
        RECT 252.150 530.700 254.100 531.600 ;
        RECT 248.100 526.050 249.900 527.850 ;
        RECT 202.950 523.950 205.050 526.050 ;
        RECT 205.950 523.950 208.050 526.050 ;
        RECT 220.950 523.950 223.050 526.050 ;
        RECT 223.950 523.950 226.050 526.050 ;
        RECT 226.950 523.950 229.050 526.050 ;
        RECT 229.950 523.950 232.050 526.050 ;
        RECT 247.950 523.950 250.050 526.050 ;
        RECT 184.950 514.500 187.050 516.600 ;
        RECT 175.200 513.600 176.250 514.500 ;
        RECT 184.950 513.600 186.000 514.500 ;
        RECT 166.650 510.600 168.450 513.600 ;
        RECT 174.450 510.600 176.250 513.600 ;
        RECT 182.250 512.700 186.000 513.600 ;
        RECT 182.250 510.600 184.050 512.700 ;
        RECT 190.050 510.600 191.850 516.600 ;
        RECT 206.400 513.600 207.600 523.950 ;
        RECT 224.100 522.150 225.900 523.950 ;
        RECT 227.850 519.750 229.050 523.950 ;
        RECT 230.100 522.150 231.900 523.950 ;
        RECT 227.850 518.700 231.600 519.750 ;
        RECT 221.400 515.700 229.200 517.050 ;
        RECT 206.400 510.600 208.200 513.600 ;
        RECT 221.400 510.600 223.200 515.700 ;
        RECT 227.400 510.600 229.200 515.700 ;
        RECT 230.400 516.600 231.600 518.700 ;
        RECT 252.150 519.300 253.050 530.700 ;
        RECT 255.000 526.050 256.200 533.400 ;
        RECT 272.400 539.400 274.200 545.400 ;
        RECT 293.400 539.400 295.200 545.400 ;
        RECT 272.400 526.050 273.600 539.400 ;
        RECT 290.100 526.050 291.900 527.850 ;
        RECT 293.400 526.050 294.600 539.400 ;
        RECT 311.700 534.600 313.500 545.400 ;
        RECT 311.700 533.400 315.300 534.600 ;
        RECT 301.950 531.450 304.050 532.050 ;
        RECT 310.950 531.450 313.050 532.050 ;
        RECT 301.950 530.550 313.050 531.450 ;
        RECT 301.950 529.950 304.050 530.550 ;
        RECT 310.950 529.950 313.050 530.550 ;
        RECT 311.100 526.050 312.900 527.850 ;
        RECT 314.400 526.050 315.300 533.400 ;
        RECT 320.550 533.400 322.350 545.400 ;
        RECT 328.050 539.400 329.850 545.400 ;
        RECT 325.950 537.300 329.850 539.400 ;
        RECT 335.850 538.500 337.650 545.400 ;
        RECT 343.650 539.400 345.450 545.400 ;
        RECT 344.250 538.500 345.450 539.400 ;
        RECT 334.950 537.450 341.550 538.500 ;
        RECT 334.950 536.700 336.750 537.450 ;
        RECT 339.750 536.700 341.550 537.450 ;
        RECT 344.250 536.400 349.050 538.500 ;
        RECT 327.150 534.600 329.850 536.400 ;
        RECT 330.750 535.800 332.550 536.400 ;
        RECT 330.750 534.900 337.050 535.800 ;
        RECT 344.250 535.500 345.450 536.400 ;
        RECT 330.750 534.600 332.550 534.900 ;
        RECT 328.950 533.700 329.850 534.600 ;
        RECT 317.100 526.050 318.900 527.850 ;
        RECT 320.550 526.050 321.750 533.400 ;
        RECT 325.950 532.800 328.050 533.700 ;
        RECT 328.950 532.800 334.050 533.700 ;
        RECT 323.850 531.600 328.050 532.800 ;
        RECT 322.950 529.800 324.750 531.600 ;
        RECT 253.950 523.950 256.200 526.050 ;
        RECT 268.950 523.950 271.050 526.050 ;
        RECT 271.950 523.950 274.050 526.050 ;
        RECT 274.950 523.950 277.050 526.050 ;
        RECT 289.950 523.950 292.050 526.050 ;
        RECT 292.950 523.950 295.050 526.050 ;
        RECT 310.950 523.950 313.050 526.050 ;
        RECT 313.950 523.950 316.050 526.050 ;
        RECT 316.950 523.950 319.050 526.050 ;
        RECT 320.550 525.750 325.050 526.050 ;
        RECT 320.550 523.950 326.850 525.750 ;
        RECT 252.150 518.400 254.100 519.300 ;
        RECT 248.400 517.500 254.100 518.400 ;
        RECT 230.400 510.600 232.200 516.600 ;
        RECT 248.400 513.600 249.600 517.500 ;
        RECT 255.000 516.600 256.200 523.950 ;
        RECT 269.100 522.150 270.900 523.950 ;
        RECT 272.400 518.700 273.600 523.950 ;
        RECT 275.100 522.150 276.900 523.950 ;
        RECT 280.950 519.450 283.050 520.050 ;
        RECT 289.950 519.450 292.050 520.050 ;
        RECT 272.400 517.800 276.600 518.700 ;
        RECT 280.950 518.550 292.050 519.450 ;
        RECT 280.950 517.950 283.050 518.550 ;
        RECT 289.950 517.950 292.050 518.550 ;
        RECT 248.400 510.600 250.200 513.600 ;
        RECT 254.400 510.600 256.200 516.600 ;
        RECT 274.800 510.600 276.600 517.800 ;
        RECT 293.400 513.600 294.600 523.950 ;
        RECT 314.400 513.600 315.300 523.950 ;
        RECT 320.550 516.600 321.750 523.950 ;
        RECT 333.150 520.200 334.050 532.800 ;
        RECT 336.150 532.800 337.050 534.900 ;
        RECT 337.950 534.300 345.450 535.500 ;
        RECT 337.950 533.700 339.750 534.300 ;
        RECT 352.050 533.400 353.850 545.400 ;
        RECT 370.800 539.400 372.600 545.400 ;
        RECT 336.150 532.500 344.550 532.800 ;
        RECT 352.950 532.500 353.850 533.400 ;
        RECT 336.150 531.900 353.850 532.500 ;
        RECT 342.750 531.300 353.850 531.900 ;
        RECT 342.750 531.000 344.550 531.300 ;
        RECT 340.950 524.400 343.050 526.050 ;
        RECT 340.950 523.200 348.900 524.400 ;
        RECT 349.950 523.950 352.050 526.050 ;
        RECT 347.100 522.600 348.900 523.200 ;
        RECT 350.100 522.150 351.900 523.950 ;
        RECT 344.100 521.400 345.900 522.000 ;
        RECT 350.100 521.400 351.000 522.150 ;
        RECT 344.100 520.200 351.000 521.400 ;
        RECT 333.150 519.000 345.150 520.200 ;
        RECT 333.150 518.400 334.950 519.000 ;
        RECT 344.100 517.200 345.150 519.000 ;
        RECT 293.400 510.600 295.200 513.600 ;
        RECT 313.800 510.600 315.600 513.600 ;
        RECT 320.550 510.600 322.350 516.600 ;
        RECT 325.950 515.700 328.050 516.600 ;
        RECT 325.950 514.500 329.700 515.700 ;
        RECT 340.350 515.550 342.150 516.300 ;
        RECT 328.650 513.600 329.700 514.500 ;
        RECT 337.200 514.500 342.150 515.550 ;
        RECT 343.650 515.400 345.450 517.200 ;
        RECT 352.950 516.600 353.850 531.300 ;
        RECT 371.400 526.050 372.600 539.400 ;
        RECT 388.800 533.400 390.600 545.400 ;
        RECT 410.400 539.400 412.200 545.400 ;
        RECT 389.400 526.050 390.600 533.400 ;
        RECT 410.850 526.050 412.050 539.400 ;
        RECT 420.150 533.400 421.950 545.400 ;
        RECT 428.550 539.400 430.350 545.400 ;
        RECT 428.550 538.500 429.750 539.400 ;
        RECT 436.350 538.500 438.150 545.400 ;
        RECT 444.150 539.400 445.950 545.400 ;
        RECT 424.950 536.400 429.750 538.500 ;
        RECT 432.450 537.450 439.050 538.500 ;
        RECT 432.450 536.700 434.250 537.450 ;
        RECT 437.250 536.700 439.050 537.450 ;
        RECT 444.150 537.300 448.050 539.400 ;
        RECT 428.550 535.500 429.750 536.400 ;
        RECT 441.450 535.800 443.250 536.400 ;
        RECT 428.550 534.300 436.050 535.500 ;
        RECT 434.250 533.700 436.050 534.300 ;
        RECT 436.950 534.900 443.250 535.800 ;
        RECT 420.150 532.500 421.050 533.400 ;
        RECT 436.950 532.800 437.850 534.900 ;
        RECT 441.450 534.600 443.250 534.900 ;
        RECT 444.150 534.600 446.850 536.400 ;
        RECT 444.150 533.700 445.050 534.600 ;
        RECT 429.450 532.500 437.850 532.800 ;
        RECT 420.150 531.900 437.850 532.500 ;
        RECT 439.950 532.800 445.050 533.700 ;
        RECT 445.950 532.800 448.050 533.700 ;
        RECT 451.650 533.400 453.450 545.400 ;
        RECT 420.150 531.300 431.250 531.900 ;
        RECT 416.100 526.050 417.900 527.850 ;
        RECT 367.950 523.950 370.050 526.050 ;
        RECT 370.950 523.950 373.050 526.050 ;
        RECT 373.950 523.950 376.050 526.050 ;
        RECT 388.950 523.950 391.050 526.050 ;
        RECT 391.950 523.950 394.050 526.050 ;
        RECT 406.950 523.950 409.050 526.050 ;
        RECT 409.950 523.950 412.050 526.050 ;
        RECT 412.950 523.950 415.050 526.050 ;
        RECT 415.950 523.950 418.050 526.050 ;
        RECT 368.100 522.150 369.900 523.950 ;
        RECT 371.400 518.700 372.600 523.950 ;
        RECT 374.100 522.150 375.900 523.950 ;
        RECT 346.950 514.500 349.050 516.600 ;
        RECT 337.200 513.600 338.250 514.500 ;
        RECT 346.950 513.600 348.000 514.500 ;
        RECT 328.650 510.600 330.450 513.600 ;
        RECT 336.450 510.600 338.250 513.600 ;
        RECT 344.250 512.700 348.000 513.600 ;
        RECT 344.250 510.600 346.050 512.700 ;
        RECT 352.050 510.600 353.850 516.600 ;
        RECT 368.400 517.800 372.600 518.700 ;
        RECT 373.950 519.450 376.050 520.050 ;
        RECT 382.950 519.450 385.050 520.050 ;
        RECT 373.950 518.550 385.050 519.450 ;
        RECT 373.950 517.950 376.050 518.550 ;
        RECT 382.950 517.950 385.050 518.550 ;
        RECT 368.400 510.600 370.200 517.800 ;
        RECT 389.400 516.600 390.600 523.950 ;
        RECT 392.100 522.150 393.900 523.950 ;
        RECT 407.100 522.150 408.900 523.950 ;
        RECT 409.950 519.750 411.150 523.950 ;
        RECT 413.100 522.150 414.900 523.950 ;
        RECT 407.400 518.700 411.150 519.750 ;
        RECT 407.400 516.600 408.600 518.700 ;
        RECT 388.800 510.600 390.600 516.600 ;
        RECT 406.800 510.600 408.600 516.600 ;
        RECT 409.800 515.700 417.600 517.050 ;
        RECT 409.800 510.600 411.600 515.700 ;
        RECT 415.800 510.600 417.600 515.700 ;
        RECT 420.150 516.600 421.050 531.300 ;
        RECT 429.450 531.000 431.250 531.300 ;
        RECT 421.950 523.950 424.050 526.050 ;
        RECT 430.950 524.400 433.050 526.050 ;
        RECT 422.100 522.150 423.900 523.950 ;
        RECT 425.100 523.200 433.050 524.400 ;
        RECT 425.100 522.600 426.900 523.200 ;
        RECT 423.000 521.400 423.900 522.150 ;
        RECT 428.100 521.400 429.900 522.000 ;
        RECT 423.000 520.200 429.900 521.400 ;
        RECT 439.950 520.200 440.850 532.800 ;
        RECT 445.950 531.600 450.150 532.800 ;
        RECT 449.250 529.800 451.050 531.600 ;
        RECT 452.250 526.050 453.450 533.400 ;
        RECT 467.400 539.400 469.200 545.400 ;
        RECT 490.800 539.400 492.600 545.400 ;
        RECT 512.400 539.400 514.200 545.400 ;
        RECT 467.400 526.050 468.600 539.400 ;
        RECT 491.400 526.050 492.600 539.400 ;
        RECT 493.950 531.450 496.050 532.200 ;
        RECT 508.950 531.450 511.050 532.050 ;
        RECT 493.950 530.550 511.050 531.450 ;
        RECT 493.950 530.100 496.050 530.550 ;
        RECT 508.950 529.950 511.050 530.550 ;
        RECT 496.950 528.450 501.000 529.050 ;
        RECT 496.950 526.950 501.450 528.450 ;
        RECT 448.950 525.750 453.450 526.050 ;
        RECT 447.150 523.950 453.450 525.750 ;
        RECT 463.950 523.950 466.050 526.050 ;
        RECT 466.950 523.950 469.050 526.050 ;
        RECT 469.950 523.950 472.050 526.050 ;
        RECT 487.950 523.950 490.050 526.050 ;
        RECT 490.950 523.950 493.050 526.050 ;
        RECT 493.950 523.950 496.050 526.050 ;
        RECT 428.850 519.000 440.850 520.200 ;
        RECT 428.850 517.200 429.900 519.000 ;
        RECT 439.050 518.400 440.850 519.000 ;
        RECT 420.150 510.600 421.950 516.600 ;
        RECT 424.950 514.500 427.050 516.600 ;
        RECT 428.550 515.400 430.350 517.200 ;
        RECT 452.250 516.600 453.450 523.950 ;
        RECT 464.100 522.150 465.900 523.950 ;
        RECT 467.400 518.700 468.600 523.950 ;
        RECT 470.100 522.150 471.900 523.950 ;
        RECT 488.100 522.150 489.900 523.950 ;
        RECT 491.400 518.700 492.600 523.950 ;
        RECT 494.100 522.150 495.900 523.950 ;
        RECT 500.550 523.050 501.450 526.950 ;
        RECT 512.850 526.050 514.050 539.400 ;
        RECT 522.150 533.400 523.950 545.400 ;
        RECT 530.550 539.400 532.350 545.400 ;
        RECT 530.550 538.500 531.750 539.400 ;
        RECT 538.350 538.500 540.150 545.400 ;
        RECT 546.150 539.400 547.950 545.400 ;
        RECT 526.950 536.400 531.750 538.500 ;
        RECT 534.450 537.450 541.050 538.500 ;
        RECT 534.450 536.700 536.250 537.450 ;
        RECT 539.250 536.700 541.050 537.450 ;
        RECT 546.150 537.300 550.050 539.400 ;
        RECT 530.550 535.500 531.750 536.400 ;
        RECT 543.450 535.800 545.250 536.400 ;
        RECT 530.550 534.300 538.050 535.500 ;
        RECT 536.250 533.700 538.050 534.300 ;
        RECT 538.950 534.900 545.250 535.800 ;
        RECT 522.150 532.500 523.050 533.400 ;
        RECT 538.950 532.800 539.850 534.900 ;
        RECT 543.450 534.600 545.250 534.900 ;
        RECT 546.150 534.600 548.850 536.400 ;
        RECT 546.150 533.700 547.050 534.600 ;
        RECT 531.450 532.500 539.850 532.800 ;
        RECT 522.150 531.900 539.850 532.500 ;
        RECT 541.950 532.800 547.050 533.700 ;
        RECT 547.950 532.800 550.050 533.700 ;
        RECT 553.650 533.400 555.450 545.400 ;
        RECT 571.800 539.400 573.600 545.400 ;
        RECT 522.150 531.300 533.250 531.900 ;
        RECT 518.100 526.050 519.900 527.850 ;
        RECT 508.950 523.950 511.050 526.050 ;
        RECT 511.950 523.950 514.050 526.050 ;
        RECT 514.950 523.950 517.050 526.050 ;
        RECT 517.950 523.950 520.050 526.050 ;
        RECT 496.950 521.550 501.450 523.050 ;
        RECT 509.100 522.150 510.900 523.950 ;
        RECT 496.950 520.950 501.000 521.550 ;
        RECT 511.950 519.750 513.150 523.950 ;
        RECT 515.100 522.150 516.900 523.950 ;
        RECT 467.400 517.800 471.600 518.700 ;
        RECT 431.850 515.550 433.650 516.300 ;
        RECT 445.950 515.700 448.050 516.600 ;
        RECT 431.850 514.500 436.800 515.550 ;
        RECT 426.000 513.600 427.050 514.500 ;
        RECT 435.750 513.600 436.800 514.500 ;
        RECT 444.300 514.500 448.050 515.700 ;
        RECT 444.300 513.600 445.350 514.500 ;
        RECT 426.000 512.700 429.750 513.600 ;
        RECT 427.950 510.600 429.750 512.700 ;
        RECT 435.750 510.600 437.550 513.600 ;
        RECT 443.550 510.600 445.350 513.600 ;
        RECT 451.650 510.600 453.450 516.600 ;
        RECT 469.800 510.600 471.600 517.800 ;
        RECT 488.400 517.800 492.600 518.700 ;
        RECT 509.400 518.700 513.150 519.750 ;
        RECT 475.950 513.450 478.050 517.050 ;
        RECT 481.950 513.450 484.050 514.050 ;
        RECT 475.950 513.000 484.050 513.450 ;
        RECT 476.550 512.550 484.050 513.000 ;
        RECT 481.950 511.950 484.050 512.550 ;
        RECT 488.400 510.600 490.200 517.800 ;
        RECT 509.400 516.600 510.600 518.700 ;
        RECT 508.800 510.600 510.600 516.600 ;
        RECT 511.800 515.700 519.600 517.050 ;
        RECT 511.800 510.600 513.600 515.700 ;
        RECT 517.800 510.600 519.600 515.700 ;
        RECT 522.150 516.600 523.050 531.300 ;
        RECT 531.450 531.000 533.250 531.300 ;
        RECT 523.950 523.950 526.050 526.050 ;
        RECT 532.950 524.400 535.050 526.050 ;
        RECT 524.100 522.150 525.900 523.950 ;
        RECT 527.100 523.200 535.050 524.400 ;
        RECT 527.100 522.600 528.900 523.200 ;
        RECT 525.000 521.400 525.900 522.150 ;
        RECT 530.100 521.400 531.900 522.000 ;
        RECT 525.000 520.200 531.900 521.400 ;
        RECT 541.950 520.200 542.850 532.800 ;
        RECT 547.950 531.600 552.150 532.800 ;
        RECT 551.250 529.800 553.050 531.600 ;
        RECT 554.250 526.050 555.450 533.400 ;
        RECT 566.100 526.050 567.900 527.850 ;
        RECT 571.950 526.050 573.150 539.400 ;
        RECT 592.800 533.400 594.600 545.400 ;
        RECT 598.800 539.400 600.600 545.400 ;
        RECT 616.800 539.400 618.600 545.400 ;
        RECT 577.950 528.450 580.050 529.050 ;
        RECT 589.950 528.450 592.050 529.050 ;
        RECT 577.950 527.550 592.050 528.450 ;
        RECT 577.950 526.950 580.050 527.550 ;
        RECT 550.950 525.750 555.450 526.050 ;
        RECT 549.150 523.950 555.450 525.750 ;
        RECT 565.950 523.950 568.050 526.050 ;
        RECT 568.950 523.950 571.050 526.050 ;
        RECT 571.950 523.950 574.050 526.050 ;
        RECT 574.950 523.950 577.050 526.050 ;
        RECT 530.850 519.000 542.850 520.200 ;
        RECT 530.850 517.200 531.900 519.000 ;
        RECT 541.050 518.400 542.850 519.000 ;
        RECT 522.150 510.600 523.950 516.600 ;
        RECT 526.950 514.500 529.050 516.600 ;
        RECT 530.550 515.400 532.350 517.200 ;
        RECT 554.250 516.600 555.450 523.950 ;
        RECT 569.100 522.150 570.900 523.950 ;
        RECT 572.850 519.750 574.050 523.950 ;
        RECT 575.100 522.150 576.900 523.950 ;
        RECT 587.550 523.050 588.450 527.550 ;
        RECT 589.950 526.950 592.050 527.550 ;
        RECT 593.400 526.050 594.300 533.400 ;
        RECT 596.100 526.050 597.900 527.850 ;
        RECT 592.950 523.950 595.050 526.050 ;
        RECT 595.950 523.950 598.050 526.050 ;
        RECT 587.550 521.550 592.050 523.050 ;
        RECT 588.000 520.950 592.050 521.550 ;
        RECT 572.850 518.700 576.600 519.750 ;
        RECT 533.850 515.550 535.650 516.300 ;
        RECT 547.950 515.700 550.050 516.600 ;
        RECT 533.850 514.500 538.800 515.550 ;
        RECT 528.000 513.600 529.050 514.500 ;
        RECT 537.750 513.600 538.800 514.500 ;
        RECT 546.300 514.500 550.050 515.700 ;
        RECT 546.300 513.600 547.350 514.500 ;
        RECT 528.000 512.700 531.750 513.600 ;
        RECT 529.950 510.600 531.750 512.700 ;
        RECT 537.750 510.600 539.550 513.600 ;
        RECT 545.550 510.600 547.350 513.600 ;
        RECT 553.650 510.600 555.450 516.600 ;
        RECT 566.400 515.700 574.200 517.050 ;
        RECT 566.400 510.600 568.200 515.700 ;
        RECT 572.400 510.600 574.200 515.700 ;
        RECT 575.400 516.600 576.600 518.700 ;
        RECT 593.400 516.600 594.300 523.950 ;
        RECT 599.700 519.300 600.600 539.400 ;
        RECT 617.700 539.100 618.600 539.400 ;
        RECT 622.800 539.400 624.600 545.400 ;
        RECT 641.400 539.400 643.200 545.400 ;
        RECT 661.800 539.400 663.600 545.400 ;
        RECT 682.800 539.400 684.600 545.400 ;
        RECT 701.400 539.400 703.200 545.400 ;
        RECT 622.800 539.100 624.300 539.400 ;
        RECT 617.700 538.200 624.300 539.100 ;
        RECT 601.950 534.450 604.050 535.050 ;
        RECT 610.950 534.450 613.050 535.050 ;
        RECT 601.950 533.550 613.050 534.450 ;
        RECT 601.950 532.950 604.050 533.550 ;
        RECT 610.950 532.950 613.050 533.550 ;
        RECT 617.700 526.050 618.600 538.200 ;
        RECT 623.100 526.050 624.900 527.850 ;
        RECT 638.100 526.050 639.900 527.850 ;
        RECT 641.400 526.050 642.600 539.400 ;
        RECT 662.400 526.050 663.600 539.400 ;
        RECT 677.100 526.050 678.900 527.850 ;
        RECT 682.950 526.050 684.150 539.400 ;
        RECT 701.400 532.500 702.600 539.400 ;
        RECT 707.400 533.400 709.200 545.400 ;
        RECT 727.800 539.400 729.600 545.400 ;
        RECT 749.400 539.400 751.200 545.400 ;
        RECT 685.950 531.450 688.050 532.050 ;
        RECT 691.950 531.450 694.050 532.050 ;
        RECT 701.400 531.600 707.100 532.500 ;
        RECT 685.950 530.550 694.050 531.450 ;
        RECT 685.950 529.950 688.050 530.550 ;
        RECT 691.950 529.950 694.050 530.550 ;
        RECT 705.150 530.700 707.100 531.600 ;
        RECT 701.100 526.050 702.900 527.850 ;
        RECT 601.950 523.950 604.050 526.050 ;
        RECT 616.950 523.950 619.050 526.050 ;
        RECT 619.950 523.950 622.050 526.050 ;
        RECT 622.950 523.950 625.050 526.050 ;
        RECT 625.950 523.950 628.050 526.050 ;
        RECT 637.950 523.950 640.050 526.050 ;
        RECT 640.950 523.950 643.050 526.050 ;
        RECT 658.950 523.950 661.050 526.050 ;
        RECT 661.950 523.950 664.050 526.050 ;
        RECT 664.950 523.950 667.050 526.050 ;
        RECT 676.950 523.950 679.050 526.050 ;
        RECT 679.950 523.950 682.050 526.050 ;
        RECT 682.950 523.950 685.050 526.050 ;
        RECT 685.950 523.950 688.050 526.050 ;
        RECT 700.950 523.950 703.050 526.050 ;
        RECT 602.100 522.150 603.900 523.950 ;
        RECT 617.700 520.200 618.600 523.950 ;
        RECT 620.100 522.150 621.900 523.950 ;
        RECT 626.100 522.150 627.900 523.950 ;
        RECT 596.100 518.400 603.600 519.300 ;
        RECT 617.700 519.000 621.000 520.200 ;
        RECT 596.100 517.500 597.900 518.400 ;
        RECT 575.400 510.600 577.200 516.600 ;
        RECT 593.400 514.800 596.100 516.600 ;
        RECT 594.300 510.600 596.100 514.800 ;
        RECT 601.800 510.600 603.600 518.400 ;
        RECT 619.200 510.600 621.000 519.000 ;
        RECT 641.400 513.600 642.600 523.950 ;
        RECT 659.100 522.150 660.900 523.950 ;
        RECT 662.400 518.700 663.600 523.950 ;
        RECT 665.100 522.150 666.900 523.950 ;
        RECT 680.100 522.150 681.900 523.950 ;
        RECT 683.850 519.750 685.050 523.950 ;
        RECT 686.100 522.150 687.900 523.950 ;
        RECT 683.850 518.700 687.600 519.750 ;
        RECT 659.400 517.800 663.600 518.700 ;
        RECT 641.400 510.600 643.200 513.600 ;
        RECT 659.400 510.600 661.200 517.800 ;
        RECT 677.400 515.700 685.200 517.050 ;
        RECT 677.400 510.600 679.200 515.700 ;
        RECT 683.400 510.600 685.200 515.700 ;
        RECT 686.400 516.600 687.600 518.700 ;
        RECT 705.150 519.300 706.050 530.700 ;
        RECT 708.000 526.050 709.200 533.400 ;
        RECT 722.100 526.050 723.900 527.850 ;
        RECT 727.950 526.050 729.150 539.400 ;
        RECT 706.950 523.950 709.200 526.050 ;
        RECT 721.950 523.950 724.050 526.050 ;
        RECT 724.950 523.950 727.050 526.050 ;
        RECT 727.950 523.950 730.050 526.050 ;
        RECT 730.950 523.950 733.050 526.050 ;
        RECT 745.950 523.950 748.050 526.050 ;
        RECT 705.150 518.400 707.100 519.300 ;
        RECT 701.400 517.500 707.100 518.400 ;
        RECT 686.400 510.600 688.200 516.600 ;
        RECT 701.400 513.600 702.600 517.500 ;
        RECT 708.000 516.600 709.200 523.950 ;
        RECT 725.100 522.150 726.900 523.950 ;
        RECT 728.850 519.750 730.050 523.950 ;
        RECT 731.100 522.150 732.900 523.950 ;
        RECT 746.100 522.150 747.900 523.950 ;
        RECT 728.850 518.700 732.600 519.750 ;
        RECT 749.400 519.300 750.300 539.400 ;
        RECT 755.400 533.400 757.200 545.400 ;
        RECT 775.800 539.400 777.600 545.400 ;
        RECT 796.800 539.400 798.600 545.400 ;
        RECT 752.100 526.050 753.900 527.850 ;
        RECT 755.700 526.050 756.600 533.400 ;
        RECT 776.400 526.050 777.600 539.400 ;
        RECT 781.950 528.450 786.000 529.050 ;
        RECT 781.950 526.950 786.450 528.450 ;
        RECT 751.950 523.950 754.050 526.050 ;
        RECT 754.950 523.950 757.050 526.050 ;
        RECT 772.950 523.950 775.050 526.050 ;
        RECT 775.950 523.950 778.050 526.050 ;
        RECT 778.950 523.950 781.050 526.050 ;
        RECT 701.400 510.600 703.200 513.600 ;
        RECT 707.400 510.600 709.200 516.600 ;
        RECT 722.400 515.700 730.200 517.050 ;
        RECT 722.400 510.600 724.200 515.700 ;
        RECT 728.400 510.600 730.200 515.700 ;
        RECT 731.400 516.600 732.600 518.700 ;
        RECT 746.400 518.400 753.900 519.300 ;
        RECT 731.400 510.600 733.200 516.600 ;
        RECT 746.400 510.600 748.200 518.400 ;
        RECT 752.100 517.500 753.900 518.400 ;
        RECT 755.700 516.600 756.600 523.950 ;
        RECT 773.100 522.150 774.900 523.950 ;
        RECT 776.400 518.700 777.600 523.950 ;
        RECT 779.100 522.150 780.900 523.950 ;
        RECT 785.550 523.050 786.450 526.950 ;
        RECT 797.400 526.050 798.600 539.400 ;
        RECT 815.400 539.400 817.200 545.400 ;
        RECT 793.950 523.950 796.050 526.050 ;
        RECT 796.950 523.950 799.050 526.050 ;
        RECT 799.950 523.950 802.050 526.050 ;
        RECT 811.950 523.950 814.050 526.050 ;
        RECT 781.950 521.550 786.450 523.050 ;
        RECT 794.100 522.150 795.900 523.950 ;
        RECT 781.950 520.950 786.000 521.550 ;
        RECT 797.400 518.700 798.600 523.950 ;
        RECT 800.100 522.150 801.900 523.950 ;
        RECT 753.900 514.800 756.600 516.600 ;
        RECT 773.400 517.800 777.600 518.700 ;
        RECT 794.400 517.800 798.600 518.700 ;
        RECT 799.950 519.450 802.050 520.050 ;
        RECT 808.950 519.450 811.050 523.050 ;
        RECT 812.100 522.150 813.900 523.950 ;
        RECT 799.950 519.000 811.050 519.450 ;
        RECT 815.400 519.300 816.300 539.400 ;
        RECT 821.400 533.400 823.200 545.400 ;
        RECT 838.800 533.400 840.600 545.400 ;
        RECT 841.800 534.300 843.600 545.400 ;
        RECT 847.800 534.300 849.600 545.400 ;
        RECT 865.800 539.400 867.600 545.400 ;
        RECT 841.800 533.400 849.600 534.300 ;
        RECT 818.100 526.050 819.900 527.850 ;
        RECT 821.700 526.050 822.600 533.400 ;
        RECT 839.400 526.050 840.300 533.400 ;
        RECT 845.100 526.050 846.900 527.850 ;
        RECT 860.100 526.050 861.900 527.850 ;
        RECT 865.950 526.050 867.150 539.400 ;
        RECT 817.950 523.950 820.050 526.050 ;
        RECT 820.950 523.950 823.050 526.050 ;
        RECT 838.950 523.950 841.050 526.050 ;
        RECT 841.950 523.950 844.050 526.050 ;
        RECT 844.950 523.950 847.050 526.050 ;
        RECT 847.950 523.950 850.050 526.050 ;
        RECT 859.950 523.950 862.050 526.050 ;
        RECT 862.950 523.950 865.050 526.050 ;
        RECT 865.950 523.950 868.050 526.050 ;
        RECT 868.950 523.950 871.050 526.050 ;
        RECT 799.950 518.550 810.450 519.000 ;
        RECT 799.950 517.950 802.050 518.550 ;
        RECT 812.400 518.400 819.900 519.300 ;
        RECT 753.900 510.600 755.700 514.800 ;
        RECT 773.400 510.600 775.200 517.800 ;
        RECT 794.400 510.600 796.200 517.800 ;
        RECT 812.400 510.600 814.200 518.400 ;
        RECT 818.100 517.500 819.900 518.400 ;
        RECT 821.700 516.600 822.600 523.950 ;
        RECT 819.900 514.800 822.600 516.600 ;
        RECT 839.400 516.600 840.300 523.950 ;
        RECT 842.100 522.150 843.900 523.950 ;
        RECT 848.100 522.150 849.900 523.950 ;
        RECT 863.100 522.150 864.900 523.950 ;
        RECT 841.950 519.450 844.050 520.050 ;
        RECT 853.950 519.450 856.050 520.050 ;
        RECT 841.950 518.550 856.050 519.450 ;
        RECT 866.850 519.750 868.050 523.950 ;
        RECT 869.100 522.150 870.900 523.950 ;
        RECT 866.850 518.700 870.600 519.750 ;
        RECT 841.950 517.950 844.050 518.550 ;
        RECT 853.950 517.950 856.050 518.550 ;
        RECT 839.400 515.400 844.500 516.600 ;
        RECT 819.900 510.600 821.700 514.800 ;
        RECT 842.700 510.600 844.500 515.400 ;
        RECT 860.400 515.700 868.200 517.050 ;
        RECT 860.400 510.600 862.200 515.700 ;
        RECT 866.400 510.600 868.200 515.700 ;
        RECT 869.400 516.600 870.600 518.700 ;
        RECT 869.400 510.600 871.200 516.600 ;
        RECT 3.150 500.400 4.950 506.400 ;
        RECT 10.950 504.300 12.750 506.400 ;
        RECT 9.000 503.400 12.750 504.300 ;
        RECT 18.750 503.400 20.550 506.400 ;
        RECT 26.550 503.400 28.350 506.400 ;
        RECT 9.000 502.500 10.050 503.400 ;
        RECT 18.750 502.500 19.800 503.400 ;
        RECT 7.950 500.400 10.050 502.500 ;
        RECT 3.150 485.700 4.050 500.400 ;
        RECT 11.550 499.800 13.350 501.600 ;
        RECT 14.850 501.450 19.800 502.500 ;
        RECT 27.300 502.500 28.350 503.400 ;
        RECT 14.850 500.700 16.650 501.450 ;
        RECT 27.300 501.300 31.050 502.500 ;
        RECT 28.950 500.400 31.050 501.300 ;
        RECT 34.650 500.400 36.450 506.400 ;
        RECT 11.850 498.000 12.900 499.800 ;
        RECT 22.050 498.000 23.850 498.600 ;
        RECT 11.850 496.800 23.850 498.000 ;
        RECT 6.000 495.600 12.900 496.800 ;
        RECT 6.000 494.850 6.900 495.600 ;
        RECT 11.100 495.000 12.900 495.600 ;
        RECT 5.100 493.050 6.900 494.850 ;
        RECT 8.100 493.800 9.900 494.400 ;
        RECT 4.950 490.950 7.050 493.050 ;
        RECT 8.100 492.600 16.050 493.800 ;
        RECT 13.950 490.950 16.050 492.600 ;
        RECT 12.450 485.700 14.250 486.000 ;
        RECT 3.150 485.100 14.250 485.700 ;
        RECT 3.150 484.500 20.850 485.100 ;
        RECT 3.150 483.600 4.050 484.500 ;
        RECT 12.450 484.200 20.850 484.500 ;
        RECT 3.150 471.600 4.950 483.600 ;
        RECT 17.250 482.700 19.050 483.300 ;
        RECT 11.550 481.500 19.050 482.700 ;
        RECT 19.950 482.100 20.850 484.200 ;
        RECT 22.950 484.200 23.850 496.800 ;
        RECT 35.250 493.050 36.450 500.400 ;
        RECT 52.800 499.200 54.600 506.400 ;
        RECT 50.400 498.300 54.600 499.200 ;
        RECT 71.400 499.200 73.200 506.400 ;
        RECT 80.550 500.400 82.350 506.400 ;
        RECT 88.650 503.400 90.450 506.400 ;
        RECT 96.450 503.400 98.250 506.400 ;
        RECT 104.250 504.300 106.050 506.400 ;
        RECT 104.250 503.400 108.000 504.300 ;
        RECT 88.650 502.500 89.700 503.400 ;
        RECT 85.950 501.300 89.700 502.500 ;
        RECT 97.200 502.500 98.250 503.400 ;
        RECT 106.950 502.500 108.000 503.400 ;
        RECT 97.200 501.450 102.150 502.500 ;
        RECT 85.950 500.400 88.050 501.300 ;
        RECT 100.350 500.700 102.150 501.450 ;
        RECT 71.400 498.300 75.600 499.200 ;
        RECT 47.100 493.050 48.900 494.850 ;
        RECT 50.400 493.050 51.600 498.300 ;
        RECT 53.100 493.050 54.900 494.850 ;
        RECT 71.100 493.050 72.900 494.850 ;
        RECT 74.400 493.050 75.600 498.300 ;
        RECT 77.100 493.050 78.900 494.850 ;
        RECT 80.550 493.050 81.750 500.400 ;
        RECT 103.650 499.800 105.450 501.600 ;
        RECT 106.950 500.400 109.050 502.500 ;
        RECT 112.050 500.400 113.850 506.400 ;
        RECT 131.700 501.600 133.500 506.400 ;
        RECT 152.400 503.400 154.200 506.400 ;
        RECT 173.400 503.400 175.200 506.400 ;
        RECT 93.150 498.000 94.950 498.600 ;
        RECT 104.100 498.000 105.150 499.800 ;
        RECT 93.150 496.800 105.150 498.000 ;
        RECT 30.150 491.250 36.450 493.050 ;
        RECT 31.950 490.950 36.450 491.250 ;
        RECT 46.950 490.950 49.050 493.050 ;
        RECT 49.950 490.950 52.050 493.050 ;
        RECT 52.950 490.950 55.050 493.050 ;
        RECT 70.950 490.950 73.050 493.050 ;
        RECT 73.950 490.950 76.050 493.050 ;
        RECT 76.950 490.950 79.050 493.050 ;
        RECT 80.550 491.250 86.850 493.050 ;
        RECT 80.550 490.950 85.050 491.250 ;
        RECT 32.250 485.400 34.050 487.200 ;
        RECT 28.950 484.200 33.150 485.400 ;
        RECT 22.950 483.300 28.050 484.200 ;
        RECT 28.950 483.300 31.050 484.200 ;
        RECT 35.250 483.600 36.450 490.950 ;
        RECT 27.150 482.400 28.050 483.300 ;
        RECT 24.450 482.100 26.250 482.400 ;
        RECT 11.550 480.600 12.750 481.500 ;
        RECT 19.950 481.200 26.250 482.100 ;
        RECT 24.450 480.600 26.250 481.200 ;
        RECT 27.150 480.600 29.850 482.400 ;
        RECT 7.950 478.500 12.750 480.600 ;
        RECT 15.450 479.550 17.250 480.300 ;
        RECT 20.250 479.550 22.050 480.300 ;
        RECT 15.450 478.500 22.050 479.550 ;
        RECT 11.550 477.600 12.750 478.500 ;
        RECT 11.550 471.600 13.350 477.600 ;
        RECT 19.350 471.600 21.150 478.500 ;
        RECT 27.150 477.600 31.050 479.700 ;
        RECT 27.150 471.600 28.950 477.600 ;
        RECT 34.650 471.600 36.450 483.600 ;
        RECT 50.400 477.600 51.600 490.950 ;
        RECT 74.400 477.600 75.600 490.950 ;
        RECT 50.400 471.600 52.200 477.600 ;
        RECT 73.800 471.600 75.600 477.600 ;
        RECT 80.550 483.600 81.750 490.950 ;
        RECT 82.950 485.400 84.750 487.200 ;
        RECT 83.850 484.200 88.050 485.400 ;
        RECT 93.150 484.200 94.050 496.800 ;
        RECT 104.100 495.600 111.000 496.800 ;
        RECT 104.100 495.000 105.900 495.600 ;
        RECT 110.100 494.850 111.000 495.600 ;
        RECT 107.100 493.800 108.900 494.400 ;
        RECT 100.950 492.600 108.900 493.800 ;
        RECT 110.100 493.050 111.900 494.850 ;
        RECT 100.950 490.950 103.050 492.600 ;
        RECT 109.950 490.950 112.050 493.050 ;
        RECT 102.750 485.700 104.550 486.000 ;
        RECT 112.950 485.700 113.850 500.400 ;
        RECT 128.400 500.400 133.500 501.600 ;
        RECT 128.400 493.050 129.300 500.400 ;
        RECT 131.100 493.050 132.900 494.850 ;
        RECT 137.100 493.050 138.900 494.850 ;
        RECT 152.700 493.050 153.600 503.400 ;
        RECT 173.400 493.050 174.600 503.400 ;
        RECT 196.800 499.200 198.600 506.400 ;
        RECT 216.300 502.200 218.100 506.400 ;
        RECT 194.400 498.300 198.600 499.200 ;
        RECT 215.400 500.400 218.100 502.200 ;
        RECT 191.100 493.050 192.900 494.850 ;
        RECT 194.400 493.050 195.600 498.300 ;
        RECT 199.950 495.450 202.050 499.050 ;
        RECT 211.950 495.450 214.050 499.050 ;
        RECT 199.950 495.000 214.050 495.450 ;
        RECT 197.100 493.050 198.900 494.850 ;
        RECT 200.550 494.550 213.450 495.000 ;
        RECT 215.400 493.050 216.300 500.400 ;
        RECT 218.100 498.600 219.900 499.500 ;
        RECT 223.800 498.600 225.600 506.400 ;
        RECT 241.800 499.200 243.600 506.400 ;
        RECT 259.800 500.400 261.600 506.400 ;
        RECT 218.100 497.700 225.600 498.600 ;
        RECT 239.400 498.300 243.600 499.200 ;
        RECT 260.400 498.300 261.600 500.400 ;
        RECT 262.800 501.300 264.600 506.400 ;
        RECT 268.800 501.300 270.600 506.400 ;
        RECT 262.800 499.950 270.600 501.300 ;
        RECT 272.550 500.400 274.350 506.400 ;
        RECT 280.650 503.400 282.450 506.400 ;
        RECT 288.450 503.400 290.250 506.400 ;
        RECT 296.250 504.300 298.050 506.400 ;
        RECT 296.250 503.400 300.000 504.300 ;
        RECT 280.650 502.500 281.700 503.400 ;
        RECT 277.950 501.300 281.700 502.500 ;
        RECT 289.200 502.500 290.250 503.400 ;
        RECT 298.950 502.500 300.000 503.400 ;
        RECT 289.200 501.450 294.150 502.500 ;
        RECT 277.950 500.400 280.050 501.300 ;
        RECT 292.350 500.700 294.150 501.450 ;
        RECT 127.950 490.950 130.050 493.050 ;
        RECT 130.950 490.950 133.050 493.050 ;
        RECT 133.950 490.950 136.050 493.050 ;
        RECT 136.950 490.950 139.050 493.050 ;
        RECT 148.950 490.950 151.050 493.050 ;
        RECT 151.950 490.950 154.050 493.050 ;
        RECT 154.950 490.950 157.050 493.050 ;
        RECT 169.950 490.950 172.050 493.050 ;
        RECT 172.950 490.950 175.050 493.050 ;
        RECT 190.950 490.950 193.050 493.050 ;
        RECT 193.950 490.950 196.050 493.050 ;
        RECT 196.950 490.950 199.050 493.050 ;
        RECT 214.950 490.950 217.050 493.050 ;
        RECT 217.950 490.950 220.050 493.050 ;
        RECT 102.750 485.100 113.850 485.700 ;
        RECT 80.550 471.600 82.350 483.600 ;
        RECT 85.950 483.300 88.050 484.200 ;
        RECT 88.950 483.300 94.050 484.200 ;
        RECT 96.150 484.500 113.850 485.100 ;
        RECT 96.150 484.200 104.550 484.500 ;
        RECT 88.950 482.400 89.850 483.300 ;
        RECT 87.150 480.600 89.850 482.400 ;
        RECT 90.750 482.100 92.550 482.400 ;
        RECT 96.150 482.100 97.050 484.200 ;
        RECT 112.950 483.600 113.850 484.500 ;
        RECT 128.400 483.600 129.300 490.950 ;
        RECT 134.100 489.150 135.900 490.950 ;
        RECT 149.100 489.150 150.900 490.950 ;
        RECT 152.700 483.600 153.600 490.950 ;
        RECT 155.100 489.150 156.900 490.950 ;
        RECT 170.100 489.150 171.900 490.950 ;
        RECT 90.750 481.200 97.050 482.100 ;
        RECT 97.950 482.700 99.750 483.300 ;
        RECT 97.950 481.500 105.450 482.700 ;
        RECT 90.750 480.600 92.550 481.200 ;
        RECT 104.250 480.600 105.450 481.500 ;
        RECT 85.950 477.600 89.850 479.700 ;
        RECT 94.950 479.550 96.750 480.300 ;
        RECT 99.750 479.550 101.550 480.300 ;
        RECT 94.950 478.500 101.550 479.550 ;
        RECT 104.250 478.500 109.050 480.600 ;
        RECT 88.050 471.600 89.850 477.600 ;
        RECT 95.850 471.600 97.650 478.500 ;
        RECT 104.250 477.600 105.450 478.500 ;
        RECT 103.650 471.600 105.450 477.600 ;
        RECT 112.050 471.600 113.850 483.600 ;
        RECT 127.800 471.600 129.600 483.600 ;
        RECT 130.800 482.700 138.600 483.600 ;
        RECT 130.800 471.600 132.600 482.700 ;
        RECT 136.800 471.600 138.600 482.700 ;
        RECT 152.700 482.400 156.300 483.600 ;
        RECT 154.500 471.600 156.300 482.400 ;
        RECT 173.400 477.600 174.600 490.950 ;
        RECT 178.950 489.450 181.050 490.050 ;
        RECT 187.950 489.450 190.050 490.050 ;
        RECT 178.950 488.550 190.050 489.450 ;
        RECT 178.950 487.950 181.050 488.550 ;
        RECT 187.950 487.950 190.050 488.550 ;
        RECT 194.400 477.600 195.600 490.950 ;
        RECT 215.400 483.600 216.300 490.950 ;
        RECT 218.100 489.150 219.900 490.950 ;
        RECT 173.400 471.600 175.200 477.600 ;
        RECT 194.400 471.600 196.200 477.600 ;
        RECT 214.800 471.600 216.600 483.600 ;
        RECT 221.700 477.600 222.600 497.700 ;
        RECT 224.100 493.050 225.900 494.850 ;
        RECT 236.100 493.050 237.900 494.850 ;
        RECT 239.400 493.050 240.600 498.300 ;
        RECT 260.400 497.250 264.150 498.300 ;
        RECT 242.100 493.050 243.900 494.850 ;
        RECT 260.100 493.050 261.900 494.850 ;
        RECT 262.950 493.050 264.150 497.250 ;
        RECT 266.100 493.050 267.900 494.850 ;
        RECT 272.550 493.050 273.750 500.400 ;
        RECT 295.650 499.800 297.450 501.600 ;
        RECT 298.950 500.400 301.050 502.500 ;
        RECT 304.050 500.400 305.850 506.400 ;
        RECT 285.150 498.000 286.950 498.600 ;
        RECT 296.100 498.000 297.150 499.800 ;
        RECT 285.150 496.800 297.150 498.000 ;
        RECT 223.950 490.950 226.050 493.050 ;
        RECT 235.950 490.950 238.050 493.050 ;
        RECT 238.950 490.950 241.050 493.050 ;
        RECT 241.950 490.950 244.050 493.050 ;
        RECT 259.950 490.950 262.050 493.050 ;
        RECT 262.950 490.950 265.050 493.050 ;
        RECT 265.950 490.950 268.050 493.050 ;
        RECT 268.950 490.950 271.050 493.050 ;
        RECT 272.550 491.250 278.850 493.050 ;
        RECT 272.550 490.950 277.050 491.250 ;
        RECT 220.800 471.600 222.600 477.600 ;
        RECT 239.400 477.600 240.600 490.950 ;
        RECT 263.850 477.600 265.050 490.950 ;
        RECT 269.100 489.150 270.900 490.950 ;
        RECT 272.550 483.600 273.750 490.950 ;
        RECT 274.950 485.400 276.750 487.200 ;
        RECT 275.850 484.200 280.050 485.400 ;
        RECT 285.150 484.200 286.050 496.800 ;
        RECT 296.100 495.600 303.000 496.800 ;
        RECT 296.100 495.000 297.900 495.600 ;
        RECT 302.100 494.850 303.000 495.600 ;
        RECT 299.100 493.800 300.900 494.400 ;
        RECT 292.950 492.600 300.900 493.800 ;
        RECT 302.100 493.050 303.900 494.850 ;
        RECT 292.950 490.950 295.050 492.600 ;
        RECT 301.950 490.950 304.050 493.050 ;
        RECT 294.750 485.700 296.550 486.000 ;
        RECT 304.950 485.700 305.850 500.400 ;
        RECT 317.400 501.300 319.200 506.400 ;
        RECT 323.400 501.300 325.200 506.400 ;
        RECT 317.400 499.950 325.200 501.300 ;
        RECT 326.400 500.400 328.200 506.400 ;
        RECT 331.950 501.450 334.050 502.050 ;
        RECT 337.950 501.450 340.050 502.050 ;
        RECT 331.950 500.550 340.050 501.450 ;
        RECT 326.400 498.300 327.600 500.400 ;
        RECT 331.950 499.950 334.050 500.550 ;
        RECT 337.950 499.950 340.050 500.550 ;
        RECT 343.800 500.400 345.600 506.400 ;
        RECT 323.850 497.250 327.600 498.300 ;
        RECT 344.400 498.300 345.600 500.400 ;
        RECT 346.800 501.300 348.600 506.400 ;
        RECT 352.800 501.300 354.600 506.400 ;
        RECT 346.800 499.950 354.600 501.300 ;
        RECT 356.550 500.400 358.350 506.400 ;
        RECT 364.650 503.400 366.450 506.400 ;
        RECT 372.450 503.400 374.250 506.400 ;
        RECT 380.250 504.300 382.050 506.400 ;
        RECT 380.250 503.400 384.000 504.300 ;
        RECT 364.650 502.500 365.700 503.400 ;
        RECT 361.950 501.300 365.700 502.500 ;
        RECT 373.200 502.500 374.250 503.400 ;
        RECT 382.950 502.500 384.000 503.400 ;
        RECT 373.200 501.450 378.150 502.500 ;
        RECT 361.950 500.400 364.050 501.300 ;
        RECT 376.350 500.700 378.150 501.450 ;
        RECT 344.400 497.250 348.150 498.300 ;
        RECT 320.100 493.050 321.900 494.850 ;
        RECT 323.850 493.050 325.050 497.250 ;
        RECT 326.100 493.050 327.900 494.850 ;
        RECT 344.100 493.050 345.900 494.850 ;
        RECT 346.950 493.050 348.150 497.250 ;
        RECT 350.100 493.050 351.900 494.850 ;
        RECT 356.550 493.050 357.750 500.400 ;
        RECT 379.650 499.800 381.450 501.600 ;
        RECT 382.950 500.400 385.050 502.500 ;
        RECT 388.050 500.400 389.850 506.400 ;
        RECT 369.150 498.000 370.950 498.600 ;
        RECT 380.100 498.000 381.150 499.800 ;
        RECT 369.150 496.800 381.150 498.000 ;
        RECT 316.950 490.950 319.050 493.050 ;
        RECT 319.950 490.950 322.050 493.050 ;
        RECT 322.950 490.950 325.050 493.050 ;
        RECT 325.950 490.950 328.050 493.050 ;
        RECT 343.950 490.950 346.050 493.050 ;
        RECT 346.950 490.950 349.050 493.050 ;
        RECT 349.950 490.950 352.050 493.050 ;
        RECT 352.950 490.950 355.050 493.050 ;
        RECT 356.550 491.250 362.850 493.050 ;
        RECT 356.550 490.950 361.050 491.250 ;
        RECT 317.100 489.150 318.900 490.950 ;
        RECT 294.750 485.100 305.850 485.700 ;
        RECT 239.400 471.600 241.200 477.600 ;
        RECT 263.400 471.600 265.200 477.600 ;
        RECT 272.550 471.600 274.350 483.600 ;
        RECT 277.950 483.300 280.050 484.200 ;
        RECT 280.950 483.300 286.050 484.200 ;
        RECT 288.150 484.500 305.850 485.100 ;
        RECT 288.150 484.200 296.550 484.500 ;
        RECT 280.950 482.400 281.850 483.300 ;
        RECT 279.150 480.600 281.850 482.400 ;
        RECT 282.750 482.100 284.550 482.400 ;
        RECT 288.150 482.100 289.050 484.200 ;
        RECT 304.950 483.600 305.850 484.500 ;
        RECT 282.750 481.200 289.050 482.100 ;
        RECT 289.950 482.700 291.750 483.300 ;
        RECT 289.950 481.500 297.450 482.700 ;
        RECT 282.750 480.600 284.550 481.200 ;
        RECT 296.250 480.600 297.450 481.500 ;
        RECT 277.950 477.600 281.850 479.700 ;
        RECT 286.950 479.550 288.750 480.300 ;
        RECT 291.750 479.550 293.550 480.300 ;
        RECT 286.950 478.500 293.550 479.550 ;
        RECT 296.250 478.500 301.050 480.600 ;
        RECT 280.050 471.600 281.850 477.600 ;
        RECT 287.850 471.600 289.650 478.500 ;
        RECT 296.250 477.600 297.450 478.500 ;
        RECT 295.650 471.600 297.450 477.600 ;
        RECT 304.050 471.600 305.850 483.600 ;
        RECT 322.950 477.600 324.150 490.950 ;
        RECT 347.850 477.600 349.050 490.950 ;
        RECT 353.100 489.150 354.900 490.950 ;
        RECT 356.550 483.600 357.750 490.950 ;
        RECT 358.950 485.400 360.750 487.200 ;
        RECT 359.850 484.200 364.050 485.400 ;
        RECT 369.150 484.200 370.050 496.800 ;
        RECT 380.100 495.600 387.000 496.800 ;
        RECT 380.100 495.000 381.900 495.600 ;
        RECT 386.100 494.850 387.000 495.600 ;
        RECT 383.100 493.800 384.900 494.400 ;
        RECT 376.950 492.600 384.900 493.800 ;
        RECT 386.100 493.050 387.900 494.850 ;
        RECT 376.950 490.950 379.050 492.600 ;
        RECT 385.950 490.950 388.050 493.050 ;
        RECT 378.750 485.700 380.550 486.000 ;
        RECT 388.950 485.700 389.850 500.400 ;
        RECT 404.400 499.200 406.200 506.400 ;
        RECT 424.800 500.400 426.600 506.400 ;
        RECT 404.400 498.300 408.600 499.200 ;
        RECT 404.100 493.050 405.900 494.850 ;
        RECT 407.400 493.050 408.600 498.300 ;
        RECT 425.400 498.300 426.600 500.400 ;
        RECT 427.800 501.300 429.600 506.400 ;
        RECT 433.800 501.300 435.600 506.400 ;
        RECT 427.800 499.950 435.600 501.300 ;
        RECT 448.800 500.400 450.600 506.400 ;
        RECT 449.400 498.300 450.600 500.400 ;
        RECT 451.800 501.300 453.600 506.400 ;
        RECT 457.800 501.300 459.600 506.400 ;
        RECT 451.800 499.950 459.600 501.300 ;
        RECT 462.150 500.400 463.950 506.400 ;
        RECT 469.950 504.300 471.750 506.400 ;
        RECT 468.000 503.400 471.750 504.300 ;
        RECT 477.750 503.400 479.550 506.400 ;
        RECT 485.550 503.400 487.350 506.400 ;
        RECT 468.000 502.500 469.050 503.400 ;
        RECT 477.750 502.500 478.800 503.400 ;
        RECT 466.950 500.400 469.050 502.500 ;
        RECT 425.400 497.250 429.150 498.300 ;
        RECT 449.400 497.250 453.150 498.300 ;
        RECT 410.100 493.050 411.900 494.850 ;
        RECT 425.100 493.050 426.900 494.850 ;
        RECT 427.950 493.050 429.150 497.250 ;
        RECT 431.100 493.050 432.900 494.850 ;
        RECT 449.100 493.050 450.900 494.850 ;
        RECT 451.950 493.050 453.150 497.250 ;
        RECT 455.100 493.050 456.900 494.850 ;
        RECT 403.950 490.950 406.050 493.050 ;
        RECT 406.950 490.950 409.050 493.050 ;
        RECT 409.950 490.950 412.050 493.050 ;
        RECT 424.950 490.950 427.050 493.050 ;
        RECT 427.950 490.950 430.050 493.050 ;
        RECT 430.950 490.950 433.050 493.050 ;
        RECT 433.950 490.950 436.050 493.050 ;
        RECT 448.950 490.950 451.050 493.050 ;
        RECT 451.950 490.950 454.050 493.050 ;
        RECT 454.950 490.950 457.050 493.050 ;
        RECT 457.950 490.950 460.050 493.050 ;
        RECT 378.750 485.100 389.850 485.700 ;
        RECT 322.800 471.600 324.600 477.600 ;
        RECT 347.400 471.600 349.200 477.600 ;
        RECT 356.550 471.600 358.350 483.600 ;
        RECT 361.950 483.300 364.050 484.200 ;
        RECT 364.950 483.300 370.050 484.200 ;
        RECT 372.150 484.500 389.850 485.100 ;
        RECT 372.150 484.200 380.550 484.500 ;
        RECT 364.950 482.400 365.850 483.300 ;
        RECT 363.150 480.600 365.850 482.400 ;
        RECT 366.750 482.100 368.550 482.400 ;
        RECT 372.150 482.100 373.050 484.200 ;
        RECT 388.950 483.600 389.850 484.500 ;
        RECT 366.750 481.200 373.050 482.100 ;
        RECT 373.950 482.700 375.750 483.300 ;
        RECT 373.950 481.500 381.450 482.700 ;
        RECT 366.750 480.600 368.550 481.200 ;
        RECT 380.250 480.600 381.450 481.500 ;
        RECT 361.950 477.600 365.850 479.700 ;
        RECT 370.950 479.550 372.750 480.300 ;
        RECT 375.750 479.550 377.550 480.300 ;
        RECT 370.950 478.500 377.550 479.550 ;
        RECT 380.250 478.500 385.050 480.600 ;
        RECT 364.050 471.600 365.850 477.600 ;
        RECT 371.850 471.600 373.650 478.500 ;
        RECT 380.250 477.600 381.450 478.500 ;
        RECT 379.650 471.600 381.450 477.600 ;
        RECT 388.050 471.600 389.850 483.600 ;
        RECT 407.400 477.600 408.600 490.950 ;
        RECT 409.950 483.450 412.050 484.050 ;
        RECT 424.950 483.450 427.050 484.050 ;
        RECT 409.950 482.550 427.050 483.450 ;
        RECT 409.950 481.950 412.050 482.550 ;
        RECT 424.950 481.950 427.050 482.550 ;
        RECT 428.850 477.600 430.050 490.950 ;
        RECT 434.100 489.150 435.900 490.950 ;
        RECT 452.850 477.600 454.050 490.950 ;
        RECT 458.100 489.150 459.900 490.950 ;
        RECT 462.150 485.700 463.050 500.400 ;
        RECT 470.550 499.800 472.350 501.600 ;
        RECT 473.850 501.450 478.800 502.500 ;
        RECT 486.300 502.500 487.350 503.400 ;
        RECT 473.850 500.700 475.650 501.450 ;
        RECT 486.300 501.300 490.050 502.500 ;
        RECT 487.950 500.400 490.050 501.300 ;
        RECT 493.650 500.400 495.450 506.400 ;
        RECT 470.850 498.000 471.900 499.800 ;
        RECT 481.050 498.000 482.850 498.600 ;
        RECT 470.850 496.800 482.850 498.000 ;
        RECT 465.000 495.600 471.900 496.800 ;
        RECT 465.000 494.850 465.900 495.600 ;
        RECT 470.100 495.000 471.900 495.600 ;
        RECT 464.100 493.050 465.900 494.850 ;
        RECT 467.100 493.800 468.900 494.400 ;
        RECT 463.950 490.950 466.050 493.050 ;
        RECT 467.100 492.600 475.050 493.800 ;
        RECT 472.950 490.950 475.050 492.600 ;
        RECT 471.450 485.700 473.250 486.000 ;
        RECT 462.150 485.100 473.250 485.700 ;
        RECT 462.150 484.500 479.850 485.100 ;
        RECT 462.150 483.600 463.050 484.500 ;
        RECT 471.450 484.200 479.850 484.500 ;
        RECT 406.800 471.600 408.600 477.600 ;
        RECT 428.400 471.600 430.200 477.600 ;
        RECT 452.400 471.600 454.200 477.600 ;
        RECT 462.150 471.600 463.950 483.600 ;
        RECT 476.250 482.700 478.050 483.300 ;
        RECT 470.550 481.500 478.050 482.700 ;
        RECT 478.950 482.100 479.850 484.200 ;
        RECT 481.950 484.200 482.850 496.800 ;
        RECT 494.250 493.050 495.450 500.400 ;
        RECT 506.400 501.300 508.200 506.400 ;
        RECT 512.400 501.300 514.200 506.400 ;
        RECT 506.400 499.950 514.200 501.300 ;
        RECT 515.400 500.400 517.200 506.400 ;
        RECT 533.400 500.400 535.200 506.400 ;
        RECT 548.400 503.400 550.200 506.400 ;
        RECT 515.400 498.300 516.600 500.400 ;
        RECT 512.850 497.250 516.600 498.300 ;
        RECT 509.100 493.050 510.900 494.850 ;
        RECT 512.850 493.050 514.050 497.250 ;
        RECT 515.100 493.050 516.900 494.850 ;
        RECT 530.100 493.050 531.900 494.850 ;
        RECT 533.400 493.050 534.600 500.400 ;
        RECT 548.400 499.500 549.600 503.400 ;
        RECT 554.400 500.400 556.200 506.400 ;
        RECT 548.400 498.600 554.100 499.500 ;
        RECT 552.150 497.700 554.100 498.600 ;
        RECT 489.150 491.250 495.450 493.050 ;
        RECT 490.950 490.950 495.450 491.250 ;
        RECT 505.950 490.950 508.050 493.050 ;
        RECT 508.950 490.950 511.050 493.050 ;
        RECT 511.950 490.950 514.050 493.050 ;
        RECT 514.950 490.950 517.050 493.050 ;
        RECT 529.950 490.950 532.050 493.050 ;
        RECT 532.950 490.950 535.050 493.050 ;
        RECT 547.950 490.950 550.050 493.050 ;
        RECT 491.250 485.400 493.050 487.200 ;
        RECT 487.950 484.200 492.150 485.400 ;
        RECT 481.950 483.300 487.050 484.200 ;
        RECT 487.950 483.300 490.050 484.200 ;
        RECT 494.250 483.600 495.450 490.950 ;
        RECT 506.100 489.150 507.900 490.950 ;
        RECT 486.150 482.400 487.050 483.300 ;
        RECT 483.450 482.100 485.250 482.400 ;
        RECT 470.550 480.600 471.750 481.500 ;
        RECT 478.950 481.200 485.250 482.100 ;
        RECT 483.450 480.600 485.250 481.200 ;
        RECT 486.150 480.600 488.850 482.400 ;
        RECT 466.950 478.500 471.750 480.600 ;
        RECT 474.450 479.550 476.250 480.300 ;
        RECT 479.250 479.550 481.050 480.300 ;
        RECT 474.450 478.500 481.050 479.550 ;
        RECT 470.550 477.600 471.750 478.500 ;
        RECT 470.550 471.600 472.350 477.600 ;
        RECT 478.350 471.600 480.150 478.500 ;
        RECT 486.150 477.600 490.050 479.700 ;
        RECT 486.150 471.600 487.950 477.600 ;
        RECT 493.650 471.600 495.450 483.600 ;
        RECT 511.950 477.600 513.150 490.950 ;
        RECT 533.400 483.600 534.600 490.950 ;
        RECT 548.100 489.150 549.900 490.950 ;
        RECT 552.150 486.300 553.050 497.700 ;
        RECT 555.000 493.050 556.200 500.400 ;
        RECT 572.400 499.200 574.200 506.400 ;
        RECT 592.800 500.400 594.600 506.400 ;
        RECT 572.400 498.300 576.600 499.200 ;
        RECT 572.100 493.050 573.900 494.850 ;
        RECT 575.400 493.050 576.600 498.300 ;
        RECT 580.950 495.450 583.050 499.050 ;
        RECT 593.400 498.300 594.600 500.400 ;
        RECT 595.800 501.300 597.600 506.400 ;
        RECT 601.800 501.300 603.600 506.400 ;
        RECT 595.800 499.950 603.600 501.300 ;
        RECT 614.400 501.300 616.200 506.400 ;
        RECT 620.400 501.300 622.200 506.400 ;
        RECT 614.400 499.950 622.200 501.300 ;
        RECT 623.400 500.400 625.200 506.400 ;
        RECT 623.400 498.300 624.600 500.400 ;
        RECT 643.800 499.200 645.600 506.400 ;
        RECT 593.400 497.250 597.150 498.300 ;
        RECT 580.950 495.000 588.450 495.450 ;
        RECT 578.100 493.050 579.900 494.850 ;
        RECT 581.550 494.550 588.450 495.000 ;
        RECT 553.950 490.950 556.200 493.050 ;
        RECT 571.950 490.950 574.050 493.050 ;
        RECT 574.950 490.950 577.050 493.050 ;
        RECT 577.950 490.950 580.050 493.050 ;
        RECT 552.150 485.400 554.100 486.300 ;
        RECT 548.400 484.500 554.100 485.400 ;
        RECT 511.800 471.600 513.600 477.600 ;
        RECT 533.400 471.600 535.200 483.600 ;
        RECT 548.400 477.600 549.600 484.500 ;
        RECT 555.000 483.600 556.200 490.950 ;
        RECT 548.400 471.600 550.200 477.600 ;
        RECT 554.400 471.600 556.200 483.600 ;
        RECT 575.400 477.600 576.600 490.950 ;
        RECT 587.550 490.050 588.450 494.550 ;
        RECT 593.100 493.050 594.900 494.850 ;
        RECT 595.950 493.050 597.150 497.250 ;
        RECT 620.850 497.250 624.600 498.300 ;
        RECT 641.400 498.300 645.600 499.200 ;
        RECT 604.950 495.450 609.000 496.050 ;
        RECT 599.100 493.050 600.900 494.850 ;
        RECT 604.950 493.950 609.450 495.450 ;
        RECT 592.950 490.950 595.050 493.050 ;
        RECT 595.950 490.950 598.050 493.050 ;
        RECT 598.950 490.950 601.050 493.050 ;
        RECT 601.950 490.950 604.050 493.050 ;
        RECT 587.550 488.550 592.050 490.050 ;
        RECT 588.000 487.950 592.050 488.550 ;
        RECT 586.950 486.450 589.050 487.050 ;
        RECT 592.950 486.450 595.050 487.050 ;
        RECT 586.950 485.550 595.050 486.450 ;
        RECT 586.950 484.950 589.050 485.550 ;
        RECT 592.950 484.950 595.050 485.550 ;
        RECT 583.950 483.450 586.050 484.050 ;
        RECT 589.950 483.450 592.050 484.050 ;
        RECT 583.950 482.550 592.050 483.450 ;
        RECT 583.950 481.950 586.050 482.550 ;
        RECT 589.950 481.950 592.050 482.550 ;
        RECT 596.850 477.600 598.050 490.950 ;
        RECT 602.100 489.150 603.900 490.950 ;
        RECT 608.550 490.050 609.450 493.950 ;
        RECT 617.100 493.050 618.900 494.850 ;
        RECT 620.850 493.050 622.050 497.250 ;
        RECT 623.100 493.050 624.900 494.850 ;
        RECT 638.100 493.050 639.900 494.850 ;
        RECT 641.400 493.050 642.600 498.300 ;
        RECT 666.000 498.000 667.800 506.400 ;
        RECT 688.800 499.200 690.600 506.400 ;
        RECT 694.950 504.450 697.050 505.050 ;
        RECT 694.950 504.000 705.450 504.450 ;
        RECT 694.950 503.550 706.050 504.000 ;
        RECT 694.950 502.950 697.050 503.550 ;
        RECT 703.950 499.950 706.050 503.550 ;
        RECT 707.400 501.300 709.200 506.400 ;
        RECT 713.400 501.300 715.200 506.400 ;
        RECT 707.400 499.950 715.200 501.300 ;
        RECT 716.400 500.400 718.200 506.400 ;
        RECT 736.500 501.600 738.300 506.400 ;
        RECT 759.300 502.200 761.100 506.400 ;
        RECT 736.500 500.400 741.600 501.600 ;
        RECT 676.950 498.450 679.050 499.050 ;
        RECT 682.950 498.450 685.050 499.050 ;
        RECT 666.000 496.800 669.300 498.000 ;
        RECT 676.950 497.550 685.050 498.450 ;
        RECT 676.950 496.950 679.050 497.550 ;
        RECT 682.950 496.950 685.050 497.550 ;
        RECT 686.400 498.300 690.600 499.200 ;
        RECT 716.400 498.300 717.600 500.400 ;
        RECT 644.100 493.050 645.900 494.850 ;
        RECT 659.100 493.050 660.900 494.850 ;
        RECT 665.100 493.050 666.900 494.850 ;
        RECT 668.400 493.050 669.300 496.800 ;
        RECT 683.100 493.050 684.900 494.850 ;
        RECT 686.400 493.050 687.600 498.300 ;
        RECT 713.850 497.250 717.600 498.300 ;
        RECT 724.950 498.450 727.050 499.050 ;
        RECT 736.950 498.450 739.050 499.050 ;
        RECT 724.950 497.550 739.050 498.450 ;
        RECT 689.100 493.050 690.900 494.850 ;
        RECT 710.100 493.050 711.900 494.850 ;
        RECT 713.850 493.050 715.050 497.250 ;
        RECT 724.950 496.950 727.050 497.550 ;
        RECT 736.950 496.950 739.050 497.550 ;
        RECT 716.100 493.050 717.900 494.850 ;
        RECT 731.100 493.050 732.900 494.850 ;
        RECT 737.100 493.050 738.900 494.850 ;
        RECT 740.700 493.050 741.600 500.400 ;
        RECT 758.400 500.400 761.100 502.200 ;
        RECT 758.400 493.050 759.300 500.400 ;
        RECT 761.100 498.600 762.900 499.500 ;
        RECT 766.800 498.600 768.600 506.400 ;
        RECT 784.200 500.400 786.000 506.400 ;
        RECT 809.400 503.400 811.200 506.400 ;
        RECT 761.100 497.700 768.600 498.600 ;
        RECT 613.950 490.950 616.050 493.050 ;
        RECT 616.950 490.950 619.050 493.050 ;
        RECT 619.950 490.950 622.050 493.050 ;
        RECT 622.950 490.950 625.050 493.050 ;
        RECT 637.950 490.950 640.050 493.050 ;
        RECT 640.950 490.950 643.050 493.050 ;
        RECT 643.950 490.950 646.050 493.050 ;
        RECT 658.950 490.950 661.050 493.050 ;
        RECT 661.950 490.950 664.050 493.050 ;
        RECT 664.950 490.950 667.050 493.050 ;
        RECT 667.950 490.950 670.050 493.050 ;
        RECT 682.950 490.950 685.050 493.050 ;
        RECT 685.950 490.950 688.050 493.050 ;
        RECT 688.950 490.950 691.050 493.050 ;
        RECT 706.950 490.950 709.050 493.050 ;
        RECT 709.950 490.950 712.050 493.050 ;
        RECT 712.950 490.950 715.050 493.050 ;
        RECT 715.950 490.950 718.050 493.050 ;
        RECT 730.950 490.950 733.050 493.050 ;
        RECT 733.950 490.950 736.050 493.050 ;
        RECT 736.950 490.950 739.050 493.050 ;
        RECT 739.950 490.950 742.050 493.050 ;
        RECT 757.950 490.950 760.050 493.050 ;
        RECT 760.950 490.950 763.050 493.050 ;
        RECT 608.550 488.550 613.050 490.050 ;
        RECT 614.100 489.150 615.900 490.950 ;
        RECT 609.000 487.950 613.050 488.550 ;
        RECT 619.950 477.600 621.150 490.950 ;
        RECT 622.950 486.450 625.050 487.050 ;
        RECT 637.950 486.450 640.050 486.750 ;
        RECT 622.950 485.550 640.050 486.450 ;
        RECT 622.950 484.950 625.050 485.550 ;
        RECT 637.950 484.650 640.050 485.550 ;
        RECT 641.400 477.600 642.600 490.950 ;
        RECT 662.100 489.150 663.900 490.950 ;
        RECT 668.400 478.800 669.300 490.950 ;
        RECT 662.700 477.900 669.300 478.800 ;
        RECT 662.700 477.600 664.200 477.900 ;
        RECT 574.800 471.600 576.600 477.600 ;
        RECT 596.400 471.600 598.200 477.600 ;
        RECT 619.800 471.600 621.600 477.600 ;
        RECT 641.400 471.600 643.200 477.600 ;
        RECT 662.400 471.600 664.200 477.600 ;
        RECT 668.400 477.600 669.300 477.900 ;
        RECT 686.400 477.600 687.600 490.950 ;
        RECT 707.100 489.150 708.900 490.950 ;
        RECT 694.950 486.450 697.050 487.050 ;
        RECT 706.950 486.450 709.050 487.050 ;
        RECT 694.950 485.550 709.050 486.450 ;
        RECT 694.950 484.950 697.050 485.550 ;
        RECT 706.950 484.950 709.050 485.550 ;
        RECT 712.950 477.600 714.150 490.950 ;
        RECT 734.100 489.150 735.900 490.950 ;
        RECT 740.700 483.600 741.600 490.950 ;
        RECT 758.400 483.600 759.300 490.950 ;
        RECT 761.100 489.150 762.900 490.950 ;
        RECT 731.400 482.700 739.200 483.600 ;
        RECT 668.400 471.600 670.200 477.600 ;
        RECT 686.400 471.600 688.200 477.600 ;
        RECT 712.800 471.600 714.600 477.600 ;
        RECT 731.400 471.600 733.200 482.700 ;
        RECT 737.400 471.600 739.200 482.700 ;
        RECT 740.400 471.600 742.200 483.600 ;
        RECT 757.800 471.600 759.600 483.600 ;
        RECT 764.700 477.600 765.600 497.700 ;
        RECT 767.100 493.050 768.900 494.850 ;
        RECT 779.100 493.050 780.900 494.850 ;
        RECT 784.950 493.050 786.000 500.400 ;
        RECT 790.950 498.450 793.050 499.050 ;
        RECT 805.950 498.450 808.050 499.050 ;
        RECT 790.950 497.550 808.050 498.450 ;
        RECT 790.950 496.950 793.050 497.550 ;
        RECT 805.950 496.950 808.050 497.550 ;
        RECT 791.100 493.050 792.900 494.850 ;
        RECT 809.700 493.050 810.600 503.400 ;
        RECT 832.800 499.200 834.600 506.400 ;
        RECT 850.800 500.400 852.600 506.400 ;
        RECT 830.400 498.300 834.600 499.200 ;
        RECT 851.400 498.300 852.600 500.400 ;
        RECT 853.800 501.300 855.600 506.400 ;
        RECT 859.800 501.300 861.600 506.400 ;
        RECT 853.800 499.950 861.600 501.300 ;
        RECT 827.100 493.050 828.900 494.850 ;
        RECT 830.400 493.050 831.600 498.300 ;
        RECT 851.400 497.250 855.150 498.300 ;
        RECT 833.100 493.050 834.900 494.850 ;
        RECT 851.100 493.050 852.900 494.850 ;
        RECT 853.950 493.050 855.150 497.250 ;
        RECT 879.000 498.000 880.800 506.400 ;
        RECT 879.000 496.800 882.300 498.000 ;
        RECT 867.000 495.450 871.050 496.050 ;
        RECT 857.100 493.050 858.900 494.850 ;
        RECT 866.550 493.950 871.050 495.450 ;
        RECT 766.950 490.950 769.050 493.050 ;
        RECT 778.950 490.950 781.050 493.050 ;
        RECT 781.950 490.950 784.050 493.050 ;
        RECT 784.950 490.950 787.050 493.050 ;
        RECT 787.950 490.950 790.050 493.050 ;
        RECT 790.950 490.950 793.050 493.050 ;
        RECT 805.950 490.950 808.050 493.050 ;
        RECT 808.950 490.950 811.050 493.050 ;
        RECT 811.950 490.950 814.050 493.050 ;
        RECT 826.950 490.950 829.050 493.050 ;
        RECT 829.950 490.950 832.050 493.050 ;
        RECT 832.950 490.950 835.050 493.050 ;
        RECT 850.950 490.950 853.050 493.050 ;
        RECT 853.950 490.950 856.050 493.050 ;
        RECT 856.950 490.950 859.050 493.050 ;
        RECT 859.950 490.950 862.050 493.050 ;
        RECT 782.100 489.150 783.900 490.950 ;
        RECT 766.950 486.450 769.050 487.050 ;
        RECT 781.950 486.450 784.050 487.050 ;
        RECT 766.950 485.550 784.050 486.450 ;
        RECT 766.950 484.950 769.050 485.550 ;
        RECT 781.950 484.950 784.050 485.550 ;
        RECT 785.100 485.400 786.000 490.950 ;
        RECT 788.100 489.150 789.900 490.950 ;
        RECT 806.100 489.150 807.900 490.950 ;
        RECT 785.100 484.500 790.200 485.400 ;
        RECT 766.950 483.450 769.050 483.900 ;
        RECT 772.950 483.450 775.050 484.050 ;
        RECT 766.950 482.550 775.050 483.450 ;
        RECT 766.950 481.800 769.050 482.550 ;
        RECT 772.950 481.950 775.050 482.550 ;
        RECT 779.400 482.400 787.200 483.300 ;
        RECT 763.800 471.600 765.600 477.600 ;
        RECT 779.400 471.600 781.200 482.400 ;
        RECT 785.400 472.500 787.200 482.400 ;
        RECT 788.400 473.400 790.200 484.500 ;
        RECT 809.700 483.600 810.600 490.950 ;
        RECT 812.100 489.150 813.900 490.950 ;
        RECT 817.950 486.450 820.050 487.050 ;
        RECT 826.950 486.450 829.050 487.050 ;
        RECT 817.950 485.550 829.050 486.450 ;
        RECT 817.950 484.950 820.050 485.550 ;
        RECT 826.950 484.950 829.050 485.550 ;
        RECT 791.400 472.500 793.200 483.600 ;
        RECT 809.700 482.400 813.300 483.600 ;
        RECT 785.400 471.600 793.200 472.500 ;
        RECT 811.500 471.600 813.300 482.400 ;
        RECT 830.400 477.600 831.600 490.950 ;
        RECT 854.850 477.600 856.050 490.950 ;
        RECT 860.100 489.150 861.900 490.950 ;
        RECT 866.550 490.050 867.450 493.950 ;
        RECT 872.100 493.050 873.900 494.850 ;
        RECT 878.100 493.050 879.900 494.850 ;
        RECT 881.400 493.050 882.300 496.800 ;
        RECT 883.950 495.450 888.000 496.050 ;
        RECT 883.950 493.950 888.450 495.450 ;
        RECT 871.950 490.950 874.050 493.050 ;
        RECT 874.950 490.950 877.050 493.050 ;
        RECT 877.950 490.950 880.050 493.050 ;
        RECT 880.950 490.950 883.050 493.050 ;
        RECT 866.550 488.550 871.050 490.050 ;
        RECT 875.100 489.150 876.900 490.950 ;
        RECT 867.000 487.950 871.050 488.550 ;
        RECT 881.400 478.800 882.300 490.950 ;
        RECT 887.550 490.050 888.450 493.950 ;
        RECT 883.950 488.550 888.450 490.050 ;
        RECT 883.950 487.950 888.000 488.550 ;
        RECT 875.700 477.900 882.300 478.800 ;
        RECT 875.700 477.600 877.200 477.900 ;
        RECT 830.400 471.600 832.200 477.600 ;
        RECT 854.400 471.600 856.200 477.600 ;
        RECT 875.400 471.600 877.200 477.600 ;
        RECT 881.400 477.600 882.300 477.900 ;
        RECT 881.400 471.600 883.200 477.600 ;
        RECT 3.150 455.400 4.950 467.400 ;
        RECT 11.550 461.400 13.350 467.400 ;
        RECT 11.550 460.500 12.750 461.400 ;
        RECT 19.350 460.500 21.150 467.400 ;
        RECT 27.150 461.400 28.950 467.400 ;
        RECT 7.950 458.400 12.750 460.500 ;
        RECT 15.450 459.450 22.050 460.500 ;
        RECT 15.450 458.700 17.250 459.450 ;
        RECT 20.250 458.700 22.050 459.450 ;
        RECT 27.150 459.300 31.050 461.400 ;
        RECT 11.550 457.500 12.750 458.400 ;
        RECT 24.450 457.800 26.250 458.400 ;
        RECT 11.550 456.300 19.050 457.500 ;
        RECT 17.250 455.700 19.050 456.300 ;
        RECT 19.950 456.900 26.250 457.800 ;
        RECT 3.150 454.500 4.050 455.400 ;
        RECT 19.950 454.800 20.850 456.900 ;
        RECT 24.450 456.600 26.250 456.900 ;
        RECT 27.150 456.600 29.850 458.400 ;
        RECT 27.150 455.700 28.050 456.600 ;
        RECT 12.450 454.500 20.850 454.800 ;
        RECT 3.150 453.900 20.850 454.500 ;
        RECT 22.950 454.800 28.050 455.700 ;
        RECT 28.950 454.800 31.050 455.700 ;
        RECT 34.650 455.400 36.450 467.400 ;
        RECT 53.400 461.400 55.200 467.400 ;
        RECT 3.150 453.300 14.250 453.900 ;
        RECT 3.150 438.600 4.050 453.300 ;
        RECT 12.450 453.000 14.250 453.300 ;
        RECT 4.950 445.950 7.050 448.050 ;
        RECT 13.950 446.400 16.050 448.050 ;
        RECT 5.100 444.150 6.900 445.950 ;
        RECT 8.100 445.200 16.050 446.400 ;
        RECT 8.100 444.600 9.900 445.200 ;
        RECT 6.000 443.400 6.900 444.150 ;
        RECT 11.100 443.400 12.900 444.000 ;
        RECT 6.000 442.200 12.900 443.400 ;
        RECT 22.950 442.200 23.850 454.800 ;
        RECT 28.950 453.600 33.150 454.800 ;
        RECT 32.250 451.800 34.050 453.600 ;
        RECT 35.250 448.050 36.450 455.400 ;
        RECT 53.850 448.050 55.050 461.400 ;
        RECT 73.800 455.400 75.600 467.400 ;
        RECT 79.800 461.400 81.600 467.400 ;
        RECT 59.100 448.050 60.900 449.850 ;
        RECT 73.800 448.050 75.000 455.400 ;
        RECT 80.400 454.500 81.600 461.400 ;
        RECT 92.400 456.300 94.200 467.400 ;
        RECT 99.900 456.300 101.700 467.400 ;
        RECT 107.400 456.600 109.200 467.400 ;
        RECT 92.400 455.100 97.200 456.300 ;
        RECT 99.900 455.400 103.200 456.300 ;
        RECT 75.900 453.600 81.600 454.500 ;
        RECT 95.100 454.200 97.200 455.100 ;
        RECT 75.900 452.700 77.850 453.600 ;
        RECT 95.100 453.300 100.500 454.200 ;
        RECT 31.950 447.750 36.450 448.050 ;
        RECT 30.150 445.950 36.450 447.750 ;
        RECT 49.950 445.950 52.050 448.050 ;
        RECT 52.950 445.950 55.050 448.050 ;
        RECT 55.950 445.950 58.050 448.050 ;
        RECT 58.950 445.950 61.050 448.050 ;
        RECT 73.800 445.950 76.050 448.050 ;
        RECT 11.850 441.000 23.850 442.200 ;
        RECT 11.850 439.200 12.900 441.000 ;
        RECT 22.050 440.400 23.850 441.000 ;
        RECT 3.150 432.600 4.950 438.600 ;
        RECT 7.950 436.500 10.050 438.600 ;
        RECT 11.550 437.400 13.350 439.200 ;
        RECT 35.250 438.600 36.450 445.950 ;
        RECT 50.100 444.150 51.900 445.950 ;
        RECT 52.950 441.750 54.150 445.950 ;
        RECT 56.100 444.150 57.900 445.950 ;
        RECT 50.400 440.700 54.150 441.750 ;
        RECT 50.400 438.600 51.600 440.700 ;
        RECT 14.850 437.550 16.650 438.300 ;
        RECT 28.950 437.700 31.050 438.600 ;
        RECT 14.850 436.500 19.800 437.550 ;
        RECT 9.000 435.600 10.050 436.500 ;
        RECT 18.750 435.600 19.800 436.500 ;
        RECT 27.300 436.500 31.050 437.700 ;
        RECT 27.300 435.600 28.350 436.500 ;
        RECT 9.000 434.700 12.750 435.600 ;
        RECT 10.950 432.600 12.750 434.700 ;
        RECT 18.750 432.600 20.550 435.600 ;
        RECT 26.550 432.600 28.350 435.600 ;
        RECT 34.650 432.600 36.450 438.600 ;
        RECT 49.800 432.600 51.600 438.600 ;
        RECT 52.800 437.700 60.600 439.050 ;
        RECT 52.800 432.600 54.600 437.700 ;
        RECT 58.800 432.600 60.600 437.700 ;
        RECT 73.800 438.600 75.000 445.950 ;
        RECT 76.950 441.300 77.850 452.700 ;
        RECT 98.700 451.200 100.500 453.300 ;
        RECT 102.000 450.900 103.200 455.400 ;
        RECT 104.100 455.400 109.200 456.600 ;
        RECT 124.800 456.600 126.600 467.400 ;
        RECT 124.800 455.400 129.600 456.600 ;
        RECT 104.100 454.500 106.200 455.400 ;
        RECT 127.500 454.500 129.600 455.400 ;
        RECT 132.300 455.400 134.100 467.400 ;
        RECT 139.800 456.300 141.600 467.400 ;
        RECT 154.800 461.400 156.600 467.400 ;
        RECT 137.100 455.400 141.600 456.300 ;
        RECT 132.300 453.900 133.500 455.400 ;
        RECT 132.000 453.000 133.500 453.900 ;
        RECT 137.100 453.300 139.200 455.400 ;
        RECT 101.400 450.300 103.500 450.900 ;
        RECT 112.950 450.450 115.050 451.050 ;
        RECT 132.000 450.900 132.900 453.000 ;
        RECT 80.100 448.050 81.900 449.850 ;
        RECT 97.200 448.200 99.000 450.000 ;
        RECT 100.350 448.800 103.500 450.300 ;
        RECT 107.550 449.700 115.050 450.450 ;
        RECT 107.100 449.550 115.050 449.700 ;
        RECT 79.950 445.950 82.050 448.050 ;
        RECT 92.400 445.800 94.500 447.900 ;
        RECT 97.200 446.100 99.300 448.200 ;
        RECT 92.700 445.200 94.500 445.800 ;
        RECT 92.700 444.000 99.300 445.200 ;
        RECT 97.200 443.100 99.300 444.000 ;
        RECT 75.900 440.400 77.850 441.300 ;
        RECT 94.650 441.000 96.750 441.600 ;
        RECT 97.650 441.300 99.450 443.100 ;
        RECT 100.350 442.200 101.250 448.800 ;
        RECT 107.100 447.900 108.900 449.550 ;
        RECT 112.950 448.950 115.050 449.550 ;
        RECT 125.100 448.050 126.900 449.850 ;
        RECT 130.800 448.800 132.900 450.900 ;
        RECT 133.800 451.500 135.900 451.800 ;
        RECT 133.800 449.700 137.700 451.500 ;
        RECT 102.300 446.100 104.100 447.900 ;
        RECT 102.150 444.000 104.250 446.100 ;
        RECT 106.950 445.800 109.050 447.900 ;
        RECT 118.950 447.450 123.000 448.050 ;
        RECT 124.950 447.450 127.050 448.050 ;
        RECT 131.400 447.900 133.800 448.800 ;
        RECT 118.950 446.550 127.050 447.450 ;
        RECT 118.950 445.950 123.000 446.550 ;
        RECT 124.950 445.950 127.050 446.550 ;
        RECT 129.600 445.200 131.400 447.000 ;
        RECT 129.750 443.100 131.850 445.200 ;
        RECT 132.750 442.200 133.800 447.900 ;
        RECT 134.700 447.900 136.500 448.500 ;
        RECT 155.400 448.050 156.600 461.400 ;
        RECT 170.400 461.400 172.200 467.400 ;
        RECT 170.400 454.500 171.600 461.400 ;
        RECT 176.400 455.400 178.200 467.400 ;
        RECT 197.400 461.400 199.200 467.400 ;
        RECT 218.400 461.400 220.200 467.400 ;
        RECT 170.400 453.600 176.100 454.500 ;
        RECT 174.150 452.700 176.100 453.600 ;
        RECT 158.100 448.050 159.900 449.850 ;
        RECT 170.100 448.050 171.900 449.850 ;
        RECT 139.500 447.900 141.600 448.050 ;
        RECT 134.700 446.700 141.600 447.900 ;
        RECT 139.500 445.950 141.600 446.700 ;
        RECT 154.950 445.950 157.050 448.050 ;
        RECT 157.950 445.950 160.050 448.050 ;
        RECT 169.950 445.950 172.050 448.050 ;
        RECT 75.900 439.500 81.600 440.400 ;
        RECT 73.800 432.600 75.600 438.600 ;
        RECT 80.400 435.600 81.600 439.500 ;
        RECT 79.800 432.600 81.600 435.600 ;
        RECT 92.400 439.500 96.750 441.000 ;
        RECT 100.350 440.100 103.500 442.200 ;
        RECT 92.400 438.600 93.900 439.500 ;
        RECT 92.400 432.600 94.200 438.600 ;
        RECT 100.350 438.000 101.400 440.100 ;
        RECT 104.700 439.800 106.800 441.900 ;
        RECT 104.700 438.600 109.200 439.800 ;
        RECT 127.500 439.500 129.600 440.700 ;
        RECT 130.800 440.100 133.800 442.200 ;
        RECT 134.700 443.400 136.500 445.200 ;
        RECT 139.800 444.150 141.600 445.950 ;
        RECT 134.700 441.300 136.800 443.400 ;
        RECT 134.700 440.400 141.000 441.300 ;
        RECT 99.600 432.600 101.400 438.000 ;
        RECT 107.400 432.600 109.200 438.600 ;
        RECT 124.800 438.600 129.600 439.500 ;
        RECT 132.600 438.600 133.800 440.100 ;
        RECT 139.800 438.600 141.000 440.400 ;
        RECT 124.800 432.600 126.600 438.600 ;
        RECT 132.300 432.600 134.100 438.600 ;
        RECT 139.800 432.600 141.600 438.600 ;
        RECT 155.400 435.600 156.600 445.950 ;
        RECT 174.150 441.300 175.050 452.700 ;
        RECT 177.000 448.050 178.200 455.400 ;
        RECT 197.850 448.050 199.050 461.400 ;
        RECT 203.100 448.050 204.900 449.850 ;
        RECT 218.400 448.050 219.600 461.400 ;
        RECT 227.550 455.400 229.350 467.400 ;
        RECT 235.050 461.400 236.850 467.400 ;
        RECT 232.950 459.300 236.850 461.400 ;
        RECT 242.850 460.500 244.650 467.400 ;
        RECT 250.650 461.400 252.450 467.400 ;
        RECT 251.250 460.500 252.450 461.400 ;
        RECT 241.950 459.450 248.550 460.500 ;
        RECT 241.950 458.700 243.750 459.450 ;
        RECT 246.750 458.700 248.550 459.450 ;
        RECT 251.250 458.400 256.050 460.500 ;
        RECT 234.150 456.600 236.850 458.400 ;
        RECT 237.750 457.800 239.550 458.400 ;
        RECT 237.750 456.900 244.050 457.800 ;
        RECT 251.250 457.500 252.450 458.400 ;
        RECT 237.750 456.600 239.550 456.900 ;
        RECT 235.950 455.700 236.850 456.600 ;
        RECT 227.550 448.050 228.750 455.400 ;
        RECT 232.950 454.800 235.050 455.700 ;
        RECT 235.950 454.800 241.050 455.700 ;
        RECT 230.850 453.600 235.050 454.800 ;
        RECT 229.950 451.800 231.750 453.600 ;
        RECT 175.950 445.950 178.200 448.050 ;
        RECT 193.950 445.950 196.050 448.050 ;
        RECT 196.950 445.950 199.050 448.050 ;
        RECT 199.950 445.950 202.050 448.050 ;
        RECT 202.950 445.950 205.050 448.050 ;
        RECT 214.950 445.950 217.050 448.050 ;
        RECT 217.950 445.950 220.050 448.050 ;
        RECT 220.950 445.950 223.050 448.050 ;
        RECT 227.550 447.750 232.050 448.050 ;
        RECT 227.550 445.950 233.850 447.750 ;
        RECT 174.150 440.400 176.100 441.300 ;
        RECT 154.800 432.600 156.600 435.600 ;
        RECT 170.400 439.500 176.100 440.400 ;
        RECT 170.400 435.600 171.600 439.500 ;
        RECT 177.000 438.600 178.200 445.950 ;
        RECT 194.100 444.150 195.900 445.950 ;
        RECT 196.950 441.750 198.150 445.950 ;
        RECT 200.100 444.150 201.900 445.950 ;
        RECT 215.100 444.150 216.900 445.950 ;
        RECT 194.400 440.700 198.150 441.750 ;
        RECT 218.400 440.700 219.600 445.950 ;
        RECT 221.100 444.150 222.900 445.950 ;
        RECT 194.400 438.600 195.600 440.700 ;
        RECT 218.400 439.800 222.600 440.700 ;
        RECT 170.400 432.600 172.200 435.600 ;
        RECT 176.400 432.600 178.200 438.600 ;
        RECT 193.800 432.600 195.600 438.600 ;
        RECT 196.800 437.700 204.600 439.050 ;
        RECT 196.800 432.600 198.600 437.700 ;
        RECT 202.800 432.600 204.600 437.700 ;
        RECT 220.800 432.600 222.600 439.800 ;
        RECT 227.550 438.600 228.750 445.950 ;
        RECT 240.150 442.200 241.050 454.800 ;
        RECT 243.150 454.800 244.050 456.900 ;
        RECT 244.950 456.300 252.450 457.500 ;
        RECT 244.950 455.700 246.750 456.300 ;
        RECT 259.050 455.400 260.850 467.400 ;
        RECT 243.150 454.500 251.550 454.800 ;
        RECT 259.950 454.500 260.850 455.400 ;
        RECT 243.150 453.900 260.850 454.500 ;
        RECT 249.750 453.300 260.850 453.900 ;
        RECT 249.750 453.000 251.550 453.300 ;
        RECT 247.950 446.400 250.050 448.050 ;
        RECT 247.950 445.200 255.900 446.400 ;
        RECT 256.950 445.950 259.050 448.050 ;
        RECT 254.100 444.600 255.900 445.200 ;
        RECT 257.100 444.150 258.900 445.950 ;
        RECT 251.100 443.400 252.900 444.000 ;
        RECT 257.100 443.400 258.000 444.150 ;
        RECT 251.100 442.200 258.000 443.400 ;
        RECT 240.150 441.000 252.150 442.200 ;
        RECT 240.150 440.400 241.950 441.000 ;
        RECT 251.100 439.200 252.150 441.000 ;
        RECT 227.550 432.600 229.350 438.600 ;
        RECT 232.950 437.700 235.050 438.600 ;
        RECT 232.950 436.500 236.700 437.700 ;
        RECT 247.350 437.550 249.150 438.300 ;
        RECT 235.650 435.600 236.700 436.500 ;
        RECT 244.200 436.500 249.150 437.550 ;
        RECT 250.650 437.400 252.450 439.200 ;
        RECT 259.950 438.600 260.850 453.300 ;
        RECT 275.400 461.400 277.200 467.400 ;
        RECT 275.400 448.050 276.600 461.400 ;
        RECT 284.550 455.400 286.350 467.400 ;
        RECT 292.050 461.400 293.850 467.400 ;
        RECT 289.950 459.300 293.850 461.400 ;
        RECT 299.850 460.500 301.650 467.400 ;
        RECT 307.650 461.400 309.450 467.400 ;
        RECT 308.250 460.500 309.450 461.400 ;
        RECT 298.950 459.450 305.550 460.500 ;
        RECT 298.950 458.700 300.750 459.450 ;
        RECT 303.750 458.700 305.550 459.450 ;
        RECT 308.250 458.400 313.050 460.500 ;
        RECT 291.150 456.600 293.850 458.400 ;
        RECT 294.750 457.800 296.550 458.400 ;
        RECT 294.750 456.900 301.050 457.800 ;
        RECT 308.250 457.500 309.450 458.400 ;
        RECT 294.750 456.600 296.550 456.900 ;
        RECT 292.950 455.700 293.850 456.600 ;
        RECT 284.550 448.050 285.750 455.400 ;
        RECT 289.950 454.800 292.050 455.700 ;
        RECT 292.950 454.800 298.050 455.700 ;
        RECT 287.850 453.600 292.050 454.800 ;
        RECT 286.950 451.800 288.750 453.600 ;
        RECT 271.950 445.950 274.050 448.050 ;
        RECT 274.950 445.950 277.050 448.050 ;
        RECT 277.950 445.950 280.050 448.050 ;
        RECT 284.550 447.750 289.050 448.050 ;
        RECT 284.550 445.950 290.850 447.750 ;
        RECT 272.100 444.150 273.900 445.950 ;
        RECT 275.400 440.700 276.600 445.950 ;
        RECT 278.100 444.150 279.900 445.950 ;
        RECT 275.400 439.800 279.600 440.700 ;
        RECT 253.950 436.500 256.050 438.600 ;
        RECT 244.200 435.600 245.250 436.500 ;
        RECT 253.950 435.600 255.000 436.500 ;
        RECT 235.650 432.600 237.450 435.600 ;
        RECT 243.450 432.600 245.250 435.600 ;
        RECT 251.250 434.700 255.000 435.600 ;
        RECT 251.250 432.600 253.050 434.700 ;
        RECT 259.050 432.600 260.850 438.600 ;
        RECT 277.800 432.600 279.600 439.800 ;
        RECT 284.550 438.600 285.750 445.950 ;
        RECT 297.150 442.200 298.050 454.800 ;
        RECT 300.150 454.800 301.050 456.900 ;
        RECT 301.950 456.300 309.450 457.500 ;
        RECT 301.950 455.700 303.750 456.300 ;
        RECT 316.050 455.400 317.850 467.400 ;
        RECT 335.400 461.400 337.200 467.400 ;
        RECT 359.400 461.400 361.200 467.400 ;
        RECT 300.150 454.500 308.550 454.800 ;
        RECT 316.950 454.500 317.850 455.400 ;
        RECT 300.150 453.900 317.850 454.500 ;
        RECT 306.750 453.300 317.850 453.900 ;
        RECT 306.750 453.000 308.550 453.300 ;
        RECT 304.950 446.400 307.050 448.050 ;
        RECT 304.950 445.200 312.900 446.400 ;
        RECT 313.950 445.950 316.050 448.050 ;
        RECT 311.100 444.600 312.900 445.200 ;
        RECT 314.100 444.150 315.900 445.950 ;
        RECT 308.100 443.400 309.900 444.000 ;
        RECT 314.100 443.400 315.000 444.150 ;
        RECT 308.100 442.200 315.000 443.400 ;
        RECT 297.150 441.000 309.150 442.200 ;
        RECT 297.150 440.400 298.950 441.000 ;
        RECT 308.100 439.200 309.150 441.000 ;
        RECT 284.550 432.600 286.350 438.600 ;
        RECT 289.950 437.700 292.050 438.600 ;
        RECT 289.950 436.500 293.700 437.700 ;
        RECT 304.350 437.550 306.150 438.300 ;
        RECT 292.650 435.600 293.700 436.500 ;
        RECT 301.200 436.500 306.150 437.550 ;
        RECT 307.650 437.400 309.450 439.200 ;
        RECT 316.950 438.600 317.850 453.300 ;
        RECT 335.850 448.050 337.050 461.400 ;
        RECT 341.100 448.050 342.900 449.850 ;
        RECT 359.850 448.050 361.050 461.400 ;
        RECT 380.700 456.600 382.500 467.400 ;
        RECT 380.700 455.400 384.300 456.600 ;
        RECT 365.100 448.050 366.900 449.850 ;
        RECT 380.100 448.050 381.900 449.850 ;
        RECT 383.400 448.050 384.300 455.400 ;
        RECT 389.550 455.400 391.350 467.400 ;
        RECT 397.050 461.400 398.850 467.400 ;
        RECT 394.950 459.300 398.850 461.400 ;
        RECT 404.850 460.500 406.650 467.400 ;
        RECT 412.650 461.400 414.450 467.400 ;
        RECT 413.250 460.500 414.450 461.400 ;
        RECT 403.950 459.450 410.550 460.500 ;
        RECT 403.950 458.700 405.750 459.450 ;
        RECT 408.750 458.700 410.550 459.450 ;
        RECT 413.250 458.400 418.050 460.500 ;
        RECT 396.150 456.600 398.850 458.400 ;
        RECT 399.750 457.800 401.550 458.400 ;
        RECT 399.750 456.900 406.050 457.800 ;
        RECT 413.250 457.500 414.450 458.400 ;
        RECT 399.750 456.600 401.550 456.900 ;
        RECT 397.950 455.700 398.850 456.600 ;
        RECT 386.100 448.050 387.900 449.850 ;
        RECT 389.550 448.050 390.750 455.400 ;
        RECT 394.950 454.800 397.050 455.700 ;
        RECT 397.950 454.800 403.050 455.700 ;
        RECT 392.850 453.600 397.050 454.800 ;
        RECT 391.950 451.800 393.750 453.600 ;
        RECT 331.950 445.950 334.050 448.050 ;
        RECT 334.950 445.950 337.050 448.050 ;
        RECT 337.950 445.950 340.050 448.050 ;
        RECT 340.950 445.950 343.050 448.050 ;
        RECT 355.950 445.950 358.050 448.050 ;
        RECT 358.950 445.950 361.050 448.050 ;
        RECT 361.950 445.950 364.050 448.050 ;
        RECT 364.950 445.950 367.050 448.050 ;
        RECT 379.950 445.950 382.050 448.050 ;
        RECT 382.950 445.950 385.050 448.050 ;
        RECT 385.950 445.950 388.050 448.050 ;
        RECT 389.550 447.750 394.050 448.050 ;
        RECT 389.550 445.950 395.850 447.750 ;
        RECT 332.100 444.150 333.900 445.950 ;
        RECT 334.950 441.750 336.150 445.950 ;
        RECT 338.100 444.150 339.900 445.950 ;
        RECT 356.100 444.150 357.900 445.950 ;
        RECT 358.950 441.750 360.150 445.950 ;
        RECT 362.100 444.150 363.900 445.950 ;
        RECT 332.400 440.700 336.150 441.750 ;
        RECT 356.400 440.700 360.150 441.750 ;
        RECT 332.400 438.600 333.600 440.700 ;
        RECT 310.950 436.500 313.050 438.600 ;
        RECT 301.200 435.600 302.250 436.500 ;
        RECT 310.950 435.600 312.000 436.500 ;
        RECT 292.650 432.600 294.450 435.600 ;
        RECT 300.450 432.600 302.250 435.600 ;
        RECT 308.250 434.700 312.000 435.600 ;
        RECT 308.250 432.600 310.050 434.700 ;
        RECT 316.050 432.600 317.850 438.600 ;
        RECT 331.800 432.600 333.600 438.600 ;
        RECT 334.800 437.700 342.600 439.050 ;
        RECT 356.400 438.600 357.600 440.700 ;
        RECT 334.800 432.600 336.600 437.700 ;
        RECT 340.800 432.600 342.600 437.700 ;
        RECT 355.800 432.600 357.600 438.600 ;
        RECT 358.800 437.700 366.600 439.050 ;
        RECT 358.800 432.600 360.600 437.700 ;
        RECT 364.800 432.600 366.600 437.700 ;
        RECT 383.400 435.600 384.300 445.950 ;
        RECT 389.550 438.600 390.750 445.950 ;
        RECT 402.150 442.200 403.050 454.800 ;
        RECT 405.150 454.800 406.050 456.900 ;
        RECT 406.950 456.300 414.450 457.500 ;
        RECT 406.950 455.700 408.750 456.300 ;
        RECT 421.050 455.400 422.850 467.400 ;
        RECT 405.150 454.500 413.550 454.800 ;
        RECT 421.950 454.500 422.850 455.400 ;
        RECT 405.150 453.900 422.850 454.500 ;
        RECT 411.750 453.300 422.850 453.900 ;
        RECT 411.750 453.000 413.550 453.300 ;
        RECT 409.950 446.400 412.050 448.050 ;
        RECT 409.950 445.200 417.900 446.400 ;
        RECT 418.950 445.950 421.050 448.050 ;
        RECT 416.100 444.600 417.900 445.200 ;
        RECT 419.100 444.150 420.900 445.950 ;
        RECT 413.100 443.400 414.900 444.000 ;
        RECT 419.100 443.400 420.000 444.150 ;
        RECT 413.100 442.200 420.000 443.400 ;
        RECT 402.150 441.000 414.150 442.200 ;
        RECT 402.150 440.400 403.950 441.000 ;
        RECT 413.100 439.200 414.150 441.000 ;
        RECT 382.800 432.600 384.600 435.600 ;
        RECT 389.550 432.600 391.350 438.600 ;
        RECT 394.950 437.700 397.050 438.600 ;
        RECT 394.950 436.500 398.700 437.700 ;
        RECT 409.350 437.550 411.150 438.300 ;
        RECT 397.650 435.600 398.700 436.500 ;
        RECT 406.200 436.500 411.150 437.550 ;
        RECT 412.650 437.400 414.450 439.200 ;
        RECT 421.950 438.600 422.850 453.300 ;
        RECT 415.950 436.500 418.050 438.600 ;
        RECT 406.200 435.600 407.250 436.500 ;
        RECT 415.950 435.600 417.000 436.500 ;
        RECT 397.650 432.600 399.450 435.600 ;
        RECT 405.450 432.600 407.250 435.600 ;
        RECT 413.250 434.700 417.000 435.600 ;
        RECT 413.250 432.600 415.050 434.700 ;
        RECT 421.050 432.600 422.850 438.600 ;
        RECT 436.800 455.400 438.600 467.400 ;
        RECT 442.800 461.400 444.600 467.400 ;
        RECT 436.800 448.050 438.000 455.400 ;
        RECT 443.400 454.500 444.600 461.400 ;
        RECT 438.900 453.600 444.600 454.500 ;
        RECT 446.550 455.400 448.350 467.400 ;
        RECT 454.050 461.400 455.850 467.400 ;
        RECT 451.950 459.300 455.850 461.400 ;
        RECT 461.850 460.500 463.650 467.400 ;
        RECT 469.650 461.400 471.450 467.400 ;
        RECT 470.250 460.500 471.450 461.400 ;
        RECT 460.950 459.450 467.550 460.500 ;
        RECT 460.950 458.700 462.750 459.450 ;
        RECT 465.750 458.700 467.550 459.450 ;
        RECT 470.250 458.400 475.050 460.500 ;
        RECT 453.150 456.600 455.850 458.400 ;
        RECT 456.750 457.800 458.550 458.400 ;
        RECT 456.750 456.900 463.050 457.800 ;
        RECT 470.250 457.500 471.450 458.400 ;
        RECT 456.750 456.600 458.550 456.900 ;
        RECT 454.950 455.700 455.850 456.600 ;
        RECT 438.900 452.700 440.850 453.600 ;
        RECT 436.800 445.950 439.050 448.050 ;
        RECT 436.800 438.600 438.000 445.950 ;
        RECT 439.950 441.300 440.850 452.700 ;
        RECT 443.100 448.050 444.900 449.850 ;
        RECT 446.550 448.050 447.750 455.400 ;
        RECT 451.950 454.800 454.050 455.700 ;
        RECT 454.950 454.800 460.050 455.700 ;
        RECT 449.850 453.600 454.050 454.800 ;
        RECT 448.950 451.800 450.750 453.600 ;
        RECT 442.950 445.950 445.050 448.050 ;
        RECT 446.550 447.750 451.050 448.050 ;
        RECT 446.550 445.950 452.850 447.750 ;
        RECT 438.900 440.400 440.850 441.300 ;
        RECT 438.900 439.500 444.600 440.400 ;
        RECT 436.800 432.600 438.600 438.600 ;
        RECT 443.400 435.600 444.600 439.500 ;
        RECT 442.800 432.600 444.600 435.600 ;
        RECT 446.550 438.600 447.750 445.950 ;
        RECT 459.150 442.200 460.050 454.800 ;
        RECT 462.150 454.800 463.050 456.900 ;
        RECT 463.950 456.300 471.450 457.500 ;
        RECT 463.950 455.700 465.750 456.300 ;
        RECT 478.050 455.400 479.850 467.400 ;
        RECT 462.150 454.500 470.550 454.800 ;
        RECT 478.950 454.500 479.850 455.400 ;
        RECT 462.150 453.900 479.850 454.500 ;
        RECT 468.750 453.300 479.850 453.900 ;
        RECT 491.400 461.400 493.200 467.400 ;
        RECT 491.400 454.500 492.600 461.400 ;
        RECT 497.400 455.400 499.200 467.400 ;
        RECT 491.400 453.600 497.100 454.500 ;
        RECT 468.750 453.000 470.550 453.300 ;
        RECT 466.950 446.400 469.050 448.050 ;
        RECT 466.950 445.200 474.900 446.400 ;
        RECT 475.950 445.950 478.050 448.050 ;
        RECT 473.100 444.600 474.900 445.200 ;
        RECT 476.100 444.150 477.900 445.950 ;
        RECT 470.100 443.400 471.900 444.000 ;
        RECT 476.100 443.400 477.000 444.150 ;
        RECT 470.100 442.200 477.000 443.400 ;
        RECT 459.150 441.000 471.150 442.200 ;
        RECT 459.150 440.400 460.950 441.000 ;
        RECT 470.100 439.200 471.150 441.000 ;
        RECT 446.550 432.600 448.350 438.600 ;
        RECT 451.950 437.700 454.050 438.600 ;
        RECT 451.950 436.500 455.700 437.700 ;
        RECT 466.350 437.550 468.150 438.300 ;
        RECT 454.650 435.600 455.700 436.500 ;
        RECT 463.200 436.500 468.150 437.550 ;
        RECT 469.650 437.400 471.450 439.200 ;
        RECT 478.950 438.600 479.850 453.300 ;
        RECT 495.150 452.700 497.100 453.600 ;
        RECT 491.100 448.050 492.900 449.850 ;
        RECT 490.950 445.950 493.050 448.050 ;
        RECT 495.150 441.300 496.050 452.700 ;
        RECT 498.000 448.050 499.200 455.400 ;
        RECT 515.400 455.400 517.200 467.400 ;
        RECT 535.800 461.400 537.600 467.400 ;
        RECT 515.400 448.050 516.600 455.400 ;
        RECT 536.400 448.050 537.600 461.400 ;
        RECT 556.800 455.400 558.600 467.400 ;
        RECT 574.800 455.400 576.600 467.400 ;
        RECT 557.400 448.050 558.600 455.400 ;
        RECT 575.400 448.050 576.600 455.400 ;
        RECT 593.400 461.400 595.200 467.400 ;
        RECT 593.400 448.050 594.600 461.400 ;
        RECT 614.700 456.600 616.500 467.400 ;
        RECT 635.400 461.400 637.200 467.400 ;
        RECT 614.700 455.400 618.300 456.600 ;
        RECT 595.950 453.450 598.050 454.200 ;
        RECT 607.950 453.450 610.050 453.900 ;
        RECT 595.950 452.550 610.050 453.450 ;
        RECT 595.950 452.100 598.050 452.550 ;
        RECT 607.950 451.800 610.050 452.550 ;
        RECT 614.100 448.050 615.900 449.850 ;
        RECT 617.400 448.050 618.300 455.400 ;
        RECT 620.100 448.050 621.900 449.850 ;
        RECT 496.950 445.950 499.200 448.050 ;
        RECT 511.950 445.950 514.050 448.050 ;
        RECT 514.950 445.950 517.050 448.050 ;
        RECT 532.950 445.950 535.050 448.050 ;
        RECT 535.950 445.950 538.050 448.050 ;
        RECT 538.950 445.950 541.050 448.050 ;
        RECT 556.950 445.950 559.050 448.050 ;
        RECT 559.950 445.950 562.050 448.050 ;
        RECT 574.950 445.950 577.050 448.050 ;
        RECT 577.950 445.950 580.050 448.050 ;
        RECT 589.950 445.950 592.050 448.050 ;
        RECT 592.950 445.950 595.050 448.050 ;
        RECT 595.950 445.950 598.050 448.050 ;
        RECT 613.950 445.950 616.050 448.050 ;
        RECT 616.950 445.950 619.050 448.050 ;
        RECT 619.950 445.950 622.050 448.050 ;
        RECT 631.950 445.950 634.050 448.050 ;
        RECT 495.150 440.400 497.100 441.300 ;
        RECT 472.950 436.500 475.050 438.600 ;
        RECT 463.200 435.600 464.250 436.500 ;
        RECT 472.950 435.600 474.000 436.500 ;
        RECT 454.650 432.600 456.450 435.600 ;
        RECT 462.450 432.600 464.250 435.600 ;
        RECT 470.250 434.700 474.000 435.600 ;
        RECT 470.250 432.600 472.050 434.700 ;
        RECT 478.050 432.600 479.850 438.600 ;
        RECT 491.400 439.500 497.100 440.400 ;
        RECT 491.400 435.600 492.600 439.500 ;
        RECT 498.000 438.600 499.200 445.950 ;
        RECT 512.100 444.150 513.900 445.950 ;
        RECT 491.400 432.600 493.200 435.600 ;
        RECT 497.400 432.600 499.200 438.600 ;
        RECT 515.400 438.600 516.600 445.950 ;
        RECT 533.100 444.150 534.900 445.950 ;
        RECT 536.400 440.700 537.600 445.950 ;
        RECT 539.100 444.150 540.900 445.950 ;
        RECT 533.400 439.800 537.600 440.700 ;
        RECT 515.400 432.600 517.200 438.600 ;
        RECT 533.400 432.600 535.200 439.800 ;
        RECT 557.400 438.600 558.600 445.950 ;
        RECT 560.100 444.150 561.900 445.950 ;
        RECT 575.400 438.600 576.600 445.950 ;
        RECT 578.100 444.150 579.900 445.950 ;
        RECT 590.100 444.150 591.900 445.950 ;
        RECT 593.400 440.700 594.600 445.950 ;
        RECT 596.100 444.150 597.900 445.950 ;
        RECT 593.400 439.800 597.600 440.700 ;
        RECT 556.800 432.600 558.600 438.600 ;
        RECT 574.800 432.600 576.600 438.600 ;
        RECT 595.800 432.600 597.600 439.800 ;
        RECT 617.400 435.600 618.300 445.950 ;
        RECT 632.100 444.150 633.900 445.950 ;
        RECT 635.400 441.300 636.300 461.400 ;
        RECT 641.400 455.400 643.200 467.400 ;
        RECT 658.800 466.500 666.600 467.400 ;
        RECT 658.800 455.400 660.600 466.500 ;
        RECT 638.100 448.050 639.900 449.850 ;
        RECT 641.700 448.050 642.600 455.400 ;
        RECT 661.800 454.500 663.600 465.600 ;
        RECT 664.800 456.600 666.600 466.500 ;
        RECT 670.800 456.600 672.600 467.400 ;
        RECT 688.800 461.400 690.600 467.400 ;
        RECT 709.800 461.400 711.600 467.400 ;
        RECT 731.400 461.400 733.200 467.400 ;
        RECT 754.800 461.400 756.600 467.400 ;
        RECT 775.800 461.400 777.600 467.400 ;
        RECT 664.800 455.700 672.600 456.600 ;
        RECT 661.800 453.600 666.900 454.500 ;
        RECT 662.100 448.050 663.900 449.850 ;
        RECT 666.000 448.050 666.900 453.600 ;
        RECT 668.100 448.050 669.900 449.850 ;
        RECT 689.400 448.050 690.600 461.400 ;
        RECT 704.100 448.050 705.900 449.850 ;
        RECT 709.950 448.050 711.150 461.400 ;
        RECT 731.400 448.050 732.600 461.400 ;
        RECT 755.400 448.050 756.600 461.400 ;
        RECT 776.400 448.050 777.600 461.400 ;
        RECT 793.800 456.600 795.600 467.400 ;
        RECT 793.800 455.400 798.600 456.600 ;
        RECT 796.500 454.500 798.600 455.400 ;
        RECT 801.300 455.400 803.100 467.400 ;
        RECT 808.800 456.300 810.600 467.400 ;
        RECT 826.800 461.400 828.600 467.400 ;
        RECT 847.800 461.400 849.600 467.400 ;
        RECT 806.100 455.400 810.600 456.300 ;
        RECT 786.000 453.450 790.050 454.050 ;
        RECT 801.300 453.900 802.500 455.400 ;
        RECT 785.550 451.950 790.050 453.450 ;
        RECT 801.000 453.000 802.500 453.900 ;
        RECT 806.100 453.300 808.200 455.400 ;
        RECT 637.950 445.950 640.050 448.050 ;
        RECT 640.950 445.950 643.050 448.050 ;
        RECT 658.950 445.950 661.050 448.050 ;
        RECT 661.950 445.950 664.050 448.050 ;
        RECT 664.950 445.950 667.050 448.050 ;
        RECT 667.950 445.950 670.050 448.050 ;
        RECT 670.950 445.950 673.050 448.050 ;
        RECT 685.950 445.950 688.050 448.050 ;
        RECT 688.950 445.950 691.050 448.050 ;
        RECT 691.950 445.950 694.050 448.050 ;
        RECT 703.950 445.950 706.050 448.050 ;
        RECT 706.950 445.950 709.050 448.050 ;
        RECT 709.950 445.950 712.050 448.050 ;
        RECT 712.950 445.950 715.050 448.050 ;
        RECT 727.950 445.950 730.050 448.050 ;
        RECT 730.950 445.950 733.050 448.050 ;
        RECT 733.950 445.950 736.050 448.050 ;
        RECT 751.950 445.950 754.050 448.050 ;
        RECT 754.950 445.950 757.050 448.050 ;
        RECT 757.950 445.950 760.050 448.050 ;
        RECT 772.950 445.950 775.050 448.050 ;
        RECT 775.950 445.950 778.050 448.050 ;
        RECT 778.950 445.950 781.050 448.050 ;
        RECT 632.400 440.400 639.900 441.300 ;
        RECT 616.800 432.600 618.600 435.600 ;
        RECT 632.400 432.600 634.200 440.400 ;
        RECT 638.100 439.500 639.900 440.400 ;
        RECT 641.700 438.600 642.600 445.950 ;
        RECT 659.100 444.150 660.900 445.950 ;
        RECT 639.900 436.800 642.600 438.600 ;
        RECT 666.000 438.600 667.050 445.950 ;
        RECT 671.100 444.150 672.900 445.950 ;
        RECT 686.100 444.150 687.900 445.950 ;
        RECT 689.400 440.700 690.600 445.950 ;
        RECT 692.100 444.150 693.900 445.950 ;
        RECT 707.100 444.150 708.900 445.950 ;
        RECT 710.850 441.750 712.050 445.950 ;
        RECT 713.100 444.150 714.900 445.950 ;
        RECT 728.100 444.150 729.900 445.950 ;
        RECT 710.850 440.700 714.600 441.750 ;
        RECT 686.400 439.800 690.600 440.700 ;
        RECT 639.900 432.600 641.700 436.800 ;
        RECT 666.000 432.600 667.800 438.600 ;
        RECT 686.400 432.600 688.200 439.800 ;
        RECT 704.400 437.700 712.200 439.050 ;
        RECT 704.400 432.600 706.200 437.700 ;
        RECT 710.400 432.600 712.200 437.700 ;
        RECT 713.400 438.600 714.600 440.700 ;
        RECT 731.400 440.700 732.600 445.950 ;
        RECT 734.100 444.150 735.900 445.950 ;
        RECT 752.100 444.150 753.900 445.950 ;
        RECT 755.400 440.700 756.600 445.950 ;
        RECT 758.100 444.150 759.900 445.950 ;
        RECT 773.100 444.150 774.900 445.950 ;
        RECT 776.400 440.700 777.600 445.950 ;
        RECT 779.100 444.150 780.900 445.950 ;
        RECT 785.550 444.450 786.450 451.950 ;
        RECT 801.000 450.900 801.900 453.000 ;
        RECT 794.100 448.050 795.900 449.850 ;
        RECT 799.800 448.800 801.900 450.900 ;
        RECT 802.800 451.500 804.900 451.800 ;
        RECT 802.800 449.700 806.700 451.500 ;
        RECT 787.950 447.450 792.000 448.050 ;
        RECT 793.950 447.450 796.050 448.050 ;
        RECT 800.400 447.900 802.800 448.800 ;
        RECT 787.950 446.550 796.050 447.450 ;
        RECT 787.950 445.950 792.000 446.550 ;
        RECT 793.950 445.950 796.050 446.550 ;
        RECT 798.600 445.200 800.400 447.000 ;
        RECT 782.550 443.550 786.450 444.450 ;
        RECT 782.550 442.050 783.450 443.550 ;
        RECT 798.750 443.100 800.850 445.200 ;
        RECT 801.750 442.200 802.800 447.900 ;
        RECT 803.700 447.900 805.500 448.500 ;
        RECT 821.100 448.050 822.900 449.850 ;
        RECT 826.950 448.050 828.150 461.400 ;
        RECT 832.950 450.450 835.050 451.050 ;
        RECT 841.950 450.450 844.050 451.050 ;
        RECT 832.950 449.550 844.050 450.450 ;
        RECT 832.950 448.950 835.050 449.550 ;
        RECT 841.950 448.950 844.050 449.550 ;
        RECT 848.400 448.050 849.600 461.400 ;
        RECT 866.400 461.400 868.200 467.400 ;
        RECT 850.950 459.450 853.050 460.050 ;
        RECT 856.950 459.450 859.050 460.050 ;
        RECT 850.950 458.550 859.050 459.450 ;
        RECT 850.950 457.950 853.050 458.550 ;
        RECT 856.950 457.950 859.050 458.550 ;
        RECT 853.950 450.450 858.000 451.050 ;
        RECT 851.100 448.050 852.900 449.850 ;
        RECT 853.950 448.950 858.450 450.450 ;
        RECT 808.500 447.900 810.600 448.050 ;
        RECT 803.700 446.700 810.600 447.900 ;
        RECT 808.500 445.950 810.600 446.700 ;
        RECT 820.950 445.950 823.050 448.050 ;
        RECT 823.950 445.950 826.050 448.050 ;
        RECT 826.950 445.950 829.050 448.050 ;
        RECT 829.950 445.950 832.050 448.050 ;
        RECT 847.950 445.950 850.050 448.050 ;
        RECT 850.950 445.950 853.050 448.050 ;
        RECT 731.400 439.800 735.600 440.700 ;
        RECT 713.400 432.600 715.200 438.600 ;
        RECT 733.800 432.600 735.600 439.800 ;
        RECT 752.400 439.800 756.600 440.700 ;
        RECT 773.400 439.800 777.600 440.700 ;
        RECT 778.950 440.550 783.450 442.050 ;
        RECT 778.950 439.950 783.000 440.550 ;
        RECT 752.400 432.600 754.200 439.800 ;
        RECT 773.400 432.600 775.200 439.800 ;
        RECT 796.500 439.500 798.600 440.700 ;
        RECT 799.800 440.100 802.800 442.200 ;
        RECT 803.700 443.400 805.500 445.200 ;
        RECT 808.800 444.450 810.600 445.950 ;
        RECT 814.950 444.450 817.050 445.050 ;
        RECT 808.800 444.150 817.050 444.450 ;
        RECT 824.100 444.150 825.900 445.950 ;
        RECT 809.550 443.550 817.050 444.150 ;
        RECT 803.700 441.300 805.800 443.400 ;
        RECT 814.950 442.950 817.050 443.550 ;
        RECT 827.850 441.750 829.050 445.950 ;
        RECT 830.100 444.150 831.900 445.950 ;
        RECT 803.700 440.400 810.000 441.300 ;
        RECT 827.850 440.700 831.600 441.750 ;
        RECT 793.800 438.600 798.600 439.500 ;
        RECT 801.600 438.600 802.800 440.100 ;
        RECT 808.800 438.600 810.000 440.400 ;
        RECT 793.800 432.600 795.600 438.600 ;
        RECT 801.300 432.600 803.100 438.600 ;
        RECT 808.800 432.600 810.600 438.600 ;
        RECT 821.400 437.700 829.200 439.050 ;
        RECT 821.400 432.600 823.200 437.700 ;
        RECT 827.400 432.600 829.200 437.700 ;
        RECT 830.400 438.600 831.600 440.700 ;
        RECT 830.400 432.600 832.200 438.600 ;
        RECT 848.400 435.600 849.600 445.950 ;
        RECT 857.550 444.450 858.450 448.950 ;
        RECT 863.100 448.050 864.900 449.850 ;
        RECT 866.400 448.050 867.600 461.400 ;
        RECT 881.400 456.300 883.200 467.400 ;
        RECT 887.400 456.300 889.200 467.400 ;
        RECT 881.400 455.400 889.200 456.300 ;
        RECT 890.400 455.400 892.200 467.400 ;
        RECT 883.950 453.450 886.050 454.050 ;
        RECT 875.550 452.550 886.050 453.450 ;
        RECT 862.950 445.950 865.050 448.050 ;
        RECT 865.950 445.950 868.050 448.050 ;
        RECT 857.550 443.550 861.450 444.450 ;
        RECT 860.550 442.050 861.450 443.550 ;
        RECT 860.550 440.550 865.050 442.050 ;
        RECT 861.000 439.950 865.050 440.550 ;
        RECT 847.800 432.600 849.600 435.600 ;
        RECT 866.400 435.600 867.600 445.950 ;
        RECT 875.550 444.450 876.450 452.550 ;
        RECT 883.950 451.950 886.050 452.550 ;
        RECT 884.100 448.050 885.900 449.850 ;
        RECT 890.700 448.050 891.600 455.400 ;
        RECT 880.950 445.950 883.050 448.050 ;
        RECT 883.950 445.950 886.050 448.050 ;
        RECT 886.950 445.950 889.050 448.050 ;
        RECT 889.950 445.950 892.050 448.050 ;
        RECT 875.550 443.550 879.450 444.450 ;
        RECT 881.100 444.150 882.900 445.950 ;
        RECT 887.100 444.150 888.900 445.950 ;
        RECT 878.550 441.450 879.450 443.550 ;
        RECT 886.950 441.450 889.050 442.050 ;
        RECT 878.550 440.550 889.050 441.450 ;
        RECT 886.950 439.950 889.050 440.550 ;
        RECT 890.700 438.600 891.600 445.950 ;
        RECT 886.500 437.400 891.600 438.600 ;
        RECT 866.400 432.600 868.200 435.600 ;
        RECT 886.500 432.600 888.300 437.400 ;
        RECT 3.150 422.400 4.950 428.400 ;
        RECT 10.950 426.300 12.750 428.400 ;
        RECT 9.000 425.400 12.750 426.300 ;
        RECT 18.750 425.400 20.550 428.400 ;
        RECT 26.550 425.400 28.350 428.400 ;
        RECT 9.000 424.500 10.050 425.400 ;
        RECT 18.750 424.500 19.800 425.400 ;
        RECT 7.950 422.400 10.050 424.500 ;
        RECT 3.150 407.700 4.050 422.400 ;
        RECT 11.550 421.800 13.350 423.600 ;
        RECT 14.850 423.450 19.800 424.500 ;
        RECT 27.300 424.500 28.350 425.400 ;
        RECT 14.850 422.700 16.650 423.450 ;
        RECT 27.300 423.300 31.050 424.500 ;
        RECT 28.950 422.400 31.050 423.300 ;
        RECT 34.650 422.400 36.450 428.400 ;
        RECT 11.850 420.000 12.900 421.800 ;
        RECT 22.050 420.000 23.850 420.600 ;
        RECT 11.850 418.800 23.850 420.000 ;
        RECT 6.000 417.600 12.900 418.800 ;
        RECT 6.000 416.850 6.900 417.600 ;
        RECT 11.100 417.000 12.900 417.600 ;
        RECT 5.100 415.050 6.900 416.850 ;
        RECT 8.100 415.800 9.900 416.400 ;
        RECT 4.950 412.950 7.050 415.050 ;
        RECT 8.100 414.600 16.050 415.800 ;
        RECT 13.950 412.950 16.050 414.600 ;
        RECT 12.450 407.700 14.250 408.000 ;
        RECT 3.150 407.100 14.250 407.700 ;
        RECT 3.150 406.500 20.850 407.100 ;
        RECT 3.150 405.600 4.050 406.500 ;
        RECT 12.450 406.200 20.850 406.500 ;
        RECT 3.150 393.600 4.950 405.600 ;
        RECT 17.250 404.700 19.050 405.300 ;
        RECT 11.550 403.500 19.050 404.700 ;
        RECT 19.950 404.100 20.850 406.200 ;
        RECT 22.950 406.200 23.850 418.800 ;
        RECT 35.250 415.050 36.450 422.400 ;
        RECT 52.800 421.200 54.600 428.400 ;
        RECT 68.400 423.300 70.200 428.400 ;
        RECT 74.400 423.300 76.200 428.400 ;
        RECT 68.400 421.950 76.200 423.300 ;
        RECT 77.400 422.400 79.200 428.400 ;
        RECT 94.800 422.400 96.600 428.400 ;
        RECT 50.400 420.300 54.600 421.200 ;
        RECT 77.400 420.300 78.600 422.400 ;
        RECT 42.000 417.450 46.050 418.050 ;
        RECT 30.150 413.250 36.450 415.050 ;
        RECT 31.950 412.950 36.450 413.250 ;
        RECT 32.250 407.400 34.050 409.200 ;
        RECT 28.950 406.200 33.150 407.400 ;
        RECT 22.950 405.300 28.050 406.200 ;
        RECT 28.950 405.300 31.050 406.200 ;
        RECT 35.250 405.600 36.450 412.950 ;
        RECT 41.550 415.950 46.050 417.450 ;
        RECT 41.550 408.900 42.450 415.950 ;
        RECT 47.100 415.050 48.900 416.850 ;
        RECT 50.400 415.050 51.600 420.300 ;
        RECT 74.850 419.250 78.600 420.300 ;
        RECT 53.100 415.050 54.900 416.850 ;
        RECT 71.100 415.050 72.900 416.850 ;
        RECT 74.850 415.050 76.050 419.250 ;
        RECT 91.950 417.450 94.050 421.050 ;
        RECT 95.400 420.300 96.600 422.400 ;
        RECT 97.800 423.300 99.600 428.400 ;
        RECT 103.800 423.300 105.600 428.400 ;
        RECT 97.800 421.950 105.600 423.300 ;
        RECT 124.800 421.200 126.600 428.400 ;
        RECT 106.950 420.450 109.050 421.050 ;
        RECT 118.950 420.450 121.050 421.050 ;
        RECT 95.400 419.250 99.150 420.300 ;
        RECT 89.550 417.000 94.050 417.450 ;
        RECT 77.100 415.050 78.900 416.850 ;
        RECT 89.550 416.550 93.450 417.000 ;
        RECT 46.950 412.950 49.050 415.050 ;
        RECT 49.950 412.950 52.050 415.050 ;
        RECT 52.950 412.950 55.050 415.050 ;
        RECT 67.950 412.950 70.050 415.050 ;
        RECT 70.950 412.950 73.050 415.050 ;
        RECT 73.950 412.950 76.050 415.050 ;
        RECT 76.950 412.950 79.050 415.050 ;
        RECT 40.950 406.800 43.050 408.900 ;
        RECT 27.150 404.400 28.050 405.300 ;
        RECT 24.450 404.100 26.250 404.400 ;
        RECT 11.550 402.600 12.750 403.500 ;
        RECT 19.950 403.200 26.250 404.100 ;
        RECT 24.450 402.600 26.250 403.200 ;
        RECT 27.150 402.600 29.850 404.400 ;
        RECT 7.950 400.500 12.750 402.600 ;
        RECT 15.450 401.550 17.250 402.300 ;
        RECT 20.250 401.550 22.050 402.300 ;
        RECT 15.450 400.500 22.050 401.550 ;
        RECT 11.550 399.600 12.750 400.500 ;
        RECT 11.550 393.600 13.350 399.600 ;
        RECT 19.350 393.600 21.150 400.500 ;
        RECT 27.150 399.600 31.050 401.700 ;
        RECT 27.150 393.600 28.950 399.600 ;
        RECT 34.650 393.600 36.450 405.600 ;
        RECT 50.400 399.600 51.600 412.950 ;
        RECT 68.100 411.150 69.900 412.950 ;
        RECT 73.950 399.600 75.150 412.950 ;
        RECT 89.550 405.900 90.450 416.550 ;
        RECT 95.100 415.050 96.900 416.850 ;
        RECT 97.950 415.050 99.150 419.250 ;
        RECT 106.950 419.550 121.050 420.450 ;
        RECT 106.950 418.950 109.050 419.550 ;
        RECT 118.950 418.950 121.050 419.550 ;
        RECT 122.400 420.300 126.600 421.200 ;
        RECT 132.150 422.400 133.950 428.400 ;
        RECT 139.950 426.300 141.750 428.400 ;
        RECT 138.000 425.400 141.750 426.300 ;
        RECT 147.750 425.400 149.550 428.400 ;
        RECT 155.550 425.400 157.350 428.400 ;
        RECT 138.000 424.500 139.050 425.400 ;
        RECT 147.750 424.500 148.800 425.400 ;
        RECT 136.950 422.400 139.050 424.500 ;
        RECT 101.100 415.050 102.900 416.850 ;
        RECT 119.100 415.050 120.900 416.850 ;
        RECT 122.400 415.050 123.600 420.300 ;
        RECT 125.100 415.050 126.900 416.850 ;
        RECT 94.950 412.950 97.050 415.050 ;
        RECT 97.950 412.950 100.050 415.050 ;
        RECT 100.950 412.950 103.050 415.050 ;
        RECT 103.950 412.950 106.050 415.050 ;
        RECT 118.950 412.950 121.050 415.050 ;
        RECT 121.950 412.950 124.050 415.050 ;
        RECT 124.950 412.950 127.050 415.050 ;
        RECT 88.950 403.800 91.050 405.900 ;
        RECT 98.850 399.600 100.050 412.950 ;
        RECT 104.100 411.150 105.900 412.950 ;
        RECT 122.400 399.600 123.600 412.950 ;
        RECT 132.150 407.700 133.050 422.400 ;
        RECT 140.550 421.800 142.350 423.600 ;
        RECT 143.850 423.450 148.800 424.500 ;
        RECT 156.300 424.500 157.350 425.400 ;
        RECT 143.850 422.700 145.650 423.450 ;
        RECT 156.300 423.300 160.050 424.500 ;
        RECT 157.950 422.400 160.050 423.300 ;
        RECT 163.650 422.400 165.450 428.400 ;
        RECT 178.800 422.400 180.600 428.400 ;
        RECT 140.850 420.000 141.900 421.800 ;
        RECT 151.050 420.000 152.850 420.600 ;
        RECT 140.850 418.800 152.850 420.000 ;
        RECT 135.000 417.600 141.900 418.800 ;
        RECT 135.000 416.850 135.900 417.600 ;
        RECT 140.100 417.000 141.900 417.600 ;
        RECT 134.100 415.050 135.900 416.850 ;
        RECT 137.100 415.800 138.900 416.400 ;
        RECT 133.950 412.950 136.050 415.050 ;
        RECT 137.100 414.600 145.050 415.800 ;
        RECT 142.950 412.950 145.050 414.600 ;
        RECT 141.450 407.700 143.250 408.000 ;
        RECT 132.150 407.100 143.250 407.700 ;
        RECT 132.150 406.500 149.850 407.100 ;
        RECT 132.150 405.600 133.050 406.500 ;
        RECT 141.450 406.200 149.850 406.500 ;
        RECT 50.400 393.600 52.200 399.600 ;
        RECT 73.800 393.600 75.600 399.600 ;
        RECT 98.400 393.600 100.200 399.600 ;
        RECT 122.400 393.600 124.200 399.600 ;
        RECT 132.150 393.600 133.950 405.600 ;
        RECT 146.250 404.700 148.050 405.300 ;
        RECT 140.550 403.500 148.050 404.700 ;
        RECT 148.950 404.100 149.850 406.200 ;
        RECT 151.950 406.200 152.850 418.800 ;
        RECT 164.250 415.050 165.450 422.400 ;
        RECT 179.400 420.300 180.600 422.400 ;
        RECT 181.800 423.300 183.600 428.400 ;
        RECT 187.800 423.300 189.600 428.400 ;
        RECT 205.800 425.400 207.600 428.400 ;
        RECT 223.800 425.400 225.600 428.400 ;
        RECT 241.800 425.400 243.600 428.400 ;
        RECT 181.800 421.950 189.600 423.300 ;
        RECT 179.400 419.250 183.150 420.300 ;
        RECT 179.100 415.050 180.900 416.850 ;
        RECT 181.950 415.050 183.150 419.250 ;
        RECT 185.100 415.050 186.900 416.850 ;
        RECT 206.400 415.050 207.300 425.400 ;
        RECT 224.400 415.050 225.600 425.400 ;
        RECT 242.400 415.050 243.600 425.400 ;
        RECT 248.550 422.400 250.350 428.400 ;
        RECT 256.650 425.400 258.450 428.400 ;
        RECT 264.450 425.400 266.250 428.400 ;
        RECT 272.250 426.300 274.050 428.400 ;
        RECT 272.250 425.400 276.000 426.300 ;
        RECT 256.650 424.500 257.700 425.400 ;
        RECT 253.950 423.300 257.700 424.500 ;
        RECT 265.200 424.500 266.250 425.400 ;
        RECT 274.950 424.500 276.000 425.400 ;
        RECT 265.200 423.450 270.150 424.500 ;
        RECT 253.950 422.400 256.050 423.300 ;
        RECT 268.350 422.700 270.150 423.450 ;
        RECT 248.550 415.050 249.750 422.400 ;
        RECT 271.650 421.800 273.450 423.600 ;
        RECT 274.950 422.400 277.050 424.500 ;
        RECT 280.050 422.400 281.850 428.400 ;
        RECT 261.150 420.000 262.950 420.600 ;
        RECT 272.100 420.000 273.150 421.800 ;
        RECT 261.150 418.800 273.150 420.000 ;
        RECT 159.150 413.250 165.450 415.050 ;
        RECT 160.950 412.950 165.450 413.250 ;
        RECT 178.950 412.950 181.050 415.050 ;
        RECT 181.950 412.950 184.050 415.050 ;
        RECT 184.950 412.950 187.050 415.050 ;
        RECT 187.950 412.950 190.050 415.050 ;
        RECT 202.950 412.950 205.050 415.050 ;
        RECT 205.950 412.950 208.050 415.050 ;
        RECT 208.950 412.950 211.050 415.050 ;
        RECT 223.950 412.950 226.050 415.050 ;
        RECT 226.950 412.950 229.050 415.050 ;
        RECT 241.950 412.950 244.050 415.050 ;
        RECT 244.950 412.950 247.050 415.050 ;
        RECT 248.550 413.250 254.850 415.050 ;
        RECT 248.550 412.950 253.050 413.250 ;
        RECT 161.250 407.400 163.050 409.200 ;
        RECT 157.950 406.200 162.150 407.400 ;
        RECT 151.950 405.300 157.050 406.200 ;
        RECT 157.950 405.300 160.050 406.200 ;
        RECT 164.250 405.600 165.450 412.950 ;
        RECT 156.150 404.400 157.050 405.300 ;
        RECT 153.450 404.100 155.250 404.400 ;
        RECT 140.550 402.600 141.750 403.500 ;
        RECT 148.950 403.200 155.250 404.100 ;
        RECT 153.450 402.600 155.250 403.200 ;
        RECT 156.150 402.600 158.850 404.400 ;
        RECT 136.950 400.500 141.750 402.600 ;
        RECT 144.450 401.550 146.250 402.300 ;
        RECT 149.250 401.550 151.050 402.300 ;
        RECT 144.450 400.500 151.050 401.550 ;
        RECT 140.550 399.600 141.750 400.500 ;
        RECT 140.550 393.600 142.350 399.600 ;
        RECT 148.350 393.600 150.150 400.500 ;
        RECT 156.150 399.600 160.050 401.700 ;
        RECT 156.150 393.600 157.950 399.600 ;
        RECT 163.650 393.600 165.450 405.600 ;
        RECT 182.850 399.600 184.050 412.950 ;
        RECT 188.100 411.150 189.900 412.950 ;
        RECT 203.100 411.150 204.900 412.950 ;
        RECT 206.400 405.600 207.300 412.950 ;
        RECT 209.100 411.150 210.900 412.950 ;
        RECT 203.700 404.400 207.300 405.600 ;
        RECT 182.400 393.600 184.200 399.600 ;
        RECT 203.700 393.600 205.500 404.400 ;
        RECT 224.400 399.600 225.600 412.950 ;
        RECT 227.100 411.150 228.900 412.950 ;
        RECT 242.400 399.600 243.600 412.950 ;
        RECT 245.100 411.150 246.900 412.950 ;
        RECT 223.800 393.600 225.600 399.600 ;
        RECT 241.800 393.600 243.600 399.600 ;
        RECT 248.550 405.600 249.750 412.950 ;
        RECT 250.950 407.400 252.750 409.200 ;
        RECT 251.850 406.200 256.050 407.400 ;
        RECT 261.150 406.200 262.050 418.800 ;
        RECT 272.100 417.600 279.000 418.800 ;
        RECT 272.100 417.000 273.900 417.600 ;
        RECT 278.100 416.850 279.000 417.600 ;
        RECT 275.100 415.800 276.900 416.400 ;
        RECT 268.950 414.600 276.900 415.800 ;
        RECT 278.100 415.050 279.900 416.850 ;
        RECT 268.950 412.950 271.050 414.600 ;
        RECT 277.950 412.950 280.050 415.050 ;
        RECT 270.750 407.700 272.550 408.000 ;
        RECT 280.950 407.700 281.850 422.400 ;
        RECT 298.800 421.200 300.600 428.400 ;
        RECT 314.400 423.300 316.200 428.400 ;
        RECT 320.400 423.300 322.200 428.400 ;
        RECT 314.400 421.950 322.200 423.300 ;
        RECT 323.400 422.400 325.200 428.400 ;
        RECT 343.800 422.400 345.600 428.400 ;
        RECT 296.400 420.300 300.600 421.200 ;
        RECT 323.400 420.300 324.600 422.400 ;
        RECT 293.100 415.050 294.900 416.850 ;
        RECT 296.400 415.050 297.600 420.300 ;
        RECT 320.850 419.250 324.600 420.300 ;
        RECT 344.400 420.300 345.600 422.400 ;
        RECT 346.800 423.300 348.600 428.400 ;
        RECT 352.800 423.300 354.600 428.400 ;
        RECT 346.800 421.950 354.600 423.300 ;
        RECT 365.400 423.300 367.200 428.400 ;
        RECT 371.400 423.300 373.200 428.400 ;
        RECT 365.400 421.950 373.200 423.300 ;
        RECT 374.400 422.400 376.200 428.400 ;
        RECT 394.500 423.600 396.300 428.400 ;
        RECT 394.500 422.400 399.600 423.600 ;
        RECT 415.800 422.400 417.600 428.400 ;
        RECT 374.400 420.300 375.600 422.400 ;
        RECT 344.400 419.250 348.150 420.300 ;
        RECT 299.100 415.050 300.900 416.850 ;
        RECT 317.100 415.050 318.900 416.850 ;
        RECT 320.850 415.050 322.050 419.250 ;
        RECT 323.100 415.050 324.900 416.850 ;
        RECT 344.100 415.050 345.900 416.850 ;
        RECT 346.950 415.050 348.150 419.250 ;
        RECT 371.850 419.250 375.600 420.300 ;
        RECT 350.100 415.050 351.900 416.850 ;
        RECT 368.100 415.050 369.900 416.850 ;
        RECT 371.850 415.050 373.050 419.250 ;
        RECT 374.100 415.050 375.900 416.850 ;
        RECT 389.100 415.050 390.900 416.850 ;
        RECT 395.100 415.050 396.900 416.850 ;
        RECT 398.700 415.050 399.600 422.400 ;
        RECT 416.400 420.300 417.600 422.400 ;
        RECT 418.800 423.300 420.600 428.400 ;
        RECT 424.800 423.300 426.600 428.400 ;
        RECT 418.800 421.950 426.600 423.300 ;
        RECT 429.150 422.400 430.950 428.400 ;
        RECT 436.950 426.300 438.750 428.400 ;
        RECT 435.000 425.400 438.750 426.300 ;
        RECT 444.750 425.400 446.550 428.400 ;
        RECT 452.550 425.400 454.350 428.400 ;
        RECT 435.000 424.500 436.050 425.400 ;
        RECT 444.750 424.500 445.800 425.400 ;
        RECT 433.950 422.400 436.050 424.500 ;
        RECT 416.400 419.250 420.150 420.300 ;
        RECT 416.100 415.050 417.900 416.850 ;
        RECT 418.950 415.050 420.150 419.250 ;
        RECT 422.100 415.050 423.900 416.850 ;
        RECT 292.950 412.950 295.050 415.050 ;
        RECT 295.950 412.950 298.050 415.050 ;
        RECT 298.950 412.950 301.050 415.050 ;
        RECT 313.950 412.950 316.050 415.050 ;
        RECT 316.950 412.950 319.050 415.050 ;
        RECT 319.950 412.950 322.050 415.050 ;
        RECT 322.950 412.950 325.050 415.050 ;
        RECT 343.950 412.950 346.050 415.050 ;
        RECT 346.950 412.950 349.050 415.050 ;
        RECT 349.950 412.950 352.050 415.050 ;
        RECT 352.950 412.950 355.050 415.050 ;
        RECT 364.950 412.950 367.050 415.050 ;
        RECT 367.950 412.950 370.050 415.050 ;
        RECT 370.950 412.950 373.050 415.050 ;
        RECT 373.950 412.950 376.050 415.050 ;
        RECT 388.950 412.950 391.050 415.050 ;
        RECT 391.950 412.950 394.050 415.050 ;
        RECT 394.950 412.950 397.050 415.050 ;
        RECT 397.950 412.950 400.050 415.050 ;
        RECT 415.950 412.950 418.050 415.050 ;
        RECT 418.950 412.950 421.050 415.050 ;
        RECT 421.950 412.950 424.050 415.050 ;
        RECT 424.950 412.950 427.050 415.050 ;
        RECT 270.750 407.100 281.850 407.700 ;
        RECT 248.550 393.600 250.350 405.600 ;
        RECT 253.950 405.300 256.050 406.200 ;
        RECT 256.950 405.300 262.050 406.200 ;
        RECT 264.150 406.500 281.850 407.100 ;
        RECT 264.150 406.200 272.550 406.500 ;
        RECT 256.950 404.400 257.850 405.300 ;
        RECT 255.150 402.600 257.850 404.400 ;
        RECT 258.750 404.100 260.550 404.400 ;
        RECT 264.150 404.100 265.050 406.200 ;
        RECT 280.950 405.600 281.850 406.500 ;
        RECT 258.750 403.200 265.050 404.100 ;
        RECT 265.950 404.700 267.750 405.300 ;
        RECT 265.950 403.500 273.450 404.700 ;
        RECT 258.750 402.600 260.550 403.200 ;
        RECT 272.250 402.600 273.450 403.500 ;
        RECT 253.950 399.600 257.850 401.700 ;
        RECT 262.950 401.550 264.750 402.300 ;
        RECT 267.750 401.550 269.550 402.300 ;
        RECT 262.950 400.500 269.550 401.550 ;
        RECT 272.250 400.500 277.050 402.600 ;
        RECT 256.050 393.600 257.850 399.600 ;
        RECT 263.850 393.600 265.650 400.500 ;
        RECT 272.250 399.600 273.450 400.500 ;
        RECT 271.650 393.600 273.450 399.600 ;
        RECT 280.050 393.600 281.850 405.600 ;
        RECT 296.400 399.600 297.600 412.950 ;
        RECT 314.100 411.150 315.900 412.950 ;
        RECT 319.950 399.600 321.150 412.950 ;
        RECT 347.850 399.600 349.050 412.950 ;
        RECT 353.100 411.150 354.900 412.950 ;
        RECT 365.100 411.150 366.900 412.950 ;
        RECT 370.950 399.600 372.150 412.950 ;
        RECT 379.950 411.450 382.050 412.050 ;
        RECT 385.950 411.450 388.050 412.050 ;
        RECT 379.950 410.550 388.050 411.450 ;
        RECT 392.100 411.150 393.900 412.950 ;
        RECT 379.950 409.950 382.050 410.550 ;
        RECT 385.950 409.950 388.050 410.550 ;
        RECT 398.700 405.600 399.600 412.950 ;
        RECT 389.400 404.700 397.200 405.600 ;
        RECT 296.400 393.600 298.200 399.600 ;
        RECT 319.800 393.600 321.600 399.600 ;
        RECT 347.400 393.600 349.200 399.600 ;
        RECT 370.800 393.600 372.600 399.600 ;
        RECT 389.400 393.600 391.200 404.700 ;
        RECT 395.400 393.600 397.200 404.700 ;
        RECT 398.400 393.600 400.200 405.600 ;
        RECT 419.850 399.600 421.050 412.950 ;
        RECT 425.100 411.150 426.900 412.950 ;
        RECT 429.150 407.700 430.050 422.400 ;
        RECT 437.550 421.800 439.350 423.600 ;
        RECT 440.850 423.450 445.800 424.500 ;
        RECT 453.300 424.500 454.350 425.400 ;
        RECT 440.850 422.700 442.650 423.450 ;
        RECT 453.300 423.300 457.050 424.500 ;
        RECT 454.950 422.400 457.050 423.300 ;
        RECT 460.650 422.400 462.450 428.400 ;
        RECT 437.850 420.000 438.900 421.800 ;
        RECT 448.050 420.000 449.850 420.600 ;
        RECT 437.850 418.800 449.850 420.000 ;
        RECT 432.000 417.600 438.900 418.800 ;
        RECT 432.000 416.850 432.900 417.600 ;
        RECT 437.100 417.000 438.900 417.600 ;
        RECT 431.100 415.050 432.900 416.850 ;
        RECT 434.100 415.800 435.900 416.400 ;
        RECT 430.950 412.950 433.050 415.050 ;
        RECT 434.100 414.600 442.050 415.800 ;
        RECT 439.950 412.950 442.050 414.600 ;
        RECT 438.450 407.700 440.250 408.000 ;
        RECT 429.150 407.100 440.250 407.700 ;
        RECT 429.150 406.500 446.850 407.100 ;
        RECT 429.150 405.600 430.050 406.500 ;
        RECT 438.450 406.200 446.850 406.500 ;
        RECT 419.400 393.600 421.200 399.600 ;
        RECT 429.150 393.600 430.950 405.600 ;
        RECT 443.250 404.700 445.050 405.300 ;
        RECT 437.550 403.500 445.050 404.700 ;
        RECT 445.950 404.100 446.850 406.200 ;
        RECT 448.950 406.200 449.850 418.800 ;
        RECT 461.250 415.050 462.450 422.400 ;
        RECT 456.150 413.250 462.450 415.050 ;
        RECT 457.950 412.950 462.450 413.250 ;
        RECT 458.250 407.400 460.050 409.200 ;
        RECT 454.950 406.200 459.150 407.400 ;
        RECT 448.950 405.300 454.050 406.200 ;
        RECT 454.950 405.300 457.050 406.200 ;
        RECT 461.250 405.600 462.450 412.950 ;
        RECT 453.150 404.400 454.050 405.300 ;
        RECT 450.450 404.100 452.250 404.400 ;
        RECT 437.550 402.600 438.750 403.500 ;
        RECT 445.950 403.200 452.250 404.100 ;
        RECT 450.450 402.600 452.250 403.200 ;
        RECT 453.150 402.600 455.850 404.400 ;
        RECT 433.950 400.500 438.750 402.600 ;
        RECT 441.450 401.550 443.250 402.300 ;
        RECT 446.250 401.550 448.050 402.300 ;
        RECT 441.450 400.500 448.050 401.550 ;
        RECT 437.550 399.600 438.750 400.500 ;
        RECT 437.550 393.600 439.350 399.600 ;
        RECT 445.350 393.600 447.150 400.500 ;
        RECT 453.150 399.600 457.050 401.700 ;
        RECT 453.150 393.600 454.950 399.600 ;
        RECT 460.650 393.600 462.450 405.600 ;
        RECT 475.800 422.400 477.600 428.400 ;
        RECT 481.800 425.400 483.600 428.400 ;
        RECT 475.800 415.050 477.000 422.400 ;
        RECT 482.400 421.500 483.600 425.400 ;
        RECT 477.900 420.600 483.600 421.500 ;
        RECT 499.800 421.200 501.600 428.400 ;
        RECT 517.800 422.400 519.600 428.400 ;
        RECT 477.900 419.700 479.850 420.600 ;
        RECT 475.800 412.950 478.050 415.050 ;
        RECT 475.800 405.600 477.000 412.950 ;
        RECT 478.950 408.300 479.850 419.700 ;
        RECT 497.400 420.300 501.600 421.200 ;
        RECT 494.100 415.050 495.900 416.850 ;
        RECT 497.400 415.050 498.600 420.300 ;
        RECT 502.950 417.450 505.050 420.900 ;
        RECT 518.400 420.300 519.600 422.400 ;
        RECT 520.800 423.300 522.600 428.400 ;
        RECT 526.800 423.300 528.600 428.400 ;
        RECT 520.800 421.950 528.600 423.300 ;
        RECT 539.400 423.300 541.200 428.400 ;
        RECT 545.400 423.300 547.200 428.400 ;
        RECT 539.400 421.950 547.200 423.300 ;
        RECT 548.400 422.400 550.200 428.400 ;
        RECT 566.400 425.400 568.200 428.400 ;
        RECT 548.400 420.300 549.600 422.400 ;
        RECT 518.400 419.250 522.150 420.300 ;
        RECT 502.950 417.000 513.450 417.450 ;
        RECT 500.100 415.050 501.900 416.850 ;
        RECT 503.550 416.550 513.450 417.000 ;
        RECT 481.950 412.950 484.050 415.050 ;
        RECT 493.950 412.950 496.050 415.050 ;
        RECT 496.950 412.950 499.050 415.050 ;
        RECT 499.950 412.950 502.050 415.050 ;
        RECT 482.100 411.150 483.900 412.950 ;
        RECT 477.900 407.400 479.850 408.300 ;
        RECT 477.900 406.500 483.600 407.400 ;
        RECT 475.800 393.600 477.600 405.600 ;
        RECT 482.400 399.600 483.600 406.500 ;
        RECT 481.800 393.600 483.600 399.600 ;
        RECT 497.400 399.600 498.600 412.950 ;
        RECT 512.550 412.050 513.450 416.550 ;
        RECT 518.100 415.050 519.900 416.850 ;
        RECT 520.950 415.050 522.150 419.250 ;
        RECT 545.850 419.250 549.600 420.300 ;
        RECT 550.950 420.450 553.050 421.050 ;
        RECT 556.950 420.450 559.050 421.050 ;
        RECT 550.950 419.550 559.050 420.450 ;
        RECT 534.000 417.450 538.050 418.050 ;
        RECT 524.100 415.050 525.900 416.850 ;
        RECT 533.550 415.950 538.050 417.450 ;
        RECT 517.950 412.950 520.050 415.050 ;
        RECT 520.950 412.950 523.050 415.050 ;
        RECT 523.950 412.950 526.050 415.050 ;
        RECT 526.950 412.950 529.050 415.050 ;
        RECT 512.550 410.550 517.050 412.050 ;
        RECT 513.000 409.950 517.050 410.550 ;
        RECT 521.850 399.600 523.050 412.950 ;
        RECT 527.100 411.150 528.900 412.950 ;
        RECT 533.550 412.050 534.450 415.950 ;
        RECT 542.100 415.050 543.900 416.850 ;
        RECT 545.850 415.050 547.050 419.250 ;
        RECT 550.950 418.950 553.050 419.550 ;
        RECT 556.950 418.950 559.050 419.550 ;
        RECT 548.100 415.050 549.900 416.850 ;
        RECT 566.700 415.050 567.600 425.400 ;
        RECT 586.800 422.400 588.600 428.400 ;
        RECT 587.400 420.300 588.600 422.400 ;
        RECT 589.800 423.300 591.600 428.400 ;
        RECT 595.800 423.300 597.600 428.400 ;
        RECT 589.800 421.950 597.600 423.300 ;
        RECT 613.800 421.200 615.600 428.400 ;
        RECT 632.400 425.400 634.200 428.400 ;
        RECT 611.400 420.300 615.600 421.200 ;
        RECT 587.400 419.250 591.150 420.300 ;
        RECT 571.950 417.450 574.050 418.050 ;
        RECT 577.950 417.450 580.050 418.050 ;
        RECT 571.950 416.550 580.050 417.450 ;
        RECT 571.950 415.950 574.050 416.550 ;
        RECT 577.950 415.950 580.050 416.550 ;
        RECT 587.100 415.050 588.900 416.850 ;
        RECT 589.950 415.050 591.150 419.250 ;
        RECT 593.100 415.050 594.900 416.850 ;
        RECT 608.100 415.050 609.900 416.850 ;
        RECT 611.400 415.050 612.600 420.300 ;
        RECT 616.950 417.450 621.000 418.050 ;
        RECT 624.000 417.450 628.050 418.050 ;
        RECT 616.950 417.000 621.450 417.450 ;
        RECT 614.100 415.050 615.900 416.850 ;
        RECT 616.950 415.950 622.050 417.000 ;
        RECT 538.950 412.950 541.050 415.050 ;
        RECT 541.950 412.950 544.050 415.050 ;
        RECT 544.950 412.950 547.050 415.050 ;
        RECT 547.950 412.950 550.050 415.050 ;
        RECT 562.950 412.950 565.050 415.050 ;
        RECT 565.950 412.950 568.050 415.050 ;
        RECT 568.950 412.950 571.050 415.050 ;
        RECT 586.950 412.950 589.050 415.050 ;
        RECT 589.950 412.950 592.050 415.050 ;
        RECT 592.950 412.950 595.050 415.050 ;
        RECT 595.950 412.950 598.050 415.050 ;
        RECT 607.950 412.950 610.050 415.050 ;
        RECT 610.950 412.950 613.050 415.050 ;
        RECT 613.950 412.950 616.050 415.050 ;
        RECT 533.550 410.550 538.050 412.050 ;
        RECT 539.100 411.150 540.900 412.950 ;
        RECT 534.000 409.950 538.050 410.550 ;
        RECT 544.950 399.600 546.150 412.950 ;
        RECT 563.100 411.150 564.900 412.950 ;
        RECT 566.700 405.600 567.600 412.950 ;
        RECT 569.100 411.150 570.900 412.950 ;
        RECT 566.700 404.400 570.300 405.600 ;
        RECT 497.400 393.600 499.200 399.600 ;
        RECT 521.400 393.600 523.200 399.600 ;
        RECT 544.800 393.600 546.600 399.600 ;
        RECT 568.500 393.600 570.300 404.400 ;
        RECT 590.850 399.600 592.050 412.950 ;
        RECT 596.100 411.150 597.900 412.950 ;
        RECT 611.400 399.600 612.600 412.950 ;
        RECT 619.950 412.800 622.050 415.950 ;
        RECT 623.550 415.950 628.050 417.450 ;
        RECT 623.550 412.050 624.450 415.950 ;
        RECT 632.700 415.050 633.600 425.400 ;
        RECT 634.950 420.450 637.050 424.050 ;
        RECT 655.800 421.200 657.600 428.400 ;
        RECT 676.500 423.600 678.300 428.400 ;
        RECT 676.500 422.400 681.600 423.600 ;
        RECT 700.200 422.400 702.000 428.400 ;
        RECT 726.300 424.200 728.100 428.400 ;
        RECT 640.950 420.450 643.050 421.050 ;
        RECT 649.950 420.450 652.050 421.050 ;
        RECT 634.950 420.000 639.450 420.450 ;
        RECT 635.550 419.550 639.450 420.000 ;
        RECT 638.550 417.450 639.450 419.550 ;
        RECT 640.950 419.550 652.050 420.450 ;
        RECT 640.950 418.950 643.050 419.550 ;
        RECT 649.950 418.950 652.050 419.550 ;
        RECT 653.400 420.300 657.600 421.200 ;
        RECT 676.950 420.450 679.050 421.050 ;
        RECT 638.550 416.550 642.450 417.450 ;
        RECT 628.950 412.950 631.050 415.050 ;
        RECT 631.950 412.950 634.050 415.050 ;
        RECT 634.950 412.950 637.050 415.050 ;
        RECT 623.550 410.550 628.050 412.050 ;
        RECT 629.100 411.150 630.900 412.950 ;
        RECT 624.000 409.950 628.050 410.550 ;
        RECT 632.700 405.600 633.600 412.950 ;
        RECT 635.100 411.150 636.900 412.950 ;
        RECT 641.550 411.450 642.450 416.550 ;
        RECT 650.100 415.050 651.900 416.850 ;
        RECT 653.400 415.050 654.600 420.300 ;
        RECT 665.550 419.550 679.050 420.450 ;
        RECT 656.100 415.050 657.900 416.850 ;
        RECT 649.950 412.950 652.050 415.050 ;
        RECT 652.950 412.950 655.050 415.050 ;
        RECT 655.950 412.950 658.050 415.050 ;
        RECT 638.550 410.550 642.450 411.450 ;
        RECT 638.550 406.050 639.450 410.550 ;
        RECT 640.950 408.450 643.050 409.050 ;
        RECT 649.950 408.450 652.050 409.050 ;
        RECT 640.950 407.550 652.050 408.450 ;
        RECT 640.950 406.950 643.050 407.550 ;
        RECT 649.950 406.950 652.050 407.550 ;
        RECT 632.700 404.400 636.300 405.600 ;
        RECT 590.400 393.600 592.200 399.600 ;
        RECT 611.400 393.600 613.200 399.600 ;
        RECT 634.500 393.600 636.300 404.400 ;
        RECT 637.950 403.950 640.050 406.050 ;
        RECT 653.400 399.600 654.600 412.950 ;
        RECT 665.550 412.050 666.450 419.550 ;
        RECT 676.950 418.950 679.050 419.550 ;
        RECT 671.100 415.050 672.900 416.850 ;
        RECT 677.100 415.050 678.900 416.850 ;
        RECT 680.700 415.050 681.600 422.400 ;
        RECT 695.100 415.050 696.900 416.850 ;
        RECT 700.950 415.050 702.000 422.400 ;
        RECT 725.400 422.400 728.100 424.200 ;
        RECT 707.100 415.050 708.900 416.850 ;
        RECT 725.400 415.050 726.300 422.400 ;
        RECT 728.100 420.600 729.900 421.500 ;
        RECT 733.800 420.600 735.600 428.400 ;
        RECT 748.800 422.400 750.600 428.400 ;
        RECT 728.100 419.700 735.600 420.600 ;
        RECT 749.400 420.300 750.600 422.400 ;
        RECT 751.800 423.300 753.600 428.400 ;
        RECT 757.800 423.300 759.600 428.400 ;
        RECT 751.800 421.950 759.600 423.300 ;
        RECT 775.800 421.200 777.600 428.400 ;
        RECT 794.400 425.400 796.200 428.400 ;
        RECT 769.950 420.450 772.050 421.050 ;
        RECT 670.950 412.950 673.050 415.050 ;
        RECT 673.950 412.950 676.050 415.050 ;
        RECT 676.950 412.950 679.050 415.050 ;
        RECT 679.950 412.950 682.050 415.050 ;
        RECT 694.950 412.950 697.050 415.050 ;
        RECT 697.950 412.950 700.050 415.050 ;
        RECT 700.950 412.950 703.050 415.050 ;
        RECT 703.950 412.950 706.050 415.050 ;
        RECT 706.950 412.950 709.050 415.050 ;
        RECT 724.950 412.950 727.050 415.050 ;
        RECT 727.950 412.950 730.050 415.050 ;
        RECT 665.550 410.550 670.050 412.050 ;
        RECT 674.100 411.150 675.900 412.950 ;
        RECT 666.000 409.950 670.050 410.550 ;
        RECT 661.950 408.450 664.050 409.050 ;
        RECT 670.950 408.450 673.050 409.050 ;
        RECT 661.950 407.550 673.050 408.450 ;
        RECT 661.950 406.950 664.050 407.550 ;
        RECT 670.950 406.950 673.050 407.550 ;
        RECT 680.700 405.600 681.600 412.950 ;
        RECT 698.100 411.150 699.900 412.950 ;
        RECT 701.100 407.400 702.000 412.950 ;
        RECT 704.100 411.150 705.900 412.950 ;
        RECT 701.100 406.500 706.200 407.400 ;
        RECT 671.400 404.700 679.200 405.600 ;
        RECT 653.400 393.600 655.200 399.600 ;
        RECT 671.400 393.600 673.200 404.700 ;
        RECT 677.400 393.600 679.200 404.700 ;
        RECT 680.400 393.600 682.200 405.600 ;
        RECT 695.400 404.400 703.200 405.300 ;
        RECT 695.400 393.600 697.200 404.400 ;
        RECT 701.400 394.500 703.200 404.400 ;
        RECT 704.400 395.400 706.200 406.500 ;
        RECT 725.400 405.600 726.300 412.950 ;
        RECT 728.100 411.150 729.900 412.950 ;
        RECT 707.400 394.500 709.200 405.600 ;
        RECT 701.400 393.600 709.200 394.500 ;
        RECT 724.800 393.600 726.600 405.600 ;
        RECT 731.700 399.600 732.600 419.700 ;
        RECT 749.400 419.250 753.150 420.300 ;
        RECT 736.950 417.450 739.050 418.050 ;
        RECT 734.100 415.050 735.900 416.850 ;
        RECT 736.950 416.550 744.450 417.450 ;
        RECT 736.950 415.950 739.050 416.550 ;
        RECT 733.950 412.950 736.050 415.050 ;
        RECT 743.550 412.050 744.450 416.550 ;
        RECT 749.100 415.050 750.900 416.850 ;
        RECT 751.950 415.050 753.150 419.250 ;
        RECT 764.550 419.550 772.050 420.450 ;
        RECT 755.100 415.050 756.900 416.850 ;
        RECT 748.950 412.950 751.050 415.050 ;
        RECT 751.950 412.950 754.050 415.050 ;
        RECT 754.950 412.950 757.050 415.050 ;
        RECT 757.950 412.950 760.050 415.050 ;
        RECT 743.550 410.550 748.050 412.050 ;
        RECT 744.000 409.950 748.050 410.550 ;
        RECT 752.850 399.600 754.050 412.950 ;
        RECT 758.100 411.150 759.900 412.950 ;
        RECT 764.550 412.050 765.450 419.550 ;
        RECT 769.950 418.950 772.050 419.550 ;
        RECT 773.400 420.300 777.600 421.200 ;
        RECT 795.300 421.200 796.200 425.400 ;
        RECT 800.400 422.400 802.200 428.400 ;
        RECT 817.800 422.400 819.600 428.400 ;
        RECT 795.300 420.300 798.600 421.200 ;
        RECT 770.100 415.050 771.900 416.850 ;
        RECT 773.400 415.050 774.600 420.300 ;
        RECT 796.800 419.400 798.600 420.300 ;
        RECT 776.100 415.050 777.900 416.850 ;
        RECT 791.100 415.050 792.900 416.850 ;
        RECT 769.950 412.950 772.050 415.050 ;
        RECT 772.950 412.950 775.050 415.050 ;
        RECT 775.950 412.950 778.050 415.050 ;
        RECT 790.950 412.950 793.050 415.050 ;
        RECT 793.950 412.950 796.050 415.050 ;
        RECT 764.550 410.550 769.050 412.050 ;
        RECT 765.000 409.950 769.050 410.550 ;
        RECT 773.400 399.600 774.600 412.950 ;
        RECT 794.100 411.150 795.900 412.950 ;
        RECT 797.700 408.900 798.600 419.400 ;
        RECT 801.000 415.050 802.050 422.400 ;
        RECT 818.400 420.300 819.600 422.400 ;
        RECT 820.800 423.300 822.600 428.400 ;
        RECT 826.800 423.300 828.600 428.400 ;
        RECT 842.400 425.400 844.200 428.400 ;
        RECT 820.800 421.950 828.600 423.300 ;
        RECT 818.400 419.250 822.150 420.300 ;
        RECT 813.000 417.450 817.050 418.050 ;
        RECT 796.800 408.300 798.600 408.900 ;
        RECT 791.400 407.100 798.600 408.300 ;
        RECT 799.950 412.950 802.050 415.050 ;
        RECT 812.550 415.950 817.050 417.450 ;
        RECT 791.400 405.600 792.600 407.100 ;
        RECT 799.950 405.600 801.300 412.950 ;
        RECT 812.550 412.050 813.450 415.950 ;
        RECT 818.100 415.050 819.900 416.850 ;
        RECT 820.950 415.050 822.150 419.250 ;
        RECT 824.100 415.050 825.900 416.850 ;
        RECT 842.700 415.050 843.600 425.400 ;
        RECT 860.400 423.300 862.200 428.400 ;
        RECT 866.400 423.300 868.200 428.400 ;
        RECT 860.400 421.950 868.200 423.300 ;
        RECT 869.400 422.400 871.200 428.400 ;
        RECT 869.400 420.300 870.600 422.400 ;
        RECT 889.800 421.200 891.600 428.400 ;
        RECT 866.850 419.250 870.600 420.300 ;
        RECT 887.400 420.300 891.600 421.200 ;
        RECT 863.100 415.050 864.900 416.850 ;
        RECT 866.850 415.050 868.050 419.250 ;
        RECT 871.950 417.450 876.000 418.050 ;
        RECT 869.100 415.050 870.900 416.850 ;
        RECT 871.950 415.950 876.450 417.450 ;
        RECT 817.950 412.950 820.050 415.050 ;
        RECT 820.950 412.950 823.050 415.050 ;
        RECT 823.950 412.950 826.050 415.050 ;
        RECT 826.950 412.950 829.050 415.050 ;
        RECT 838.950 412.950 841.050 415.050 ;
        RECT 841.950 412.950 844.050 415.050 ;
        RECT 844.950 412.950 847.050 415.050 ;
        RECT 859.950 412.950 862.050 415.050 ;
        RECT 862.950 412.950 865.050 415.050 ;
        RECT 865.950 412.950 868.050 415.050 ;
        RECT 868.950 412.950 871.050 415.050 ;
        RECT 812.550 410.550 817.050 412.050 ;
        RECT 813.000 409.950 817.050 410.550 ;
        RECT 805.950 408.450 808.050 409.050 ;
        RECT 817.950 408.450 820.050 409.050 ;
        RECT 805.950 407.550 820.050 408.450 ;
        RECT 805.950 406.950 808.050 407.550 ;
        RECT 817.950 406.950 820.050 407.550 ;
        RECT 730.800 393.600 732.600 399.600 ;
        RECT 752.400 393.600 754.200 399.600 ;
        RECT 773.400 393.600 775.200 399.600 ;
        RECT 791.400 393.600 793.200 405.600 ;
        RECT 798.900 404.100 801.300 405.600 ;
        RECT 798.900 393.600 800.700 404.100 ;
        RECT 821.850 399.600 823.050 412.950 ;
        RECT 827.100 411.150 828.900 412.950 ;
        RECT 839.100 411.150 840.900 412.950 ;
        RECT 842.700 405.600 843.600 412.950 ;
        RECT 845.100 411.150 846.900 412.950 ;
        RECT 860.100 411.150 861.900 412.950 ;
        RECT 842.700 404.400 846.300 405.600 ;
        RECT 821.400 393.600 823.200 399.600 ;
        RECT 844.500 393.600 846.300 404.400 ;
        RECT 865.950 399.600 867.150 412.950 ;
        RECT 875.550 408.450 876.450 415.950 ;
        RECT 884.100 415.050 885.900 416.850 ;
        RECT 887.400 415.050 888.600 420.300 ;
        RECT 890.100 415.050 891.900 416.850 ;
        RECT 883.950 412.950 886.050 415.050 ;
        RECT 886.950 412.950 889.050 415.050 ;
        RECT 889.950 412.950 892.050 415.050 ;
        RECT 883.950 408.450 886.050 408.750 ;
        RECT 875.550 407.550 886.050 408.450 ;
        RECT 883.950 406.650 886.050 407.550 ;
        RECT 887.400 399.600 888.600 412.950 ;
        RECT 865.800 393.600 867.600 399.600 ;
        RECT 887.400 393.600 889.200 399.600 ;
        RECT 3.150 377.400 4.950 389.400 ;
        RECT 11.550 383.400 13.350 389.400 ;
        RECT 11.550 382.500 12.750 383.400 ;
        RECT 19.350 382.500 21.150 389.400 ;
        RECT 27.150 383.400 28.950 389.400 ;
        RECT 7.950 380.400 12.750 382.500 ;
        RECT 15.450 381.450 22.050 382.500 ;
        RECT 15.450 380.700 17.250 381.450 ;
        RECT 20.250 380.700 22.050 381.450 ;
        RECT 27.150 381.300 31.050 383.400 ;
        RECT 11.550 379.500 12.750 380.400 ;
        RECT 24.450 379.800 26.250 380.400 ;
        RECT 11.550 378.300 19.050 379.500 ;
        RECT 17.250 377.700 19.050 378.300 ;
        RECT 19.950 378.900 26.250 379.800 ;
        RECT 3.150 376.500 4.050 377.400 ;
        RECT 19.950 376.800 20.850 378.900 ;
        RECT 24.450 378.600 26.250 378.900 ;
        RECT 27.150 378.600 29.850 380.400 ;
        RECT 27.150 377.700 28.050 378.600 ;
        RECT 12.450 376.500 20.850 376.800 ;
        RECT 3.150 375.900 20.850 376.500 ;
        RECT 22.950 376.800 28.050 377.700 ;
        RECT 28.950 376.800 31.050 377.700 ;
        RECT 34.650 377.400 36.450 389.400 ;
        RECT 53.400 383.400 55.200 389.400 ;
        RECT 76.800 383.400 78.600 389.400 ;
        RECT 3.150 375.300 14.250 375.900 ;
        RECT 3.150 360.600 4.050 375.300 ;
        RECT 12.450 375.000 14.250 375.300 ;
        RECT 4.950 367.950 7.050 370.050 ;
        RECT 13.950 368.400 16.050 370.050 ;
        RECT 5.100 366.150 6.900 367.950 ;
        RECT 8.100 367.200 16.050 368.400 ;
        RECT 8.100 366.600 9.900 367.200 ;
        RECT 6.000 365.400 6.900 366.150 ;
        RECT 11.100 365.400 12.900 366.000 ;
        RECT 6.000 364.200 12.900 365.400 ;
        RECT 22.950 364.200 23.850 376.800 ;
        RECT 28.950 375.600 33.150 376.800 ;
        RECT 32.250 373.800 34.050 375.600 ;
        RECT 35.250 370.050 36.450 377.400 ;
        RECT 53.850 370.050 55.050 383.400 ;
        RECT 69.000 372.450 73.050 373.050 ;
        RECT 59.100 370.050 60.900 371.850 ;
        RECT 68.550 370.950 73.050 372.450 ;
        RECT 31.950 369.750 36.450 370.050 ;
        RECT 30.150 367.950 36.450 369.750 ;
        RECT 49.950 367.950 52.050 370.050 ;
        RECT 52.950 367.950 55.050 370.050 ;
        RECT 55.950 367.950 58.050 370.050 ;
        RECT 58.950 367.950 61.050 370.050 ;
        RECT 11.850 363.000 23.850 364.200 ;
        RECT 11.850 361.200 12.900 363.000 ;
        RECT 22.050 362.400 23.850 363.000 ;
        RECT 3.150 354.600 4.950 360.600 ;
        RECT 7.950 358.500 10.050 360.600 ;
        RECT 11.550 359.400 13.350 361.200 ;
        RECT 35.250 360.600 36.450 367.950 ;
        RECT 50.100 366.150 51.900 367.950 ;
        RECT 52.950 363.750 54.150 367.950 ;
        RECT 56.100 366.150 57.900 367.950 ;
        RECT 68.550 363.900 69.450 370.950 ;
        RECT 77.400 370.050 78.600 383.400 ;
        RECT 83.550 377.400 85.350 389.400 ;
        RECT 91.050 383.400 92.850 389.400 ;
        RECT 88.950 381.300 92.850 383.400 ;
        RECT 98.850 382.500 100.650 389.400 ;
        RECT 106.650 383.400 108.450 389.400 ;
        RECT 107.250 382.500 108.450 383.400 ;
        RECT 97.950 381.450 104.550 382.500 ;
        RECT 97.950 380.700 99.750 381.450 ;
        RECT 102.750 380.700 104.550 381.450 ;
        RECT 107.250 380.400 112.050 382.500 ;
        RECT 90.150 378.600 92.850 380.400 ;
        RECT 93.750 379.800 95.550 380.400 ;
        RECT 93.750 378.900 100.050 379.800 ;
        RECT 107.250 379.500 108.450 380.400 ;
        RECT 93.750 378.600 95.550 378.900 ;
        RECT 91.950 377.700 92.850 378.600 ;
        RECT 83.550 370.050 84.750 377.400 ;
        RECT 88.950 376.800 91.050 377.700 ;
        RECT 91.950 376.800 97.050 377.700 ;
        RECT 86.850 375.600 91.050 376.800 ;
        RECT 85.950 373.800 87.750 375.600 ;
        RECT 73.950 367.950 76.050 370.050 ;
        RECT 76.950 367.950 79.050 370.050 ;
        RECT 79.950 367.950 82.050 370.050 ;
        RECT 83.550 369.750 88.050 370.050 ;
        RECT 83.550 367.950 89.850 369.750 ;
        RECT 74.100 366.150 75.900 367.950 ;
        RECT 50.400 362.700 54.150 363.750 ;
        RECT 50.400 360.600 51.600 362.700 ;
        RECT 67.950 361.800 70.050 363.900 ;
        RECT 77.400 362.700 78.600 367.950 ;
        RECT 80.100 366.150 81.900 367.950 ;
        RECT 74.400 361.800 78.600 362.700 ;
        RECT 14.850 359.550 16.650 360.300 ;
        RECT 28.950 359.700 31.050 360.600 ;
        RECT 14.850 358.500 19.800 359.550 ;
        RECT 9.000 357.600 10.050 358.500 ;
        RECT 18.750 357.600 19.800 358.500 ;
        RECT 27.300 358.500 31.050 359.700 ;
        RECT 27.300 357.600 28.350 358.500 ;
        RECT 9.000 356.700 12.750 357.600 ;
        RECT 10.950 354.600 12.750 356.700 ;
        RECT 18.750 354.600 20.550 357.600 ;
        RECT 26.550 354.600 28.350 357.600 ;
        RECT 34.650 354.600 36.450 360.600 ;
        RECT 49.800 354.600 51.600 360.600 ;
        RECT 52.800 359.700 60.600 361.050 ;
        RECT 52.800 354.600 54.600 359.700 ;
        RECT 58.800 354.600 60.600 359.700 ;
        RECT 74.400 354.600 76.200 361.800 ;
        RECT 83.550 360.600 84.750 367.950 ;
        RECT 96.150 364.200 97.050 376.800 ;
        RECT 99.150 376.800 100.050 378.900 ;
        RECT 100.950 378.300 108.450 379.500 ;
        RECT 100.950 377.700 102.750 378.300 ;
        RECT 115.050 377.400 116.850 389.400 ;
        RECT 99.150 376.500 107.550 376.800 ;
        RECT 115.950 376.500 116.850 377.400 ;
        RECT 99.150 375.900 116.850 376.500 ;
        RECT 105.750 375.300 116.850 375.900 ;
        RECT 105.750 375.000 107.550 375.300 ;
        RECT 103.950 368.400 106.050 370.050 ;
        RECT 103.950 367.200 111.900 368.400 ;
        RECT 112.950 367.950 115.050 370.050 ;
        RECT 110.100 366.600 111.900 367.200 ;
        RECT 113.100 366.150 114.900 367.950 ;
        RECT 107.100 365.400 108.900 366.000 ;
        RECT 113.100 365.400 114.000 366.150 ;
        RECT 107.100 364.200 114.000 365.400 ;
        RECT 96.150 363.000 108.150 364.200 ;
        RECT 96.150 362.400 97.950 363.000 ;
        RECT 107.100 361.200 108.150 363.000 ;
        RECT 83.550 354.600 85.350 360.600 ;
        RECT 88.950 359.700 91.050 360.600 ;
        RECT 88.950 358.500 92.700 359.700 ;
        RECT 103.350 359.550 105.150 360.300 ;
        RECT 91.650 357.600 92.700 358.500 ;
        RECT 100.200 358.500 105.150 359.550 ;
        RECT 106.650 359.400 108.450 361.200 ;
        RECT 115.950 360.600 116.850 375.300 ;
        RECT 109.950 358.500 112.050 360.600 ;
        RECT 100.200 357.600 101.250 358.500 ;
        RECT 109.950 357.600 111.000 358.500 ;
        RECT 91.650 354.600 93.450 357.600 ;
        RECT 99.450 354.600 101.250 357.600 ;
        RECT 107.250 356.700 111.000 357.600 ;
        RECT 107.250 354.600 109.050 356.700 ;
        RECT 115.050 354.600 116.850 360.600 ;
        RECT 130.800 377.400 132.600 389.400 ;
        RECT 136.800 383.400 138.600 389.400 ;
        RECT 130.800 370.050 132.000 377.400 ;
        RECT 137.400 376.500 138.600 383.400 ;
        RECT 152.700 378.600 154.500 389.400 ;
        RECT 175.800 383.400 177.600 389.400 ;
        RECT 152.700 377.400 156.300 378.600 ;
        RECT 132.900 375.600 138.600 376.500 ;
        RECT 132.900 374.700 134.850 375.600 ;
        RECT 130.800 367.950 133.050 370.050 ;
        RECT 130.800 360.600 132.000 367.950 ;
        RECT 133.950 363.300 134.850 374.700 ;
        RECT 137.100 370.050 138.900 371.850 ;
        RECT 152.100 370.050 153.900 371.850 ;
        RECT 155.400 370.050 156.300 377.400 ;
        RECT 158.100 370.050 159.900 371.850 ;
        RECT 170.100 370.050 171.900 371.850 ;
        RECT 175.950 370.050 177.150 383.400 ;
        RECT 197.700 378.600 199.500 389.400 ;
        RECT 197.700 377.400 201.300 378.600 ;
        RECT 197.100 370.050 198.900 371.850 ;
        RECT 200.400 370.050 201.300 377.400 ;
        RECT 206.550 377.400 208.350 389.400 ;
        RECT 214.050 383.400 215.850 389.400 ;
        RECT 211.950 381.300 215.850 383.400 ;
        RECT 221.850 382.500 223.650 389.400 ;
        RECT 229.650 383.400 231.450 389.400 ;
        RECT 230.250 382.500 231.450 383.400 ;
        RECT 220.950 381.450 227.550 382.500 ;
        RECT 220.950 380.700 222.750 381.450 ;
        RECT 225.750 380.700 227.550 381.450 ;
        RECT 230.250 380.400 235.050 382.500 ;
        RECT 213.150 378.600 215.850 380.400 ;
        RECT 216.750 379.800 218.550 380.400 ;
        RECT 216.750 378.900 223.050 379.800 ;
        RECT 230.250 379.500 231.450 380.400 ;
        RECT 216.750 378.600 218.550 378.900 ;
        RECT 214.950 377.700 215.850 378.600 ;
        RECT 203.100 370.050 204.900 371.850 ;
        RECT 206.550 370.050 207.750 377.400 ;
        RECT 211.950 376.800 214.050 377.700 ;
        RECT 214.950 376.800 220.050 377.700 ;
        RECT 209.850 375.600 214.050 376.800 ;
        RECT 208.950 373.800 210.750 375.600 ;
        RECT 136.950 367.950 139.050 370.050 ;
        RECT 151.950 367.950 154.050 370.050 ;
        RECT 154.950 367.950 157.050 370.050 ;
        RECT 157.950 367.950 160.050 370.050 ;
        RECT 169.950 367.950 172.050 370.050 ;
        RECT 172.950 367.950 175.050 370.050 ;
        RECT 175.950 367.950 178.050 370.050 ;
        RECT 178.950 367.950 181.050 370.050 ;
        RECT 196.950 367.950 199.050 370.050 ;
        RECT 199.950 367.950 202.050 370.050 ;
        RECT 202.950 367.950 205.050 370.050 ;
        RECT 206.550 369.750 211.050 370.050 ;
        RECT 206.550 367.950 212.850 369.750 ;
        RECT 132.900 362.400 134.850 363.300 ;
        RECT 132.900 361.500 138.600 362.400 ;
        RECT 130.800 354.600 132.600 360.600 ;
        RECT 137.400 357.600 138.600 361.500 ;
        RECT 155.400 357.600 156.300 367.950 ;
        RECT 173.100 366.150 174.900 367.950 ;
        RECT 176.850 363.750 178.050 367.950 ;
        RECT 179.100 366.150 180.900 367.950 ;
        RECT 176.850 362.700 180.600 363.750 ;
        RECT 170.400 359.700 178.200 361.050 ;
        RECT 136.800 354.600 138.600 357.600 ;
        RECT 154.800 354.600 156.600 357.600 ;
        RECT 170.400 354.600 172.200 359.700 ;
        RECT 176.400 354.600 178.200 359.700 ;
        RECT 179.400 360.600 180.600 362.700 ;
        RECT 179.400 354.600 181.200 360.600 ;
        RECT 200.400 357.600 201.300 367.950 ;
        RECT 206.550 360.600 207.750 367.950 ;
        RECT 219.150 364.200 220.050 376.800 ;
        RECT 222.150 376.800 223.050 378.900 ;
        RECT 223.950 378.300 231.450 379.500 ;
        RECT 223.950 377.700 225.750 378.300 ;
        RECT 238.050 377.400 239.850 389.400 ;
        RECT 256.800 383.400 258.600 389.400 ;
        RECT 281.400 383.400 283.200 389.400 ;
        RECT 222.150 376.500 230.550 376.800 ;
        RECT 238.950 376.500 239.850 377.400 ;
        RECT 222.150 375.900 239.850 376.500 ;
        RECT 228.750 375.300 239.850 375.900 ;
        RECT 228.750 375.000 230.550 375.300 ;
        RECT 226.950 368.400 229.050 370.050 ;
        RECT 226.950 367.200 234.900 368.400 ;
        RECT 235.950 367.950 238.050 370.050 ;
        RECT 233.100 366.600 234.900 367.200 ;
        RECT 236.100 366.150 237.900 367.950 ;
        RECT 230.100 365.400 231.900 366.000 ;
        RECT 236.100 365.400 237.000 366.150 ;
        RECT 230.100 364.200 237.000 365.400 ;
        RECT 219.150 363.000 231.150 364.200 ;
        RECT 219.150 362.400 220.950 363.000 ;
        RECT 230.100 361.200 231.150 363.000 ;
        RECT 199.800 354.600 201.600 357.600 ;
        RECT 206.550 354.600 208.350 360.600 ;
        RECT 211.950 359.700 214.050 360.600 ;
        RECT 211.950 358.500 215.700 359.700 ;
        RECT 226.350 359.550 228.150 360.300 ;
        RECT 214.650 357.600 215.700 358.500 ;
        RECT 223.200 358.500 228.150 359.550 ;
        RECT 229.650 359.400 231.450 361.200 ;
        RECT 238.950 360.600 239.850 375.300 ;
        RECT 251.100 370.050 252.900 371.850 ;
        RECT 256.950 370.050 258.150 383.400 ;
        RECT 259.950 378.450 262.050 379.050 ;
        RECT 277.950 378.450 280.050 379.050 ;
        RECT 259.950 377.550 280.050 378.450 ;
        RECT 259.950 376.950 262.050 377.550 ;
        RECT 277.950 376.950 280.050 377.550 ;
        RECT 281.400 370.050 282.600 383.400 ;
        RECT 302.400 377.400 304.200 389.400 ;
        RECT 322.800 383.400 324.600 389.400 ;
        RECT 343.800 383.400 345.600 389.400 ;
        RECT 302.400 370.050 303.600 377.400 ;
        RECT 323.400 370.050 324.600 383.400 ;
        RECT 326.100 370.050 327.900 371.850 ;
        RECT 338.100 370.050 339.900 371.850 ;
        RECT 343.950 370.050 345.150 383.400 ;
        RECT 353.550 377.400 355.350 389.400 ;
        RECT 361.050 383.400 362.850 389.400 ;
        RECT 358.950 381.300 362.850 383.400 ;
        RECT 368.850 382.500 370.650 389.400 ;
        RECT 376.650 383.400 378.450 389.400 ;
        RECT 377.250 382.500 378.450 383.400 ;
        RECT 367.950 381.450 374.550 382.500 ;
        RECT 367.950 380.700 369.750 381.450 ;
        RECT 372.750 380.700 374.550 381.450 ;
        RECT 377.250 380.400 382.050 382.500 ;
        RECT 360.150 378.600 362.850 380.400 ;
        RECT 363.750 379.800 365.550 380.400 ;
        RECT 363.750 378.900 370.050 379.800 ;
        RECT 377.250 379.500 378.450 380.400 ;
        RECT 363.750 378.600 365.550 378.900 ;
        RECT 361.950 377.700 362.850 378.600 ;
        RECT 353.550 370.050 354.750 377.400 ;
        RECT 358.950 376.800 361.050 377.700 ;
        RECT 361.950 376.800 367.050 377.700 ;
        RECT 356.850 375.600 361.050 376.800 ;
        RECT 355.950 373.800 357.750 375.600 ;
        RECT 250.950 367.950 253.050 370.050 ;
        RECT 253.950 367.950 256.050 370.050 ;
        RECT 256.950 367.950 259.050 370.050 ;
        RECT 259.950 367.950 262.050 370.050 ;
        RECT 277.950 367.950 280.050 370.050 ;
        RECT 280.950 367.950 283.050 370.050 ;
        RECT 283.950 367.950 286.050 370.050 ;
        RECT 298.950 367.950 301.050 370.050 ;
        RECT 301.950 367.950 304.050 370.050 ;
        RECT 322.950 367.950 325.050 370.050 ;
        RECT 325.950 367.950 328.050 370.050 ;
        RECT 337.950 367.950 340.050 370.050 ;
        RECT 340.950 367.950 343.050 370.050 ;
        RECT 343.950 367.950 346.050 370.050 ;
        RECT 346.950 367.950 349.050 370.050 ;
        RECT 353.550 369.750 358.050 370.050 ;
        RECT 353.550 367.950 359.850 369.750 ;
        RECT 254.100 366.150 255.900 367.950 ;
        RECT 257.850 363.750 259.050 367.950 ;
        RECT 260.100 366.150 261.900 367.950 ;
        RECT 278.100 366.150 279.900 367.950 ;
        RECT 257.850 362.700 261.600 363.750 ;
        RECT 232.950 358.500 235.050 360.600 ;
        RECT 223.200 357.600 224.250 358.500 ;
        RECT 232.950 357.600 234.000 358.500 ;
        RECT 214.650 354.600 216.450 357.600 ;
        RECT 222.450 354.600 224.250 357.600 ;
        RECT 230.250 356.700 234.000 357.600 ;
        RECT 230.250 354.600 232.050 356.700 ;
        RECT 238.050 354.600 239.850 360.600 ;
        RECT 251.400 359.700 259.200 361.050 ;
        RECT 251.400 354.600 253.200 359.700 ;
        RECT 257.400 354.600 259.200 359.700 ;
        RECT 260.400 360.600 261.600 362.700 ;
        RECT 281.400 362.700 282.600 367.950 ;
        RECT 284.100 366.150 285.900 367.950 ;
        RECT 299.100 366.150 300.900 367.950 ;
        RECT 281.400 361.800 285.600 362.700 ;
        RECT 260.400 354.600 262.200 360.600 ;
        RECT 283.800 354.600 285.600 361.800 ;
        RECT 302.400 360.600 303.600 367.950 ;
        RECT 302.400 354.600 304.200 360.600 ;
        RECT 323.400 357.600 324.600 367.950 ;
        RECT 341.100 366.150 342.900 367.950 ;
        RECT 344.850 363.750 346.050 367.950 ;
        RECT 347.100 366.150 348.900 367.950 ;
        RECT 344.850 362.700 348.600 363.750 ;
        RECT 322.800 354.600 324.600 357.600 ;
        RECT 338.400 359.700 346.200 361.050 ;
        RECT 338.400 354.600 340.200 359.700 ;
        RECT 344.400 354.600 346.200 359.700 ;
        RECT 347.400 360.600 348.600 362.700 ;
        RECT 353.550 360.600 354.750 367.950 ;
        RECT 366.150 364.200 367.050 376.800 ;
        RECT 369.150 376.800 370.050 378.900 ;
        RECT 370.950 378.300 378.450 379.500 ;
        RECT 370.950 377.700 372.750 378.300 ;
        RECT 385.050 377.400 386.850 389.400 ;
        RECT 369.150 376.500 377.550 376.800 ;
        RECT 385.950 376.500 386.850 377.400 ;
        RECT 369.150 375.900 386.850 376.500 ;
        RECT 375.750 375.300 386.850 375.900 ;
        RECT 375.750 375.000 377.550 375.300 ;
        RECT 373.950 368.400 376.050 370.050 ;
        RECT 373.950 367.200 381.900 368.400 ;
        RECT 382.950 367.950 385.050 370.050 ;
        RECT 380.100 366.600 381.900 367.200 ;
        RECT 383.100 366.150 384.900 367.950 ;
        RECT 377.100 365.400 378.900 366.000 ;
        RECT 383.100 365.400 384.000 366.150 ;
        RECT 377.100 364.200 384.000 365.400 ;
        RECT 366.150 363.000 378.150 364.200 ;
        RECT 366.150 362.400 367.950 363.000 ;
        RECT 377.100 361.200 378.150 363.000 ;
        RECT 347.400 354.600 349.200 360.600 ;
        RECT 353.550 354.600 355.350 360.600 ;
        RECT 358.950 359.700 361.050 360.600 ;
        RECT 358.950 358.500 362.700 359.700 ;
        RECT 373.350 359.550 375.150 360.300 ;
        RECT 361.650 357.600 362.700 358.500 ;
        RECT 370.200 358.500 375.150 359.550 ;
        RECT 376.650 359.400 378.450 361.200 ;
        RECT 385.950 360.600 386.850 375.300 ;
        RECT 379.950 358.500 382.050 360.600 ;
        RECT 370.200 357.600 371.250 358.500 ;
        RECT 379.950 357.600 381.000 358.500 ;
        RECT 361.650 354.600 363.450 357.600 ;
        RECT 369.450 354.600 371.250 357.600 ;
        RECT 377.250 356.700 381.000 357.600 ;
        RECT 377.250 354.600 379.050 356.700 ;
        RECT 385.050 354.600 386.850 360.600 ;
        RECT 389.550 377.400 391.350 389.400 ;
        RECT 397.050 383.400 398.850 389.400 ;
        RECT 394.950 381.300 398.850 383.400 ;
        RECT 404.850 382.500 406.650 389.400 ;
        RECT 412.650 383.400 414.450 389.400 ;
        RECT 413.250 382.500 414.450 383.400 ;
        RECT 403.950 381.450 410.550 382.500 ;
        RECT 403.950 380.700 405.750 381.450 ;
        RECT 408.750 380.700 410.550 381.450 ;
        RECT 413.250 380.400 418.050 382.500 ;
        RECT 396.150 378.600 398.850 380.400 ;
        RECT 399.750 379.800 401.550 380.400 ;
        RECT 399.750 378.900 406.050 379.800 ;
        RECT 413.250 379.500 414.450 380.400 ;
        RECT 399.750 378.600 401.550 378.900 ;
        RECT 397.950 377.700 398.850 378.600 ;
        RECT 389.550 370.050 390.750 377.400 ;
        RECT 394.950 376.800 397.050 377.700 ;
        RECT 397.950 376.800 403.050 377.700 ;
        RECT 392.850 375.600 397.050 376.800 ;
        RECT 391.950 373.800 393.750 375.600 ;
        RECT 389.550 369.750 394.050 370.050 ;
        RECT 389.550 367.950 395.850 369.750 ;
        RECT 389.550 360.600 390.750 367.950 ;
        RECT 402.150 364.200 403.050 376.800 ;
        RECT 405.150 376.800 406.050 378.900 ;
        RECT 406.950 378.300 414.450 379.500 ;
        RECT 406.950 377.700 408.750 378.300 ;
        RECT 421.050 377.400 422.850 389.400 ;
        RECT 405.150 376.500 413.550 376.800 ;
        RECT 421.950 376.500 422.850 377.400 ;
        RECT 405.150 375.900 422.850 376.500 ;
        RECT 411.750 375.300 422.850 375.900 ;
        RECT 411.750 375.000 413.550 375.300 ;
        RECT 409.950 368.400 412.050 370.050 ;
        RECT 409.950 367.200 417.900 368.400 ;
        RECT 418.950 367.950 421.050 370.050 ;
        RECT 416.100 366.600 417.900 367.200 ;
        RECT 419.100 366.150 420.900 367.950 ;
        RECT 413.100 365.400 414.900 366.000 ;
        RECT 419.100 365.400 420.000 366.150 ;
        RECT 413.100 364.200 420.000 365.400 ;
        RECT 402.150 363.000 414.150 364.200 ;
        RECT 402.150 362.400 403.950 363.000 ;
        RECT 413.100 361.200 414.150 363.000 ;
        RECT 389.550 354.600 391.350 360.600 ;
        RECT 394.950 359.700 397.050 360.600 ;
        RECT 394.950 358.500 398.700 359.700 ;
        RECT 409.350 359.550 411.150 360.300 ;
        RECT 397.650 357.600 398.700 358.500 ;
        RECT 406.200 358.500 411.150 359.550 ;
        RECT 412.650 359.400 414.450 361.200 ;
        RECT 421.950 360.600 422.850 375.300 ;
        RECT 415.950 358.500 418.050 360.600 ;
        RECT 406.200 357.600 407.250 358.500 ;
        RECT 415.950 357.600 417.000 358.500 ;
        RECT 397.650 354.600 399.450 357.600 ;
        RECT 405.450 354.600 407.250 357.600 ;
        RECT 413.250 356.700 417.000 357.600 ;
        RECT 413.250 354.600 415.050 356.700 ;
        RECT 421.050 354.600 422.850 360.600 ;
        RECT 426.150 377.400 427.950 389.400 ;
        RECT 434.550 383.400 436.350 389.400 ;
        RECT 434.550 382.500 435.750 383.400 ;
        RECT 442.350 382.500 444.150 389.400 ;
        RECT 450.150 383.400 451.950 389.400 ;
        RECT 430.950 380.400 435.750 382.500 ;
        RECT 438.450 381.450 445.050 382.500 ;
        RECT 438.450 380.700 440.250 381.450 ;
        RECT 443.250 380.700 445.050 381.450 ;
        RECT 450.150 381.300 454.050 383.400 ;
        RECT 434.550 379.500 435.750 380.400 ;
        RECT 447.450 379.800 449.250 380.400 ;
        RECT 434.550 378.300 442.050 379.500 ;
        RECT 440.250 377.700 442.050 378.300 ;
        RECT 442.950 378.900 449.250 379.800 ;
        RECT 426.150 376.500 427.050 377.400 ;
        RECT 442.950 376.800 443.850 378.900 ;
        RECT 447.450 378.600 449.250 378.900 ;
        RECT 450.150 378.600 452.850 380.400 ;
        RECT 450.150 377.700 451.050 378.600 ;
        RECT 435.450 376.500 443.850 376.800 ;
        RECT 426.150 375.900 443.850 376.500 ;
        RECT 445.950 376.800 451.050 377.700 ;
        RECT 451.950 376.800 454.050 377.700 ;
        RECT 457.650 377.400 459.450 389.400 ;
        RECT 475.500 378.600 477.300 389.400 ;
        RECT 426.150 375.300 437.250 375.900 ;
        RECT 426.150 360.600 427.050 375.300 ;
        RECT 435.450 375.000 437.250 375.300 ;
        RECT 427.950 367.950 430.050 370.050 ;
        RECT 436.950 368.400 439.050 370.050 ;
        RECT 428.100 366.150 429.900 367.950 ;
        RECT 431.100 367.200 439.050 368.400 ;
        RECT 431.100 366.600 432.900 367.200 ;
        RECT 429.000 365.400 429.900 366.150 ;
        RECT 434.100 365.400 435.900 366.000 ;
        RECT 429.000 364.200 435.900 365.400 ;
        RECT 445.950 364.200 446.850 376.800 ;
        RECT 451.950 375.600 456.150 376.800 ;
        RECT 455.250 373.800 457.050 375.600 ;
        RECT 458.250 370.050 459.450 377.400 ;
        RECT 473.700 377.400 477.300 378.600 ;
        RECT 494.400 378.300 496.200 389.400 ;
        RECT 500.400 378.300 502.200 389.400 ;
        RECT 494.400 377.400 502.200 378.300 ;
        RECT 503.400 377.400 505.200 389.400 ;
        RECT 525.300 378.900 527.100 389.400 ;
        RECT 524.700 377.400 527.100 378.900 ;
        RECT 532.800 377.400 534.600 389.400 ;
        RECT 553.800 383.400 555.600 389.400 ;
        RECT 577.800 383.400 579.600 389.400 ;
        RECT 470.100 370.050 471.900 371.850 ;
        RECT 473.700 370.050 474.600 377.400 ;
        RECT 476.100 370.050 477.900 371.850 ;
        RECT 497.100 370.050 498.900 371.850 ;
        RECT 503.700 370.050 504.600 377.400 ;
        RECT 524.700 370.050 526.050 377.400 ;
        RECT 533.400 375.900 534.600 377.400 ;
        RECT 454.950 369.750 459.450 370.050 ;
        RECT 453.150 367.950 459.450 369.750 ;
        RECT 469.950 367.950 472.050 370.050 ;
        RECT 472.950 367.950 475.050 370.050 ;
        RECT 475.950 367.950 478.050 370.050 ;
        RECT 493.950 367.950 496.050 370.050 ;
        RECT 496.950 367.950 499.050 370.050 ;
        RECT 499.950 367.950 502.050 370.050 ;
        RECT 502.950 367.950 505.050 370.050 ;
        RECT 523.950 367.950 526.050 370.050 ;
        RECT 527.400 374.700 534.600 375.900 ;
        RECT 527.400 374.100 529.200 374.700 ;
        RECT 434.850 363.000 446.850 364.200 ;
        RECT 434.850 361.200 435.900 363.000 ;
        RECT 445.050 362.400 446.850 363.000 ;
        RECT 426.150 354.600 427.950 360.600 ;
        RECT 430.950 358.500 433.050 360.600 ;
        RECT 434.550 359.400 436.350 361.200 ;
        RECT 458.250 360.600 459.450 367.950 ;
        RECT 437.850 359.550 439.650 360.300 ;
        RECT 451.950 359.700 454.050 360.600 ;
        RECT 437.850 358.500 442.800 359.550 ;
        RECT 432.000 357.600 433.050 358.500 ;
        RECT 441.750 357.600 442.800 358.500 ;
        RECT 450.300 358.500 454.050 359.700 ;
        RECT 450.300 357.600 451.350 358.500 ;
        RECT 432.000 356.700 435.750 357.600 ;
        RECT 433.950 354.600 435.750 356.700 ;
        RECT 441.750 354.600 443.550 357.600 ;
        RECT 449.550 354.600 451.350 357.600 ;
        RECT 457.650 354.600 459.450 360.600 ;
        RECT 473.700 357.600 474.600 367.950 ;
        RECT 494.100 366.150 495.900 367.950 ;
        RECT 500.100 366.150 501.900 367.950 ;
        RECT 503.700 360.600 504.600 367.950 ;
        RECT 523.950 360.600 525.000 367.950 ;
        RECT 527.400 363.600 528.300 374.100 ;
        RECT 530.100 370.050 531.900 371.850 ;
        RECT 548.100 370.050 549.900 371.850 ;
        RECT 553.950 370.050 555.150 383.400 ;
        RECT 556.950 375.450 559.050 376.050 ;
        RECT 565.950 375.450 568.050 376.050 ;
        RECT 556.950 374.550 568.050 375.450 ;
        RECT 556.950 373.950 559.050 374.550 ;
        RECT 565.950 373.950 568.050 374.550 ;
        RECT 572.100 370.050 573.900 371.850 ;
        RECT 577.950 370.050 579.150 383.400 ;
        RECT 600.900 377.400 604.200 389.400 ;
        RECT 626.400 383.400 628.200 389.400 ;
        RECT 647.400 383.400 649.200 389.400 ;
        RECT 668.400 383.400 670.200 389.400 ;
        RECT 613.950 378.450 616.050 379.050 ;
        RECT 619.950 378.450 622.050 379.050 ;
        RECT 613.950 377.550 622.050 378.450 ;
        RECT 596.100 370.050 597.900 371.850 ;
        RECT 602.100 370.050 603.300 377.400 ;
        RECT 613.950 376.950 616.050 377.550 ;
        RECT 619.950 376.950 622.050 377.550 ;
        RECT 619.950 372.450 622.050 375.900 ;
        RECT 614.550 372.000 622.050 372.450 ;
        RECT 608.100 370.050 609.900 371.850 ;
        RECT 614.550 371.550 621.450 372.000 ;
        RECT 529.950 367.950 532.050 370.050 ;
        RECT 532.950 367.950 535.050 370.050 ;
        RECT 547.950 367.950 550.050 370.050 ;
        RECT 550.950 367.950 553.050 370.050 ;
        RECT 553.950 367.950 556.050 370.050 ;
        RECT 556.950 367.950 559.050 370.050 ;
        RECT 571.950 367.950 574.050 370.050 ;
        RECT 574.950 367.950 577.050 370.050 ;
        RECT 577.950 367.950 580.050 370.050 ;
        RECT 580.950 367.950 583.050 370.050 ;
        RECT 595.950 367.950 598.050 370.050 ;
        RECT 598.950 367.950 601.050 370.050 ;
        RECT 601.950 367.950 604.050 370.050 ;
        RECT 604.950 367.950 607.050 370.050 ;
        RECT 607.950 367.950 610.050 370.050 ;
        RECT 533.100 366.150 534.900 367.950 ;
        RECT 551.100 366.150 552.900 367.950 ;
        RECT 554.850 363.750 556.050 367.950 ;
        RECT 557.100 366.150 558.900 367.950 ;
        RECT 575.100 366.150 576.900 367.950 ;
        RECT 578.850 363.750 580.050 367.950 ;
        RECT 581.100 366.150 582.900 367.950 ;
        RECT 599.100 366.150 600.900 367.950 ;
        RECT 527.400 362.700 529.200 363.600 ;
        RECT 554.850 362.700 558.600 363.750 ;
        RECT 578.850 362.700 582.600 363.750 ;
        RECT 527.400 361.800 530.700 362.700 ;
        RECT 499.500 359.400 504.600 360.600 ;
        RECT 473.400 354.600 475.200 357.600 ;
        RECT 499.500 354.600 501.300 359.400 ;
        RECT 523.800 354.600 525.600 360.600 ;
        RECT 529.800 357.600 530.700 361.800 ;
        RECT 548.400 359.700 556.200 361.050 ;
        RECT 529.800 354.600 531.600 357.600 ;
        RECT 548.400 354.600 550.200 359.700 ;
        RECT 554.400 354.600 556.200 359.700 ;
        RECT 557.400 360.600 558.600 362.700 ;
        RECT 557.400 354.600 559.200 360.600 ;
        RECT 572.400 359.700 580.200 361.050 ;
        RECT 572.400 354.600 574.200 359.700 ;
        RECT 578.400 354.600 580.200 359.700 ;
        RECT 581.400 360.600 582.600 362.700 ;
        RECT 601.950 363.300 603.300 367.950 ;
        RECT 605.100 366.150 606.900 367.950 ;
        RECT 614.550 367.050 615.450 371.550 ;
        RECT 623.100 370.050 624.900 371.850 ;
        RECT 626.400 370.050 627.600 383.400 ;
        RECT 647.850 370.050 649.050 383.400 ;
        RECT 653.100 370.050 654.900 371.850 ;
        RECT 668.400 370.050 669.600 383.400 ;
        RECT 689.400 378.300 691.200 389.400 ;
        RECT 696.900 378.300 698.700 389.400 ;
        RECT 704.400 378.600 706.200 389.400 ;
        RECT 725.400 383.400 727.200 389.400 ;
        RECT 689.400 377.100 694.200 378.300 ;
        RECT 696.900 377.400 700.200 378.300 ;
        RECT 692.100 376.200 694.200 377.100 ;
        RECT 692.100 375.300 697.500 376.200 ;
        RECT 695.700 373.200 697.500 375.300 ;
        RECT 699.000 372.900 700.200 377.400 ;
        RECT 701.100 377.400 706.200 378.600 ;
        RECT 701.100 376.500 703.200 377.400 ;
        RECT 698.400 372.300 700.500 372.900 ;
        RECT 705.000 372.450 709.050 373.050 ;
        RECT 694.200 370.200 696.000 372.000 ;
        RECT 697.350 370.800 700.500 372.300 ;
        RECT 704.550 371.700 709.050 372.450 ;
        RECT 704.100 370.950 709.050 371.700 ;
        RECT 622.950 367.950 625.050 370.050 ;
        RECT 625.950 367.950 628.050 370.050 ;
        RECT 643.950 367.950 646.050 370.050 ;
        RECT 646.950 367.950 649.050 370.050 ;
        RECT 649.950 367.950 652.050 370.050 ;
        RECT 652.950 367.950 655.050 370.050 ;
        RECT 664.950 367.950 667.050 370.050 ;
        RECT 667.950 367.950 670.050 370.050 ;
        RECT 670.950 367.950 673.050 370.050 ;
        RECT 679.950 369.450 682.050 370.050 ;
        RECT 689.400 369.450 691.500 369.900 ;
        RECT 679.950 368.550 691.500 369.450 ;
        RECT 679.950 367.950 682.050 368.550 ;
        RECT 610.950 365.550 615.450 367.050 ;
        RECT 610.950 364.950 615.000 365.550 ;
        RECT 601.950 362.100 606.600 363.300 ;
        RECT 581.400 354.600 583.200 360.600 ;
        RECT 596.400 360.000 604.200 360.900 ;
        RECT 605.700 360.600 606.600 362.100 ;
        RECT 596.400 354.600 598.200 360.000 ;
        RECT 602.400 355.500 604.200 360.000 ;
        RECT 605.400 356.400 607.200 360.600 ;
        RECT 608.400 355.500 610.200 360.600 ;
        RECT 602.400 354.600 610.200 355.500 ;
        RECT 626.400 357.600 627.600 367.950 ;
        RECT 644.100 366.150 645.900 367.950 ;
        RECT 646.950 363.750 648.150 367.950 ;
        RECT 650.100 366.150 651.900 367.950 ;
        RECT 665.100 366.150 666.900 367.950 ;
        RECT 644.400 362.700 648.150 363.750 ;
        RECT 668.400 362.700 669.600 367.950 ;
        RECT 671.100 366.150 672.900 367.950 ;
        RECT 689.400 367.800 691.500 368.550 ;
        RECT 694.200 368.100 696.300 370.200 ;
        RECT 689.700 367.200 691.500 367.800 ;
        RECT 689.700 366.000 696.300 367.200 ;
        RECT 694.200 365.100 696.300 366.000 ;
        RECT 691.650 363.000 693.750 363.600 ;
        RECT 694.650 363.300 696.450 365.100 ;
        RECT 697.350 364.200 698.250 370.800 ;
        RECT 704.100 369.900 705.900 370.950 ;
        RECT 725.850 370.050 727.050 383.400 ;
        RECT 748.500 378.600 750.300 389.400 ;
        RECT 746.700 377.400 750.300 378.600 ;
        RECT 764.400 378.300 766.200 389.400 ;
        RECT 764.400 377.400 768.900 378.300 ;
        RECT 771.900 377.400 773.700 389.400 ;
        RECT 779.400 378.600 781.200 389.400 ;
        RECT 800.400 383.400 802.200 389.400 ;
        RECT 821.400 383.400 823.200 389.400 ;
        RECT 844.800 383.400 846.600 389.400 ;
        RECT 733.950 372.450 738.000 373.050 ;
        RECT 731.100 370.050 732.900 371.850 ;
        RECT 733.950 370.950 738.450 372.450 ;
        RECT 699.300 368.100 701.100 369.900 ;
        RECT 699.150 366.000 701.250 368.100 ;
        RECT 703.950 367.800 706.050 369.900 ;
        RECT 721.950 367.950 724.050 370.050 ;
        RECT 724.950 367.950 727.050 370.050 ;
        RECT 727.950 367.950 730.050 370.050 ;
        RECT 730.950 367.950 733.050 370.050 ;
        RECT 722.100 366.150 723.900 367.950 ;
        RECT 644.400 360.600 645.600 362.700 ;
        RECT 668.400 361.800 672.600 362.700 ;
        RECT 626.400 354.600 628.200 357.600 ;
        RECT 643.800 354.600 645.600 360.600 ;
        RECT 646.800 359.700 654.600 361.050 ;
        RECT 646.800 354.600 648.600 359.700 ;
        RECT 652.800 354.600 654.600 359.700 ;
        RECT 670.800 354.600 672.600 361.800 ;
        RECT 689.400 361.500 693.750 363.000 ;
        RECT 697.350 362.100 700.500 364.200 ;
        RECT 689.400 360.600 690.900 361.500 ;
        RECT 689.400 354.600 691.200 360.600 ;
        RECT 697.350 360.000 698.400 362.100 ;
        RECT 701.700 361.800 703.800 363.900 ;
        RECT 724.950 363.750 726.150 367.950 ;
        RECT 728.100 366.150 729.900 367.950 ;
        RECT 737.550 367.050 738.450 370.950 ;
        RECT 743.100 370.050 744.900 371.850 ;
        RECT 746.700 370.050 747.600 377.400 ;
        RECT 748.950 375.450 751.050 376.050 ;
        RECT 748.950 374.550 762.450 375.450 ;
        RECT 766.800 375.300 768.900 377.400 ;
        RECT 772.500 375.900 773.700 377.400 ;
        RECT 776.400 377.400 781.200 378.600 ;
        RECT 776.400 376.500 778.500 377.400 ;
        RECT 772.500 375.000 774.000 375.900 ;
        RECT 748.950 373.950 751.050 374.550 ;
        RECT 751.950 372.450 756.000 373.050 ;
        RECT 749.100 370.050 750.900 371.850 ;
        RECT 751.950 370.950 756.450 372.450 ;
        RECT 742.950 367.950 745.050 370.050 ;
        RECT 745.950 367.950 748.050 370.050 ;
        RECT 748.950 367.950 751.050 370.050 ;
        RECT 733.950 365.550 738.450 367.050 ;
        RECT 733.950 364.950 738.000 365.550 ;
        RECT 722.400 362.700 726.150 363.750 ;
        RECT 701.700 360.600 706.200 361.800 ;
        RECT 722.400 360.600 723.600 362.700 ;
        RECT 696.600 354.600 698.400 360.000 ;
        RECT 704.400 354.600 706.200 360.600 ;
        RECT 721.800 354.600 723.600 360.600 ;
        RECT 724.800 359.700 732.600 361.050 ;
        RECT 724.800 354.600 726.600 359.700 ;
        RECT 730.800 354.600 732.600 359.700 ;
        RECT 746.700 357.600 747.600 367.950 ;
        RECT 755.550 367.050 756.450 370.950 ;
        RECT 761.550 369.450 762.450 374.550 ;
        RECT 770.100 373.500 772.200 373.800 ;
        RECT 768.300 371.700 772.200 373.500 ;
        RECT 773.100 372.900 774.000 375.000 ;
        RECT 773.100 370.800 775.200 372.900 ;
        RECT 764.400 369.900 766.500 370.050 ;
        RECT 769.500 369.900 771.300 370.500 ;
        RECT 764.400 369.450 771.300 369.900 ;
        RECT 761.550 368.700 771.300 369.450 ;
        RECT 772.200 369.900 774.600 370.800 ;
        RECT 779.100 370.050 780.900 371.850 ;
        RECT 800.850 370.050 802.050 383.400 ;
        RECT 808.950 375.450 811.050 376.050 ;
        RECT 817.950 375.450 820.050 376.050 ;
        RECT 808.950 374.550 820.050 375.450 ;
        RECT 808.950 373.950 811.050 374.550 ;
        RECT 817.950 373.950 820.050 374.550 ;
        RECT 809.550 372.450 810.450 373.950 ;
        RECT 806.100 370.050 807.900 371.850 ;
        RECT 809.550 371.550 813.450 372.450 ;
        RECT 761.550 368.550 766.500 368.700 ;
        RECT 751.950 365.550 756.450 367.050 ;
        RECT 764.400 367.950 766.500 368.550 ;
        RECT 764.400 366.150 766.200 367.950 ;
        RECT 751.950 364.950 756.000 365.550 ;
        RECT 769.500 365.400 771.300 367.200 ;
        RECT 769.200 363.300 771.300 365.400 ;
        RECT 765.000 362.400 771.300 363.300 ;
        RECT 772.200 364.200 773.250 369.900 ;
        RECT 778.950 369.450 781.050 370.050 ;
        RECT 787.950 369.450 790.050 370.050 ;
        RECT 774.600 367.200 776.400 369.000 ;
        RECT 778.950 368.550 790.050 369.450 ;
        RECT 778.950 367.950 781.050 368.550 ;
        RECT 787.950 367.950 790.050 368.550 ;
        RECT 796.950 367.950 799.050 370.050 ;
        RECT 799.950 367.950 802.050 370.050 ;
        RECT 802.950 367.950 805.050 370.050 ;
        RECT 805.950 367.950 808.050 370.050 ;
        RECT 774.150 365.100 776.250 367.200 ;
        RECT 797.100 366.150 798.900 367.950 ;
        RECT 765.000 360.600 766.200 362.400 ;
        RECT 772.200 362.100 775.200 364.200 ;
        RECT 799.950 363.750 801.150 367.950 ;
        RECT 803.100 366.150 804.900 367.950 ;
        RECT 812.550 367.050 813.450 371.550 ;
        RECT 821.400 370.050 822.600 383.400 ;
        RECT 839.100 370.050 840.900 371.850 ;
        RECT 844.950 370.050 846.150 383.400 ;
        RECT 863.400 378.300 865.200 389.400 ;
        RECT 869.400 378.300 871.200 389.400 ;
        RECT 863.400 377.400 871.200 378.300 ;
        RECT 872.400 377.400 874.200 389.400 ;
        RECT 847.950 375.450 850.050 376.050 ;
        RECT 868.950 375.450 871.050 376.050 ;
        RECT 847.950 374.550 871.050 375.450 ;
        RECT 847.950 373.950 850.050 374.550 ;
        RECT 868.950 373.950 871.050 374.550 ;
        RECT 866.100 370.050 867.900 371.850 ;
        RECT 872.700 370.050 873.600 377.400 ;
        RECT 817.950 367.950 820.050 370.050 ;
        RECT 820.950 367.950 823.050 370.050 ;
        RECT 823.950 367.950 826.050 370.050 ;
        RECT 838.950 367.950 841.050 370.050 ;
        RECT 841.950 367.950 844.050 370.050 ;
        RECT 844.950 367.950 847.050 370.050 ;
        RECT 847.950 367.950 850.050 370.050 ;
        RECT 862.950 367.950 865.050 370.050 ;
        RECT 865.950 367.950 868.050 370.050 ;
        RECT 868.950 367.950 871.050 370.050 ;
        RECT 871.950 367.950 874.050 370.050 ;
        RECT 812.550 365.550 817.050 367.050 ;
        RECT 818.100 366.150 819.900 367.950 ;
        RECT 813.000 364.950 817.050 365.550 ;
        RECT 797.400 362.700 801.150 363.750 ;
        RECT 821.400 362.700 822.600 367.950 ;
        RECT 824.100 366.150 825.900 367.950 ;
        RECT 842.100 366.150 843.900 367.950 ;
        RECT 845.850 363.750 847.050 367.950 ;
        RECT 848.100 366.150 849.900 367.950 ;
        RECT 863.100 366.150 864.900 367.950 ;
        RECT 869.100 366.150 870.900 367.950 ;
        RECT 845.850 362.700 849.600 363.750 ;
        RECT 772.200 360.600 773.400 362.100 ;
        RECT 776.400 361.500 778.500 362.700 ;
        RECT 776.400 360.600 781.200 361.500 ;
        RECT 797.400 360.600 798.600 362.700 ;
        RECT 821.400 361.800 825.600 362.700 ;
        RECT 746.400 354.600 748.200 357.600 ;
        RECT 764.400 354.600 766.200 360.600 ;
        RECT 771.900 354.600 773.700 360.600 ;
        RECT 779.400 354.600 781.200 360.600 ;
        RECT 796.800 354.600 798.600 360.600 ;
        RECT 799.800 359.700 807.600 361.050 ;
        RECT 799.800 354.600 801.600 359.700 ;
        RECT 805.800 354.600 807.600 359.700 ;
        RECT 823.800 354.600 825.600 361.800 ;
        RECT 839.400 359.700 847.200 361.050 ;
        RECT 839.400 354.600 841.200 359.700 ;
        RECT 845.400 354.600 847.200 359.700 ;
        RECT 848.400 360.600 849.600 362.700 ;
        RECT 872.700 360.600 873.600 367.950 ;
        RECT 848.400 354.600 850.200 360.600 ;
        RECT 868.500 359.400 873.600 360.600 ;
        RECT 868.500 354.600 870.300 359.400 ;
        RECT 3.150 344.400 4.950 350.400 ;
        RECT 10.950 348.300 12.750 350.400 ;
        RECT 9.000 347.400 12.750 348.300 ;
        RECT 18.750 347.400 20.550 350.400 ;
        RECT 26.550 347.400 28.350 350.400 ;
        RECT 9.000 346.500 10.050 347.400 ;
        RECT 18.750 346.500 19.800 347.400 ;
        RECT 7.950 344.400 10.050 346.500 ;
        RECT 3.150 329.700 4.050 344.400 ;
        RECT 11.550 343.800 13.350 345.600 ;
        RECT 14.850 345.450 19.800 346.500 ;
        RECT 27.300 346.500 28.350 347.400 ;
        RECT 14.850 344.700 16.650 345.450 ;
        RECT 27.300 345.300 31.050 346.500 ;
        RECT 28.950 344.400 31.050 345.300 ;
        RECT 34.650 344.400 36.450 350.400 ;
        RECT 11.850 342.000 12.900 343.800 ;
        RECT 22.050 342.000 23.850 342.600 ;
        RECT 11.850 340.800 23.850 342.000 ;
        RECT 6.000 339.600 12.900 340.800 ;
        RECT 6.000 338.850 6.900 339.600 ;
        RECT 11.100 339.000 12.900 339.600 ;
        RECT 5.100 337.050 6.900 338.850 ;
        RECT 8.100 337.800 9.900 338.400 ;
        RECT 4.950 334.950 7.050 337.050 ;
        RECT 8.100 336.600 16.050 337.800 ;
        RECT 13.950 334.950 16.050 336.600 ;
        RECT 12.450 329.700 14.250 330.000 ;
        RECT 3.150 329.100 14.250 329.700 ;
        RECT 3.150 328.500 20.850 329.100 ;
        RECT 3.150 327.600 4.050 328.500 ;
        RECT 12.450 328.200 20.850 328.500 ;
        RECT 3.150 315.600 4.950 327.600 ;
        RECT 17.250 326.700 19.050 327.300 ;
        RECT 11.550 325.500 19.050 326.700 ;
        RECT 19.950 326.100 20.850 328.200 ;
        RECT 22.950 328.200 23.850 340.800 ;
        RECT 35.250 337.050 36.450 344.400 ;
        RECT 52.800 343.200 54.600 350.400 ;
        RECT 50.400 342.300 54.600 343.200 ;
        RECT 81.000 344.400 82.800 350.400 ;
        RECT 47.100 337.050 48.900 338.850 ;
        RECT 50.400 337.050 51.600 342.300 ;
        RECT 53.100 337.050 54.900 338.850 ;
        RECT 74.100 337.050 75.900 338.850 ;
        RECT 81.000 337.050 82.050 344.400 ;
        RECT 106.800 343.200 108.600 350.400 ;
        RECT 124.800 344.400 126.600 350.400 ;
        RECT 104.400 342.300 108.600 343.200 ;
        RECT 125.400 342.300 126.600 344.400 ;
        RECT 127.800 345.300 129.600 350.400 ;
        RECT 133.800 345.300 135.600 350.400 ;
        RECT 127.800 343.950 135.600 345.300 ;
        RECT 149.400 343.200 151.200 350.400 ;
        RECT 170.400 343.200 172.200 350.400 ;
        RECT 191.400 347.400 193.200 350.400 ;
        RECT 206.400 347.400 208.200 350.400 ;
        RECT 149.400 342.300 153.600 343.200 ;
        RECT 170.400 342.300 174.600 343.200 ;
        RECT 86.100 337.050 87.900 338.850 ;
        RECT 101.100 337.050 102.900 338.850 ;
        RECT 104.400 337.050 105.600 342.300 ;
        RECT 125.400 341.250 129.150 342.300 ;
        RECT 112.950 339.450 115.050 340.050 ;
        RECT 121.950 339.450 124.050 340.050 ;
        RECT 107.100 337.050 108.900 338.850 ;
        RECT 112.950 338.550 124.050 339.450 ;
        RECT 112.950 337.950 115.050 338.550 ;
        RECT 121.950 337.950 124.050 338.550 ;
        RECT 125.100 337.050 126.900 338.850 ;
        RECT 127.950 337.050 129.150 341.250 ;
        RECT 131.100 337.050 132.900 338.850 ;
        RECT 149.100 337.050 150.900 338.850 ;
        RECT 152.400 337.050 153.600 342.300 ;
        RECT 155.100 337.050 156.900 338.850 ;
        RECT 170.100 337.050 171.900 338.850 ;
        RECT 173.400 337.050 174.600 342.300 ;
        RECT 176.100 337.050 177.900 338.850 ;
        RECT 191.400 337.050 192.600 347.400 ;
        RECT 206.400 343.500 207.600 347.400 ;
        RECT 212.400 344.400 214.200 350.400 ;
        RECT 232.800 347.400 234.600 350.400 ;
        RECT 206.400 342.600 212.100 343.500 ;
        RECT 210.150 341.700 212.100 342.600 ;
        RECT 30.150 335.250 36.450 337.050 ;
        RECT 31.950 334.950 36.450 335.250 ;
        RECT 46.950 334.950 49.050 337.050 ;
        RECT 49.950 334.950 52.050 337.050 ;
        RECT 52.950 334.950 55.050 337.050 ;
        RECT 73.950 334.950 76.050 337.050 ;
        RECT 76.950 334.950 79.050 337.050 ;
        RECT 79.950 334.950 82.050 337.050 ;
        RECT 82.950 334.950 85.050 337.050 ;
        RECT 85.950 334.950 88.050 337.050 ;
        RECT 100.950 334.950 103.050 337.050 ;
        RECT 103.950 334.950 106.050 337.050 ;
        RECT 106.950 334.950 109.050 337.050 ;
        RECT 124.950 334.950 127.050 337.050 ;
        RECT 127.950 334.950 130.050 337.050 ;
        RECT 130.950 334.950 133.050 337.050 ;
        RECT 133.950 334.950 136.050 337.050 ;
        RECT 148.950 334.950 151.050 337.050 ;
        RECT 151.950 334.950 154.050 337.050 ;
        RECT 154.950 334.950 157.050 337.050 ;
        RECT 169.950 334.950 172.050 337.050 ;
        RECT 172.950 334.950 175.050 337.050 ;
        RECT 175.950 334.950 178.050 337.050 ;
        RECT 187.950 334.950 190.050 337.050 ;
        RECT 190.950 334.950 193.050 337.050 ;
        RECT 205.950 334.950 208.050 337.050 ;
        RECT 32.250 329.400 34.050 331.200 ;
        RECT 28.950 328.200 33.150 329.400 ;
        RECT 22.950 327.300 28.050 328.200 ;
        RECT 28.950 327.300 31.050 328.200 ;
        RECT 35.250 327.600 36.450 334.950 ;
        RECT 27.150 326.400 28.050 327.300 ;
        RECT 24.450 326.100 26.250 326.400 ;
        RECT 11.550 324.600 12.750 325.500 ;
        RECT 19.950 325.200 26.250 326.100 ;
        RECT 24.450 324.600 26.250 325.200 ;
        RECT 27.150 324.600 29.850 326.400 ;
        RECT 7.950 322.500 12.750 324.600 ;
        RECT 15.450 323.550 17.250 324.300 ;
        RECT 20.250 323.550 22.050 324.300 ;
        RECT 15.450 322.500 22.050 323.550 ;
        RECT 11.550 321.600 12.750 322.500 ;
        RECT 11.550 315.600 13.350 321.600 ;
        RECT 19.350 315.600 21.150 322.500 ;
        RECT 27.150 321.600 31.050 323.700 ;
        RECT 27.150 315.600 28.950 321.600 ;
        RECT 34.650 315.600 36.450 327.600 ;
        RECT 50.400 321.600 51.600 334.950 ;
        RECT 77.100 333.150 78.900 334.950 ;
        RECT 81.000 329.400 81.900 334.950 ;
        RECT 83.100 333.150 84.900 334.950 ;
        RECT 76.800 328.500 81.900 329.400 ;
        RECT 50.400 315.600 52.200 321.600 ;
        RECT 73.800 316.500 75.600 327.600 ;
        RECT 76.800 317.400 78.600 328.500 ;
        RECT 79.800 326.400 87.600 327.300 ;
        RECT 79.800 316.500 81.600 326.400 ;
        RECT 73.800 315.600 81.600 316.500 ;
        RECT 85.800 315.600 87.600 326.400 ;
        RECT 104.400 321.600 105.600 334.950 ;
        RECT 128.850 321.600 130.050 334.950 ;
        RECT 134.100 333.150 135.900 334.950 ;
        RECT 152.400 321.600 153.600 334.950 ;
        RECT 160.950 330.450 163.050 331.050 ;
        RECT 169.950 330.450 172.050 331.050 ;
        RECT 160.950 329.550 172.050 330.450 ;
        RECT 160.950 328.950 163.050 329.550 ;
        RECT 169.950 328.950 172.050 329.550 ;
        RECT 173.400 321.600 174.600 334.950 ;
        RECT 188.100 333.150 189.900 334.950 ;
        RECT 104.400 315.600 106.200 321.600 ;
        RECT 128.400 315.600 130.200 321.600 ;
        RECT 151.800 315.600 153.600 321.600 ;
        RECT 172.800 315.600 174.600 321.600 ;
        RECT 191.400 321.600 192.600 334.950 ;
        RECT 206.100 333.150 207.900 334.950 ;
        RECT 210.150 330.300 211.050 341.700 ;
        RECT 213.000 337.050 214.200 344.400 ;
        RECT 233.400 337.050 234.300 347.400 ;
        RECT 253.500 345.600 255.300 350.400 ;
        RECT 275.400 347.400 277.200 350.400 ;
        RECT 253.500 344.400 258.600 345.600 ;
        RECT 248.100 337.050 249.900 338.850 ;
        RECT 254.100 337.050 255.900 338.850 ;
        RECT 257.700 337.050 258.600 344.400 ;
        RECT 275.700 337.050 276.600 347.400 ;
        RECT 285.150 344.400 286.950 350.400 ;
        RECT 292.950 348.300 294.750 350.400 ;
        RECT 291.000 347.400 294.750 348.300 ;
        RECT 300.750 347.400 302.550 350.400 ;
        RECT 308.550 347.400 310.350 350.400 ;
        RECT 291.000 346.500 292.050 347.400 ;
        RECT 300.750 346.500 301.800 347.400 ;
        RECT 289.950 344.400 292.050 346.500 ;
        RECT 211.950 334.950 214.200 337.050 ;
        RECT 229.950 334.950 232.050 337.050 ;
        RECT 232.950 334.950 235.050 337.050 ;
        RECT 235.950 334.950 238.050 337.050 ;
        RECT 247.950 334.950 250.050 337.050 ;
        RECT 250.950 334.950 253.050 337.050 ;
        RECT 253.950 334.950 256.050 337.050 ;
        RECT 256.950 334.950 259.050 337.050 ;
        RECT 271.950 334.950 274.050 337.050 ;
        RECT 274.950 334.950 277.050 337.050 ;
        RECT 277.950 334.950 280.050 337.050 ;
        RECT 210.150 329.400 212.100 330.300 ;
        RECT 206.400 328.500 212.100 329.400 ;
        RECT 206.400 321.600 207.600 328.500 ;
        RECT 213.000 327.600 214.200 334.950 ;
        RECT 230.100 333.150 231.900 334.950 ;
        RECT 233.400 327.600 234.300 334.950 ;
        RECT 236.100 333.150 237.900 334.950 ;
        RECT 251.100 333.150 252.900 334.950 ;
        RECT 257.700 327.600 258.600 334.950 ;
        RECT 272.100 333.150 273.900 334.950 ;
        RECT 275.700 327.600 276.600 334.950 ;
        RECT 278.100 333.150 279.900 334.950 ;
        RECT 285.150 329.700 286.050 344.400 ;
        RECT 293.550 343.800 295.350 345.600 ;
        RECT 296.850 345.450 301.800 346.500 ;
        RECT 309.300 346.500 310.350 347.400 ;
        RECT 296.850 344.700 298.650 345.450 ;
        RECT 309.300 345.300 313.050 346.500 ;
        RECT 310.950 344.400 313.050 345.300 ;
        RECT 316.650 344.400 318.450 350.400 ;
        RECT 293.850 342.000 294.900 343.800 ;
        RECT 304.050 342.000 305.850 342.600 ;
        RECT 293.850 340.800 305.850 342.000 ;
        RECT 288.000 339.600 294.900 340.800 ;
        RECT 288.000 338.850 288.900 339.600 ;
        RECT 293.100 339.000 294.900 339.600 ;
        RECT 287.100 337.050 288.900 338.850 ;
        RECT 290.100 337.800 291.900 338.400 ;
        RECT 286.950 334.950 289.050 337.050 ;
        RECT 290.100 336.600 298.050 337.800 ;
        RECT 295.950 334.950 298.050 336.600 ;
        RECT 294.450 329.700 296.250 330.000 ;
        RECT 285.150 329.100 296.250 329.700 ;
        RECT 285.150 328.500 302.850 329.100 ;
        RECT 285.150 327.600 286.050 328.500 ;
        RECT 294.450 328.200 302.850 328.500 ;
        RECT 191.400 315.600 193.200 321.600 ;
        RECT 206.400 315.600 208.200 321.600 ;
        RECT 212.400 315.600 214.200 327.600 ;
        RECT 230.700 326.400 234.300 327.600 ;
        RECT 248.400 326.700 256.200 327.600 ;
        RECT 230.700 315.600 232.500 326.400 ;
        RECT 248.400 315.600 250.200 326.700 ;
        RECT 254.400 315.600 256.200 326.700 ;
        RECT 257.400 315.600 259.200 327.600 ;
        RECT 275.700 326.400 279.300 327.600 ;
        RECT 277.500 315.600 279.300 326.400 ;
        RECT 285.150 315.600 286.950 327.600 ;
        RECT 299.250 326.700 301.050 327.300 ;
        RECT 293.550 325.500 301.050 326.700 ;
        RECT 301.950 326.100 302.850 328.200 ;
        RECT 304.950 328.200 305.850 340.800 ;
        RECT 317.250 337.050 318.450 344.400 ;
        RECT 332.400 347.400 334.200 350.400 ;
        RECT 332.400 337.050 333.600 347.400 ;
        RECT 350.400 343.500 352.200 350.400 ;
        RECT 356.400 343.500 358.200 350.400 ;
        RECT 362.400 343.500 364.200 350.400 ;
        RECT 368.400 343.500 370.200 350.400 ;
        RECT 391.800 347.400 393.600 350.400 ;
        RECT 350.400 342.300 354.300 343.500 ;
        RECT 356.400 342.300 360.300 343.500 ;
        RECT 362.400 342.300 366.300 343.500 ;
        RECT 368.400 342.300 371.100 343.500 ;
        RECT 353.100 341.400 354.300 342.300 ;
        RECT 359.100 341.400 360.300 342.300 ;
        RECT 365.100 341.400 366.300 342.300 ;
        RECT 353.100 340.200 357.300 341.400 ;
        RECT 350.100 337.050 351.900 338.850 ;
        RECT 312.150 335.250 318.450 337.050 ;
        RECT 313.950 334.950 318.450 335.250 ;
        RECT 328.950 334.950 331.050 337.050 ;
        RECT 331.950 334.950 334.050 337.050 ;
        RECT 349.950 334.950 352.050 337.050 ;
        RECT 314.250 329.400 316.050 331.200 ;
        RECT 310.950 328.200 315.150 329.400 ;
        RECT 304.950 327.300 310.050 328.200 ;
        RECT 310.950 327.300 313.050 328.200 ;
        RECT 317.250 327.600 318.450 334.950 ;
        RECT 329.100 333.150 330.900 334.950 ;
        RECT 309.150 326.400 310.050 327.300 ;
        RECT 306.450 326.100 308.250 326.400 ;
        RECT 293.550 324.600 294.750 325.500 ;
        RECT 301.950 325.200 308.250 326.100 ;
        RECT 306.450 324.600 308.250 325.200 ;
        RECT 309.150 324.600 311.850 326.400 ;
        RECT 289.950 322.500 294.750 324.600 ;
        RECT 297.450 323.550 299.250 324.300 ;
        RECT 302.250 323.550 304.050 324.300 ;
        RECT 297.450 322.500 304.050 323.550 ;
        RECT 293.550 321.600 294.750 322.500 ;
        RECT 293.550 315.600 295.350 321.600 ;
        RECT 301.350 315.600 303.150 322.500 ;
        RECT 309.150 321.600 313.050 323.700 ;
        RECT 309.150 315.600 310.950 321.600 ;
        RECT 316.650 315.600 318.450 327.600 ;
        RECT 332.400 321.600 333.600 334.950 ;
        RECT 353.100 329.700 354.300 340.200 ;
        RECT 355.500 339.600 357.300 340.200 ;
        RECT 359.100 340.200 363.300 341.400 ;
        RECT 359.100 329.700 360.300 340.200 ;
        RECT 361.500 339.600 363.300 340.200 ;
        RECT 365.100 340.200 369.300 341.400 ;
        RECT 365.100 329.700 366.300 340.200 ;
        RECT 367.500 339.600 369.300 340.200 ;
        RECT 370.200 337.050 371.100 342.300 ;
        RECT 392.400 337.050 393.300 347.400 ;
        RECT 413.700 345.600 415.500 350.400 ;
        RECT 410.400 344.400 415.500 345.600 ;
        RECT 433.800 344.400 435.600 350.400 ;
        RECT 439.800 347.400 441.600 350.400 ;
        RECT 410.400 337.050 411.300 344.400 ;
        RECT 413.100 337.050 414.900 338.850 ;
        RECT 419.100 337.050 420.900 338.850 ;
        RECT 433.800 337.050 435.000 344.400 ;
        RECT 440.400 343.500 441.600 347.400 ;
        RECT 435.900 342.600 441.600 343.500 ;
        RECT 452.400 347.400 454.200 350.400 ;
        RECT 452.400 343.500 453.600 347.400 ;
        RECT 458.400 344.400 460.200 350.400 ;
        RECT 478.800 347.400 480.600 350.400 ;
        RECT 452.400 342.600 458.100 343.500 ;
        RECT 435.900 341.700 437.850 342.600 ;
        RECT 370.200 334.950 373.050 337.050 ;
        RECT 388.950 334.950 391.050 337.050 ;
        RECT 391.950 334.950 394.050 337.050 ;
        RECT 394.950 334.950 397.050 337.050 ;
        RECT 409.950 334.950 412.050 337.050 ;
        RECT 412.950 334.950 415.050 337.050 ;
        RECT 415.950 334.950 418.050 337.050 ;
        RECT 418.950 334.950 421.050 337.050 ;
        RECT 433.800 334.950 436.050 337.050 ;
        RECT 370.200 329.700 371.100 334.950 ;
        RECT 389.100 333.150 390.900 334.950 ;
        RECT 350.400 328.500 354.300 329.700 ;
        RECT 356.400 328.500 360.300 329.700 ;
        RECT 362.400 328.500 366.300 329.700 ;
        RECT 368.400 328.500 371.100 329.700 ;
        RECT 332.400 315.600 334.200 321.600 ;
        RECT 350.400 315.600 352.200 328.500 ;
        RECT 356.400 315.600 358.200 328.500 ;
        RECT 362.400 315.600 364.200 328.500 ;
        RECT 368.400 315.600 370.200 328.500 ;
        RECT 392.400 327.600 393.300 334.950 ;
        RECT 395.100 333.150 396.900 334.950 ;
        RECT 410.400 327.600 411.300 334.950 ;
        RECT 416.100 333.150 417.900 334.950 ;
        RECT 433.800 327.600 435.000 334.950 ;
        RECT 436.950 330.300 437.850 341.700 ;
        RECT 456.150 341.700 458.100 342.600 ;
        RECT 439.950 334.950 442.050 337.050 ;
        RECT 451.950 334.950 454.050 337.050 ;
        RECT 440.100 333.150 441.900 334.950 ;
        RECT 452.100 333.150 453.900 334.950 ;
        RECT 435.900 329.400 437.850 330.300 ;
        RECT 456.150 330.300 457.050 341.700 ;
        RECT 459.000 337.050 460.200 344.400 ;
        RECT 479.400 337.050 480.300 347.400 ;
        RECT 481.950 342.450 484.050 343.050 ;
        RECT 490.950 342.450 493.050 343.050 ;
        RECT 481.950 341.550 493.050 342.450 ;
        RECT 481.950 340.950 484.050 341.550 ;
        RECT 490.950 340.950 493.050 341.550 ;
        RECT 501.000 342.000 502.800 350.400 ;
        RECT 518.400 345.300 520.200 350.400 ;
        RECT 524.400 345.300 526.200 350.400 ;
        RECT 518.400 343.950 526.200 345.300 ;
        RECT 527.400 344.400 529.200 350.400 ;
        RECT 542.400 345.300 544.200 350.400 ;
        RECT 548.400 345.300 550.200 350.400 ;
        RECT 527.400 342.300 528.600 344.400 ;
        RECT 542.400 343.950 550.200 345.300 ;
        RECT 551.400 344.400 553.200 350.400 ;
        RECT 551.400 342.300 552.600 344.400 ;
        RECT 569.400 343.200 571.200 350.400 ;
        RECT 590.400 344.400 592.200 350.400 ;
        RECT 597.900 344.400 599.700 350.400 ;
        RECT 605.400 344.400 607.200 350.400 ;
        RECT 622.800 344.400 624.600 350.400 ;
        RECT 569.400 342.300 573.600 343.200 ;
        RECT 501.000 340.800 504.300 342.000 ;
        RECT 494.100 337.050 495.900 338.850 ;
        RECT 500.100 337.050 501.900 338.850 ;
        RECT 503.400 337.050 504.300 340.800 ;
        RECT 524.850 341.250 528.600 342.300 ;
        RECT 548.850 341.250 552.600 342.300 ;
        RECT 513.000 339.450 517.050 340.050 ;
        RECT 512.550 337.950 517.050 339.450 ;
        RECT 457.950 334.950 460.200 337.050 ;
        RECT 475.950 334.950 478.050 337.050 ;
        RECT 478.950 334.950 481.050 337.050 ;
        RECT 481.950 334.950 484.050 337.050 ;
        RECT 493.950 334.950 496.050 337.050 ;
        RECT 496.950 334.950 499.050 337.050 ;
        RECT 499.950 334.950 502.050 337.050 ;
        RECT 502.950 334.950 505.050 337.050 ;
        RECT 456.150 329.400 458.100 330.300 ;
        RECT 435.900 328.500 441.600 329.400 ;
        RECT 389.700 326.400 393.300 327.600 ;
        RECT 389.700 315.600 391.500 326.400 ;
        RECT 409.800 315.600 411.600 327.600 ;
        RECT 412.800 326.700 420.600 327.600 ;
        RECT 412.800 315.600 414.600 326.700 ;
        RECT 418.800 315.600 420.600 326.700 ;
        RECT 433.800 315.600 435.600 327.600 ;
        RECT 440.400 321.600 441.600 328.500 ;
        RECT 439.800 315.600 441.600 321.600 ;
        RECT 452.400 328.500 458.100 329.400 ;
        RECT 452.400 321.600 453.600 328.500 ;
        RECT 459.000 327.600 460.200 334.950 ;
        RECT 476.100 333.150 477.900 334.950 ;
        RECT 479.400 327.600 480.300 334.950 ;
        RECT 482.100 333.150 483.900 334.950 ;
        RECT 497.100 333.150 498.900 334.950 ;
        RECT 452.400 315.600 454.200 321.600 ;
        RECT 458.400 315.600 460.200 327.600 ;
        RECT 476.700 326.400 480.300 327.600 ;
        RECT 476.700 315.600 478.500 326.400 ;
        RECT 503.400 322.800 504.300 334.950 ;
        RECT 512.550 334.050 513.450 337.950 ;
        RECT 521.100 337.050 522.900 338.850 ;
        RECT 524.850 337.050 526.050 341.250 ;
        RECT 527.100 337.050 528.900 338.850 ;
        RECT 545.100 337.050 546.900 338.850 ;
        RECT 548.850 337.050 550.050 341.250 ;
        RECT 553.950 339.450 558.000 340.050 ;
        RECT 551.100 337.050 552.900 338.850 ;
        RECT 553.950 337.950 558.450 339.450 ;
        RECT 517.950 334.950 520.050 337.050 ;
        RECT 520.950 334.950 523.050 337.050 ;
        RECT 523.950 334.950 526.050 337.050 ;
        RECT 526.950 334.950 529.050 337.050 ;
        RECT 541.950 334.950 544.050 337.050 ;
        RECT 544.950 334.950 547.050 337.050 ;
        RECT 547.950 334.950 550.050 337.050 ;
        RECT 550.950 334.950 553.050 337.050 ;
        RECT 512.550 332.550 517.050 334.050 ;
        RECT 518.100 333.150 519.900 334.950 ;
        RECT 513.000 331.950 517.050 332.550 ;
        RECT 497.700 321.900 504.300 322.800 ;
        RECT 497.700 321.600 499.200 321.900 ;
        RECT 497.400 315.600 499.200 321.600 ;
        RECT 503.400 321.600 504.300 321.900 ;
        RECT 523.950 321.600 525.150 334.950 ;
        RECT 542.100 333.150 543.900 334.950 ;
        RECT 526.950 330.450 529.050 331.050 ;
        RECT 541.950 330.450 544.050 331.050 ;
        RECT 526.950 329.550 544.050 330.450 ;
        RECT 526.950 328.950 529.050 329.550 ;
        RECT 541.950 328.950 544.050 329.550 ;
        RECT 532.950 327.900 537.000 328.050 ;
        RECT 532.950 325.950 538.050 327.900 ;
        RECT 535.950 325.800 538.050 325.950 ;
        RECT 547.950 321.600 549.150 334.950 ;
        RECT 557.550 330.900 558.450 337.950 ;
        RECT 569.100 337.050 570.900 338.850 ;
        RECT 572.400 337.050 573.600 342.300 ;
        RECT 591.000 342.600 592.200 344.400 ;
        RECT 598.200 342.900 599.400 344.400 ;
        RECT 602.400 343.500 607.200 344.400 ;
        RECT 591.000 341.700 597.300 342.600 ;
        RECT 577.950 339.450 580.050 340.050 ;
        RECT 595.200 339.600 597.300 341.700 ;
        RECT 577.950 338.850 591.450 339.450 ;
        RECT 575.100 337.050 576.900 338.850 ;
        RECT 577.950 338.550 592.200 338.850 ;
        RECT 577.950 337.950 580.050 338.550 ;
        RECT 590.400 337.050 592.200 338.550 ;
        RECT 595.500 337.800 597.300 339.600 ;
        RECT 598.200 340.800 601.200 342.900 ;
        RECT 602.400 342.300 604.500 343.500 ;
        RECT 623.400 342.300 624.600 344.400 ;
        RECT 625.800 345.300 627.600 350.400 ;
        RECT 631.800 345.300 633.600 350.400 ;
        RECT 625.800 343.950 633.600 345.300 ;
        RECT 623.400 341.250 627.150 342.300 ;
        RECT 649.200 342.000 651.000 350.400 ;
        RECT 673.500 345.600 675.300 350.400 ;
        RECT 673.500 344.400 678.600 345.600 ;
        RECT 568.950 334.950 571.050 337.050 ;
        RECT 571.950 334.950 574.050 337.050 ;
        RECT 574.950 334.950 577.050 337.050 ;
        RECT 590.400 336.300 592.500 337.050 ;
        RECT 590.400 335.100 597.300 336.300 ;
        RECT 590.400 334.950 592.500 335.100 ;
        RECT 556.950 328.800 559.050 330.900 ;
        RECT 572.400 321.600 573.600 334.950 ;
        RECT 595.500 334.500 597.300 335.100 ;
        RECT 598.200 335.100 599.250 340.800 ;
        RECT 600.150 337.800 602.250 339.900 ;
        RECT 600.600 336.000 602.400 337.800 ;
        RECT 623.100 337.050 624.900 338.850 ;
        RECT 625.950 337.050 627.150 341.250 ;
        RECT 647.700 340.800 651.000 342.000 ;
        RECT 629.100 337.050 630.900 338.850 ;
        RECT 647.700 337.050 648.600 340.800 ;
        RECT 658.950 339.450 663.000 340.050 ;
        RECT 650.100 337.050 651.900 338.850 ;
        RECT 656.100 337.050 657.900 338.850 ;
        RECT 658.950 337.950 663.450 339.450 ;
        RECT 604.950 336.450 607.050 337.050 ;
        RECT 609.000 336.450 613.050 337.050 ;
        RECT 604.950 335.550 613.050 336.450 ;
        RECT 598.200 334.200 600.600 335.100 ;
        RECT 604.950 334.950 607.050 335.550 ;
        RECT 609.000 334.950 613.050 335.550 ;
        RECT 622.950 334.950 625.050 337.050 ;
        RECT 625.950 334.950 628.050 337.050 ;
        RECT 628.950 334.950 631.050 337.050 ;
        RECT 631.950 334.950 634.050 337.050 ;
        RECT 646.950 334.950 649.050 337.050 ;
        RECT 649.950 334.950 652.050 337.050 ;
        RECT 652.950 334.950 655.050 337.050 ;
        RECT 655.950 334.950 658.050 337.050 ;
        RECT 594.300 331.500 598.200 333.300 ;
        RECT 596.100 331.200 598.200 331.500 ;
        RECT 599.100 332.100 601.200 334.200 ;
        RECT 605.100 333.150 606.900 334.950 ;
        RECT 599.100 330.000 600.000 332.100 ;
        RECT 592.800 327.600 594.900 329.700 ;
        RECT 598.500 329.100 600.000 330.000 ;
        RECT 598.500 327.600 599.700 329.100 ;
        RECT 503.400 315.600 505.200 321.600 ;
        RECT 523.800 315.600 525.600 321.600 ;
        RECT 547.800 315.600 549.600 321.600 ;
        RECT 571.800 315.600 573.600 321.600 ;
        RECT 590.400 326.700 594.900 327.600 ;
        RECT 590.400 315.600 592.200 326.700 ;
        RECT 597.900 319.050 599.700 327.600 ;
        RECT 602.400 327.600 604.500 328.500 ;
        RECT 602.400 326.400 607.200 327.600 ;
        RECT 597.900 316.950 601.050 319.050 ;
        RECT 597.900 315.600 599.700 316.950 ;
        RECT 605.400 315.600 607.200 326.400 ;
        RECT 626.850 321.600 628.050 334.950 ;
        RECT 632.100 333.150 633.900 334.950 ;
        RECT 647.700 322.800 648.600 334.950 ;
        RECT 653.100 333.150 654.900 334.950 ;
        RECT 662.550 333.450 663.450 337.950 ;
        RECT 668.100 337.050 669.900 338.850 ;
        RECT 674.100 337.050 675.900 338.850 ;
        RECT 677.700 337.050 678.600 344.400 ;
        RECT 697.200 342.000 699.000 350.400 ;
        RECT 695.700 340.800 699.000 342.000 ;
        RECT 723.000 342.000 724.800 350.400 ;
        RECT 746.700 345.600 748.500 350.400 ;
        RECT 743.400 344.400 748.500 345.600 ;
        RECT 723.000 340.800 726.300 342.000 ;
        RECT 682.950 339.450 685.050 340.050 ;
        RECT 691.950 339.450 694.050 340.050 ;
        RECT 682.950 338.550 694.050 339.450 ;
        RECT 682.950 337.950 685.050 338.550 ;
        RECT 691.950 337.950 694.050 338.550 ;
        RECT 695.700 337.050 696.600 340.800 ;
        RECT 706.950 339.450 711.000 340.050 ;
        RECT 698.100 337.050 699.900 338.850 ;
        RECT 704.100 337.050 705.900 338.850 ;
        RECT 706.950 337.950 711.450 339.450 ;
        RECT 667.950 334.950 670.050 337.050 ;
        RECT 670.950 334.950 673.050 337.050 ;
        RECT 673.950 334.950 676.050 337.050 ;
        RECT 676.950 334.950 679.050 337.050 ;
        RECT 694.950 334.950 697.050 337.050 ;
        RECT 697.950 334.950 700.050 337.050 ;
        RECT 700.950 334.950 703.050 337.050 ;
        RECT 703.950 334.950 706.050 337.050 ;
        RECT 662.550 332.550 666.450 333.450 ;
        RECT 671.100 333.150 672.900 334.950 ;
        RECT 655.950 330.450 658.050 331.050 ;
        RECT 661.950 330.450 664.050 331.050 ;
        RECT 655.950 329.550 664.050 330.450 ;
        RECT 655.950 328.950 658.050 329.550 ;
        RECT 661.950 328.950 664.050 329.550 ;
        RECT 665.550 328.050 666.450 332.550 ;
        RECT 663.000 327.900 666.450 328.050 ;
        RECT 661.950 326.550 666.450 327.900 ;
        RECT 677.700 327.600 678.600 334.950 ;
        RECT 668.400 326.700 676.200 327.600 ;
        RECT 661.950 325.950 666.000 326.550 ;
        RECT 661.950 325.800 664.050 325.950 ;
        RECT 647.700 321.900 654.300 322.800 ;
        RECT 647.700 321.600 648.600 321.900 ;
        RECT 626.400 315.600 628.200 321.600 ;
        RECT 646.800 315.600 648.600 321.600 ;
        RECT 652.800 321.600 654.300 321.900 ;
        RECT 652.800 315.600 654.600 321.600 ;
        RECT 668.400 315.600 670.200 326.700 ;
        RECT 674.400 315.600 676.200 326.700 ;
        RECT 677.400 315.600 679.200 327.600 ;
        RECT 695.700 322.800 696.600 334.950 ;
        RECT 701.100 333.150 702.900 334.950 ;
        RECT 710.550 334.050 711.450 337.950 ;
        RECT 716.100 337.050 717.900 338.850 ;
        RECT 722.100 337.050 723.900 338.850 ;
        RECT 725.400 337.050 726.300 340.800 ;
        RECT 727.950 339.450 732.000 340.050 ;
        RECT 727.950 337.950 732.450 339.450 ;
        RECT 715.950 334.950 718.050 337.050 ;
        RECT 718.950 334.950 721.050 337.050 ;
        RECT 721.950 334.950 724.050 337.050 ;
        RECT 724.950 334.950 727.050 337.050 ;
        RECT 706.950 332.550 711.450 334.050 ;
        RECT 719.100 333.150 720.900 334.950 ;
        RECT 706.950 331.950 711.000 332.550 ;
        RECT 725.400 322.800 726.300 334.950 ;
        RECT 731.550 334.050 732.450 337.950 ;
        RECT 743.400 337.050 744.300 344.400 ;
        RECT 774.000 342.000 775.800 350.400 ;
        RECT 796.500 345.600 798.300 350.400 ;
        RECT 796.500 344.400 801.600 345.600 ;
        RECT 817.800 344.400 819.600 350.400 ;
        RECT 781.950 342.450 784.050 343.050 ;
        RECT 793.950 342.450 796.050 343.200 ;
        RECT 774.000 340.800 777.300 342.000 ;
        RECT 781.950 341.550 796.050 342.450 ;
        RECT 781.950 340.950 784.050 341.550 ;
        RECT 793.950 341.100 796.050 341.550 ;
        RECT 762.000 339.450 766.050 340.050 ;
        RECT 746.100 337.050 747.900 338.850 ;
        RECT 752.100 337.050 753.900 338.850 ;
        RECT 761.550 337.950 766.050 339.450 ;
        RECT 742.950 334.950 745.050 337.050 ;
        RECT 745.950 334.950 748.050 337.050 ;
        RECT 748.950 334.950 751.050 337.050 ;
        RECT 751.950 334.950 754.050 337.050 ;
        RECT 727.950 332.550 732.450 334.050 ;
        RECT 727.950 331.950 732.000 332.550 ;
        RECT 743.400 327.600 744.300 334.950 ;
        RECT 749.100 333.150 750.900 334.950 ;
        RECT 761.550 334.050 762.450 337.950 ;
        RECT 767.100 337.050 768.900 338.850 ;
        RECT 773.100 337.050 774.900 338.850 ;
        RECT 776.400 337.050 777.300 340.800 ;
        RECT 778.950 339.450 783.000 340.050 ;
        RECT 778.950 337.950 783.450 339.450 ;
        RECT 766.950 334.950 769.050 337.050 ;
        RECT 769.950 334.950 772.050 337.050 ;
        RECT 772.950 334.950 775.050 337.050 ;
        RECT 775.950 334.950 778.050 337.050 ;
        RECT 761.550 332.550 766.050 334.050 ;
        RECT 770.100 333.150 771.900 334.950 ;
        RECT 762.000 331.950 766.050 332.550 ;
        RECT 695.700 321.900 702.300 322.800 ;
        RECT 695.700 321.600 696.600 321.900 ;
        RECT 694.800 315.600 696.600 321.600 ;
        RECT 700.800 321.600 702.300 321.900 ;
        RECT 719.700 321.900 726.300 322.800 ;
        RECT 719.700 321.600 721.200 321.900 ;
        RECT 700.800 315.600 702.600 321.600 ;
        RECT 719.400 315.600 721.200 321.600 ;
        RECT 725.400 321.600 726.300 321.900 ;
        RECT 725.400 315.600 727.200 321.600 ;
        RECT 742.800 315.600 744.600 327.600 ;
        RECT 745.800 326.700 753.600 327.600 ;
        RECT 745.800 315.600 747.600 326.700 ;
        RECT 751.800 315.600 753.600 326.700 ;
        RECT 776.400 322.800 777.300 334.950 ;
        RECT 782.550 334.050 783.450 337.950 ;
        RECT 791.100 337.050 792.900 338.850 ;
        RECT 797.100 337.050 798.900 338.850 ;
        RECT 800.700 337.050 801.600 344.400 ;
        RECT 818.400 342.300 819.600 344.400 ;
        RECT 820.800 345.300 822.600 350.400 ;
        RECT 826.800 345.300 828.600 350.400 ;
        RECT 820.800 343.950 828.600 345.300 ;
        RECT 839.400 345.300 841.200 350.400 ;
        RECT 845.400 345.300 847.200 350.400 ;
        RECT 839.400 343.950 847.200 345.300 ;
        RECT 848.400 344.400 850.200 350.400 ;
        RECT 848.400 342.300 849.600 344.400 ;
        RECT 818.400 341.250 822.150 342.300 ;
        RECT 818.100 337.050 819.900 338.850 ;
        RECT 820.950 337.050 822.150 341.250 ;
        RECT 845.850 341.250 849.600 342.300 ;
        RECT 870.000 342.000 871.800 350.400 ;
        RECT 824.100 337.050 825.900 338.850 ;
        RECT 842.100 337.050 843.900 338.850 ;
        RECT 845.850 337.050 847.050 341.250 ;
        RECT 870.000 340.800 873.300 342.000 ;
        RECT 848.100 337.050 849.900 338.850 ;
        RECT 863.100 337.050 864.900 338.850 ;
        RECT 869.100 337.050 870.900 338.850 ;
        RECT 872.400 337.050 873.300 340.800 ;
        RECT 790.950 334.950 793.050 337.050 ;
        RECT 793.950 334.950 796.050 337.050 ;
        RECT 796.950 334.950 799.050 337.050 ;
        RECT 799.950 334.950 802.050 337.050 ;
        RECT 817.950 334.950 820.050 337.050 ;
        RECT 820.950 334.950 823.050 337.050 ;
        RECT 823.950 334.950 826.050 337.050 ;
        RECT 826.950 334.950 829.050 337.050 ;
        RECT 838.950 334.950 841.050 337.050 ;
        RECT 841.950 334.950 844.050 337.050 ;
        RECT 844.950 334.950 847.050 337.050 ;
        RECT 847.950 334.950 850.050 337.050 ;
        RECT 862.950 334.950 865.050 337.050 ;
        RECT 865.950 334.950 868.050 337.050 ;
        RECT 868.950 334.950 871.050 337.050 ;
        RECT 871.950 334.950 874.050 337.050 ;
        RECT 778.950 332.550 783.450 334.050 ;
        RECT 794.100 333.150 795.900 334.950 ;
        RECT 778.950 331.950 783.000 332.550 ;
        RECT 800.700 327.600 801.600 334.950 ;
        RECT 770.700 321.900 777.300 322.800 ;
        RECT 770.700 321.600 772.200 321.900 ;
        RECT 770.400 315.600 772.200 321.600 ;
        RECT 776.400 321.600 777.300 321.900 ;
        RECT 791.400 326.700 799.200 327.600 ;
        RECT 776.400 315.600 778.200 321.600 ;
        RECT 791.400 315.600 793.200 326.700 ;
        RECT 797.400 315.600 799.200 326.700 ;
        RECT 800.400 315.600 802.200 327.600 ;
        RECT 821.850 321.600 823.050 334.950 ;
        RECT 827.100 333.150 828.900 334.950 ;
        RECT 839.100 333.150 840.900 334.950 ;
        RECT 844.950 321.600 846.150 334.950 ;
        RECT 866.100 333.150 867.900 334.950 ;
        RECT 847.950 330.450 850.050 331.050 ;
        RECT 859.950 330.450 862.050 331.050 ;
        RECT 847.950 329.550 862.050 330.450 ;
        RECT 847.950 328.950 850.050 329.550 ;
        RECT 859.950 328.950 862.050 329.550 ;
        RECT 872.400 322.800 873.300 334.950 ;
        RECT 866.700 321.900 873.300 322.800 ;
        RECT 866.700 321.600 868.200 321.900 ;
        RECT 821.400 315.600 823.200 321.600 ;
        RECT 844.800 315.600 846.600 321.600 ;
        RECT 866.400 315.600 868.200 321.600 ;
        RECT 872.400 321.600 873.300 321.900 ;
        RECT 872.400 315.600 874.200 321.600 ;
        RECT 16.800 298.500 18.600 311.400 ;
        RECT 22.800 298.500 24.600 311.400 ;
        RECT 28.800 298.500 30.600 311.400 ;
        RECT 34.800 298.500 36.600 311.400 ;
        RECT 52.800 310.500 60.600 311.400 ;
        RECT 52.800 299.400 54.600 310.500 ;
        RECT 15.900 297.300 18.600 298.500 ;
        RECT 20.700 297.300 24.600 298.500 ;
        RECT 26.700 297.300 30.600 298.500 ;
        RECT 32.700 297.300 36.600 298.500 ;
        RECT 55.800 298.500 57.600 309.600 ;
        RECT 58.800 300.600 60.600 310.500 ;
        RECT 64.800 300.600 66.600 311.400 ;
        RECT 58.800 299.700 66.600 300.600 ;
        RECT 79.800 310.500 87.600 311.400 ;
        RECT 79.800 299.400 81.600 310.500 ;
        RECT 82.800 298.500 84.600 309.600 ;
        RECT 85.800 300.600 87.600 310.500 ;
        RECT 91.800 300.600 93.600 311.400 ;
        RECT 85.800 299.700 93.600 300.600 ;
        RECT 95.550 299.400 97.350 311.400 ;
        RECT 103.050 305.400 104.850 311.400 ;
        RECT 100.950 303.300 104.850 305.400 ;
        RECT 110.850 304.500 112.650 311.400 ;
        RECT 118.650 305.400 120.450 311.400 ;
        RECT 119.250 304.500 120.450 305.400 ;
        RECT 109.950 303.450 116.550 304.500 ;
        RECT 109.950 302.700 111.750 303.450 ;
        RECT 114.750 302.700 116.550 303.450 ;
        RECT 119.250 302.400 124.050 304.500 ;
        RECT 102.150 300.600 104.850 302.400 ;
        RECT 105.750 301.800 107.550 302.400 ;
        RECT 105.750 300.900 112.050 301.800 ;
        RECT 119.250 301.500 120.450 302.400 ;
        RECT 105.750 300.600 107.550 300.900 ;
        RECT 103.950 299.700 104.850 300.600 ;
        RECT 55.800 297.600 60.900 298.500 ;
        RECT 15.900 292.050 16.800 297.300 ;
        RECT 13.950 289.950 16.800 292.050 ;
        RECT 15.900 284.700 16.800 289.950 ;
        RECT 17.700 286.800 19.500 287.400 ;
        RECT 20.700 286.800 21.900 297.300 ;
        RECT 17.700 285.600 21.900 286.800 ;
        RECT 23.700 286.800 25.500 287.400 ;
        RECT 26.700 286.800 27.900 297.300 ;
        RECT 23.700 285.600 27.900 286.800 ;
        RECT 29.700 286.800 31.500 287.400 ;
        RECT 32.700 286.800 33.900 297.300 ;
        RECT 48.000 294.450 52.050 295.050 ;
        RECT 47.550 292.950 52.050 294.450 ;
        RECT 34.950 289.950 37.050 292.050 ;
        RECT 35.100 288.150 36.900 289.950 ;
        RECT 47.550 288.900 48.450 292.950 ;
        RECT 56.100 292.050 57.900 293.850 ;
        RECT 60.000 292.050 60.900 297.600 ;
        RECT 70.950 295.950 73.050 298.050 ;
        RECT 82.800 297.600 87.900 298.500 ;
        RECT 62.100 292.050 63.900 293.850 ;
        RECT 52.950 289.950 55.050 292.050 ;
        RECT 55.950 289.950 58.050 292.050 ;
        RECT 58.950 289.950 61.050 292.050 ;
        RECT 61.950 289.950 64.050 292.050 ;
        RECT 64.950 289.950 67.050 292.050 ;
        RECT 46.950 286.800 49.050 288.900 ;
        RECT 53.100 288.150 54.900 289.950 ;
        RECT 29.700 285.600 33.900 286.800 ;
        RECT 20.700 284.700 21.900 285.600 ;
        RECT 26.700 284.700 27.900 285.600 ;
        RECT 32.700 284.700 33.900 285.600 ;
        RECT 15.900 283.500 18.600 284.700 ;
        RECT 20.700 283.500 24.600 284.700 ;
        RECT 26.700 283.500 30.600 284.700 ;
        RECT 32.700 283.500 36.600 284.700 ;
        RECT 16.800 276.600 18.600 283.500 ;
        RECT 22.800 276.600 24.600 283.500 ;
        RECT 28.800 276.600 30.600 283.500 ;
        RECT 34.800 276.600 36.600 283.500 ;
        RECT 60.000 282.600 61.050 289.950 ;
        RECT 65.100 288.150 66.900 289.950 ;
        RECT 71.550 288.450 72.450 295.950 ;
        RECT 75.000 294.450 79.050 295.050 ;
        RECT 68.550 287.550 72.450 288.450 ;
        RECT 74.550 292.950 79.050 294.450 ;
        RECT 74.550 289.050 75.450 292.950 ;
        RECT 83.100 292.050 84.900 293.850 ;
        RECT 87.000 292.050 87.900 297.600 ;
        RECT 89.100 292.050 90.900 293.850 ;
        RECT 95.550 292.050 96.750 299.400 ;
        RECT 100.950 298.800 103.050 299.700 ;
        RECT 103.950 298.800 109.050 299.700 ;
        RECT 98.850 297.600 103.050 298.800 ;
        RECT 97.950 295.800 99.750 297.600 ;
        RECT 79.950 289.950 82.050 292.050 ;
        RECT 82.950 289.950 85.050 292.050 ;
        RECT 85.950 289.950 88.050 292.050 ;
        RECT 88.950 289.950 91.050 292.050 ;
        RECT 91.950 289.950 94.050 292.050 ;
        RECT 95.550 291.750 100.050 292.050 ;
        RECT 95.550 289.950 101.850 291.750 ;
        RECT 74.550 287.550 79.050 289.050 ;
        RECT 80.100 288.150 81.900 289.950 ;
        RECT 68.550 283.050 69.450 287.550 ;
        RECT 75.000 286.950 79.050 287.550 ;
        RECT 70.950 285.450 73.050 286.050 ;
        RECT 82.950 285.450 85.050 286.050 ;
        RECT 70.950 284.550 85.050 285.450 ;
        RECT 70.950 283.950 73.050 284.550 ;
        RECT 82.950 283.950 85.050 284.550 ;
        RECT 60.000 276.600 61.800 282.600 ;
        RECT 67.950 280.950 70.050 283.050 ;
        RECT 87.000 282.600 88.050 289.950 ;
        RECT 92.100 288.150 93.900 289.950 ;
        RECT 95.550 282.600 96.750 289.950 ;
        RECT 108.150 286.200 109.050 298.800 ;
        RECT 111.150 298.800 112.050 300.900 ;
        RECT 112.950 300.300 120.450 301.500 ;
        RECT 112.950 299.700 114.750 300.300 ;
        RECT 127.050 299.400 128.850 311.400 ;
        RECT 111.150 298.500 119.550 298.800 ;
        RECT 127.950 298.500 128.850 299.400 ;
        RECT 111.150 297.900 128.850 298.500 ;
        RECT 117.750 297.300 128.850 297.900 ;
        RECT 117.750 297.000 119.550 297.300 ;
        RECT 115.950 290.400 118.050 292.050 ;
        RECT 115.950 289.200 123.900 290.400 ;
        RECT 124.950 289.950 127.050 292.050 ;
        RECT 122.100 288.600 123.900 289.200 ;
        RECT 125.100 288.150 126.900 289.950 ;
        RECT 119.100 287.400 120.900 288.000 ;
        RECT 125.100 287.400 126.000 288.150 ;
        RECT 119.100 286.200 126.000 287.400 ;
        RECT 108.150 285.000 120.150 286.200 ;
        RECT 108.150 284.400 109.950 285.000 ;
        RECT 119.100 283.200 120.150 285.000 ;
        RECT 87.000 276.600 88.800 282.600 ;
        RECT 95.550 276.600 97.350 282.600 ;
        RECT 100.950 281.700 103.050 282.600 ;
        RECT 100.950 280.500 104.700 281.700 ;
        RECT 115.350 281.550 117.150 282.300 ;
        RECT 103.650 279.600 104.700 280.500 ;
        RECT 112.200 280.500 117.150 281.550 ;
        RECT 118.650 281.400 120.450 283.200 ;
        RECT 127.950 282.600 128.850 297.300 ;
        RECT 121.950 280.500 124.050 282.600 ;
        RECT 112.200 279.600 113.250 280.500 ;
        RECT 121.950 279.600 123.000 280.500 ;
        RECT 103.650 276.600 105.450 279.600 ;
        RECT 111.450 276.600 113.250 279.600 ;
        RECT 119.250 278.700 123.000 279.600 ;
        RECT 119.250 276.600 121.050 278.700 ;
        RECT 127.050 276.600 128.850 282.600 ;
        RECT 132.150 299.400 133.950 311.400 ;
        RECT 140.550 305.400 142.350 311.400 ;
        RECT 140.550 304.500 141.750 305.400 ;
        RECT 148.350 304.500 150.150 311.400 ;
        RECT 156.150 305.400 157.950 311.400 ;
        RECT 136.950 302.400 141.750 304.500 ;
        RECT 144.450 303.450 151.050 304.500 ;
        RECT 144.450 302.700 146.250 303.450 ;
        RECT 149.250 302.700 151.050 303.450 ;
        RECT 156.150 303.300 160.050 305.400 ;
        RECT 140.550 301.500 141.750 302.400 ;
        RECT 153.450 301.800 155.250 302.400 ;
        RECT 140.550 300.300 148.050 301.500 ;
        RECT 146.250 299.700 148.050 300.300 ;
        RECT 148.950 300.900 155.250 301.800 ;
        RECT 132.150 298.500 133.050 299.400 ;
        RECT 148.950 298.800 149.850 300.900 ;
        RECT 153.450 300.600 155.250 300.900 ;
        RECT 156.150 300.600 158.850 302.400 ;
        RECT 156.150 299.700 157.050 300.600 ;
        RECT 141.450 298.500 149.850 298.800 ;
        RECT 132.150 297.900 149.850 298.500 ;
        RECT 151.950 298.800 157.050 299.700 ;
        RECT 157.950 298.800 160.050 299.700 ;
        RECT 163.650 299.400 165.450 311.400 ;
        RECT 132.150 297.300 143.250 297.900 ;
        RECT 132.150 282.600 133.050 297.300 ;
        RECT 141.450 297.000 143.250 297.300 ;
        RECT 133.950 289.950 136.050 292.050 ;
        RECT 142.950 290.400 145.050 292.050 ;
        RECT 134.100 288.150 135.900 289.950 ;
        RECT 137.100 289.200 145.050 290.400 ;
        RECT 137.100 288.600 138.900 289.200 ;
        RECT 135.000 287.400 135.900 288.150 ;
        RECT 140.100 287.400 141.900 288.000 ;
        RECT 135.000 286.200 141.900 287.400 ;
        RECT 151.950 286.200 152.850 298.800 ;
        RECT 157.950 297.600 162.150 298.800 ;
        RECT 161.250 295.800 163.050 297.600 ;
        RECT 164.250 292.050 165.450 299.400 ;
        RECT 160.950 291.750 165.450 292.050 ;
        RECT 159.150 289.950 165.450 291.750 ;
        RECT 140.850 285.000 152.850 286.200 ;
        RECT 140.850 283.200 141.900 285.000 ;
        RECT 151.050 284.400 152.850 285.000 ;
        RECT 132.150 276.600 133.950 282.600 ;
        RECT 136.950 280.500 139.050 282.600 ;
        RECT 140.550 281.400 142.350 283.200 ;
        RECT 164.250 282.600 165.450 289.950 ;
        RECT 143.850 281.550 145.650 282.300 ;
        RECT 157.950 281.700 160.050 282.600 ;
        RECT 143.850 280.500 148.800 281.550 ;
        RECT 138.000 279.600 139.050 280.500 ;
        RECT 147.750 279.600 148.800 280.500 ;
        RECT 156.300 280.500 160.050 281.700 ;
        RECT 156.300 279.600 157.350 280.500 ;
        RECT 138.000 278.700 141.750 279.600 ;
        RECT 139.950 276.600 141.750 278.700 ;
        RECT 147.750 276.600 149.550 279.600 ;
        RECT 155.550 276.600 157.350 279.600 ;
        RECT 163.650 276.600 165.450 282.600 ;
        RECT 168.150 299.400 169.950 311.400 ;
        RECT 176.550 305.400 178.350 311.400 ;
        RECT 176.550 304.500 177.750 305.400 ;
        RECT 184.350 304.500 186.150 311.400 ;
        RECT 192.150 305.400 193.950 311.400 ;
        RECT 172.950 302.400 177.750 304.500 ;
        RECT 180.450 303.450 187.050 304.500 ;
        RECT 180.450 302.700 182.250 303.450 ;
        RECT 185.250 302.700 187.050 303.450 ;
        RECT 192.150 303.300 196.050 305.400 ;
        RECT 176.550 301.500 177.750 302.400 ;
        RECT 189.450 301.800 191.250 302.400 ;
        RECT 176.550 300.300 184.050 301.500 ;
        RECT 182.250 299.700 184.050 300.300 ;
        RECT 184.950 300.900 191.250 301.800 ;
        RECT 168.150 298.500 169.050 299.400 ;
        RECT 184.950 298.800 185.850 300.900 ;
        RECT 189.450 300.600 191.250 300.900 ;
        RECT 192.150 300.600 194.850 302.400 ;
        RECT 192.150 299.700 193.050 300.600 ;
        RECT 177.450 298.500 185.850 298.800 ;
        RECT 168.150 297.900 185.850 298.500 ;
        RECT 187.950 298.800 193.050 299.700 ;
        RECT 193.950 298.800 196.050 299.700 ;
        RECT 199.650 299.400 201.450 311.400 ;
        RECT 217.800 305.400 219.600 311.400 ;
        RECT 238.800 305.400 240.600 311.400 ;
        RECT 168.150 297.300 179.250 297.900 ;
        RECT 168.150 282.600 169.050 297.300 ;
        RECT 177.450 297.000 179.250 297.300 ;
        RECT 169.950 289.950 172.050 292.050 ;
        RECT 178.950 290.400 181.050 292.050 ;
        RECT 170.100 288.150 171.900 289.950 ;
        RECT 173.100 289.200 181.050 290.400 ;
        RECT 173.100 288.600 174.900 289.200 ;
        RECT 171.000 287.400 171.900 288.150 ;
        RECT 176.100 287.400 177.900 288.000 ;
        RECT 171.000 286.200 177.900 287.400 ;
        RECT 187.950 286.200 188.850 298.800 ;
        RECT 193.950 297.600 198.150 298.800 ;
        RECT 197.250 295.800 199.050 297.600 ;
        RECT 200.250 292.050 201.450 299.400 ;
        RECT 218.400 292.050 219.600 305.400 ;
        RECT 239.400 292.050 240.600 305.400 ;
        RECT 245.550 299.400 247.350 311.400 ;
        RECT 253.050 305.400 254.850 311.400 ;
        RECT 250.950 303.300 254.850 305.400 ;
        RECT 260.850 304.500 262.650 311.400 ;
        RECT 268.650 305.400 270.450 311.400 ;
        RECT 269.250 304.500 270.450 305.400 ;
        RECT 259.950 303.450 266.550 304.500 ;
        RECT 259.950 302.700 261.750 303.450 ;
        RECT 264.750 302.700 266.550 303.450 ;
        RECT 269.250 302.400 274.050 304.500 ;
        RECT 252.150 300.600 254.850 302.400 ;
        RECT 255.750 301.800 257.550 302.400 ;
        RECT 255.750 300.900 262.050 301.800 ;
        RECT 269.250 301.500 270.450 302.400 ;
        RECT 255.750 300.600 257.550 300.900 ;
        RECT 253.950 299.700 254.850 300.600 ;
        RECT 245.550 292.050 246.750 299.400 ;
        RECT 250.950 298.800 253.050 299.700 ;
        RECT 253.950 298.800 259.050 299.700 ;
        RECT 248.850 297.600 253.050 298.800 ;
        RECT 247.950 295.800 249.750 297.600 ;
        RECT 196.950 291.750 201.450 292.050 ;
        RECT 195.150 289.950 201.450 291.750 ;
        RECT 214.950 289.950 217.050 292.050 ;
        RECT 217.950 289.950 220.050 292.050 ;
        RECT 220.950 289.950 223.050 292.050 ;
        RECT 235.950 289.950 238.050 292.050 ;
        RECT 238.950 289.950 241.050 292.050 ;
        RECT 241.950 289.950 244.050 292.050 ;
        RECT 245.550 291.750 250.050 292.050 ;
        RECT 245.550 289.950 251.850 291.750 ;
        RECT 176.850 285.000 188.850 286.200 ;
        RECT 176.850 283.200 177.900 285.000 ;
        RECT 187.050 284.400 188.850 285.000 ;
        RECT 168.150 276.600 169.950 282.600 ;
        RECT 172.950 280.500 175.050 282.600 ;
        RECT 176.550 281.400 178.350 283.200 ;
        RECT 200.250 282.600 201.450 289.950 ;
        RECT 215.100 288.150 216.900 289.950 ;
        RECT 218.400 284.700 219.600 289.950 ;
        RECT 221.100 288.150 222.900 289.950 ;
        RECT 236.100 288.150 237.900 289.950 ;
        RECT 239.400 284.700 240.600 289.950 ;
        RECT 242.100 288.150 243.900 289.950 ;
        RECT 179.850 281.550 181.650 282.300 ;
        RECT 193.950 281.700 196.050 282.600 ;
        RECT 179.850 280.500 184.800 281.550 ;
        RECT 174.000 279.600 175.050 280.500 ;
        RECT 183.750 279.600 184.800 280.500 ;
        RECT 192.300 280.500 196.050 281.700 ;
        RECT 192.300 279.600 193.350 280.500 ;
        RECT 174.000 278.700 177.750 279.600 ;
        RECT 175.950 276.600 177.750 278.700 ;
        RECT 183.750 276.600 185.550 279.600 ;
        RECT 191.550 276.600 193.350 279.600 ;
        RECT 199.650 276.600 201.450 282.600 ;
        RECT 215.400 283.800 219.600 284.700 ;
        RECT 236.400 283.800 240.600 284.700 ;
        RECT 215.400 276.600 217.200 283.800 ;
        RECT 236.400 276.600 238.200 283.800 ;
        RECT 245.550 282.600 246.750 289.950 ;
        RECT 258.150 286.200 259.050 298.800 ;
        RECT 261.150 298.800 262.050 300.900 ;
        RECT 262.950 300.300 270.450 301.500 ;
        RECT 262.950 299.700 264.750 300.300 ;
        RECT 277.050 299.400 278.850 311.400 ;
        RECT 295.800 305.400 297.600 311.400 ;
        RECT 319.800 305.400 321.600 311.400 ;
        RECT 261.150 298.500 269.550 298.800 ;
        RECT 277.950 298.500 278.850 299.400 ;
        RECT 261.150 297.900 278.850 298.500 ;
        RECT 267.750 297.300 278.850 297.900 ;
        RECT 267.750 297.000 269.550 297.300 ;
        RECT 265.950 290.400 268.050 292.050 ;
        RECT 265.950 289.200 273.900 290.400 ;
        RECT 274.950 289.950 277.050 292.050 ;
        RECT 272.100 288.600 273.900 289.200 ;
        RECT 275.100 288.150 276.900 289.950 ;
        RECT 269.100 287.400 270.900 288.000 ;
        RECT 275.100 287.400 276.000 288.150 ;
        RECT 269.100 286.200 276.000 287.400 ;
        RECT 258.150 285.000 270.150 286.200 ;
        RECT 258.150 284.400 259.950 285.000 ;
        RECT 269.100 283.200 270.150 285.000 ;
        RECT 245.550 276.600 247.350 282.600 ;
        RECT 250.950 281.700 253.050 282.600 ;
        RECT 250.950 280.500 254.700 281.700 ;
        RECT 265.350 281.550 267.150 282.300 ;
        RECT 253.650 279.600 254.700 280.500 ;
        RECT 262.200 280.500 267.150 281.550 ;
        RECT 268.650 281.400 270.450 283.200 ;
        RECT 277.950 282.600 278.850 297.300 ;
        RECT 290.100 292.050 291.900 293.850 ;
        RECT 295.950 292.050 297.150 305.400 ;
        RECT 301.950 294.450 304.050 295.050 ;
        RECT 310.950 294.450 313.050 295.050 ;
        RECT 301.950 293.550 313.050 294.450 ;
        RECT 301.950 292.950 304.050 293.550 ;
        RECT 310.950 292.950 313.050 293.550 ;
        RECT 320.400 292.050 321.600 305.400 ;
        RECT 338.700 300.600 340.500 311.400 ;
        RECT 338.700 299.400 342.300 300.600 ;
        RECT 338.100 292.050 339.900 293.850 ;
        RECT 341.400 292.050 342.300 299.400 ;
        RECT 347.550 299.400 349.350 311.400 ;
        RECT 355.050 305.400 356.850 311.400 ;
        RECT 352.950 303.300 356.850 305.400 ;
        RECT 362.850 304.500 364.650 311.400 ;
        RECT 370.650 305.400 372.450 311.400 ;
        RECT 371.250 304.500 372.450 305.400 ;
        RECT 361.950 303.450 368.550 304.500 ;
        RECT 361.950 302.700 363.750 303.450 ;
        RECT 366.750 302.700 368.550 303.450 ;
        RECT 371.250 302.400 376.050 304.500 ;
        RECT 354.150 300.600 356.850 302.400 ;
        RECT 357.750 301.800 359.550 302.400 ;
        RECT 357.750 300.900 364.050 301.800 ;
        RECT 371.250 301.500 372.450 302.400 ;
        RECT 357.750 300.600 359.550 300.900 ;
        RECT 355.950 299.700 356.850 300.600 ;
        RECT 344.100 292.050 345.900 293.850 ;
        RECT 347.550 292.050 348.750 299.400 ;
        RECT 352.950 298.800 355.050 299.700 ;
        RECT 355.950 298.800 361.050 299.700 ;
        RECT 350.850 297.600 355.050 298.800 ;
        RECT 349.950 295.800 351.750 297.600 ;
        RECT 289.950 289.950 292.050 292.050 ;
        RECT 292.950 289.950 295.050 292.050 ;
        RECT 295.950 289.950 298.050 292.050 ;
        RECT 298.950 289.950 301.050 292.050 ;
        RECT 316.950 289.950 319.050 292.050 ;
        RECT 319.950 289.950 322.050 292.050 ;
        RECT 322.950 289.950 325.050 292.050 ;
        RECT 337.950 289.950 340.050 292.050 ;
        RECT 340.950 289.950 343.050 292.050 ;
        RECT 343.950 289.950 346.050 292.050 ;
        RECT 347.550 291.750 352.050 292.050 ;
        RECT 347.550 289.950 353.850 291.750 ;
        RECT 293.100 288.150 294.900 289.950 ;
        RECT 296.850 285.750 298.050 289.950 ;
        RECT 299.100 288.150 300.900 289.950 ;
        RECT 317.100 288.150 318.900 289.950 ;
        RECT 296.850 284.700 300.600 285.750 ;
        RECT 320.400 284.700 321.600 289.950 ;
        RECT 323.100 288.150 324.900 289.950 ;
        RECT 271.950 280.500 274.050 282.600 ;
        RECT 262.200 279.600 263.250 280.500 ;
        RECT 271.950 279.600 273.000 280.500 ;
        RECT 253.650 276.600 255.450 279.600 ;
        RECT 261.450 276.600 263.250 279.600 ;
        RECT 269.250 278.700 273.000 279.600 ;
        RECT 269.250 276.600 271.050 278.700 ;
        RECT 277.050 276.600 278.850 282.600 ;
        RECT 290.400 281.700 298.200 283.050 ;
        RECT 290.400 276.600 292.200 281.700 ;
        RECT 296.400 276.600 298.200 281.700 ;
        RECT 299.400 282.600 300.600 284.700 ;
        RECT 317.400 283.800 321.600 284.700 ;
        RECT 299.400 276.600 301.200 282.600 ;
        RECT 317.400 276.600 319.200 283.800 ;
        RECT 341.400 279.600 342.300 289.950 ;
        RECT 347.550 282.600 348.750 289.950 ;
        RECT 360.150 286.200 361.050 298.800 ;
        RECT 363.150 298.800 364.050 300.900 ;
        RECT 364.950 300.300 372.450 301.500 ;
        RECT 364.950 299.700 366.750 300.300 ;
        RECT 379.050 299.400 380.850 311.400 ;
        RECT 394.800 299.400 396.600 311.400 ;
        RECT 397.800 300.300 399.600 311.400 ;
        RECT 403.800 300.300 405.600 311.400 ;
        RECT 397.800 299.400 405.600 300.300 ;
        RECT 416.400 305.400 418.200 311.400 ;
        RECT 363.150 298.500 371.550 298.800 ;
        RECT 379.950 298.500 380.850 299.400 ;
        RECT 363.150 297.900 380.850 298.500 ;
        RECT 369.750 297.300 380.850 297.900 ;
        RECT 369.750 297.000 371.550 297.300 ;
        RECT 367.950 290.400 370.050 292.050 ;
        RECT 367.950 289.200 375.900 290.400 ;
        RECT 376.950 289.950 379.050 292.050 ;
        RECT 374.100 288.600 375.900 289.200 ;
        RECT 377.100 288.150 378.900 289.950 ;
        RECT 371.100 287.400 372.900 288.000 ;
        RECT 377.100 287.400 378.000 288.150 ;
        RECT 371.100 286.200 378.000 287.400 ;
        RECT 360.150 285.000 372.150 286.200 ;
        RECT 360.150 284.400 361.950 285.000 ;
        RECT 371.100 283.200 372.150 285.000 ;
        RECT 340.800 276.600 342.600 279.600 ;
        RECT 347.550 276.600 349.350 282.600 ;
        RECT 352.950 281.700 355.050 282.600 ;
        RECT 352.950 280.500 356.700 281.700 ;
        RECT 367.350 281.550 369.150 282.300 ;
        RECT 355.650 279.600 356.700 280.500 ;
        RECT 364.200 280.500 369.150 281.550 ;
        RECT 370.650 281.400 372.450 283.200 ;
        RECT 379.950 282.600 380.850 297.300 ;
        RECT 395.400 292.050 396.300 299.400 ;
        RECT 416.400 298.500 417.600 305.400 ;
        RECT 422.400 299.400 424.200 311.400 ;
        RECT 416.400 297.600 422.100 298.500 ;
        RECT 420.150 296.700 422.100 297.600 ;
        RECT 401.100 292.050 402.900 293.850 ;
        RECT 416.100 292.050 417.900 293.850 ;
        RECT 394.950 289.950 397.050 292.050 ;
        RECT 397.950 289.950 400.050 292.050 ;
        RECT 400.950 289.950 403.050 292.050 ;
        RECT 403.950 289.950 406.050 292.050 ;
        RECT 415.950 289.950 418.050 292.050 ;
        RECT 373.950 280.500 376.050 282.600 ;
        RECT 364.200 279.600 365.250 280.500 ;
        RECT 373.950 279.600 375.000 280.500 ;
        RECT 355.650 276.600 357.450 279.600 ;
        RECT 363.450 276.600 365.250 279.600 ;
        RECT 371.250 278.700 375.000 279.600 ;
        RECT 371.250 276.600 373.050 278.700 ;
        RECT 379.050 276.600 380.850 282.600 ;
        RECT 395.400 282.600 396.300 289.950 ;
        RECT 398.100 288.150 399.900 289.950 ;
        RECT 404.100 288.150 405.900 289.950 ;
        RECT 420.150 285.300 421.050 296.700 ;
        RECT 423.000 292.050 424.200 299.400 ;
        RECT 440.400 305.400 442.200 311.400 ;
        RECT 427.950 297.450 430.050 298.050 ;
        RECT 436.950 297.450 439.050 298.050 ;
        RECT 427.950 296.550 439.050 297.450 ;
        RECT 427.950 295.950 430.050 296.550 ;
        RECT 436.950 295.950 439.050 296.550 ;
        RECT 440.400 292.050 441.600 305.400 ;
        RECT 461.700 300.600 463.500 311.400 ;
        RECT 461.700 299.400 465.300 300.600 ;
        RECT 479.400 300.300 481.200 311.400 ;
        RECT 485.400 300.300 487.200 311.400 ;
        RECT 479.400 299.400 487.200 300.300 ;
        RECT 488.400 299.400 490.200 311.400 ;
        RECT 495.150 299.400 496.950 311.400 ;
        RECT 503.550 305.400 505.350 311.400 ;
        RECT 503.550 304.500 504.750 305.400 ;
        RECT 511.350 304.500 513.150 311.400 ;
        RECT 519.150 305.400 520.950 311.400 ;
        RECT 499.950 302.400 504.750 304.500 ;
        RECT 507.450 303.450 514.050 304.500 ;
        RECT 507.450 302.700 509.250 303.450 ;
        RECT 512.250 302.700 514.050 303.450 ;
        RECT 519.150 303.300 523.050 305.400 ;
        RECT 503.550 301.500 504.750 302.400 ;
        RECT 516.450 301.800 518.250 302.400 ;
        RECT 503.550 300.300 511.050 301.500 ;
        RECT 509.250 299.700 511.050 300.300 ;
        RECT 511.950 300.900 518.250 301.800 ;
        RECT 461.100 292.050 462.900 293.850 ;
        RECT 464.400 292.050 465.300 299.400 ;
        RECT 466.950 297.450 469.050 298.050 ;
        RECT 484.950 297.450 487.050 298.050 ;
        RECT 466.950 296.550 487.050 297.450 ;
        RECT 466.950 295.950 469.050 296.550 ;
        RECT 484.950 295.950 487.050 296.550 ;
        RECT 467.100 292.050 468.900 293.850 ;
        RECT 482.100 292.050 483.900 293.850 ;
        RECT 488.700 292.050 489.600 299.400 ;
        RECT 495.150 298.500 496.050 299.400 ;
        RECT 511.950 298.800 512.850 300.900 ;
        RECT 516.450 300.600 518.250 300.900 ;
        RECT 519.150 300.600 521.850 302.400 ;
        RECT 519.150 299.700 520.050 300.600 ;
        RECT 504.450 298.500 512.850 298.800 ;
        RECT 495.150 297.900 512.850 298.500 ;
        RECT 514.950 298.800 520.050 299.700 ;
        RECT 520.950 298.800 523.050 299.700 ;
        RECT 526.650 299.400 528.450 311.400 ;
        RECT 541.800 299.400 543.600 311.400 ;
        RECT 547.800 305.400 549.600 311.400 ;
        RECT 565.800 305.400 567.600 311.400 ;
        RECT 495.150 297.300 506.250 297.900 ;
        RECT 421.950 289.950 424.200 292.050 ;
        RECT 436.950 289.950 439.050 292.050 ;
        RECT 439.950 289.950 442.050 292.050 ;
        RECT 442.950 289.950 445.050 292.050 ;
        RECT 460.950 289.950 463.050 292.050 ;
        RECT 463.950 289.950 466.050 292.050 ;
        RECT 466.950 289.950 469.050 292.050 ;
        RECT 478.950 289.950 481.050 292.050 ;
        RECT 481.950 289.950 484.050 292.050 ;
        RECT 484.950 289.950 487.050 292.050 ;
        RECT 487.950 289.950 490.050 292.050 ;
        RECT 420.150 284.400 422.100 285.300 ;
        RECT 416.400 283.500 422.100 284.400 ;
        RECT 395.400 281.400 400.500 282.600 ;
        RECT 398.700 276.600 400.500 281.400 ;
        RECT 416.400 279.600 417.600 283.500 ;
        RECT 423.000 282.600 424.200 289.950 ;
        RECT 437.100 288.150 438.900 289.950 ;
        RECT 440.400 284.700 441.600 289.950 ;
        RECT 443.100 288.150 444.900 289.950 ;
        RECT 445.950 285.450 448.050 286.050 ;
        RECT 460.950 285.450 463.050 286.050 ;
        RECT 440.400 283.800 444.600 284.700 ;
        RECT 445.950 284.550 463.050 285.450 ;
        RECT 445.950 283.950 448.050 284.550 ;
        RECT 460.950 283.950 463.050 284.550 ;
        RECT 416.400 276.600 418.200 279.600 ;
        RECT 422.400 276.600 424.200 282.600 ;
        RECT 442.800 276.600 444.600 283.800 ;
        RECT 464.400 279.600 465.300 289.950 ;
        RECT 479.100 288.150 480.900 289.950 ;
        RECT 485.100 288.150 486.900 289.950 ;
        RECT 488.700 282.600 489.600 289.950 ;
        RECT 484.500 281.400 489.600 282.600 ;
        RECT 495.150 282.600 496.050 297.300 ;
        RECT 504.450 297.000 506.250 297.300 ;
        RECT 496.950 289.950 499.050 292.050 ;
        RECT 505.950 290.400 508.050 292.050 ;
        RECT 497.100 288.150 498.900 289.950 ;
        RECT 500.100 289.200 508.050 290.400 ;
        RECT 500.100 288.600 501.900 289.200 ;
        RECT 498.000 287.400 498.900 288.150 ;
        RECT 503.100 287.400 504.900 288.000 ;
        RECT 498.000 286.200 504.900 287.400 ;
        RECT 514.950 286.200 515.850 298.800 ;
        RECT 520.950 297.600 525.150 298.800 ;
        RECT 524.250 295.800 526.050 297.600 ;
        RECT 527.250 292.050 528.450 299.400 ;
        RECT 542.400 292.050 543.300 299.400 ;
        RECT 545.100 292.050 546.900 293.850 ;
        RECT 523.950 291.750 528.450 292.050 ;
        RECT 522.150 289.950 528.450 291.750 ;
        RECT 541.950 289.950 544.050 292.050 ;
        RECT 544.950 289.950 547.050 292.050 ;
        RECT 503.850 285.000 515.850 286.200 ;
        RECT 503.850 283.200 504.900 285.000 ;
        RECT 514.050 284.400 515.850 285.000 ;
        RECT 463.800 276.600 465.600 279.600 ;
        RECT 484.500 276.600 486.300 281.400 ;
        RECT 495.150 276.600 496.950 282.600 ;
        RECT 499.950 280.500 502.050 282.600 ;
        RECT 503.550 281.400 505.350 283.200 ;
        RECT 527.250 282.600 528.450 289.950 ;
        RECT 506.850 281.550 508.650 282.300 ;
        RECT 520.950 281.700 523.050 282.600 ;
        RECT 506.850 280.500 511.800 281.550 ;
        RECT 501.000 279.600 502.050 280.500 ;
        RECT 510.750 279.600 511.800 280.500 ;
        RECT 519.300 280.500 523.050 281.700 ;
        RECT 519.300 279.600 520.350 280.500 ;
        RECT 501.000 278.700 504.750 279.600 ;
        RECT 502.950 276.600 504.750 278.700 ;
        RECT 510.750 276.600 512.550 279.600 ;
        RECT 518.550 276.600 520.350 279.600 ;
        RECT 526.650 276.600 528.450 282.600 ;
        RECT 542.400 282.600 543.300 289.950 ;
        RECT 548.700 285.300 549.600 305.400 ;
        RECT 566.400 292.050 567.600 305.400 ;
        RECT 581.400 299.400 583.200 311.400 ;
        RECT 588.900 300.900 590.700 311.400 ;
        RECT 608.400 305.400 610.200 311.400 ;
        RECT 588.900 299.400 591.300 300.900 ;
        RECT 581.400 297.900 582.600 299.400 ;
        RECT 581.400 296.700 588.600 297.900 ;
        RECT 586.800 296.100 588.600 296.700 ;
        RECT 569.100 292.050 570.900 293.850 ;
        RECT 584.100 292.050 585.900 293.850 ;
        RECT 550.950 289.950 553.050 292.050 ;
        RECT 565.950 289.950 568.050 292.050 ;
        RECT 568.950 289.950 571.050 292.050 ;
        RECT 580.950 289.950 583.050 292.050 ;
        RECT 583.950 289.950 586.050 292.050 ;
        RECT 551.100 288.150 552.900 289.950 ;
        RECT 545.100 284.400 552.600 285.300 ;
        RECT 545.100 283.500 546.900 284.400 ;
        RECT 542.400 280.800 545.100 282.600 ;
        RECT 543.300 276.600 545.100 280.800 ;
        RECT 550.800 276.600 552.600 284.400 ;
        RECT 566.400 279.600 567.600 289.950 ;
        RECT 581.100 288.150 582.900 289.950 ;
        RECT 587.700 285.600 588.600 296.100 ;
        RECT 589.950 292.050 591.300 299.400 ;
        RECT 605.100 292.050 606.900 293.850 ;
        RECT 608.400 292.050 609.600 305.400 ;
        RECT 626.400 300.300 628.200 311.400 ;
        RECT 632.400 300.300 634.200 311.400 ;
        RECT 626.400 299.400 634.200 300.300 ;
        RECT 635.400 299.400 637.200 311.400 ;
        RECT 652.800 305.400 654.600 311.400 ;
        RECT 629.100 292.050 630.900 293.850 ;
        RECT 635.700 292.050 636.600 299.400 ;
        RECT 637.950 294.450 640.050 295.050 ;
        RECT 646.950 294.450 649.050 295.050 ;
        RECT 637.950 293.550 649.050 294.450 ;
        RECT 637.950 292.950 640.050 293.550 ;
        RECT 646.950 292.950 649.050 293.550 ;
        RECT 653.400 292.050 654.600 305.400 ;
        RECT 671.400 305.400 673.200 311.400 ;
        RECT 689.400 305.400 691.200 311.400 ;
        RECT 656.100 292.050 657.900 293.850 ;
        RECT 668.100 292.050 669.900 293.850 ;
        RECT 671.400 292.050 672.600 305.400 ;
        RECT 689.700 305.100 691.200 305.400 ;
        RECT 695.400 305.400 697.200 311.400 ;
        RECT 718.800 305.400 720.600 311.400 ;
        RECT 742.800 305.400 744.600 311.400 ;
        RECT 764.400 305.400 766.200 311.400 ;
        RECT 695.400 305.100 696.300 305.400 ;
        RECT 689.700 304.200 696.300 305.100 ;
        RECT 689.100 292.050 690.900 293.850 ;
        RECT 695.400 292.050 696.300 304.200 ;
        RECT 713.100 292.050 714.900 293.850 ;
        RECT 718.950 292.050 720.150 305.400 ;
        RECT 727.950 297.450 730.050 298.050 ;
        RECT 733.950 297.450 736.050 298.050 ;
        RECT 727.950 296.550 736.050 297.450 ;
        RECT 727.950 295.950 730.050 296.550 ;
        RECT 733.950 295.950 736.050 296.550 ;
        RECT 724.950 294.450 727.050 295.050 ;
        RECT 730.950 294.450 733.050 295.050 ;
        RECT 724.950 293.550 733.050 294.450 ;
        RECT 724.950 292.950 727.050 293.550 ;
        RECT 730.950 292.950 733.050 293.550 ;
        RECT 737.100 292.050 738.900 293.850 ;
        RECT 742.950 292.050 744.150 305.400 ;
        RECT 764.700 305.100 766.200 305.400 ;
        RECT 770.400 305.400 772.200 311.400 ;
        RECT 788.400 305.400 790.200 311.400 ;
        RECT 770.400 305.100 771.300 305.400 ;
        RECT 764.700 304.200 771.300 305.100 ;
        RECT 788.700 305.100 790.200 305.400 ;
        RECT 794.400 305.400 796.200 311.400 ;
        RECT 815.400 305.400 817.200 311.400 ;
        RECT 794.400 305.100 795.300 305.400 ;
        RECT 788.700 304.200 795.300 305.100 ;
        RECT 757.950 297.450 760.050 298.050 ;
        RECT 766.950 297.450 769.050 298.050 ;
        RECT 757.950 296.550 769.050 297.450 ;
        RECT 757.950 295.950 760.050 296.550 ;
        RECT 766.950 295.950 769.050 296.550 ;
        RECT 764.100 292.050 765.900 293.850 ;
        RECT 770.400 292.050 771.300 304.200 ;
        RECT 788.100 292.050 789.900 293.850 ;
        RECT 794.400 292.050 795.300 304.200 ;
        RECT 812.100 292.050 813.900 293.850 ;
        RECT 815.400 292.050 816.600 305.400 ;
        RECT 830.400 300.300 832.200 311.400 ;
        RECT 836.400 300.300 838.200 311.400 ;
        RECT 830.400 299.400 838.200 300.300 ;
        RECT 839.400 299.400 841.200 311.400 ;
        RECT 856.800 305.400 858.600 311.400 ;
        RECT 857.700 305.100 858.600 305.400 ;
        RECT 862.800 305.400 864.600 311.400 ;
        RECT 862.800 305.100 864.300 305.400 ;
        RECT 857.700 304.200 864.300 305.100 ;
        RECT 826.950 297.450 829.050 298.050 ;
        RECT 835.950 297.450 838.050 298.050 ;
        RECT 826.950 296.550 838.050 297.450 ;
        RECT 826.950 295.950 829.050 296.550 ;
        RECT 835.950 295.950 838.050 296.550 ;
        RECT 817.950 294.450 820.050 295.050 ;
        RECT 817.950 293.550 825.450 294.450 ;
        RECT 817.950 292.950 820.050 293.550 ;
        RECT 589.950 289.950 592.050 292.050 ;
        RECT 604.950 289.950 607.050 292.050 ;
        RECT 607.950 289.950 610.050 292.050 ;
        RECT 625.950 289.950 628.050 292.050 ;
        RECT 628.950 289.950 631.050 292.050 ;
        RECT 631.950 289.950 634.050 292.050 ;
        RECT 634.950 289.950 637.050 292.050 ;
        RECT 652.950 289.950 655.050 292.050 ;
        RECT 655.950 289.950 658.050 292.050 ;
        RECT 667.950 289.950 670.050 292.050 ;
        RECT 670.950 289.950 673.050 292.050 ;
        RECT 685.950 289.950 688.050 292.050 ;
        RECT 688.950 289.950 691.050 292.050 ;
        RECT 691.950 289.950 694.050 292.050 ;
        RECT 694.950 289.950 697.050 292.050 ;
        RECT 712.950 289.950 715.050 292.050 ;
        RECT 715.950 289.950 718.050 292.050 ;
        RECT 718.950 289.950 721.050 292.050 ;
        RECT 721.950 289.950 724.050 292.050 ;
        RECT 736.950 289.950 739.050 292.050 ;
        RECT 739.950 289.950 742.050 292.050 ;
        RECT 742.950 289.950 745.050 292.050 ;
        RECT 745.950 289.950 748.050 292.050 ;
        RECT 760.950 289.950 763.050 292.050 ;
        RECT 763.950 289.950 766.050 292.050 ;
        RECT 766.950 289.950 769.050 292.050 ;
        RECT 769.950 289.950 772.050 292.050 ;
        RECT 784.950 289.950 787.050 292.050 ;
        RECT 787.950 289.950 790.050 292.050 ;
        RECT 790.950 289.950 793.050 292.050 ;
        RECT 793.950 289.950 796.050 292.050 ;
        RECT 811.950 289.950 814.050 292.050 ;
        RECT 814.950 289.950 817.050 292.050 ;
        RECT 586.800 284.700 588.600 285.600 ;
        RECT 585.300 283.800 588.600 284.700 ;
        RECT 585.300 279.600 586.200 283.800 ;
        RECT 591.000 282.600 592.050 289.950 ;
        RECT 565.800 276.600 567.600 279.600 ;
        RECT 584.400 276.600 586.200 279.600 ;
        RECT 590.400 276.600 592.200 282.600 ;
        RECT 608.400 279.600 609.600 289.950 ;
        RECT 626.100 288.150 627.900 289.950 ;
        RECT 632.100 288.150 633.900 289.950 ;
        RECT 613.950 285.450 616.050 286.050 ;
        RECT 628.950 285.450 631.050 286.050 ;
        RECT 613.950 284.550 631.050 285.450 ;
        RECT 613.950 283.950 616.050 284.550 ;
        RECT 628.950 283.950 631.050 284.550 ;
        RECT 635.700 282.600 636.600 289.950 ;
        RECT 631.500 281.400 636.600 282.600 ;
        RECT 608.400 276.600 610.200 279.600 ;
        RECT 631.500 276.600 633.300 281.400 ;
        RECT 653.400 279.600 654.600 289.950 ;
        RECT 652.800 276.600 654.600 279.600 ;
        RECT 671.400 279.600 672.600 289.950 ;
        RECT 686.100 288.150 687.900 289.950 ;
        RECT 692.100 288.150 693.900 289.950 ;
        RECT 695.400 286.200 696.300 289.950 ;
        RECT 700.950 288.450 703.050 289.050 ;
        RECT 709.950 288.450 712.050 289.050 ;
        RECT 700.950 287.550 712.050 288.450 ;
        RECT 716.100 288.150 717.900 289.950 ;
        RECT 700.950 286.950 703.050 287.550 ;
        RECT 709.950 286.950 712.050 287.550 ;
        RECT 693.000 285.000 696.300 286.200 ;
        RECT 719.850 285.750 721.050 289.950 ;
        RECT 722.100 288.150 723.900 289.950 ;
        RECT 740.100 288.150 741.900 289.950 ;
        RECT 743.850 285.750 745.050 289.950 ;
        RECT 746.100 288.150 747.900 289.950 ;
        RECT 761.100 288.150 762.900 289.950 ;
        RECT 767.100 288.150 768.900 289.950 ;
        RECT 770.400 286.200 771.300 289.950 ;
        RECT 785.100 288.150 786.900 289.950 ;
        RECT 791.100 288.150 792.900 289.950 ;
        RECT 794.400 286.200 795.300 289.950 ;
        RECT 671.400 276.600 673.200 279.600 ;
        RECT 693.000 276.600 694.800 285.000 ;
        RECT 719.850 284.700 723.600 285.750 ;
        RECT 743.850 284.700 747.600 285.750 ;
        RECT 713.400 281.700 721.200 283.050 ;
        RECT 713.400 276.600 715.200 281.700 ;
        RECT 719.400 276.600 721.200 281.700 ;
        RECT 722.400 282.600 723.600 284.700 ;
        RECT 722.400 276.600 724.200 282.600 ;
        RECT 737.400 281.700 745.200 283.050 ;
        RECT 737.400 276.600 739.200 281.700 ;
        RECT 743.400 276.600 745.200 281.700 ;
        RECT 746.400 282.600 747.600 284.700 ;
        RECT 768.000 285.000 771.300 286.200 ;
        RECT 792.000 285.000 795.300 286.200 ;
        RECT 746.400 276.600 748.200 282.600 ;
        RECT 768.000 276.600 769.800 285.000 ;
        RECT 792.000 276.600 793.800 285.000 ;
        RECT 815.400 279.600 816.600 289.950 ;
        RECT 824.550 289.050 825.450 293.550 ;
        RECT 833.100 292.050 834.900 293.850 ;
        RECT 839.700 292.050 840.600 299.400 ;
        RECT 844.950 294.450 847.050 295.050 ;
        RECT 853.950 294.450 856.050 295.050 ;
        RECT 844.950 293.550 856.050 294.450 ;
        RECT 844.950 292.950 847.050 293.550 ;
        RECT 853.950 292.950 856.050 293.550 ;
        RECT 857.700 292.050 858.600 304.200 ;
        RECT 878.400 300.300 880.200 311.400 ;
        RECT 884.400 300.300 886.200 311.400 ;
        RECT 878.400 299.400 886.200 300.300 ;
        RECT 887.400 299.400 889.200 311.400 ;
        RECT 862.950 297.450 865.050 298.050 ;
        RECT 877.950 297.450 880.050 298.050 ;
        RECT 862.950 296.550 880.050 297.450 ;
        RECT 862.950 295.950 865.050 296.550 ;
        RECT 877.950 295.950 880.050 296.550 ;
        RECT 868.950 294.450 873.000 295.050 ;
        RECT 863.100 292.050 864.900 293.850 ;
        RECT 868.950 292.950 873.450 294.450 ;
        RECT 829.950 289.950 832.050 292.050 ;
        RECT 832.950 289.950 835.050 292.050 ;
        RECT 835.950 289.950 838.050 292.050 ;
        RECT 838.950 289.950 841.050 292.050 ;
        RECT 856.950 289.950 859.050 292.050 ;
        RECT 859.950 289.950 862.050 292.050 ;
        RECT 862.950 289.950 865.050 292.050 ;
        RECT 865.950 289.950 868.050 292.050 ;
        RECT 824.550 287.550 829.050 289.050 ;
        RECT 830.100 288.150 831.900 289.950 ;
        RECT 836.100 288.150 837.900 289.950 ;
        RECT 825.000 286.950 829.050 287.550 ;
        RECT 839.700 282.600 840.600 289.950 ;
        RECT 857.700 286.200 858.600 289.950 ;
        RECT 860.100 288.150 861.900 289.950 ;
        RECT 866.100 288.150 867.900 289.950 ;
        RECT 872.550 288.450 873.450 292.950 ;
        RECT 881.100 292.050 882.900 293.850 ;
        RECT 887.700 292.050 888.600 299.400 ;
        RECT 877.950 289.950 880.050 292.050 ;
        RECT 880.950 289.950 883.050 292.050 ;
        RECT 883.950 289.950 886.050 292.050 ;
        RECT 886.950 289.950 889.050 292.050 ;
        RECT 869.550 287.550 873.450 288.450 ;
        RECT 878.100 288.150 879.900 289.950 ;
        RECT 884.100 288.150 885.900 289.950 ;
        RECT 857.700 285.000 861.000 286.200 ;
        RECT 835.500 281.400 840.600 282.600 ;
        RECT 815.400 276.600 817.200 279.600 ;
        RECT 835.500 276.600 837.300 281.400 ;
        RECT 859.200 276.600 861.000 285.000 ;
        RECT 869.550 283.050 870.450 287.550 ;
        RECT 871.950 285.450 874.050 286.050 ;
        RECT 880.950 285.450 883.050 286.050 ;
        RECT 871.950 284.550 883.050 285.450 ;
        RECT 871.950 283.950 874.050 284.550 ;
        RECT 880.950 283.950 883.050 284.550 ;
        RECT 868.950 280.950 871.050 283.050 ;
        RECT 887.700 282.600 888.600 289.950 ;
        RECT 883.500 281.400 888.600 282.600 ;
        RECT 883.500 276.600 885.300 281.400 ;
        RECT 16.800 265.500 18.600 272.400 ;
        RECT 22.800 265.500 24.600 272.400 ;
        RECT 28.800 265.500 30.600 272.400 ;
        RECT 34.800 265.500 36.600 272.400 ;
        RECT 52.800 266.400 54.600 272.400 ;
        RECT 15.900 264.300 18.600 265.500 ;
        RECT 20.700 264.300 24.600 265.500 ;
        RECT 26.700 264.300 30.600 265.500 ;
        RECT 32.700 264.300 36.600 265.500 ;
        RECT 53.400 264.300 54.600 266.400 ;
        RECT 55.800 267.300 57.600 272.400 ;
        RECT 61.800 267.300 63.600 272.400 ;
        RECT 55.800 265.950 63.600 267.300 ;
        RECT 79.800 266.400 81.600 272.400 ;
        RECT 85.800 269.400 87.600 272.400 ;
        RECT 15.900 259.050 16.800 264.300 ;
        RECT 20.700 263.400 21.900 264.300 ;
        RECT 26.700 263.400 27.900 264.300 ;
        RECT 32.700 263.400 33.900 264.300 ;
        RECT 17.700 262.200 21.900 263.400 ;
        RECT 17.700 261.600 19.500 262.200 ;
        RECT 13.950 256.950 16.800 259.050 ;
        RECT 15.900 251.700 16.800 256.950 ;
        RECT 20.700 251.700 21.900 262.200 ;
        RECT 23.700 262.200 27.900 263.400 ;
        RECT 23.700 261.600 25.500 262.200 ;
        RECT 26.700 251.700 27.900 262.200 ;
        RECT 29.700 262.200 33.900 263.400 ;
        RECT 53.400 263.250 57.150 264.300 ;
        RECT 29.700 261.600 31.500 262.200 ;
        RECT 32.700 251.700 33.900 262.200 ;
        RECT 35.100 259.050 36.900 260.850 ;
        RECT 53.100 259.050 54.900 260.850 ;
        RECT 55.950 259.050 57.150 263.250 ;
        RECT 59.100 259.050 60.900 260.850 ;
        RECT 79.800 259.050 81.000 266.400 ;
        RECT 86.400 265.500 87.600 269.400 ;
        RECT 100.800 266.400 102.600 272.400 ;
        RECT 81.900 264.600 87.600 265.500 ;
        RECT 81.900 263.700 83.850 264.600 ;
        RECT 34.950 256.950 37.050 259.050 ;
        RECT 52.950 256.950 55.050 259.050 ;
        RECT 55.950 256.950 58.050 259.050 ;
        RECT 58.950 256.950 61.050 259.050 ;
        RECT 61.950 256.950 64.050 259.050 ;
        RECT 79.800 256.950 82.050 259.050 ;
        RECT 15.900 250.500 18.600 251.700 ;
        RECT 20.700 250.500 24.600 251.700 ;
        RECT 26.700 250.500 30.600 251.700 ;
        RECT 32.700 250.500 36.600 251.700 ;
        RECT 16.800 237.600 18.600 250.500 ;
        RECT 22.800 237.600 24.600 250.500 ;
        RECT 28.800 237.600 30.600 250.500 ;
        RECT 34.800 237.600 36.600 250.500 ;
        RECT 56.850 243.600 58.050 256.950 ;
        RECT 62.100 255.150 63.900 256.950 ;
        RECT 79.800 249.600 81.000 256.950 ;
        RECT 82.950 252.300 83.850 263.700 ;
        RECT 101.400 259.050 102.600 266.400 ;
        RECT 126.000 266.400 127.800 272.400 ;
        RECT 106.950 261.450 109.050 262.050 ;
        RECT 112.950 261.450 115.050 262.050 ;
        RECT 104.100 259.050 105.900 260.850 ;
        RECT 106.950 260.550 115.050 261.450 ;
        RECT 106.950 259.950 109.050 260.550 ;
        RECT 112.950 259.950 115.050 260.550 ;
        RECT 119.100 259.050 120.900 260.850 ;
        RECT 126.000 259.050 127.050 266.400 ;
        RECT 146.400 265.200 148.200 272.400 ;
        RECT 155.550 266.400 157.350 272.400 ;
        RECT 163.650 269.400 165.450 272.400 ;
        RECT 171.450 269.400 173.250 272.400 ;
        RECT 179.250 270.300 181.050 272.400 ;
        RECT 179.250 269.400 183.000 270.300 ;
        RECT 163.650 268.500 164.700 269.400 ;
        RECT 160.950 267.300 164.700 268.500 ;
        RECT 172.200 268.500 173.250 269.400 ;
        RECT 181.950 268.500 183.000 269.400 ;
        RECT 172.200 267.450 177.150 268.500 ;
        RECT 160.950 266.400 163.050 267.300 ;
        RECT 175.350 266.700 177.150 267.450 ;
        RECT 146.400 264.300 150.600 265.200 ;
        RECT 131.100 259.050 132.900 260.850 ;
        RECT 146.100 259.050 147.900 260.850 ;
        RECT 149.400 259.050 150.600 264.300 ;
        RECT 152.100 259.050 153.900 260.850 ;
        RECT 155.550 259.050 156.750 266.400 ;
        RECT 178.650 265.800 180.450 267.600 ;
        RECT 181.950 266.400 184.050 268.500 ;
        RECT 187.050 266.400 188.850 272.400 ;
        RECT 202.800 266.400 204.600 272.400 ;
        RECT 168.150 264.000 169.950 264.600 ;
        RECT 179.100 264.000 180.150 265.800 ;
        RECT 168.150 262.800 180.150 264.000 ;
        RECT 85.950 256.950 88.050 259.050 ;
        RECT 100.950 256.950 103.050 259.050 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 118.950 256.950 121.050 259.050 ;
        RECT 121.950 256.950 124.050 259.050 ;
        RECT 124.950 256.950 127.050 259.050 ;
        RECT 127.950 256.950 130.050 259.050 ;
        RECT 130.950 256.950 133.050 259.050 ;
        RECT 145.950 256.950 148.050 259.050 ;
        RECT 148.950 256.950 151.050 259.050 ;
        RECT 151.950 256.950 154.050 259.050 ;
        RECT 155.550 257.250 161.850 259.050 ;
        RECT 155.550 256.950 160.050 257.250 ;
        RECT 86.100 255.150 87.900 256.950 ;
        RECT 81.900 251.400 83.850 252.300 ;
        RECT 81.900 250.500 87.600 251.400 ;
        RECT 56.400 237.600 58.200 243.600 ;
        RECT 79.800 237.600 81.600 249.600 ;
        RECT 86.400 243.600 87.600 250.500 ;
        RECT 101.400 249.600 102.600 256.950 ;
        RECT 122.100 255.150 123.900 256.950 ;
        RECT 126.000 251.400 126.900 256.950 ;
        RECT 128.100 255.150 129.900 256.950 ;
        RECT 121.800 250.500 126.900 251.400 ;
        RECT 85.800 237.600 87.600 243.600 ;
        RECT 100.800 237.600 102.600 249.600 ;
        RECT 118.800 238.500 120.600 249.600 ;
        RECT 121.800 239.400 123.600 250.500 ;
        RECT 124.800 248.400 132.600 249.300 ;
        RECT 124.800 238.500 126.600 248.400 ;
        RECT 118.800 237.600 126.600 238.500 ;
        RECT 130.800 237.600 132.600 248.400 ;
        RECT 149.400 243.600 150.600 256.950 ;
        RECT 148.800 237.600 150.600 243.600 ;
        RECT 155.550 249.600 156.750 256.950 ;
        RECT 157.950 251.400 159.750 253.200 ;
        RECT 158.850 250.200 163.050 251.400 ;
        RECT 168.150 250.200 169.050 262.800 ;
        RECT 179.100 261.600 186.000 262.800 ;
        RECT 179.100 261.000 180.900 261.600 ;
        RECT 185.100 260.850 186.000 261.600 ;
        RECT 182.100 259.800 183.900 260.400 ;
        RECT 175.950 258.600 183.900 259.800 ;
        RECT 185.100 259.050 186.900 260.850 ;
        RECT 175.950 256.950 178.050 258.600 ;
        RECT 184.950 256.950 187.050 259.050 ;
        RECT 177.750 251.700 179.550 252.000 ;
        RECT 187.950 251.700 188.850 266.400 ;
        RECT 203.400 264.300 204.600 266.400 ;
        RECT 205.800 267.300 207.600 272.400 ;
        RECT 211.800 267.300 213.600 272.400 ;
        RECT 205.800 265.950 213.600 267.300 ;
        RECT 203.400 263.250 207.150 264.300 ;
        RECT 203.100 259.050 204.900 260.850 ;
        RECT 205.950 259.050 207.150 263.250 ;
        RECT 231.000 264.000 232.800 272.400 ;
        RECT 253.800 269.400 255.600 272.400 ;
        RECT 231.000 262.800 234.300 264.000 ;
        RECT 209.100 259.050 210.900 260.850 ;
        RECT 224.100 259.050 225.900 260.850 ;
        RECT 230.100 259.050 231.900 260.850 ;
        RECT 233.400 259.050 234.300 262.800 ;
        RECT 254.400 259.050 255.300 269.400 ;
        RECT 260.550 266.400 262.350 272.400 ;
        RECT 268.650 269.400 270.450 272.400 ;
        RECT 276.450 269.400 278.250 272.400 ;
        RECT 284.250 270.300 286.050 272.400 ;
        RECT 284.250 269.400 288.000 270.300 ;
        RECT 268.650 268.500 269.700 269.400 ;
        RECT 265.950 267.300 269.700 268.500 ;
        RECT 277.200 268.500 278.250 269.400 ;
        RECT 286.950 268.500 288.000 269.400 ;
        RECT 277.200 267.450 282.150 268.500 ;
        RECT 265.950 266.400 268.050 267.300 ;
        RECT 280.350 266.700 282.150 267.450 ;
        RECT 260.550 259.050 261.750 266.400 ;
        RECT 283.650 265.800 285.450 267.600 ;
        RECT 286.950 266.400 289.050 268.500 ;
        RECT 292.050 266.400 293.850 272.400 ;
        RECT 273.150 264.000 274.950 264.600 ;
        RECT 284.100 264.000 285.150 265.800 ;
        RECT 273.150 262.800 285.150 264.000 ;
        RECT 202.950 256.950 205.050 259.050 ;
        RECT 205.950 256.950 208.050 259.050 ;
        RECT 208.950 256.950 211.050 259.050 ;
        RECT 211.950 256.950 214.050 259.050 ;
        RECT 223.950 256.950 226.050 259.050 ;
        RECT 226.950 256.950 229.050 259.050 ;
        RECT 229.950 256.950 232.050 259.050 ;
        RECT 232.950 256.950 235.050 259.050 ;
        RECT 250.950 256.950 253.050 259.050 ;
        RECT 253.950 256.950 256.050 259.050 ;
        RECT 256.950 256.950 259.050 259.050 ;
        RECT 260.550 257.250 266.850 259.050 ;
        RECT 260.550 256.950 265.050 257.250 ;
        RECT 177.750 251.100 188.850 251.700 ;
        RECT 155.550 237.600 157.350 249.600 ;
        RECT 160.950 249.300 163.050 250.200 ;
        RECT 163.950 249.300 169.050 250.200 ;
        RECT 171.150 250.500 188.850 251.100 ;
        RECT 171.150 250.200 179.550 250.500 ;
        RECT 163.950 248.400 164.850 249.300 ;
        RECT 162.150 246.600 164.850 248.400 ;
        RECT 165.750 248.100 167.550 248.400 ;
        RECT 171.150 248.100 172.050 250.200 ;
        RECT 187.950 249.600 188.850 250.500 ;
        RECT 165.750 247.200 172.050 248.100 ;
        RECT 172.950 248.700 174.750 249.300 ;
        RECT 172.950 247.500 180.450 248.700 ;
        RECT 165.750 246.600 167.550 247.200 ;
        RECT 179.250 246.600 180.450 247.500 ;
        RECT 160.950 243.600 164.850 245.700 ;
        RECT 169.950 245.550 171.750 246.300 ;
        RECT 174.750 245.550 176.550 246.300 ;
        RECT 169.950 244.500 176.550 245.550 ;
        RECT 179.250 244.500 184.050 246.600 ;
        RECT 163.050 237.600 164.850 243.600 ;
        RECT 170.850 237.600 172.650 244.500 ;
        RECT 179.250 243.600 180.450 244.500 ;
        RECT 178.650 237.600 180.450 243.600 ;
        RECT 187.050 237.600 188.850 249.600 ;
        RECT 206.850 243.600 208.050 256.950 ;
        RECT 212.100 255.150 213.900 256.950 ;
        RECT 227.100 255.150 228.900 256.950 ;
        RECT 233.400 244.800 234.300 256.950 ;
        RECT 251.100 255.150 252.900 256.950 ;
        RECT 254.400 249.600 255.300 256.950 ;
        RECT 257.100 255.150 258.900 256.950 ;
        RECT 227.700 243.900 234.300 244.800 ;
        RECT 227.700 243.600 229.200 243.900 ;
        RECT 206.400 237.600 208.200 243.600 ;
        RECT 227.400 237.600 229.200 243.600 ;
        RECT 233.400 243.600 234.300 243.900 ;
        RECT 251.700 248.400 255.300 249.600 ;
        RECT 260.550 249.600 261.750 256.950 ;
        RECT 262.950 251.400 264.750 253.200 ;
        RECT 263.850 250.200 268.050 251.400 ;
        RECT 273.150 250.200 274.050 262.800 ;
        RECT 284.100 261.600 291.000 262.800 ;
        RECT 284.100 261.000 285.900 261.600 ;
        RECT 290.100 260.850 291.000 261.600 ;
        RECT 287.100 259.800 288.900 260.400 ;
        RECT 280.950 258.600 288.900 259.800 ;
        RECT 290.100 259.050 291.900 260.850 ;
        RECT 280.950 256.950 283.050 258.600 ;
        RECT 289.950 256.950 292.050 259.050 ;
        RECT 282.750 251.700 284.550 252.000 ;
        RECT 292.950 251.700 293.850 266.400 ;
        RECT 308.400 266.400 310.200 272.400 ;
        RECT 314.400 266.400 316.200 272.400 ;
        RECT 335.400 269.400 337.200 272.400 ;
        RECT 350.400 269.400 352.200 272.400 ;
        RECT 308.400 265.500 309.600 266.400 ;
        RECT 314.400 265.500 315.600 266.400 ;
        RECT 308.400 264.300 315.600 265.500 ;
        RECT 314.400 259.050 315.600 264.300 ;
        RECT 335.400 259.050 336.600 269.400 ;
        RECT 350.400 265.500 351.600 269.400 ;
        RECT 356.400 266.400 358.200 272.400 ;
        RECT 350.400 264.600 356.100 265.500 ;
        RECT 354.150 263.700 356.100 264.600 ;
        RECT 307.950 256.950 310.050 259.050 ;
        RECT 313.950 256.950 316.050 259.050 ;
        RECT 331.950 256.950 334.050 259.050 ;
        RECT 334.950 256.950 337.050 259.050 ;
        RECT 349.950 256.950 352.050 259.050 ;
        RECT 308.100 255.150 309.900 256.950 ;
        RECT 282.750 251.100 293.850 251.700 ;
        RECT 314.400 251.400 315.600 256.950 ;
        RECT 332.100 255.150 333.900 256.950 ;
        RECT 233.400 237.600 235.200 243.600 ;
        RECT 251.700 237.600 253.500 248.400 ;
        RECT 260.550 237.600 262.350 249.600 ;
        RECT 265.950 249.300 268.050 250.200 ;
        RECT 268.950 249.300 274.050 250.200 ;
        RECT 276.150 250.500 293.850 251.100 ;
        RECT 276.150 250.200 284.550 250.500 ;
        RECT 268.950 248.400 269.850 249.300 ;
        RECT 267.150 246.600 269.850 248.400 ;
        RECT 270.750 248.100 272.550 248.400 ;
        RECT 276.150 248.100 277.050 250.200 ;
        RECT 292.950 249.600 293.850 250.500 ;
        RECT 270.750 247.200 277.050 248.100 ;
        RECT 277.950 248.700 279.750 249.300 ;
        RECT 277.950 247.500 285.450 248.700 ;
        RECT 270.750 246.600 272.550 247.200 ;
        RECT 284.250 246.600 285.450 247.500 ;
        RECT 265.950 243.600 269.850 245.700 ;
        RECT 274.950 245.550 276.750 246.300 ;
        RECT 279.750 245.550 281.550 246.300 ;
        RECT 274.950 244.500 281.550 245.550 ;
        RECT 284.250 244.500 289.050 246.600 ;
        RECT 268.050 237.600 269.850 243.600 ;
        RECT 275.850 237.600 277.650 244.500 ;
        RECT 284.250 243.600 285.450 244.500 ;
        RECT 283.650 237.600 285.450 243.600 ;
        RECT 292.050 237.600 293.850 249.600 ;
        RECT 308.400 250.500 315.600 251.400 ;
        RECT 308.400 237.600 310.200 250.500 ;
        RECT 314.400 249.600 315.600 250.500 ;
        RECT 314.400 237.600 316.200 249.600 ;
        RECT 335.400 243.600 336.600 256.950 ;
        RECT 350.100 255.150 351.900 256.950 ;
        RECT 354.150 252.300 355.050 263.700 ;
        RECT 357.000 259.050 358.200 266.400 ;
        RECT 355.950 256.950 358.200 259.050 ;
        RECT 354.150 251.400 356.100 252.300 ;
        RECT 350.400 250.500 356.100 251.400 ;
        RECT 350.400 243.600 351.600 250.500 ;
        RECT 357.000 249.600 358.200 256.950 ;
        RECT 335.400 237.600 337.200 243.600 ;
        RECT 350.400 237.600 352.200 243.600 ;
        RECT 356.400 237.600 358.200 249.600 ;
        RECT 363.150 266.400 364.950 272.400 ;
        RECT 370.950 270.300 372.750 272.400 ;
        RECT 369.000 269.400 372.750 270.300 ;
        RECT 378.750 269.400 380.550 272.400 ;
        RECT 386.550 269.400 388.350 272.400 ;
        RECT 369.000 268.500 370.050 269.400 ;
        RECT 378.750 268.500 379.800 269.400 ;
        RECT 367.950 266.400 370.050 268.500 ;
        RECT 363.150 251.700 364.050 266.400 ;
        RECT 371.550 265.800 373.350 267.600 ;
        RECT 374.850 267.450 379.800 268.500 ;
        RECT 387.300 268.500 388.350 269.400 ;
        RECT 374.850 266.700 376.650 267.450 ;
        RECT 387.300 267.300 391.050 268.500 ;
        RECT 388.950 266.400 391.050 267.300 ;
        RECT 394.650 266.400 396.450 272.400 ;
        RECT 371.850 264.000 372.900 265.800 ;
        RECT 382.050 264.000 383.850 264.600 ;
        RECT 371.850 262.800 383.850 264.000 ;
        RECT 366.000 261.600 372.900 262.800 ;
        RECT 366.000 260.850 366.900 261.600 ;
        RECT 371.100 261.000 372.900 261.600 ;
        RECT 365.100 259.050 366.900 260.850 ;
        RECT 368.100 259.800 369.900 260.400 ;
        RECT 364.950 256.950 367.050 259.050 ;
        RECT 368.100 258.600 376.050 259.800 ;
        RECT 373.950 256.950 376.050 258.600 ;
        RECT 372.450 251.700 374.250 252.000 ;
        RECT 363.150 251.100 374.250 251.700 ;
        RECT 363.150 250.500 380.850 251.100 ;
        RECT 363.150 249.600 364.050 250.500 ;
        RECT 372.450 250.200 380.850 250.500 ;
        RECT 363.150 237.600 364.950 249.600 ;
        RECT 377.250 248.700 379.050 249.300 ;
        RECT 371.550 247.500 379.050 248.700 ;
        RECT 379.950 248.100 380.850 250.200 ;
        RECT 382.950 250.200 383.850 262.800 ;
        RECT 395.250 259.050 396.450 266.400 ;
        RECT 410.400 269.400 412.200 272.400 ;
        RECT 410.400 259.050 411.600 269.400 ;
        RECT 425.400 267.300 427.200 272.400 ;
        RECT 431.400 267.300 433.200 272.400 ;
        RECT 425.400 265.950 433.200 267.300 ;
        RECT 434.400 266.400 436.200 272.400 ;
        RECT 449.400 269.400 451.200 272.400 ;
        RECT 434.400 264.300 435.600 266.400 ;
        RECT 449.400 265.500 450.600 269.400 ;
        RECT 455.400 266.400 457.200 272.400 ;
        RECT 449.400 264.600 455.100 265.500 ;
        RECT 431.850 263.250 435.600 264.300 ;
        RECT 453.150 263.700 455.100 264.600 ;
        RECT 428.100 259.050 429.900 260.850 ;
        RECT 431.850 259.050 433.050 263.250 ;
        RECT 444.000 261.450 448.050 262.050 ;
        RECT 434.100 259.050 435.900 260.850 ;
        RECT 443.550 259.950 448.050 261.450 ;
        RECT 390.150 257.250 396.450 259.050 ;
        RECT 391.950 256.950 396.450 257.250 ;
        RECT 406.950 256.950 409.050 259.050 ;
        RECT 409.950 256.950 412.050 259.050 ;
        RECT 424.950 256.950 427.050 259.050 ;
        RECT 427.950 256.950 430.050 259.050 ;
        RECT 430.950 256.950 433.050 259.050 ;
        RECT 433.950 256.950 436.050 259.050 ;
        RECT 392.250 251.400 394.050 253.200 ;
        RECT 388.950 250.200 393.150 251.400 ;
        RECT 382.950 249.300 388.050 250.200 ;
        RECT 388.950 249.300 391.050 250.200 ;
        RECT 395.250 249.600 396.450 256.950 ;
        RECT 407.100 255.150 408.900 256.950 ;
        RECT 387.150 248.400 388.050 249.300 ;
        RECT 384.450 248.100 386.250 248.400 ;
        RECT 371.550 246.600 372.750 247.500 ;
        RECT 379.950 247.200 386.250 248.100 ;
        RECT 384.450 246.600 386.250 247.200 ;
        RECT 387.150 246.600 389.850 248.400 ;
        RECT 367.950 244.500 372.750 246.600 ;
        RECT 375.450 245.550 377.250 246.300 ;
        RECT 380.250 245.550 382.050 246.300 ;
        RECT 375.450 244.500 382.050 245.550 ;
        RECT 371.550 243.600 372.750 244.500 ;
        RECT 371.550 237.600 373.350 243.600 ;
        RECT 379.350 237.600 381.150 244.500 ;
        RECT 387.150 243.600 391.050 245.700 ;
        RECT 387.150 237.600 388.950 243.600 ;
        RECT 394.650 237.600 396.450 249.600 ;
        RECT 410.400 243.600 411.600 256.950 ;
        RECT 425.100 255.150 426.900 256.950 ;
        RECT 430.950 243.600 432.150 256.950 ;
        RECT 443.550 256.050 444.450 259.950 ;
        RECT 448.950 256.950 451.050 259.050 ;
        RECT 443.550 254.550 448.050 256.050 ;
        RECT 449.100 255.150 450.900 256.950 ;
        RECT 444.000 253.950 448.050 254.550 ;
        RECT 453.150 252.300 454.050 263.700 ;
        RECT 456.000 259.050 457.200 266.400 ;
        RECT 454.950 256.950 457.200 259.050 ;
        RECT 453.150 251.400 455.100 252.300 ;
        RECT 449.400 250.500 455.100 251.400 ;
        RECT 449.400 243.600 450.600 250.500 ;
        RECT 456.000 249.600 457.200 256.950 ;
        RECT 410.400 237.600 412.200 243.600 ;
        RECT 430.800 237.600 432.600 243.600 ;
        RECT 449.400 237.600 451.200 243.600 ;
        RECT 455.400 237.600 457.200 249.600 ;
        RECT 462.150 266.400 463.950 272.400 ;
        RECT 469.950 270.300 471.750 272.400 ;
        RECT 468.000 269.400 471.750 270.300 ;
        RECT 477.750 269.400 479.550 272.400 ;
        RECT 485.550 269.400 487.350 272.400 ;
        RECT 468.000 268.500 469.050 269.400 ;
        RECT 477.750 268.500 478.800 269.400 ;
        RECT 466.950 266.400 469.050 268.500 ;
        RECT 462.150 251.700 463.050 266.400 ;
        RECT 470.550 265.800 472.350 267.600 ;
        RECT 473.850 267.450 478.800 268.500 ;
        RECT 486.300 268.500 487.350 269.400 ;
        RECT 473.850 266.700 475.650 267.450 ;
        RECT 486.300 267.300 490.050 268.500 ;
        RECT 487.950 266.400 490.050 267.300 ;
        RECT 493.650 266.400 495.450 272.400 ;
        RECT 470.850 264.000 471.900 265.800 ;
        RECT 481.050 264.000 482.850 264.600 ;
        RECT 470.850 262.800 482.850 264.000 ;
        RECT 465.000 261.600 471.900 262.800 ;
        RECT 465.000 260.850 465.900 261.600 ;
        RECT 470.100 261.000 471.900 261.600 ;
        RECT 464.100 259.050 465.900 260.850 ;
        RECT 467.100 259.800 468.900 260.400 ;
        RECT 463.950 256.950 466.050 259.050 ;
        RECT 467.100 258.600 475.050 259.800 ;
        RECT 472.950 256.950 475.050 258.600 ;
        RECT 471.450 251.700 473.250 252.000 ;
        RECT 462.150 251.100 473.250 251.700 ;
        RECT 462.150 250.500 479.850 251.100 ;
        RECT 462.150 249.600 463.050 250.500 ;
        RECT 471.450 250.200 479.850 250.500 ;
        RECT 462.150 237.600 463.950 249.600 ;
        RECT 476.250 248.700 478.050 249.300 ;
        RECT 470.550 247.500 478.050 248.700 ;
        RECT 478.950 248.100 479.850 250.200 ;
        RECT 481.950 250.200 482.850 262.800 ;
        RECT 494.250 259.050 495.450 266.400 ;
        RECT 506.400 267.300 508.200 272.400 ;
        RECT 512.400 267.300 514.200 272.400 ;
        RECT 506.400 265.950 514.200 267.300 ;
        RECT 515.400 266.400 517.200 272.400 ;
        RECT 515.400 264.300 516.600 266.400 ;
        RECT 535.800 265.200 537.600 272.400 ;
        RECT 512.850 263.250 516.600 264.300 ;
        RECT 533.400 264.300 537.600 265.200 ;
        RECT 554.400 265.200 556.200 272.400 ;
        RECT 574.800 266.400 576.600 272.400 ;
        RECT 580.800 269.400 582.600 272.400 ;
        RECT 589.950 270.450 592.050 271.050 ;
        RECT 595.950 270.450 598.050 271.050 ;
        RECT 589.950 269.550 598.050 270.450 ;
        RECT 554.400 264.300 558.600 265.200 ;
        RECT 509.100 259.050 510.900 260.850 ;
        RECT 512.850 259.050 514.050 263.250 ;
        RECT 515.100 259.050 516.900 260.850 ;
        RECT 530.100 259.050 531.900 260.850 ;
        RECT 533.400 259.050 534.600 264.300 ;
        RECT 536.100 259.050 537.900 260.850 ;
        RECT 554.100 259.050 555.900 260.850 ;
        RECT 557.400 259.050 558.600 264.300 ;
        RECT 560.100 259.050 561.900 260.850 ;
        RECT 574.950 259.050 576.000 266.400 ;
        RECT 580.800 265.200 581.700 269.400 ;
        RECT 589.950 268.950 592.050 269.550 ;
        RECT 595.950 268.950 598.050 269.550 ;
        RECT 578.400 264.300 581.700 265.200 ;
        RECT 599.400 265.200 601.200 272.400 ;
        RECT 617.400 267.300 619.200 272.400 ;
        RECT 623.400 267.300 625.200 272.400 ;
        RECT 617.400 265.950 625.200 267.300 ;
        RECT 626.400 266.400 628.200 272.400 ;
        RECT 646.800 266.400 648.600 272.400 ;
        RECT 654.600 267.000 656.400 272.400 ;
        RECT 599.400 264.300 603.600 265.200 ;
        RECT 626.400 264.300 627.600 266.400 ;
        RECT 646.800 265.200 651.300 266.400 ;
        RECT 578.400 263.400 580.200 264.300 ;
        RECT 489.150 257.250 495.450 259.050 ;
        RECT 490.950 256.950 495.450 257.250 ;
        RECT 505.950 256.950 508.050 259.050 ;
        RECT 508.950 256.950 511.050 259.050 ;
        RECT 511.950 256.950 514.050 259.050 ;
        RECT 514.950 256.950 517.050 259.050 ;
        RECT 529.950 256.950 532.050 259.050 ;
        RECT 532.950 256.950 535.050 259.050 ;
        RECT 535.950 256.950 538.050 259.050 ;
        RECT 553.950 256.950 556.050 259.050 ;
        RECT 556.950 256.950 559.050 259.050 ;
        RECT 559.950 256.950 562.050 259.050 ;
        RECT 574.950 256.950 577.050 259.050 ;
        RECT 491.250 251.400 493.050 253.200 ;
        RECT 487.950 250.200 492.150 251.400 ;
        RECT 481.950 249.300 487.050 250.200 ;
        RECT 487.950 249.300 490.050 250.200 ;
        RECT 494.250 249.600 495.450 256.950 ;
        RECT 506.100 255.150 507.900 256.950 ;
        RECT 486.150 248.400 487.050 249.300 ;
        RECT 483.450 248.100 485.250 248.400 ;
        RECT 470.550 246.600 471.750 247.500 ;
        RECT 478.950 247.200 485.250 248.100 ;
        RECT 483.450 246.600 485.250 247.200 ;
        RECT 486.150 246.600 488.850 248.400 ;
        RECT 466.950 244.500 471.750 246.600 ;
        RECT 474.450 245.550 476.250 246.300 ;
        RECT 479.250 245.550 481.050 246.300 ;
        RECT 474.450 244.500 481.050 245.550 ;
        RECT 470.550 243.600 471.750 244.500 ;
        RECT 470.550 237.600 472.350 243.600 ;
        RECT 478.350 237.600 480.150 244.500 ;
        RECT 486.150 243.600 490.050 245.700 ;
        RECT 486.150 237.600 487.950 243.600 ;
        RECT 493.650 237.600 495.450 249.600 ;
        RECT 511.950 243.600 513.150 256.950 ;
        RECT 533.400 243.600 534.600 256.950 ;
        RECT 557.400 243.600 558.600 256.950 ;
        RECT 575.700 249.600 577.050 256.950 ;
        RECT 578.400 252.900 579.300 263.400 ;
        RECT 584.100 259.050 585.900 260.850 ;
        RECT 599.100 259.050 600.900 260.850 ;
        RECT 602.400 259.050 603.600 264.300 ;
        RECT 623.850 263.250 627.600 264.300 ;
        RECT 605.100 259.050 606.900 260.850 ;
        RECT 620.100 259.050 621.900 260.850 ;
        RECT 623.850 259.050 625.050 263.250 ;
        RECT 649.200 263.100 651.300 265.200 ;
        RECT 654.600 264.900 655.650 267.000 ;
        RECT 661.800 266.400 663.600 272.400 ;
        RECT 662.100 265.500 663.600 266.400 ;
        RECT 652.500 262.800 655.650 264.900 ;
        RECT 659.250 264.000 663.600 265.500 ;
        RECT 677.400 265.200 679.200 272.400 ;
        RECT 701.700 267.600 703.500 272.400 ;
        RECT 698.400 266.400 703.500 267.600 ;
        RECT 677.400 264.300 681.600 265.200 ;
        RECT 626.100 259.050 627.900 260.850 ;
        RECT 580.950 256.950 583.050 259.050 ;
        RECT 583.950 256.950 586.050 259.050 ;
        RECT 598.950 256.950 601.050 259.050 ;
        RECT 601.950 256.950 604.050 259.050 ;
        RECT 604.950 256.950 607.050 259.050 ;
        RECT 616.950 256.950 619.050 259.050 ;
        RECT 619.950 256.950 622.050 259.050 ;
        RECT 622.950 256.950 625.050 259.050 ;
        RECT 625.950 256.950 628.050 259.050 ;
        RECT 646.950 257.100 649.050 259.200 ;
        RECT 651.750 258.900 653.850 261.000 ;
        RECT 651.900 257.100 653.700 258.900 ;
        RECT 581.100 255.150 582.900 256.950 ;
        RECT 578.400 252.300 580.200 252.900 ;
        RECT 578.400 251.100 585.600 252.300 ;
        RECT 584.400 249.600 585.600 251.100 ;
        RECT 575.700 248.100 578.100 249.600 ;
        RECT 511.800 237.600 513.600 243.600 ;
        RECT 533.400 237.600 535.200 243.600 ;
        RECT 556.800 237.600 558.600 243.600 ;
        RECT 576.300 237.600 578.100 248.100 ;
        RECT 583.800 237.600 585.600 249.600 ;
        RECT 602.400 243.600 603.600 256.950 ;
        RECT 617.100 255.150 618.900 256.950 ;
        RECT 622.950 243.600 624.150 256.950 ;
        RECT 631.950 255.450 634.050 256.050 ;
        RECT 647.100 255.450 648.900 257.100 ;
        RECT 654.750 256.200 655.650 262.800 ;
        RECT 656.550 261.900 658.350 263.700 ;
        RECT 659.250 263.400 661.350 264.000 ;
        RECT 656.700 261.000 658.800 261.900 ;
        RECT 656.700 259.800 663.300 261.000 ;
        RECT 661.500 259.200 663.300 259.800 ;
        RECT 656.700 256.800 658.800 258.900 ;
        RECT 661.500 257.100 663.600 259.200 ;
        RECT 677.100 259.050 678.900 260.850 ;
        RECT 680.400 259.050 681.600 264.300 ;
        RECT 685.950 261.450 690.000 262.050 ;
        RECT 683.100 259.050 684.900 260.850 ;
        RECT 685.950 259.950 690.450 261.450 ;
        RECT 676.950 256.950 679.050 259.050 ;
        RECT 679.950 256.950 682.050 259.050 ;
        RECT 682.950 256.950 685.050 259.050 ;
        RECT 631.950 255.300 648.900 255.450 ;
        RECT 631.950 254.550 648.450 255.300 ;
        RECT 652.500 254.700 655.650 256.200 ;
        RECT 657.000 255.000 658.800 256.800 ;
        RECT 631.950 253.950 634.050 254.550 ;
        RECT 652.500 254.100 654.600 254.700 ;
        RECT 649.800 249.600 651.900 250.500 ;
        RECT 646.800 248.400 651.900 249.600 ;
        RECT 652.800 249.600 654.000 254.100 ;
        RECT 655.500 251.700 657.300 253.800 ;
        RECT 655.500 250.800 660.900 251.700 ;
        RECT 658.800 249.900 660.900 250.800 ;
        RECT 652.800 248.700 656.100 249.600 ;
        RECT 658.800 248.700 663.600 249.900 ;
        RECT 601.800 237.600 603.600 243.600 ;
        RECT 622.800 237.600 624.600 243.600 ;
        RECT 646.800 237.600 648.600 248.400 ;
        RECT 654.300 237.600 656.100 248.700 ;
        RECT 661.800 237.600 663.600 248.700 ;
        RECT 680.400 243.600 681.600 256.950 ;
        RECT 689.550 256.050 690.450 259.950 ;
        RECT 698.400 259.050 699.300 266.400 ;
        RECT 726.000 264.000 727.800 272.400 ;
        RECT 748.200 264.000 750.000 272.400 ;
        RECT 770.400 265.200 772.200 272.400 ;
        RECT 770.400 264.300 774.600 265.200 ;
        RECT 726.000 262.800 729.300 264.000 ;
        RECT 701.100 259.050 702.900 260.850 ;
        RECT 707.100 259.050 708.900 260.850 ;
        RECT 719.100 259.050 720.900 260.850 ;
        RECT 725.100 259.050 726.900 260.850 ;
        RECT 728.400 259.050 729.300 262.800 ;
        RECT 746.700 262.800 750.000 264.000 ;
        RECT 730.950 261.450 733.050 262.050 ;
        RECT 739.950 261.450 742.050 262.050 ;
        RECT 730.950 260.550 742.050 261.450 ;
        RECT 730.950 259.950 733.050 260.550 ;
        RECT 739.950 259.950 742.050 260.550 ;
        RECT 746.700 259.050 747.600 262.800 ;
        RECT 749.100 259.050 750.900 260.850 ;
        RECT 755.100 259.050 756.900 260.850 ;
        RECT 770.100 259.050 771.900 260.850 ;
        RECT 773.400 259.050 774.600 264.300 ;
        RECT 795.000 264.000 796.800 272.400 ;
        RECT 814.800 266.400 816.600 272.400 ;
        RECT 815.400 264.300 816.600 266.400 ;
        RECT 817.800 267.300 819.600 272.400 ;
        RECT 823.800 267.300 825.600 272.400 ;
        RECT 817.800 265.950 825.600 267.300 ;
        RECT 795.000 262.800 798.300 264.000 ;
        RECT 815.400 263.250 819.150 264.300 ;
        RECT 776.100 259.050 777.900 260.850 ;
        RECT 788.100 259.050 789.900 260.850 ;
        RECT 794.100 259.050 795.900 260.850 ;
        RECT 797.400 259.050 798.300 262.800 ;
        RECT 811.950 261.450 814.050 262.050 ;
        RECT 803.550 260.550 814.050 261.450 ;
        RECT 697.950 256.950 700.050 259.050 ;
        RECT 700.950 256.950 703.050 259.050 ;
        RECT 703.950 256.950 706.050 259.050 ;
        RECT 706.950 256.950 709.050 259.050 ;
        RECT 718.950 256.950 721.050 259.050 ;
        RECT 721.950 256.950 724.050 259.050 ;
        RECT 724.950 256.950 727.050 259.050 ;
        RECT 727.950 256.950 730.050 259.050 ;
        RECT 745.950 256.950 748.050 259.050 ;
        RECT 748.950 256.950 751.050 259.050 ;
        RECT 751.950 256.950 754.050 259.050 ;
        RECT 754.950 256.950 757.050 259.050 ;
        RECT 769.950 256.950 772.050 259.050 ;
        RECT 772.950 256.950 775.050 259.050 ;
        RECT 775.950 256.950 778.050 259.050 ;
        RECT 787.950 256.950 790.050 259.050 ;
        RECT 790.950 256.950 793.050 259.050 ;
        RECT 793.950 256.950 796.050 259.050 ;
        RECT 796.950 256.950 799.050 259.050 ;
        RECT 685.950 254.550 690.450 256.050 ;
        RECT 685.950 253.950 690.000 254.550 ;
        RECT 698.400 249.600 699.300 256.950 ;
        RECT 704.100 255.150 705.900 256.950 ;
        RECT 722.100 255.150 723.900 256.950 ;
        RECT 700.950 252.450 703.050 253.050 ;
        RECT 712.950 252.450 715.050 253.050 ;
        RECT 724.950 252.450 727.050 253.050 ;
        RECT 700.950 251.550 727.050 252.450 ;
        RECT 700.950 250.950 703.050 251.550 ;
        RECT 712.950 250.950 715.050 251.550 ;
        RECT 724.950 250.950 727.050 251.550 ;
        RECT 679.800 237.600 681.600 243.600 ;
        RECT 697.800 237.600 699.600 249.600 ;
        RECT 700.800 248.700 708.600 249.600 ;
        RECT 700.800 237.600 702.600 248.700 ;
        RECT 706.800 237.600 708.600 248.700 ;
        RECT 728.400 244.800 729.300 256.950 ;
        RECT 722.700 243.900 729.300 244.800 ;
        RECT 722.700 243.600 724.200 243.900 ;
        RECT 722.400 237.600 724.200 243.600 ;
        RECT 728.400 243.600 729.300 243.900 ;
        RECT 746.700 244.800 747.600 256.950 ;
        RECT 752.100 255.150 753.900 256.950 ;
        RECT 757.950 252.450 760.050 253.050 ;
        RECT 769.950 252.450 772.050 252.750 ;
        RECT 757.950 251.550 772.050 252.450 ;
        RECT 757.950 250.950 760.050 251.550 ;
        RECT 769.950 250.650 772.050 251.550 ;
        RECT 746.700 243.900 753.300 244.800 ;
        RECT 746.700 243.600 747.600 243.900 ;
        RECT 728.400 237.600 730.200 243.600 ;
        RECT 745.800 237.600 747.600 243.600 ;
        RECT 751.800 243.600 753.300 243.900 ;
        RECT 773.400 243.600 774.600 256.950 ;
        RECT 791.100 255.150 792.900 256.950 ;
        RECT 781.950 252.450 784.050 253.050 ;
        RECT 793.950 252.450 796.050 253.050 ;
        RECT 781.950 251.550 796.050 252.450 ;
        RECT 781.950 250.950 784.050 251.550 ;
        RECT 793.950 250.950 796.050 251.550 ;
        RECT 797.400 244.800 798.300 256.950 ;
        RECT 803.550 256.050 804.450 260.550 ;
        RECT 811.950 259.950 814.050 260.550 ;
        RECT 815.100 259.050 816.900 260.850 ;
        RECT 817.950 259.050 819.150 263.250 ;
        RECT 843.000 264.000 844.800 272.400 ;
        RECT 847.950 270.450 850.050 271.050 ;
        RECT 853.950 270.450 856.050 271.050 ;
        RECT 847.950 269.550 856.050 270.450 ;
        RECT 847.950 268.950 850.050 269.550 ;
        RECT 853.950 268.950 856.050 269.550 ;
        RECT 866.700 267.600 868.500 272.400 ;
        RECT 863.400 266.400 868.500 267.600 ;
        RECT 843.000 262.800 846.300 264.000 ;
        RECT 831.000 261.450 835.050 262.050 ;
        RECT 821.100 259.050 822.900 260.850 ;
        RECT 830.550 259.950 835.050 261.450 ;
        RECT 814.950 256.950 817.050 259.050 ;
        RECT 817.950 256.950 820.050 259.050 ;
        RECT 820.950 256.950 823.050 259.050 ;
        RECT 823.950 256.950 826.050 259.050 ;
        RECT 799.950 254.550 804.450 256.050 ;
        RECT 799.950 253.950 804.000 254.550 ;
        RECT 791.700 243.900 798.300 244.800 ;
        RECT 791.700 243.600 793.200 243.900 ;
        RECT 751.800 237.600 753.600 243.600 ;
        RECT 772.800 237.600 774.600 243.600 ;
        RECT 791.400 237.600 793.200 243.600 ;
        RECT 797.400 243.600 798.300 243.900 ;
        RECT 818.850 243.600 820.050 256.950 ;
        RECT 824.100 255.150 825.900 256.950 ;
        RECT 830.550 255.450 831.450 259.950 ;
        RECT 836.100 259.050 837.900 260.850 ;
        RECT 842.100 259.050 843.900 260.850 ;
        RECT 845.400 259.050 846.300 262.800 ;
        RECT 863.400 259.050 864.300 266.400 ;
        RECT 866.100 259.050 867.900 260.850 ;
        RECT 872.100 259.050 873.900 260.850 ;
        RECT 835.950 256.950 838.050 259.050 ;
        RECT 838.950 256.950 841.050 259.050 ;
        RECT 841.950 256.950 844.050 259.050 ;
        RECT 844.950 256.950 847.050 259.050 ;
        RECT 862.950 256.950 865.050 259.050 ;
        RECT 865.950 256.950 868.050 259.050 ;
        RECT 868.950 256.950 871.050 259.050 ;
        RECT 871.950 256.950 874.050 259.050 ;
        RECT 830.550 254.550 834.450 255.450 ;
        RECT 839.100 255.150 840.900 256.950 ;
        RECT 833.550 252.450 834.450 254.550 ;
        RECT 838.950 252.450 841.050 253.050 ;
        RECT 833.550 251.550 841.050 252.450 ;
        RECT 838.950 250.950 841.050 251.550 ;
        RECT 845.400 244.800 846.300 256.950 ;
        RECT 863.400 249.600 864.300 256.950 ;
        RECT 869.100 255.150 870.900 256.950 ;
        RECT 839.700 243.900 846.300 244.800 ;
        RECT 839.700 243.600 841.200 243.900 ;
        RECT 797.400 237.600 799.200 243.600 ;
        RECT 818.400 237.600 820.200 243.600 ;
        RECT 839.400 237.600 841.200 243.600 ;
        RECT 845.400 243.600 846.300 243.900 ;
        RECT 845.400 237.600 847.200 243.600 ;
        RECT 862.800 237.600 864.600 249.600 ;
        RECT 865.800 248.700 873.600 249.600 ;
        RECT 865.800 237.600 867.600 248.700 ;
        RECT 871.800 237.600 873.600 248.700 ;
        RECT 3.150 221.400 4.950 233.400 ;
        RECT 11.550 227.400 13.350 233.400 ;
        RECT 11.550 226.500 12.750 227.400 ;
        RECT 19.350 226.500 21.150 233.400 ;
        RECT 27.150 227.400 28.950 233.400 ;
        RECT 7.950 224.400 12.750 226.500 ;
        RECT 15.450 225.450 22.050 226.500 ;
        RECT 15.450 224.700 17.250 225.450 ;
        RECT 20.250 224.700 22.050 225.450 ;
        RECT 27.150 225.300 31.050 227.400 ;
        RECT 11.550 223.500 12.750 224.400 ;
        RECT 24.450 223.800 26.250 224.400 ;
        RECT 11.550 222.300 19.050 223.500 ;
        RECT 17.250 221.700 19.050 222.300 ;
        RECT 19.950 222.900 26.250 223.800 ;
        RECT 3.150 220.500 4.050 221.400 ;
        RECT 19.950 220.800 20.850 222.900 ;
        RECT 24.450 222.600 26.250 222.900 ;
        RECT 27.150 222.600 29.850 224.400 ;
        RECT 27.150 221.700 28.050 222.600 ;
        RECT 12.450 220.500 20.850 220.800 ;
        RECT 3.150 219.900 20.850 220.500 ;
        RECT 22.950 220.800 28.050 221.700 ;
        RECT 28.950 220.800 31.050 221.700 ;
        RECT 34.650 221.400 36.450 233.400 ;
        RECT 53.400 227.400 55.200 233.400 ;
        RECT 74.400 227.400 76.200 233.400 ;
        RECT 95.400 227.400 97.200 233.400 ;
        RECT 3.150 219.300 14.250 219.900 ;
        RECT 3.150 204.600 4.050 219.300 ;
        RECT 12.450 219.000 14.250 219.300 ;
        RECT 4.950 211.950 7.050 214.050 ;
        RECT 13.950 212.400 16.050 214.050 ;
        RECT 5.100 210.150 6.900 211.950 ;
        RECT 8.100 211.200 16.050 212.400 ;
        RECT 8.100 210.600 9.900 211.200 ;
        RECT 6.000 209.400 6.900 210.150 ;
        RECT 11.100 209.400 12.900 210.000 ;
        RECT 6.000 208.200 12.900 209.400 ;
        RECT 22.950 208.200 23.850 220.800 ;
        RECT 28.950 219.600 33.150 220.800 ;
        RECT 32.250 217.800 34.050 219.600 ;
        RECT 35.250 214.050 36.450 221.400 ;
        RECT 53.850 214.050 55.050 227.400 ;
        RECT 59.100 214.050 60.900 215.850 ;
        RECT 71.100 214.050 72.900 215.850 ;
        RECT 74.400 214.050 75.600 227.400 ;
        RECT 95.850 214.050 97.050 227.400 ;
        RECT 118.500 222.600 120.300 233.400 ;
        RECT 116.700 221.400 120.300 222.600 ;
        RECT 137.700 222.600 139.500 233.400 ;
        RECT 161.400 227.400 163.200 233.400 ;
        RECT 137.700 221.400 141.300 222.600 ;
        RECT 101.100 214.050 102.900 215.850 ;
        RECT 113.100 214.050 114.900 215.850 ;
        RECT 116.700 214.050 117.600 221.400 ;
        RECT 119.100 214.050 120.900 215.850 ;
        RECT 137.100 214.050 138.900 215.850 ;
        RECT 140.400 214.050 141.300 221.400 ;
        RECT 143.100 214.050 144.900 215.850 ;
        RECT 161.850 214.050 163.050 227.400 ;
        RECT 184.500 222.600 186.300 233.400 ;
        RECT 209.400 227.400 211.200 233.400 ;
        RECT 182.700 221.400 186.300 222.600 ;
        RECT 169.950 216.450 172.050 220.050 ;
        RECT 169.950 216.000 174.450 216.450 ;
        RECT 167.100 214.050 168.900 215.850 ;
        RECT 170.550 215.550 174.450 216.000 ;
        RECT 31.950 213.750 36.450 214.050 ;
        RECT 30.150 211.950 36.450 213.750 ;
        RECT 49.950 211.950 52.050 214.050 ;
        RECT 52.950 211.950 55.050 214.050 ;
        RECT 55.950 211.950 58.050 214.050 ;
        RECT 58.950 211.950 61.050 214.050 ;
        RECT 70.950 211.950 73.050 214.050 ;
        RECT 73.950 211.950 76.050 214.050 ;
        RECT 91.950 211.950 94.050 214.050 ;
        RECT 94.950 211.950 97.050 214.050 ;
        RECT 97.950 211.950 100.050 214.050 ;
        RECT 100.950 211.950 103.050 214.050 ;
        RECT 112.950 211.950 115.050 214.050 ;
        RECT 115.950 211.950 118.050 214.050 ;
        RECT 118.950 211.950 121.050 214.050 ;
        RECT 136.950 211.950 139.050 214.050 ;
        RECT 139.950 211.950 142.050 214.050 ;
        RECT 142.950 211.950 145.050 214.050 ;
        RECT 157.950 211.950 160.050 214.050 ;
        RECT 160.950 211.950 163.050 214.050 ;
        RECT 163.950 211.950 166.050 214.050 ;
        RECT 166.950 211.950 169.050 214.050 ;
        RECT 11.850 207.000 23.850 208.200 ;
        RECT 11.850 205.200 12.900 207.000 ;
        RECT 22.050 206.400 23.850 207.000 ;
        RECT 3.150 198.600 4.950 204.600 ;
        RECT 7.950 202.500 10.050 204.600 ;
        RECT 11.550 203.400 13.350 205.200 ;
        RECT 35.250 204.600 36.450 211.950 ;
        RECT 50.100 210.150 51.900 211.950 ;
        RECT 52.950 207.750 54.150 211.950 ;
        RECT 56.100 210.150 57.900 211.950 ;
        RECT 50.400 206.700 54.150 207.750 ;
        RECT 64.950 207.450 67.050 208.050 ;
        RECT 70.950 207.450 73.050 208.050 ;
        RECT 50.400 204.600 51.600 206.700 ;
        RECT 64.950 206.550 73.050 207.450 ;
        RECT 64.950 205.950 67.050 206.550 ;
        RECT 70.950 205.950 73.050 206.550 ;
        RECT 14.850 203.550 16.650 204.300 ;
        RECT 28.950 203.700 31.050 204.600 ;
        RECT 14.850 202.500 19.800 203.550 ;
        RECT 9.000 201.600 10.050 202.500 ;
        RECT 18.750 201.600 19.800 202.500 ;
        RECT 27.300 202.500 31.050 203.700 ;
        RECT 27.300 201.600 28.350 202.500 ;
        RECT 9.000 200.700 12.750 201.600 ;
        RECT 10.950 198.600 12.750 200.700 ;
        RECT 18.750 198.600 20.550 201.600 ;
        RECT 26.550 198.600 28.350 201.600 ;
        RECT 34.650 198.600 36.450 204.600 ;
        RECT 49.800 198.600 51.600 204.600 ;
        RECT 52.800 203.700 60.600 205.050 ;
        RECT 52.800 198.600 54.600 203.700 ;
        RECT 58.800 198.600 60.600 203.700 ;
        RECT 74.400 201.600 75.600 211.950 ;
        RECT 92.100 210.150 93.900 211.950 ;
        RECT 94.950 207.750 96.150 211.950 ;
        RECT 98.100 210.150 99.900 211.950 ;
        RECT 92.400 206.700 96.150 207.750 ;
        RECT 92.400 204.600 93.600 206.700 ;
        RECT 74.400 198.600 76.200 201.600 ;
        RECT 91.800 198.600 93.600 204.600 ;
        RECT 94.800 203.700 102.600 205.050 ;
        RECT 94.800 198.600 96.600 203.700 ;
        RECT 100.800 198.600 102.600 203.700 ;
        RECT 116.700 201.600 117.600 211.950 ;
        RECT 140.400 201.600 141.300 211.950 ;
        RECT 158.100 210.150 159.900 211.950 ;
        RECT 160.950 207.750 162.150 211.950 ;
        RECT 164.100 210.150 165.900 211.950 ;
        RECT 158.400 206.700 162.150 207.750 ;
        RECT 173.550 207.450 174.450 215.550 ;
        RECT 179.100 214.050 180.900 215.850 ;
        RECT 182.700 214.050 183.600 221.400 ;
        RECT 185.100 214.050 186.900 215.850 ;
        RECT 209.850 214.050 211.050 227.400 ;
        RECT 218.550 221.400 220.350 233.400 ;
        RECT 226.050 227.400 227.850 233.400 ;
        RECT 223.950 225.300 227.850 227.400 ;
        RECT 233.850 226.500 235.650 233.400 ;
        RECT 241.650 227.400 243.450 233.400 ;
        RECT 242.250 226.500 243.450 227.400 ;
        RECT 232.950 225.450 239.550 226.500 ;
        RECT 232.950 224.700 234.750 225.450 ;
        RECT 237.750 224.700 239.550 225.450 ;
        RECT 242.250 224.400 247.050 226.500 ;
        RECT 225.150 222.600 227.850 224.400 ;
        RECT 228.750 223.800 230.550 224.400 ;
        RECT 228.750 222.900 235.050 223.800 ;
        RECT 242.250 223.500 243.450 224.400 ;
        RECT 228.750 222.600 230.550 222.900 ;
        RECT 226.950 221.700 227.850 222.600 ;
        RECT 215.100 214.050 216.900 215.850 ;
        RECT 218.550 214.050 219.750 221.400 ;
        RECT 223.950 220.800 226.050 221.700 ;
        RECT 226.950 220.800 232.050 221.700 ;
        RECT 221.850 219.600 226.050 220.800 ;
        RECT 220.950 217.800 222.750 219.600 ;
        RECT 178.950 211.950 181.050 214.050 ;
        RECT 181.950 211.950 184.050 214.050 ;
        RECT 184.950 211.950 187.050 214.050 ;
        RECT 205.950 211.950 208.050 214.050 ;
        RECT 208.950 211.950 211.050 214.050 ;
        RECT 211.950 211.950 214.050 214.050 ;
        RECT 214.950 211.950 217.050 214.050 ;
        RECT 218.550 213.750 223.050 214.050 ;
        RECT 218.550 211.950 224.850 213.750 ;
        RECT 178.950 207.450 181.050 207.750 ;
        RECT 158.400 204.600 159.600 206.700 ;
        RECT 173.550 206.550 181.050 207.450 ;
        RECT 178.950 205.650 181.050 206.550 ;
        RECT 116.400 198.600 118.200 201.600 ;
        RECT 139.800 198.600 141.600 201.600 ;
        RECT 157.800 198.600 159.600 204.600 ;
        RECT 160.800 203.700 168.600 205.050 ;
        RECT 160.800 198.600 162.600 203.700 ;
        RECT 166.800 198.600 168.600 203.700 ;
        RECT 182.700 201.600 183.600 211.950 ;
        RECT 206.100 210.150 207.900 211.950 ;
        RECT 208.950 207.750 210.150 211.950 ;
        RECT 212.100 210.150 213.900 211.950 ;
        RECT 206.400 206.700 210.150 207.750 ;
        RECT 206.400 204.600 207.600 206.700 ;
        RECT 182.400 198.600 184.200 201.600 ;
        RECT 205.800 198.600 207.600 204.600 ;
        RECT 208.800 203.700 216.600 205.050 ;
        RECT 208.800 198.600 210.600 203.700 ;
        RECT 214.800 198.600 216.600 203.700 ;
        RECT 218.550 204.600 219.750 211.950 ;
        RECT 231.150 208.200 232.050 220.800 ;
        RECT 234.150 220.800 235.050 222.900 ;
        RECT 235.950 222.300 243.450 223.500 ;
        RECT 235.950 221.700 237.750 222.300 ;
        RECT 250.050 221.400 251.850 233.400 ;
        RECT 234.150 220.500 242.550 220.800 ;
        RECT 250.950 220.500 251.850 221.400 ;
        RECT 234.150 219.900 251.850 220.500 ;
        RECT 240.750 219.300 251.850 219.900 ;
        RECT 240.750 219.000 242.550 219.300 ;
        RECT 238.950 212.400 241.050 214.050 ;
        RECT 238.950 211.200 246.900 212.400 ;
        RECT 247.950 211.950 250.050 214.050 ;
        RECT 245.100 210.600 246.900 211.200 ;
        RECT 248.100 210.150 249.900 211.950 ;
        RECT 242.100 209.400 243.900 210.000 ;
        RECT 248.100 209.400 249.000 210.150 ;
        RECT 242.100 208.200 249.000 209.400 ;
        RECT 231.150 207.000 243.150 208.200 ;
        RECT 231.150 206.400 232.950 207.000 ;
        RECT 242.100 205.200 243.150 207.000 ;
        RECT 218.550 198.600 220.350 204.600 ;
        RECT 223.950 203.700 226.050 204.600 ;
        RECT 223.950 202.500 227.700 203.700 ;
        RECT 238.350 203.550 240.150 204.300 ;
        RECT 226.650 201.600 227.700 202.500 ;
        RECT 235.200 202.500 240.150 203.550 ;
        RECT 241.650 203.400 243.450 205.200 ;
        RECT 250.950 204.600 251.850 219.300 ;
        RECT 266.400 227.400 268.200 233.400 ;
        RECT 290.400 227.400 292.200 233.400 ;
        RECT 314.400 227.400 316.200 233.400 ;
        RECT 266.400 214.050 267.600 227.400 ;
        RECT 290.850 214.050 292.050 227.400 ;
        RECT 296.100 214.050 297.900 215.850 ;
        RECT 314.850 214.050 316.050 227.400 ;
        RECT 335.700 222.600 337.500 233.400 ;
        RECT 355.800 227.400 357.600 233.400 ;
        RECT 335.700 221.400 339.300 222.600 ;
        RECT 320.100 214.050 321.900 215.850 ;
        RECT 335.100 214.050 336.900 215.850 ;
        RECT 338.400 214.050 339.300 221.400 ;
        RECT 341.100 214.050 342.900 215.850 ;
        RECT 356.400 214.050 357.600 227.400 ;
        RECT 373.800 221.400 375.600 233.400 ;
        RECT 379.800 227.400 381.600 233.400 ;
        RECT 359.100 214.050 360.900 215.850 ;
        RECT 374.400 214.050 375.300 221.400 ;
        RECT 377.100 214.050 378.900 215.850 ;
        RECT 262.950 211.950 265.050 214.050 ;
        RECT 265.950 211.950 268.050 214.050 ;
        RECT 268.950 211.950 271.050 214.050 ;
        RECT 286.950 211.950 289.050 214.050 ;
        RECT 289.950 211.950 292.050 214.050 ;
        RECT 292.950 211.950 295.050 214.050 ;
        RECT 295.950 211.950 298.050 214.050 ;
        RECT 310.950 211.950 313.050 214.050 ;
        RECT 313.950 211.950 316.050 214.050 ;
        RECT 316.950 211.950 319.050 214.050 ;
        RECT 319.950 211.950 322.050 214.050 ;
        RECT 334.950 211.950 337.050 214.050 ;
        RECT 337.950 211.950 340.050 214.050 ;
        RECT 340.950 211.950 343.050 214.050 ;
        RECT 355.950 211.950 358.050 214.050 ;
        RECT 358.950 211.950 361.050 214.050 ;
        RECT 373.950 211.950 376.050 214.050 ;
        RECT 376.950 211.950 379.050 214.050 ;
        RECT 263.100 210.150 264.900 211.950 ;
        RECT 266.400 206.700 267.600 211.950 ;
        RECT 269.100 210.150 270.900 211.950 ;
        RECT 287.100 210.150 288.900 211.950 ;
        RECT 289.950 207.750 291.150 211.950 ;
        RECT 293.100 210.150 294.900 211.950 ;
        RECT 311.100 210.150 312.900 211.950 ;
        RECT 313.950 207.750 315.150 211.950 ;
        RECT 317.100 210.150 318.900 211.950 ;
        RECT 287.400 206.700 291.150 207.750 ;
        RECT 311.400 206.700 315.150 207.750 ;
        RECT 266.400 205.800 270.600 206.700 ;
        RECT 244.950 202.500 247.050 204.600 ;
        RECT 235.200 201.600 236.250 202.500 ;
        RECT 244.950 201.600 246.000 202.500 ;
        RECT 226.650 198.600 228.450 201.600 ;
        RECT 234.450 198.600 236.250 201.600 ;
        RECT 242.250 200.700 246.000 201.600 ;
        RECT 242.250 198.600 244.050 200.700 ;
        RECT 250.050 198.600 251.850 204.600 ;
        RECT 268.800 198.600 270.600 205.800 ;
        RECT 287.400 204.600 288.600 206.700 ;
        RECT 286.800 198.600 288.600 204.600 ;
        RECT 289.800 203.700 297.600 205.050 ;
        RECT 311.400 204.600 312.600 206.700 ;
        RECT 289.800 198.600 291.600 203.700 ;
        RECT 295.800 198.600 297.600 203.700 ;
        RECT 310.800 198.600 312.600 204.600 ;
        RECT 313.800 203.700 321.600 205.050 ;
        RECT 313.800 198.600 315.600 203.700 ;
        RECT 319.800 198.600 321.600 203.700 ;
        RECT 338.400 201.600 339.300 211.950 ;
        RECT 356.400 201.600 357.600 211.950 ;
        RECT 374.400 204.600 375.300 211.950 ;
        RECT 380.700 207.300 381.600 227.400 ;
        RECT 399.300 222.900 401.100 233.400 ;
        RECT 398.700 221.400 401.100 222.900 ;
        RECT 406.800 221.400 408.600 233.400 ;
        RECT 398.700 214.050 400.050 221.400 ;
        RECT 407.400 219.900 408.600 221.400 ;
        RECT 422.400 227.400 424.200 233.400 ;
        RECT 382.950 211.950 385.050 214.050 ;
        RECT 397.950 211.950 400.050 214.050 ;
        RECT 401.400 218.700 408.600 219.900 ;
        RECT 412.950 219.450 415.050 220.050 ;
        RECT 418.950 219.450 421.050 220.200 ;
        RECT 401.400 218.100 403.200 218.700 ;
        RECT 412.950 218.550 421.050 219.450 ;
        RECT 383.100 210.150 384.900 211.950 ;
        RECT 377.100 206.400 384.600 207.300 ;
        RECT 377.100 205.500 378.900 206.400 ;
        RECT 374.400 202.800 377.100 204.600 ;
        RECT 337.800 198.600 339.600 201.600 ;
        RECT 355.800 198.600 357.600 201.600 ;
        RECT 375.300 198.600 377.100 202.800 ;
        RECT 382.800 198.600 384.600 206.400 ;
        RECT 397.950 204.600 399.000 211.950 ;
        RECT 401.400 207.600 402.300 218.100 ;
        RECT 412.950 217.950 415.050 218.550 ;
        RECT 418.950 218.100 421.050 218.550 ;
        RECT 404.100 214.050 405.900 215.850 ;
        RECT 422.400 214.050 423.600 227.400 ;
        RECT 432.150 221.400 433.950 233.400 ;
        RECT 440.550 227.400 442.350 233.400 ;
        RECT 440.550 226.500 441.750 227.400 ;
        RECT 448.350 226.500 450.150 233.400 ;
        RECT 456.150 227.400 457.950 233.400 ;
        RECT 436.950 224.400 441.750 226.500 ;
        RECT 444.450 225.450 451.050 226.500 ;
        RECT 444.450 224.700 446.250 225.450 ;
        RECT 449.250 224.700 451.050 225.450 ;
        RECT 456.150 225.300 460.050 227.400 ;
        RECT 440.550 223.500 441.750 224.400 ;
        RECT 453.450 223.800 455.250 224.400 ;
        RECT 440.550 222.300 448.050 223.500 ;
        RECT 446.250 221.700 448.050 222.300 ;
        RECT 448.950 222.900 455.250 223.800 ;
        RECT 432.150 220.500 433.050 221.400 ;
        RECT 448.950 220.800 449.850 222.900 ;
        RECT 453.450 222.600 455.250 222.900 ;
        RECT 456.150 222.600 458.850 224.400 ;
        RECT 456.150 221.700 457.050 222.600 ;
        RECT 441.450 220.500 449.850 220.800 ;
        RECT 432.150 219.900 449.850 220.500 ;
        RECT 451.950 220.800 457.050 221.700 ;
        RECT 457.950 220.800 460.050 221.700 ;
        RECT 463.650 221.400 465.450 233.400 ;
        RECT 432.150 219.300 443.250 219.900 ;
        RECT 403.950 211.950 406.050 214.050 ;
        RECT 406.950 211.950 409.050 214.050 ;
        RECT 418.950 211.950 421.050 214.050 ;
        RECT 421.950 211.950 424.050 214.050 ;
        RECT 424.950 211.950 427.050 214.050 ;
        RECT 407.100 210.150 408.900 211.950 ;
        RECT 419.100 210.150 420.900 211.950 ;
        RECT 401.400 206.700 403.200 207.600 ;
        RECT 422.400 206.700 423.600 211.950 ;
        RECT 425.100 210.150 426.900 211.950 ;
        RECT 401.400 205.800 404.700 206.700 ;
        RECT 422.400 205.800 426.600 206.700 ;
        RECT 397.800 198.600 399.600 204.600 ;
        RECT 403.800 201.600 404.700 205.800 ;
        RECT 403.800 198.600 405.600 201.600 ;
        RECT 424.800 198.600 426.600 205.800 ;
        RECT 432.150 204.600 433.050 219.300 ;
        RECT 441.450 219.000 443.250 219.300 ;
        RECT 433.950 211.950 436.050 214.050 ;
        RECT 442.950 212.400 445.050 214.050 ;
        RECT 434.100 210.150 435.900 211.950 ;
        RECT 437.100 211.200 445.050 212.400 ;
        RECT 437.100 210.600 438.900 211.200 ;
        RECT 435.000 209.400 435.900 210.150 ;
        RECT 440.100 209.400 441.900 210.000 ;
        RECT 435.000 208.200 441.900 209.400 ;
        RECT 451.950 208.200 452.850 220.800 ;
        RECT 457.950 219.600 462.150 220.800 ;
        RECT 461.250 217.800 463.050 219.600 ;
        RECT 464.250 214.050 465.450 221.400 ;
        RECT 479.400 227.400 481.200 233.400 ;
        RECT 499.800 227.400 501.600 233.400 ;
        RECT 521.400 227.400 523.200 233.400 ;
        RECT 476.100 214.050 477.900 215.850 ;
        RECT 479.400 214.050 480.600 227.400 ;
        RECT 494.100 214.050 495.900 215.850 ;
        RECT 499.950 214.050 501.150 227.400 ;
        RECT 505.950 216.450 510.000 217.050 ;
        RECT 505.950 214.950 510.450 216.450 ;
        RECT 460.950 213.750 465.450 214.050 ;
        RECT 459.150 211.950 465.450 213.750 ;
        RECT 475.950 211.950 478.050 214.050 ;
        RECT 478.950 211.950 481.050 214.050 ;
        RECT 493.950 211.950 496.050 214.050 ;
        RECT 496.950 211.950 499.050 214.050 ;
        RECT 499.950 211.950 502.050 214.050 ;
        RECT 502.950 211.950 505.050 214.050 ;
        RECT 440.850 207.000 452.850 208.200 ;
        RECT 440.850 205.200 441.900 207.000 ;
        RECT 451.050 206.400 452.850 207.000 ;
        RECT 432.150 198.600 433.950 204.600 ;
        RECT 436.950 202.500 439.050 204.600 ;
        RECT 440.550 203.400 442.350 205.200 ;
        RECT 464.250 204.600 465.450 211.950 ;
        RECT 443.850 203.550 445.650 204.300 ;
        RECT 457.950 203.700 460.050 204.600 ;
        RECT 443.850 202.500 448.800 203.550 ;
        RECT 438.000 201.600 439.050 202.500 ;
        RECT 447.750 201.600 448.800 202.500 ;
        RECT 456.300 202.500 460.050 203.700 ;
        RECT 456.300 201.600 457.350 202.500 ;
        RECT 438.000 200.700 441.750 201.600 ;
        RECT 439.950 198.600 441.750 200.700 ;
        RECT 447.750 198.600 449.550 201.600 ;
        RECT 455.550 198.600 457.350 201.600 ;
        RECT 463.650 198.600 465.450 204.600 ;
        RECT 479.400 201.600 480.600 211.950 ;
        RECT 497.100 210.150 498.900 211.950 ;
        RECT 484.950 207.450 487.050 207.900 ;
        RECT 490.950 207.450 493.050 208.050 ;
        RECT 484.950 206.550 493.050 207.450 ;
        RECT 500.850 207.750 502.050 211.950 ;
        RECT 503.100 210.150 504.900 211.950 ;
        RECT 509.550 210.450 510.450 214.950 ;
        RECT 521.400 214.050 522.600 227.400 ;
        RECT 530.550 221.400 532.350 233.400 ;
        RECT 538.050 227.400 539.850 233.400 ;
        RECT 535.950 225.300 539.850 227.400 ;
        RECT 545.850 226.500 547.650 233.400 ;
        RECT 553.650 227.400 555.450 233.400 ;
        RECT 554.250 226.500 555.450 227.400 ;
        RECT 544.950 225.450 551.550 226.500 ;
        RECT 544.950 224.700 546.750 225.450 ;
        RECT 549.750 224.700 551.550 225.450 ;
        RECT 554.250 224.400 559.050 226.500 ;
        RECT 537.150 222.600 539.850 224.400 ;
        RECT 540.750 223.800 542.550 224.400 ;
        RECT 540.750 222.900 547.050 223.800 ;
        RECT 554.250 223.500 555.450 224.400 ;
        RECT 540.750 222.600 542.550 222.900 ;
        RECT 538.950 221.700 539.850 222.600 ;
        RECT 530.550 214.050 531.750 221.400 ;
        RECT 535.950 220.800 538.050 221.700 ;
        RECT 538.950 220.800 544.050 221.700 ;
        RECT 533.850 219.600 538.050 220.800 ;
        RECT 532.950 217.800 534.750 219.600 ;
        RECT 517.950 211.950 520.050 214.050 ;
        RECT 520.950 211.950 523.050 214.050 ;
        RECT 523.950 211.950 526.050 214.050 ;
        RECT 530.550 213.750 535.050 214.050 ;
        RECT 530.550 211.950 536.850 213.750 ;
        RECT 514.950 210.450 517.050 211.050 ;
        RECT 509.550 209.550 517.050 210.450 ;
        RECT 518.100 210.150 519.900 211.950 ;
        RECT 514.950 208.950 517.050 209.550 ;
        RECT 500.850 206.700 504.600 207.750 ;
        RECT 484.950 205.800 487.050 206.550 ;
        RECT 490.950 205.950 493.050 206.550 ;
        RECT 494.400 203.700 502.200 205.050 ;
        RECT 479.400 198.600 481.200 201.600 ;
        RECT 494.400 198.600 496.200 203.700 ;
        RECT 500.400 198.600 502.200 203.700 ;
        RECT 503.400 204.600 504.600 206.700 ;
        RECT 521.400 206.700 522.600 211.950 ;
        RECT 524.100 210.150 525.900 211.950 ;
        RECT 521.400 205.800 525.600 206.700 ;
        RECT 503.400 198.600 505.200 204.600 ;
        RECT 523.800 198.600 525.600 205.800 ;
        RECT 530.550 204.600 531.750 211.950 ;
        RECT 543.150 208.200 544.050 220.800 ;
        RECT 546.150 220.800 547.050 222.900 ;
        RECT 547.950 222.300 555.450 223.500 ;
        RECT 547.950 221.700 549.750 222.300 ;
        RECT 562.050 221.400 563.850 233.400 ;
        RECT 546.150 220.500 554.550 220.800 ;
        RECT 562.950 220.500 563.850 221.400 ;
        RECT 546.150 219.900 563.850 220.500 ;
        RECT 552.750 219.300 563.850 219.900 ;
        RECT 552.750 219.000 554.550 219.300 ;
        RECT 550.950 212.400 553.050 214.050 ;
        RECT 550.950 211.200 558.900 212.400 ;
        RECT 559.950 211.950 562.050 214.050 ;
        RECT 557.100 210.600 558.900 211.200 ;
        RECT 560.100 210.150 561.900 211.950 ;
        RECT 554.100 209.400 555.900 210.000 ;
        RECT 560.100 209.400 561.000 210.150 ;
        RECT 554.100 208.200 561.000 209.400 ;
        RECT 543.150 207.000 555.150 208.200 ;
        RECT 543.150 206.400 544.950 207.000 ;
        RECT 554.100 205.200 555.150 207.000 ;
        RECT 530.550 198.600 532.350 204.600 ;
        RECT 535.950 203.700 538.050 204.600 ;
        RECT 535.950 202.500 539.700 203.700 ;
        RECT 550.350 203.550 552.150 204.300 ;
        RECT 538.650 201.600 539.700 202.500 ;
        RECT 547.200 202.500 552.150 203.550 ;
        RECT 553.650 203.400 555.450 205.200 ;
        RECT 562.950 204.600 563.850 219.300 ;
        RECT 581.400 227.400 583.200 233.400 ;
        RECT 605.400 227.400 607.200 233.400 ;
        RECT 626.400 227.400 628.200 233.400 ;
        RECT 581.400 214.050 582.600 227.400 ;
        RECT 605.850 214.050 607.050 227.400 ;
        RECT 610.950 219.450 613.050 220.050 ;
        RECT 616.950 219.450 619.050 220.050 ;
        RECT 610.950 218.550 619.050 219.450 ;
        RECT 610.950 217.950 613.050 218.550 ;
        RECT 616.950 217.950 619.050 218.550 ;
        RECT 611.100 214.050 612.900 215.850 ;
        RECT 577.950 211.950 580.050 214.050 ;
        RECT 580.950 211.950 583.050 214.050 ;
        RECT 583.950 211.950 586.050 214.050 ;
        RECT 601.950 211.950 604.050 214.050 ;
        RECT 604.950 211.950 607.050 214.050 ;
        RECT 607.950 211.950 610.050 214.050 ;
        RECT 610.950 211.950 613.050 214.050 ;
        RECT 622.950 211.950 625.050 214.050 ;
        RECT 578.100 210.150 579.900 211.950 ;
        RECT 581.400 206.700 582.600 211.950 ;
        RECT 584.100 210.150 585.900 211.950 ;
        RECT 602.100 210.150 603.900 211.950 ;
        RECT 604.950 207.750 606.150 211.950 ;
        RECT 608.100 210.150 609.900 211.950 ;
        RECT 623.100 210.150 624.900 211.950 ;
        RECT 602.400 206.700 606.150 207.750 ;
        RECT 626.400 207.300 627.300 227.400 ;
        RECT 632.400 221.400 634.200 233.400 ;
        RECT 650.400 227.400 652.200 233.400 ;
        RECT 629.100 214.050 630.900 215.850 ;
        RECT 632.700 214.050 633.600 221.400 ;
        RECT 628.950 211.950 631.050 214.050 ;
        RECT 631.950 211.950 634.050 214.050 ;
        RECT 646.950 211.950 649.050 214.050 ;
        RECT 581.400 205.800 585.600 206.700 ;
        RECT 556.950 202.500 559.050 204.600 ;
        RECT 547.200 201.600 548.250 202.500 ;
        RECT 556.950 201.600 558.000 202.500 ;
        RECT 538.650 198.600 540.450 201.600 ;
        RECT 546.450 198.600 548.250 201.600 ;
        RECT 554.250 200.700 558.000 201.600 ;
        RECT 554.250 198.600 556.050 200.700 ;
        RECT 562.050 198.600 563.850 204.600 ;
        RECT 583.800 198.600 585.600 205.800 ;
        RECT 602.400 204.600 603.600 206.700 ;
        RECT 623.400 206.400 630.900 207.300 ;
        RECT 601.800 198.600 603.600 204.600 ;
        RECT 604.800 203.700 612.600 205.050 ;
        RECT 604.800 198.600 606.600 203.700 ;
        RECT 610.800 198.600 612.600 203.700 ;
        RECT 623.400 198.600 625.200 206.400 ;
        RECT 629.100 205.500 630.900 206.400 ;
        RECT 632.700 204.600 633.600 211.950 ;
        RECT 647.100 210.150 648.900 211.950 ;
        RECT 650.400 207.300 651.300 227.400 ;
        RECT 656.400 221.400 658.200 233.400 ;
        RECT 673.800 221.400 675.600 233.400 ;
        RECT 676.800 222.300 678.600 233.400 ;
        RECT 682.800 222.300 684.600 233.400 ;
        RECT 676.800 221.400 684.600 222.300 ;
        RECT 695.400 222.300 697.200 233.400 ;
        RECT 695.400 221.400 699.900 222.300 ;
        RECT 702.900 221.400 704.700 233.400 ;
        RECT 710.400 222.600 712.200 233.400 ;
        RECT 653.100 214.050 654.900 215.850 ;
        RECT 656.700 214.050 657.600 221.400 ;
        RECT 674.400 214.050 675.300 221.400 ;
        RECT 697.800 219.300 699.900 221.400 ;
        RECT 703.500 219.900 704.700 221.400 ;
        RECT 707.400 221.400 712.200 222.600 ;
        RECT 727.800 222.600 729.600 233.400 ;
        RECT 727.800 221.400 732.600 222.600 ;
        RECT 707.400 220.500 709.500 221.400 ;
        RECT 730.500 220.500 732.600 221.400 ;
        RECT 735.300 221.400 737.100 233.400 ;
        RECT 742.800 222.300 744.600 233.400 ;
        RECT 740.100 221.400 744.600 222.300 ;
        RECT 757.800 221.400 759.600 233.400 ;
        RECT 760.800 222.300 762.600 233.400 ;
        RECT 766.800 222.300 768.600 233.400 ;
        RECT 781.800 227.400 783.600 233.400 ;
        RECT 760.800 221.400 768.600 222.300 ;
        RECT 735.300 219.900 736.500 221.400 ;
        RECT 703.500 219.000 705.000 219.900 ;
        RECT 701.100 217.500 703.200 217.800 ;
        RECT 685.950 216.450 688.050 217.050 ;
        RECT 680.100 214.050 681.900 215.850 ;
        RECT 685.950 215.550 693.450 216.450 ;
        RECT 699.300 215.700 703.200 217.500 ;
        RECT 704.100 216.900 705.000 219.000 ;
        RECT 735.000 219.000 736.500 219.900 ;
        RECT 740.100 219.300 742.200 221.400 ;
        RECT 735.000 216.900 735.900 219.000 ;
        RECT 685.950 214.950 688.050 215.550 ;
        RECT 652.950 211.950 655.050 214.050 ;
        RECT 655.950 211.950 658.050 214.050 ;
        RECT 673.950 211.950 676.050 214.050 ;
        RECT 676.950 211.950 679.050 214.050 ;
        RECT 679.950 211.950 682.050 214.050 ;
        RECT 682.950 211.950 685.050 214.050 ;
        RECT 692.550 213.450 693.450 215.550 ;
        RECT 704.100 214.800 706.200 216.900 ;
        RECT 695.400 213.900 697.500 214.050 ;
        RECT 700.500 213.900 702.300 214.500 ;
        RECT 695.400 213.450 702.300 213.900 ;
        RECT 692.550 212.700 702.300 213.450 ;
        RECT 703.200 213.900 705.600 214.800 ;
        RECT 710.100 214.050 711.900 215.850 ;
        RECT 728.100 214.050 729.900 215.850 ;
        RECT 733.800 214.800 735.900 216.900 ;
        RECT 736.800 217.500 738.900 217.800 ;
        RECT 736.800 215.700 740.700 217.500 ;
        RECT 692.550 212.550 697.500 212.700 ;
        RECT 695.400 211.950 697.500 212.550 ;
        RECT 630.900 202.800 633.600 204.600 ;
        RECT 647.400 206.400 654.900 207.300 ;
        RECT 630.900 198.600 632.700 202.800 ;
        RECT 634.950 201.450 637.050 202.050 ;
        RECT 643.950 201.450 646.050 202.050 ;
        RECT 634.950 200.550 646.050 201.450 ;
        RECT 634.950 199.950 637.050 200.550 ;
        RECT 643.950 199.950 646.050 200.550 ;
        RECT 647.400 198.600 649.200 206.400 ;
        RECT 653.100 205.500 654.900 206.400 ;
        RECT 656.700 204.600 657.600 211.950 ;
        RECT 654.900 202.800 657.600 204.600 ;
        RECT 674.400 204.600 675.300 211.950 ;
        RECT 677.100 210.150 678.900 211.950 ;
        RECT 683.100 210.150 684.900 211.950 ;
        RECT 695.400 210.150 697.200 211.950 ;
        RECT 700.500 209.400 702.300 211.200 ;
        RECT 700.200 207.300 702.300 209.400 ;
        RECT 696.000 206.400 702.300 207.300 ;
        RECT 703.200 208.200 704.250 213.900 ;
        RECT 709.950 213.450 712.050 214.050 ;
        RECT 714.000 213.450 717.900 214.050 ;
        RECT 705.600 211.200 707.400 213.000 ;
        RECT 709.950 212.550 717.900 213.450 ;
        RECT 709.950 211.950 712.050 212.550 ;
        RECT 714.000 211.950 717.900 212.550 ;
        RECT 718.950 213.450 721.050 214.050 ;
        RECT 727.950 213.450 730.050 214.050 ;
        RECT 734.400 213.900 736.800 214.800 ;
        RECT 718.950 212.550 730.050 213.450 ;
        RECT 718.950 211.950 721.050 212.550 ;
        RECT 727.950 211.950 730.050 212.550 ;
        RECT 732.600 211.200 734.400 213.000 ;
        RECT 705.150 209.100 707.250 211.200 ;
        RECT 732.750 209.100 734.850 211.200 ;
        RECT 735.750 208.200 736.800 213.900 ;
        RECT 737.700 213.900 739.500 214.500 ;
        RECT 758.400 214.050 759.300 221.400 ;
        RECT 760.950 219.450 763.050 220.200 ;
        RECT 772.950 219.450 775.050 220.050 ;
        RECT 760.950 218.550 775.050 219.450 ;
        RECT 760.950 218.100 763.050 218.550 ;
        RECT 772.950 217.950 775.050 218.550 ;
        RECT 764.100 214.050 765.900 215.850 ;
        RECT 782.400 214.050 783.600 227.400 ;
        RECT 800.400 227.400 802.200 233.400 ;
        RECT 787.950 216.450 792.000 217.050 ;
        RECT 785.100 214.050 786.900 215.850 ;
        RECT 787.950 214.950 792.450 216.450 ;
        RECT 742.500 213.900 744.600 214.050 ;
        RECT 737.700 212.700 744.600 213.900 ;
        RECT 742.500 211.950 744.600 212.700 ;
        RECT 757.950 211.950 760.050 214.050 ;
        RECT 760.950 211.950 763.050 214.050 ;
        RECT 763.950 211.950 766.050 214.050 ;
        RECT 766.950 211.950 769.050 214.050 ;
        RECT 781.950 211.950 784.050 214.050 ;
        RECT 784.950 211.950 787.050 214.050 ;
        RECT 696.000 204.600 697.200 206.400 ;
        RECT 703.200 206.100 706.200 208.200 ;
        RECT 703.200 204.600 704.400 206.100 ;
        RECT 707.400 205.500 709.500 206.700 ;
        RECT 730.500 205.500 732.600 206.700 ;
        RECT 733.800 206.100 736.800 208.200 ;
        RECT 737.700 209.400 739.500 211.200 ;
        RECT 742.800 210.450 744.600 211.950 ;
        RECT 754.950 210.450 757.050 211.050 ;
        RECT 742.800 210.150 757.050 210.450 ;
        RECT 743.550 209.550 757.050 210.150 ;
        RECT 737.700 207.300 739.800 209.400 ;
        RECT 754.950 208.950 757.050 209.550 ;
        RECT 737.700 206.400 744.000 207.300 ;
        RECT 707.400 204.600 712.200 205.500 ;
        RECT 674.400 203.400 679.500 204.600 ;
        RECT 654.900 198.600 656.700 202.800 ;
        RECT 677.700 198.600 679.500 203.400 ;
        RECT 695.400 198.600 697.200 204.600 ;
        RECT 702.900 198.600 704.700 204.600 ;
        RECT 710.400 198.600 712.200 204.600 ;
        RECT 727.800 204.600 732.600 205.500 ;
        RECT 735.600 204.600 736.800 206.100 ;
        RECT 742.800 204.600 744.000 206.400 ;
        RECT 758.400 204.600 759.300 211.950 ;
        RECT 761.100 210.150 762.900 211.950 ;
        RECT 767.100 210.150 768.900 211.950 ;
        RECT 760.950 207.450 763.050 208.050 ;
        RECT 769.950 207.450 772.050 208.050 ;
        RECT 760.950 206.550 772.050 207.450 ;
        RECT 760.950 205.950 763.050 206.550 ;
        RECT 769.950 205.950 772.050 206.550 ;
        RECT 727.800 198.600 729.600 204.600 ;
        RECT 735.300 198.600 737.100 204.600 ;
        RECT 742.800 198.600 744.600 204.600 ;
        RECT 758.400 203.400 763.500 204.600 ;
        RECT 761.700 198.600 763.500 203.400 ;
        RECT 782.400 201.600 783.600 211.950 ;
        RECT 791.550 211.050 792.450 214.950 ;
        RECT 800.400 214.050 801.600 227.400 ;
        RECT 820.800 221.400 822.600 233.400 ;
        RECT 826.800 227.400 828.600 233.400 ;
        RECT 845.400 227.400 847.200 233.400 ;
        RECT 821.400 214.050 822.300 221.400 ;
        RECT 824.100 214.050 825.900 215.850 ;
        RECT 796.950 211.950 799.050 214.050 ;
        RECT 799.950 211.950 802.050 214.050 ;
        RECT 802.950 211.950 805.050 214.050 ;
        RECT 820.950 211.950 823.050 214.050 ;
        RECT 823.950 211.950 826.050 214.050 ;
        RECT 791.550 209.550 796.050 211.050 ;
        RECT 797.100 210.150 798.900 211.950 ;
        RECT 792.000 208.950 796.050 209.550 ;
        RECT 800.400 206.700 801.600 211.950 ;
        RECT 803.100 210.150 804.900 211.950 ;
        RECT 800.400 205.800 804.600 206.700 ;
        RECT 781.800 198.600 783.600 201.600 ;
        RECT 802.800 198.600 804.600 205.800 ;
        RECT 821.400 204.600 822.300 211.950 ;
        RECT 827.700 207.300 828.600 227.400 ;
        RECT 845.700 227.100 847.200 227.400 ;
        RECT 851.400 227.400 853.200 233.400 ;
        RECT 872.400 227.400 874.200 233.400 ;
        RECT 851.400 227.100 852.300 227.400 ;
        RECT 845.700 226.200 852.300 227.100 ;
        RECT 845.100 214.050 846.900 215.850 ;
        RECT 851.400 214.050 852.300 226.200 ;
        RECT 864.000 216.450 868.050 217.050 ;
        RECT 863.550 214.950 868.050 216.450 ;
        RECT 829.950 211.950 832.050 214.050 ;
        RECT 841.950 211.950 844.050 214.050 ;
        RECT 844.950 211.950 847.050 214.050 ;
        RECT 847.950 211.950 850.050 214.050 ;
        RECT 850.950 211.950 853.050 214.050 ;
        RECT 830.100 210.150 831.900 211.950 ;
        RECT 842.100 210.150 843.900 211.950 ;
        RECT 848.100 210.150 849.900 211.950 ;
        RECT 851.400 208.200 852.300 211.950 ;
        RECT 863.550 211.050 864.450 214.950 ;
        RECT 872.850 214.050 874.050 227.400 ;
        RECT 878.100 214.050 879.900 215.850 ;
        RECT 868.950 211.950 871.050 214.050 ;
        RECT 871.950 211.950 874.050 214.050 ;
        RECT 874.950 211.950 877.050 214.050 ;
        RECT 877.950 211.950 880.050 214.050 ;
        RECT 863.550 209.550 868.050 211.050 ;
        RECT 869.100 210.150 870.900 211.950 ;
        RECT 864.000 208.950 868.050 209.550 ;
        RECT 824.100 206.400 831.600 207.300 ;
        RECT 824.100 205.500 825.900 206.400 ;
        RECT 821.400 202.800 824.100 204.600 ;
        RECT 822.300 198.600 824.100 202.800 ;
        RECT 829.800 198.600 831.600 206.400 ;
        RECT 849.000 207.000 852.300 208.200 ;
        RECT 871.950 207.750 873.150 211.950 ;
        RECT 875.100 210.150 876.900 211.950 ;
        RECT 849.000 198.600 850.800 207.000 ;
        RECT 869.400 206.700 873.150 207.750 ;
        RECT 869.400 204.600 870.600 206.700 ;
        RECT 868.800 198.600 870.600 204.600 ;
        RECT 871.800 203.700 879.600 205.050 ;
        RECT 871.800 198.600 873.600 203.700 ;
        RECT 877.800 198.600 879.600 203.700 ;
        RECT 13.800 188.400 15.600 194.400 ;
        RECT 14.400 186.300 15.600 188.400 ;
        RECT 16.800 189.300 18.600 194.400 ;
        RECT 22.800 189.300 24.600 194.400 ;
        RECT 16.800 187.950 24.600 189.300 ;
        RECT 40.800 187.200 42.600 194.400 ;
        RECT 58.800 188.400 60.600 194.400 ;
        RECT 38.400 186.300 42.600 187.200 ;
        RECT 59.400 186.300 60.600 188.400 ;
        RECT 61.800 189.300 63.600 194.400 ;
        RECT 67.800 189.300 69.600 194.400 ;
        RECT 61.800 187.950 69.600 189.300 ;
        RECT 80.400 189.300 82.200 194.400 ;
        RECT 86.400 189.300 88.200 194.400 ;
        RECT 80.400 187.950 88.200 189.300 ;
        RECT 89.400 188.400 91.200 194.400 ;
        RECT 95.550 188.400 97.350 194.400 ;
        RECT 103.650 191.400 105.450 194.400 ;
        RECT 111.450 191.400 113.250 194.400 ;
        RECT 119.250 192.300 121.050 194.400 ;
        RECT 119.250 191.400 123.000 192.300 ;
        RECT 103.650 190.500 104.700 191.400 ;
        RECT 100.950 189.300 104.700 190.500 ;
        RECT 112.200 190.500 113.250 191.400 ;
        RECT 121.950 190.500 123.000 191.400 ;
        RECT 112.200 189.450 117.150 190.500 ;
        RECT 100.950 188.400 103.050 189.300 ;
        RECT 115.350 188.700 117.150 189.450 ;
        RECT 89.400 186.300 90.600 188.400 ;
        RECT 14.400 185.250 18.150 186.300 ;
        RECT 14.100 181.050 15.900 182.850 ;
        RECT 16.950 181.050 18.150 185.250 ;
        RECT 20.100 181.050 21.900 182.850 ;
        RECT 35.100 181.050 36.900 182.850 ;
        RECT 38.400 181.050 39.600 186.300 ;
        RECT 59.400 185.250 63.150 186.300 ;
        RECT 41.100 181.050 42.900 182.850 ;
        RECT 59.100 181.050 60.900 182.850 ;
        RECT 61.950 181.050 63.150 185.250 ;
        RECT 86.850 185.250 90.600 186.300 ;
        RECT 65.100 181.050 66.900 182.850 ;
        RECT 83.100 181.050 84.900 182.850 ;
        RECT 86.850 181.050 88.050 185.250 ;
        RECT 89.100 181.050 90.900 182.850 ;
        RECT 95.550 181.050 96.750 188.400 ;
        RECT 118.650 187.800 120.450 189.600 ;
        RECT 121.950 188.400 124.050 190.500 ;
        RECT 127.050 188.400 128.850 194.400 ;
        RECT 108.150 186.000 109.950 186.600 ;
        RECT 119.100 186.000 120.150 187.800 ;
        RECT 108.150 184.800 120.150 186.000 ;
        RECT 13.950 178.950 16.050 181.050 ;
        RECT 16.950 178.950 19.050 181.050 ;
        RECT 19.950 178.950 22.050 181.050 ;
        RECT 22.950 178.950 25.050 181.050 ;
        RECT 34.950 178.950 37.050 181.050 ;
        RECT 37.950 178.950 40.050 181.050 ;
        RECT 40.950 178.950 43.050 181.050 ;
        RECT 58.950 178.950 61.050 181.050 ;
        RECT 61.950 178.950 64.050 181.050 ;
        RECT 64.950 178.950 67.050 181.050 ;
        RECT 67.950 178.950 70.050 181.050 ;
        RECT 79.950 178.950 82.050 181.050 ;
        RECT 82.950 178.950 85.050 181.050 ;
        RECT 85.950 178.950 88.050 181.050 ;
        RECT 88.950 178.950 91.050 181.050 ;
        RECT 95.550 179.250 101.850 181.050 ;
        RECT 95.550 178.950 100.050 179.250 ;
        RECT 17.850 165.600 19.050 178.950 ;
        RECT 23.100 177.150 24.900 178.950 ;
        RECT 38.400 165.600 39.600 178.950 ;
        RECT 62.850 165.600 64.050 178.950 ;
        RECT 68.100 177.150 69.900 178.950 ;
        RECT 80.100 177.150 81.900 178.950 ;
        RECT 85.950 165.600 87.150 178.950 ;
        RECT 95.550 171.600 96.750 178.950 ;
        RECT 97.950 173.400 99.750 175.200 ;
        RECT 98.850 172.200 103.050 173.400 ;
        RECT 108.150 172.200 109.050 184.800 ;
        RECT 119.100 183.600 126.000 184.800 ;
        RECT 119.100 183.000 120.900 183.600 ;
        RECT 125.100 182.850 126.000 183.600 ;
        RECT 122.100 181.800 123.900 182.400 ;
        RECT 115.950 180.600 123.900 181.800 ;
        RECT 125.100 181.050 126.900 182.850 ;
        RECT 115.950 178.950 118.050 180.600 ;
        RECT 124.950 178.950 127.050 181.050 ;
        RECT 117.750 173.700 119.550 174.000 ;
        RECT 127.950 173.700 128.850 188.400 ;
        RECT 145.800 187.200 147.600 194.400 ;
        RECT 163.800 188.400 165.600 194.400 ;
        RECT 143.400 186.300 147.600 187.200 ;
        RECT 164.400 186.300 165.600 188.400 ;
        RECT 166.800 189.300 168.600 194.400 ;
        RECT 172.800 189.300 174.600 194.400 ;
        RECT 166.800 187.950 174.600 189.300 ;
        RECT 190.800 187.200 192.600 194.400 ;
        RECT 188.400 186.300 192.600 187.200 ;
        RECT 209.400 187.200 211.200 194.400 ;
        RECT 218.550 188.400 220.350 194.400 ;
        RECT 226.650 191.400 228.450 194.400 ;
        RECT 234.450 191.400 236.250 194.400 ;
        RECT 242.250 192.300 244.050 194.400 ;
        RECT 242.250 191.400 246.000 192.300 ;
        RECT 226.650 190.500 227.700 191.400 ;
        RECT 223.950 189.300 227.700 190.500 ;
        RECT 235.200 190.500 236.250 191.400 ;
        RECT 244.950 190.500 246.000 191.400 ;
        RECT 235.200 189.450 240.150 190.500 ;
        RECT 223.950 188.400 226.050 189.300 ;
        RECT 238.350 188.700 240.150 189.450 ;
        RECT 209.400 186.300 213.600 187.200 ;
        RECT 140.100 181.050 141.900 182.850 ;
        RECT 143.400 181.050 144.600 186.300 ;
        RECT 164.400 185.250 168.150 186.300 ;
        RECT 146.100 181.050 147.900 182.850 ;
        RECT 164.100 181.050 165.900 182.850 ;
        RECT 166.950 181.050 168.150 185.250 ;
        RECT 180.000 183.450 184.050 184.050 ;
        RECT 170.100 181.050 171.900 182.850 ;
        RECT 179.550 181.950 184.050 183.450 ;
        RECT 139.950 178.950 142.050 181.050 ;
        RECT 142.950 178.950 145.050 181.050 ;
        RECT 145.950 178.950 148.050 181.050 ;
        RECT 163.950 178.950 166.050 181.050 ;
        RECT 166.950 178.950 169.050 181.050 ;
        RECT 169.950 178.950 172.050 181.050 ;
        RECT 172.950 178.950 175.050 181.050 ;
        RECT 117.750 173.100 128.850 173.700 ;
        RECT 17.400 159.600 19.200 165.600 ;
        RECT 38.400 159.600 40.200 165.600 ;
        RECT 62.400 159.600 64.200 165.600 ;
        RECT 85.800 159.600 87.600 165.600 ;
        RECT 95.550 159.600 97.350 171.600 ;
        RECT 100.950 171.300 103.050 172.200 ;
        RECT 103.950 171.300 109.050 172.200 ;
        RECT 111.150 172.500 128.850 173.100 ;
        RECT 130.950 174.450 133.050 175.050 ;
        RECT 136.950 174.450 139.050 175.050 ;
        RECT 130.950 173.550 139.050 174.450 ;
        RECT 130.950 172.950 133.050 173.550 ;
        RECT 136.950 172.950 139.050 173.550 ;
        RECT 111.150 172.200 119.550 172.500 ;
        RECT 103.950 170.400 104.850 171.300 ;
        RECT 102.150 168.600 104.850 170.400 ;
        RECT 105.750 170.100 107.550 170.400 ;
        RECT 111.150 170.100 112.050 172.200 ;
        RECT 127.950 171.600 128.850 172.500 ;
        RECT 105.750 169.200 112.050 170.100 ;
        RECT 112.950 170.700 114.750 171.300 ;
        RECT 112.950 169.500 120.450 170.700 ;
        RECT 105.750 168.600 107.550 169.200 ;
        RECT 119.250 168.600 120.450 169.500 ;
        RECT 100.950 165.600 104.850 167.700 ;
        RECT 109.950 167.550 111.750 168.300 ;
        RECT 114.750 167.550 116.550 168.300 ;
        RECT 109.950 166.500 116.550 167.550 ;
        RECT 119.250 166.500 124.050 168.600 ;
        RECT 103.050 159.600 104.850 165.600 ;
        RECT 110.850 159.600 112.650 166.500 ;
        RECT 119.250 165.600 120.450 166.500 ;
        RECT 118.650 159.600 120.450 165.600 ;
        RECT 127.050 159.600 128.850 171.600 ;
        RECT 143.400 165.600 144.600 178.950 ;
        RECT 167.850 165.600 169.050 178.950 ;
        RECT 173.100 177.150 174.900 178.950 ;
        RECT 179.550 177.450 180.450 181.950 ;
        RECT 185.100 181.050 186.900 182.850 ;
        RECT 188.400 181.050 189.600 186.300 ;
        RECT 191.100 181.050 192.900 182.850 ;
        RECT 209.100 181.050 210.900 182.850 ;
        RECT 212.400 181.050 213.600 186.300 ;
        RECT 215.100 181.050 216.900 182.850 ;
        RECT 218.550 181.050 219.750 188.400 ;
        RECT 241.650 187.800 243.450 189.600 ;
        RECT 244.950 188.400 247.050 190.500 ;
        RECT 250.050 188.400 251.850 194.400 ;
        RECT 265.800 188.400 267.600 194.400 ;
        RECT 231.150 186.000 232.950 186.600 ;
        RECT 242.100 186.000 243.150 187.800 ;
        RECT 231.150 184.800 243.150 186.000 ;
        RECT 184.950 178.950 187.050 181.050 ;
        RECT 187.950 178.950 190.050 181.050 ;
        RECT 190.950 178.950 193.050 181.050 ;
        RECT 208.950 178.950 211.050 181.050 ;
        RECT 211.950 178.950 214.050 181.050 ;
        RECT 214.950 178.950 217.050 181.050 ;
        RECT 218.550 179.250 224.850 181.050 ;
        RECT 218.550 178.950 223.050 179.250 ;
        RECT 176.550 177.000 180.450 177.450 ;
        RECT 175.950 176.550 180.450 177.000 ;
        RECT 175.950 172.950 178.050 176.550 ;
        RECT 188.400 165.600 189.600 178.950 ;
        RECT 199.950 174.450 202.050 175.050 ;
        RECT 208.950 174.450 211.050 175.050 ;
        RECT 199.950 173.550 211.050 174.450 ;
        RECT 199.950 172.950 202.050 173.550 ;
        RECT 208.950 172.950 211.050 173.550 ;
        RECT 212.400 165.600 213.600 178.950 ;
        RECT 143.400 159.600 145.200 165.600 ;
        RECT 167.400 159.600 169.200 165.600 ;
        RECT 188.400 159.600 190.200 165.600 ;
        RECT 211.800 159.600 213.600 165.600 ;
        RECT 218.550 171.600 219.750 178.950 ;
        RECT 220.950 173.400 222.750 175.200 ;
        RECT 221.850 172.200 226.050 173.400 ;
        RECT 231.150 172.200 232.050 184.800 ;
        RECT 242.100 183.600 249.000 184.800 ;
        RECT 242.100 183.000 243.900 183.600 ;
        RECT 248.100 182.850 249.000 183.600 ;
        RECT 245.100 181.800 246.900 182.400 ;
        RECT 238.950 180.600 246.900 181.800 ;
        RECT 248.100 181.050 249.900 182.850 ;
        RECT 238.950 178.950 241.050 180.600 ;
        RECT 247.950 178.950 250.050 181.050 ;
        RECT 240.750 173.700 242.550 174.000 ;
        RECT 250.950 173.700 251.850 188.400 ;
        RECT 266.400 186.300 267.600 188.400 ;
        RECT 268.800 189.300 270.600 194.400 ;
        RECT 274.800 189.300 276.600 194.400 ;
        RECT 293.700 189.600 295.500 194.400 ;
        RECT 316.800 191.400 318.600 194.400 ;
        RECT 268.800 187.950 276.600 189.300 ;
        RECT 290.400 188.400 295.500 189.600 ;
        RECT 266.400 185.250 270.150 186.300 ;
        RECT 266.100 181.050 267.900 182.850 ;
        RECT 268.950 181.050 270.150 185.250 ;
        RECT 272.100 181.050 273.900 182.850 ;
        RECT 290.400 181.050 291.300 188.400 ;
        RECT 293.100 181.050 294.900 182.850 ;
        RECT 299.100 181.050 300.900 182.850 ;
        RECT 317.400 181.050 318.300 191.400 ;
        RECT 334.800 188.400 336.600 194.400 ;
        RECT 342.300 188.400 344.100 194.400 ;
        RECT 349.800 188.400 351.600 194.400 ;
        RECT 362.400 189.300 364.200 194.400 ;
        RECT 368.400 189.300 370.200 194.400 ;
        RECT 334.800 187.500 339.600 188.400 ;
        RECT 337.500 186.300 339.600 187.500 ;
        RECT 342.600 186.900 343.800 188.400 ;
        RECT 340.800 184.800 343.800 186.900 ;
        RECT 349.800 186.600 351.000 188.400 ;
        RECT 362.400 187.950 370.200 189.300 ;
        RECT 371.400 188.400 373.200 194.400 ;
        RECT 388.800 191.400 390.600 194.400 ;
        RECT 339.750 181.800 341.850 183.900 ;
        RECT 265.950 178.950 268.050 181.050 ;
        RECT 268.950 178.950 271.050 181.050 ;
        RECT 271.950 178.950 274.050 181.050 ;
        RECT 274.950 178.950 277.050 181.050 ;
        RECT 289.950 178.950 292.050 181.050 ;
        RECT 292.950 178.950 295.050 181.050 ;
        RECT 295.950 178.950 298.050 181.050 ;
        RECT 298.950 178.950 301.050 181.050 ;
        RECT 313.950 178.950 316.050 181.050 ;
        RECT 316.950 178.950 319.050 181.050 ;
        RECT 319.950 178.950 322.050 181.050 ;
        RECT 325.950 180.450 328.050 181.050 ;
        RECT 334.950 180.450 337.050 181.050 ;
        RECT 325.950 179.550 337.050 180.450 ;
        RECT 339.600 180.000 341.400 181.800 ;
        RECT 325.950 178.950 328.050 179.550 ;
        RECT 334.950 178.950 337.050 179.550 ;
        RECT 342.750 179.100 343.800 184.800 ;
        RECT 344.700 185.700 351.000 186.600 ;
        RECT 371.400 186.300 372.600 188.400 ;
        RECT 344.700 183.600 346.800 185.700 ;
        RECT 368.850 185.250 372.600 186.300 ;
        RECT 344.700 181.800 346.500 183.600 ;
        RECT 355.950 183.450 358.050 184.050 ;
        RECT 350.550 182.850 358.050 183.450 ;
        RECT 349.800 182.550 358.050 182.850 ;
        RECT 349.800 181.050 351.600 182.550 ;
        RECT 355.950 181.950 358.050 182.550 ;
        RECT 365.100 181.050 366.900 182.850 ;
        RECT 368.850 181.050 370.050 185.250 ;
        RECT 371.100 181.050 372.900 182.850 ;
        RECT 389.400 181.050 390.600 191.400 ;
        RECT 406.800 188.400 408.600 194.400 ;
        RECT 407.400 186.300 408.600 188.400 ;
        RECT 409.800 189.300 411.600 194.400 ;
        RECT 415.800 189.300 417.600 194.400 ;
        RECT 434.400 191.400 436.200 194.400 ;
        RECT 455.400 191.400 457.200 194.400 ;
        RECT 472.800 191.400 474.600 194.400 ;
        RECT 409.800 187.950 417.600 189.300 ;
        RECT 407.400 185.250 411.150 186.300 ;
        RECT 407.100 181.050 408.900 182.850 ;
        RECT 409.950 181.050 411.150 185.250 ;
        RECT 413.100 181.050 414.900 182.850 ;
        RECT 434.700 181.050 435.600 191.400 ;
        RECT 455.400 181.050 456.600 191.400 ;
        RECT 473.400 181.050 474.600 191.400 ;
        RECT 479.550 188.400 481.350 194.400 ;
        RECT 487.650 191.400 489.450 194.400 ;
        RECT 495.450 191.400 497.250 194.400 ;
        RECT 503.250 192.300 505.050 194.400 ;
        RECT 503.250 191.400 507.000 192.300 ;
        RECT 487.650 190.500 488.700 191.400 ;
        RECT 484.950 189.300 488.700 190.500 ;
        RECT 496.200 190.500 497.250 191.400 ;
        RECT 505.950 190.500 507.000 191.400 ;
        RECT 496.200 189.450 501.150 190.500 ;
        RECT 484.950 188.400 487.050 189.300 ;
        RECT 499.350 188.700 501.150 189.450 ;
        RECT 479.550 181.050 480.750 188.400 ;
        RECT 502.650 187.800 504.450 189.600 ;
        RECT 505.950 188.400 508.050 190.500 ;
        RECT 511.050 188.400 512.850 194.400 ;
        RECT 527.400 191.400 529.200 194.400 ;
        RECT 492.150 186.000 493.950 186.600 ;
        RECT 503.100 186.000 504.150 187.800 ;
        RECT 492.150 184.800 504.150 186.000 ;
        RECT 349.500 180.300 351.600 181.050 ;
        RECT 240.750 173.100 251.850 173.700 ;
        RECT 218.550 159.600 220.350 171.600 ;
        RECT 223.950 171.300 226.050 172.200 ;
        RECT 226.950 171.300 232.050 172.200 ;
        RECT 234.150 172.500 251.850 173.100 ;
        RECT 234.150 172.200 242.550 172.500 ;
        RECT 226.950 170.400 227.850 171.300 ;
        RECT 225.150 168.600 227.850 170.400 ;
        RECT 228.750 170.100 230.550 170.400 ;
        RECT 234.150 170.100 235.050 172.200 ;
        RECT 250.950 171.600 251.850 172.500 ;
        RECT 228.750 169.200 235.050 170.100 ;
        RECT 235.950 170.700 237.750 171.300 ;
        RECT 235.950 169.500 243.450 170.700 ;
        RECT 228.750 168.600 230.550 169.200 ;
        RECT 242.250 168.600 243.450 169.500 ;
        RECT 223.950 165.600 227.850 167.700 ;
        RECT 232.950 167.550 234.750 168.300 ;
        RECT 237.750 167.550 239.550 168.300 ;
        RECT 232.950 166.500 239.550 167.550 ;
        RECT 242.250 166.500 247.050 168.600 ;
        RECT 226.050 159.600 227.850 165.600 ;
        RECT 233.850 159.600 235.650 166.500 ;
        RECT 242.250 165.600 243.450 166.500 ;
        RECT 241.650 159.600 243.450 165.600 ;
        RECT 250.050 159.600 251.850 171.600 ;
        RECT 269.850 165.600 271.050 178.950 ;
        RECT 275.100 177.150 276.900 178.950 ;
        RECT 274.950 174.450 277.050 175.050 ;
        RECT 283.950 174.450 286.050 175.050 ;
        RECT 274.950 173.550 286.050 174.450 ;
        RECT 274.950 172.950 277.050 173.550 ;
        RECT 283.950 172.950 286.050 173.550 ;
        RECT 290.400 171.600 291.300 178.950 ;
        RECT 296.100 177.150 297.900 178.950 ;
        RECT 314.100 177.150 315.900 178.950 ;
        RECT 292.950 174.450 295.050 175.050 ;
        RECT 307.950 174.450 310.050 175.050 ;
        RECT 292.950 173.550 310.050 174.450 ;
        RECT 292.950 172.950 295.050 173.550 ;
        RECT 307.950 172.950 310.050 173.550 ;
        RECT 317.400 171.600 318.300 178.950 ;
        RECT 320.100 177.150 321.900 178.950 ;
        RECT 335.100 177.150 336.900 178.950 ;
        RECT 341.400 178.200 343.800 179.100 ;
        RECT 344.700 179.100 351.600 180.300 ;
        RECT 344.700 178.500 346.500 179.100 ;
        RECT 349.500 178.950 351.600 179.100 ;
        RECT 361.950 178.950 364.050 181.050 ;
        RECT 364.950 178.950 367.050 181.050 ;
        RECT 367.950 178.950 370.050 181.050 ;
        RECT 370.950 178.950 373.050 181.050 ;
        RECT 388.950 178.950 391.050 181.050 ;
        RECT 391.950 178.950 394.050 181.050 ;
        RECT 406.950 178.950 409.050 181.050 ;
        RECT 409.950 178.950 412.050 181.050 ;
        RECT 412.950 178.950 415.050 181.050 ;
        RECT 415.950 178.950 418.050 181.050 ;
        RECT 430.950 178.950 433.050 181.050 ;
        RECT 433.950 178.950 436.050 181.050 ;
        RECT 436.950 178.950 439.050 181.050 ;
        RECT 451.950 178.950 454.050 181.050 ;
        RECT 454.950 178.950 457.050 181.050 ;
        RECT 472.950 178.950 475.050 181.050 ;
        RECT 475.950 178.950 478.050 181.050 ;
        RECT 479.550 179.250 485.850 181.050 ;
        RECT 479.550 178.950 484.050 179.250 ;
        RECT 340.800 176.100 342.900 178.200 ;
        RECT 342.000 174.000 342.900 176.100 ;
        RECT 343.800 175.500 347.700 177.300 ;
        RECT 362.100 177.150 363.900 178.950 ;
        RECT 343.800 175.200 345.900 175.500 ;
        RECT 342.000 173.100 343.500 174.000 ;
        RECT 337.500 171.600 339.600 172.500 ;
        RECT 269.400 159.600 271.200 165.600 ;
        RECT 289.800 159.600 291.600 171.600 ;
        RECT 292.800 170.700 300.600 171.600 ;
        RECT 292.800 159.600 294.600 170.700 ;
        RECT 298.800 159.600 300.600 170.700 ;
        RECT 314.700 170.400 318.300 171.600 ;
        RECT 334.800 170.400 339.600 171.600 ;
        RECT 342.300 171.600 343.500 173.100 ;
        RECT 347.100 171.600 349.200 173.700 ;
        RECT 314.700 159.600 316.500 170.400 ;
        RECT 334.800 159.600 336.600 170.400 ;
        RECT 342.300 163.050 344.100 171.600 ;
        RECT 347.100 170.700 351.600 171.600 ;
        RECT 340.950 160.950 344.100 163.050 ;
        RECT 342.300 159.600 344.100 160.950 ;
        RECT 349.800 159.600 351.600 170.700 ;
        RECT 367.950 165.600 369.150 178.950 ;
        RECT 389.400 165.600 390.600 178.950 ;
        RECT 392.100 177.150 393.900 178.950 ;
        RECT 410.850 165.600 412.050 178.950 ;
        RECT 416.100 177.150 417.900 178.950 ;
        RECT 431.100 177.150 432.900 178.950 ;
        RECT 434.700 171.600 435.600 178.950 ;
        RECT 437.100 177.150 438.900 178.950 ;
        RECT 452.100 177.150 453.900 178.950 ;
        RECT 434.700 170.400 438.300 171.600 ;
        RECT 367.800 159.600 369.600 165.600 ;
        RECT 388.800 159.600 390.600 165.600 ;
        RECT 410.400 159.600 412.200 165.600 ;
        RECT 436.500 159.600 438.300 170.400 ;
        RECT 455.400 165.600 456.600 178.950 ;
        RECT 473.400 165.600 474.600 178.950 ;
        RECT 476.100 177.150 477.900 178.950 ;
        RECT 455.400 159.600 457.200 165.600 ;
        RECT 472.800 159.600 474.600 165.600 ;
        RECT 479.550 171.600 480.750 178.950 ;
        RECT 481.950 173.400 483.750 175.200 ;
        RECT 482.850 172.200 487.050 173.400 ;
        RECT 492.150 172.200 493.050 184.800 ;
        RECT 503.100 183.600 510.000 184.800 ;
        RECT 503.100 183.000 504.900 183.600 ;
        RECT 509.100 182.850 510.000 183.600 ;
        RECT 506.100 181.800 507.900 182.400 ;
        RECT 499.950 180.600 507.900 181.800 ;
        RECT 509.100 181.050 510.900 182.850 ;
        RECT 499.950 178.950 502.050 180.600 ;
        RECT 508.950 178.950 511.050 181.050 ;
        RECT 501.750 173.700 503.550 174.000 ;
        RECT 511.950 173.700 512.850 188.400 ;
        RECT 527.700 181.050 528.600 191.400 ;
        RECT 550.800 187.200 552.600 194.400 ;
        RECT 548.400 186.300 552.600 187.200 ;
        RECT 558.150 188.400 559.950 194.400 ;
        RECT 565.950 192.300 567.750 194.400 ;
        RECT 564.000 191.400 567.750 192.300 ;
        RECT 573.750 191.400 575.550 194.400 ;
        RECT 581.550 191.400 583.350 194.400 ;
        RECT 564.000 190.500 565.050 191.400 ;
        RECT 573.750 190.500 574.800 191.400 ;
        RECT 562.950 188.400 565.050 190.500 ;
        RECT 545.100 181.050 546.900 182.850 ;
        RECT 548.400 181.050 549.600 186.300 ;
        RECT 551.100 181.050 552.900 182.850 ;
        RECT 523.950 178.950 526.050 181.050 ;
        RECT 526.950 178.950 529.050 181.050 ;
        RECT 529.950 178.950 532.050 181.050 ;
        RECT 544.950 178.950 547.050 181.050 ;
        RECT 547.950 178.950 550.050 181.050 ;
        RECT 550.950 178.950 553.050 181.050 ;
        RECT 524.100 177.150 525.900 178.950 ;
        RECT 501.750 173.100 512.850 173.700 ;
        RECT 479.550 159.600 481.350 171.600 ;
        RECT 484.950 171.300 487.050 172.200 ;
        RECT 487.950 171.300 493.050 172.200 ;
        RECT 495.150 172.500 512.850 173.100 ;
        RECT 495.150 172.200 503.550 172.500 ;
        RECT 487.950 170.400 488.850 171.300 ;
        RECT 486.150 168.600 488.850 170.400 ;
        RECT 489.750 170.100 491.550 170.400 ;
        RECT 495.150 170.100 496.050 172.200 ;
        RECT 511.950 171.600 512.850 172.500 ;
        RECT 489.750 169.200 496.050 170.100 ;
        RECT 496.950 170.700 498.750 171.300 ;
        RECT 496.950 169.500 504.450 170.700 ;
        RECT 489.750 168.600 491.550 169.200 ;
        RECT 503.250 168.600 504.450 169.500 ;
        RECT 484.950 165.600 488.850 167.700 ;
        RECT 493.950 167.550 495.750 168.300 ;
        RECT 498.750 167.550 500.550 168.300 ;
        RECT 493.950 166.500 500.550 167.550 ;
        RECT 503.250 166.500 508.050 168.600 ;
        RECT 487.050 159.600 488.850 165.600 ;
        RECT 494.850 159.600 496.650 166.500 ;
        RECT 503.250 165.600 504.450 166.500 ;
        RECT 502.650 159.600 504.450 165.600 ;
        RECT 511.050 159.600 512.850 171.600 ;
        RECT 527.700 171.600 528.600 178.950 ;
        RECT 530.100 177.150 531.900 178.950 ;
        RECT 527.700 170.400 531.300 171.600 ;
        RECT 529.500 159.600 531.300 170.400 ;
        RECT 548.400 165.600 549.600 178.950 ;
        RECT 558.150 173.700 559.050 188.400 ;
        RECT 566.550 187.800 568.350 189.600 ;
        RECT 569.850 189.450 574.800 190.500 ;
        RECT 582.300 190.500 583.350 191.400 ;
        RECT 569.850 188.700 571.650 189.450 ;
        RECT 582.300 189.300 586.050 190.500 ;
        RECT 583.950 188.400 586.050 189.300 ;
        RECT 589.650 188.400 591.450 194.400 ;
        RECT 604.800 188.400 606.600 194.400 ;
        RECT 566.850 186.000 567.900 187.800 ;
        RECT 577.050 186.000 578.850 186.600 ;
        RECT 566.850 184.800 578.850 186.000 ;
        RECT 561.000 183.600 567.900 184.800 ;
        RECT 561.000 182.850 561.900 183.600 ;
        RECT 566.100 183.000 567.900 183.600 ;
        RECT 560.100 181.050 561.900 182.850 ;
        RECT 563.100 181.800 564.900 182.400 ;
        RECT 559.950 178.950 562.050 181.050 ;
        RECT 563.100 180.600 571.050 181.800 ;
        RECT 568.950 178.950 571.050 180.600 ;
        RECT 567.450 173.700 569.250 174.000 ;
        RECT 558.150 173.100 569.250 173.700 ;
        RECT 558.150 172.500 575.850 173.100 ;
        RECT 558.150 171.600 559.050 172.500 ;
        RECT 567.450 172.200 575.850 172.500 ;
        RECT 548.400 159.600 550.200 165.600 ;
        RECT 558.150 159.600 559.950 171.600 ;
        RECT 572.250 170.700 574.050 171.300 ;
        RECT 566.550 169.500 574.050 170.700 ;
        RECT 574.950 170.100 575.850 172.200 ;
        RECT 577.950 172.200 578.850 184.800 ;
        RECT 590.250 181.050 591.450 188.400 ;
        RECT 605.400 186.300 606.600 188.400 ;
        RECT 607.800 189.300 609.600 194.400 ;
        RECT 613.800 189.300 615.600 194.400 ;
        RECT 607.800 187.950 615.600 189.300 ;
        RECT 631.800 187.200 633.600 194.400 ;
        RECT 649.800 188.400 651.600 194.400 ;
        RECT 629.400 186.300 633.600 187.200 ;
        RECT 650.400 186.300 651.600 188.400 ;
        RECT 652.800 189.300 654.600 194.400 ;
        RECT 658.800 189.300 660.600 194.400 ;
        RECT 652.800 187.950 660.600 189.300 ;
        RECT 679.200 188.400 681.000 194.400 ;
        RECT 704.400 191.400 706.200 194.400 ;
        RECT 725.400 191.400 727.200 194.400 ;
        RECT 605.400 185.250 609.150 186.300 ;
        RECT 605.100 181.050 606.900 182.850 ;
        RECT 607.950 181.050 609.150 185.250 ;
        RECT 611.100 181.050 612.900 182.850 ;
        RECT 626.100 181.050 627.900 182.850 ;
        RECT 629.400 181.050 630.600 186.300 ;
        RECT 650.400 185.250 654.150 186.300 ;
        RECT 632.100 181.050 633.900 182.850 ;
        RECT 650.100 181.050 651.900 182.850 ;
        RECT 652.950 181.050 654.150 185.250 ;
        RECT 656.100 181.050 657.900 182.850 ;
        RECT 674.100 181.050 675.900 182.850 ;
        RECT 679.950 181.050 681.000 188.400 ;
        RECT 686.100 181.050 687.900 182.850 ;
        RECT 704.700 181.050 705.600 191.400 ;
        RECT 725.400 181.050 726.600 191.400 ;
        RECT 740.400 189.300 742.200 194.400 ;
        RECT 746.400 189.300 748.200 194.400 ;
        RECT 740.400 187.950 748.200 189.300 ;
        RECT 749.400 188.400 751.200 194.400 ;
        RECT 767.400 191.400 769.200 194.400 ;
        RECT 749.400 186.300 750.600 188.400 ;
        RECT 746.850 185.250 750.600 186.300 ;
        RECT 743.100 181.050 744.900 182.850 ;
        RECT 746.850 181.050 748.050 185.250 ;
        RECT 749.100 181.050 750.900 182.850 ;
        RECT 767.400 181.050 768.600 191.400 ;
        RECT 787.500 189.600 789.300 194.400 ;
        RECT 811.800 191.400 813.600 194.400 ;
        RECT 787.500 188.400 792.600 189.600 ;
        RECT 784.950 186.450 787.050 187.050 ;
        RECT 779.550 185.550 787.050 186.450 ;
        RECT 769.950 183.450 774.000 184.050 ;
        RECT 779.550 183.450 780.450 185.550 ;
        RECT 784.950 184.950 787.050 185.550 ;
        RECT 769.950 181.950 774.450 183.450 ;
        RECT 585.150 179.250 591.450 181.050 ;
        RECT 586.950 178.950 591.450 179.250 ;
        RECT 604.950 178.950 607.050 181.050 ;
        RECT 607.950 178.950 610.050 181.050 ;
        RECT 610.950 178.950 613.050 181.050 ;
        RECT 613.950 178.950 616.050 181.050 ;
        RECT 625.950 178.950 628.050 181.050 ;
        RECT 628.950 178.950 631.050 181.050 ;
        RECT 631.950 178.950 634.050 181.050 ;
        RECT 649.950 178.950 652.050 181.050 ;
        RECT 652.950 178.950 655.050 181.050 ;
        RECT 655.950 178.950 658.050 181.050 ;
        RECT 658.950 178.950 661.050 181.050 ;
        RECT 673.950 178.950 676.050 181.050 ;
        RECT 676.950 178.950 679.050 181.050 ;
        RECT 679.950 178.950 682.050 181.050 ;
        RECT 682.950 178.950 685.050 181.050 ;
        RECT 685.950 178.950 688.050 181.050 ;
        RECT 700.950 178.950 703.050 181.050 ;
        RECT 703.950 178.950 706.050 181.050 ;
        RECT 706.950 178.950 709.050 181.050 ;
        RECT 721.950 178.950 724.050 181.050 ;
        RECT 724.950 178.950 727.050 181.050 ;
        RECT 739.950 178.950 742.050 181.050 ;
        RECT 742.950 178.950 745.050 181.050 ;
        RECT 745.950 178.950 748.050 181.050 ;
        RECT 748.950 178.950 751.050 181.050 ;
        RECT 763.950 178.950 766.050 181.050 ;
        RECT 766.950 178.950 769.050 181.050 ;
        RECT 587.250 173.400 589.050 175.200 ;
        RECT 583.950 172.200 588.150 173.400 ;
        RECT 577.950 171.300 583.050 172.200 ;
        RECT 583.950 171.300 586.050 172.200 ;
        RECT 590.250 171.600 591.450 178.950 ;
        RECT 582.150 170.400 583.050 171.300 ;
        RECT 579.450 170.100 581.250 170.400 ;
        RECT 566.550 168.600 567.750 169.500 ;
        RECT 574.950 169.200 581.250 170.100 ;
        RECT 579.450 168.600 581.250 169.200 ;
        RECT 582.150 168.600 584.850 170.400 ;
        RECT 562.950 166.500 567.750 168.600 ;
        RECT 570.450 167.550 572.250 168.300 ;
        RECT 575.250 167.550 577.050 168.300 ;
        RECT 570.450 166.500 577.050 167.550 ;
        RECT 566.550 165.600 567.750 166.500 ;
        RECT 566.550 159.600 568.350 165.600 ;
        RECT 574.350 159.600 576.150 166.500 ;
        RECT 582.150 165.600 586.050 167.700 ;
        RECT 582.150 159.600 583.950 165.600 ;
        RECT 589.650 159.600 591.450 171.600 ;
        RECT 608.850 165.600 610.050 178.950 ;
        RECT 614.100 177.150 615.900 178.950 ;
        RECT 629.400 165.600 630.600 178.950 ;
        RECT 643.950 174.450 646.050 175.050 ;
        RECT 649.950 174.450 652.050 175.050 ;
        RECT 643.950 173.550 652.050 174.450 ;
        RECT 643.950 172.950 646.050 173.550 ;
        RECT 649.950 172.950 652.050 173.550 ;
        RECT 653.850 165.600 655.050 178.950 ;
        RECT 659.100 177.150 660.900 178.950 ;
        RECT 677.100 177.150 678.900 178.950 ;
        RECT 680.100 173.400 681.000 178.950 ;
        RECT 683.100 177.150 684.900 178.950 ;
        RECT 701.100 177.150 702.900 178.950 ;
        RECT 680.100 172.500 685.200 173.400 ;
        RECT 674.400 170.400 682.200 171.300 ;
        RECT 608.400 159.600 610.200 165.600 ;
        RECT 629.400 159.600 631.200 165.600 ;
        RECT 653.400 159.600 655.200 165.600 ;
        RECT 674.400 159.600 676.200 170.400 ;
        RECT 680.400 160.500 682.200 170.400 ;
        RECT 683.400 161.400 685.200 172.500 ;
        RECT 704.700 171.600 705.600 178.950 ;
        RECT 707.100 177.150 708.900 178.950 ;
        RECT 722.100 177.150 723.900 178.950 ;
        RECT 686.400 160.500 688.200 171.600 ;
        RECT 704.700 170.400 708.300 171.600 ;
        RECT 680.400 159.600 688.200 160.500 ;
        RECT 706.500 159.600 708.300 170.400 ;
        RECT 725.400 165.600 726.600 178.950 ;
        RECT 740.100 177.150 741.900 178.950 ;
        RECT 745.950 165.600 747.150 178.950 ;
        RECT 764.100 177.150 765.900 178.950 ;
        RECT 767.400 165.600 768.600 178.950 ;
        RECT 773.550 178.050 774.450 181.950 ;
        RECT 769.950 176.550 774.450 178.050 ;
        RECT 776.550 182.550 780.450 183.450 ;
        RECT 776.550 178.050 777.450 182.550 ;
        RECT 782.100 181.050 783.900 182.850 ;
        RECT 788.100 181.050 789.900 182.850 ;
        RECT 791.700 181.050 792.600 188.400 ;
        RECT 799.950 186.450 802.050 187.050 ;
        RECT 805.950 186.450 808.050 187.050 ;
        RECT 799.950 185.550 808.050 186.450 ;
        RECT 799.950 184.950 802.050 185.550 ;
        RECT 805.950 184.950 808.050 185.550 ;
        RECT 793.950 183.450 798.000 184.050 ;
        RECT 793.950 181.950 798.450 183.450 ;
        RECT 781.950 178.950 784.050 181.050 ;
        RECT 784.950 178.950 787.050 181.050 ;
        RECT 787.950 178.950 790.050 181.050 ;
        RECT 790.950 178.950 793.050 181.050 ;
        RECT 776.550 176.550 781.050 178.050 ;
        RECT 785.100 177.150 786.900 178.950 ;
        RECT 769.950 175.950 774.000 176.550 ;
        RECT 777.000 175.950 781.050 176.550 ;
        RECT 775.950 174.450 778.050 175.050 ;
        RECT 781.950 174.450 784.050 174.750 ;
        RECT 775.950 173.550 784.050 174.450 ;
        RECT 775.950 172.950 778.050 173.550 ;
        RECT 781.950 172.650 784.050 173.550 ;
        RECT 791.700 171.600 792.600 178.950 ;
        RECT 797.550 178.050 798.450 181.950 ;
        RECT 812.400 181.050 813.300 191.400 ;
        RECT 832.800 187.200 834.600 194.400 ;
        RECT 853.800 187.200 855.600 194.400 ;
        RECT 874.800 187.200 876.600 194.400 ;
        RECT 814.950 186.450 817.050 187.200 ;
        RECT 820.950 186.450 823.050 187.050 ;
        RECT 814.950 185.550 823.050 186.450 ;
        RECT 814.950 185.100 817.050 185.550 ;
        RECT 820.950 184.950 823.050 185.550 ;
        RECT 830.400 186.300 834.600 187.200 ;
        RECT 840.000 186.450 844.050 187.050 ;
        RECT 827.100 181.050 828.900 182.850 ;
        RECT 830.400 181.050 831.600 186.300 ;
        RECT 839.550 184.950 844.050 186.450 ;
        RECT 851.400 186.300 855.600 187.200 ;
        RECT 872.400 186.300 876.600 187.200 ;
        RECT 833.100 181.050 834.900 182.850 ;
        RECT 808.950 178.950 811.050 181.050 ;
        RECT 811.950 178.950 814.050 181.050 ;
        RECT 814.950 178.950 817.050 181.050 ;
        RECT 826.950 178.950 829.050 181.050 ;
        RECT 829.950 178.950 832.050 181.050 ;
        RECT 832.950 178.950 835.050 181.050 ;
        RECT 793.950 176.550 798.450 178.050 ;
        RECT 809.100 177.150 810.900 178.950 ;
        RECT 793.950 175.950 798.000 176.550 ;
        RECT 812.400 171.600 813.300 178.950 ;
        RECT 815.100 177.150 816.900 178.950 ;
        RECT 782.400 170.700 790.200 171.600 ;
        RECT 769.950 168.450 772.050 169.050 ;
        RECT 775.950 168.450 778.050 169.050 ;
        RECT 769.950 167.550 778.050 168.450 ;
        RECT 769.950 166.950 772.050 167.550 ;
        RECT 775.950 166.950 778.050 167.550 ;
        RECT 725.400 159.600 727.200 165.600 ;
        RECT 745.800 159.600 747.600 165.600 ;
        RECT 767.400 159.600 769.200 165.600 ;
        RECT 782.400 159.600 784.200 170.700 ;
        RECT 788.400 159.600 790.200 170.700 ;
        RECT 791.400 159.600 793.200 171.600 ;
        RECT 809.700 170.400 813.300 171.600 ;
        RECT 809.700 159.600 811.500 170.400 ;
        RECT 830.400 165.600 831.600 178.950 ;
        RECT 839.550 178.050 840.450 184.950 ;
        RECT 848.100 181.050 849.900 182.850 ;
        RECT 851.400 181.050 852.600 186.300 ;
        RECT 856.950 183.450 859.050 184.050 ;
        RECT 854.100 181.050 855.900 182.850 ;
        RECT 856.950 182.550 864.450 183.450 ;
        RECT 856.950 181.950 859.050 182.550 ;
        RECT 847.950 178.950 850.050 181.050 ;
        RECT 850.950 178.950 853.050 181.050 ;
        RECT 853.950 178.950 856.050 181.050 ;
        RECT 835.950 176.550 840.450 178.050 ;
        RECT 835.950 175.950 840.000 176.550 ;
        RECT 851.400 165.600 852.600 178.950 ;
        RECT 863.550 177.450 864.450 182.550 ;
        RECT 869.100 181.050 870.900 182.850 ;
        RECT 872.400 181.050 873.600 186.300 ;
        RECT 875.100 181.050 876.900 182.850 ;
        RECT 868.950 178.950 871.050 181.050 ;
        RECT 871.950 178.950 874.050 181.050 ;
        RECT 874.950 178.950 877.050 181.050 ;
        RECT 863.550 176.550 867.450 177.450 ;
        RECT 866.550 175.050 867.450 176.550 ;
        RECT 866.550 173.550 871.050 175.050 ;
        RECT 867.000 172.950 871.050 173.550 ;
        RECT 872.400 165.600 873.600 178.950 ;
        RECT 830.400 159.600 832.200 165.600 ;
        RECT 851.400 159.600 853.200 165.600 ;
        RECT 872.400 159.600 874.200 165.600 ;
        RECT 13.800 143.400 15.600 155.400 ;
        RECT 19.800 149.400 21.600 155.400 ;
        RECT 13.800 136.050 15.000 143.400 ;
        RECT 20.400 142.500 21.600 149.400 ;
        RECT 15.900 141.600 21.600 142.500 ;
        RECT 35.400 142.500 37.200 155.400 ;
        RECT 41.400 142.500 43.200 155.400 ;
        RECT 47.400 142.500 49.200 155.400 ;
        RECT 53.400 142.500 55.200 155.400 ;
        RECT 76.800 149.400 78.600 155.400 ;
        RECT 15.900 140.700 17.850 141.600 ;
        RECT 35.400 141.300 39.300 142.500 ;
        RECT 41.400 141.300 45.300 142.500 ;
        RECT 47.400 141.300 51.300 142.500 ;
        RECT 53.400 141.300 56.100 142.500 ;
        RECT 13.800 133.950 16.050 136.050 ;
        RECT 13.800 126.600 15.000 133.950 ;
        RECT 16.950 129.300 17.850 140.700 ;
        RECT 20.100 136.050 21.900 137.850 ;
        RECT 19.950 133.950 22.050 136.050 ;
        RECT 34.950 133.950 37.050 136.050 ;
        RECT 35.100 132.150 36.900 133.950 ;
        RECT 15.900 128.400 17.850 129.300 ;
        RECT 38.100 130.800 39.300 141.300 ;
        RECT 40.500 130.800 42.300 131.400 ;
        RECT 38.100 129.600 42.300 130.800 ;
        RECT 44.100 130.800 45.300 141.300 ;
        RECT 46.500 130.800 48.300 131.400 ;
        RECT 44.100 129.600 48.300 130.800 ;
        RECT 50.100 130.800 51.300 141.300 ;
        RECT 55.200 136.050 56.100 141.300 ;
        RECT 77.400 136.050 78.600 149.400 ;
        RECT 95.400 149.400 97.200 155.400 ;
        RECT 79.950 141.450 82.050 145.050 ;
        RECT 85.950 141.450 88.050 142.050 ;
        RECT 91.950 141.450 94.050 142.200 ;
        RECT 79.950 141.000 84.450 141.450 ;
        RECT 80.550 140.550 84.450 141.000 ;
        RECT 83.550 138.450 84.450 140.550 ;
        RECT 85.950 140.550 94.050 141.450 ;
        RECT 85.950 139.950 88.050 140.550 ;
        RECT 91.950 140.100 94.050 140.550 ;
        RECT 83.550 137.550 87.450 138.450 ;
        RECT 55.200 133.950 58.050 136.050 ;
        RECT 73.950 133.950 76.050 136.050 ;
        RECT 76.950 133.950 79.050 136.050 ;
        RECT 79.950 133.950 82.050 136.050 ;
        RECT 52.500 130.800 54.300 131.400 ;
        RECT 50.100 129.600 54.300 130.800 ;
        RECT 38.100 128.700 39.300 129.600 ;
        RECT 44.100 128.700 45.300 129.600 ;
        RECT 50.100 128.700 51.300 129.600 ;
        RECT 55.200 128.700 56.100 133.950 ;
        RECT 74.100 132.150 75.900 133.950 ;
        RECT 77.400 128.700 78.600 133.950 ;
        RECT 80.100 132.150 81.900 133.950 ;
        RECT 15.900 127.500 21.600 128.400 ;
        RECT 13.800 120.600 15.600 126.600 ;
        RECT 20.400 123.600 21.600 127.500 ;
        RECT 19.800 120.600 21.600 123.600 ;
        RECT 35.400 127.500 39.300 128.700 ;
        RECT 41.400 127.500 45.300 128.700 ;
        RECT 47.400 127.500 51.300 128.700 ;
        RECT 53.400 127.500 56.100 128.700 ;
        RECT 74.400 127.800 78.600 128.700 ;
        RECT 79.950 129.450 82.050 130.050 ;
        RECT 86.550 129.450 87.450 137.550 ;
        RECT 91.950 133.950 94.050 136.050 ;
        RECT 92.100 132.150 93.900 133.950 ;
        RECT 79.950 128.550 87.450 129.450 ;
        RECT 95.400 129.300 96.300 149.400 ;
        RECT 101.400 143.400 103.200 155.400 ;
        RECT 125.400 149.400 127.200 155.400 ;
        RECT 148.800 149.400 150.600 155.400 ;
        RECT 98.100 136.050 99.900 137.850 ;
        RECT 101.700 136.050 102.600 143.400 ;
        RECT 103.950 141.450 106.050 142.050 ;
        RECT 121.950 141.450 124.050 142.050 ;
        RECT 103.950 140.550 124.050 141.450 ;
        RECT 103.950 139.950 106.050 140.550 ;
        RECT 121.950 139.950 124.050 140.550 ;
        RECT 125.850 136.050 127.050 149.400 ;
        RECT 131.100 136.050 132.900 137.850 ;
        RECT 143.100 136.050 144.900 137.850 ;
        RECT 148.950 136.050 150.150 149.400 ;
        RECT 169.800 143.400 171.600 155.400 ;
        RECT 175.800 149.400 177.600 155.400 ;
        RECT 190.800 149.400 192.600 155.400 ;
        RECT 169.800 136.050 171.000 143.400 ;
        RECT 176.400 142.500 177.600 149.400 ;
        RECT 171.900 141.600 177.600 142.500 ;
        RECT 171.900 140.700 173.850 141.600 ;
        RECT 97.950 133.950 100.050 136.050 ;
        RECT 100.950 133.950 103.050 136.050 ;
        RECT 121.950 133.950 124.050 136.050 ;
        RECT 124.950 133.950 127.050 136.050 ;
        RECT 127.950 133.950 130.050 136.050 ;
        RECT 130.950 133.950 133.050 136.050 ;
        RECT 142.950 133.950 145.050 136.050 ;
        RECT 145.950 133.950 148.050 136.050 ;
        RECT 148.950 133.950 151.050 136.050 ;
        RECT 151.950 133.950 154.050 136.050 ;
        RECT 169.800 133.950 172.050 136.050 ;
        RECT 79.950 127.950 82.050 128.550 ;
        RECT 92.400 128.400 99.900 129.300 ;
        RECT 35.400 120.600 37.200 127.500 ;
        RECT 41.400 120.600 43.200 127.500 ;
        RECT 47.400 120.600 49.200 127.500 ;
        RECT 53.400 120.600 55.200 127.500 ;
        RECT 74.400 120.600 76.200 127.800 ;
        RECT 92.400 120.600 94.200 128.400 ;
        RECT 98.100 127.500 99.900 128.400 ;
        RECT 101.700 126.600 102.600 133.950 ;
        RECT 122.100 132.150 123.900 133.950 ;
        RECT 124.950 129.750 126.150 133.950 ;
        RECT 128.100 132.150 129.900 133.950 ;
        RECT 146.100 132.150 147.900 133.950 ;
        RECT 122.400 128.700 126.150 129.750 ;
        RECT 149.850 129.750 151.050 133.950 ;
        RECT 152.100 132.150 153.900 133.950 ;
        RECT 149.850 128.700 153.600 129.750 ;
        RECT 122.400 126.600 123.600 128.700 ;
        RECT 99.900 124.800 102.600 126.600 ;
        RECT 99.900 120.600 101.700 124.800 ;
        RECT 121.800 120.600 123.600 126.600 ;
        RECT 124.800 125.700 132.600 127.050 ;
        RECT 124.800 120.600 126.600 125.700 ;
        RECT 130.800 120.600 132.600 125.700 ;
        RECT 143.400 125.700 151.200 127.050 ;
        RECT 143.400 120.600 145.200 125.700 ;
        RECT 149.400 120.600 151.200 125.700 ;
        RECT 152.400 126.600 153.600 128.700 ;
        RECT 169.800 126.600 171.000 133.950 ;
        RECT 172.950 129.300 173.850 140.700 ;
        RECT 176.100 136.050 177.900 137.850 ;
        RECT 191.400 136.050 192.600 149.400 ;
        RECT 197.550 143.400 199.350 155.400 ;
        RECT 205.050 149.400 206.850 155.400 ;
        RECT 202.950 147.300 206.850 149.400 ;
        RECT 212.850 148.500 214.650 155.400 ;
        RECT 220.650 149.400 222.450 155.400 ;
        RECT 221.250 148.500 222.450 149.400 ;
        RECT 211.950 147.450 218.550 148.500 ;
        RECT 211.950 146.700 213.750 147.450 ;
        RECT 216.750 146.700 218.550 147.450 ;
        RECT 221.250 146.400 226.050 148.500 ;
        RECT 204.150 144.600 206.850 146.400 ;
        RECT 207.750 145.800 209.550 146.400 ;
        RECT 207.750 144.900 214.050 145.800 ;
        RECT 221.250 145.500 222.450 146.400 ;
        RECT 207.750 144.600 209.550 144.900 ;
        RECT 205.950 143.700 206.850 144.600 ;
        RECT 194.100 136.050 195.900 137.850 ;
        RECT 197.550 136.050 198.750 143.400 ;
        RECT 202.950 142.800 205.050 143.700 ;
        RECT 205.950 142.800 211.050 143.700 ;
        RECT 200.850 141.600 205.050 142.800 ;
        RECT 199.950 139.800 201.750 141.600 ;
        RECT 175.950 133.950 178.050 136.050 ;
        RECT 190.950 133.950 193.050 136.050 ;
        RECT 193.950 133.950 196.050 136.050 ;
        RECT 197.550 135.750 202.050 136.050 ;
        RECT 197.550 133.950 203.850 135.750 ;
        RECT 171.900 128.400 173.850 129.300 ;
        RECT 171.900 127.500 177.600 128.400 ;
        RECT 152.400 120.600 154.200 126.600 ;
        RECT 169.800 120.600 171.600 126.600 ;
        RECT 176.400 123.600 177.600 127.500 ;
        RECT 191.400 123.600 192.600 133.950 ;
        RECT 175.800 120.600 177.600 123.600 ;
        RECT 190.800 120.600 192.600 123.600 ;
        RECT 197.550 126.600 198.750 133.950 ;
        RECT 210.150 130.200 211.050 142.800 ;
        RECT 213.150 142.800 214.050 144.900 ;
        RECT 214.950 144.300 222.450 145.500 ;
        RECT 214.950 143.700 216.750 144.300 ;
        RECT 229.050 143.400 230.850 155.400 ;
        RECT 247.800 149.400 249.600 155.400 ;
        RECT 271.800 149.400 273.600 155.400 ;
        RECT 293.400 149.400 295.200 155.400 ;
        RECT 213.150 142.500 221.550 142.800 ;
        RECT 229.950 142.500 230.850 143.400 ;
        RECT 213.150 141.900 230.850 142.500 ;
        RECT 219.750 141.300 230.850 141.900 ;
        RECT 219.750 141.000 221.550 141.300 ;
        RECT 217.950 134.400 220.050 136.050 ;
        RECT 217.950 133.200 225.900 134.400 ;
        RECT 226.950 133.950 229.050 136.050 ;
        RECT 224.100 132.600 225.900 133.200 ;
        RECT 227.100 132.150 228.900 133.950 ;
        RECT 221.100 131.400 222.900 132.000 ;
        RECT 227.100 131.400 228.000 132.150 ;
        RECT 221.100 130.200 228.000 131.400 ;
        RECT 210.150 129.000 222.150 130.200 ;
        RECT 210.150 128.400 211.950 129.000 ;
        RECT 221.100 127.200 222.150 129.000 ;
        RECT 197.550 120.600 199.350 126.600 ;
        RECT 202.950 125.700 205.050 126.600 ;
        RECT 202.950 124.500 206.700 125.700 ;
        RECT 217.350 125.550 219.150 126.300 ;
        RECT 205.650 123.600 206.700 124.500 ;
        RECT 214.200 124.500 219.150 125.550 ;
        RECT 220.650 125.400 222.450 127.200 ;
        RECT 229.950 126.600 230.850 141.300 ;
        RECT 242.100 136.050 243.900 137.850 ;
        RECT 247.950 136.050 249.150 149.400 ;
        RECT 272.400 136.050 273.600 149.400 ;
        RECT 274.950 141.450 277.050 142.050 ;
        RECT 280.950 141.450 283.050 142.050 ;
        RECT 274.950 140.550 283.050 141.450 ;
        RECT 274.950 139.950 277.050 140.550 ;
        RECT 280.950 139.950 283.050 140.550 ;
        RECT 293.850 136.050 295.050 149.400 ;
        RECT 302.550 143.400 304.350 155.400 ;
        RECT 310.050 149.400 311.850 155.400 ;
        RECT 307.950 147.300 311.850 149.400 ;
        RECT 317.850 148.500 319.650 155.400 ;
        RECT 325.650 149.400 327.450 155.400 ;
        RECT 326.250 148.500 327.450 149.400 ;
        RECT 316.950 147.450 323.550 148.500 ;
        RECT 316.950 146.700 318.750 147.450 ;
        RECT 321.750 146.700 323.550 147.450 ;
        RECT 326.250 146.400 331.050 148.500 ;
        RECT 309.150 144.600 311.850 146.400 ;
        RECT 312.750 145.800 314.550 146.400 ;
        RECT 312.750 144.900 319.050 145.800 ;
        RECT 326.250 145.500 327.450 146.400 ;
        RECT 312.750 144.600 314.550 144.900 ;
        RECT 310.950 143.700 311.850 144.600 ;
        RECT 299.100 136.050 300.900 137.850 ;
        RECT 302.550 136.050 303.750 143.400 ;
        RECT 307.950 142.800 310.050 143.700 ;
        RECT 310.950 142.800 316.050 143.700 ;
        RECT 305.850 141.600 310.050 142.800 ;
        RECT 304.950 139.800 306.750 141.600 ;
        RECT 241.950 133.950 244.050 136.050 ;
        RECT 244.950 133.950 247.050 136.050 ;
        RECT 247.950 133.950 250.050 136.050 ;
        RECT 250.950 133.950 253.050 136.050 ;
        RECT 268.950 133.950 271.050 136.050 ;
        RECT 271.950 133.950 274.050 136.050 ;
        RECT 274.950 133.950 277.050 136.050 ;
        RECT 289.950 133.950 292.050 136.050 ;
        RECT 292.950 133.950 295.050 136.050 ;
        RECT 295.950 133.950 298.050 136.050 ;
        RECT 298.950 133.950 301.050 136.050 ;
        RECT 302.550 135.750 307.050 136.050 ;
        RECT 302.550 133.950 308.850 135.750 ;
        RECT 245.100 132.150 246.900 133.950 ;
        RECT 248.850 129.750 250.050 133.950 ;
        RECT 251.100 132.150 252.900 133.950 ;
        RECT 269.100 132.150 270.900 133.950 ;
        RECT 248.850 128.700 252.600 129.750 ;
        RECT 272.400 128.700 273.600 133.950 ;
        RECT 275.100 132.150 276.900 133.950 ;
        RECT 290.100 132.150 291.900 133.950 ;
        RECT 292.950 129.750 294.150 133.950 ;
        RECT 296.100 132.150 297.900 133.950 ;
        RECT 223.950 124.500 226.050 126.600 ;
        RECT 214.200 123.600 215.250 124.500 ;
        RECT 223.950 123.600 225.000 124.500 ;
        RECT 205.650 120.600 207.450 123.600 ;
        RECT 213.450 120.600 215.250 123.600 ;
        RECT 221.250 122.700 225.000 123.600 ;
        RECT 221.250 120.600 223.050 122.700 ;
        RECT 229.050 120.600 230.850 126.600 ;
        RECT 242.400 125.700 250.200 127.050 ;
        RECT 242.400 120.600 244.200 125.700 ;
        RECT 248.400 120.600 250.200 125.700 ;
        RECT 251.400 126.600 252.600 128.700 ;
        RECT 269.400 127.800 273.600 128.700 ;
        RECT 290.400 128.700 294.150 129.750 ;
        RECT 251.400 120.600 253.200 126.600 ;
        RECT 269.400 120.600 271.200 127.800 ;
        RECT 290.400 126.600 291.600 128.700 ;
        RECT 289.800 120.600 291.600 126.600 ;
        RECT 292.800 125.700 300.600 127.050 ;
        RECT 292.800 120.600 294.600 125.700 ;
        RECT 298.800 120.600 300.600 125.700 ;
        RECT 302.550 126.600 303.750 133.950 ;
        RECT 315.150 130.200 316.050 142.800 ;
        RECT 318.150 142.800 319.050 144.900 ;
        RECT 319.950 144.300 327.450 145.500 ;
        RECT 319.950 143.700 321.750 144.300 ;
        RECT 334.050 143.400 335.850 155.400 ;
        RECT 318.150 142.500 326.550 142.800 ;
        RECT 334.950 142.500 335.850 143.400 ;
        RECT 318.150 141.900 335.850 142.500 ;
        RECT 324.750 141.300 335.850 141.900 ;
        RECT 324.750 141.000 326.550 141.300 ;
        RECT 322.950 134.400 325.050 136.050 ;
        RECT 322.950 133.200 330.900 134.400 ;
        RECT 331.950 133.950 334.050 136.050 ;
        RECT 329.100 132.600 330.900 133.200 ;
        RECT 332.100 132.150 333.900 133.950 ;
        RECT 326.100 131.400 327.900 132.000 ;
        RECT 332.100 131.400 333.000 132.150 ;
        RECT 326.100 130.200 333.000 131.400 ;
        RECT 315.150 129.000 327.150 130.200 ;
        RECT 315.150 128.400 316.950 129.000 ;
        RECT 326.100 127.200 327.150 129.000 ;
        RECT 302.550 120.600 304.350 126.600 ;
        RECT 307.950 125.700 310.050 126.600 ;
        RECT 307.950 124.500 311.700 125.700 ;
        RECT 322.350 125.550 324.150 126.300 ;
        RECT 310.650 123.600 311.700 124.500 ;
        RECT 319.200 124.500 324.150 125.550 ;
        RECT 325.650 125.400 327.450 127.200 ;
        RECT 334.950 126.600 335.850 141.300 ;
        RECT 328.950 124.500 331.050 126.600 ;
        RECT 319.200 123.600 320.250 124.500 ;
        RECT 328.950 123.600 330.000 124.500 ;
        RECT 310.650 120.600 312.450 123.600 ;
        RECT 318.450 120.600 320.250 123.600 ;
        RECT 326.250 122.700 330.000 123.600 ;
        RECT 326.250 120.600 328.050 122.700 ;
        RECT 334.050 120.600 335.850 126.600 ;
        RECT 349.800 143.400 351.600 155.400 ;
        RECT 355.800 149.400 357.600 155.400 ;
        RECT 349.800 136.050 351.000 143.400 ;
        RECT 356.400 142.500 357.600 149.400 ;
        RECT 351.900 141.600 357.600 142.500 ;
        RECT 371.400 149.400 373.200 155.400 ;
        RECT 351.900 140.700 353.850 141.600 ;
        RECT 349.800 133.950 352.050 136.050 ;
        RECT 349.800 126.600 351.000 133.950 ;
        RECT 352.950 129.300 353.850 140.700 ;
        RECT 356.100 136.050 357.900 137.850 ;
        RECT 371.400 136.050 372.600 149.400 ;
        RECT 392.400 142.500 394.200 155.400 ;
        RECT 398.400 142.500 400.200 155.400 ;
        RECT 404.400 142.500 406.200 155.400 ;
        RECT 410.400 142.500 412.200 155.400 ;
        RECT 433.800 149.400 435.600 155.400 ;
        RECT 455.400 149.400 457.200 155.400 ;
        RECT 392.400 141.300 396.300 142.500 ;
        RECT 398.400 141.300 402.300 142.500 ;
        RECT 404.400 141.300 408.300 142.500 ;
        RECT 410.400 141.300 413.100 142.500 ;
        RECT 355.950 133.950 358.050 136.050 ;
        RECT 367.950 133.950 370.050 136.050 ;
        RECT 370.950 133.950 373.050 136.050 ;
        RECT 373.950 133.950 376.050 136.050 ;
        RECT 391.950 133.950 394.050 136.050 ;
        RECT 368.100 132.150 369.900 133.950 ;
        RECT 351.900 128.400 353.850 129.300 ;
        RECT 371.400 128.700 372.600 133.950 ;
        RECT 374.100 132.150 375.900 133.950 ;
        RECT 392.100 132.150 393.900 133.950 ;
        RECT 395.100 130.800 396.300 141.300 ;
        RECT 397.500 130.800 399.300 131.400 ;
        RECT 395.100 129.600 399.300 130.800 ;
        RECT 401.100 130.800 402.300 141.300 ;
        RECT 403.500 130.800 405.300 131.400 ;
        RECT 401.100 129.600 405.300 130.800 ;
        RECT 407.100 130.800 408.300 141.300 ;
        RECT 412.200 136.050 413.100 141.300 ;
        RECT 434.400 136.050 435.600 149.400 ;
        RECT 455.850 136.050 457.050 149.400 ;
        RECT 464.550 143.400 466.350 155.400 ;
        RECT 472.050 149.400 473.850 155.400 ;
        RECT 469.950 147.300 473.850 149.400 ;
        RECT 479.850 148.500 481.650 155.400 ;
        RECT 487.650 149.400 489.450 155.400 ;
        RECT 488.250 148.500 489.450 149.400 ;
        RECT 478.950 147.450 485.550 148.500 ;
        RECT 478.950 146.700 480.750 147.450 ;
        RECT 483.750 146.700 485.550 147.450 ;
        RECT 488.250 146.400 493.050 148.500 ;
        RECT 471.150 144.600 473.850 146.400 ;
        RECT 474.750 145.800 476.550 146.400 ;
        RECT 474.750 144.900 481.050 145.800 ;
        RECT 488.250 145.500 489.450 146.400 ;
        RECT 474.750 144.600 476.550 144.900 ;
        RECT 472.950 143.700 473.850 144.600 ;
        RECT 461.100 136.050 462.900 137.850 ;
        RECT 464.550 136.050 465.750 143.400 ;
        RECT 469.950 142.800 472.050 143.700 ;
        RECT 472.950 142.800 478.050 143.700 ;
        RECT 467.850 141.600 472.050 142.800 ;
        RECT 466.950 139.800 468.750 141.600 ;
        RECT 412.200 133.950 415.050 136.050 ;
        RECT 430.950 133.950 433.050 136.050 ;
        RECT 433.950 133.950 436.050 136.050 ;
        RECT 436.950 133.950 439.050 136.050 ;
        RECT 451.950 133.950 454.050 136.050 ;
        RECT 454.950 133.950 457.050 136.050 ;
        RECT 457.950 133.950 460.050 136.050 ;
        RECT 460.950 133.950 463.050 136.050 ;
        RECT 464.550 135.750 469.050 136.050 ;
        RECT 464.550 133.950 470.850 135.750 ;
        RECT 409.500 130.800 411.300 131.400 ;
        RECT 407.100 129.600 411.300 130.800 ;
        RECT 395.100 128.700 396.300 129.600 ;
        RECT 401.100 128.700 402.300 129.600 ;
        RECT 407.100 128.700 408.300 129.600 ;
        RECT 412.200 128.700 413.100 133.950 ;
        RECT 431.100 132.150 432.900 133.950 ;
        RECT 434.400 128.700 435.600 133.950 ;
        RECT 437.100 132.150 438.900 133.950 ;
        RECT 452.100 132.150 453.900 133.950 ;
        RECT 454.950 129.750 456.150 133.950 ;
        RECT 458.100 132.150 459.900 133.950 ;
        RECT 351.900 127.500 357.600 128.400 ;
        RECT 371.400 127.800 375.600 128.700 ;
        RECT 349.800 120.600 351.600 126.600 ;
        RECT 356.400 123.600 357.600 127.500 ;
        RECT 355.800 120.600 357.600 123.600 ;
        RECT 373.800 120.600 375.600 127.800 ;
        RECT 392.400 127.500 396.300 128.700 ;
        RECT 398.400 127.500 402.300 128.700 ;
        RECT 404.400 127.500 408.300 128.700 ;
        RECT 410.400 127.500 413.100 128.700 ;
        RECT 431.400 127.800 435.600 128.700 ;
        RECT 452.400 128.700 456.150 129.750 ;
        RECT 392.400 120.600 394.200 127.500 ;
        RECT 398.400 120.600 400.200 127.500 ;
        RECT 404.400 120.600 406.200 127.500 ;
        RECT 410.400 120.600 412.200 127.500 ;
        RECT 431.400 120.600 433.200 127.800 ;
        RECT 452.400 126.600 453.600 128.700 ;
        RECT 451.800 120.600 453.600 126.600 ;
        RECT 454.800 125.700 462.600 127.050 ;
        RECT 454.800 120.600 456.600 125.700 ;
        RECT 460.800 120.600 462.600 125.700 ;
        RECT 464.550 126.600 465.750 133.950 ;
        RECT 477.150 130.200 478.050 142.800 ;
        RECT 480.150 142.800 481.050 144.900 ;
        RECT 481.950 144.300 489.450 145.500 ;
        RECT 481.950 143.700 483.750 144.300 ;
        RECT 496.050 143.400 497.850 155.400 ;
        RECT 509.400 144.600 511.200 155.400 ;
        RECT 515.400 154.500 523.200 155.400 ;
        RECT 515.400 144.600 517.200 154.500 ;
        RECT 509.400 143.700 517.200 144.600 ;
        RECT 480.150 142.500 488.550 142.800 ;
        RECT 496.950 142.500 497.850 143.400 ;
        RECT 518.400 142.500 520.200 153.600 ;
        RECT 521.400 143.400 523.200 154.500 ;
        RECT 540.300 144.900 542.100 155.400 ;
        RECT 539.700 143.400 542.100 144.900 ;
        RECT 547.800 143.400 549.600 155.400 ;
        RECT 563.400 144.300 565.200 155.400 ;
        RECT 569.400 144.300 571.200 155.400 ;
        RECT 563.400 143.400 571.200 144.300 ;
        RECT 572.400 143.400 574.200 155.400 ;
        RECT 590.400 149.400 592.200 155.400 ;
        RECT 607.800 149.400 609.600 155.400 ;
        RECT 480.150 141.900 497.850 142.500 ;
        RECT 486.750 141.300 497.850 141.900 ;
        RECT 486.750 141.000 488.550 141.300 ;
        RECT 484.950 134.400 487.050 136.050 ;
        RECT 484.950 133.200 492.900 134.400 ;
        RECT 493.950 133.950 496.050 136.050 ;
        RECT 491.100 132.600 492.900 133.200 ;
        RECT 494.100 132.150 495.900 133.950 ;
        RECT 488.100 131.400 489.900 132.000 ;
        RECT 494.100 131.400 495.000 132.150 ;
        RECT 488.100 130.200 495.000 131.400 ;
        RECT 477.150 129.000 489.150 130.200 ;
        RECT 477.150 128.400 478.950 129.000 ;
        RECT 488.100 127.200 489.150 129.000 ;
        RECT 464.550 120.600 466.350 126.600 ;
        RECT 469.950 125.700 472.050 126.600 ;
        RECT 469.950 124.500 473.700 125.700 ;
        RECT 484.350 125.550 486.150 126.300 ;
        RECT 472.650 123.600 473.700 124.500 ;
        RECT 481.200 124.500 486.150 125.550 ;
        RECT 487.650 125.400 489.450 127.200 ;
        RECT 496.950 126.600 497.850 141.300 ;
        RECT 515.100 141.600 520.200 142.500 ;
        RECT 512.100 136.050 513.900 137.850 ;
        RECT 515.100 136.050 516.000 141.600 ;
        RECT 518.100 136.050 519.900 137.850 ;
        RECT 539.700 136.050 541.050 143.400 ;
        RECT 548.400 141.900 549.600 143.400 ;
        RECT 508.950 133.950 511.050 136.050 ;
        RECT 511.950 133.950 514.050 136.050 ;
        RECT 514.950 133.950 517.050 136.050 ;
        RECT 517.950 133.950 520.050 136.050 ;
        RECT 520.950 133.950 523.050 136.050 ;
        RECT 538.950 133.950 541.050 136.050 ;
        RECT 542.400 140.700 549.600 141.900 ;
        RECT 542.400 140.100 544.200 140.700 ;
        RECT 509.100 132.150 510.900 133.950 ;
        RECT 514.950 126.600 516.000 133.950 ;
        RECT 521.100 132.150 522.900 133.950 ;
        RECT 517.950 129.450 520.050 130.050 ;
        RECT 523.950 129.450 526.050 130.050 ;
        RECT 517.950 128.550 526.050 129.450 ;
        RECT 517.950 127.950 520.050 128.550 ;
        RECT 523.950 127.950 526.050 128.550 ;
        RECT 538.950 126.600 540.000 133.950 ;
        RECT 542.400 129.600 543.300 140.100 ;
        RECT 545.100 136.050 546.900 137.850 ;
        RECT 566.100 136.050 567.900 137.850 ;
        RECT 572.700 136.050 573.600 143.400 ;
        RECT 587.100 136.050 588.900 137.850 ;
        RECT 590.400 136.050 591.600 149.400 ;
        RECT 592.950 138.450 595.050 139.050 ;
        RECT 598.950 138.450 601.050 139.050 ;
        RECT 592.950 137.550 601.050 138.450 ;
        RECT 592.950 136.950 595.050 137.550 ;
        RECT 598.950 136.950 601.050 137.550 ;
        RECT 608.400 136.050 609.600 149.400 ;
        RECT 614.550 143.400 616.350 155.400 ;
        RECT 622.050 149.400 623.850 155.400 ;
        RECT 619.950 147.300 623.850 149.400 ;
        RECT 629.850 148.500 631.650 155.400 ;
        RECT 637.650 149.400 639.450 155.400 ;
        RECT 638.250 148.500 639.450 149.400 ;
        RECT 628.950 147.450 635.550 148.500 ;
        RECT 628.950 146.700 630.750 147.450 ;
        RECT 633.750 146.700 635.550 147.450 ;
        RECT 638.250 146.400 643.050 148.500 ;
        RECT 621.150 144.600 623.850 146.400 ;
        RECT 624.750 145.800 626.550 146.400 ;
        RECT 624.750 144.900 631.050 145.800 ;
        RECT 638.250 145.500 639.450 146.400 ;
        RECT 624.750 144.600 626.550 144.900 ;
        RECT 622.950 143.700 623.850 144.600 ;
        RECT 611.100 136.050 612.900 137.850 ;
        RECT 614.550 136.050 615.750 143.400 ;
        RECT 619.950 142.800 622.050 143.700 ;
        RECT 622.950 142.800 628.050 143.700 ;
        RECT 617.850 141.600 622.050 142.800 ;
        RECT 616.950 139.800 618.750 141.600 ;
        RECT 544.950 133.950 547.050 136.050 ;
        RECT 547.950 133.950 550.050 136.050 ;
        RECT 562.950 133.950 565.050 136.050 ;
        RECT 565.950 133.950 568.050 136.050 ;
        RECT 568.950 133.950 571.050 136.050 ;
        RECT 571.950 133.950 574.050 136.050 ;
        RECT 586.950 133.950 589.050 136.050 ;
        RECT 589.950 133.950 592.050 136.050 ;
        RECT 607.950 133.950 610.050 136.050 ;
        RECT 610.950 133.950 613.050 136.050 ;
        RECT 614.550 135.750 619.050 136.050 ;
        RECT 614.550 133.950 620.850 135.750 ;
        RECT 548.100 132.150 549.900 133.950 ;
        RECT 563.100 132.150 564.900 133.950 ;
        RECT 569.100 132.150 570.900 133.950 ;
        RECT 542.400 128.700 544.200 129.600 ;
        RECT 547.950 129.450 550.050 130.050 ;
        RECT 568.950 129.450 571.050 130.050 ;
        RECT 542.400 127.800 545.700 128.700 ;
        RECT 547.950 128.550 571.050 129.450 ;
        RECT 547.950 127.950 550.050 128.550 ;
        RECT 568.950 127.950 571.050 128.550 ;
        RECT 490.950 124.500 493.050 126.600 ;
        RECT 481.200 123.600 482.250 124.500 ;
        RECT 490.950 123.600 492.000 124.500 ;
        RECT 472.650 120.600 474.450 123.600 ;
        RECT 480.450 120.600 482.250 123.600 ;
        RECT 488.250 122.700 492.000 123.600 ;
        RECT 488.250 120.600 490.050 122.700 ;
        RECT 496.050 120.600 497.850 126.600 ;
        RECT 514.200 120.600 516.000 126.600 ;
        RECT 538.800 120.600 540.600 126.600 ;
        RECT 544.800 123.600 545.700 127.800 ;
        RECT 572.700 126.600 573.600 133.950 ;
        RECT 568.500 125.400 573.600 126.600 ;
        RECT 544.800 120.600 546.600 123.600 ;
        RECT 568.500 120.600 570.300 125.400 ;
        RECT 590.400 123.600 591.600 133.950 ;
        RECT 608.400 123.600 609.600 133.950 ;
        RECT 590.400 120.600 592.200 123.600 ;
        RECT 607.800 120.600 609.600 123.600 ;
        RECT 614.550 126.600 615.750 133.950 ;
        RECT 627.150 130.200 628.050 142.800 ;
        RECT 630.150 142.800 631.050 144.900 ;
        RECT 631.950 144.300 639.450 145.500 ;
        RECT 631.950 143.700 633.750 144.300 ;
        RECT 646.050 143.400 647.850 155.400 ;
        RECT 661.800 149.400 663.600 155.400 ;
        RECT 630.150 142.500 638.550 142.800 ;
        RECT 646.950 142.500 647.850 143.400 ;
        RECT 630.150 141.900 647.850 142.500 ;
        RECT 636.750 141.300 647.850 141.900 ;
        RECT 636.750 141.000 638.550 141.300 ;
        RECT 634.950 134.400 637.050 136.050 ;
        RECT 634.950 133.200 642.900 134.400 ;
        RECT 643.950 133.950 646.050 136.050 ;
        RECT 641.100 132.600 642.900 133.200 ;
        RECT 644.100 132.150 645.900 133.950 ;
        RECT 638.100 131.400 639.900 132.000 ;
        RECT 644.100 131.400 645.000 132.150 ;
        RECT 638.100 130.200 645.000 131.400 ;
        RECT 627.150 129.000 639.150 130.200 ;
        RECT 627.150 128.400 628.950 129.000 ;
        RECT 638.100 127.200 639.150 129.000 ;
        RECT 614.550 120.600 616.350 126.600 ;
        RECT 619.950 125.700 622.050 126.600 ;
        RECT 619.950 124.500 623.700 125.700 ;
        RECT 634.350 125.550 636.150 126.300 ;
        RECT 622.650 123.600 623.700 124.500 ;
        RECT 631.200 124.500 636.150 125.550 ;
        RECT 637.650 125.400 639.450 127.200 ;
        RECT 646.950 126.600 647.850 141.300 ;
        RECT 662.400 136.050 663.600 149.400 ;
        RECT 668.550 143.400 670.350 155.400 ;
        RECT 676.050 149.400 677.850 155.400 ;
        RECT 673.950 147.300 677.850 149.400 ;
        RECT 683.850 148.500 685.650 155.400 ;
        RECT 691.650 149.400 693.450 155.400 ;
        RECT 692.250 148.500 693.450 149.400 ;
        RECT 682.950 147.450 689.550 148.500 ;
        RECT 682.950 146.700 684.750 147.450 ;
        RECT 687.750 146.700 689.550 147.450 ;
        RECT 692.250 146.400 697.050 148.500 ;
        RECT 675.150 144.600 677.850 146.400 ;
        RECT 678.750 145.800 680.550 146.400 ;
        RECT 678.750 144.900 685.050 145.800 ;
        RECT 692.250 145.500 693.450 146.400 ;
        RECT 678.750 144.600 680.550 144.900 ;
        RECT 676.950 143.700 677.850 144.600 ;
        RECT 665.100 136.050 666.900 137.850 ;
        RECT 668.550 136.050 669.750 143.400 ;
        RECT 673.950 142.800 676.050 143.700 ;
        RECT 676.950 142.800 682.050 143.700 ;
        RECT 671.850 141.600 676.050 142.800 ;
        RECT 670.950 139.800 672.750 141.600 ;
        RECT 661.950 133.950 664.050 136.050 ;
        RECT 664.950 133.950 667.050 136.050 ;
        RECT 668.550 135.750 673.050 136.050 ;
        RECT 668.550 133.950 674.850 135.750 ;
        RECT 640.950 124.500 643.050 126.600 ;
        RECT 631.200 123.600 632.250 124.500 ;
        RECT 640.950 123.600 642.000 124.500 ;
        RECT 622.650 120.600 624.450 123.600 ;
        RECT 630.450 120.600 632.250 123.600 ;
        RECT 638.250 122.700 642.000 123.600 ;
        RECT 638.250 120.600 640.050 122.700 ;
        RECT 646.050 120.600 647.850 126.600 ;
        RECT 662.400 123.600 663.600 133.950 ;
        RECT 661.800 120.600 663.600 123.600 ;
        RECT 668.550 126.600 669.750 133.950 ;
        RECT 681.150 130.200 682.050 142.800 ;
        RECT 684.150 142.800 685.050 144.900 ;
        RECT 685.950 144.300 693.450 145.500 ;
        RECT 685.950 143.700 687.750 144.300 ;
        RECT 700.050 143.400 701.850 155.400 ;
        RECT 717.900 143.400 721.200 155.400 ;
        RECT 745.800 149.400 747.600 155.400 ;
        RECT 684.150 142.500 692.550 142.800 ;
        RECT 700.950 142.500 701.850 143.400 ;
        RECT 684.150 141.900 701.850 142.500 ;
        RECT 690.750 141.300 701.850 141.900 ;
        RECT 690.750 141.000 692.550 141.300 ;
        RECT 688.950 134.400 691.050 136.050 ;
        RECT 688.950 133.200 696.900 134.400 ;
        RECT 697.950 133.950 700.050 136.050 ;
        RECT 695.100 132.600 696.900 133.200 ;
        RECT 698.100 132.150 699.900 133.950 ;
        RECT 692.100 131.400 693.900 132.000 ;
        RECT 698.100 131.400 699.000 132.150 ;
        RECT 692.100 130.200 699.000 131.400 ;
        RECT 681.150 129.000 693.150 130.200 ;
        RECT 681.150 128.400 682.950 129.000 ;
        RECT 692.100 127.200 693.150 129.000 ;
        RECT 668.550 120.600 670.350 126.600 ;
        RECT 673.950 125.700 676.050 126.600 ;
        RECT 673.950 124.500 677.700 125.700 ;
        RECT 688.350 125.550 690.150 126.300 ;
        RECT 676.650 123.600 677.700 124.500 ;
        RECT 685.200 124.500 690.150 125.550 ;
        RECT 691.650 125.400 693.450 127.200 ;
        RECT 700.950 126.600 701.850 141.300 ;
        RECT 713.100 136.050 714.900 137.850 ;
        RECT 719.100 136.050 720.300 143.400 ;
        RECT 724.950 141.450 727.050 142.050 ;
        RECT 724.950 140.550 735.450 141.450 ;
        RECT 724.950 139.950 727.050 140.550 ;
        RECT 725.100 136.050 726.900 137.850 ;
        RECT 712.950 133.950 715.050 136.050 ;
        RECT 715.950 133.950 718.050 136.050 ;
        RECT 718.950 133.950 721.050 136.050 ;
        RECT 721.950 133.950 724.050 136.050 ;
        RECT 724.950 133.950 727.050 136.050 ;
        RECT 716.100 132.150 717.900 133.950 ;
        RECT 718.950 129.300 720.300 133.950 ;
        RECT 722.100 132.150 723.900 133.950 ;
        RECT 734.550 133.050 735.450 140.550 ;
        RECT 740.100 136.050 741.900 137.850 ;
        RECT 745.950 136.050 747.150 149.400 ;
        RECT 766.800 143.400 768.600 155.400 ;
        RECT 769.800 144.300 771.600 155.400 ;
        RECT 775.800 144.300 777.600 155.400 ;
        RECT 793.800 149.400 795.600 155.400 ;
        RECT 814.800 149.400 816.600 155.400 ;
        RECT 836.400 149.400 838.200 155.400 ;
        RECT 856.800 149.400 858.600 155.400 ;
        RECT 875.400 149.400 877.200 155.400 ;
        RECT 769.800 143.400 777.600 144.300 ;
        RECT 751.950 138.450 754.050 139.050 ;
        RECT 751.950 137.550 762.450 138.450 ;
        RECT 751.950 136.950 754.050 137.550 ;
        RECT 739.950 133.950 742.050 136.050 ;
        RECT 742.950 133.950 745.050 136.050 ;
        RECT 745.950 133.950 748.050 136.050 ;
        RECT 748.950 133.950 751.050 136.050 ;
        RECT 734.550 131.550 739.050 133.050 ;
        RECT 743.100 132.150 744.900 133.950 ;
        RECT 735.000 130.950 739.050 131.550 ;
        RECT 746.850 129.750 748.050 133.950 ;
        RECT 749.100 132.150 750.900 133.950 ;
        RECT 761.550 133.050 762.450 137.550 ;
        RECT 767.400 136.050 768.300 143.400 ;
        RECT 783.000 138.450 787.050 139.050 ;
        RECT 773.100 136.050 774.900 137.850 ;
        RECT 782.550 136.950 787.050 138.450 ;
        RECT 766.950 133.950 769.050 136.050 ;
        RECT 769.950 133.950 772.050 136.050 ;
        RECT 772.950 133.950 775.050 136.050 ;
        RECT 775.950 133.950 778.050 136.050 ;
        RECT 761.550 131.550 766.050 133.050 ;
        RECT 762.000 130.950 766.050 131.550 ;
        RECT 718.950 128.100 723.600 129.300 ;
        RECT 746.850 128.700 750.600 129.750 ;
        RECT 694.950 124.500 697.050 126.600 ;
        RECT 685.200 123.600 686.250 124.500 ;
        RECT 694.950 123.600 696.000 124.500 ;
        RECT 676.650 120.600 678.450 123.600 ;
        RECT 684.450 120.600 686.250 123.600 ;
        RECT 692.250 122.700 696.000 123.600 ;
        RECT 692.250 120.600 694.050 122.700 ;
        RECT 700.050 120.600 701.850 126.600 ;
        RECT 713.400 126.000 721.200 126.900 ;
        RECT 722.700 126.600 723.600 128.100 ;
        RECT 713.400 120.600 715.200 126.000 ;
        RECT 719.400 121.500 721.200 126.000 ;
        RECT 722.400 122.400 724.200 126.600 ;
        RECT 725.400 121.500 727.200 126.600 ;
        RECT 719.400 120.600 727.200 121.500 ;
        RECT 740.400 125.700 748.200 127.050 ;
        RECT 740.400 120.600 742.200 125.700 ;
        RECT 746.400 120.600 748.200 125.700 ;
        RECT 749.400 126.600 750.600 128.700 ;
        RECT 767.400 126.600 768.300 133.950 ;
        RECT 770.100 132.150 771.900 133.950 ;
        RECT 776.100 132.150 777.900 133.950 ;
        RECT 782.550 133.050 783.450 136.950 ;
        RECT 788.100 136.050 789.900 137.850 ;
        RECT 793.950 136.050 795.150 149.400 ;
        RECT 796.950 141.450 799.050 141.900 ;
        RECT 811.950 141.450 814.050 142.050 ;
        RECT 796.950 140.550 814.050 141.450 ;
        RECT 796.950 139.800 799.050 140.550 ;
        RECT 811.950 139.950 814.050 140.550 ;
        RECT 815.400 136.050 816.600 149.400 ;
        RECT 828.000 138.450 832.050 139.050 ;
        RECT 818.100 136.050 819.900 137.850 ;
        RECT 827.550 136.950 832.050 138.450 ;
        RECT 787.950 133.950 790.050 136.050 ;
        RECT 790.950 133.950 793.050 136.050 ;
        RECT 793.950 133.950 796.050 136.050 ;
        RECT 796.950 133.950 799.050 136.050 ;
        RECT 814.950 133.950 817.050 136.050 ;
        RECT 817.950 133.950 820.050 136.050 ;
        RECT 778.950 130.950 787.050 133.050 ;
        RECT 791.100 132.150 792.900 133.950 ;
        RECT 794.850 129.750 796.050 133.950 ;
        RECT 797.100 132.150 798.900 133.950 ;
        RECT 794.850 128.700 798.600 129.750 ;
        RECT 749.400 120.600 751.200 126.600 ;
        RECT 767.400 125.400 772.500 126.600 ;
        RECT 770.700 120.600 772.500 125.400 ;
        RECT 788.400 125.700 796.200 127.050 ;
        RECT 788.400 120.600 790.200 125.700 ;
        RECT 794.400 120.600 796.200 125.700 ;
        RECT 797.400 126.600 798.600 128.700 ;
        RECT 797.400 120.600 799.200 126.600 ;
        RECT 815.400 123.600 816.600 133.950 ;
        RECT 827.550 133.050 828.450 136.950 ;
        RECT 836.850 136.050 838.050 149.400 ;
        RECT 842.100 136.050 843.900 137.850 ;
        RECT 857.400 136.050 858.600 149.400 ;
        RECT 875.700 149.100 877.200 149.400 ;
        RECT 881.400 149.400 883.200 155.400 ;
        RECT 881.400 149.100 882.300 149.400 ;
        RECT 875.700 148.200 882.300 149.100 ;
        RECT 859.950 141.450 862.050 142.050 ;
        RECT 877.950 141.450 880.050 142.050 ;
        RECT 859.950 140.550 880.050 141.450 ;
        RECT 859.950 139.950 862.050 140.550 ;
        RECT 877.950 139.950 880.050 140.550 ;
        RECT 860.100 136.050 861.900 137.850 ;
        RECT 875.100 136.050 876.900 137.850 ;
        RECT 881.400 136.050 882.300 148.200 ;
        RECT 832.950 133.950 835.050 136.050 ;
        RECT 835.950 133.950 838.050 136.050 ;
        RECT 838.950 133.950 841.050 136.050 ;
        RECT 841.950 133.950 844.050 136.050 ;
        RECT 856.950 133.950 859.050 136.050 ;
        RECT 859.950 133.950 862.050 136.050 ;
        RECT 871.950 133.950 874.050 136.050 ;
        RECT 874.950 133.950 877.050 136.050 ;
        RECT 877.950 133.950 880.050 136.050 ;
        RECT 880.950 133.950 883.050 136.050 ;
        RECT 827.550 131.550 832.050 133.050 ;
        RECT 833.100 132.150 834.900 133.950 ;
        RECT 828.000 130.950 832.050 131.550 ;
        RECT 835.950 129.750 837.150 133.950 ;
        RECT 839.100 132.150 840.900 133.950 ;
        RECT 844.950 132.450 847.050 133.050 ;
        RECT 850.950 132.450 853.050 133.050 ;
        RECT 844.950 131.550 853.050 132.450 ;
        RECT 844.950 130.950 847.050 131.550 ;
        RECT 850.950 130.950 853.050 131.550 ;
        RECT 833.400 128.700 837.150 129.750 ;
        RECT 833.400 126.600 834.600 128.700 ;
        RECT 814.800 120.600 816.600 123.600 ;
        RECT 832.800 120.600 834.600 126.600 ;
        RECT 835.800 125.700 843.600 127.050 ;
        RECT 835.800 120.600 837.600 125.700 ;
        RECT 841.800 120.600 843.600 125.700 ;
        RECT 857.400 123.600 858.600 133.950 ;
        RECT 872.100 132.150 873.900 133.950 ;
        RECT 878.100 132.150 879.900 133.950 ;
        RECT 881.400 130.200 882.300 133.950 ;
        RECT 883.950 132.450 886.050 133.050 ;
        RECT 889.950 132.450 892.050 133.050 ;
        RECT 883.950 131.550 892.050 132.450 ;
        RECT 883.950 130.950 886.050 131.550 ;
        RECT 889.950 130.950 892.050 131.550 ;
        RECT 856.800 120.600 858.600 123.600 ;
        RECT 879.000 129.000 882.300 130.200 ;
        RECT 879.000 120.600 880.800 129.000 ;
        RECT 13.800 110.400 15.600 116.400 ;
        RECT 21.300 110.400 23.100 116.400 ;
        RECT 28.800 110.400 30.600 116.400 ;
        RECT 46.800 113.400 48.600 116.400 ;
        RECT 13.800 109.500 18.600 110.400 ;
        RECT 16.500 108.300 18.600 109.500 ;
        RECT 21.600 108.900 22.800 110.400 ;
        RECT 19.800 106.800 22.800 108.900 ;
        RECT 28.800 108.600 30.000 110.400 ;
        RECT 18.750 103.800 20.850 105.900 ;
        RECT 4.950 102.450 7.050 103.050 ;
        RECT 13.950 102.450 16.050 103.050 ;
        RECT 4.950 101.550 16.050 102.450 ;
        RECT 18.600 102.000 20.400 103.800 ;
        RECT 4.950 100.950 7.050 101.550 ;
        RECT 13.950 100.950 16.050 101.550 ;
        RECT 21.750 101.100 22.800 106.800 ;
        RECT 23.700 107.700 30.000 108.600 ;
        RECT 23.700 105.600 25.800 107.700 ;
        RECT 23.700 103.800 25.500 105.600 ;
        RECT 28.800 103.050 30.600 104.850 ;
        RECT 47.400 103.050 48.300 113.400 ;
        RECT 65.400 109.200 67.200 116.400 ;
        RECT 88.800 113.400 90.600 116.400 ;
        RECT 107.400 113.400 109.200 116.400 ;
        RECT 127.800 113.400 129.600 116.400 ;
        RECT 143.400 113.400 145.200 116.400 ;
        RECT 65.400 108.300 69.600 109.200 ;
        RECT 65.100 103.050 66.900 104.850 ;
        RECT 68.400 103.050 69.600 108.300 ;
        RECT 71.100 103.050 72.900 104.850 ;
        RECT 89.400 103.050 90.300 113.400 ;
        RECT 107.400 103.050 108.600 113.400 ;
        RECT 128.400 103.050 129.300 113.400 ;
        RECT 143.400 109.500 144.600 113.400 ;
        RECT 149.400 110.400 151.200 116.400 ;
        RECT 169.800 113.400 171.600 116.400 ;
        RECT 190.800 113.400 192.600 116.400 ;
        RECT 211.800 113.400 213.600 116.400 ;
        RECT 143.400 108.600 149.100 109.500 ;
        RECT 147.150 107.700 149.100 108.600 ;
        RECT 28.500 102.300 34.050 103.050 ;
        RECT 14.100 99.150 15.900 100.950 ;
        RECT 20.400 100.200 22.800 101.100 ;
        RECT 23.700 101.100 34.050 102.300 ;
        RECT 23.700 100.500 25.500 101.100 ;
        RECT 28.500 100.950 34.050 101.100 ;
        RECT 43.950 100.950 46.050 103.050 ;
        RECT 46.950 100.950 49.050 103.050 ;
        RECT 49.950 100.950 52.050 103.050 ;
        RECT 64.950 100.950 67.050 103.050 ;
        RECT 67.950 100.950 70.050 103.050 ;
        RECT 70.950 100.950 73.050 103.050 ;
        RECT 85.950 100.950 88.050 103.050 ;
        RECT 88.950 100.950 91.050 103.050 ;
        RECT 91.950 100.950 94.050 103.050 ;
        RECT 103.950 100.950 106.050 103.050 ;
        RECT 106.950 100.950 109.050 103.050 ;
        RECT 124.950 100.950 127.050 103.050 ;
        RECT 127.950 100.950 130.050 103.050 ;
        RECT 130.950 100.950 133.050 103.050 ;
        RECT 142.950 100.950 145.050 103.050 ;
        RECT 19.800 98.100 21.900 100.200 ;
        RECT 21.000 96.000 21.900 98.100 ;
        RECT 22.800 97.500 26.700 99.300 ;
        RECT 44.100 99.150 45.900 100.950 ;
        RECT 22.800 97.200 24.900 97.500 ;
        RECT 21.000 95.100 22.500 96.000 ;
        RECT 16.500 93.600 18.600 94.500 ;
        RECT 13.800 92.400 18.600 93.600 ;
        RECT 21.300 93.600 22.500 95.100 ;
        RECT 26.100 93.600 28.200 95.700 ;
        RECT 47.400 93.600 48.300 100.950 ;
        RECT 50.100 99.150 51.900 100.950 ;
        RECT 13.800 81.600 15.600 92.400 ;
        RECT 21.300 81.600 23.100 93.600 ;
        RECT 26.100 92.700 30.600 93.600 ;
        RECT 28.800 81.600 30.600 92.700 ;
        RECT 44.700 92.400 48.300 93.600 ;
        RECT 44.700 81.600 46.500 92.400 ;
        RECT 68.400 87.600 69.600 100.950 ;
        RECT 86.100 99.150 87.900 100.950 ;
        RECT 89.400 93.600 90.300 100.950 ;
        RECT 92.100 99.150 93.900 100.950 ;
        RECT 104.100 99.150 105.900 100.950 ;
        RECT 67.800 81.600 69.600 87.600 ;
        RECT 86.700 92.400 90.300 93.600 ;
        RECT 86.700 81.600 88.500 92.400 ;
        RECT 107.400 87.600 108.600 100.950 ;
        RECT 125.100 99.150 126.900 100.950 ;
        RECT 128.400 93.600 129.300 100.950 ;
        RECT 131.100 99.150 132.900 100.950 ;
        RECT 143.100 99.150 144.900 100.950 ;
        RECT 147.150 96.300 148.050 107.700 ;
        RECT 150.000 103.050 151.200 110.400 ;
        RECT 170.400 103.050 171.300 113.400 ;
        RECT 191.400 103.050 192.300 113.400 ;
        RECT 212.400 103.050 213.600 113.400 ;
        RECT 218.550 110.400 220.350 116.400 ;
        RECT 226.650 113.400 228.450 116.400 ;
        RECT 234.450 113.400 236.250 116.400 ;
        RECT 242.250 114.300 244.050 116.400 ;
        RECT 242.250 113.400 246.000 114.300 ;
        RECT 226.650 112.500 227.700 113.400 ;
        RECT 223.950 111.300 227.700 112.500 ;
        RECT 235.200 112.500 236.250 113.400 ;
        RECT 244.950 112.500 246.000 113.400 ;
        RECT 235.200 111.450 240.150 112.500 ;
        RECT 223.950 110.400 226.050 111.300 ;
        RECT 238.350 110.700 240.150 111.450 ;
        RECT 218.550 103.050 219.750 110.400 ;
        RECT 241.650 109.800 243.450 111.600 ;
        RECT 244.950 110.400 247.050 112.500 ;
        RECT 250.050 110.400 251.850 116.400 ;
        RECT 231.150 108.000 232.950 108.600 ;
        RECT 242.100 108.000 243.150 109.800 ;
        RECT 231.150 106.800 243.150 108.000 ;
        RECT 148.950 100.950 151.200 103.050 ;
        RECT 166.950 100.950 169.050 103.050 ;
        RECT 169.950 100.950 172.050 103.050 ;
        RECT 172.950 100.950 175.050 103.050 ;
        RECT 187.950 100.950 190.050 103.050 ;
        RECT 190.950 100.950 193.050 103.050 ;
        RECT 193.950 100.950 196.050 103.050 ;
        RECT 211.950 100.950 214.050 103.050 ;
        RECT 214.950 100.950 217.050 103.050 ;
        RECT 218.550 101.250 224.850 103.050 ;
        RECT 218.550 100.950 223.050 101.250 ;
        RECT 147.150 95.400 149.100 96.300 ;
        RECT 125.700 92.400 129.300 93.600 ;
        RECT 143.400 94.500 149.100 95.400 ;
        RECT 107.400 81.600 109.200 87.600 ;
        RECT 125.700 81.600 127.500 92.400 ;
        RECT 143.400 87.600 144.600 94.500 ;
        RECT 150.000 93.600 151.200 100.950 ;
        RECT 167.100 99.150 168.900 100.950 ;
        RECT 170.400 93.600 171.300 100.950 ;
        RECT 173.100 99.150 174.900 100.950 ;
        RECT 188.100 99.150 189.900 100.950 ;
        RECT 191.400 93.600 192.300 100.950 ;
        RECT 194.100 99.150 195.900 100.950 ;
        RECT 143.400 81.600 145.200 87.600 ;
        RECT 149.400 81.600 151.200 93.600 ;
        RECT 167.700 92.400 171.300 93.600 ;
        RECT 188.700 92.400 192.300 93.600 ;
        RECT 167.700 81.600 169.500 92.400 ;
        RECT 188.700 81.600 190.500 92.400 ;
        RECT 212.400 87.600 213.600 100.950 ;
        RECT 215.100 99.150 216.900 100.950 ;
        RECT 211.800 81.600 213.600 87.600 ;
        RECT 218.550 93.600 219.750 100.950 ;
        RECT 220.950 95.400 222.750 97.200 ;
        RECT 221.850 94.200 226.050 95.400 ;
        RECT 231.150 94.200 232.050 106.800 ;
        RECT 242.100 105.600 249.000 106.800 ;
        RECT 242.100 105.000 243.900 105.600 ;
        RECT 248.100 104.850 249.000 105.600 ;
        RECT 245.100 103.800 246.900 104.400 ;
        RECT 238.950 102.600 246.900 103.800 ;
        RECT 248.100 103.050 249.900 104.850 ;
        RECT 238.950 100.950 241.050 102.600 ;
        RECT 247.950 100.950 250.050 103.050 ;
        RECT 240.750 95.700 242.550 96.000 ;
        RECT 250.950 95.700 251.850 110.400 ;
        RECT 263.400 111.300 265.200 116.400 ;
        RECT 269.400 111.300 271.200 116.400 ;
        RECT 263.400 109.950 271.200 111.300 ;
        RECT 272.400 110.400 274.200 116.400 ;
        RECT 289.800 113.400 291.600 116.400 ;
        RECT 272.400 108.300 273.600 110.400 ;
        RECT 269.850 107.250 273.600 108.300 ;
        RECT 266.100 103.050 267.900 104.850 ;
        RECT 269.850 103.050 271.050 107.250 ;
        RECT 272.100 103.050 273.900 104.850 ;
        RECT 290.400 103.050 291.600 113.400 ;
        RECT 296.550 110.400 298.350 116.400 ;
        RECT 304.650 113.400 306.450 116.400 ;
        RECT 312.450 113.400 314.250 116.400 ;
        RECT 320.250 114.300 322.050 116.400 ;
        RECT 320.250 113.400 324.000 114.300 ;
        RECT 304.650 112.500 305.700 113.400 ;
        RECT 301.950 111.300 305.700 112.500 ;
        RECT 313.200 112.500 314.250 113.400 ;
        RECT 322.950 112.500 324.000 113.400 ;
        RECT 313.200 111.450 318.150 112.500 ;
        RECT 301.950 110.400 304.050 111.300 ;
        RECT 316.350 110.700 318.150 111.450 ;
        RECT 296.550 103.050 297.750 110.400 ;
        RECT 319.650 109.800 321.450 111.600 ;
        RECT 322.950 110.400 325.050 112.500 ;
        RECT 328.050 110.400 329.850 116.400 ;
        RECT 309.150 108.000 310.950 108.600 ;
        RECT 320.100 108.000 321.150 109.800 ;
        RECT 309.150 106.800 321.150 108.000 ;
        RECT 262.950 100.950 265.050 103.050 ;
        RECT 265.950 100.950 268.050 103.050 ;
        RECT 268.950 100.950 271.050 103.050 ;
        RECT 271.950 100.950 274.050 103.050 ;
        RECT 289.950 100.950 292.050 103.050 ;
        RECT 292.950 100.950 295.050 103.050 ;
        RECT 296.550 101.250 302.850 103.050 ;
        RECT 296.550 100.950 301.050 101.250 ;
        RECT 263.100 99.150 264.900 100.950 ;
        RECT 240.750 95.100 251.850 95.700 ;
        RECT 218.550 81.600 220.350 93.600 ;
        RECT 223.950 93.300 226.050 94.200 ;
        RECT 226.950 93.300 232.050 94.200 ;
        RECT 234.150 94.500 251.850 95.100 ;
        RECT 234.150 94.200 242.550 94.500 ;
        RECT 226.950 92.400 227.850 93.300 ;
        RECT 225.150 90.600 227.850 92.400 ;
        RECT 228.750 92.100 230.550 92.400 ;
        RECT 234.150 92.100 235.050 94.200 ;
        RECT 250.950 93.600 251.850 94.500 ;
        RECT 228.750 91.200 235.050 92.100 ;
        RECT 235.950 92.700 237.750 93.300 ;
        RECT 235.950 91.500 243.450 92.700 ;
        RECT 228.750 90.600 230.550 91.200 ;
        RECT 242.250 90.600 243.450 91.500 ;
        RECT 223.950 87.600 227.850 89.700 ;
        RECT 232.950 89.550 234.750 90.300 ;
        RECT 237.750 89.550 239.550 90.300 ;
        RECT 232.950 88.500 239.550 89.550 ;
        RECT 242.250 88.500 247.050 90.600 ;
        RECT 226.050 81.600 227.850 87.600 ;
        RECT 233.850 81.600 235.650 88.500 ;
        RECT 242.250 87.600 243.450 88.500 ;
        RECT 241.650 81.600 243.450 87.600 ;
        RECT 250.050 81.600 251.850 93.600 ;
        RECT 268.950 87.600 270.150 100.950 ;
        RECT 290.400 87.600 291.600 100.950 ;
        RECT 293.100 99.150 294.900 100.950 ;
        RECT 268.800 81.600 270.600 87.600 ;
        RECT 289.800 81.600 291.600 87.600 ;
        RECT 296.550 93.600 297.750 100.950 ;
        RECT 298.950 95.400 300.750 97.200 ;
        RECT 299.850 94.200 304.050 95.400 ;
        RECT 309.150 94.200 310.050 106.800 ;
        RECT 320.100 105.600 327.000 106.800 ;
        RECT 320.100 105.000 321.900 105.600 ;
        RECT 326.100 104.850 327.000 105.600 ;
        RECT 323.100 103.800 324.900 104.400 ;
        RECT 316.950 102.600 324.900 103.800 ;
        RECT 326.100 103.050 327.900 104.850 ;
        RECT 316.950 100.950 319.050 102.600 ;
        RECT 325.950 100.950 328.050 103.050 ;
        RECT 318.750 95.700 320.550 96.000 ;
        RECT 328.950 95.700 329.850 110.400 ;
        RECT 341.400 111.000 343.200 116.400 ;
        RECT 347.400 115.500 355.200 116.400 ;
        RECT 347.400 111.000 349.200 115.500 ;
        RECT 341.400 110.100 349.200 111.000 ;
        RECT 350.400 110.400 352.200 114.600 ;
        RECT 353.400 110.400 355.200 115.500 ;
        RECT 373.800 113.400 375.600 116.400 ;
        RECT 350.700 108.900 351.600 110.400 ;
        RECT 346.950 107.700 351.600 108.900 ;
        RECT 344.100 103.050 345.900 104.850 ;
        RECT 346.950 103.050 348.300 107.700 ;
        RECT 350.100 103.050 351.900 104.850 ;
        RECT 374.400 103.050 375.300 113.400 ;
        RECT 380.550 110.400 382.350 116.400 ;
        RECT 388.650 113.400 390.450 116.400 ;
        RECT 396.450 113.400 398.250 116.400 ;
        RECT 404.250 114.300 406.050 116.400 ;
        RECT 404.250 113.400 408.000 114.300 ;
        RECT 388.650 112.500 389.700 113.400 ;
        RECT 385.950 111.300 389.700 112.500 ;
        RECT 397.200 112.500 398.250 113.400 ;
        RECT 406.950 112.500 408.000 113.400 ;
        RECT 397.200 111.450 402.150 112.500 ;
        RECT 385.950 110.400 388.050 111.300 ;
        RECT 400.350 110.700 402.150 111.450 ;
        RECT 380.550 103.050 381.750 110.400 ;
        RECT 403.650 109.800 405.450 111.600 ;
        RECT 406.950 110.400 409.050 112.500 ;
        RECT 412.050 110.400 413.850 116.400 ;
        RECT 431.700 111.600 433.500 116.400 ;
        RECT 454.800 113.400 456.600 116.400 ;
        RECT 393.150 108.000 394.950 108.600 ;
        RECT 404.100 108.000 405.150 109.800 ;
        RECT 393.150 106.800 405.150 108.000 ;
        RECT 340.950 100.950 343.050 103.050 ;
        RECT 343.950 100.950 346.050 103.050 ;
        RECT 346.950 100.950 349.050 103.050 ;
        RECT 349.950 100.950 352.050 103.050 ;
        RECT 352.950 100.950 355.050 103.050 ;
        RECT 370.950 100.950 373.050 103.050 ;
        RECT 373.950 100.950 376.050 103.050 ;
        RECT 376.950 100.950 379.050 103.050 ;
        RECT 380.550 101.250 386.850 103.050 ;
        RECT 380.550 100.950 385.050 101.250 ;
        RECT 341.100 99.150 342.900 100.950 ;
        RECT 318.750 95.100 329.850 95.700 ;
        RECT 296.550 81.600 298.350 93.600 ;
        RECT 301.950 93.300 304.050 94.200 ;
        RECT 304.950 93.300 310.050 94.200 ;
        RECT 312.150 94.500 329.850 95.100 ;
        RECT 312.150 94.200 320.550 94.500 ;
        RECT 304.950 92.400 305.850 93.300 ;
        RECT 303.150 90.600 305.850 92.400 ;
        RECT 306.750 92.100 308.550 92.400 ;
        RECT 312.150 92.100 313.050 94.200 ;
        RECT 328.950 93.600 329.850 94.500 ;
        RECT 347.100 93.600 348.300 100.950 ;
        RECT 353.100 99.150 354.900 100.950 ;
        RECT 371.100 99.150 372.900 100.950 ;
        RECT 374.400 93.600 375.300 100.950 ;
        RECT 377.100 99.150 378.900 100.950 ;
        RECT 306.750 91.200 313.050 92.100 ;
        RECT 313.950 92.700 315.750 93.300 ;
        RECT 313.950 91.500 321.450 92.700 ;
        RECT 306.750 90.600 308.550 91.200 ;
        RECT 320.250 90.600 321.450 91.500 ;
        RECT 301.950 87.600 305.850 89.700 ;
        RECT 310.950 89.550 312.750 90.300 ;
        RECT 315.750 89.550 317.550 90.300 ;
        RECT 310.950 88.500 317.550 89.550 ;
        RECT 320.250 88.500 325.050 90.600 ;
        RECT 304.050 81.600 305.850 87.600 ;
        RECT 311.850 81.600 313.650 88.500 ;
        RECT 320.250 87.600 321.450 88.500 ;
        RECT 319.650 81.600 321.450 87.600 ;
        RECT 328.050 81.600 329.850 93.600 ;
        RECT 345.900 81.600 349.200 93.600 ;
        RECT 371.700 92.400 375.300 93.600 ;
        RECT 380.550 93.600 381.750 100.950 ;
        RECT 382.950 95.400 384.750 97.200 ;
        RECT 383.850 94.200 388.050 95.400 ;
        RECT 393.150 94.200 394.050 106.800 ;
        RECT 404.100 105.600 411.000 106.800 ;
        RECT 404.100 105.000 405.900 105.600 ;
        RECT 410.100 104.850 411.000 105.600 ;
        RECT 407.100 103.800 408.900 104.400 ;
        RECT 400.950 102.600 408.900 103.800 ;
        RECT 410.100 103.050 411.900 104.850 ;
        RECT 400.950 100.950 403.050 102.600 ;
        RECT 409.950 100.950 412.050 103.050 ;
        RECT 402.750 95.700 404.550 96.000 ;
        RECT 412.950 95.700 413.850 110.400 ;
        RECT 428.400 110.400 433.500 111.600 ;
        RECT 428.400 103.050 429.300 110.400 ;
        RECT 431.100 103.050 432.900 104.850 ;
        RECT 437.100 103.050 438.900 104.850 ;
        RECT 455.400 103.050 456.300 113.400 ;
        RECT 472.800 110.400 474.600 116.400 ;
        RECT 473.400 108.300 474.600 110.400 ;
        RECT 475.800 111.300 477.600 116.400 ;
        RECT 481.800 111.300 483.600 116.400 ;
        RECT 475.800 109.950 483.600 111.300 ;
        RECT 497.400 113.400 499.200 116.400 ;
        RECT 517.800 113.400 519.600 116.400 ;
        RECT 473.400 107.250 477.150 108.300 ;
        RECT 473.100 103.050 474.900 104.850 ;
        RECT 475.950 103.050 477.150 107.250 ;
        RECT 479.100 103.050 480.900 104.850 ;
        RECT 497.400 103.050 498.600 113.400 ;
        RECT 518.400 103.050 519.300 113.400 ;
        RECT 533.400 111.300 535.200 116.400 ;
        RECT 539.400 111.300 541.200 116.400 ;
        RECT 533.400 109.950 541.200 111.300 ;
        RECT 542.400 110.400 544.200 116.400 ;
        RECT 559.800 113.400 561.600 116.400 ;
        RECT 542.400 108.300 543.600 110.400 ;
        RECT 539.850 107.250 543.600 108.300 ;
        RECT 536.100 103.050 537.900 104.850 ;
        RECT 539.850 103.050 541.050 107.250 ;
        RECT 542.100 103.050 543.900 104.850 ;
        RECT 560.400 103.050 561.600 113.400 ;
        RECT 575.400 108.600 577.200 116.400 ;
        RECT 582.900 112.200 584.700 116.400 ;
        RECT 589.950 112.950 595.050 115.050 ;
        RECT 582.900 110.400 585.600 112.200 ;
        RECT 581.100 108.600 582.900 109.500 ;
        RECT 575.400 107.700 582.900 108.600 ;
        RECT 575.100 103.050 576.900 104.850 ;
        RECT 427.950 100.950 430.050 103.050 ;
        RECT 430.950 100.950 433.050 103.050 ;
        RECT 433.950 100.950 436.050 103.050 ;
        RECT 436.950 100.950 439.050 103.050 ;
        RECT 451.950 100.950 454.050 103.050 ;
        RECT 454.950 100.950 457.050 103.050 ;
        RECT 457.950 100.950 460.050 103.050 ;
        RECT 472.950 100.950 475.050 103.050 ;
        RECT 475.950 100.950 478.050 103.050 ;
        RECT 478.950 100.950 481.050 103.050 ;
        RECT 481.950 100.950 484.050 103.050 ;
        RECT 493.950 100.950 496.050 103.050 ;
        RECT 496.950 100.950 499.050 103.050 ;
        RECT 514.950 100.950 517.050 103.050 ;
        RECT 517.950 100.950 520.050 103.050 ;
        RECT 520.950 100.950 523.050 103.050 ;
        RECT 532.950 100.950 535.050 103.050 ;
        RECT 535.950 100.950 538.050 103.050 ;
        RECT 538.950 100.950 541.050 103.050 ;
        RECT 541.950 100.950 544.050 103.050 ;
        RECT 559.950 100.950 562.050 103.050 ;
        RECT 562.950 100.950 565.050 103.050 ;
        RECT 574.950 100.950 577.050 103.050 ;
        RECT 402.750 95.100 413.850 95.700 ;
        RECT 371.700 81.600 373.500 92.400 ;
        RECT 380.550 81.600 382.350 93.600 ;
        RECT 385.950 93.300 388.050 94.200 ;
        RECT 388.950 93.300 394.050 94.200 ;
        RECT 396.150 94.500 413.850 95.100 ;
        RECT 396.150 94.200 404.550 94.500 ;
        RECT 388.950 92.400 389.850 93.300 ;
        RECT 387.150 90.600 389.850 92.400 ;
        RECT 390.750 92.100 392.550 92.400 ;
        RECT 396.150 92.100 397.050 94.200 ;
        RECT 412.950 93.600 413.850 94.500 ;
        RECT 428.400 93.600 429.300 100.950 ;
        RECT 434.100 99.150 435.900 100.950 ;
        RECT 452.100 99.150 453.900 100.950 ;
        RECT 455.400 93.600 456.300 100.950 ;
        RECT 458.100 99.150 459.900 100.950 ;
        RECT 390.750 91.200 397.050 92.100 ;
        RECT 397.950 92.700 399.750 93.300 ;
        RECT 397.950 91.500 405.450 92.700 ;
        RECT 390.750 90.600 392.550 91.200 ;
        RECT 404.250 90.600 405.450 91.500 ;
        RECT 385.950 87.600 389.850 89.700 ;
        RECT 394.950 89.550 396.750 90.300 ;
        RECT 399.750 89.550 401.550 90.300 ;
        RECT 394.950 88.500 401.550 89.550 ;
        RECT 404.250 88.500 409.050 90.600 ;
        RECT 388.050 81.600 389.850 87.600 ;
        RECT 395.850 81.600 397.650 88.500 ;
        RECT 404.250 87.600 405.450 88.500 ;
        RECT 403.650 81.600 405.450 87.600 ;
        RECT 412.050 81.600 413.850 93.600 ;
        RECT 427.800 81.600 429.600 93.600 ;
        RECT 430.800 92.700 438.600 93.600 ;
        RECT 430.800 81.600 432.600 92.700 ;
        RECT 436.800 81.600 438.600 92.700 ;
        RECT 452.700 92.400 456.300 93.600 ;
        RECT 452.700 81.600 454.500 92.400 ;
        RECT 476.850 87.600 478.050 100.950 ;
        RECT 482.100 99.150 483.900 100.950 ;
        RECT 494.100 99.150 495.900 100.950 ;
        RECT 497.400 87.600 498.600 100.950 ;
        RECT 505.950 99.450 508.050 100.050 ;
        RECT 511.950 99.450 514.050 100.050 ;
        RECT 505.950 98.550 514.050 99.450 ;
        RECT 515.100 99.150 516.900 100.950 ;
        RECT 505.950 97.950 508.050 98.550 ;
        RECT 511.950 97.950 514.050 98.550 ;
        RECT 518.400 93.600 519.300 100.950 ;
        RECT 521.100 99.150 522.900 100.950 ;
        RECT 533.100 99.150 534.900 100.950 ;
        RECT 515.700 92.400 519.300 93.600 ;
        RECT 476.400 81.600 478.200 87.600 ;
        RECT 497.400 81.600 499.200 87.600 ;
        RECT 515.700 81.600 517.500 92.400 ;
        RECT 538.950 87.600 540.150 100.950 ;
        RECT 560.400 87.600 561.600 100.950 ;
        RECT 563.100 99.150 564.900 100.950 ;
        RECT 538.800 81.600 540.600 87.600 ;
        RECT 559.800 81.600 561.600 87.600 ;
        RECT 578.400 87.600 579.300 107.700 ;
        RECT 584.700 103.050 585.600 110.400 ;
        RECT 602.400 109.200 604.200 116.400 ;
        RECT 626.400 113.400 628.200 116.400 ;
        RECT 646.800 113.400 648.600 116.400 ;
        RECT 602.400 108.300 606.600 109.200 ;
        RECT 602.100 103.050 603.900 104.850 ;
        RECT 605.400 103.050 606.600 108.300 ;
        RECT 608.100 103.050 609.900 104.850 ;
        RECT 626.700 103.050 627.600 113.400 ;
        RECT 647.400 103.050 648.600 113.400 ;
        RECT 653.550 110.400 655.350 116.400 ;
        RECT 661.650 113.400 663.450 116.400 ;
        RECT 669.450 113.400 671.250 116.400 ;
        RECT 677.250 114.300 679.050 116.400 ;
        RECT 677.250 113.400 681.000 114.300 ;
        RECT 661.650 112.500 662.700 113.400 ;
        RECT 658.950 111.300 662.700 112.500 ;
        RECT 670.200 112.500 671.250 113.400 ;
        RECT 679.950 112.500 681.000 113.400 ;
        RECT 670.200 111.450 675.150 112.500 ;
        RECT 658.950 110.400 661.050 111.300 ;
        RECT 673.350 110.700 675.150 111.450 ;
        RECT 653.550 103.050 654.750 110.400 ;
        RECT 676.650 109.800 678.450 111.600 ;
        RECT 679.950 110.400 682.050 112.500 ;
        RECT 685.050 110.400 686.850 116.400 ;
        RECT 666.150 108.000 667.950 108.600 ;
        RECT 677.100 108.000 678.150 109.800 ;
        RECT 666.150 106.800 678.150 108.000 ;
        RECT 580.950 100.950 583.050 103.050 ;
        RECT 583.950 100.950 586.050 103.050 ;
        RECT 601.950 100.950 604.050 103.050 ;
        RECT 604.950 100.950 607.050 103.050 ;
        RECT 607.950 100.950 610.050 103.050 ;
        RECT 622.950 100.950 625.050 103.050 ;
        RECT 625.950 100.950 628.050 103.050 ;
        RECT 628.950 100.950 631.050 103.050 ;
        RECT 646.950 100.950 649.050 103.050 ;
        RECT 649.950 100.950 652.050 103.050 ;
        RECT 653.550 101.250 659.850 103.050 ;
        RECT 653.550 100.950 658.050 101.250 ;
        RECT 581.100 99.150 582.900 100.950 ;
        RECT 584.700 93.600 585.600 100.950 ;
        RECT 578.400 81.600 580.200 87.600 ;
        RECT 584.400 81.600 586.200 93.600 ;
        RECT 605.400 87.600 606.600 100.950 ;
        RECT 623.100 99.150 624.900 100.950 ;
        RECT 626.700 93.600 627.600 100.950 ;
        RECT 629.100 99.150 630.900 100.950 ;
        RECT 626.700 92.400 630.300 93.600 ;
        RECT 604.800 81.600 606.600 87.600 ;
        RECT 628.500 81.600 630.300 92.400 ;
        RECT 647.400 87.600 648.600 100.950 ;
        RECT 650.100 99.150 651.900 100.950 ;
        RECT 646.800 81.600 648.600 87.600 ;
        RECT 653.550 93.600 654.750 100.950 ;
        RECT 655.950 95.400 657.750 97.200 ;
        RECT 656.850 94.200 661.050 95.400 ;
        RECT 666.150 94.200 667.050 106.800 ;
        RECT 677.100 105.600 684.000 106.800 ;
        RECT 677.100 105.000 678.900 105.600 ;
        RECT 683.100 104.850 684.000 105.600 ;
        RECT 680.100 103.800 681.900 104.400 ;
        RECT 673.950 102.600 681.900 103.800 ;
        RECT 683.100 103.050 684.900 104.850 ;
        RECT 673.950 100.950 676.050 102.600 ;
        RECT 682.950 100.950 685.050 103.050 ;
        RECT 675.750 95.700 677.550 96.000 ;
        RECT 685.950 95.700 686.850 110.400 ;
        RECT 703.200 108.000 705.000 116.400 ;
        RECT 727.800 109.200 729.600 116.400 ;
        RECT 743.400 110.400 745.200 116.400 ;
        RECT 750.900 110.400 752.700 116.400 ;
        RECT 758.400 110.400 760.200 116.400 ;
        RECT 778.500 111.600 780.300 116.400 ;
        RECT 778.500 110.400 783.600 111.600 ;
        RECT 701.700 106.800 705.000 108.000 ;
        RECT 725.400 108.300 729.600 109.200 ;
        RECT 744.000 108.600 745.200 110.400 ;
        RECT 751.200 108.900 752.400 110.400 ;
        RECT 755.400 109.500 760.200 110.400 ;
        RECT 701.700 103.050 702.600 106.800 ;
        RECT 704.100 103.050 705.900 104.850 ;
        RECT 710.100 103.050 711.900 104.850 ;
        RECT 722.100 103.050 723.900 104.850 ;
        RECT 725.400 103.050 726.600 108.300 ;
        RECT 744.000 107.700 750.300 108.600 ;
        RECT 730.950 105.450 735.000 106.050 ;
        RECT 748.200 105.600 750.300 107.700 ;
        RECT 728.100 103.050 729.900 104.850 ;
        RECT 730.950 103.950 735.450 105.450 ;
        RECT 700.950 100.950 703.050 103.050 ;
        RECT 703.950 100.950 706.050 103.050 ;
        RECT 706.950 100.950 709.050 103.050 ;
        RECT 709.950 100.950 712.050 103.050 ;
        RECT 721.950 100.950 724.050 103.050 ;
        RECT 724.950 100.950 727.050 103.050 ;
        RECT 727.950 100.950 730.050 103.050 ;
        RECT 675.750 95.100 686.850 95.700 ;
        RECT 653.550 81.600 655.350 93.600 ;
        RECT 658.950 93.300 661.050 94.200 ;
        RECT 661.950 93.300 667.050 94.200 ;
        RECT 669.150 94.500 686.850 95.100 ;
        RECT 669.150 94.200 677.550 94.500 ;
        RECT 661.950 92.400 662.850 93.300 ;
        RECT 660.150 90.600 662.850 92.400 ;
        RECT 663.750 92.100 665.550 92.400 ;
        RECT 669.150 92.100 670.050 94.200 ;
        RECT 685.950 93.600 686.850 94.500 ;
        RECT 663.750 91.200 670.050 92.100 ;
        RECT 670.950 92.700 672.750 93.300 ;
        RECT 670.950 91.500 678.450 92.700 ;
        RECT 663.750 90.600 665.550 91.200 ;
        RECT 677.250 90.600 678.450 91.500 ;
        RECT 658.950 87.600 662.850 89.700 ;
        RECT 667.950 89.550 669.750 90.300 ;
        RECT 672.750 89.550 674.550 90.300 ;
        RECT 667.950 88.500 674.550 89.550 ;
        RECT 677.250 88.500 682.050 90.600 ;
        RECT 661.050 81.600 662.850 87.600 ;
        RECT 668.850 81.600 670.650 88.500 ;
        RECT 677.250 87.600 678.450 88.500 ;
        RECT 676.650 81.600 678.450 87.600 ;
        RECT 685.050 81.600 686.850 93.600 ;
        RECT 701.700 88.800 702.600 100.950 ;
        RECT 707.100 99.150 708.900 100.950 ;
        RECT 701.700 87.900 708.300 88.800 ;
        RECT 701.700 87.600 702.600 87.900 ;
        RECT 700.800 81.600 702.600 87.600 ;
        RECT 706.800 87.600 708.300 87.900 ;
        RECT 725.400 87.600 726.600 100.950 ;
        RECT 734.550 100.050 735.450 103.950 ;
        RECT 743.400 103.050 745.200 104.850 ;
        RECT 748.500 103.800 750.300 105.600 ;
        RECT 751.200 106.800 754.200 108.900 ;
        RECT 755.400 108.300 757.500 109.500 ;
        RECT 743.400 102.300 745.500 103.050 ;
        RECT 743.400 101.100 750.300 102.300 ;
        RECT 743.400 100.950 745.500 101.100 ;
        RECT 748.500 100.500 750.300 101.100 ;
        RECT 751.200 101.100 752.250 106.800 ;
        RECT 753.150 103.800 755.250 105.900 ;
        RECT 769.950 105.450 772.050 106.050 ;
        RECT 764.550 104.550 772.050 105.450 ;
        RECT 753.600 102.000 755.400 103.800 ;
        RECT 757.950 102.450 760.050 103.050 ;
        RECT 764.550 102.450 765.450 104.550 ;
        RECT 769.950 103.950 772.050 104.550 ;
        RECT 773.100 103.050 774.900 104.850 ;
        RECT 779.100 103.050 780.900 104.850 ;
        RECT 782.700 103.050 783.600 110.400 ;
        RECT 784.950 111.450 787.050 112.050 ;
        RECT 802.500 111.600 804.300 116.400 ;
        RECT 826.800 113.400 828.600 116.400 ;
        RECT 845.400 113.400 847.200 116.400 ;
        RECT 866.400 113.400 868.200 116.400 ;
        RECT 887.400 113.400 889.200 116.400 ;
        RECT 784.950 110.550 792.450 111.450 ;
        RECT 784.950 109.950 787.050 110.550 ;
        RECT 757.950 101.550 765.450 102.450 ;
        RECT 751.200 100.200 753.600 101.100 ;
        RECT 757.950 100.950 760.050 101.550 ;
        RECT 772.950 100.950 775.050 103.050 ;
        RECT 775.950 100.950 778.050 103.050 ;
        RECT 778.950 100.950 781.050 103.050 ;
        RECT 781.950 100.950 784.050 103.050 ;
        RECT 730.950 98.550 735.450 100.050 ;
        RECT 730.950 97.950 735.000 98.550 ;
        RECT 747.300 97.500 751.200 99.300 ;
        RECT 749.100 97.200 751.200 97.500 ;
        RECT 752.100 98.100 754.200 100.200 ;
        RECT 758.100 99.150 759.900 100.950 ;
        RECT 776.100 99.150 777.900 100.950 ;
        RECT 752.100 96.000 753.000 98.100 ;
        RECT 745.800 93.600 747.900 95.700 ;
        RECT 751.500 95.100 753.000 96.000 ;
        RECT 763.950 96.450 766.050 97.050 ;
        RECT 778.950 96.450 781.050 97.050 ;
        RECT 763.950 95.550 781.050 96.450 ;
        RECT 751.500 93.600 752.700 95.100 ;
        RECT 763.950 94.950 766.050 95.550 ;
        RECT 778.950 94.950 781.050 95.550 ;
        RECT 743.400 92.700 747.900 93.600 ;
        RECT 706.800 81.600 708.600 87.600 ;
        RECT 725.400 81.600 727.200 87.600 ;
        RECT 743.400 81.600 745.200 92.700 ;
        RECT 750.900 85.050 752.700 93.600 ;
        RECT 755.400 93.600 757.500 94.500 ;
        RECT 782.700 93.600 783.600 100.950 ;
        RECT 791.550 99.450 792.450 110.550 ;
        RECT 802.500 110.400 807.600 111.600 ;
        RECT 797.100 103.050 798.900 104.850 ;
        RECT 803.100 103.050 804.900 104.850 ;
        RECT 806.700 103.050 807.600 110.400 ;
        RECT 817.950 111.450 820.050 112.050 ;
        RECT 823.950 111.450 826.050 112.050 ;
        RECT 817.950 110.550 826.050 111.450 ;
        RECT 817.950 109.950 820.050 110.550 ;
        RECT 823.950 109.950 826.050 110.550 ;
        RECT 827.400 103.050 828.300 113.400 ;
        RECT 829.950 108.450 832.050 109.200 ;
        RECT 829.950 107.550 837.450 108.450 ;
        RECT 829.950 107.100 832.050 107.550 ;
        RECT 796.950 100.950 799.050 103.050 ;
        RECT 799.950 100.950 802.050 103.050 ;
        RECT 802.950 100.950 805.050 103.050 ;
        RECT 805.950 100.950 808.050 103.050 ;
        RECT 823.950 100.950 826.050 103.050 ;
        RECT 826.950 100.950 829.050 103.050 ;
        RECT 829.950 100.950 832.050 103.050 ;
        RECT 791.550 98.550 795.450 99.450 ;
        RECT 800.100 99.150 801.900 100.950 ;
        RECT 784.950 96.450 787.050 97.050 ;
        RECT 790.950 96.450 793.050 97.050 ;
        RECT 784.950 95.550 793.050 96.450 ;
        RECT 794.550 96.450 795.450 98.550 ;
        RECT 799.950 96.450 802.050 97.050 ;
        RECT 794.550 95.550 802.050 96.450 ;
        RECT 784.950 94.950 787.050 95.550 ;
        RECT 790.950 94.950 793.050 95.550 ;
        RECT 799.950 94.950 802.050 95.550 ;
        RECT 806.700 93.600 807.600 100.950 ;
        RECT 824.100 99.150 825.900 100.950 ;
        RECT 827.400 93.600 828.300 100.950 ;
        RECT 830.100 99.150 831.900 100.950 ;
        RECT 836.550 99.450 837.450 107.550 ;
        RECT 845.700 103.050 846.600 113.400 ;
        RECT 853.950 108.450 856.050 109.050 ;
        RECT 862.950 108.450 865.050 109.050 ;
        RECT 853.950 107.550 865.050 108.450 ;
        RECT 853.950 106.950 856.050 107.550 ;
        RECT 862.950 106.950 865.050 107.550 ;
        RECT 866.700 103.050 867.600 113.400 ;
        RECT 879.000 105.450 883.050 106.050 ;
        RECT 878.550 103.950 883.050 105.450 ;
        RECT 841.950 100.950 844.050 103.050 ;
        RECT 844.950 100.950 847.050 103.050 ;
        RECT 847.950 100.950 850.050 103.050 ;
        RECT 862.950 100.950 865.050 103.050 ;
        RECT 865.950 100.950 868.050 103.050 ;
        RECT 868.950 100.950 871.050 103.050 ;
        RECT 836.550 98.550 840.450 99.450 ;
        RECT 842.100 99.150 843.900 100.950 ;
        RECT 839.550 97.050 840.450 98.550 ;
        RECT 839.550 95.550 844.050 97.050 ;
        RECT 840.000 94.950 844.050 95.550 ;
        RECT 755.400 92.400 760.200 93.600 ;
        RECT 750.900 82.950 754.050 85.050 ;
        RECT 750.900 81.600 752.700 82.950 ;
        RECT 758.400 81.600 760.200 92.400 ;
        RECT 773.400 92.700 781.200 93.600 ;
        RECT 773.400 81.600 775.200 92.700 ;
        RECT 779.400 81.600 781.200 92.700 ;
        RECT 782.400 81.600 784.200 93.600 ;
        RECT 797.400 92.700 805.200 93.600 ;
        RECT 797.400 81.600 799.200 92.700 ;
        RECT 803.400 81.600 805.200 92.700 ;
        RECT 806.400 81.600 808.200 93.600 ;
        RECT 824.700 92.400 828.300 93.600 ;
        RECT 845.700 93.600 846.600 100.950 ;
        RECT 848.100 99.150 849.900 100.950 ;
        RECT 863.100 99.150 864.900 100.950 ;
        RECT 866.700 93.600 867.600 100.950 ;
        RECT 869.100 99.150 870.900 100.950 ;
        RECT 878.550 96.450 879.450 103.950 ;
        RECT 887.400 103.050 888.600 113.400 ;
        RECT 883.950 100.950 886.050 103.050 ;
        RECT 886.950 100.950 889.050 103.050 ;
        RECT 884.100 99.150 885.900 100.950 ;
        RECT 883.950 96.450 886.050 97.050 ;
        RECT 878.550 95.550 886.050 96.450 ;
        RECT 883.950 94.950 886.050 95.550 ;
        RECT 845.700 92.400 849.300 93.600 ;
        RECT 866.700 92.400 870.300 93.600 ;
        RECT 824.700 81.600 826.500 92.400 ;
        RECT 847.500 81.600 849.300 92.400 ;
        RECT 868.500 81.600 870.300 92.400 ;
        RECT 887.400 87.600 888.600 100.950 ;
        RECT 887.400 81.600 889.200 87.600 ;
        RECT 14.700 66.600 16.500 77.400 ;
        RECT 37.500 66.600 39.300 77.400 ;
        RECT 14.700 65.400 18.300 66.600 ;
        RECT 14.100 58.050 15.900 59.850 ;
        RECT 17.400 58.050 18.300 65.400 ;
        RECT 35.700 65.400 39.300 66.600 ;
        RECT 53.400 66.300 55.200 77.400 ;
        RECT 59.400 66.300 61.200 77.400 ;
        RECT 53.400 65.400 61.200 66.300 ;
        RECT 62.400 65.400 64.200 77.400 ;
        RECT 83.400 71.400 85.200 77.400 ;
        RECT 104.400 71.400 106.200 77.400 ;
        RECT 125.400 71.400 127.200 77.400 ;
        RECT 20.100 58.050 21.900 59.850 ;
        RECT 32.100 58.050 33.900 59.850 ;
        RECT 35.700 58.050 36.600 65.400 ;
        RECT 38.100 58.050 39.900 59.850 ;
        RECT 56.100 58.050 57.900 59.850 ;
        RECT 62.700 58.050 63.600 65.400 ;
        RECT 83.850 58.050 85.050 71.400 ;
        RECT 89.100 58.050 90.900 59.850 ;
        RECT 104.400 58.050 105.600 71.400 ;
        RECT 125.400 58.050 126.600 71.400 ;
        RECT 134.550 65.400 136.350 77.400 ;
        RECT 142.050 71.400 143.850 77.400 ;
        RECT 139.950 69.300 143.850 71.400 ;
        RECT 149.850 70.500 151.650 77.400 ;
        RECT 157.650 71.400 159.450 77.400 ;
        RECT 158.250 70.500 159.450 71.400 ;
        RECT 148.950 69.450 155.550 70.500 ;
        RECT 148.950 68.700 150.750 69.450 ;
        RECT 153.750 68.700 155.550 69.450 ;
        RECT 158.250 68.400 163.050 70.500 ;
        RECT 141.150 66.600 143.850 68.400 ;
        RECT 144.750 67.800 146.550 68.400 ;
        RECT 144.750 66.900 151.050 67.800 ;
        RECT 158.250 67.500 159.450 68.400 ;
        RECT 144.750 66.600 146.550 66.900 ;
        RECT 142.950 65.700 143.850 66.600 ;
        RECT 134.550 58.050 135.750 65.400 ;
        RECT 139.950 64.800 142.050 65.700 ;
        RECT 142.950 64.800 148.050 65.700 ;
        RECT 137.850 63.600 142.050 64.800 ;
        RECT 136.950 61.800 138.750 63.600 ;
        RECT 13.950 55.950 16.050 58.050 ;
        RECT 16.950 55.950 19.050 58.050 ;
        RECT 19.950 55.950 22.050 58.050 ;
        RECT 31.950 55.950 34.050 58.050 ;
        RECT 34.950 55.950 37.050 58.050 ;
        RECT 37.950 55.950 40.050 58.050 ;
        RECT 52.950 55.950 55.050 58.050 ;
        RECT 55.950 55.950 58.050 58.050 ;
        RECT 58.950 55.950 61.050 58.050 ;
        RECT 61.950 55.950 64.050 58.050 ;
        RECT 79.950 55.950 82.050 58.050 ;
        RECT 82.950 55.950 85.050 58.050 ;
        RECT 85.950 55.950 88.050 58.050 ;
        RECT 88.950 55.950 91.050 58.050 ;
        RECT 100.950 55.950 103.050 58.050 ;
        RECT 103.950 55.950 106.050 58.050 ;
        RECT 106.950 55.950 109.050 58.050 ;
        RECT 121.950 55.950 124.050 58.050 ;
        RECT 124.950 55.950 127.050 58.050 ;
        RECT 127.950 55.950 130.050 58.050 ;
        RECT 134.550 57.750 139.050 58.050 ;
        RECT 134.550 55.950 140.850 57.750 ;
        RECT 17.400 45.600 18.300 55.950 ;
        RECT 35.700 45.600 36.600 55.950 ;
        RECT 53.100 54.150 54.900 55.950 ;
        RECT 59.100 54.150 60.900 55.950 ;
        RECT 62.700 48.600 63.600 55.950 ;
        RECT 80.100 54.150 81.900 55.950 ;
        RECT 82.950 51.750 84.150 55.950 ;
        RECT 86.100 54.150 87.900 55.950 ;
        RECT 101.100 54.150 102.900 55.950 ;
        RECT 80.400 50.700 84.150 51.750 ;
        RECT 104.400 50.700 105.600 55.950 ;
        RECT 107.100 54.150 108.900 55.950 ;
        RECT 122.100 54.150 123.900 55.950 ;
        RECT 125.400 50.700 126.600 55.950 ;
        RECT 128.100 54.150 129.900 55.950 ;
        RECT 80.400 48.600 81.600 50.700 ;
        RECT 104.400 49.800 108.600 50.700 ;
        RECT 125.400 49.800 129.600 50.700 ;
        RECT 58.500 47.400 63.600 48.600 ;
        RECT 16.800 42.600 18.600 45.600 ;
        RECT 35.400 42.600 37.200 45.600 ;
        RECT 58.500 42.600 60.300 47.400 ;
        RECT 79.800 42.600 81.600 48.600 ;
        RECT 82.800 47.700 90.600 49.050 ;
        RECT 82.800 42.600 84.600 47.700 ;
        RECT 88.800 42.600 90.600 47.700 ;
        RECT 106.800 42.600 108.600 49.800 ;
        RECT 127.800 42.600 129.600 49.800 ;
        RECT 134.550 48.600 135.750 55.950 ;
        RECT 147.150 52.200 148.050 64.800 ;
        RECT 150.150 64.800 151.050 66.900 ;
        RECT 151.950 66.300 159.450 67.500 ;
        RECT 151.950 65.700 153.750 66.300 ;
        RECT 166.050 65.400 167.850 77.400 ;
        RECT 184.500 66.600 186.300 77.400 ;
        RECT 150.150 64.500 158.550 64.800 ;
        RECT 166.950 64.500 167.850 65.400 ;
        RECT 150.150 63.900 167.850 64.500 ;
        RECT 156.750 63.300 167.850 63.900 ;
        RECT 156.750 63.000 158.550 63.300 ;
        RECT 154.950 56.400 157.050 58.050 ;
        RECT 154.950 55.200 162.900 56.400 ;
        RECT 163.950 55.950 166.050 58.050 ;
        RECT 161.100 54.600 162.900 55.200 ;
        RECT 164.100 54.150 165.900 55.950 ;
        RECT 158.100 53.400 159.900 54.000 ;
        RECT 164.100 53.400 165.000 54.150 ;
        RECT 158.100 52.200 165.000 53.400 ;
        RECT 147.150 51.000 159.150 52.200 ;
        RECT 147.150 50.400 148.950 51.000 ;
        RECT 158.100 49.200 159.150 51.000 ;
        RECT 134.550 42.600 136.350 48.600 ;
        RECT 139.950 47.700 142.050 48.600 ;
        RECT 139.950 46.500 143.700 47.700 ;
        RECT 154.350 47.550 156.150 48.300 ;
        RECT 142.650 45.600 143.700 46.500 ;
        RECT 151.200 46.500 156.150 47.550 ;
        RECT 157.650 47.400 159.450 49.200 ;
        RECT 166.950 48.600 167.850 63.300 ;
        RECT 182.700 65.400 186.300 66.600 ;
        RECT 202.800 65.400 204.600 77.400 ;
        RECT 205.800 66.300 207.600 77.400 ;
        RECT 211.800 66.300 213.600 77.400 ;
        RECT 229.800 71.400 231.600 77.400 ;
        RECT 205.800 65.400 213.600 66.300 ;
        RECT 179.100 58.050 180.900 59.850 ;
        RECT 182.700 58.050 183.600 65.400 ;
        RECT 185.100 58.050 186.900 59.850 ;
        RECT 203.400 58.050 204.300 65.400 ;
        RECT 209.100 58.050 210.900 59.850 ;
        RECT 224.100 58.050 225.900 59.850 ;
        RECT 229.950 58.050 231.150 71.400 ;
        RECT 239.550 65.400 241.350 77.400 ;
        RECT 247.050 71.400 248.850 77.400 ;
        RECT 244.950 69.300 248.850 71.400 ;
        RECT 254.850 70.500 256.650 77.400 ;
        RECT 262.650 71.400 264.450 77.400 ;
        RECT 263.250 70.500 264.450 71.400 ;
        RECT 253.950 69.450 260.550 70.500 ;
        RECT 253.950 68.700 255.750 69.450 ;
        RECT 258.750 68.700 260.550 69.450 ;
        RECT 263.250 68.400 268.050 70.500 ;
        RECT 246.150 66.600 248.850 68.400 ;
        RECT 249.750 67.800 251.550 68.400 ;
        RECT 249.750 66.900 256.050 67.800 ;
        RECT 263.250 67.500 264.450 68.400 ;
        RECT 249.750 66.600 251.550 66.900 ;
        RECT 247.950 65.700 248.850 66.600 ;
        RECT 239.550 58.050 240.750 65.400 ;
        RECT 244.950 64.800 247.050 65.700 ;
        RECT 247.950 64.800 253.050 65.700 ;
        RECT 242.850 63.600 247.050 64.800 ;
        RECT 241.950 61.800 243.750 63.600 ;
        RECT 178.950 55.950 181.050 58.050 ;
        RECT 181.950 55.950 184.050 58.050 ;
        RECT 184.950 55.950 187.050 58.050 ;
        RECT 202.950 55.950 205.050 58.050 ;
        RECT 205.950 55.950 208.050 58.050 ;
        RECT 208.950 55.950 211.050 58.050 ;
        RECT 211.950 55.950 214.050 58.050 ;
        RECT 223.950 55.950 226.050 58.050 ;
        RECT 226.950 55.950 229.050 58.050 ;
        RECT 229.950 55.950 232.050 58.050 ;
        RECT 232.950 55.950 235.050 58.050 ;
        RECT 239.550 57.750 244.050 58.050 ;
        RECT 239.550 55.950 245.850 57.750 ;
        RECT 160.950 46.500 163.050 48.600 ;
        RECT 151.200 45.600 152.250 46.500 ;
        RECT 160.950 45.600 162.000 46.500 ;
        RECT 142.650 42.600 144.450 45.600 ;
        RECT 150.450 42.600 152.250 45.600 ;
        RECT 158.250 44.700 162.000 45.600 ;
        RECT 158.250 42.600 160.050 44.700 ;
        RECT 166.050 42.600 167.850 48.600 ;
        RECT 182.700 45.600 183.600 55.950 ;
        RECT 203.400 48.600 204.300 55.950 ;
        RECT 206.100 54.150 207.900 55.950 ;
        RECT 212.100 54.150 213.900 55.950 ;
        RECT 227.100 54.150 228.900 55.950 ;
        RECT 230.850 51.750 232.050 55.950 ;
        RECT 233.100 54.150 234.900 55.950 ;
        RECT 230.850 50.700 234.600 51.750 ;
        RECT 203.400 47.400 208.500 48.600 ;
        RECT 182.400 42.600 184.200 45.600 ;
        RECT 206.700 42.600 208.500 47.400 ;
        RECT 224.400 47.700 232.200 49.050 ;
        RECT 224.400 42.600 226.200 47.700 ;
        RECT 230.400 42.600 232.200 47.700 ;
        RECT 233.400 48.600 234.600 50.700 ;
        RECT 239.550 48.600 240.750 55.950 ;
        RECT 252.150 52.200 253.050 64.800 ;
        RECT 255.150 64.800 256.050 66.900 ;
        RECT 256.950 66.300 264.450 67.500 ;
        RECT 256.950 65.700 258.750 66.300 ;
        RECT 271.050 65.400 272.850 77.400 ;
        RECT 255.150 64.500 263.550 64.800 ;
        RECT 271.950 64.500 272.850 65.400 ;
        RECT 255.150 63.900 272.850 64.500 ;
        RECT 261.750 63.300 272.850 63.900 ;
        RECT 261.750 63.000 263.550 63.300 ;
        RECT 259.950 56.400 262.050 58.050 ;
        RECT 259.950 55.200 267.900 56.400 ;
        RECT 268.950 55.950 271.050 58.050 ;
        RECT 266.100 54.600 267.900 55.200 ;
        RECT 269.100 54.150 270.900 55.950 ;
        RECT 263.100 53.400 264.900 54.000 ;
        RECT 269.100 53.400 270.000 54.150 ;
        RECT 263.100 52.200 270.000 53.400 ;
        RECT 252.150 51.000 264.150 52.200 ;
        RECT 252.150 50.400 253.950 51.000 ;
        RECT 263.100 49.200 264.150 51.000 ;
        RECT 233.400 42.600 235.200 48.600 ;
        RECT 239.550 42.600 241.350 48.600 ;
        RECT 244.950 47.700 247.050 48.600 ;
        RECT 244.950 46.500 248.700 47.700 ;
        RECT 259.350 47.550 261.150 48.300 ;
        RECT 247.650 45.600 248.700 46.500 ;
        RECT 256.200 46.500 261.150 47.550 ;
        RECT 262.650 47.400 264.450 49.200 ;
        RECT 271.950 48.600 272.850 63.300 ;
        RECT 287.400 71.400 289.200 77.400 ;
        RECT 307.800 71.400 309.600 77.400 ;
        RECT 325.800 71.400 327.600 77.400 ;
        RECT 284.100 58.050 285.900 59.850 ;
        RECT 287.400 58.050 288.600 71.400 ;
        RECT 308.400 58.050 309.600 71.400 ;
        RECT 326.700 71.100 327.600 71.400 ;
        RECT 331.800 71.400 333.600 77.400 ;
        RECT 331.800 71.100 333.300 71.400 ;
        RECT 326.700 70.200 333.300 71.100 ;
        RECT 326.700 58.050 327.600 70.200 ;
        RECT 352.500 66.600 354.300 77.400 ;
        RECT 374.400 71.400 376.200 77.400 ;
        RECT 394.800 71.400 396.600 77.400 ;
        RECT 415.800 71.400 417.600 77.400 ;
        RECT 437.400 71.400 439.200 77.400 ;
        RECT 457.800 71.400 459.600 77.400 ;
        RECT 478.800 71.400 480.600 77.400 ;
        RECT 350.700 65.400 354.300 66.600 ;
        RECT 332.100 58.050 333.900 59.850 ;
        RECT 347.100 58.050 348.900 59.850 ;
        RECT 350.700 58.050 351.600 65.400 ;
        RECT 353.100 58.050 354.900 59.850 ;
        RECT 374.850 58.050 376.050 71.400 ;
        RECT 385.950 60.450 388.050 61.050 ;
        RECT 391.950 60.450 394.050 61.050 ;
        RECT 380.100 58.050 381.900 59.850 ;
        RECT 385.950 59.550 394.050 60.450 ;
        RECT 385.950 58.950 388.050 59.550 ;
        RECT 391.950 58.950 394.050 59.550 ;
        RECT 395.400 58.050 396.600 71.400 ;
        RECT 398.100 58.050 399.900 59.850 ;
        RECT 410.100 58.050 411.900 59.850 ;
        RECT 415.950 58.050 417.150 71.400 ;
        RECT 434.100 58.050 435.900 59.850 ;
        RECT 437.400 58.050 438.600 71.400 ;
        RECT 452.100 58.050 453.900 59.850 ;
        RECT 457.950 58.050 459.150 71.400 ;
        RECT 479.400 58.050 480.600 71.400 ;
        RECT 496.800 65.400 498.600 77.400 ;
        RECT 499.800 66.300 501.600 77.400 ;
        RECT 505.800 66.300 507.600 77.400 ;
        RECT 523.800 71.400 525.600 77.400 ;
        RECT 541.800 71.400 543.600 77.400 ;
        RECT 499.800 65.400 507.600 66.300 ;
        RECT 482.100 58.050 483.900 59.850 ;
        RECT 497.400 58.050 498.300 65.400 ;
        RECT 503.100 58.050 504.900 59.850 ;
        RECT 524.400 58.050 525.600 71.400 ;
        RECT 527.100 58.050 528.900 59.850 ;
        RECT 542.400 58.050 543.600 71.400 ;
        RECT 559.800 65.400 561.600 77.400 ;
        RECT 562.800 66.300 564.600 77.400 ;
        RECT 568.800 66.300 570.600 77.400 ;
        RECT 562.800 65.400 570.600 66.300 ;
        RECT 584.700 66.600 586.500 77.400 ;
        RECT 605.700 66.600 607.500 77.400 ;
        RECT 625.800 71.400 627.600 77.400 ;
        RECT 584.700 65.400 588.300 66.600 ;
        RECT 605.700 65.400 609.300 66.600 ;
        RECT 545.100 58.050 546.900 59.850 ;
        RECT 560.400 58.050 561.300 65.400 ;
        RECT 562.950 63.450 565.050 64.050 ;
        RECT 580.950 63.450 583.050 64.050 ;
        RECT 562.950 62.550 583.050 63.450 ;
        RECT 562.950 61.950 565.050 62.550 ;
        RECT 580.950 61.950 583.050 62.550 ;
        RECT 566.100 58.050 567.900 59.850 ;
        RECT 584.100 58.050 585.900 59.850 ;
        RECT 587.400 58.050 588.300 65.400 ;
        RECT 590.100 58.050 591.900 59.850 ;
        RECT 605.100 58.050 606.900 59.850 ;
        RECT 608.400 58.050 609.300 65.400 ;
        RECT 611.100 58.050 612.900 59.850 ;
        RECT 626.400 58.050 627.600 71.400 ;
        RECT 646.500 66.600 648.300 77.400 ;
        RECT 664.800 71.400 666.600 77.400 ;
        RECT 644.700 65.400 648.300 66.600 ;
        RECT 665.700 71.100 666.600 71.400 ;
        RECT 670.800 71.400 672.600 77.400 ;
        RECT 688.800 71.400 690.600 77.400 ;
        RECT 670.800 71.100 672.300 71.400 ;
        RECT 665.700 70.200 672.300 71.100 ;
        RECT 689.700 71.100 690.600 71.400 ;
        RECT 694.800 71.400 696.600 77.400 ;
        RECT 713.400 71.400 715.200 77.400 ;
        RECT 731.400 71.400 733.200 77.400 ;
        RECT 694.800 71.100 696.300 71.400 ;
        RECT 689.700 70.200 696.300 71.100 ;
        RECT 629.100 58.050 630.900 59.850 ;
        RECT 641.100 58.050 642.900 59.850 ;
        RECT 644.700 58.050 645.600 65.400 ;
        RECT 647.100 58.050 648.900 59.850 ;
        RECT 665.700 58.050 666.600 70.200 ;
        RECT 671.100 58.050 672.900 59.850 ;
        RECT 689.700 58.050 690.600 70.200 ;
        RECT 697.950 63.450 700.050 64.050 ;
        RECT 703.950 63.450 706.050 64.050 ;
        RECT 697.950 62.550 706.050 63.450 ;
        RECT 697.950 61.950 700.050 62.550 ;
        RECT 703.950 61.950 706.050 62.550 ;
        RECT 695.100 58.050 696.900 59.850 ;
        RECT 710.100 58.050 711.900 59.850 ;
        RECT 713.400 58.050 714.600 71.400 ;
        RECT 731.700 71.100 733.200 71.400 ;
        RECT 737.400 71.400 739.200 77.400 ;
        RECT 757.800 71.400 759.600 77.400 ;
        RECT 776.400 71.400 778.200 77.400 ;
        RECT 737.400 71.100 738.300 71.400 ;
        RECT 731.700 70.200 738.300 71.100 ;
        RECT 731.100 58.050 732.900 59.850 ;
        RECT 737.400 58.050 738.300 70.200 ;
        RECT 758.400 58.050 759.600 71.400 ;
        RECT 776.700 71.100 778.200 71.400 ;
        RECT 782.400 71.400 784.200 77.400 ;
        RECT 800.400 71.400 802.200 77.400 ;
        RECT 818.400 71.400 820.200 77.400 ;
        RECT 833.400 71.400 835.200 77.400 ;
        RECT 782.400 71.100 783.300 71.400 ;
        RECT 776.700 70.200 783.300 71.100 ;
        RECT 776.100 58.050 777.900 59.850 ;
        RECT 782.400 58.050 783.300 70.200 ;
        RECT 797.100 58.050 798.900 59.850 ;
        RECT 800.400 58.050 801.600 71.400 ;
        RECT 815.100 58.050 816.900 59.850 ;
        RECT 818.400 58.050 819.600 71.400 ;
        RECT 833.400 64.500 834.600 71.400 ;
        RECT 839.400 65.400 841.200 77.400 ;
        RECT 857.400 71.400 859.200 77.400 ;
        RECT 857.700 71.100 859.200 71.400 ;
        RECT 863.400 71.400 865.200 77.400 ;
        RECT 881.400 71.400 883.200 77.400 ;
        RECT 863.400 71.100 864.300 71.400 ;
        RECT 857.700 70.200 864.300 71.100 ;
        RECT 833.400 63.600 839.100 64.500 ;
        RECT 837.150 62.700 839.100 63.600 ;
        RECT 833.100 58.050 834.900 59.850 ;
        RECT 283.950 55.950 286.050 58.050 ;
        RECT 286.950 55.950 289.050 58.050 ;
        RECT 304.950 55.950 307.050 58.050 ;
        RECT 307.950 55.950 310.050 58.050 ;
        RECT 310.950 55.950 313.050 58.050 ;
        RECT 325.950 55.950 328.050 58.050 ;
        RECT 328.950 55.950 331.050 58.050 ;
        RECT 331.950 55.950 334.050 58.050 ;
        RECT 334.950 55.950 337.050 58.050 ;
        RECT 346.950 55.950 349.050 58.050 ;
        RECT 349.950 55.950 352.050 58.050 ;
        RECT 352.950 55.950 355.050 58.050 ;
        RECT 370.950 55.950 373.050 58.050 ;
        RECT 373.950 55.950 376.050 58.050 ;
        RECT 376.950 55.950 379.050 58.050 ;
        RECT 379.950 55.950 382.050 58.050 ;
        RECT 394.950 55.950 397.050 58.050 ;
        RECT 397.950 55.950 400.050 58.050 ;
        RECT 409.950 55.950 412.050 58.050 ;
        RECT 412.950 55.950 415.050 58.050 ;
        RECT 415.950 55.950 418.050 58.050 ;
        RECT 418.950 55.950 421.050 58.050 ;
        RECT 433.950 55.950 436.050 58.050 ;
        RECT 436.950 55.950 439.050 58.050 ;
        RECT 451.950 55.950 454.050 58.050 ;
        RECT 454.950 55.950 457.050 58.050 ;
        RECT 457.950 55.950 460.050 58.050 ;
        RECT 460.950 55.950 463.050 58.050 ;
        RECT 478.950 55.950 481.050 58.050 ;
        RECT 481.950 55.950 484.050 58.050 ;
        RECT 496.950 55.950 499.050 58.050 ;
        RECT 499.950 55.950 502.050 58.050 ;
        RECT 502.950 55.950 505.050 58.050 ;
        RECT 505.950 55.950 508.050 58.050 ;
        RECT 523.950 55.950 526.050 58.050 ;
        RECT 526.950 55.950 529.050 58.050 ;
        RECT 541.950 55.950 544.050 58.050 ;
        RECT 544.950 55.950 547.050 58.050 ;
        RECT 559.950 55.950 562.050 58.050 ;
        RECT 562.950 55.950 565.050 58.050 ;
        RECT 565.950 55.950 568.050 58.050 ;
        RECT 568.950 55.950 571.050 58.050 ;
        RECT 583.950 55.950 586.050 58.050 ;
        RECT 586.950 55.950 589.050 58.050 ;
        RECT 589.950 55.950 592.050 58.050 ;
        RECT 604.950 55.950 607.050 58.050 ;
        RECT 607.950 55.950 610.050 58.050 ;
        RECT 610.950 55.950 613.050 58.050 ;
        RECT 625.950 55.950 628.050 58.050 ;
        RECT 628.950 55.950 631.050 58.050 ;
        RECT 640.950 55.950 643.050 58.050 ;
        RECT 643.950 55.950 646.050 58.050 ;
        RECT 646.950 55.950 649.050 58.050 ;
        RECT 664.950 55.950 667.050 58.050 ;
        RECT 667.950 55.950 670.050 58.050 ;
        RECT 670.950 55.950 673.050 58.050 ;
        RECT 673.950 55.950 676.050 58.050 ;
        RECT 688.950 55.950 691.050 58.050 ;
        RECT 691.950 55.950 694.050 58.050 ;
        RECT 694.950 55.950 697.050 58.050 ;
        RECT 697.950 55.950 700.050 58.050 ;
        RECT 709.950 55.950 712.050 58.050 ;
        RECT 712.950 55.950 715.050 58.050 ;
        RECT 727.950 55.950 730.050 58.050 ;
        RECT 730.950 55.950 733.050 58.050 ;
        RECT 733.950 55.950 736.050 58.050 ;
        RECT 736.950 55.950 739.050 58.050 ;
        RECT 754.950 55.950 757.050 58.050 ;
        RECT 757.950 55.950 760.050 58.050 ;
        RECT 760.950 55.950 763.050 58.050 ;
        RECT 772.950 55.950 775.050 58.050 ;
        RECT 775.950 55.950 778.050 58.050 ;
        RECT 778.950 55.950 781.050 58.050 ;
        RECT 781.950 55.950 784.050 58.050 ;
        RECT 796.950 55.950 799.050 58.050 ;
        RECT 799.950 55.950 802.050 58.050 ;
        RECT 814.950 55.950 817.050 58.050 ;
        RECT 817.950 55.950 820.050 58.050 ;
        RECT 832.950 55.950 835.050 58.050 ;
        RECT 265.950 46.500 268.050 48.600 ;
        RECT 256.200 45.600 257.250 46.500 ;
        RECT 265.950 45.600 267.000 46.500 ;
        RECT 247.650 42.600 249.450 45.600 ;
        RECT 255.450 42.600 257.250 45.600 ;
        RECT 263.250 44.700 267.000 45.600 ;
        RECT 263.250 42.600 265.050 44.700 ;
        RECT 271.050 42.600 272.850 48.600 ;
        RECT 287.400 45.600 288.600 55.950 ;
        RECT 305.100 54.150 306.900 55.950 ;
        RECT 308.400 50.700 309.600 55.950 ;
        RECT 311.100 54.150 312.900 55.950 ;
        RECT 326.700 52.200 327.600 55.950 ;
        RECT 329.100 54.150 330.900 55.950 ;
        RECT 335.100 54.150 336.900 55.950 ;
        RECT 326.700 51.000 330.000 52.200 ;
        RECT 305.400 49.800 309.600 50.700 ;
        RECT 287.400 42.600 289.200 45.600 ;
        RECT 305.400 42.600 307.200 49.800 ;
        RECT 328.200 42.600 330.000 51.000 ;
        RECT 350.700 45.600 351.600 55.950 ;
        RECT 371.100 54.150 372.900 55.950 ;
        RECT 373.950 51.750 375.150 55.950 ;
        RECT 377.100 54.150 378.900 55.950 ;
        RECT 371.400 50.700 375.150 51.750 ;
        RECT 371.400 48.600 372.600 50.700 ;
        RECT 350.400 42.600 352.200 45.600 ;
        RECT 370.800 42.600 372.600 48.600 ;
        RECT 373.800 47.700 381.600 49.050 ;
        RECT 373.800 42.600 375.600 47.700 ;
        RECT 379.800 42.600 381.600 47.700 ;
        RECT 395.400 45.600 396.600 55.950 ;
        RECT 413.100 54.150 414.900 55.950 ;
        RECT 416.850 51.750 418.050 55.950 ;
        RECT 419.100 54.150 420.900 55.950 ;
        RECT 416.850 50.700 420.600 51.750 ;
        RECT 394.800 42.600 396.600 45.600 ;
        RECT 410.400 47.700 418.200 49.050 ;
        RECT 410.400 42.600 412.200 47.700 ;
        RECT 416.400 42.600 418.200 47.700 ;
        RECT 419.400 48.600 420.600 50.700 ;
        RECT 419.400 42.600 421.200 48.600 ;
        RECT 437.400 45.600 438.600 55.950 ;
        RECT 455.100 54.150 456.900 55.950 ;
        RECT 458.850 51.750 460.050 55.950 ;
        RECT 461.100 54.150 462.900 55.950 ;
        RECT 458.850 50.700 462.600 51.750 ;
        RECT 452.400 47.700 460.200 49.050 ;
        RECT 437.400 42.600 439.200 45.600 ;
        RECT 452.400 42.600 454.200 47.700 ;
        RECT 458.400 42.600 460.200 47.700 ;
        RECT 461.400 48.600 462.600 50.700 ;
        RECT 461.400 42.600 463.200 48.600 ;
        RECT 479.400 45.600 480.600 55.950 ;
        RECT 497.400 48.600 498.300 55.950 ;
        RECT 500.100 54.150 501.900 55.950 ;
        RECT 506.100 54.150 507.900 55.950 ;
        RECT 497.400 47.400 502.500 48.600 ;
        RECT 478.800 42.600 480.600 45.600 ;
        RECT 500.700 42.600 502.500 47.400 ;
        RECT 524.400 45.600 525.600 55.950 ;
        RECT 542.400 45.600 543.600 55.950 ;
        RECT 560.400 48.600 561.300 55.950 ;
        RECT 563.100 54.150 564.900 55.950 ;
        RECT 569.100 54.150 570.900 55.950 ;
        RECT 560.400 47.400 565.500 48.600 ;
        RECT 523.800 42.600 525.600 45.600 ;
        RECT 541.800 42.600 543.600 45.600 ;
        RECT 563.700 42.600 565.500 47.400 ;
        RECT 587.400 45.600 588.300 55.950 ;
        RECT 608.400 45.600 609.300 55.950 ;
        RECT 626.400 45.600 627.600 55.950 ;
        RECT 644.700 45.600 645.600 55.950 ;
        RECT 665.700 52.200 666.600 55.950 ;
        RECT 668.100 54.150 669.900 55.950 ;
        RECT 674.100 54.150 675.900 55.950 ;
        RECT 689.700 52.200 690.600 55.950 ;
        RECT 692.100 54.150 693.900 55.950 ;
        RECT 698.100 54.150 699.900 55.950 ;
        RECT 665.700 51.000 669.000 52.200 ;
        RECT 689.700 51.000 693.000 52.200 ;
        RECT 586.800 42.600 588.600 45.600 ;
        RECT 607.800 42.600 609.600 45.600 ;
        RECT 625.800 42.600 627.600 45.600 ;
        RECT 644.400 42.600 646.200 45.600 ;
        RECT 667.200 42.600 669.000 51.000 ;
        RECT 691.200 42.600 693.000 51.000 ;
        RECT 713.400 45.600 714.600 55.950 ;
        RECT 728.100 54.150 729.900 55.950 ;
        RECT 734.100 54.150 735.900 55.950 ;
        RECT 737.400 52.200 738.300 55.950 ;
        RECT 755.100 54.150 756.900 55.950 ;
        RECT 735.000 51.000 738.300 52.200 ;
        RECT 713.400 42.600 715.200 45.600 ;
        RECT 735.000 42.600 736.800 51.000 ;
        RECT 758.400 50.700 759.600 55.950 ;
        RECT 761.100 54.150 762.900 55.950 ;
        RECT 773.100 54.150 774.900 55.950 ;
        RECT 779.100 54.150 780.900 55.950 ;
        RECT 782.400 52.200 783.300 55.950 ;
        RECT 793.950 54.450 796.050 55.050 ;
        RECT 785.550 54.000 796.050 54.450 ;
        RECT 755.400 49.800 759.600 50.700 ;
        RECT 780.000 51.000 783.300 52.200 ;
        RECT 784.950 53.550 796.050 54.000 ;
        RECT 755.400 42.600 757.200 49.800 ;
        RECT 780.000 42.600 781.800 51.000 ;
        RECT 784.950 49.950 787.050 53.550 ;
        RECT 793.950 52.950 796.050 53.550 ;
        RECT 800.400 45.600 801.600 55.950 ;
        RECT 818.400 45.600 819.600 55.950 ;
        RECT 837.150 51.300 838.050 62.700 ;
        RECT 840.000 58.050 841.200 65.400 ;
        RECT 847.950 63.450 850.050 64.050 ;
        RECT 856.950 63.450 859.050 64.050 ;
        RECT 847.950 62.550 859.050 63.450 ;
        RECT 847.950 61.950 850.050 62.550 ;
        RECT 856.950 61.950 859.050 62.550 ;
        RECT 857.100 58.050 858.900 59.850 ;
        RECT 863.400 58.050 864.300 70.200 ;
        RECT 865.950 60.450 870.000 61.050 ;
        RECT 865.950 58.950 870.450 60.450 ;
        RECT 838.950 55.950 841.200 58.050 ;
        RECT 853.950 55.950 856.050 58.050 ;
        RECT 856.950 55.950 859.050 58.050 ;
        RECT 859.950 55.950 862.050 58.050 ;
        RECT 862.950 55.950 865.050 58.050 ;
        RECT 837.150 50.400 839.100 51.300 ;
        RECT 833.400 49.500 839.100 50.400 ;
        RECT 833.400 45.600 834.600 49.500 ;
        RECT 840.000 48.600 841.200 55.950 ;
        RECT 854.100 54.150 855.900 55.950 ;
        RECT 860.100 54.150 861.900 55.950 ;
        RECT 863.400 52.200 864.300 55.950 ;
        RECT 869.550 55.050 870.450 58.950 ;
        RECT 878.100 58.050 879.900 59.850 ;
        RECT 881.400 58.050 882.600 71.400 ;
        RECT 877.950 55.950 880.050 58.050 ;
        RECT 880.950 55.950 883.050 58.050 ;
        RECT 865.950 53.550 870.450 55.050 ;
        RECT 865.950 52.950 870.000 53.550 ;
        RECT 800.400 42.600 802.200 45.600 ;
        RECT 818.400 42.600 820.200 45.600 ;
        RECT 833.400 42.600 835.200 45.600 ;
        RECT 839.400 42.600 841.200 48.600 ;
        RECT 861.000 51.000 864.300 52.200 ;
        RECT 861.000 42.600 862.800 51.000 ;
        RECT 881.400 45.600 882.600 55.950 ;
        RECT 881.400 42.600 883.200 45.600 ;
        RECT 13.800 35.400 15.600 38.400 ;
        RECT 14.400 25.050 15.600 35.400 ;
        RECT 34.800 31.200 36.600 38.400 ;
        RECT 32.400 30.300 36.600 31.200 ;
        RECT 52.800 32.400 54.600 38.400 ;
        RECT 58.800 35.400 60.600 38.400 ;
        RECT 29.100 25.050 30.900 26.850 ;
        RECT 32.400 25.050 33.600 30.300 ;
        RECT 35.100 25.050 36.900 26.850 ;
        RECT 52.800 25.050 54.000 32.400 ;
        RECT 59.400 31.500 60.600 35.400 ;
        RECT 54.900 30.600 60.600 31.500 ;
        RECT 73.800 32.400 75.600 38.400 ;
        RECT 79.800 35.400 81.600 38.400 ;
        RECT 54.900 29.700 56.850 30.600 ;
        RECT 13.950 22.950 16.050 25.050 ;
        RECT 16.950 22.950 19.050 25.050 ;
        RECT 28.950 22.950 31.050 25.050 ;
        RECT 31.950 22.950 34.050 25.050 ;
        RECT 34.950 22.950 37.050 25.050 ;
        RECT 52.800 22.950 55.050 25.050 ;
        RECT 14.400 9.600 15.600 22.950 ;
        RECT 17.100 21.150 18.900 22.950 ;
        RECT 13.800 3.600 15.600 9.600 ;
        RECT 32.400 9.600 33.600 22.950 ;
        RECT 52.800 15.600 54.000 22.950 ;
        RECT 55.950 18.300 56.850 29.700 ;
        RECT 73.800 25.050 75.000 32.400 ;
        RECT 80.400 31.500 81.600 35.400 ;
        RECT 75.900 30.600 81.600 31.500 ;
        RECT 83.550 32.400 85.350 38.400 ;
        RECT 91.650 35.400 93.450 38.400 ;
        RECT 99.450 35.400 101.250 38.400 ;
        RECT 107.250 36.300 109.050 38.400 ;
        RECT 107.250 35.400 111.000 36.300 ;
        RECT 91.650 34.500 92.700 35.400 ;
        RECT 88.950 33.300 92.700 34.500 ;
        RECT 100.200 34.500 101.250 35.400 ;
        RECT 109.950 34.500 111.000 35.400 ;
        RECT 100.200 33.450 105.150 34.500 ;
        RECT 88.950 32.400 91.050 33.300 ;
        RECT 103.350 32.700 105.150 33.450 ;
        RECT 75.900 29.700 77.850 30.600 ;
        RECT 58.950 22.950 61.050 25.050 ;
        RECT 73.800 22.950 76.050 25.050 ;
        RECT 59.100 21.150 60.900 22.950 ;
        RECT 54.900 17.400 56.850 18.300 ;
        RECT 54.900 16.500 60.600 17.400 ;
        RECT 32.400 3.600 34.200 9.600 ;
        RECT 52.800 3.600 54.600 15.600 ;
        RECT 59.400 9.600 60.600 16.500 ;
        RECT 58.800 3.600 60.600 9.600 ;
        RECT 73.800 15.600 75.000 22.950 ;
        RECT 76.950 18.300 77.850 29.700 ;
        RECT 83.550 25.050 84.750 32.400 ;
        RECT 106.650 31.800 108.450 33.600 ;
        RECT 109.950 32.400 112.050 34.500 ;
        RECT 115.050 32.400 116.850 38.400 ;
        RECT 96.150 30.000 97.950 30.600 ;
        RECT 107.100 30.000 108.150 31.800 ;
        RECT 96.150 28.800 108.150 30.000 ;
        RECT 79.950 22.950 82.050 25.050 ;
        RECT 83.550 23.250 89.850 25.050 ;
        RECT 83.550 22.950 88.050 23.250 ;
        RECT 80.100 21.150 81.900 22.950 ;
        RECT 75.900 17.400 77.850 18.300 ;
        RECT 75.900 16.500 81.600 17.400 ;
        RECT 73.800 3.600 75.600 15.600 ;
        RECT 80.400 9.600 81.600 16.500 ;
        RECT 79.800 3.600 81.600 9.600 ;
        RECT 83.550 15.600 84.750 22.950 ;
        RECT 85.950 17.400 87.750 19.200 ;
        RECT 86.850 16.200 91.050 17.400 ;
        RECT 96.150 16.200 97.050 28.800 ;
        RECT 107.100 27.600 114.000 28.800 ;
        RECT 107.100 27.000 108.900 27.600 ;
        RECT 113.100 26.850 114.000 27.600 ;
        RECT 110.100 25.800 111.900 26.400 ;
        RECT 103.950 24.600 111.900 25.800 ;
        RECT 113.100 25.050 114.900 26.850 ;
        RECT 103.950 22.950 106.050 24.600 ;
        RECT 112.950 22.950 115.050 25.050 ;
        RECT 105.750 17.700 107.550 18.000 ;
        RECT 115.950 17.700 116.850 32.400 ;
        RECT 134.400 35.400 136.200 38.400 ;
        RECT 134.400 25.050 135.600 35.400 ;
        RECT 149.400 33.300 151.200 38.400 ;
        RECT 155.400 33.300 157.200 38.400 ;
        RECT 149.400 31.950 157.200 33.300 ;
        RECT 158.400 32.400 160.200 38.400 ;
        RECT 158.400 30.300 159.600 32.400 ;
        RECT 178.800 31.200 180.600 38.400 ;
        RECT 155.850 29.250 159.600 30.300 ;
        RECT 163.950 30.450 166.050 31.050 ;
        RECT 172.950 30.450 175.050 31.050 ;
        RECT 163.950 29.550 175.050 30.450 ;
        RECT 152.100 25.050 153.900 26.850 ;
        RECT 155.850 25.050 157.050 29.250 ;
        RECT 163.950 28.950 166.050 29.550 ;
        RECT 172.950 28.950 175.050 29.550 ;
        RECT 176.400 30.300 180.600 31.200 ;
        RECT 185.550 32.400 187.350 38.400 ;
        RECT 193.650 35.400 195.450 38.400 ;
        RECT 201.450 35.400 203.250 38.400 ;
        RECT 209.250 36.300 211.050 38.400 ;
        RECT 209.250 35.400 213.000 36.300 ;
        RECT 193.650 34.500 194.700 35.400 ;
        RECT 190.950 33.300 194.700 34.500 ;
        RECT 202.200 34.500 203.250 35.400 ;
        RECT 211.950 34.500 213.000 35.400 ;
        RECT 202.200 33.450 207.150 34.500 ;
        RECT 190.950 32.400 193.050 33.300 ;
        RECT 205.350 32.700 207.150 33.450 ;
        RECT 158.100 25.050 159.900 26.850 ;
        RECT 173.100 25.050 174.900 26.850 ;
        RECT 176.400 25.050 177.600 30.300 ;
        RECT 179.100 25.050 180.900 26.850 ;
        RECT 185.550 25.050 186.750 32.400 ;
        RECT 208.650 31.800 210.450 33.600 ;
        RECT 211.950 32.400 214.050 34.500 ;
        RECT 217.050 32.400 218.850 38.400 ;
        RECT 198.150 30.000 199.950 30.600 ;
        RECT 209.100 30.000 210.150 31.800 ;
        RECT 198.150 28.800 210.150 30.000 ;
        RECT 130.950 22.950 133.050 25.050 ;
        RECT 133.950 22.950 136.050 25.050 ;
        RECT 148.950 22.950 151.050 25.050 ;
        RECT 151.950 22.950 154.050 25.050 ;
        RECT 154.950 22.950 157.050 25.050 ;
        RECT 157.950 22.950 160.050 25.050 ;
        RECT 172.950 22.950 175.050 25.050 ;
        RECT 175.950 22.950 178.050 25.050 ;
        RECT 178.950 22.950 181.050 25.050 ;
        RECT 185.550 23.250 191.850 25.050 ;
        RECT 185.550 22.950 190.050 23.250 ;
        RECT 131.100 21.150 132.900 22.950 ;
        RECT 105.750 17.100 116.850 17.700 ;
        RECT 83.550 3.600 85.350 15.600 ;
        RECT 88.950 15.300 91.050 16.200 ;
        RECT 91.950 15.300 97.050 16.200 ;
        RECT 99.150 16.500 116.850 17.100 ;
        RECT 99.150 16.200 107.550 16.500 ;
        RECT 91.950 14.400 92.850 15.300 ;
        RECT 90.150 12.600 92.850 14.400 ;
        RECT 93.750 14.100 95.550 14.400 ;
        RECT 99.150 14.100 100.050 16.200 ;
        RECT 115.950 15.600 116.850 16.500 ;
        RECT 93.750 13.200 100.050 14.100 ;
        RECT 100.950 14.700 102.750 15.300 ;
        RECT 100.950 13.500 108.450 14.700 ;
        RECT 93.750 12.600 95.550 13.200 ;
        RECT 107.250 12.600 108.450 13.500 ;
        RECT 88.950 9.600 92.850 11.700 ;
        RECT 97.950 11.550 99.750 12.300 ;
        RECT 102.750 11.550 104.550 12.300 ;
        RECT 97.950 10.500 104.550 11.550 ;
        RECT 107.250 10.500 112.050 12.600 ;
        RECT 91.050 3.600 92.850 9.600 ;
        RECT 98.850 3.600 100.650 10.500 ;
        RECT 107.250 9.600 108.450 10.500 ;
        RECT 106.650 3.600 108.450 9.600 ;
        RECT 115.050 3.600 116.850 15.600 ;
        RECT 134.400 9.600 135.600 22.950 ;
        RECT 149.100 21.150 150.900 22.950 ;
        RECT 154.950 9.600 156.150 22.950 ;
        RECT 176.400 9.600 177.600 22.950 ;
        RECT 185.550 15.600 186.750 22.950 ;
        RECT 187.950 17.400 189.750 19.200 ;
        RECT 188.850 16.200 193.050 17.400 ;
        RECT 198.150 16.200 199.050 28.800 ;
        RECT 209.100 27.600 216.000 28.800 ;
        RECT 209.100 27.000 210.900 27.600 ;
        RECT 215.100 26.850 216.000 27.600 ;
        RECT 212.100 25.800 213.900 26.400 ;
        RECT 205.950 24.600 213.900 25.800 ;
        RECT 215.100 25.050 216.900 26.850 ;
        RECT 205.950 22.950 208.050 24.600 ;
        RECT 214.950 22.950 217.050 25.050 ;
        RECT 207.750 17.700 209.550 18.000 ;
        RECT 217.950 17.700 218.850 32.400 ;
        RECT 233.400 31.200 235.200 38.400 ;
        RECT 254.400 31.200 256.200 38.400 ;
        RECT 274.800 32.400 276.600 38.400 ;
        RECT 233.400 30.300 237.600 31.200 ;
        RECT 254.400 30.300 258.600 31.200 ;
        RECT 233.100 25.050 234.900 26.850 ;
        RECT 236.400 25.050 237.600 30.300 ;
        RECT 239.100 25.050 240.900 26.850 ;
        RECT 254.100 25.050 255.900 26.850 ;
        RECT 257.400 25.050 258.600 30.300 ;
        RECT 275.400 30.300 276.600 32.400 ;
        RECT 277.800 33.300 279.600 38.400 ;
        RECT 283.800 33.300 285.600 38.400 ;
        RECT 277.800 31.950 285.600 33.300 ;
        RECT 288.150 32.400 289.950 38.400 ;
        RECT 295.950 36.300 297.750 38.400 ;
        RECT 294.000 35.400 297.750 36.300 ;
        RECT 303.750 35.400 305.550 38.400 ;
        RECT 311.550 35.400 313.350 38.400 ;
        RECT 294.000 34.500 295.050 35.400 ;
        RECT 303.750 34.500 304.800 35.400 ;
        RECT 292.950 32.400 295.050 34.500 ;
        RECT 275.400 29.250 279.150 30.300 ;
        RECT 260.100 25.050 261.900 26.850 ;
        RECT 275.100 25.050 276.900 26.850 ;
        RECT 277.950 25.050 279.150 29.250 ;
        RECT 281.100 25.050 282.900 26.850 ;
        RECT 232.950 22.950 235.050 25.050 ;
        RECT 235.950 22.950 238.050 25.050 ;
        RECT 238.950 22.950 241.050 25.050 ;
        RECT 253.950 22.950 256.050 25.050 ;
        RECT 256.950 22.950 259.050 25.050 ;
        RECT 259.950 22.950 262.050 25.050 ;
        RECT 274.950 22.950 277.050 25.050 ;
        RECT 277.950 22.950 280.050 25.050 ;
        RECT 280.950 22.950 283.050 25.050 ;
        RECT 283.950 22.950 286.050 25.050 ;
        RECT 207.750 17.100 218.850 17.700 ;
        RECT 134.400 3.600 136.200 9.600 ;
        RECT 154.800 3.600 156.600 9.600 ;
        RECT 176.400 3.600 178.200 9.600 ;
        RECT 185.550 3.600 187.350 15.600 ;
        RECT 190.950 15.300 193.050 16.200 ;
        RECT 193.950 15.300 199.050 16.200 ;
        RECT 201.150 16.500 218.850 17.100 ;
        RECT 201.150 16.200 209.550 16.500 ;
        RECT 193.950 14.400 194.850 15.300 ;
        RECT 192.150 12.600 194.850 14.400 ;
        RECT 195.750 14.100 197.550 14.400 ;
        RECT 201.150 14.100 202.050 16.200 ;
        RECT 217.950 15.600 218.850 16.500 ;
        RECT 195.750 13.200 202.050 14.100 ;
        RECT 202.950 14.700 204.750 15.300 ;
        RECT 202.950 13.500 210.450 14.700 ;
        RECT 195.750 12.600 197.550 13.200 ;
        RECT 209.250 12.600 210.450 13.500 ;
        RECT 190.950 9.600 194.850 11.700 ;
        RECT 199.950 11.550 201.750 12.300 ;
        RECT 204.750 11.550 206.550 12.300 ;
        RECT 199.950 10.500 206.550 11.550 ;
        RECT 209.250 10.500 214.050 12.600 ;
        RECT 193.050 3.600 194.850 9.600 ;
        RECT 200.850 3.600 202.650 10.500 ;
        RECT 209.250 9.600 210.450 10.500 ;
        RECT 208.650 3.600 210.450 9.600 ;
        RECT 217.050 3.600 218.850 15.600 ;
        RECT 236.400 9.600 237.600 22.950 ;
        RECT 257.400 9.600 258.600 22.950 ;
        RECT 268.950 18.450 271.050 19.050 ;
        RECT 274.950 18.450 277.050 19.050 ;
        RECT 268.950 17.550 277.050 18.450 ;
        RECT 268.950 16.950 271.050 17.550 ;
        RECT 274.950 16.950 277.050 17.550 ;
        RECT 278.850 9.600 280.050 22.950 ;
        RECT 284.100 21.150 285.900 22.950 ;
        RECT 288.150 17.700 289.050 32.400 ;
        RECT 296.550 31.800 298.350 33.600 ;
        RECT 299.850 33.450 304.800 34.500 ;
        RECT 312.300 34.500 313.350 35.400 ;
        RECT 299.850 32.700 301.650 33.450 ;
        RECT 312.300 33.300 316.050 34.500 ;
        RECT 313.950 32.400 316.050 33.300 ;
        RECT 319.650 32.400 321.450 38.400 ;
        RECT 296.850 30.000 297.900 31.800 ;
        RECT 307.050 30.000 308.850 30.600 ;
        RECT 296.850 28.800 308.850 30.000 ;
        RECT 291.000 27.600 297.900 28.800 ;
        RECT 291.000 26.850 291.900 27.600 ;
        RECT 296.100 27.000 297.900 27.600 ;
        RECT 290.100 25.050 291.900 26.850 ;
        RECT 293.100 25.800 294.900 26.400 ;
        RECT 289.950 22.950 292.050 25.050 ;
        RECT 293.100 24.600 301.050 25.800 ;
        RECT 298.950 22.950 301.050 24.600 ;
        RECT 297.450 17.700 299.250 18.000 ;
        RECT 288.150 17.100 299.250 17.700 ;
        RECT 288.150 16.500 305.850 17.100 ;
        RECT 288.150 15.600 289.050 16.500 ;
        RECT 297.450 16.200 305.850 16.500 ;
        RECT 235.800 3.600 237.600 9.600 ;
        RECT 256.800 3.600 258.600 9.600 ;
        RECT 278.400 3.600 280.200 9.600 ;
        RECT 288.150 3.600 289.950 15.600 ;
        RECT 302.250 14.700 304.050 15.300 ;
        RECT 296.550 13.500 304.050 14.700 ;
        RECT 304.950 14.100 305.850 16.200 ;
        RECT 307.950 16.200 308.850 28.800 ;
        RECT 320.250 25.050 321.450 32.400 ;
        RECT 335.400 35.400 337.200 38.400 ;
        RECT 352.800 35.400 354.600 38.400 ;
        RECT 335.400 25.050 336.600 35.400 ;
        RECT 353.400 25.050 354.600 35.400 ;
        RECT 359.550 32.400 361.350 38.400 ;
        RECT 367.650 35.400 369.450 38.400 ;
        RECT 375.450 35.400 377.250 38.400 ;
        RECT 383.250 36.300 385.050 38.400 ;
        RECT 383.250 35.400 387.000 36.300 ;
        RECT 367.650 34.500 368.700 35.400 ;
        RECT 364.950 33.300 368.700 34.500 ;
        RECT 376.200 34.500 377.250 35.400 ;
        RECT 385.950 34.500 387.000 35.400 ;
        RECT 376.200 33.450 381.150 34.500 ;
        RECT 364.950 32.400 367.050 33.300 ;
        RECT 379.350 32.700 381.150 33.450 ;
        RECT 359.550 25.050 360.750 32.400 ;
        RECT 382.650 31.800 384.450 33.600 ;
        RECT 385.950 32.400 388.050 34.500 ;
        RECT 391.050 32.400 392.850 38.400 ;
        RECT 372.150 30.000 373.950 30.600 ;
        RECT 383.100 30.000 384.150 31.800 ;
        RECT 372.150 28.800 384.150 30.000 ;
        RECT 315.150 23.250 321.450 25.050 ;
        RECT 316.950 22.950 321.450 23.250 ;
        RECT 331.950 22.950 334.050 25.050 ;
        RECT 334.950 22.950 337.050 25.050 ;
        RECT 352.950 22.950 355.050 25.050 ;
        RECT 355.950 22.950 358.050 25.050 ;
        RECT 359.550 23.250 365.850 25.050 ;
        RECT 359.550 22.950 364.050 23.250 ;
        RECT 317.250 17.400 319.050 19.200 ;
        RECT 313.950 16.200 318.150 17.400 ;
        RECT 307.950 15.300 313.050 16.200 ;
        RECT 313.950 15.300 316.050 16.200 ;
        RECT 320.250 15.600 321.450 22.950 ;
        RECT 332.100 21.150 333.900 22.950 ;
        RECT 312.150 14.400 313.050 15.300 ;
        RECT 309.450 14.100 311.250 14.400 ;
        RECT 296.550 12.600 297.750 13.500 ;
        RECT 304.950 13.200 311.250 14.100 ;
        RECT 309.450 12.600 311.250 13.200 ;
        RECT 312.150 12.600 314.850 14.400 ;
        RECT 292.950 10.500 297.750 12.600 ;
        RECT 300.450 11.550 302.250 12.300 ;
        RECT 305.250 11.550 307.050 12.300 ;
        RECT 300.450 10.500 307.050 11.550 ;
        RECT 296.550 9.600 297.750 10.500 ;
        RECT 296.550 3.600 298.350 9.600 ;
        RECT 304.350 3.600 306.150 10.500 ;
        RECT 312.150 9.600 316.050 11.700 ;
        RECT 312.150 3.600 313.950 9.600 ;
        RECT 319.650 3.600 321.450 15.600 ;
        RECT 335.400 9.600 336.600 22.950 ;
        RECT 353.400 9.600 354.600 22.950 ;
        RECT 356.100 21.150 357.900 22.950 ;
        RECT 335.400 3.600 337.200 9.600 ;
        RECT 352.800 3.600 354.600 9.600 ;
        RECT 359.550 15.600 360.750 22.950 ;
        RECT 361.950 17.400 363.750 19.200 ;
        RECT 362.850 16.200 367.050 17.400 ;
        RECT 372.150 16.200 373.050 28.800 ;
        RECT 383.100 27.600 390.000 28.800 ;
        RECT 383.100 27.000 384.900 27.600 ;
        RECT 389.100 26.850 390.000 27.600 ;
        RECT 386.100 25.800 387.900 26.400 ;
        RECT 379.950 24.600 387.900 25.800 ;
        RECT 389.100 25.050 390.900 26.850 ;
        RECT 379.950 22.950 382.050 24.600 ;
        RECT 388.950 22.950 391.050 25.050 ;
        RECT 381.750 17.700 383.550 18.000 ;
        RECT 391.950 17.700 392.850 32.400 ;
        RECT 404.400 33.300 406.200 38.400 ;
        RECT 410.400 33.300 412.200 38.400 ;
        RECT 404.400 31.950 412.200 33.300 ;
        RECT 413.400 32.400 415.200 38.400 ;
        RECT 413.400 30.300 414.600 32.400 ;
        RECT 433.800 31.200 435.600 38.400 ;
        RECT 454.800 31.200 456.600 38.400 ;
        RECT 410.850 29.250 414.600 30.300 ;
        RECT 431.400 30.300 435.600 31.200 ;
        RECT 452.400 30.300 456.600 31.200 ;
        RECT 461.550 32.400 463.350 38.400 ;
        RECT 469.650 35.400 471.450 38.400 ;
        RECT 477.450 35.400 479.250 38.400 ;
        RECT 485.250 36.300 487.050 38.400 ;
        RECT 485.250 35.400 489.000 36.300 ;
        RECT 469.650 34.500 470.700 35.400 ;
        RECT 466.950 33.300 470.700 34.500 ;
        RECT 478.200 34.500 479.250 35.400 ;
        RECT 487.950 34.500 489.000 35.400 ;
        RECT 478.200 33.450 483.150 34.500 ;
        RECT 466.950 32.400 469.050 33.300 ;
        RECT 481.350 32.700 483.150 33.450 ;
        RECT 407.100 25.050 408.900 26.850 ;
        RECT 410.850 25.050 412.050 29.250 ;
        RECT 413.100 25.050 414.900 26.850 ;
        RECT 428.100 25.050 429.900 26.850 ;
        RECT 431.400 25.050 432.600 30.300 ;
        RECT 434.100 25.050 435.900 26.850 ;
        RECT 449.100 25.050 450.900 26.850 ;
        RECT 452.400 25.050 453.600 30.300 ;
        RECT 455.100 25.050 456.900 26.850 ;
        RECT 461.550 25.050 462.750 32.400 ;
        RECT 484.650 31.800 486.450 33.600 ;
        RECT 487.950 32.400 490.050 34.500 ;
        RECT 493.050 32.400 494.850 38.400 ;
        RECT 474.150 30.000 475.950 30.600 ;
        RECT 485.100 30.000 486.150 31.800 ;
        RECT 474.150 28.800 486.150 30.000 ;
        RECT 403.950 22.950 406.050 25.050 ;
        RECT 406.950 22.950 409.050 25.050 ;
        RECT 409.950 22.950 412.050 25.050 ;
        RECT 412.950 22.950 415.050 25.050 ;
        RECT 427.950 22.950 430.050 25.050 ;
        RECT 430.950 22.950 433.050 25.050 ;
        RECT 433.950 22.950 436.050 25.050 ;
        RECT 448.950 22.950 451.050 25.050 ;
        RECT 451.950 22.950 454.050 25.050 ;
        RECT 454.950 22.950 457.050 25.050 ;
        RECT 461.550 23.250 467.850 25.050 ;
        RECT 461.550 22.950 466.050 23.250 ;
        RECT 404.100 21.150 405.900 22.950 ;
        RECT 381.750 17.100 392.850 17.700 ;
        RECT 359.550 3.600 361.350 15.600 ;
        RECT 364.950 15.300 367.050 16.200 ;
        RECT 367.950 15.300 373.050 16.200 ;
        RECT 375.150 16.500 392.850 17.100 ;
        RECT 375.150 16.200 383.550 16.500 ;
        RECT 367.950 14.400 368.850 15.300 ;
        RECT 366.150 12.600 368.850 14.400 ;
        RECT 369.750 14.100 371.550 14.400 ;
        RECT 375.150 14.100 376.050 16.200 ;
        RECT 391.950 15.600 392.850 16.500 ;
        RECT 369.750 13.200 376.050 14.100 ;
        RECT 376.950 14.700 378.750 15.300 ;
        RECT 376.950 13.500 384.450 14.700 ;
        RECT 369.750 12.600 371.550 13.200 ;
        RECT 383.250 12.600 384.450 13.500 ;
        RECT 364.950 9.600 368.850 11.700 ;
        RECT 373.950 11.550 375.750 12.300 ;
        RECT 378.750 11.550 380.550 12.300 ;
        RECT 373.950 10.500 380.550 11.550 ;
        RECT 383.250 10.500 388.050 12.600 ;
        RECT 367.050 3.600 368.850 9.600 ;
        RECT 374.850 3.600 376.650 10.500 ;
        RECT 383.250 9.600 384.450 10.500 ;
        RECT 382.650 3.600 384.450 9.600 ;
        RECT 391.050 3.600 392.850 15.600 ;
        RECT 409.950 9.600 411.150 22.950 ;
        RECT 431.400 9.600 432.600 22.950 ;
        RECT 452.400 9.600 453.600 22.950 ;
        RECT 461.550 15.600 462.750 22.950 ;
        RECT 463.950 17.400 465.750 19.200 ;
        RECT 464.850 16.200 469.050 17.400 ;
        RECT 474.150 16.200 475.050 28.800 ;
        RECT 485.100 27.600 492.000 28.800 ;
        RECT 485.100 27.000 486.900 27.600 ;
        RECT 491.100 26.850 492.000 27.600 ;
        RECT 488.100 25.800 489.900 26.400 ;
        RECT 481.950 24.600 489.900 25.800 ;
        RECT 491.100 25.050 492.900 26.850 ;
        RECT 481.950 22.950 484.050 24.600 ;
        RECT 490.950 22.950 493.050 25.050 ;
        RECT 483.750 17.700 485.550 18.000 ;
        RECT 493.950 17.700 494.850 32.400 ;
        RECT 509.400 35.400 511.200 38.400 ;
        RECT 509.400 25.050 510.600 35.400 ;
        RECT 524.400 33.300 526.200 38.400 ;
        RECT 530.400 33.300 532.200 38.400 ;
        RECT 524.400 31.950 532.200 33.300 ;
        RECT 533.400 32.400 535.200 38.400 ;
        RECT 533.400 30.300 534.600 32.400 ;
        RECT 551.400 31.200 553.200 38.400 ;
        RECT 561.150 32.400 562.950 38.400 ;
        RECT 568.950 36.300 570.750 38.400 ;
        RECT 567.000 35.400 570.750 36.300 ;
        RECT 576.750 35.400 578.550 38.400 ;
        RECT 584.550 35.400 586.350 38.400 ;
        RECT 567.000 34.500 568.050 35.400 ;
        RECT 576.750 34.500 577.800 35.400 ;
        RECT 565.950 32.400 568.050 34.500 ;
        RECT 551.400 30.300 555.600 31.200 ;
        RECT 530.850 29.250 534.600 30.300 ;
        RECT 527.100 25.050 528.900 26.850 ;
        RECT 530.850 25.050 532.050 29.250 ;
        RECT 533.100 25.050 534.900 26.850 ;
        RECT 551.100 25.050 552.900 26.850 ;
        RECT 554.400 25.050 555.600 30.300 ;
        RECT 557.100 25.050 558.900 26.850 ;
        RECT 505.950 22.950 508.050 25.050 ;
        RECT 508.950 22.950 511.050 25.050 ;
        RECT 523.950 22.950 526.050 25.050 ;
        RECT 526.950 22.950 529.050 25.050 ;
        RECT 529.950 22.950 532.050 25.050 ;
        RECT 532.950 22.950 535.050 25.050 ;
        RECT 550.950 22.950 553.050 25.050 ;
        RECT 553.950 22.950 556.050 25.050 ;
        RECT 556.950 22.950 559.050 25.050 ;
        RECT 506.100 21.150 507.900 22.950 ;
        RECT 483.750 17.100 494.850 17.700 ;
        RECT 409.800 3.600 411.600 9.600 ;
        RECT 431.400 3.600 433.200 9.600 ;
        RECT 452.400 3.600 454.200 9.600 ;
        RECT 461.550 3.600 463.350 15.600 ;
        RECT 466.950 15.300 469.050 16.200 ;
        RECT 469.950 15.300 475.050 16.200 ;
        RECT 477.150 16.500 494.850 17.100 ;
        RECT 477.150 16.200 485.550 16.500 ;
        RECT 469.950 14.400 470.850 15.300 ;
        RECT 468.150 12.600 470.850 14.400 ;
        RECT 471.750 14.100 473.550 14.400 ;
        RECT 477.150 14.100 478.050 16.200 ;
        RECT 493.950 15.600 494.850 16.500 ;
        RECT 471.750 13.200 478.050 14.100 ;
        RECT 478.950 14.700 480.750 15.300 ;
        RECT 478.950 13.500 486.450 14.700 ;
        RECT 471.750 12.600 473.550 13.200 ;
        RECT 485.250 12.600 486.450 13.500 ;
        RECT 466.950 9.600 470.850 11.700 ;
        RECT 475.950 11.550 477.750 12.300 ;
        RECT 480.750 11.550 482.550 12.300 ;
        RECT 475.950 10.500 482.550 11.550 ;
        RECT 485.250 10.500 490.050 12.600 ;
        RECT 469.050 3.600 470.850 9.600 ;
        RECT 476.850 3.600 478.650 10.500 ;
        RECT 485.250 9.600 486.450 10.500 ;
        RECT 484.650 3.600 486.450 9.600 ;
        RECT 493.050 3.600 494.850 15.600 ;
        RECT 509.400 9.600 510.600 22.950 ;
        RECT 524.100 21.150 525.900 22.950 ;
        RECT 529.950 9.600 531.150 22.950 ;
        RECT 554.400 9.600 555.600 22.950 ;
        RECT 509.400 3.600 511.200 9.600 ;
        RECT 529.800 3.600 531.600 9.600 ;
        RECT 553.800 3.600 555.600 9.600 ;
        RECT 561.150 17.700 562.050 32.400 ;
        RECT 569.550 31.800 571.350 33.600 ;
        RECT 572.850 33.450 577.800 34.500 ;
        RECT 585.300 34.500 586.350 35.400 ;
        RECT 572.850 32.700 574.650 33.450 ;
        RECT 585.300 33.300 589.050 34.500 ;
        RECT 586.950 32.400 589.050 33.300 ;
        RECT 592.650 32.400 594.450 38.400 ;
        RECT 569.850 30.000 570.900 31.800 ;
        RECT 580.050 30.000 581.850 30.600 ;
        RECT 569.850 28.800 581.850 30.000 ;
        RECT 564.000 27.600 570.900 28.800 ;
        RECT 564.000 26.850 564.900 27.600 ;
        RECT 569.100 27.000 570.900 27.600 ;
        RECT 563.100 25.050 564.900 26.850 ;
        RECT 566.100 25.800 567.900 26.400 ;
        RECT 562.950 22.950 565.050 25.050 ;
        RECT 566.100 24.600 574.050 25.800 ;
        RECT 571.950 22.950 574.050 24.600 ;
        RECT 570.450 17.700 572.250 18.000 ;
        RECT 561.150 17.100 572.250 17.700 ;
        RECT 561.150 16.500 578.850 17.100 ;
        RECT 561.150 15.600 562.050 16.500 ;
        RECT 570.450 16.200 578.850 16.500 ;
        RECT 561.150 3.600 562.950 15.600 ;
        RECT 575.250 14.700 577.050 15.300 ;
        RECT 569.550 13.500 577.050 14.700 ;
        RECT 577.950 14.100 578.850 16.200 ;
        RECT 580.950 16.200 581.850 28.800 ;
        RECT 593.250 25.050 594.450 32.400 ;
        RECT 608.400 31.200 610.200 38.400 ;
        RECT 626.400 33.300 628.200 38.400 ;
        RECT 632.400 33.300 634.200 38.400 ;
        RECT 626.400 31.950 634.200 33.300 ;
        RECT 635.400 32.400 637.200 38.400 ;
        RECT 641.550 32.400 643.350 38.400 ;
        RECT 649.650 35.400 651.450 38.400 ;
        RECT 657.450 35.400 659.250 38.400 ;
        RECT 665.250 36.300 667.050 38.400 ;
        RECT 665.250 35.400 669.000 36.300 ;
        RECT 649.650 34.500 650.700 35.400 ;
        RECT 646.950 33.300 650.700 34.500 ;
        RECT 658.200 34.500 659.250 35.400 ;
        RECT 667.950 34.500 669.000 35.400 ;
        RECT 658.200 33.450 663.150 34.500 ;
        RECT 646.950 32.400 649.050 33.300 ;
        RECT 661.350 32.700 663.150 33.450 ;
        RECT 608.400 30.300 612.600 31.200 ;
        RECT 608.100 25.050 609.900 26.850 ;
        RECT 611.400 25.050 612.600 30.300 ;
        RECT 613.950 30.450 616.050 31.050 ;
        RECT 613.950 29.550 621.450 30.450 ;
        RECT 635.400 30.300 636.600 32.400 ;
        RECT 613.950 28.950 616.050 29.550 ;
        RECT 614.100 25.050 615.900 26.850 ;
        RECT 588.150 23.250 594.450 25.050 ;
        RECT 589.950 22.950 594.450 23.250 ;
        RECT 607.950 22.950 610.050 25.050 ;
        RECT 610.950 22.950 613.050 25.050 ;
        RECT 613.950 22.950 616.050 25.050 ;
        RECT 590.250 17.400 592.050 19.200 ;
        RECT 586.950 16.200 591.150 17.400 ;
        RECT 580.950 15.300 586.050 16.200 ;
        RECT 586.950 15.300 589.050 16.200 ;
        RECT 593.250 15.600 594.450 22.950 ;
        RECT 585.150 14.400 586.050 15.300 ;
        RECT 582.450 14.100 584.250 14.400 ;
        RECT 569.550 12.600 570.750 13.500 ;
        RECT 577.950 13.200 584.250 14.100 ;
        RECT 582.450 12.600 584.250 13.200 ;
        RECT 585.150 12.600 587.850 14.400 ;
        RECT 565.950 10.500 570.750 12.600 ;
        RECT 573.450 11.550 575.250 12.300 ;
        RECT 578.250 11.550 580.050 12.300 ;
        RECT 573.450 10.500 580.050 11.550 ;
        RECT 569.550 9.600 570.750 10.500 ;
        RECT 569.550 3.600 571.350 9.600 ;
        RECT 577.350 3.600 579.150 10.500 ;
        RECT 585.150 9.600 589.050 11.700 ;
        RECT 585.150 3.600 586.950 9.600 ;
        RECT 592.650 3.600 594.450 15.600 ;
        RECT 611.400 9.600 612.600 22.950 ;
        RECT 620.550 22.050 621.450 29.550 ;
        RECT 632.850 29.250 636.600 30.300 ;
        RECT 629.100 25.050 630.900 26.850 ;
        RECT 632.850 25.050 634.050 29.250 ;
        RECT 635.100 25.050 636.900 26.850 ;
        RECT 641.550 25.050 642.750 32.400 ;
        RECT 664.650 31.800 666.450 33.600 ;
        RECT 667.950 32.400 670.050 34.500 ;
        RECT 673.050 32.400 674.850 38.400 ;
        RECT 654.150 30.000 655.950 30.600 ;
        RECT 665.100 30.000 666.150 31.800 ;
        RECT 654.150 28.800 666.150 30.000 ;
        RECT 625.950 22.950 628.050 25.050 ;
        RECT 628.950 22.950 631.050 25.050 ;
        RECT 631.950 22.950 634.050 25.050 ;
        RECT 634.950 22.950 637.050 25.050 ;
        RECT 641.550 23.250 647.850 25.050 ;
        RECT 641.550 22.950 646.050 23.250 ;
        RECT 620.550 20.550 625.050 22.050 ;
        RECT 626.100 21.150 627.900 22.950 ;
        RECT 621.000 19.950 625.050 20.550 ;
        RECT 631.950 9.600 633.150 22.950 ;
        RECT 641.550 15.600 642.750 22.950 ;
        RECT 643.950 17.400 645.750 19.200 ;
        RECT 644.850 16.200 649.050 17.400 ;
        RECT 654.150 16.200 655.050 28.800 ;
        RECT 665.100 27.600 672.000 28.800 ;
        RECT 665.100 27.000 666.900 27.600 ;
        RECT 671.100 26.850 672.000 27.600 ;
        RECT 668.100 25.800 669.900 26.400 ;
        RECT 661.950 24.600 669.900 25.800 ;
        RECT 671.100 25.050 672.900 26.850 ;
        RECT 661.950 22.950 664.050 24.600 ;
        RECT 670.950 22.950 673.050 25.050 ;
        RECT 663.750 17.700 665.550 18.000 ;
        RECT 673.950 17.700 674.850 32.400 ;
        RECT 689.400 31.200 691.200 38.400 ;
        RECT 709.800 32.400 711.600 38.400 ;
        RECT 689.400 30.300 693.600 31.200 ;
        RECT 689.100 25.050 690.900 26.850 ;
        RECT 692.400 25.050 693.600 30.300 ;
        RECT 710.400 30.300 711.600 32.400 ;
        RECT 712.800 33.300 714.600 38.400 ;
        RECT 718.800 33.300 720.600 38.400 ;
        RECT 712.800 31.950 720.600 33.300 ;
        RECT 736.800 31.200 738.600 38.400 ;
        RECT 739.950 36.450 742.050 37.050 ;
        RECT 745.950 36.450 748.050 36.900 ;
        RECT 739.950 35.550 748.050 36.450 ;
        RECT 739.950 34.950 742.050 35.550 ;
        RECT 745.950 34.800 748.050 35.550 ;
        RECT 754.800 32.400 756.600 38.400 ;
        RECT 760.800 35.400 762.600 38.400 ;
        RECT 734.400 30.300 738.600 31.200 ;
        RECT 710.400 29.250 714.150 30.300 ;
        RECT 695.100 25.050 696.900 26.850 ;
        RECT 710.100 25.050 711.900 26.850 ;
        RECT 712.950 25.050 714.150 29.250 ;
        RECT 716.100 25.050 717.900 26.850 ;
        RECT 731.100 25.050 732.900 26.850 ;
        RECT 734.400 25.050 735.600 30.300 ;
        RECT 737.100 25.050 738.900 26.850 ;
        RECT 754.950 25.050 756.000 32.400 ;
        RECT 760.800 31.200 761.700 35.400 ;
        RECT 780.300 34.200 782.100 38.400 ;
        RECT 758.400 30.300 761.700 31.200 ;
        RECT 779.400 32.400 782.100 34.200 ;
        RECT 758.400 29.400 760.200 30.300 ;
        RECT 688.950 22.950 691.050 25.050 ;
        RECT 691.950 22.950 694.050 25.050 ;
        RECT 694.950 22.950 697.050 25.050 ;
        RECT 709.950 22.950 712.050 25.050 ;
        RECT 712.950 22.950 715.050 25.050 ;
        RECT 715.950 22.950 718.050 25.050 ;
        RECT 718.950 22.950 721.050 25.050 ;
        RECT 730.950 22.950 733.050 25.050 ;
        RECT 733.950 22.950 736.050 25.050 ;
        RECT 736.950 22.950 739.050 25.050 ;
        RECT 754.950 22.950 757.050 25.050 ;
        RECT 663.750 17.100 674.850 17.700 ;
        RECT 610.800 3.600 612.600 9.600 ;
        RECT 631.800 3.600 633.600 9.600 ;
        RECT 641.550 3.600 643.350 15.600 ;
        RECT 646.950 15.300 649.050 16.200 ;
        RECT 649.950 15.300 655.050 16.200 ;
        RECT 657.150 16.500 674.850 17.100 ;
        RECT 657.150 16.200 665.550 16.500 ;
        RECT 649.950 14.400 650.850 15.300 ;
        RECT 648.150 12.600 650.850 14.400 ;
        RECT 651.750 14.100 653.550 14.400 ;
        RECT 657.150 14.100 658.050 16.200 ;
        RECT 673.950 15.600 674.850 16.500 ;
        RECT 651.750 13.200 658.050 14.100 ;
        RECT 658.950 14.700 660.750 15.300 ;
        RECT 658.950 13.500 666.450 14.700 ;
        RECT 651.750 12.600 653.550 13.200 ;
        RECT 665.250 12.600 666.450 13.500 ;
        RECT 646.950 9.600 650.850 11.700 ;
        RECT 655.950 11.550 657.750 12.300 ;
        RECT 660.750 11.550 662.550 12.300 ;
        RECT 655.950 10.500 662.550 11.550 ;
        RECT 665.250 10.500 670.050 12.600 ;
        RECT 649.050 3.600 650.850 9.600 ;
        RECT 656.850 3.600 658.650 10.500 ;
        RECT 665.250 9.600 666.450 10.500 ;
        RECT 664.650 3.600 666.450 9.600 ;
        RECT 673.050 3.600 674.850 15.600 ;
        RECT 692.400 9.600 693.600 22.950 ;
        RECT 703.950 18.450 706.050 19.050 ;
        RECT 709.950 18.450 712.050 19.050 ;
        RECT 703.950 17.550 712.050 18.450 ;
        RECT 703.950 16.950 706.050 17.550 ;
        RECT 709.950 16.950 712.050 17.550 ;
        RECT 713.850 9.600 715.050 22.950 ;
        RECT 719.100 21.150 720.900 22.950 ;
        RECT 734.400 9.600 735.600 22.950 ;
        RECT 755.700 15.600 757.050 22.950 ;
        RECT 758.400 18.900 759.300 29.400 ;
        RECT 764.100 25.050 765.900 26.850 ;
        RECT 779.400 25.050 780.300 32.400 ;
        RECT 782.100 30.600 783.900 31.500 ;
        RECT 787.800 30.600 789.600 38.400 ;
        RECT 800.400 33.300 802.200 38.400 ;
        RECT 806.400 33.300 808.200 38.400 ;
        RECT 800.400 31.950 808.200 33.300 ;
        RECT 809.400 32.400 811.200 38.400 ;
        RECT 827.400 35.400 829.200 38.400 ;
        RECT 782.100 29.700 789.600 30.600 ;
        RECT 809.400 30.300 810.600 32.400 ;
        RECT 760.950 22.950 763.050 25.050 ;
        RECT 763.950 22.950 766.050 25.050 ;
        RECT 778.950 22.950 781.050 25.050 ;
        RECT 781.950 22.950 784.050 25.050 ;
        RECT 761.100 21.150 762.900 22.950 ;
        RECT 758.400 18.300 760.200 18.900 ;
        RECT 758.400 17.100 765.600 18.300 ;
        RECT 764.400 15.600 765.600 17.100 ;
        RECT 779.400 15.600 780.300 22.950 ;
        RECT 782.100 21.150 783.900 22.950 ;
        RECT 755.700 14.100 758.100 15.600 ;
        RECT 691.800 3.600 693.600 9.600 ;
        RECT 713.400 3.600 715.200 9.600 ;
        RECT 734.400 3.600 736.200 9.600 ;
        RECT 756.300 3.600 758.100 14.100 ;
        RECT 763.800 3.600 765.600 15.600 ;
        RECT 778.800 3.600 780.600 15.600 ;
        RECT 785.700 9.600 786.600 29.700 ;
        RECT 806.850 29.250 810.600 30.300 ;
        RECT 788.100 25.050 789.900 26.850 ;
        RECT 803.100 25.050 804.900 26.850 ;
        RECT 806.850 25.050 808.050 29.250 ;
        RECT 809.100 25.050 810.900 26.850 ;
        RECT 827.400 25.050 828.600 35.400 ;
        RECT 847.500 33.600 849.300 38.400 ;
        RECT 847.500 32.400 852.600 33.600 ;
        RECT 868.800 32.400 870.600 38.400 ;
        RECT 842.100 25.050 843.900 26.850 ;
        RECT 848.100 25.050 849.900 26.850 ;
        RECT 851.700 25.050 852.600 32.400 ;
        RECT 869.400 30.300 870.600 32.400 ;
        RECT 871.800 33.300 873.600 38.400 ;
        RECT 877.800 33.300 879.600 38.400 ;
        RECT 871.800 31.950 879.600 33.300 ;
        RECT 869.400 29.250 873.150 30.300 ;
        RECT 869.100 25.050 870.900 26.850 ;
        RECT 871.950 25.050 873.150 29.250 ;
        RECT 875.100 25.050 876.900 26.850 ;
        RECT 787.950 22.950 790.050 25.050 ;
        RECT 799.950 22.950 802.050 25.050 ;
        RECT 802.950 22.950 805.050 25.050 ;
        RECT 805.950 22.950 808.050 25.050 ;
        RECT 808.950 22.950 811.050 25.050 ;
        RECT 823.950 22.950 826.050 25.050 ;
        RECT 826.950 22.950 829.050 25.050 ;
        RECT 841.950 22.950 844.050 25.050 ;
        RECT 844.950 22.950 847.050 25.050 ;
        RECT 847.950 22.950 850.050 25.050 ;
        RECT 850.950 22.950 853.050 25.050 ;
        RECT 868.950 22.950 871.050 25.050 ;
        RECT 871.950 22.950 874.050 25.050 ;
        RECT 874.950 22.950 877.050 25.050 ;
        RECT 877.950 22.950 880.050 25.050 ;
        RECT 800.100 21.150 801.900 22.950 ;
        RECT 805.950 9.600 807.150 22.950 ;
        RECT 824.100 21.150 825.900 22.950 ;
        RECT 827.400 9.600 828.600 22.950 ;
        RECT 845.100 21.150 846.900 22.950 ;
        RECT 851.700 15.600 852.600 22.950 ;
        RECT 842.400 14.700 850.200 15.600 ;
        RECT 784.800 3.600 786.600 9.600 ;
        RECT 805.800 3.600 807.600 9.600 ;
        RECT 827.400 3.600 829.200 9.600 ;
        RECT 842.400 3.600 844.200 14.700 ;
        RECT 848.400 3.600 850.200 14.700 ;
        RECT 851.400 3.600 853.200 15.600 ;
        RECT 872.850 9.600 874.050 22.950 ;
        RECT 878.100 21.150 879.900 22.950 ;
        RECT 872.400 3.600 874.200 9.600 ;
      LAYER metal2 ;
        RECT 256.950 892.950 259.050 895.050 ;
        RECT 268.950 892.950 271.050 895.050 ;
        RECT 310.950 892.950 313.050 895.050 ;
        RECT 322.950 892.950 325.050 895.050 ;
        RECT 334.950 892.950 337.050 895.050 ;
        RECT 364.950 894.600 367.050 895.050 ;
        RECT 370.950 894.600 373.050 895.050 ;
        RECT 364.950 893.400 373.050 894.600 ;
        RECT 364.950 892.950 367.050 893.400 ;
        RECT 370.950 892.950 373.050 893.400 ;
        RECT 394.950 892.950 397.050 895.050 ;
        RECT 562.950 892.950 565.050 895.050 ;
        RECT 679.950 892.950 682.050 895.050 ;
        RECT 688.950 892.950 691.050 895.050 ;
        RECT 778.950 892.950 781.050 895.050 ;
        RECT 46.950 890.400 49.050 892.500 ;
        RECT 67.950 890.400 70.050 892.500 ;
        RECT 82.950 890.400 85.050 892.500 ;
        RECT 103.950 890.400 106.050 892.500 ;
        RECT 22.950 886.950 25.050 889.050 ;
        RECT 16.950 884.100 19.050 886.200 ;
        RECT 17.400 883.050 18.600 884.100 ;
        RECT 13.950 880.950 16.050 883.050 ;
        RECT 16.950 880.950 19.050 883.050 ;
        RECT 14.400 879.900 15.600 880.950 ;
        RECT 13.950 877.800 16.050 879.900 ;
        RECT 10.950 839.100 13.050 841.200 ;
        RECT 19.800 839.100 21.900 841.200 ;
        RECT 23.400 841.050 24.600 886.950 ;
        RECT 31.950 885.000 34.050 889.050 ;
        RECT 32.400 883.050 33.600 885.000 ;
        RECT 43.950 884.400 46.050 886.500 ;
        RECT 44.400 883.050 45.600 884.400 ;
        RECT 28.950 880.950 31.050 883.050 ;
        RECT 31.950 880.950 34.050 883.050 ;
        RECT 34.950 880.950 37.050 883.050 ;
        RECT 43.950 880.950 46.050 883.050 ;
        RECT 29.400 879.900 30.600 880.950 ;
        RECT 35.400 879.900 36.600 880.950 ;
        RECT 25.800 877.800 27.900 879.900 ;
        RECT 28.950 877.800 31.050 879.900 ;
        RECT 34.950 877.800 37.050 879.900 ;
        RECT 11.400 838.050 12.600 839.100 ;
        RECT 20.400 838.050 21.600 839.100 ;
        RECT 22.950 838.950 25.050 841.050 ;
        RECT 10.950 835.950 13.050 838.050 ;
        RECT 16.950 835.950 19.050 838.050 ;
        RECT 19.950 835.950 22.050 838.050 ;
        RECT 7.950 832.950 10.050 835.050 ;
        RECT 13.800 832.950 15.900 835.050 ;
        RECT 17.400 834.900 18.600 835.950 ;
        RECT 8.400 826.050 9.600 832.950 ;
        RECT 14.400 829.050 15.600 832.950 ;
        RECT 16.950 832.800 19.050 834.900 ;
        RECT 22.950 832.950 25.050 835.050 ;
        RECT 13.950 826.950 16.050 829.050 ;
        RECT 19.950 826.950 22.050 829.050 ;
        RECT 7.950 823.950 10.050 826.050 ;
        RECT 13.950 823.800 16.050 825.900 ;
        RECT 4.950 806.100 7.050 808.200 ;
        RECT 1.950 766.950 4.050 769.050 ;
        RECT 2.400 631.050 3.600 766.950 ;
        RECT 5.400 670.050 6.600 806.100 ;
        RECT 14.400 805.050 15.600 823.800 ;
        RECT 20.400 808.050 21.600 826.950 ;
        RECT 19.950 805.950 22.050 808.050 ;
        RECT 10.950 802.950 13.050 805.050 ;
        RECT 13.950 802.950 16.050 805.050 ;
        RECT 16.950 802.950 19.050 805.050 ;
        RECT 11.400 801.000 12.600 802.950 ;
        RECT 10.950 796.950 13.050 801.000 ;
        RECT 17.400 781.050 18.600 802.950 ;
        RECT 16.950 778.950 19.050 781.050 ;
        RECT 7.950 760.950 10.050 763.050 ;
        RECT 13.950 761.100 16.050 763.200 ;
        RECT 8.400 730.050 9.600 760.950 ;
        RECT 14.400 760.050 15.600 761.100 ;
        RECT 13.950 757.950 16.050 760.050 ;
        RECT 16.950 757.950 19.050 760.050 ;
        RECT 17.400 756.900 18.600 757.950 ;
        RECT 16.950 754.800 19.050 756.900 ;
        RECT 13.950 748.950 16.050 751.050 ;
        RECT 7.950 727.950 10.050 730.050 ;
        RECT 14.400 727.050 15.600 748.950 ;
        RECT 10.950 724.950 13.050 727.050 ;
        RECT 13.950 724.950 16.050 727.050 ;
        RECT 16.950 724.950 19.050 727.050 ;
        RECT 11.400 723.900 12.600 724.950 ;
        RECT 17.400 723.900 18.600 724.950 ;
        RECT 10.950 723.600 13.050 723.900 ;
        RECT 8.400 722.400 13.050 723.600 ;
        RECT 4.950 667.950 7.050 670.050 ;
        RECT 4.950 661.950 7.050 664.050 ;
        RECT 1.950 628.950 4.050 631.050 ;
        RECT 5.400 544.050 6.600 661.950 ;
        RECT 8.400 658.050 9.600 722.400 ;
        RECT 10.950 721.800 13.050 722.400 ;
        RECT 16.950 721.800 19.050 723.900 ;
        RECT 19.950 697.950 22.050 700.050 ;
        RECT 13.950 691.950 16.050 694.050 ;
        RECT 14.400 682.050 15.600 691.950 ;
        RECT 20.400 682.050 21.600 697.950 ;
        RECT 23.400 688.050 24.600 832.950 ;
        RECT 26.400 799.050 27.600 877.800 ;
        RECT 47.850 875.400 49.050 890.400 ;
        RECT 55.950 884.400 58.050 886.500 ;
        RECT 56.400 880.050 57.600 884.400 ;
        RECT 61.950 880.950 64.050 883.050 ;
        RECT 55.950 877.950 58.050 880.050 ;
        RECT 46.950 873.300 49.050 875.400 ;
        RECT 47.850 869.700 49.050 873.300 ;
        RECT 46.950 867.600 49.050 869.700 ;
        RECT 49.950 849.300 52.050 851.400 ;
        RECT 50.850 845.700 52.050 849.300 ;
        RECT 49.950 843.600 52.050 845.700 ;
        RECT 28.950 838.950 31.050 841.050 ;
        RECT 37.950 839.100 40.050 841.200 ;
        RECT 29.400 834.900 30.600 838.950 ;
        RECT 38.400 838.050 39.600 839.100 ;
        RECT 34.950 835.950 37.050 838.050 ;
        RECT 37.950 835.950 40.050 838.050 ;
        RECT 46.950 835.950 49.050 838.050 ;
        RECT 28.950 832.800 31.050 834.900 ;
        RECT 35.400 820.050 36.600 835.950 ;
        RECT 43.950 832.950 46.050 835.050 ;
        RECT 47.400 834.000 48.600 835.950 ;
        RECT 37.950 829.950 40.050 832.050 ;
        RECT 34.950 817.950 37.050 820.050 ;
        RECT 31.950 806.100 34.050 808.200 ;
        RECT 38.400 808.050 39.600 829.950 ;
        RECT 40.950 823.950 43.050 826.050 ;
        RECT 32.400 805.050 33.600 806.100 ;
        RECT 37.950 805.950 40.050 808.050 ;
        RECT 31.950 802.950 34.050 805.050 ;
        RECT 34.950 802.950 37.050 805.050 ;
        RECT 28.950 799.950 31.050 802.050 ;
        RECT 35.400 801.900 36.600 802.950 ;
        RECT 41.400 802.050 42.600 823.950 ;
        RECT 25.950 796.950 28.050 799.050 ;
        RECT 29.400 763.200 30.600 799.950 ;
        RECT 34.950 799.800 37.050 801.900 ;
        RECT 40.950 799.950 43.050 802.050 ;
        RECT 35.400 769.050 36.600 799.800 ;
        RECT 40.950 796.800 43.050 798.900 ;
        RECT 34.950 766.950 37.050 769.050 ;
        RECT 28.950 761.100 31.050 763.200 ;
        RECT 34.950 761.100 37.050 763.200 ;
        RECT 29.400 760.050 30.600 761.100 ;
        RECT 35.400 760.050 36.600 761.100 ;
        RECT 28.950 757.950 31.050 760.050 ;
        RECT 31.950 757.950 34.050 760.050 ;
        RECT 34.950 757.950 37.050 760.050 ;
        RECT 32.400 756.900 33.600 757.950 ;
        RECT 31.950 754.800 34.050 756.900 ;
        RECT 31.950 729.000 34.050 733.050 ;
        RECT 32.400 727.050 33.600 729.000 ;
        RECT 31.950 724.950 34.050 727.050 ;
        RECT 34.950 724.950 37.050 727.050 ;
        RECT 35.400 723.900 36.600 724.950 ;
        RECT 41.400 724.050 42.600 796.800 ;
        RECT 44.400 781.050 45.600 832.950 ;
        RECT 46.950 829.950 49.050 834.000 ;
        RECT 50.850 828.600 52.050 843.600 ;
        RECT 49.950 826.500 52.050 828.600 ;
        RECT 56.400 820.050 57.600 877.950 ;
        RECT 62.400 840.600 63.600 880.950 ;
        RECT 68.100 870.600 69.300 890.400 ;
        RECT 79.950 884.400 82.050 886.500 ;
        RECT 80.400 883.050 81.600 884.400 ;
        RECT 70.950 880.950 73.050 883.050 ;
        RECT 79.950 880.950 82.050 883.050 ;
        RECT 71.400 879.000 72.600 880.950 ;
        RECT 70.950 874.950 73.050 879.000 ;
        RECT 76.950 874.950 79.050 877.050 ;
        RECT 83.850 875.400 85.050 890.400 ;
        RECT 97.950 880.950 100.050 883.050 ;
        RECT 67.950 868.500 70.050 870.600 ;
        RECT 70.950 848.400 73.050 850.500 ;
        RECT 59.400 839.400 63.600 840.600 ;
        RECT 64.950 839.400 67.050 841.500 ;
        RECT 55.950 817.950 58.050 820.050 ;
        RECT 59.400 810.600 60.600 839.400 ;
        RECT 65.400 838.050 66.600 839.400 ;
        RECT 64.950 835.950 67.050 838.050 ;
        RECT 71.100 828.600 72.300 848.400 ;
        RECT 77.400 844.050 78.600 874.950 ;
        RECT 82.950 873.300 85.050 875.400 ;
        RECT 83.850 869.700 85.050 873.300 ;
        RECT 82.950 867.600 85.050 869.700 ;
        RECT 98.400 862.050 99.600 880.950 ;
        RECT 104.100 870.600 105.300 890.400 ;
        RECT 166.950 889.950 169.050 892.050 ;
        RECT 163.650 887.400 165.750 889.500 ;
        RECT 106.950 880.950 109.050 883.050 ;
        RECT 145.950 880.950 148.050 883.050 ;
        RECT 161.400 881.100 163.500 883.200 ;
        RECT 107.400 880.050 108.600 880.950 ;
        RECT 107.400 879.000 112.050 880.050 ;
        RECT 146.400 879.900 147.600 880.950 ;
        RECT 106.950 877.950 112.050 879.000 ;
        RECT 106.950 874.950 109.050 877.950 ;
        RECT 145.950 877.800 148.050 879.900 ;
        RECT 161.400 878.550 162.600 881.100 ;
        RECT 164.400 874.800 165.300 887.400 ;
        RECT 167.400 885.900 168.600 889.950 ;
        RECT 170.400 888.900 171.600 891.450 ;
        RECT 196.950 889.950 199.050 892.050 ;
        RECT 226.950 889.950 229.050 892.050 ;
        RECT 244.950 889.950 247.050 892.050 ;
        RECT 170.400 886.800 172.500 888.900 ;
        RECT 173.700 887.100 175.800 889.200 ;
        RECT 166.200 885.000 168.600 885.900 ;
        RECT 166.200 883.800 173.250 885.000 ;
        RECT 171.150 882.900 173.250 883.800 ;
        RECT 166.200 882.000 168.300 882.900 ;
        RECT 174.150 882.000 175.050 887.100 ;
        RECT 176.400 883.200 177.600 885.600 ;
        RECT 181.950 883.950 184.050 886.050 ;
        RECT 166.200 881.100 175.050 882.000 ;
        RECT 175.950 881.100 178.050 883.200 ;
        RECT 166.200 880.800 168.300 881.100 ;
        RECT 170.400 878.100 172.500 880.200 ;
        RECT 164.100 872.700 166.200 874.800 ;
        RECT 103.950 868.500 106.050 870.600 ;
        RECT 97.950 859.950 100.050 862.050 ;
        RECT 106.950 859.950 109.050 862.050 ;
        RECT 97.950 853.950 100.050 856.050 ;
        RECT 76.950 841.950 79.050 844.050 ;
        RECT 82.950 841.950 85.050 844.050 ;
        RECT 77.400 840.600 78.600 841.950 ;
        RECT 74.400 839.400 78.600 840.600 ;
        RECT 74.400 838.050 75.600 839.400 ;
        RECT 73.950 835.950 76.050 838.050 ;
        RECT 70.950 826.500 73.050 828.600 ;
        RECT 70.950 812.400 73.050 814.500 ;
        RECT 56.400 809.400 60.600 810.600 ;
        RECT 56.400 805.050 57.600 809.400 ;
        RECT 61.950 806.100 64.050 808.200 ;
        RECT 62.400 805.050 63.600 806.100 ;
        RECT 52.950 802.950 55.050 805.050 ;
        RECT 55.950 802.950 58.050 805.050 ;
        RECT 58.950 802.950 61.050 805.050 ;
        RECT 61.950 802.950 64.050 805.050 ;
        RECT 67.950 802.950 70.050 805.050 ;
        RECT 53.400 801.000 54.600 802.950 ;
        RECT 59.400 801.000 60.600 802.950 ;
        RECT 68.400 801.000 69.600 802.950 ;
        RECT 46.950 796.950 49.050 799.050 ;
        RECT 52.950 796.950 55.050 801.000 ;
        RECT 58.950 796.950 61.050 801.000 ;
        RECT 67.950 796.950 70.050 801.000 ;
        RECT 43.950 778.950 46.050 781.050 ;
        RECT 43.950 761.100 46.050 763.200 ;
        RECT 47.400 763.050 48.600 796.950 ;
        RECT 71.700 792.600 72.900 812.400 ;
        RECT 76.950 802.950 79.050 805.050 ;
        RECT 77.400 793.050 78.600 802.950 ;
        RECT 83.400 799.050 84.600 841.950 ;
        RECT 91.950 839.100 94.050 841.200 ;
        RECT 92.400 838.050 93.600 839.100 ;
        RECT 98.400 838.050 99.600 853.950 ;
        RECT 88.950 835.950 91.050 838.050 ;
        RECT 91.950 835.950 94.050 838.050 ;
        RECT 94.950 835.950 97.050 838.050 ;
        RECT 97.950 835.950 100.050 838.050 ;
        RECT 100.950 835.950 103.050 838.050 ;
        RECT 89.400 826.050 90.600 835.950 ;
        RECT 95.400 834.900 96.600 835.950 ;
        RECT 94.950 832.800 97.050 834.900 ;
        RECT 101.400 834.000 102.600 835.950 ;
        RECT 107.400 834.900 108.600 859.950 ;
        RECT 151.950 853.950 154.050 856.050 ;
        RECT 148.950 847.950 151.050 850.050 ;
        RECT 109.950 839.100 112.050 841.200 ;
        RECT 118.950 839.100 121.050 841.200 ;
        RECT 124.950 840.000 127.050 844.050 ;
        RECT 133.950 841.950 136.050 844.050 ;
        RECT 100.950 829.950 103.050 834.000 ;
        RECT 106.950 832.800 109.050 834.900 ;
        RECT 88.950 823.950 91.050 826.050 ;
        RECT 85.950 811.950 88.050 814.050 ;
        RECT 91.950 812.400 94.050 814.500 ;
        RECT 110.400 814.050 111.600 839.100 ;
        RECT 119.400 838.050 120.600 839.100 ;
        RECT 125.400 838.050 126.600 840.000 ;
        RECT 115.950 835.950 118.050 838.050 ;
        RECT 118.950 835.950 121.050 838.050 ;
        RECT 121.950 835.950 124.050 838.050 ;
        RECT 124.950 835.950 127.050 838.050 ;
        RECT 127.950 835.950 130.050 838.050 ;
        RECT 116.400 831.600 117.600 835.950 ;
        RECT 122.400 834.900 123.600 835.950 ;
        RECT 121.950 832.800 124.050 834.900 ;
        RECT 116.400 830.400 120.600 831.600 ;
        RECT 86.400 808.200 87.600 811.950 ;
        RECT 85.950 806.100 88.050 808.200 ;
        RECT 82.950 796.950 85.050 799.050 ;
        RECT 91.950 797.400 93.150 812.400 ;
        RECT 109.950 811.950 112.050 814.050 ;
        RECT 94.950 806.400 97.050 808.500 ;
        RECT 95.400 805.050 96.600 806.400 ;
        RECT 103.950 806.100 106.050 808.200 ;
        RECT 109.950 806.100 112.050 808.200 ;
        RECT 94.950 802.950 97.050 805.050 ;
        RECT 104.400 801.600 105.600 806.100 ;
        RECT 110.400 805.050 111.600 806.100 ;
        RECT 109.950 802.950 112.050 805.050 ;
        RECT 112.950 802.950 115.050 805.050 ;
        RECT 113.400 801.900 114.600 802.950 ;
        RECT 104.400 800.400 108.600 801.600 ;
        RECT 70.950 790.500 73.050 792.600 ;
        RECT 76.950 790.950 79.050 793.050 ;
        RECT 52.950 778.950 55.050 781.050 ;
        RECT 44.400 757.050 45.600 761.100 ;
        RECT 46.950 760.950 49.050 763.050 ;
        RECT 53.400 760.050 54.600 778.950 ;
        RECT 83.400 769.050 84.600 796.950 ;
        RECT 91.950 795.300 94.050 797.400 ;
        RECT 91.950 791.700 93.150 795.300 ;
        RECT 91.950 789.600 94.050 791.700 ;
        RECT 82.950 766.950 85.050 769.050 ;
        RECT 58.950 761.100 61.050 763.200 ;
        RECT 73.950 761.100 76.050 763.200 ;
        RECT 79.950 762.000 82.050 766.050 ;
        RECT 85.950 763.950 88.050 766.050 ;
        RECT 59.400 760.050 60.600 761.100 ;
        RECT 74.400 760.050 75.600 761.100 ;
        RECT 80.400 760.050 81.600 762.000 ;
        RECT 49.950 757.950 52.050 760.050 ;
        RECT 52.950 757.950 55.050 760.050 ;
        RECT 55.950 757.950 58.050 760.050 ;
        RECT 58.950 757.950 61.050 760.050 ;
        RECT 64.950 757.950 67.050 760.050 ;
        RECT 73.950 757.950 76.050 760.050 ;
        RECT 76.950 757.950 79.050 760.050 ;
        RECT 79.950 757.950 82.050 760.050 ;
        RECT 50.400 757.050 51.600 757.950 ;
        RECT 43.950 754.950 46.050 757.050 ;
        RECT 46.950 755.400 51.600 757.050 ;
        RECT 46.950 754.950 51.000 755.400 ;
        RECT 56.400 730.200 57.600 757.950 ;
        RECT 65.400 733.050 66.600 757.950 ;
        RECT 77.400 736.050 78.600 757.950 ;
        RECT 86.400 751.050 87.600 763.950 ;
        RECT 88.950 760.950 91.050 763.050 ;
        RECT 97.950 761.100 100.050 763.200 ;
        RECT 85.950 748.950 88.050 751.050 ;
        RECT 79.950 739.950 82.050 742.050 ;
        RECT 76.950 733.950 79.050 736.050 ;
        RECT 64.950 730.950 67.050 733.050 ;
        RECT 55.950 728.100 58.050 730.200 ;
        RECT 56.400 727.050 57.600 728.100 ;
        RECT 61.950 727.950 64.050 730.050 ;
        RECT 52.950 724.950 55.050 727.050 ;
        RECT 55.950 724.950 58.050 727.050 ;
        RECT 34.950 721.800 37.050 723.900 ;
        RECT 40.950 721.950 43.050 724.050 ;
        RECT 49.950 721.950 52.050 724.050 ;
        RECT 43.950 697.950 46.050 700.050 ;
        RECT 44.400 688.050 45.600 697.950 ;
        RECT 46.950 691.950 49.050 694.050 ;
        RECT 22.950 685.950 25.050 688.050 ;
        RECT 43.950 685.950 46.050 688.050 ;
        RECT 28.950 683.100 31.050 685.200 ;
        RECT 37.950 683.100 40.050 685.200 ;
        RECT 47.400 685.050 48.600 691.950 ;
        RECT 45.000 684.600 49.050 685.050 ;
        RECT 13.950 679.950 16.050 682.050 ;
        RECT 16.950 679.950 19.050 682.050 ;
        RECT 19.950 679.950 22.050 682.050 ;
        RECT 22.950 679.950 25.050 682.050 ;
        RECT 17.400 658.050 18.600 679.950 ;
        RECT 23.400 678.900 24.600 679.950 ;
        RECT 29.400 679.050 30.600 683.100 ;
        RECT 38.400 682.050 39.600 683.100 ;
        RECT 44.400 682.950 49.050 684.600 ;
        RECT 44.400 682.050 45.600 682.950 ;
        RECT 34.950 679.950 37.050 682.050 ;
        RECT 37.950 679.950 40.050 682.050 ;
        RECT 40.950 679.950 43.050 682.050 ;
        RECT 43.950 679.950 46.050 682.050 ;
        RECT 35.400 679.050 36.600 679.950 ;
        RECT 22.950 676.800 25.050 678.900 ;
        RECT 28.950 676.950 31.050 679.050 ;
        RECT 31.950 677.400 36.600 679.050 ;
        RECT 31.950 676.950 36.000 677.400 ;
        RECT 7.950 655.950 10.050 658.050 ;
        RECT 13.950 655.950 16.050 658.050 ;
        RECT 16.950 655.950 19.050 658.050 ;
        RECT 14.400 649.050 15.600 655.950 ;
        RECT 19.950 650.100 22.050 652.200 ;
        RECT 23.400 652.050 24.600 676.800 ;
        RECT 28.950 667.950 31.050 670.050 ;
        RECT 25.950 655.950 28.050 658.050 ;
        RECT 20.400 649.050 21.600 650.100 ;
        RECT 22.950 649.950 25.050 652.050 ;
        RECT 13.950 646.950 16.050 649.050 ;
        RECT 16.950 646.950 19.050 649.050 ;
        RECT 19.950 646.950 22.050 649.050 ;
        RECT 17.400 640.050 18.600 646.950 ;
        RECT 16.950 637.950 19.050 640.050 ;
        RECT 7.950 628.950 10.050 631.050 ;
        RECT 22.950 628.950 25.050 631.050 ;
        RECT 8.400 562.050 9.600 628.950 ;
        RECT 13.950 619.950 16.050 622.050 ;
        RECT 14.400 604.050 15.600 619.950 ;
        RECT 23.400 610.050 24.600 628.950 ;
        RECT 22.950 607.950 25.050 610.050 ;
        RECT 23.400 604.050 24.600 607.950 ;
        RECT 26.400 607.050 27.600 655.950 ;
        RECT 29.400 652.050 30.600 667.950 ;
        RECT 31.950 655.950 34.050 658.050 ;
        RECT 28.950 649.950 31.050 652.050 ;
        RECT 32.400 649.050 33.600 655.950 ;
        RECT 31.950 646.950 34.050 649.050 ;
        RECT 34.950 646.950 37.050 649.050 ;
        RECT 28.950 643.950 31.050 646.050 ;
        RECT 35.400 645.900 36.600 646.950 ;
        RECT 25.950 604.950 28.050 607.050 ;
        RECT 13.950 601.950 16.050 604.050 ;
        RECT 16.950 601.950 19.050 604.050 ;
        RECT 22.950 601.950 25.050 604.050 ;
        RECT 13.950 595.950 16.050 598.050 ;
        RECT 14.400 574.200 15.600 595.950 ;
        RECT 17.400 592.050 18.600 601.950 ;
        RECT 25.950 598.950 28.050 601.050 ;
        RECT 16.950 589.950 19.050 592.050 ;
        RECT 19.950 589.950 22.050 592.050 ;
        RECT 13.950 572.100 16.050 574.200 ;
        RECT 14.400 571.050 15.600 572.100 ;
        RECT 20.400 571.050 21.600 589.950 ;
        RECT 13.950 568.950 16.050 571.050 ;
        RECT 16.950 568.950 19.050 571.050 ;
        RECT 19.950 568.950 22.050 571.050 ;
        RECT 7.950 559.950 10.050 562.050 ;
        RECT 4.950 541.950 7.050 544.050 ;
        RECT 17.400 532.050 18.600 568.950 ;
        RECT 26.400 541.050 27.600 598.950 ;
        RECT 29.400 595.050 30.600 643.950 ;
        RECT 34.950 643.800 37.050 645.900 ;
        RECT 31.950 634.950 34.050 637.050 ;
        RECT 32.400 601.050 33.600 634.950 ;
        RECT 41.400 625.050 42.600 679.950 ;
        RECT 43.950 673.950 46.050 676.050 ;
        RECT 44.400 645.900 45.600 673.950 ;
        RECT 50.400 670.050 51.600 721.950 ;
        RECT 53.400 700.050 54.600 724.950 ;
        RECT 52.950 697.950 55.050 700.050 ;
        RECT 62.400 690.600 63.600 727.950 ;
        RECT 65.400 694.050 66.600 730.950 ;
        RECT 73.950 729.000 76.050 733.050 ;
        RECT 74.400 727.050 75.600 729.000 ;
        RECT 80.400 727.050 81.600 739.950 ;
        RECT 85.950 733.950 88.050 736.050 ;
        RECT 70.950 724.950 73.050 727.050 ;
        RECT 73.950 724.950 76.050 727.050 ;
        RECT 76.950 724.950 79.050 727.050 ;
        RECT 79.950 724.950 82.050 727.050 ;
        RECT 71.400 723.000 72.600 724.950 ;
        RECT 70.950 718.950 73.050 723.000 ;
        RECT 77.400 720.600 78.600 724.950 ;
        RECT 77.400 719.400 81.600 720.600 ;
        RECT 64.950 691.950 67.050 694.050 ;
        RECT 76.950 691.950 79.050 694.050 ;
        RECT 59.400 689.400 63.600 690.600 ;
        RECT 52.950 685.950 55.050 688.050 ;
        RECT 49.950 667.950 52.050 670.050 ;
        RECT 53.400 658.050 54.600 685.950 ;
        RECT 59.400 685.050 60.600 689.400 ;
        RECT 55.950 682.950 58.050 685.050 ;
        RECT 58.950 682.950 61.050 685.050 ;
        RECT 61.950 684.000 64.050 688.050 ;
        RECT 72.000 684.600 76.050 685.050 ;
        RECT 56.400 673.050 57.600 682.950 ;
        RECT 62.400 682.050 63.600 684.000 ;
        RECT 71.400 682.950 76.050 684.600 ;
        RECT 71.400 682.050 72.600 682.950 ;
        RECT 61.950 679.950 64.050 682.050 ;
        RECT 64.950 679.950 67.050 682.050 ;
        RECT 70.950 679.950 73.050 682.050 ;
        RECT 58.950 676.950 61.050 679.050 ;
        RECT 55.950 670.950 58.050 673.050 ;
        RECT 55.950 661.950 58.050 664.050 ;
        RECT 52.950 655.950 55.050 658.050 ;
        RECT 49.950 650.100 52.050 652.200 ;
        RECT 50.400 649.050 51.600 650.100 ;
        RECT 56.400 649.050 57.600 661.950 ;
        RECT 59.400 658.050 60.600 676.950 ;
        RECT 65.400 673.050 66.600 679.950 ;
        RECT 67.950 676.950 70.050 679.050 ;
        RECT 64.950 670.950 67.050 673.050 ;
        RECT 58.950 655.950 61.050 658.050 ;
        RECT 64.950 655.950 67.050 658.050 ;
        RECT 49.950 646.950 52.050 649.050 ;
        RECT 52.950 646.950 55.050 649.050 ;
        RECT 55.950 646.950 58.050 649.050 ;
        RECT 58.950 646.950 61.050 649.050 ;
        RECT 53.400 645.900 54.600 646.950 ;
        RECT 43.950 643.800 46.050 645.900 ;
        RECT 52.950 643.800 55.050 645.900 ;
        RECT 59.400 645.600 60.600 646.950 ;
        RECT 65.400 645.900 66.600 655.950 ;
        RECT 59.400 644.400 63.600 645.600 ;
        RECT 58.950 640.950 61.050 643.050 ;
        RECT 40.950 622.950 43.050 625.050 ;
        RECT 40.800 610.500 42.900 612.600 ;
        RECT 40.950 603.900 41.850 610.500 ;
        RECT 49.800 610.200 51.900 612.300 ;
        RECT 44.400 606.900 45.600 609.450 ;
        RECT 43.500 604.800 45.600 606.900 ;
        RECT 47.700 603.900 49.800 604.200 ;
        RECT 37.950 601.800 40.050 603.900 ;
        RECT 40.950 603.000 49.800 603.900 ;
        RECT 31.950 598.950 34.050 601.050 ;
        RECT 38.400 599.400 39.600 601.800 ;
        RECT 40.950 597.900 41.850 603.000 ;
        RECT 47.700 602.100 49.800 603.000 ;
        RECT 42.750 601.200 44.850 602.100 ;
        RECT 42.750 600.000 49.800 601.200 ;
        RECT 47.400 599.100 49.800 600.000 ;
        RECT 40.200 595.800 42.300 597.900 ;
        RECT 43.500 596.100 45.600 598.200 ;
        RECT 28.950 592.950 31.050 595.050 ;
        RECT 44.400 580.050 45.600 596.100 ;
        RECT 28.950 577.950 31.050 580.050 ;
        RECT 43.950 577.950 46.050 580.050 ;
        RECT 25.950 538.950 28.050 541.050 ;
        RECT 16.950 529.950 19.050 532.050 ;
        RECT 13.950 527.100 16.050 529.200 ;
        RECT 19.950 527.100 22.050 529.200 ;
        RECT 25.950 527.100 28.050 529.200 ;
        RECT 14.400 526.050 15.600 527.100 ;
        RECT 20.400 526.050 21.600 527.100 ;
        RECT 10.950 523.950 13.050 526.050 ;
        RECT 13.950 523.950 16.050 526.050 ;
        RECT 16.950 523.950 19.050 526.050 ;
        RECT 19.950 523.950 22.050 526.050 ;
        RECT 11.400 522.900 12.600 523.950 ;
        RECT 10.950 520.800 13.050 522.900 ;
        RECT 7.950 500.400 10.050 502.500 ;
        RECT 4.950 490.950 7.050 493.050 ;
        RECT 5.400 489.600 6.600 490.950 ;
        RECT 2.400 489.000 6.600 489.600 ;
        RECT 2.400 488.400 7.050 489.000 ;
        RECT 2.400 456.600 3.600 488.400 ;
        RECT 4.950 484.950 7.050 488.400 ;
        RECT 8.700 480.600 9.900 500.400 ;
        RECT 17.400 495.600 18.600 523.950 ;
        RECT 26.400 517.050 27.600 527.100 ;
        RECT 25.950 514.950 28.050 517.050 ;
        RECT 29.400 508.050 30.600 577.950 ;
        RECT 37.950 572.100 40.050 574.200 ;
        RECT 47.400 574.050 48.600 599.100 ;
        RECT 50.700 597.600 51.600 610.200 ;
        RECT 53.400 603.900 54.600 606.450 ;
        RECT 52.500 601.800 54.600 603.900 ;
        RECT 55.950 601.950 58.050 604.050 ;
        RECT 50.250 595.500 52.350 597.600 ;
        RECT 56.400 595.050 57.600 601.950 ;
        RECT 55.950 592.950 58.050 595.050 ;
        RECT 49.950 589.950 52.050 592.050 ;
        RECT 38.400 571.050 39.600 572.100 ;
        RECT 46.950 571.950 49.050 574.050 ;
        RECT 34.950 568.950 37.050 571.050 ;
        RECT 37.950 568.950 40.050 571.050 ;
        RECT 40.950 568.950 43.050 571.050 ;
        RECT 35.400 567.900 36.600 568.950 ;
        RECT 41.400 567.900 42.600 568.950 ;
        RECT 46.950 568.800 49.050 570.900 ;
        RECT 34.950 565.800 37.050 567.900 ;
        RECT 40.950 565.800 43.050 567.900 ;
        RECT 47.400 565.050 48.600 568.800 ;
        RECT 50.400 567.900 51.600 589.950 ;
        RECT 59.400 586.050 60.600 640.950 ;
        RECT 62.400 610.050 63.600 644.400 ;
        RECT 64.950 643.800 67.050 645.900 ;
        RECT 68.400 637.050 69.600 676.950 ;
        RECT 70.950 667.950 73.050 670.050 ;
        RECT 71.400 643.050 72.600 667.950 ;
        RECT 77.400 658.050 78.600 691.950 ;
        RECT 80.400 679.050 81.600 719.400 ;
        RECT 86.400 684.600 87.600 733.950 ;
        RECT 89.400 691.050 90.600 760.950 ;
        RECT 98.400 760.050 99.600 761.100 ;
        RECT 94.950 757.950 97.050 760.050 ;
        RECT 97.950 757.950 100.050 760.050 ;
        RECT 100.950 757.950 103.050 760.050 ;
        RECT 95.400 756.900 96.600 757.950 ;
        RECT 94.950 754.800 97.050 756.900 ;
        RECT 95.400 742.050 96.600 754.800 ;
        RECT 94.950 739.950 97.050 742.050 ;
        RECT 101.400 739.050 102.600 757.950 ;
        RECT 107.400 757.050 108.600 800.400 ;
        RECT 112.950 799.800 115.050 801.900 ;
        RECT 119.400 781.050 120.600 830.400 ;
        RECT 128.400 823.050 129.600 835.950 ;
        RECT 134.400 826.050 135.600 841.950 ;
        RECT 142.950 839.100 145.050 841.200 ;
        RECT 143.400 838.050 144.600 839.100 ;
        RECT 149.400 838.050 150.600 847.950 ;
        RECT 152.400 847.050 153.600 853.950 ;
        RECT 170.400 853.050 171.600 878.100 ;
        RECT 174.150 874.500 175.050 881.100 ;
        RECT 182.400 880.050 183.600 883.950 ;
        RECT 197.400 883.050 198.600 889.950 ;
        RECT 217.950 884.100 220.050 886.200 ;
        RECT 218.400 883.050 219.600 884.100 ;
        RECT 193.950 880.950 196.050 883.050 ;
        RECT 196.950 880.950 199.050 883.050 ;
        RECT 199.950 880.950 202.050 883.050 ;
        RECT 214.950 880.950 217.050 883.050 ;
        RECT 217.950 880.950 220.050 883.050 ;
        RECT 220.950 880.950 223.050 883.050 ;
        RECT 181.950 877.950 184.050 880.050 ;
        RECT 173.100 872.400 175.200 874.500 ;
        RECT 194.400 868.050 195.600 880.950 ;
        RECT 200.400 874.050 201.600 880.950 ;
        RECT 215.400 879.900 216.600 880.950 ;
        RECT 214.950 877.800 217.050 879.900 ;
        RECT 199.950 871.950 202.050 874.050 ;
        RECT 172.950 865.950 175.050 868.050 ;
        RECT 193.950 865.950 196.050 868.050 ;
        RECT 160.950 850.950 163.050 853.050 ;
        RECT 169.950 850.950 172.050 853.050 ;
        RECT 151.950 844.950 154.050 847.050 ;
        RECT 142.950 835.950 145.050 838.050 ;
        RECT 145.950 835.950 148.050 838.050 ;
        RECT 148.950 835.950 151.050 838.050 ;
        RECT 146.400 834.000 147.600 835.950 ;
        RECT 145.950 829.950 148.050 834.000 ;
        RECT 148.950 826.950 151.050 829.050 ;
        RECT 133.950 823.950 136.050 826.050 ;
        RECT 127.950 820.950 130.050 823.050 ;
        RECT 127.950 811.950 130.050 814.050 ;
        RECT 128.400 808.200 129.600 811.950 ;
        RECT 127.950 806.100 130.050 808.200 ;
        RECT 133.950 806.100 136.050 808.200 ;
        RECT 142.950 806.100 145.050 808.200 ;
        RECT 128.400 805.050 129.600 806.100 ;
        RECT 134.400 805.050 135.600 806.100 ;
        RECT 127.950 802.950 130.050 805.050 ;
        RECT 130.950 802.950 133.050 805.050 ;
        RECT 133.950 802.950 136.050 805.050 ;
        RECT 136.950 802.950 139.050 805.050 ;
        RECT 131.400 801.900 132.600 802.950 ;
        RECT 130.950 799.800 133.050 801.900 ;
        RECT 127.950 793.950 130.050 796.050 ;
        RECT 118.950 778.950 121.050 781.050 ;
        RECT 109.950 766.950 112.050 769.050 ;
        RECT 106.950 754.950 109.050 757.050 ;
        RECT 110.400 741.600 111.600 766.950 ;
        RECT 118.950 761.100 121.050 763.200 ;
        RECT 119.400 760.050 120.600 761.100 ;
        RECT 115.950 757.950 118.050 760.050 ;
        RECT 118.950 757.950 121.050 760.050 ;
        RECT 121.950 757.950 124.050 760.050 ;
        RECT 116.400 756.900 117.600 757.950 ;
        RECT 115.950 754.800 118.050 756.900 ;
        RECT 122.400 751.050 123.600 757.950 ;
        RECT 121.950 748.950 124.050 751.050 ;
        RECT 128.400 748.050 129.600 793.950 ;
        RECT 131.400 757.050 132.600 799.800 ;
        RECT 137.400 796.050 138.600 802.950 ;
        RECT 136.950 793.950 139.050 796.050 ;
        RECT 143.400 793.050 144.600 806.100 ;
        RECT 149.400 802.050 150.600 826.950 ;
        RECT 157.950 807.000 160.050 811.050 ;
        RECT 161.400 807.600 162.600 850.950 ;
        RECT 166.950 839.100 169.050 841.200 ;
        RECT 167.400 838.050 168.600 839.100 ;
        RECT 173.400 838.050 174.600 865.950 ;
        RECT 200.400 841.200 201.600 871.950 ;
        RECT 221.400 856.050 222.600 880.950 ;
        RECT 227.400 879.900 228.600 889.950 ;
        RECT 229.950 883.950 232.050 886.050 ;
        RECT 238.950 884.100 241.050 886.200 ;
        RECT 226.950 877.800 229.050 879.900 ;
        RECT 230.400 874.050 231.600 883.950 ;
        RECT 239.400 883.050 240.600 884.100 ;
        RECT 245.400 883.050 246.600 889.950 ;
        RECT 235.950 880.950 238.050 883.050 ;
        RECT 238.950 880.950 241.050 883.050 ;
        RECT 241.950 880.950 244.050 883.050 ;
        RECT 244.950 880.950 247.050 883.050 ;
        RECT 247.950 880.950 250.050 883.050 ;
        RECT 229.950 871.950 232.050 874.050 ;
        RECT 236.400 868.050 237.600 880.950 ;
        RECT 242.400 874.050 243.600 880.950 ;
        RECT 241.950 871.950 244.050 874.050 ;
        RECT 226.950 865.950 229.050 868.050 ;
        RECT 235.950 865.950 238.050 868.050 ;
        RECT 220.950 853.950 223.050 856.050 ;
        RECT 223.950 850.950 226.050 853.050 ;
        RECT 224.400 847.050 225.600 850.950 ;
        RECT 223.950 844.950 226.050 847.050 ;
        RECT 193.950 839.100 196.050 841.200 ;
        RECT 199.950 839.100 202.050 841.200 ;
        RECT 211.950 839.100 214.050 841.200 ;
        RECT 217.950 839.100 220.050 841.200 ;
        RECT 194.400 838.050 195.600 839.100 ;
        RECT 200.400 838.050 201.600 839.100 ;
        RECT 212.400 838.050 213.600 839.100 ;
        RECT 218.400 838.050 219.600 839.100 ;
        RECT 166.950 835.950 169.050 838.050 ;
        RECT 169.950 835.950 172.050 838.050 ;
        RECT 172.950 835.950 175.050 838.050 ;
        RECT 184.950 835.950 187.050 838.050 ;
        RECT 190.950 835.950 193.050 838.050 ;
        RECT 193.950 835.950 196.050 838.050 ;
        RECT 196.950 835.950 199.050 838.050 ;
        RECT 199.950 835.950 202.050 838.050 ;
        RECT 205.950 835.950 208.050 838.050 ;
        RECT 211.950 835.950 214.050 838.050 ;
        RECT 214.950 835.950 217.050 838.050 ;
        RECT 217.950 835.950 220.050 838.050 ;
        RECT 220.950 835.950 223.050 838.050 ;
        RECT 170.400 826.050 171.600 835.950 ;
        RECT 185.400 829.050 186.600 835.950 ;
        RECT 184.950 826.950 187.050 829.050 ;
        RECT 169.950 823.950 172.050 826.050 ;
        RECT 191.400 823.050 192.600 835.950 ;
        RECT 197.400 834.900 198.600 835.950 ;
        RECT 196.950 832.800 199.050 834.900 ;
        RECT 206.400 829.050 207.600 835.950 ;
        RECT 215.400 834.900 216.600 835.950 ;
        RECT 221.400 834.900 222.600 835.950 ;
        RECT 227.400 835.050 228.600 865.950 ;
        RECT 248.400 856.050 249.600 880.950 ;
        RECT 247.950 853.950 250.050 856.050 ;
        RECT 253.950 841.950 256.050 844.050 ;
        RECT 229.950 839.100 232.050 841.200 ;
        RECT 235.950 839.100 238.050 841.200 ;
        RECT 241.950 839.100 244.050 841.200 ;
        RECT 250.950 839.100 253.050 841.200 ;
        RECT 214.950 832.800 217.050 834.900 ;
        RECT 220.950 832.800 223.050 834.900 ;
        RECT 226.950 832.950 229.050 835.050 ;
        RECT 230.400 834.600 231.600 839.100 ;
        RECT 236.400 838.050 237.600 839.100 ;
        RECT 242.400 838.050 243.600 839.100 ;
        RECT 235.950 835.950 238.050 838.050 ;
        RECT 238.950 835.950 241.050 838.050 ;
        RECT 241.950 835.950 244.050 838.050 ;
        RECT 244.950 835.950 247.050 838.050 ;
        RECT 230.400 833.400 234.600 834.600 ;
        RECT 239.400 834.000 240.600 835.950 ;
        RECT 245.400 834.900 246.600 835.950 ;
        RECT 215.400 829.050 216.600 832.800 ;
        RECT 229.950 829.950 232.050 832.050 ;
        RECT 205.950 826.950 208.050 829.050 ;
        RECT 214.950 826.950 217.050 829.050 ;
        RECT 190.950 820.950 193.050 823.050 ;
        RECT 184.950 808.950 187.050 811.050 ;
        RECT 158.400 805.050 159.600 807.000 ;
        RECT 161.400 806.400 165.600 807.600 ;
        RECT 154.950 802.950 157.050 805.050 ;
        RECT 157.950 802.950 160.050 805.050 ;
        RECT 148.950 799.950 151.050 802.050 ;
        RECT 155.400 801.900 156.600 802.950 ;
        RECT 154.950 799.800 157.050 801.900 ;
        RECT 142.950 790.950 145.050 793.050 ;
        RECT 164.400 769.050 165.600 806.400 ;
        RECT 166.950 805.950 169.050 808.050 ;
        RECT 175.950 806.100 178.050 808.200 ;
        RECT 167.400 772.050 168.600 805.950 ;
        RECT 176.400 805.050 177.600 806.100 ;
        RECT 172.950 802.950 175.050 805.050 ;
        RECT 175.950 802.950 178.050 805.050 ;
        RECT 178.950 802.950 181.050 805.050 ;
        RECT 173.400 790.050 174.600 802.950 ;
        RECT 179.400 801.900 180.600 802.950 ;
        RECT 178.950 799.800 181.050 801.900 ;
        RECT 172.950 787.950 175.050 790.050 ;
        RECT 166.950 769.950 169.050 772.050 ;
        RECT 151.950 766.950 154.050 769.050 ;
        RECT 163.950 766.950 166.050 769.050 ;
        RECT 139.950 761.100 142.050 763.200 ;
        RECT 140.400 760.050 141.600 761.100 ;
        RECT 148.950 760.950 151.050 763.050 ;
        RECT 136.950 757.950 139.050 760.050 ;
        RECT 139.950 757.950 142.050 760.050 ;
        RECT 142.950 757.950 145.050 760.050 ;
        RECT 130.950 754.950 133.050 757.050 ;
        RECT 137.400 756.900 138.600 757.950 ;
        RECT 143.400 756.900 144.600 757.950 ;
        RECT 136.950 754.800 139.050 756.900 ;
        RECT 142.950 754.800 145.050 756.900 ;
        RECT 127.950 745.950 130.050 748.050 ;
        RECT 142.950 745.950 145.050 748.050 ;
        RECT 110.400 740.400 114.600 741.600 ;
        RECT 97.950 736.950 100.050 739.050 ;
        RECT 100.950 736.950 103.050 739.050 ;
        RECT 98.400 727.050 99.600 736.950 ;
        RECT 106.950 734.400 109.050 736.500 ;
        RECT 103.950 728.400 106.050 730.500 ;
        RECT 104.400 727.050 105.600 728.400 ;
        RECT 94.950 724.950 97.050 727.050 ;
        RECT 97.950 724.950 100.050 727.050 ;
        RECT 103.950 724.950 106.050 727.050 ;
        RECT 95.400 723.000 96.600 724.950 ;
        RECT 94.950 718.950 97.050 723.000 ;
        RECT 107.850 719.400 109.050 734.400 ;
        RECT 106.950 717.300 109.050 719.400 ;
        RECT 113.400 718.050 114.600 740.400 ;
        RECT 115.950 733.950 118.050 736.050 ;
        RECT 127.950 734.400 130.050 736.500 ;
        RECT 116.400 724.050 117.600 733.950 ;
        RECT 121.950 724.950 124.050 727.050 ;
        RECT 115.950 721.950 118.050 724.050 ;
        RECT 122.400 723.600 123.600 724.950 ;
        RECT 121.950 721.500 124.050 723.600 ;
        RECT 107.850 713.700 109.050 717.300 ;
        RECT 112.950 715.950 115.050 718.050 ;
        RECT 121.950 715.950 124.050 718.050 ;
        RECT 106.950 711.600 109.050 713.700 ;
        RECT 88.950 688.950 91.050 691.050 ;
        RECT 103.950 688.950 106.050 691.050 ;
        RECT 83.400 683.400 87.600 684.600 ;
        RECT 79.950 676.950 82.050 679.050 ;
        RECT 76.950 655.950 79.050 658.050 ;
        RECT 83.400 655.200 84.600 683.400 ;
        RECT 88.950 683.100 91.050 685.200 ;
        RECT 97.950 683.100 100.050 685.200 ;
        RECT 89.400 682.050 90.600 683.100 ;
        RECT 98.400 682.050 99.600 683.100 ;
        RECT 88.950 679.950 91.050 682.050 ;
        RECT 94.950 679.950 97.050 682.050 ;
        RECT 97.950 679.950 100.050 682.050 ;
        RECT 95.400 678.000 96.600 679.950 ;
        RECT 94.950 673.950 97.050 678.000 ;
        RECT 76.950 651.000 79.050 654.900 ;
        RECT 82.950 653.100 85.050 655.200 ;
        RECT 104.400 655.050 105.600 688.950 ;
        RECT 109.950 683.100 112.050 685.200 ;
        RECT 115.950 683.100 118.050 685.200 ;
        RECT 110.400 682.050 111.600 683.100 ;
        RECT 116.400 682.050 117.600 683.100 ;
        RECT 109.950 679.950 112.050 682.050 ;
        RECT 112.950 679.950 115.050 682.050 ;
        RECT 115.950 679.950 118.050 682.050 ;
        RECT 113.400 673.050 114.600 679.950 ;
        RECT 118.950 676.950 121.050 679.050 ;
        RECT 112.950 670.950 115.050 673.050 ;
        RECT 119.400 670.050 120.600 676.950 ;
        RECT 118.950 667.950 121.050 670.050 ;
        RECT 106.950 658.950 109.050 661.050 ;
        RECT 115.950 658.950 118.050 661.050 ;
        RECT 88.950 652.950 91.050 655.050 ;
        RECT 103.950 652.950 106.050 655.050 ;
        RECT 77.400 649.050 78.600 651.000 ;
        RECT 82.950 649.950 85.050 652.050 ;
        RECT 83.400 649.050 84.600 649.950 ;
        RECT 76.950 646.950 79.050 649.050 ;
        RECT 79.950 646.950 82.050 649.050 ;
        RECT 82.950 646.950 85.050 649.050 ;
        RECT 70.950 640.950 73.050 643.050 ;
        RECT 67.950 634.950 70.050 637.050 ;
        RECT 80.400 616.050 81.600 646.950 ;
        RECT 85.950 622.950 88.050 625.050 ;
        RECT 86.400 619.050 87.600 622.950 ;
        RECT 85.950 616.950 88.050 619.050 ;
        RECT 79.950 613.950 82.050 616.050 ;
        RECT 85.950 613.800 88.050 615.900 ;
        RECT 70.500 610.500 72.600 612.600 ;
        RECT 61.950 607.950 64.050 610.050 ;
        RECT 58.950 583.950 61.050 586.050 ;
        RECT 62.400 577.200 63.600 607.950 ;
        RECT 67.950 601.950 70.050 604.050 ;
        RECT 70.950 603.300 72.000 610.500 ;
        RECT 74.400 606.900 75.600 609.450 ;
        RECT 80.100 609.300 82.200 611.400 ;
        RECT 73.800 604.800 75.900 606.900 ;
        RECT 76.800 605.700 78.900 607.800 ;
        RECT 76.800 603.300 77.700 605.700 ;
        RECT 70.950 602.100 77.700 603.300 ;
        RECT 68.400 599.400 69.600 601.950 ;
        RECT 70.950 596.700 71.850 602.100 ;
        RECT 72.750 600.300 74.850 601.200 ;
        RECT 80.400 600.300 81.300 609.300 ;
        RECT 83.400 604.050 84.600 606.600 ;
        RECT 82.500 601.950 84.600 604.050 ;
        RECT 72.750 599.100 81.300 600.300 ;
        RECT 70.500 594.600 72.600 596.700 ;
        RECT 73.800 596.100 75.900 598.200 ;
        RECT 77.700 597.300 79.800 599.100 ;
        RECT 74.400 594.000 75.600 596.100 ;
        RECT 73.950 589.950 76.050 594.000 ;
        RECT 79.950 586.950 82.050 589.050 ;
        RECT 52.950 574.950 55.050 577.050 ;
        RECT 61.950 575.100 64.050 577.200 ;
        RECT 49.950 565.800 52.050 567.900 ;
        RECT 46.950 562.950 49.050 565.050 ;
        RECT 47.400 556.050 48.600 562.950 ;
        RECT 37.950 553.950 40.050 556.050 ;
        RECT 46.950 553.950 49.050 556.050 ;
        RECT 38.400 526.050 39.600 553.950 ;
        RECT 53.400 553.050 54.600 574.950 ;
        RECT 61.950 571.950 64.050 574.050 ;
        RECT 67.950 572.100 70.050 574.200 ;
        RECT 62.400 571.050 63.600 571.950 ;
        RECT 68.400 571.050 69.600 572.100 ;
        RECT 80.400 571.050 81.600 586.950 ;
        RECT 83.400 583.050 84.600 601.950 ;
        RECT 86.400 589.050 87.600 613.800 ;
        RECT 85.950 586.950 88.050 589.050 ;
        RECT 82.950 580.950 85.050 583.050 ;
        RECT 85.950 577.950 88.050 580.050 ;
        RECT 86.400 571.050 87.600 577.950 ;
        RECT 89.400 577.050 90.600 652.950 ;
        RECT 91.950 650.100 94.050 652.200 ;
        RECT 100.950 650.100 103.050 652.200 ;
        RECT 92.400 622.050 93.600 650.100 ;
        RECT 101.400 649.050 102.600 650.100 ;
        RECT 107.400 649.050 108.600 658.950 ;
        RECT 112.950 652.950 115.050 655.050 ;
        RECT 97.950 646.950 100.050 649.050 ;
        RECT 100.950 646.950 103.050 649.050 ;
        RECT 103.950 646.950 106.050 649.050 ;
        RECT 106.950 646.950 109.050 649.050 ;
        RECT 98.400 640.050 99.600 646.950 ;
        RECT 104.400 645.900 105.600 646.950 ;
        RECT 103.950 643.800 106.050 645.900 ;
        RECT 97.950 637.950 100.050 640.050 ;
        RECT 94.950 628.950 97.050 631.050 ;
        RECT 91.950 619.950 94.050 622.050 ;
        RECT 92.400 607.050 93.600 619.950 ;
        RECT 95.400 619.050 96.600 628.950 ;
        RECT 94.950 616.950 97.050 619.050 ;
        RECT 91.950 604.950 94.050 607.050 ;
        RECT 94.950 606.000 97.050 610.050 ;
        RECT 95.400 604.050 96.600 606.000 ;
        RECT 100.950 605.100 103.050 607.200 ;
        RECT 109.950 605.100 112.050 607.200 ;
        RECT 101.400 604.050 102.600 605.100 ;
        RECT 94.950 601.950 97.050 604.050 ;
        RECT 97.950 601.950 100.050 604.050 ;
        RECT 100.950 601.950 103.050 604.050 ;
        RECT 103.950 601.950 106.050 604.050 ;
        RECT 98.400 600.900 99.600 601.950 ;
        RECT 104.400 600.900 105.600 601.950 ;
        RECT 97.950 598.800 100.050 600.900 ;
        RECT 103.950 598.800 106.050 600.900 ;
        RECT 103.950 592.950 106.050 595.050 ;
        RECT 100.950 580.950 103.050 583.050 ;
        RECT 97.950 577.950 100.050 580.050 ;
        RECT 88.950 574.950 91.050 577.050 ;
        RECT 94.950 574.950 97.050 577.050 ;
        RECT 58.950 568.950 61.050 571.050 ;
        RECT 61.950 568.950 64.050 571.050 ;
        RECT 64.950 568.950 67.050 571.050 ;
        RECT 67.950 568.950 70.050 571.050 ;
        RECT 79.950 568.950 82.050 571.050 ;
        RECT 82.950 568.950 85.050 571.050 ;
        RECT 85.950 568.950 88.050 571.050 ;
        RECT 88.950 568.950 91.050 571.050 ;
        RECT 55.950 565.800 58.050 567.900 ;
        RECT 59.400 567.000 60.600 568.950 ;
        RECT 65.400 567.900 66.600 568.950 ;
        RECT 56.400 562.050 57.600 565.800 ;
        RECT 58.950 562.950 61.050 567.000 ;
        RECT 64.950 565.800 67.050 567.900 ;
        RECT 55.950 559.950 58.050 562.050 ;
        RECT 43.950 550.950 46.050 553.050 ;
        RECT 52.950 550.950 55.050 553.050 ;
        RECT 44.400 526.050 45.600 550.950 ;
        RECT 52.950 547.800 55.050 549.900 ;
        RECT 53.400 526.050 54.600 547.800 ;
        RECT 83.400 544.050 84.600 568.950 ;
        RECT 82.950 541.950 85.050 544.050 ;
        RECT 76.950 538.950 79.050 541.050 ;
        RECT 61.500 532.500 63.600 534.600 ;
        RECT 37.950 523.950 40.050 526.050 ;
        RECT 40.950 523.950 43.050 526.050 ;
        RECT 43.950 523.950 46.050 526.050 ;
        RECT 52.950 523.950 55.050 526.050 ;
        RECT 58.950 523.950 61.050 526.050 ;
        RECT 61.950 525.300 63.000 532.500 ;
        RECT 65.400 528.900 66.600 531.450 ;
        RECT 71.100 531.300 73.200 533.400 ;
        RECT 64.800 526.800 66.900 528.900 ;
        RECT 67.800 527.700 69.900 529.800 ;
        RECT 67.800 525.300 68.700 527.700 ;
        RECT 61.950 524.100 68.700 525.300 ;
        RECT 41.400 522.900 42.600 523.950 ;
        RECT 40.950 520.800 43.050 522.900 ;
        RECT 59.400 521.400 60.600 523.950 ;
        RECT 61.950 518.700 62.850 524.100 ;
        RECT 63.750 522.300 65.850 523.200 ;
        RECT 71.400 522.300 72.300 531.300 ;
        RECT 77.400 529.050 78.600 538.950 ;
        RECT 82.950 537.300 85.050 539.400 ;
        RECT 89.400 538.050 90.600 568.950 ;
        RECT 95.400 567.600 96.600 574.950 ;
        RECT 92.400 566.400 96.600 567.600 ;
        RECT 83.850 533.700 85.050 537.300 ;
        RECT 88.950 535.950 91.050 538.050 ;
        RECT 92.400 535.050 93.600 566.400 ;
        RECT 94.950 562.950 97.050 565.050 ;
        RECT 82.950 531.600 85.050 533.700 ;
        RECT 91.950 532.950 94.050 535.050 ;
        RECT 74.400 526.050 75.600 528.600 ;
        RECT 76.950 526.950 79.050 529.050 ;
        RECT 73.500 525.900 75.600 526.050 ;
        RECT 73.500 523.950 76.050 525.900 ;
        RECT 79.950 523.950 82.050 526.050 ;
        RECT 73.950 523.800 76.050 523.950 ;
        RECT 80.400 522.600 81.600 523.950 ;
        RECT 63.750 521.100 72.300 522.300 ;
        RECT 49.950 514.950 52.050 517.050 ;
        RECT 61.500 516.600 63.600 518.700 ;
        RECT 64.800 518.100 66.900 520.200 ;
        RECT 68.700 519.300 70.800 521.100 ;
        RECT 79.950 520.500 82.050 522.600 ;
        RECT 28.950 505.950 31.050 508.050 ;
        RECT 37.950 505.950 40.050 508.050 ;
        RECT 28.950 500.400 31.050 502.500 ;
        RECT 17.400 494.400 21.600 495.600 ;
        RECT 13.950 490.950 16.050 493.050 ;
        RECT 14.400 489.600 15.600 490.950 ;
        RECT 20.400 489.600 21.600 494.400 ;
        RECT 13.950 487.500 16.050 489.600 ;
        RECT 19.950 487.500 22.050 489.600 ;
        RECT 28.950 485.400 30.150 500.400 ;
        RECT 31.950 494.400 34.050 496.500 ;
        RECT 32.400 493.050 33.600 494.400 ;
        RECT 31.950 490.950 34.050 493.050 ;
        RECT 28.950 483.300 31.050 485.400 ;
        RECT 7.950 478.500 10.050 480.600 ;
        RECT 28.950 479.700 30.150 483.300 ;
        RECT 28.950 477.600 31.050 479.700 ;
        RECT 7.950 458.400 10.050 460.500 ;
        RECT 28.950 459.300 31.050 461.400 ;
        RECT 4.950 456.600 7.050 457.050 ;
        RECT 2.400 455.400 7.050 456.600 ;
        RECT 4.950 454.950 7.050 455.400 ;
        RECT 5.400 448.050 6.600 454.950 ;
        RECT 4.950 445.950 7.050 448.050 ;
        RECT 8.700 438.600 9.900 458.400 ;
        RECT 22.950 454.950 25.050 457.050 ;
        RECT 28.950 455.700 30.150 459.300 ;
        RECT 13.950 449.400 16.050 451.500 ;
        RECT 19.950 449.400 22.050 451.500 ;
        RECT 14.400 448.050 15.600 449.400 ;
        RECT 13.950 445.950 16.050 448.050 ;
        RECT 7.950 436.500 10.050 438.600 ;
        RECT 20.400 436.050 21.600 449.400 ;
        RECT 19.950 433.950 22.050 436.050 ;
        RECT 7.950 422.400 10.050 424.500 ;
        RECT 4.950 412.950 7.050 415.050 ;
        RECT 5.400 406.050 6.600 412.950 ;
        RECT 4.950 403.950 7.050 406.050 ;
        RECT 8.700 402.600 9.900 422.400 ;
        RECT 19.950 421.950 22.050 424.050 ;
        RECT 13.950 412.950 16.050 415.050 ;
        RECT 14.400 411.600 15.600 412.950 ;
        RECT 20.400 411.600 21.600 421.950 ;
        RECT 13.950 409.500 16.050 411.600 ;
        RECT 19.950 409.500 22.050 411.600 ;
        RECT 23.400 406.050 24.600 454.950 ;
        RECT 28.950 453.600 31.050 455.700 ;
        RECT 28.950 438.600 30.150 453.600 ;
        RECT 31.950 445.950 34.050 448.050 ;
        RECT 32.400 444.600 33.600 445.950 ;
        RECT 31.950 442.500 34.050 444.600 ;
        RECT 28.950 436.500 31.050 438.600 ;
        RECT 28.950 422.400 31.050 424.500 ;
        RECT 28.950 407.400 30.150 422.400 ;
        RECT 31.950 416.400 34.050 418.500 ;
        RECT 32.400 415.050 33.600 416.400 ;
        RECT 31.950 412.950 34.050 415.050 ;
        RECT 22.950 403.950 25.050 406.050 ;
        RECT 28.950 405.300 31.050 407.400 ;
        RECT 38.400 406.050 39.600 505.950 ;
        RECT 40.950 494.400 43.050 496.500 ;
        RECT 41.400 490.050 42.600 494.400 ;
        RECT 50.400 493.050 51.600 514.950 ;
        RECT 61.950 511.950 64.050 514.050 ;
        RECT 46.950 490.950 49.050 493.050 ;
        RECT 49.950 490.950 52.050 493.050 ;
        RECT 52.950 490.950 55.050 493.050 ;
        RECT 40.950 487.950 43.050 490.050 ;
        RECT 47.400 489.900 48.600 490.950 ;
        RECT 53.400 489.900 54.600 490.950 ;
        RECT 46.950 489.600 49.050 489.900 ;
        RECT 44.400 488.400 49.050 489.600 ;
        RECT 40.950 442.500 43.050 444.600 ;
        RECT 41.400 412.050 42.600 442.500 ;
        RECT 44.400 418.050 45.600 488.400 ;
        RECT 46.950 487.800 49.050 488.400 ;
        RECT 52.950 487.800 55.050 489.900 ;
        RECT 49.950 449.100 52.050 451.200 ;
        RECT 55.950 450.000 58.050 454.050 ;
        RECT 62.400 450.600 63.600 511.950 ;
        RECT 65.400 454.050 66.600 518.100 ;
        RECT 73.950 517.800 76.050 519.900 ;
        RECT 70.950 514.950 73.050 517.050 ;
        RECT 71.400 510.600 72.600 514.950 ;
        RECT 74.400 514.050 75.600 517.800 ;
        RECT 83.850 516.600 85.050 531.600 ;
        RECT 95.400 529.050 96.600 562.950 ;
        RECT 98.400 544.050 99.600 577.950 ;
        RECT 101.400 565.050 102.600 580.950 ;
        RECT 104.400 574.050 105.600 592.950 ;
        RECT 110.400 592.050 111.600 605.100 ;
        RECT 109.950 589.950 112.050 592.050 ;
        RECT 106.950 580.950 109.050 583.050 ;
        RECT 103.950 571.950 106.050 574.050 ;
        RECT 107.400 571.050 108.600 580.950 ;
        RECT 113.400 573.600 114.600 652.950 ;
        RECT 116.400 622.050 117.600 658.950 ;
        RECT 122.400 652.050 123.600 715.950 ;
        RECT 128.100 714.600 129.300 734.400 ;
        RECT 136.950 728.400 139.050 730.500 ;
        RECT 130.950 724.950 133.050 727.050 ;
        RECT 131.400 718.050 132.600 724.950 ;
        RECT 130.950 715.950 133.050 718.050 ;
        RECT 127.950 712.500 130.050 714.600 ;
        RECT 137.400 709.050 138.600 728.400 ;
        RECT 130.950 706.950 133.050 709.050 ;
        RECT 136.950 706.950 139.050 709.050 ;
        RECT 131.400 685.200 132.600 706.950 ;
        RECT 124.950 683.100 127.050 685.200 ;
        RECT 130.950 683.100 133.050 685.200 ;
        RECT 136.950 683.100 139.050 685.200 ;
        RECT 125.400 676.050 126.600 683.100 ;
        RECT 131.400 682.050 132.600 683.100 ;
        RECT 137.400 682.050 138.600 683.100 ;
        RECT 130.950 679.950 133.050 682.050 ;
        RECT 133.950 679.950 136.050 682.050 ;
        RECT 136.950 679.950 139.050 682.050 ;
        RECT 134.400 678.900 135.600 679.950 ;
        RECT 133.950 676.800 136.050 678.900 ;
        RECT 124.950 673.950 127.050 676.050 ;
        RECT 127.950 667.950 130.050 670.050 ;
        RECT 128.400 655.050 129.600 667.950 ;
        RECT 136.950 656.400 139.050 658.500 ;
        RECT 127.950 652.950 130.050 655.050 ;
        RECT 121.950 649.950 124.050 652.050 ;
        RECT 128.400 649.050 129.600 652.950 ;
        RECT 133.950 651.000 136.050 655.050 ;
        RECT 134.400 649.050 135.600 651.000 ;
        RECT 124.950 646.950 127.050 649.050 ;
        RECT 127.950 646.950 130.050 649.050 ;
        RECT 133.950 646.950 136.050 649.050 ;
        RECT 125.400 637.050 126.600 646.950 ;
        RECT 137.850 641.400 139.050 656.400 ;
        RECT 136.950 639.300 139.050 641.400 ;
        RECT 124.950 634.950 127.050 637.050 ;
        RECT 137.850 635.700 139.050 639.300 ;
        RECT 136.950 633.600 139.050 635.700 ;
        RECT 143.400 631.050 144.600 745.950 ;
        RECT 145.950 739.950 148.050 742.050 ;
        RECT 146.400 730.050 147.600 739.950 ;
        RECT 149.400 739.050 150.600 760.950 ;
        RECT 152.400 742.050 153.600 766.950 ;
        RECT 179.400 763.200 180.600 799.800 ;
        RECT 185.400 790.050 186.600 808.950 ;
        RECT 196.950 806.100 199.050 808.200 ;
        RECT 197.400 805.050 198.600 806.100 ;
        RECT 208.950 805.950 211.050 808.050 ;
        RECT 214.950 806.100 217.050 808.200 ;
        RECT 220.950 806.100 223.050 808.200 ;
        RECT 193.950 802.950 196.050 805.050 ;
        RECT 196.950 802.950 199.050 805.050 ;
        RECT 194.400 796.050 195.600 802.950 ;
        RECT 193.950 793.950 196.050 796.050 ;
        RECT 184.950 787.950 187.050 790.050 ;
        RECT 196.950 787.950 199.050 790.050 ;
        RECT 184.950 769.950 187.050 772.050 ;
        RECT 160.950 761.100 163.050 763.200 ;
        RECT 166.950 761.100 169.050 763.200 ;
        RECT 178.950 761.100 181.050 763.200 ;
        RECT 161.400 760.050 162.600 761.100 ;
        RECT 157.950 757.950 160.050 760.050 ;
        RECT 160.950 757.950 163.050 760.050 ;
        RECT 158.400 751.050 159.600 757.950 ;
        RECT 167.400 757.050 168.600 761.100 ;
        RECT 179.400 760.050 180.600 761.100 ;
        RECT 185.400 760.050 186.600 769.950 ;
        RECT 193.950 766.950 196.050 769.050 ;
        RECT 175.950 757.950 178.050 760.050 ;
        RECT 178.950 757.950 181.050 760.050 ;
        RECT 181.950 757.950 184.050 760.050 ;
        RECT 184.950 757.950 187.050 760.050 ;
        RECT 187.950 757.950 190.050 760.050 ;
        RECT 166.950 754.950 169.050 757.050 ;
        RECT 176.400 756.900 177.600 757.950 ;
        RECT 175.950 754.800 178.050 756.900 ;
        RECT 157.950 750.600 160.050 751.050 ;
        RECT 157.950 749.400 162.600 750.600 ;
        RECT 157.950 748.950 160.050 749.400 ;
        RECT 151.950 739.950 154.050 742.050 ;
        RECT 148.950 736.950 151.050 739.050 ;
        RECT 148.950 732.600 151.050 735.900 ;
        RECT 148.950 732.000 153.600 732.600 ;
        RECT 149.400 731.400 153.600 732.000 ;
        RECT 145.950 727.950 148.050 730.050 ;
        RECT 152.400 727.050 153.600 731.400 ;
        RECT 157.950 728.100 160.050 730.200 ;
        RECT 161.400 729.600 162.600 749.400 ;
        RECT 175.950 748.950 178.050 751.050 ;
        RECT 166.950 734.400 169.050 736.500 ;
        RECT 161.400 728.400 165.600 729.600 ;
        RECT 158.400 727.050 159.600 728.100 ;
        RECT 164.400 727.050 165.600 728.400 ;
        RECT 148.950 724.950 151.050 727.050 ;
        RECT 151.950 724.950 154.050 727.050 ;
        RECT 154.950 724.950 157.050 727.050 ;
        RECT 157.950 724.950 160.050 727.050 ;
        RECT 163.950 724.950 166.050 727.050 ;
        RECT 149.400 679.050 150.600 724.950 ;
        RECT 155.400 723.900 156.600 724.950 ;
        RECT 154.950 721.800 157.050 723.900 ;
        RECT 157.950 718.950 160.050 721.050 ;
        RECT 167.850 719.400 169.050 734.400 ;
        RECT 154.950 712.950 157.050 715.050 ;
        RECT 155.400 682.050 156.600 712.950 ;
        RECT 158.400 685.050 159.600 718.950 ;
        RECT 166.950 717.300 169.050 719.400 ;
        RECT 167.850 713.700 169.050 717.300 ;
        RECT 176.400 715.050 177.600 748.950 ;
        RECT 182.400 733.050 183.600 757.950 ;
        RECT 188.400 745.050 189.600 757.950 ;
        RECT 194.400 753.600 195.600 766.950 ;
        RECT 197.400 757.050 198.600 787.950 ;
        RECT 209.400 763.200 210.600 805.950 ;
        RECT 215.400 805.050 216.600 806.100 ;
        RECT 221.400 805.050 222.600 806.100 ;
        RECT 214.950 802.950 217.050 805.050 ;
        RECT 217.950 802.950 220.050 805.050 ;
        RECT 220.950 802.950 223.050 805.050 ;
        RECT 223.950 802.950 226.050 805.050 ;
        RECT 218.400 799.050 219.600 802.950 ;
        RECT 224.400 802.050 225.600 802.950 ;
        RECT 224.400 800.400 229.050 802.050 ;
        RECT 225.000 799.950 229.050 800.400 ;
        RECT 230.400 799.050 231.600 829.950 ;
        RECT 233.400 814.050 234.600 833.400 ;
        RECT 238.950 829.950 241.050 834.000 ;
        RECT 244.950 832.800 247.050 834.900 ;
        RECT 251.400 834.600 252.600 839.100 ;
        RECT 254.400 835.050 255.600 841.950 ;
        RECT 248.400 833.400 252.600 834.600 ;
        RECT 232.950 811.950 235.050 814.050 ;
        RECT 233.400 801.600 234.600 811.950 ;
        RECT 241.950 806.100 244.050 808.200 ;
        RECT 242.400 805.050 243.600 806.100 ;
        RECT 238.950 802.950 241.050 805.050 ;
        RECT 241.950 802.950 244.050 805.050 ;
        RECT 239.400 802.050 240.600 802.950 ;
        RECT 235.950 801.600 240.600 802.050 ;
        RECT 233.400 800.400 240.600 801.600 ;
        RECT 235.950 799.950 240.000 800.400 ;
        RECT 217.950 796.950 220.050 799.050 ;
        RECT 229.950 796.950 232.050 799.050 ;
        RECT 218.400 783.600 219.600 796.950 ;
        RECT 248.400 796.050 249.600 833.400 ;
        RECT 253.950 832.950 256.050 835.050 ;
        RECT 257.400 834.600 258.600 892.950 ;
        RECT 262.950 884.100 265.050 886.200 ;
        RECT 263.400 883.050 264.600 884.100 ;
        RECT 269.400 883.050 270.600 892.950 ;
        RECT 289.950 884.100 292.050 886.200 ;
        RECT 304.950 884.100 307.050 886.200 ;
        RECT 290.400 883.050 291.600 884.100 ;
        RECT 305.400 883.050 306.600 884.100 ;
        RECT 311.400 883.050 312.600 892.950 ;
        RECT 316.950 889.950 319.050 892.050 ;
        RECT 317.400 886.050 318.600 889.950 ;
        RECT 316.950 883.950 319.050 886.050 ;
        RECT 262.950 880.950 265.050 883.050 ;
        RECT 265.950 880.950 268.050 883.050 ;
        RECT 268.950 880.950 271.050 883.050 ;
        RECT 271.950 880.950 274.050 883.050 ;
        RECT 286.950 880.950 289.050 883.050 ;
        RECT 289.950 880.950 292.050 883.050 ;
        RECT 304.950 880.950 307.050 883.050 ;
        RECT 307.950 880.950 310.050 883.050 ;
        RECT 310.950 880.950 313.050 883.050 ;
        RECT 313.950 880.950 316.050 883.050 ;
        RECT 266.400 862.050 267.600 880.950 ;
        RECT 272.400 879.900 273.600 880.950 ;
        RECT 271.950 877.800 274.050 879.900 ;
        RECT 265.950 859.950 268.050 862.050 ;
        RECT 287.400 847.050 288.600 880.950 ;
        RECT 308.400 879.900 309.600 880.950 ;
        RECT 314.400 879.900 315.600 880.950 ;
        RECT 295.950 877.800 298.050 879.900 ;
        RECT 307.950 877.800 310.050 879.900 ;
        RECT 313.950 877.800 316.050 879.900 ;
        RECT 268.950 844.950 271.050 847.050 ;
        RECT 286.800 844.950 288.900 847.050 ;
        RECT 289.950 844.950 292.050 847.050 ;
        RECT 262.950 840.000 265.050 844.050 ;
        RECT 263.400 838.050 264.600 840.000 ;
        RECT 269.400 838.050 270.600 844.950 ;
        RECT 280.950 839.100 283.050 841.200 ;
        RECT 262.950 835.950 265.050 838.050 ;
        RECT 265.950 835.950 268.050 838.050 ;
        RECT 268.950 835.950 271.050 838.050 ;
        RECT 271.950 835.950 274.050 838.050 ;
        RECT 257.400 833.400 261.600 834.600 ;
        RECT 253.950 806.100 256.050 808.200 ;
        RECT 254.400 805.050 255.600 806.100 ;
        RECT 260.400 805.050 261.600 833.400 ;
        RECT 266.400 829.050 267.600 835.950 ;
        RECT 272.400 834.900 273.600 835.950 ;
        RECT 271.950 832.800 274.050 834.900 ;
        RECT 265.950 826.950 268.050 829.050 ;
        RECT 268.950 806.100 271.050 808.200 ;
        RECT 253.950 802.950 256.050 805.050 ;
        RECT 256.950 802.950 259.050 805.050 ;
        RECT 259.950 802.950 262.050 805.050 ;
        RECT 262.950 802.950 265.050 805.050 ;
        RECT 247.950 793.950 250.050 796.050 ;
        RECT 257.400 790.050 258.600 802.950 ;
        RECT 263.400 801.900 264.600 802.950 ;
        RECT 262.950 799.800 265.050 801.900 ;
        RECT 263.400 796.050 264.600 799.800 ;
        RECT 262.950 793.950 265.050 796.050 ;
        RECT 256.950 787.950 259.050 790.050 ;
        RECT 218.400 782.400 222.600 783.600 ;
        RECT 214.950 766.950 217.050 769.050 ;
        RECT 199.950 760.950 202.050 763.050 ;
        RECT 208.950 761.100 211.050 763.200 ;
        RECT 196.950 754.950 199.050 757.050 ;
        RECT 194.400 752.400 198.600 753.600 ;
        RECT 187.950 742.950 190.050 745.050 ;
        RECT 187.950 734.400 190.050 736.500 ;
        RECT 181.950 730.950 184.050 733.050 ;
        RECT 181.950 724.950 184.050 727.050 ;
        RECT 182.400 723.600 183.600 724.950 ;
        RECT 181.950 721.500 184.050 723.600 ;
        RECT 166.950 711.600 169.050 713.700 ;
        RECT 175.950 712.950 178.050 715.050 ;
        RECT 188.100 714.600 189.300 734.400 ;
        RECT 190.950 724.950 193.050 727.050 ;
        RECT 191.400 718.050 192.600 724.950 ;
        RECT 197.400 718.050 198.600 752.400 ;
        RECT 200.400 730.200 201.600 760.950 ;
        RECT 209.400 760.050 210.600 761.100 ;
        RECT 215.400 760.050 216.600 766.950 ;
        RECT 205.950 757.950 208.050 760.050 ;
        RECT 208.950 757.950 211.050 760.050 ;
        RECT 211.950 757.950 214.050 760.050 ;
        RECT 214.950 757.950 217.050 760.050 ;
        RECT 206.400 756.900 207.600 757.950 ;
        RECT 205.950 754.800 208.050 756.900 ;
        RECT 212.400 748.050 213.600 757.950 ;
        RECT 211.950 745.950 214.050 748.050 ;
        RECT 208.950 742.950 211.050 745.050 ;
        RECT 199.950 728.100 202.050 730.200 ;
        RECT 209.400 727.050 210.600 742.950 ;
        RECT 221.400 739.050 222.600 782.400 ;
        RECT 269.400 769.050 270.600 806.100 ;
        RECT 281.400 805.050 282.600 839.100 ;
        RECT 290.400 838.050 291.600 844.950 ;
        RECT 296.400 841.200 297.600 877.800 ;
        RECT 301.950 865.950 304.050 868.050 ;
        RECT 295.950 839.100 298.050 841.200 ;
        RECT 296.400 838.050 297.600 839.100 ;
        RECT 286.950 835.950 289.050 838.050 ;
        RECT 289.950 835.950 292.050 838.050 ;
        RECT 292.950 835.950 295.050 838.050 ;
        RECT 295.950 835.950 298.050 838.050 ;
        RECT 287.400 834.900 288.600 835.950 ;
        RECT 293.400 834.900 294.600 835.950 ;
        RECT 302.400 834.900 303.600 865.950 ;
        RECT 314.400 847.050 315.600 877.800 ;
        RECT 323.400 868.050 324.600 892.950 ;
        RECT 331.950 885.000 334.050 889.050 ;
        RECT 335.400 886.050 336.600 892.950 ;
        RECT 367.950 889.950 370.050 892.050 ;
        RECT 337.950 886.950 340.050 889.050 ;
        RECT 332.400 883.050 333.600 885.000 ;
        RECT 334.950 883.950 337.050 886.050 ;
        RECT 328.950 880.950 331.050 883.050 ;
        RECT 331.950 880.950 334.050 883.050 ;
        RECT 329.400 879.900 330.600 880.950 ;
        RECT 328.950 877.800 331.050 879.900 ;
        RECT 322.950 865.950 325.050 868.050 ;
        RECT 325.950 859.950 328.050 862.050 ;
        RECT 313.950 844.950 316.050 847.050 ;
        RECT 319.950 844.950 322.050 847.050 ;
        RECT 307.950 839.100 310.050 841.200 ;
        RECT 313.950 840.000 316.050 843.900 ;
        RECT 320.400 841.050 321.600 844.950 ;
        RECT 322.950 841.950 325.050 844.050 ;
        RECT 308.400 838.050 309.600 839.100 ;
        RECT 314.400 838.050 315.600 840.000 ;
        RECT 319.950 838.950 322.050 841.050 ;
        RECT 307.950 835.950 310.050 838.050 ;
        RECT 310.950 835.950 313.050 838.050 ;
        RECT 313.950 835.950 316.050 838.050 ;
        RECT 316.950 835.950 319.050 838.050 ;
        RECT 311.400 834.900 312.600 835.950 ;
        RECT 286.950 832.800 289.050 834.900 ;
        RECT 292.950 832.800 295.050 834.900 ;
        RECT 301.950 832.800 304.050 834.900 ;
        RECT 310.950 832.800 313.050 834.900 ;
        RECT 317.400 826.050 318.600 835.950 ;
        RECT 316.950 823.950 319.050 826.050 ;
        RECT 286.950 820.950 289.050 823.050 ;
        RECT 295.950 820.950 298.050 823.050 ;
        RECT 287.400 805.050 288.600 820.950 ;
        RECT 280.950 802.950 283.050 805.050 ;
        RECT 283.950 802.950 286.050 805.050 ;
        RECT 286.950 802.950 289.050 805.050 ;
        RECT 289.950 802.950 292.050 805.050 ;
        RECT 284.400 801.000 285.600 802.950 ;
        RECT 290.400 801.900 291.600 802.950 ;
        RECT 296.400 801.900 297.600 820.950 ;
        RECT 304.950 806.100 307.050 811.050 ;
        RECT 310.950 806.100 313.050 808.200 ;
        RECT 323.400 808.050 324.600 841.950 ;
        RECT 326.400 835.050 327.600 859.950 ;
        RECT 334.950 843.600 337.050 844.050 ;
        RECT 338.400 843.600 339.600 886.950 ;
        RECT 340.950 883.950 343.050 886.050 ;
        RECT 346.950 884.100 349.050 886.200 ;
        RECT 352.950 884.100 355.050 886.200 ;
        RECT 358.950 884.100 361.050 886.200 ;
        RECT 341.400 874.050 342.600 883.950 ;
        RECT 347.400 883.050 348.600 884.100 ;
        RECT 353.400 883.050 354.600 884.100 ;
        RECT 346.950 880.950 349.050 883.050 ;
        RECT 349.950 880.950 352.050 883.050 ;
        RECT 352.950 880.950 355.050 883.050 ;
        RECT 340.950 871.950 343.050 874.050 ;
        RECT 350.400 853.050 351.600 880.950 ;
        RECT 352.950 868.950 355.050 871.050 ;
        RECT 349.950 850.950 352.050 853.050 ;
        RECT 334.950 842.400 339.600 843.600 ;
        RECT 334.950 840.000 337.050 842.400 ;
        RECT 349.950 841.950 352.050 844.050 ;
        RECT 335.400 838.050 336.600 840.000 ;
        RECT 340.950 839.100 343.050 841.200 ;
        RECT 341.400 838.050 342.600 839.100 ;
        RECT 334.950 835.950 337.050 838.050 ;
        RECT 337.950 835.950 340.050 838.050 ;
        RECT 340.950 835.950 343.050 838.050 ;
        RECT 343.950 835.950 346.050 838.050 ;
        RECT 325.950 832.950 328.050 835.050 ;
        RECT 338.400 834.900 339.600 835.950 ;
        RECT 344.400 834.900 345.600 835.950 ;
        RECT 337.950 832.800 340.050 834.900 ;
        RECT 343.950 832.800 346.050 834.900 ;
        RECT 350.400 831.600 351.600 841.950 ;
        RECT 353.400 835.050 354.600 868.950 ;
        RECT 359.400 862.050 360.600 884.100 ;
        RECT 368.400 883.050 369.600 889.950 ;
        RECT 373.950 884.100 376.050 886.200 ;
        RECT 374.400 883.050 375.600 884.100 ;
        RECT 388.950 883.950 391.050 886.050 ;
        RECT 367.950 880.950 370.050 883.050 ;
        RECT 370.950 880.950 373.050 883.050 ;
        RECT 373.950 880.950 376.050 883.050 ;
        RECT 376.950 880.950 379.050 883.050 ;
        RECT 371.400 871.050 372.600 880.950 ;
        RECT 370.950 868.950 373.050 871.050 ;
        RECT 377.400 868.050 378.600 880.950 ;
        RECT 389.400 879.900 390.600 883.950 ;
        RECT 395.400 883.050 396.600 892.950 ;
        RECT 490.950 889.950 493.050 892.050 ;
        RECT 541.950 889.950 544.050 892.050 ;
        RECT 400.950 884.100 403.050 886.200 ;
        RECT 409.950 884.100 412.050 886.200 ;
        RECT 415.950 884.100 418.050 886.200 ;
        RECT 439.950 884.100 442.050 886.200 ;
        RECT 445.950 884.100 448.050 886.200 ;
        RECT 454.950 884.100 457.050 886.200 ;
        RECT 463.950 884.100 466.050 886.200 ;
        RECT 469.950 884.100 472.050 886.200 ;
        RECT 401.400 883.050 402.600 884.100 ;
        RECT 394.950 880.950 397.050 883.050 ;
        RECT 397.950 880.950 400.050 883.050 ;
        RECT 400.950 880.950 403.050 883.050 ;
        RECT 403.950 880.950 406.050 883.050 ;
        RECT 388.950 877.800 391.050 879.900 ;
        RECT 398.400 879.000 399.600 880.950 ;
        RECT 397.950 874.950 400.050 879.000 ;
        RECT 404.400 871.050 405.600 880.950 ;
        RECT 406.950 874.950 409.050 877.050 ;
        RECT 403.950 868.950 406.050 871.050 ;
        RECT 407.400 868.050 408.600 874.950 ;
        RECT 410.400 871.050 411.600 884.100 ;
        RECT 416.400 883.050 417.600 884.100 ;
        RECT 440.400 883.050 441.600 884.100 ;
        RECT 446.400 883.050 447.600 884.100 ;
        RECT 415.950 880.950 418.050 883.050 ;
        RECT 418.950 880.950 421.050 883.050 ;
        RECT 439.950 880.950 442.050 883.050 ;
        RECT 442.950 880.950 445.050 883.050 ;
        RECT 445.950 880.950 448.050 883.050 ;
        RECT 448.950 880.950 451.050 883.050 ;
        RECT 419.400 880.050 420.600 880.950 ;
        RECT 419.400 878.400 424.050 880.050 ;
        RECT 420.000 877.950 424.050 878.400 ;
        RECT 430.950 877.950 433.050 880.050 ;
        RECT 443.400 879.900 444.600 880.950 ;
        RECT 449.400 879.900 450.600 880.950 ;
        RECT 409.950 868.950 412.050 871.050 ;
        RECT 421.950 868.950 424.050 871.050 ;
        RECT 376.950 865.950 379.050 868.050 ;
        RECT 406.950 865.950 409.050 868.050 ;
        RECT 358.950 859.950 361.050 862.050 ;
        RECT 367.950 844.950 370.050 847.050 ;
        RECT 361.950 840.000 364.050 844.050 ;
        RECT 362.400 838.050 363.600 840.000 ;
        RECT 368.400 838.050 369.600 844.950 ;
        RECT 373.950 841.950 376.050 844.050 ;
        RECT 358.950 835.950 361.050 838.050 ;
        RECT 361.950 835.950 364.050 838.050 ;
        RECT 364.950 835.950 367.050 838.050 ;
        RECT 367.950 835.950 370.050 838.050 ;
        RECT 352.950 832.950 355.050 835.050 ;
        RECT 359.400 834.900 360.600 835.950 ;
        RECT 358.950 832.800 361.050 834.900 ;
        RECT 365.400 834.000 366.600 835.950 ;
        RECT 347.400 830.400 351.600 831.600 ;
        RECT 343.950 814.950 346.050 817.050 ;
        RECT 305.400 805.050 306.600 806.100 ;
        RECT 311.400 805.050 312.600 806.100 ;
        RECT 322.950 805.950 325.050 808.050 ;
        RECT 328.950 807.000 331.050 811.050 ;
        RECT 344.400 808.200 345.600 814.950 ;
        RECT 329.400 805.050 330.600 807.000 ;
        RECT 334.950 806.100 337.050 808.200 ;
        RECT 343.950 806.100 346.050 808.200 ;
        RECT 335.400 805.050 336.600 806.100 ;
        RECT 301.950 802.950 304.050 805.050 ;
        RECT 304.950 802.950 307.050 805.050 ;
        RECT 307.950 802.950 310.050 805.050 ;
        RECT 310.950 802.950 313.050 805.050 ;
        RECT 328.950 802.950 331.050 805.050 ;
        RECT 331.950 802.950 334.050 805.050 ;
        RECT 334.950 802.950 337.050 805.050 ;
        RECT 337.950 802.950 340.050 805.050 ;
        RECT 302.400 801.900 303.600 802.950 ;
        RECT 283.950 796.950 286.050 801.000 ;
        RECT 289.950 799.800 292.050 801.900 ;
        RECT 295.950 799.800 298.050 801.900 ;
        RECT 301.950 799.800 304.050 801.900 ;
        RECT 308.400 799.050 309.600 802.950 ;
        RECT 307.950 796.950 310.050 799.050 ;
        RECT 274.950 787.950 277.050 790.050 ;
        RECT 238.950 766.950 241.050 769.050 ;
        RECT 268.950 766.950 271.050 769.050 ;
        RECT 232.950 761.100 235.050 763.200 ;
        RECT 233.400 760.050 234.600 761.100 ;
        RECT 239.400 760.050 240.600 766.950 ;
        RECT 244.950 761.100 247.050 763.200 ;
        RECT 259.950 761.100 262.050 763.200 ;
        RECT 265.950 761.100 268.050 763.200 ;
        RECT 271.950 761.100 274.050 763.200 ;
        RECT 229.950 757.950 232.050 760.050 ;
        RECT 232.950 757.950 235.050 760.050 ;
        RECT 235.950 757.950 238.050 760.050 ;
        RECT 238.950 757.950 241.050 760.050 ;
        RECT 230.400 748.050 231.600 757.950 ;
        RECT 236.400 756.900 237.600 757.950 ;
        RECT 235.950 754.800 238.050 756.900 ;
        RECT 245.400 748.050 246.600 761.100 ;
        RECT 260.400 760.050 261.600 761.100 ;
        RECT 266.400 760.050 267.600 761.100 ;
        RECT 247.950 757.950 250.050 760.050 ;
        RECT 256.950 757.950 259.050 760.050 ;
        RECT 259.950 757.950 262.050 760.050 ;
        RECT 262.950 757.950 265.050 760.050 ;
        RECT 265.950 757.950 268.050 760.050 ;
        RECT 223.950 745.950 226.050 748.050 ;
        RECT 229.950 745.950 232.050 748.050 ;
        RECT 244.950 745.950 247.050 748.050 ;
        RECT 220.950 736.950 223.050 739.050 ;
        RECT 214.950 728.100 217.050 730.200 ;
        RECT 215.400 727.050 216.600 728.100 ;
        RECT 208.950 724.950 211.050 727.050 ;
        RECT 211.950 724.950 214.050 727.050 ;
        RECT 214.950 724.950 217.050 727.050 ;
        RECT 217.950 724.950 220.050 727.050 ;
        RECT 212.400 718.050 213.600 724.950 ;
        RECT 218.400 723.600 219.600 724.950 ;
        RECT 224.400 723.600 225.600 745.950 ;
        RECT 235.950 736.950 238.050 739.050 ;
        RECT 236.400 727.050 237.600 736.950 ;
        RECT 241.950 728.100 244.050 730.200 ;
        RECT 242.400 727.050 243.600 728.100 ;
        RECT 232.950 724.950 235.050 727.050 ;
        RECT 235.950 724.950 238.050 727.050 ;
        RECT 238.950 724.950 241.050 727.050 ;
        RECT 241.950 724.950 244.050 727.050 ;
        RECT 218.400 722.400 225.600 723.600 ;
        RECT 190.950 715.950 193.050 718.050 ;
        RECT 196.950 715.950 199.050 718.050 ;
        RECT 211.950 715.950 214.050 718.050 ;
        RECT 187.950 712.500 190.050 714.600 ;
        RECT 212.400 693.600 213.600 715.950 ;
        RECT 233.400 714.600 234.600 724.950 ;
        RECT 239.400 723.900 240.600 724.950 ;
        RECT 238.950 721.800 241.050 723.900 ;
        RECT 248.400 718.050 249.600 757.950 ;
        RECT 257.400 756.900 258.600 757.950 ;
        RECT 256.950 754.800 259.050 756.900 ;
        RECT 263.400 751.050 264.600 757.950 ;
        RECT 268.950 754.950 271.050 757.050 ;
        RECT 262.950 748.950 265.050 751.050 ;
        RECT 269.400 748.050 270.600 754.950 ;
        RECT 259.950 745.950 262.050 748.050 ;
        RECT 268.950 745.950 271.050 748.050 ;
        RECT 253.950 728.100 256.050 730.200 ;
        RECT 254.400 727.050 255.600 728.100 ;
        RECT 260.400 727.050 261.600 745.950 ;
        RECT 268.950 733.950 271.050 736.050 ;
        RECT 253.950 724.950 256.050 727.050 ;
        RECT 256.950 724.950 259.050 727.050 ;
        RECT 259.950 724.950 262.050 727.050 ;
        RECT 262.950 724.950 265.050 727.050 ;
        RECT 257.400 723.900 258.600 724.950 ;
        RECT 263.400 723.900 264.600 724.950 ;
        RECT 256.950 721.800 259.050 723.900 ;
        RECT 262.950 721.800 265.050 723.900 ;
        RECT 257.400 720.600 258.600 721.800 ;
        RECT 257.400 719.400 261.600 720.600 ;
        RECT 235.950 714.600 238.050 718.050 ;
        RECT 247.950 715.950 250.050 718.050 ;
        RECT 233.400 714.000 238.050 714.600 ;
        RECT 233.400 713.400 237.600 714.000 ;
        RECT 209.400 692.400 213.600 693.600 ;
        RECT 202.950 688.950 205.050 691.050 ;
        RECT 157.950 682.950 160.050 685.050 ;
        RECT 166.950 683.100 169.050 685.200 ;
        RECT 175.950 683.100 178.050 685.200 ;
        RECT 154.950 679.950 157.050 682.050 ;
        RECT 160.950 679.950 163.050 682.050 ;
        RECT 148.950 676.950 151.050 679.050 ;
        RECT 161.400 664.050 162.600 679.950 ;
        RECT 167.400 679.050 168.600 683.100 ;
        RECT 176.400 682.050 177.600 683.100 ;
        RECT 187.950 682.950 190.050 685.050 ;
        RECT 196.950 684.000 199.050 688.050 ;
        RECT 175.950 679.950 178.050 682.050 ;
        RECT 178.950 679.950 181.050 682.050 ;
        RECT 166.950 676.950 169.050 679.050 ;
        RECT 179.400 670.050 180.600 679.950 ;
        RECT 188.400 676.050 189.600 682.950 ;
        RECT 197.400 682.050 198.600 684.000 ;
        RECT 203.400 682.050 204.600 688.950 ;
        RECT 193.950 679.950 196.050 682.050 ;
        RECT 196.950 679.950 199.050 682.050 ;
        RECT 199.950 679.950 202.050 682.050 ;
        RECT 202.950 679.950 205.050 682.050 ;
        RECT 187.950 673.950 190.050 676.050 ;
        RECT 178.950 667.950 181.050 670.050 ;
        RECT 160.950 661.950 163.050 664.050 ;
        RECT 190.950 661.950 193.050 664.050 ;
        RECT 145.950 655.950 148.050 658.050 ;
        RECT 157.950 656.400 160.050 658.500 ;
        RECT 146.400 646.050 147.600 655.950 ;
        RECT 151.950 646.950 154.050 649.050 ;
        RECT 145.950 643.950 148.050 646.050 ;
        RECT 152.400 645.600 153.600 646.950 ;
        RECT 151.950 643.500 154.050 645.600 ;
        RECT 158.100 636.600 159.300 656.400 ;
        RECT 181.950 655.950 184.050 658.050 ;
        RECT 166.950 650.100 169.050 652.200 ;
        RECT 175.950 650.100 178.050 652.200 ;
        RECT 160.950 646.950 163.050 649.050 ;
        RECT 161.400 645.600 162.600 646.950 ;
        RECT 167.400 645.600 168.600 650.100 ;
        RECT 176.400 649.050 177.600 650.100 ;
        RECT 182.400 649.050 183.600 655.950 ;
        RECT 175.950 646.950 178.050 649.050 ;
        RECT 178.950 646.950 181.050 649.050 ;
        RECT 181.950 646.950 184.050 649.050 ;
        RECT 184.950 646.950 187.050 649.050 ;
        RECT 160.950 643.500 163.050 645.600 ;
        RECT 164.400 644.400 168.600 645.600 ;
        RECT 161.400 640.050 162.600 643.500 ;
        RECT 160.950 637.950 163.050 640.050 ;
        RECT 157.950 634.500 160.050 636.600 ;
        RECT 136.950 628.950 139.050 631.050 ;
        RECT 142.950 628.950 145.050 631.050 ;
        RECT 115.950 619.950 118.050 622.050 ;
        RECT 124.950 619.950 127.050 622.050 ;
        RECT 118.950 605.100 121.050 607.200 ;
        RECT 119.400 604.050 120.600 605.100 ;
        RECT 125.400 604.050 126.600 619.950 ;
        RECT 118.950 601.950 121.050 604.050 ;
        RECT 121.950 601.950 124.050 604.050 ;
        RECT 124.950 601.950 127.050 604.050 ;
        RECT 122.400 600.900 123.600 601.950 ;
        RECT 121.950 598.800 124.050 600.900 ;
        RECT 133.950 598.950 136.050 601.050 ;
        RECT 137.400 600.600 138.600 628.950 ;
        RECT 164.400 622.050 165.600 644.400 ;
        RECT 179.400 642.600 180.600 646.950 ;
        RECT 185.400 642.600 186.600 646.950 ;
        RECT 176.400 641.400 180.600 642.600 ;
        RECT 182.400 641.400 186.600 642.600 ;
        RECT 176.400 637.050 177.600 641.400 ;
        RECT 182.400 639.600 183.600 641.400 ;
        RECT 179.400 638.400 183.600 639.600 ;
        RECT 175.950 634.950 178.050 637.050 ;
        RECT 175.950 628.950 178.050 631.050 ;
        RECT 163.950 619.950 166.050 622.050 ;
        RECT 145.950 616.950 148.050 619.050 ;
        RECT 157.950 616.950 160.050 619.050 ;
        RECT 146.400 604.050 147.600 616.950 ;
        RECT 154.950 610.950 157.050 613.050 ;
        RECT 142.950 601.950 145.050 604.050 ;
        RECT 145.950 601.950 148.050 604.050 ;
        RECT 148.950 601.950 151.050 604.050 ;
        RECT 137.400 599.400 141.600 600.600 ;
        RECT 127.950 577.950 130.050 580.050 ;
        RECT 113.400 572.400 117.600 573.600 ;
        RECT 106.950 568.950 109.050 571.050 ;
        RECT 109.950 568.950 112.050 571.050 ;
        RECT 110.400 567.900 111.600 568.950 ;
        RECT 109.950 565.800 112.050 567.900 ;
        RECT 100.950 562.950 103.050 565.050 ;
        RECT 97.950 541.950 100.050 544.050 ;
        RECT 103.950 536.400 106.050 538.500 ;
        RECT 110.400 538.050 111.600 565.800 ;
        RECT 116.400 550.050 117.600 572.400 ;
        RECT 128.400 571.050 129.600 577.950 ;
        RECT 134.400 573.600 135.600 598.950 ;
        RECT 134.400 572.400 138.600 573.600 ;
        RECT 124.950 568.950 127.050 571.050 ;
        RECT 127.950 568.950 130.050 571.050 ;
        RECT 130.950 568.950 133.050 571.050 ;
        RECT 125.400 567.000 126.600 568.950 ;
        RECT 131.400 567.900 132.600 568.950 ;
        RECT 124.950 562.950 127.050 567.000 ;
        RECT 130.950 565.800 133.050 567.900 ;
        RECT 115.950 547.950 118.050 550.050 ;
        RECT 112.950 541.950 115.050 544.050 ;
        RECT 88.950 528.600 93.000 529.050 ;
        RECT 88.950 526.950 93.600 528.600 ;
        RECT 94.950 526.950 97.050 529.050 ;
        RECT 99.000 528.600 103.050 529.050 ;
        RECT 98.400 526.950 103.050 528.600 ;
        RECT 82.950 514.500 85.050 516.600 ;
        RECT 73.950 511.950 76.050 514.050 ;
        RECT 71.400 509.400 75.600 510.600 ;
        RECT 74.400 493.050 75.600 509.400 ;
        RECT 85.950 500.400 88.050 502.500 ;
        RECT 82.950 494.400 85.050 496.500 ;
        RECT 83.400 493.050 84.600 494.400 ;
        RECT 70.950 490.950 73.050 493.050 ;
        RECT 73.950 490.950 76.050 493.050 ;
        RECT 76.950 490.950 79.050 493.050 ;
        RECT 82.950 490.950 85.050 493.050 ;
        RECT 71.400 489.900 72.600 490.950 ;
        RECT 77.400 489.900 78.600 490.950 ;
        RECT 70.950 487.800 73.050 489.900 ;
        RECT 76.950 487.800 79.050 489.900 ;
        RECT 71.400 486.600 72.600 487.800 ;
        RECT 71.400 485.400 75.600 486.600 ;
        RECT 64.950 451.950 67.050 454.050 ;
        RECT 74.400 451.200 75.600 485.400 ;
        RECT 77.400 454.050 78.600 487.800 ;
        RECT 86.850 485.400 88.050 500.400 ;
        RECT 92.400 493.050 93.600 526.950 ;
        RECT 98.400 526.050 99.600 526.950 ;
        RECT 97.950 523.950 100.050 526.050 ;
        RECT 104.100 516.600 105.300 536.400 ;
        RECT 109.950 535.950 112.050 538.050 ;
        RECT 109.950 532.800 112.050 534.900 ;
        RECT 110.400 528.600 111.600 532.800 ;
        RECT 107.400 527.400 111.600 528.600 ;
        RECT 107.400 526.050 108.600 527.400 ;
        RECT 106.950 523.950 109.050 526.050 ;
        RECT 103.950 514.500 106.050 516.600 ;
        RECT 106.950 500.400 109.050 502.500 ;
        RECT 94.950 493.950 97.050 496.050 ;
        RECT 91.950 490.950 94.050 493.050 ;
        RECT 95.400 489.600 96.600 493.950 ;
        RECT 100.950 490.950 103.050 493.050 ;
        RECT 101.400 489.600 102.600 490.950 ;
        RECT 94.950 487.500 97.050 489.600 ;
        RECT 100.950 487.500 103.050 489.600 ;
        RECT 85.950 483.300 88.050 485.400 ;
        RECT 86.850 479.700 88.050 483.300 ;
        RECT 107.100 480.600 108.300 500.400 ;
        RECT 113.400 496.050 114.600 541.950 ;
        RECT 137.400 538.050 138.600 572.400 ;
        RECT 124.950 535.950 127.050 538.050 ;
        RECT 136.950 535.950 139.050 538.050 ;
        RECT 115.950 526.950 118.050 529.050 ;
        RECT 116.400 517.050 117.600 526.950 ;
        RECT 125.400 526.050 126.600 535.950 ;
        RECT 130.950 528.000 133.050 532.050 ;
        RECT 136.950 529.950 139.050 532.050 ;
        RECT 131.400 526.050 132.600 528.000 ;
        RECT 121.950 523.950 124.050 526.050 ;
        RECT 124.950 523.950 127.050 526.050 ;
        RECT 127.950 523.950 130.050 526.050 ;
        RECT 130.950 523.950 133.050 526.050 ;
        RECT 122.400 522.900 123.600 523.950 ;
        RECT 121.950 520.800 124.050 522.900 ;
        RECT 128.400 517.050 129.600 523.950 ;
        RECT 137.400 523.050 138.600 529.950 ;
        RECT 136.950 520.950 139.050 523.050 ;
        RECT 140.400 517.050 141.600 599.400 ;
        RECT 143.400 574.050 144.600 601.950 ;
        RECT 149.400 600.900 150.600 601.950 ;
        RECT 155.400 600.900 156.600 610.950 ;
        RECT 148.950 598.800 151.050 600.900 ;
        RECT 154.950 598.800 157.050 600.900 ;
        RECT 151.950 589.950 154.050 592.050 ;
        RECT 145.950 577.950 148.050 580.050 ;
        RECT 142.950 571.950 145.050 574.050 ;
        RECT 146.400 571.050 147.600 577.950 ;
        RECT 152.400 571.050 153.600 589.950 ;
        RECT 158.400 574.050 159.600 616.950 ;
        RECT 164.400 610.050 165.600 619.950 ;
        RECT 163.950 607.950 166.050 610.050 ;
        RECT 164.400 604.050 165.600 607.950 ;
        RECT 163.950 601.950 166.050 604.050 ;
        RECT 169.950 601.950 172.050 604.050 ;
        RECT 160.950 598.950 163.050 601.050 ;
        RECT 170.400 600.900 171.600 601.950 ;
        RECT 176.400 601.050 177.600 628.950 ;
        RECT 157.950 571.950 160.050 574.050 ;
        RECT 145.950 568.950 148.050 571.050 ;
        RECT 148.950 568.950 151.050 571.050 ;
        RECT 151.950 568.950 154.050 571.050 ;
        RECT 154.950 568.950 157.050 571.050 ;
        RECT 149.400 567.000 150.600 568.950 ;
        RECT 155.400 567.000 156.600 568.950 ;
        RECT 148.950 562.950 151.050 567.000 ;
        RECT 154.950 562.950 157.050 567.000 ;
        RECT 161.400 565.050 162.600 598.950 ;
        RECT 169.950 598.800 172.050 600.900 ;
        RECT 175.950 598.950 178.050 601.050 ;
        RECT 166.950 574.950 169.050 577.050 ;
        RECT 163.950 571.950 166.050 574.050 ;
        RECT 160.950 562.950 163.050 565.050 ;
        RECT 164.400 550.050 165.600 571.950 ;
        RECT 167.400 565.050 168.600 574.950 ;
        RECT 175.950 573.000 178.050 577.050 ;
        RECT 179.400 574.050 180.600 638.400 ;
        RECT 184.950 637.950 187.050 640.050 ;
        RECT 185.400 619.050 186.600 637.950 ;
        RECT 191.400 631.050 192.600 661.950 ;
        RECT 194.400 640.050 195.600 679.950 ;
        RECT 200.400 678.000 201.600 679.950 ;
        RECT 199.950 673.950 202.050 678.000 ;
        RECT 205.950 676.950 208.050 679.050 ;
        RECT 206.400 664.050 207.600 676.950 ;
        RECT 205.950 661.950 208.050 664.050 ;
        RECT 205.950 651.000 208.050 655.050 ;
        RECT 209.400 652.050 210.600 692.400 ;
        RECT 232.950 691.950 235.050 694.050 ;
        RECT 229.950 688.950 232.050 691.050 ;
        RECT 214.950 683.100 217.050 685.200 ;
        RECT 220.950 683.100 223.050 685.200 ;
        RECT 215.400 682.050 216.600 683.100 ;
        RECT 221.400 682.050 222.600 683.100 ;
        RECT 214.950 679.950 217.050 682.050 ;
        RECT 217.950 679.950 220.050 682.050 ;
        RECT 220.950 679.950 223.050 682.050 ;
        RECT 223.950 679.950 226.050 682.050 ;
        RECT 211.950 676.950 214.050 679.050 ;
        RECT 206.400 649.050 207.600 651.000 ;
        RECT 208.950 649.950 211.050 652.050 ;
        RECT 202.950 646.950 205.050 649.050 ;
        RECT 205.950 646.950 208.050 649.050 ;
        RECT 203.400 645.900 204.600 646.950 ;
        RECT 202.950 643.800 205.050 645.900 ;
        RECT 193.950 637.950 196.050 640.050 ;
        RECT 190.950 628.950 193.050 631.050 ;
        RECT 184.950 616.950 187.050 619.050 ;
        RECT 185.400 610.050 186.600 616.950 ;
        RECT 199.950 614.400 202.050 616.500 ;
        RECT 187.950 610.950 190.050 613.050 ;
        RECT 184.950 607.950 187.050 610.050 ;
        RECT 188.400 604.050 189.600 610.950 ;
        RECT 196.950 606.000 199.050 610.050 ;
        RECT 197.400 604.050 198.600 606.000 ;
        RECT 184.950 601.950 187.050 604.050 ;
        RECT 187.950 601.950 190.050 604.050 ;
        RECT 190.950 601.950 193.050 604.050 ;
        RECT 196.950 601.950 199.050 604.050 ;
        RECT 181.950 580.950 184.050 583.050 ;
        RECT 176.400 571.050 177.600 573.000 ;
        RECT 178.950 571.950 181.050 574.050 ;
        RECT 172.950 568.950 175.050 571.050 ;
        RECT 175.950 568.950 178.050 571.050 ;
        RECT 173.400 567.900 174.600 568.950 ;
        RECT 172.950 565.800 175.050 567.900 ;
        RECT 182.400 565.050 183.600 580.950 ;
        RECT 185.400 574.050 186.600 601.950 ;
        RECT 191.400 583.050 192.600 601.950 ;
        RECT 200.700 594.600 201.900 614.400 ;
        RECT 205.950 605.400 208.050 607.500 ;
        RECT 206.400 604.050 207.600 605.400 ;
        RECT 205.950 601.950 208.050 604.050 ;
        RECT 208.950 598.800 211.050 600.900 ;
        RECT 209.400 594.600 210.600 598.800 ;
        RECT 212.400 598.050 213.600 676.950 ;
        RECT 218.400 667.050 219.600 679.950 ;
        RECT 224.400 678.900 225.600 679.950 ;
        RECT 223.950 676.800 226.050 678.900 ;
        RECT 220.950 673.950 223.050 676.050 ;
        RECT 217.950 664.950 220.050 667.050 ;
        RECT 214.950 658.950 217.050 661.050 ;
        RECT 215.400 655.050 216.600 658.950 ;
        RECT 221.400 658.050 222.600 673.950 ;
        RECT 230.400 667.050 231.600 688.950 ;
        RECT 229.950 664.950 232.050 667.050 ;
        RECT 220.950 655.950 223.050 658.050 ;
        RECT 214.950 652.950 217.050 655.050 ;
        RECT 214.950 649.800 217.050 651.900 ;
        RECT 223.950 650.100 226.050 652.200 ;
        RECT 229.950 650.100 232.050 652.200 ;
        RECT 233.400 651.600 234.600 691.950 ;
        RECT 236.400 679.050 237.600 713.400 ;
        RECT 247.950 694.950 250.050 697.050 ;
        RECT 241.950 683.100 244.050 685.200 ;
        RECT 242.400 682.050 243.600 683.100 ;
        RECT 248.400 682.050 249.600 694.950 ;
        RECT 256.950 683.100 259.050 685.200 ;
        RECT 241.950 679.950 244.050 682.050 ;
        RECT 244.950 679.950 247.050 682.050 ;
        RECT 247.950 679.950 250.050 682.050 ;
        RECT 250.950 679.950 253.050 682.050 ;
        RECT 235.950 676.950 238.050 679.050 ;
        RECT 245.400 678.900 246.600 679.950 ;
        RECT 244.950 676.800 247.050 678.900 ;
        RECT 251.400 670.050 252.600 679.950 ;
        RECT 250.950 667.950 253.050 670.050 ;
        RECT 257.400 667.050 258.600 683.100 ;
        RECT 260.400 676.050 261.600 719.400 ;
        RECT 263.400 685.050 264.600 721.800 ;
        RECT 262.950 682.950 265.050 685.050 ;
        RECT 269.400 682.050 270.600 733.950 ;
        RECT 272.400 724.050 273.600 761.100 ;
        RECT 275.400 757.050 276.600 787.950 ;
        RECT 308.400 775.050 309.600 796.950 ;
        RECT 332.400 796.050 333.600 802.950 ;
        RECT 313.950 793.950 316.050 796.050 ;
        RECT 331.950 793.950 334.050 796.050 ;
        RECT 307.950 772.950 310.050 775.050 ;
        RECT 283.950 761.100 286.050 766.050 ;
        RECT 295.950 762.600 298.050 763.200 ;
        RECT 290.400 761.400 298.050 762.600 ;
        RECT 301.950 762.000 304.050 766.050 ;
        RECT 284.400 760.050 285.600 761.100 ;
        RECT 290.400 760.050 291.600 761.400 ;
        RECT 295.950 761.100 298.050 761.400 ;
        RECT 280.950 757.950 283.050 760.050 ;
        RECT 283.950 757.950 286.050 760.050 ;
        RECT 286.950 757.950 289.050 760.050 ;
        RECT 289.950 757.950 292.050 760.050 ;
        RECT 274.950 754.950 277.050 757.050 ;
        RECT 281.400 756.900 282.600 757.950 ;
        RECT 287.400 756.900 288.600 757.950 ;
        RECT 280.950 754.800 283.050 756.900 ;
        RECT 286.950 754.800 289.050 756.900 ;
        RECT 287.400 748.050 288.600 754.800 ;
        RECT 296.400 751.050 297.600 761.100 ;
        RECT 302.400 760.050 303.600 762.000 ;
        RECT 307.950 761.100 310.050 763.200 ;
        RECT 314.400 763.050 315.600 793.950 ;
        RECT 325.950 784.950 328.050 787.050 ;
        RECT 316.950 772.950 319.050 775.050 ;
        RECT 308.400 760.050 309.600 761.100 ;
        RECT 313.950 760.950 316.050 763.050 ;
        RECT 301.950 757.950 304.050 760.050 ;
        RECT 304.950 757.950 307.050 760.050 ;
        RECT 307.950 757.950 310.050 760.050 ;
        RECT 310.950 757.950 313.050 760.050 ;
        RECT 305.400 756.900 306.600 757.950 ;
        RECT 311.400 756.900 312.600 757.950 ;
        RECT 304.950 754.800 307.050 756.900 ;
        RECT 310.950 754.800 313.050 756.900 ;
        RECT 295.950 748.950 298.050 751.050 ;
        RECT 286.950 745.950 289.050 748.050 ;
        RECT 274.950 739.950 277.050 742.050 ;
        RECT 271.950 721.950 274.050 724.050 ;
        RECT 275.400 694.050 276.600 739.950 ;
        RECT 280.950 728.100 283.050 730.200 ;
        RECT 286.950 728.100 289.050 730.200 ;
        RECT 281.400 727.050 282.600 728.100 ;
        RECT 287.400 727.050 288.600 728.100 ;
        RECT 305.400 727.050 306.600 754.800 ;
        RECT 317.400 748.050 318.600 772.950 ;
        RECT 319.950 763.950 322.050 766.050 ;
        RECT 316.950 745.950 319.050 748.050 ;
        RECT 310.950 728.100 313.050 730.200 ;
        RECT 311.400 727.050 312.600 728.100 ;
        RECT 280.950 724.950 283.050 727.050 ;
        RECT 283.950 724.950 286.050 727.050 ;
        RECT 286.950 724.950 289.050 727.050 ;
        RECT 289.950 724.950 292.050 727.050 ;
        RECT 304.950 724.950 307.050 727.050 ;
        RECT 307.950 724.950 310.050 727.050 ;
        RECT 310.950 724.950 313.050 727.050 ;
        RECT 313.950 724.950 316.050 727.050 ;
        RECT 284.400 723.000 285.600 724.950 ;
        RECT 290.400 723.900 291.600 724.950 ;
        RECT 308.400 723.900 309.600 724.950 ;
        RECT 314.400 723.900 315.600 724.950 ;
        RECT 283.950 718.950 286.050 723.000 ;
        RECT 289.950 721.800 292.050 723.900 ;
        RECT 307.950 718.950 310.050 723.900 ;
        RECT 313.950 718.950 316.050 723.900 ;
        RECT 320.400 721.050 321.600 763.950 ;
        RECT 326.400 760.050 327.600 784.950 ;
        RECT 338.400 781.050 339.600 802.950 ;
        RECT 344.400 802.050 345.600 806.100 ;
        RECT 343.950 799.950 346.050 802.050 ;
        RECT 347.400 793.050 348.600 830.400 ;
        RECT 364.950 829.950 367.050 834.000 ;
        RECT 370.950 829.950 373.050 834.900 ;
        RECT 364.950 817.950 367.050 820.050 ;
        RECT 355.950 806.100 358.050 808.200 ;
        RECT 356.400 805.050 357.600 806.100 ;
        RECT 352.950 802.950 355.050 805.050 ;
        RECT 355.950 802.950 358.050 805.050 ;
        RECT 353.400 801.900 354.600 802.950 ;
        RECT 352.950 799.800 355.050 801.900 ;
        RECT 346.950 790.950 349.050 793.050 ;
        RECT 361.950 784.950 364.050 787.050 ;
        RECT 337.950 778.950 340.050 781.050 ;
        RECT 358.950 769.950 361.050 772.050 ;
        RECT 343.950 760.950 346.050 763.050 ;
        RECT 349.950 761.100 352.050 763.200 ;
        RECT 325.950 757.950 328.050 760.050 ;
        RECT 328.950 757.950 331.050 760.050 ;
        RECT 329.400 736.050 330.600 757.950 ;
        RECT 328.950 733.950 331.050 736.050 ;
        RECT 334.950 733.950 337.050 736.050 ;
        RECT 329.400 732.600 330.600 733.950 ;
        RECT 326.400 731.400 330.600 732.600 ;
        RECT 326.400 727.050 327.600 731.400 ;
        RECT 325.950 724.950 328.050 727.050 ;
        RECT 328.950 724.950 331.050 727.050 ;
        RECT 329.400 723.900 330.600 724.950 ;
        RECT 328.950 721.800 331.050 723.900 ;
        RECT 319.950 718.950 322.050 721.050 ;
        RECT 274.950 691.950 277.050 694.050 ;
        RECT 308.400 690.600 309.600 718.950 ;
        RECT 335.400 718.050 336.600 733.950 ;
        RECT 344.400 732.600 345.600 760.950 ;
        RECT 350.400 760.050 351.600 761.100 ;
        RECT 349.950 757.950 352.050 760.050 ;
        RECT 352.950 757.950 355.050 760.050 ;
        RECT 353.400 756.900 354.600 757.950 ;
        RECT 359.400 756.900 360.600 769.950 ;
        RECT 352.950 754.800 355.050 756.900 ;
        RECT 358.950 754.800 361.050 756.900 ;
        RECT 352.950 745.950 355.050 748.050 ;
        RECT 344.400 731.400 348.600 732.600 ;
        RECT 347.400 730.200 348.600 731.400 ;
        RECT 346.950 728.100 349.050 730.200 ;
        RECT 347.400 727.050 348.600 728.100 ;
        RECT 353.400 727.050 354.600 745.950 ;
        RECT 359.400 730.200 360.600 754.800 ;
        RECT 358.950 728.100 361.050 730.200 ;
        RECT 343.950 724.950 346.050 727.050 ;
        RECT 346.950 724.950 349.050 727.050 ;
        RECT 349.950 724.950 352.050 727.050 ;
        RECT 352.950 724.950 355.050 727.050 ;
        RECT 344.400 723.900 345.600 724.950 ;
        RECT 350.400 723.900 351.600 724.950 ;
        RECT 343.950 721.800 346.050 723.900 ;
        RECT 349.950 721.800 352.050 723.900 ;
        RECT 334.950 715.950 337.050 718.050 ;
        RECT 355.950 700.950 358.050 703.050 ;
        RECT 328.950 697.950 331.050 700.050 ;
        RECT 322.950 694.950 325.050 697.050 ;
        RECT 310.950 691.950 313.050 694.050 ;
        RECT 305.400 689.400 309.600 690.600 ;
        RECT 274.950 683.100 277.050 685.200 ;
        RECT 283.950 683.100 286.050 685.200 ;
        RECT 295.950 683.100 298.050 685.200 ;
        RECT 301.950 683.100 304.050 685.200 ;
        RECT 275.400 682.050 276.600 683.100 ;
        RECT 265.950 679.950 268.050 682.050 ;
        RECT 268.950 679.950 271.050 682.050 ;
        RECT 271.950 679.950 274.050 682.050 ;
        RECT 274.950 679.950 277.050 682.050 ;
        RECT 266.400 678.000 267.600 679.950 ;
        RECT 272.400 678.900 273.600 679.950 ;
        RECT 259.950 673.950 262.050 676.050 ;
        RECT 265.950 673.950 268.050 678.000 ;
        RECT 271.950 676.800 274.050 678.900 ;
        RECT 280.950 676.800 283.050 678.900 ;
        RECT 256.950 664.950 259.050 667.050 ;
        RECT 281.400 661.050 282.600 676.800 ;
        RECT 274.950 658.950 277.050 661.050 ;
        RECT 280.950 658.950 283.050 661.050 ;
        RECT 238.950 652.950 241.050 655.050 ;
        RECT 233.400 650.400 237.600 651.600 ;
        RECT 215.400 613.050 216.600 649.800 ;
        RECT 224.400 649.050 225.600 650.100 ;
        RECT 230.400 649.050 231.600 650.100 ;
        RECT 220.950 646.950 223.050 649.050 ;
        RECT 223.950 646.950 226.050 649.050 ;
        RECT 226.950 646.950 229.050 649.050 ;
        RECT 229.950 646.950 232.050 649.050 ;
        RECT 221.400 622.050 222.600 646.950 ;
        RECT 227.400 645.900 228.600 646.950 ;
        RECT 226.950 643.800 229.050 645.900 ;
        RECT 220.950 619.950 223.050 622.050 ;
        RECT 232.950 619.950 235.050 622.050 ;
        RECT 220.950 615.300 223.050 617.400 ;
        RECT 214.950 610.950 217.050 613.050 ;
        RECT 220.950 611.700 222.150 615.300 ;
        RECT 220.950 609.600 223.050 611.700 ;
        RECT 229.950 610.950 232.050 613.050 ;
        RECT 214.950 605.400 217.050 607.500 ;
        RECT 215.400 601.050 216.600 605.400 ;
        RECT 214.950 598.950 217.050 601.050 ;
        RECT 211.950 595.950 214.050 598.050 ;
        RECT 220.950 594.600 222.150 609.600 ;
        RECT 223.950 601.950 226.050 604.050 ;
        RECT 224.400 600.600 225.600 601.950 ;
        RECT 224.400 599.400 228.600 600.600 ;
        RECT 227.400 595.050 228.600 599.400 ;
        RECT 199.950 592.500 202.050 594.600 ;
        RECT 209.400 593.400 213.600 594.600 ;
        RECT 190.950 580.950 193.050 583.050 ;
        RECT 199.950 580.950 202.050 583.050 ;
        RECT 184.950 571.950 187.050 574.050 ;
        RECT 190.950 573.000 193.050 577.050 ;
        RECT 200.400 573.600 201.600 580.950 ;
        RECT 205.950 578.400 208.050 580.500 ;
        RECT 191.400 571.050 192.600 573.000 ;
        RECT 200.400 572.400 204.600 573.600 ;
        RECT 203.400 571.050 204.600 572.400 ;
        RECT 187.950 568.950 190.050 571.050 ;
        RECT 190.950 568.950 193.050 571.050 ;
        RECT 193.950 568.950 196.050 571.050 ;
        RECT 202.950 568.950 205.050 571.050 ;
        RECT 188.400 567.000 189.600 568.950 ;
        RECT 194.400 567.900 195.600 568.950 ;
        RECT 166.950 562.950 169.050 565.050 ;
        RECT 175.950 562.950 178.050 565.050 ;
        RECT 181.950 562.950 184.050 565.050 ;
        RECT 187.950 562.950 190.050 567.000 ;
        RECT 193.950 565.800 196.050 567.900 ;
        RECT 206.850 563.400 208.050 578.400 ;
        RECT 163.950 547.950 166.050 550.050 ;
        RECT 176.400 544.050 177.600 562.950 ;
        RECT 188.400 550.050 189.600 562.950 ;
        RECT 205.950 561.300 208.050 563.400 ;
        RECT 206.850 557.700 208.050 561.300 ;
        RECT 205.950 555.600 208.050 557.700 ;
        RECT 212.400 556.050 213.600 593.400 ;
        RECT 220.950 592.500 223.050 594.600 ;
        RECT 226.950 592.950 229.050 595.050 ;
        RECT 230.400 589.050 231.600 610.950 ;
        RECT 214.950 586.950 217.050 589.050 ;
        RECT 229.950 586.950 232.050 589.050 ;
        RECT 211.950 553.950 214.050 556.050 ;
        RECT 178.950 547.950 181.050 550.050 ;
        RECT 187.950 547.950 190.050 550.050 ;
        RECT 196.950 547.950 199.050 550.050 ;
        RECT 175.950 541.950 178.050 544.050 ;
        RECT 145.950 538.950 148.050 541.050 ;
        RECT 146.400 529.200 147.600 538.950 ;
        RECT 163.950 537.300 166.050 539.400 ;
        RECT 164.850 533.700 166.050 537.300 ;
        RECT 179.400 535.050 180.600 547.950 ;
        RECT 184.950 536.400 187.050 538.500 ;
        RECT 163.950 531.600 166.050 533.700 ;
        RECT 178.950 532.950 181.050 535.050 ;
        RECT 145.950 527.100 148.050 529.200 ;
        RECT 151.950 527.100 154.050 529.200 ;
        RECT 146.400 526.050 147.600 527.100 ;
        RECT 152.400 526.050 153.600 527.100 ;
        RECT 145.950 523.950 148.050 526.050 ;
        RECT 148.950 523.950 151.050 526.050 ;
        RECT 151.950 523.950 154.050 526.050 ;
        RECT 160.950 523.950 163.050 526.050 ;
        RECT 149.400 522.900 150.600 523.950 ;
        RECT 148.950 520.800 151.050 522.900 ;
        RECT 161.400 522.600 162.600 523.950 ;
        RECT 158.400 521.400 162.600 522.600 ;
        RECT 115.950 514.950 118.050 517.050 ;
        RECT 127.950 514.950 130.050 517.050 ;
        RECT 139.950 514.950 142.050 517.050 ;
        RECT 158.400 502.050 159.600 521.400 ;
        RECT 164.850 516.600 166.050 531.600 ;
        RECT 169.800 527.100 171.900 529.200 ;
        RECT 163.950 514.500 166.050 516.600 ;
        RECT 170.400 508.050 171.600 527.100 ;
        RECT 172.950 526.950 175.050 529.050 ;
        RECT 178.950 527.400 181.050 529.500 ;
        RECT 169.950 505.950 172.050 508.050 ;
        RECT 173.400 505.050 174.600 526.950 ;
        RECT 179.400 526.050 180.600 527.400 ;
        RECT 178.950 523.950 181.050 526.050 ;
        RECT 178.950 514.950 181.050 517.050 ;
        RECT 185.100 516.600 186.300 536.400 ;
        RECT 193.950 535.950 196.050 538.050 ;
        RECT 187.950 532.950 190.050 535.050 ;
        RECT 188.400 526.050 189.600 532.950 ;
        RECT 187.950 523.950 190.050 526.050 ;
        RECT 172.950 502.950 175.050 505.050 ;
        RECT 118.950 499.950 121.050 502.050 ;
        RECT 157.950 499.950 160.050 502.050 ;
        RECT 169.950 499.950 172.050 502.050 ;
        RECT 115.950 496.950 118.050 499.050 ;
        RECT 112.950 493.950 115.050 496.050 ;
        RECT 109.950 490.950 112.050 493.050 ;
        RECT 110.400 489.000 111.600 490.950 ;
        RECT 109.950 484.950 112.050 489.000 ;
        RECT 85.950 477.600 88.050 479.700 ;
        RECT 106.950 478.500 109.050 480.600 ;
        RECT 95.100 454.200 97.200 456.300 ;
        RECT 104.100 454.500 106.200 456.600 ;
        RECT 76.950 451.950 79.050 454.050 ;
        RECT 85.950 451.950 88.050 454.050 ;
        RECT 50.400 448.050 51.600 449.100 ;
        RECT 56.400 448.050 57.600 450.000 ;
        RECT 62.400 449.400 66.600 450.600 ;
        RECT 49.950 445.950 52.050 448.050 ;
        RECT 52.950 445.950 55.050 448.050 ;
        RECT 55.950 445.950 58.050 448.050 ;
        RECT 58.950 445.950 61.050 448.050 ;
        RECT 49.950 439.950 52.050 442.050 ;
        RECT 43.950 415.950 46.050 418.050 ;
        RECT 50.400 415.050 51.600 439.950 ;
        RECT 53.400 436.050 54.600 445.950 ;
        RECT 59.400 444.900 60.600 445.950 ;
        RECT 58.950 442.800 61.050 444.900 ;
        RECT 52.950 433.950 55.050 436.050 ;
        RECT 46.950 412.950 49.050 415.050 ;
        RECT 49.950 412.950 52.050 415.050 ;
        RECT 52.950 412.950 55.050 415.050 ;
        RECT 40.950 409.950 43.050 412.050 ;
        RECT 47.400 411.900 48.600 412.950 ;
        RECT 53.400 411.900 54.600 412.950 ;
        RECT 59.400 411.900 60.600 442.800 ;
        RECT 65.400 417.600 66.600 449.400 ;
        RECT 67.950 448.950 70.050 451.050 ;
        RECT 73.950 449.100 76.050 451.200 ;
        RECT 68.400 444.900 69.600 448.950 ;
        RECT 74.400 448.050 75.600 449.100 ;
        RECT 73.950 445.950 76.050 448.050 ;
        RECT 79.950 445.950 82.050 448.050 ;
        RECT 67.950 442.800 70.050 444.900 ;
        RECT 80.400 444.000 81.600 445.950 ;
        RECT 62.400 416.400 66.600 417.600 ;
        RECT 62.400 411.900 63.600 416.400 ;
        RECT 68.400 415.050 69.600 442.800 ;
        RECT 79.950 439.950 82.050 444.000 ;
        RECT 73.950 421.950 76.050 424.050 ;
        RECT 82.950 421.950 85.050 424.050 ;
        RECT 74.400 415.050 75.600 421.950 ;
        RECT 67.950 412.950 70.050 415.050 ;
        RECT 70.950 412.950 73.050 415.050 ;
        RECT 73.950 412.950 76.050 415.050 ;
        RECT 76.950 412.950 79.050 415.050 ;
        RECT 71.400 411.900 72.600 412.950 ;
        RECT 77.400 411.900 78.600 412.950 ;
        RECT 83.400 411.900 84.600 421.950 ;
        RECT 46.950 411.600 49.050 411.900 ;
        RECT 44.400 410.400 49.050 411.600 ;
        RECT 40.950 406.800 43.050 408.900 ;
        RECT 7.950 400.500 10.050 402.600 ;
        RECT 7.950 380.400 10.050 382.500 ;
        RECT 4.950 372.000 7.050 376.050 ;
        RECT 5.400 370.050 6.600 372.000 ;
        RECT 4.950 367.950 7.050 370.050 ;
        RECT 8.700 360.600 9.900 380.400 ;
        RECT 23.400 376.050 24.600 403.950 ;
        RECT 28.950 401.700 30.150 405.300 ;
        RECT 37.950 403.950 40.050 406.050 ;
        RECT 28.950 399.600 31.050 401.700 ;
        RECT 37.950 394.950 40.050 397.050 ;
        RECT 28.950 381.300 31.050 383.400 ;
        RECT 28.950 377.700 30.150 381.300 ;
        RECT 22.950 373.950 25.050 376.050 ;
        RECT 28.950 375.600 31.050 377.700 ;
        RECT 13.950 371.400 16.050 373.500 ;
        RECT 19.950 371.400 22.050 373.500 ;
        RECT 14.400 370.050 15.600 371.400 ;
        RECT 13.950 367.950 16.050 370.050 ;
        RECT 7.950 358.500 10.050 360.600 ;
        RECT 20.400 358.050 21.600 371.400 ;
        RECT 19.950 355.950 22.050 358.050 ;
        RECT 7.950 344.400 10.050 346.500 ;
        RECT 4.950 334.950 7.050 337.050 ;
        RECT 5.400 333.600 6.600 334.950 ;
        RECT 4.950 331.500 7.050 333.600 ;
        RECT 5.400 330.600 6.600 331.500 ;
        RECT 2.400 329.400 6.600 330.600 ;
        RECT 2.400 307.050 3.600 329.400 ;
        RECT 8.700 324.600 9.900 344.400 ;
        RECT 23.400 334.050 24.600 373.950 ;
        RECT 28.950 360.600 30.150 375.600 ;
        RECT 31.950 367.950 34.050 370.050 ;
        RECT 32.400 366.000 33.600 367.950 ;
        RECT 31.950 361.950 34.050 366.000 ;
        RECT 38.400 363.600 39.600 394.950 ;
        RECT 35.400 362.400 39.600 363.600 ;
        RECT 28.950 358.500 31.050 360.600 ;
        RECT 28.950 344.400 31.050 346.500 ;
        RECT 22.950 331.950 25.050 334.050 ;
        RECT 28.950 329.400 30.150 344.400 ;
        RECT 35.400 339.600 36.600 362.400 ;
        RECT 37.950 358.950 40.050 361.050 ;
        RECT 32.400 338.400 36.600 339.600 ;
        RECT 32.400 337.050 33.600 338.400 ;
        RECT 31.950 334.950 34.050 337.050 ;
        RECT 38.400 331.050 39.600 358.950 ;
        RECT 41.400 343.050 42.600 406.800 ;
        RECT 40.950 340.950 43.050 343.050 ;
        RECT 44.400 339.600 45.600 410.400 ;
        RECT 46.950 409.800 49.050 410.400 ;
        RECT 52.950 409.800 55.050 411.900 ;
        RECT 58.800 409.800 60.900 411.900 ;
        RECT 61.950 409.800 64.050 411.900 ;
        RECT 70.950 409.800 73.050 411.900 ;
        RECT 76.950 409.800 79.050 411.900 ;
        RECT 82.950 409.800 85.050 411.900 ;
        RECT 55.950 403.950 58.050 406.050 ;
        RECT 49.950 371.100 52.050 373.200 ;
        RECT 50.400 370.050 51.600 371.100 ;
        RECT 56.400 370.050 57.600 403.950 ;
        RECT 59.400 403.050 60.600 409.800 ;
        RECT 64.950 403.950 67.050 406.050 ;
        RECT 58.950 400.950 61.050 403.050 ;
        RECT 49.950 367.950 52.050 370.050 ;
        RECT 52.950 367.950 55.050 370.050 ;
        RECT 55.950 367.950 58.050 370.050 ;
        RECT 58.950 367.950 61.050 370.050 ;
        RECT 49.950 361.950 52.050 364.050 ;
        RECT 41.400 338.400 45.600 339.600 ;
        RECT 28.950 327.300 31.050 329.400 ;
        RECT 37.950 328.950 40.050 331.050 ;
        RECT 7.950 322.500 10.050 324.600 ;
        RECT 28.950 323.700 30.150 327.300 ;
        RECT 28.950 321.600 31.050 323.700 ;
        RECT 41.400 321.600 42.600 338.400 ;
        RECT 50.400 337.050 51.600 361.950 ;
        RECT 53.400 358.050 54.600 367.950 ;
        RECT 59.400 366.900 60.600 367.950 ;
        RECT 58.950 364.800 61.050 366.900 ;
        RECT 52.950 355.950 55.050 358.050 ;
        RECT 46.950 334.950 49.050 337.050 ;
        RECT 49.950 334.950 52.050 337.050 ;
        RECT 52.950 334.950 55.050 337.050 ;
        RECT 47.400 331.050 48.600 334.950 ;
        RECT 53.400 333.900 54.600 334.950 ;
        RECT 59.400 333.900 60.600 364.800 ;
        RECT 65.400 358.050 66.600 403.950 ;
        RECT 86.400 388.050 87.600 451.950 ;
        RECT 92.400 447.900 93.600 450.450 ;
        RECT 92.400 445.800 94.500 447.900 ;
        RECT 95.400 441.600 96.300 454.200 ;
        RECT 101.400 450.900 102.600 453.450 ;
        RECT 101.400 448.800 103.500 450.900 ;
        RECT 97.200 447.900 99.300 448.200 ;
        RECT 105.150 447.900 106.050 454.500 ;
        RECT 112.950 450.600 115.050 451.050 ;
        RECT 116.400 450.600 117.600 496.950 ;
        RECT 112.950 449.400 117.600 450.600 ;
        RECT 112.950 448.950 115.050 449.400 ;
        RECT 97.200 447.000 106.050 447.900 ;
        RECT 97.200 446.100 99.300 447.000 ;
        RECT 102.150 445.200 104.250 446.100 ;
        RECT 97.200 444.000 104.250 445.200 ;
        RECT 97.200 443.100 99.600 444.000 ;
        RECT 94.650 439.500 96.750 441.600 ;
        RECT 98.400 433.050 99.600 443.100 ;
        RECT 101.400 440.100 103.500 442.200 ;
        RECT 105.150 441.900 106.050 447.000 ;
        RECT 106.950 445.800 109.050 447.900 ;
        RECT 107.400 443.400 108.600 445.800 ;
        RECT 97.950 430.950 100.050 433.050 ;
        RECT 101.400 427.050 102.600 440.100 ;
        RECT 104.700 439.800 106.800 441.900 ;
        RECT 113.400 439.050 114.600 448.950 ;
        RECT 119.400 448.050 120.600 499.950 ;
        RECT 127.950 494.100 130.050 496.200 ;
        RECT 133.950 495.000 136.050 499.050 ;
        RECT 128.400 493.050 129.600 494.100 ;
        RECT 134.400 493.050 135.600 495.000 ;
        RECT 142.950 493.950 145.050 496.050 ;
        RECT 148.950 494.100 151.050 496.200 ;
        RECT 154.950 494.100 157.050 496.200 ;
        RECT 127.950 490.950 130.050 493.050 ;
        RECT 130.950 490.950 133.050 493.050 ;
        RECT 133.950 490.950 136.050 493.050 ;
        RECT 136.950 490.950 139.050 493.050 ;
        RECT 131.400 489.900 132.600 490.950 ;
        RECT 130.950 487.800 133.050 489.900 ;
        RECT 137.400 460.050 138.600 490.950 ;
        RECT 136.950 457.950 139.050 460.050 ;
        RECT 127.500 454.500 129.600 456.600 ;
        RECT 118.950 445.950 121.050 448.050 ;
        RECT 124.950 445.950 127.050 448.050 ;
        RECT 127.950 447.300 129.000 454.500 ;
        RECT 131.400 450.900 132.600 453.450 ;
        RECT 137.100 453.300 139.200 455.400 ;
        RECT 130.800 448.800 132.900 450.900 ;
        RECT 133.800 449.700 135.900 451.800 ;
        RECT 133.800 447.300 134.700 449.700 ;
        RECT 127.950 446.100 134.700 447.300 ;
        RECT 125.400 443.400 126.600 445.950 ;
        RECT 127.950 440.700 128.850 446.100 ;
        RECT 129.750 444.300 131.850 445.200 ;
        RECT 137.400 444.300 138.300 453.300 ;
        RECT 143.400 451.200 144.600 493.950 ;
        RECT 149.400 493.050 150.600 494.100 ;
        RECT 155.400 493.050 156.600 494.100 ;
        RECT 160.950 493.950 163.050 496.050 ;
        RECT 148.950 490.950 151.050 493.050 ;
        RECT 151.950 490.950 154.050 493.050 ;
        RECT 154.950 490.950 157.050 493.050 ;
        RECT 152.400 489.900 153.600 490.950 ;
        RECT 161.400 489.900 162.600 493.950 ;
        RECT 170.400 493.050 171.600 499.950 ;
        RECT 169.950 490.950 172.050 493.050 ;
        RECT 172.950 490.950 175.050 493.050 ;
        RECT 173.400 489.900 174.600 490.950 ;
        RECT 179.400 490.050 180.600 514.950 ;
        RECT 184.950 514.500 187.050 516.600 ;
        RECT 194.400 514.050 195.600 535.950 ;
        RECT 197.400 522.900 198.600 547.950 ;
        RECT 211.950 541.950 214.050 544.050 ;
        RECT 205.950 532.950 208.050 535.050 ;
        RECT 206.400 526.050 207.600 532.950 ;
        RECT 202.950 523.950 205.050 526.050 ;
        RECT 205.950 523.950 208.050 526.050 ;
        RECT 203.400 522.900 204.600 523.950 ;
        RECT 196.950 520.800 199.050 522.900 ;
        RECT 202.950 520.800 205.050 522.900 ;
        RECT 212.400 517.050 213.600 541.950 ;
        RECT 202.950 514.950 205.050 517.050 ;
        RECT 211.950 514.950 214.050 517.050 ;
        RECT 193.950 511.950 196.050 514.050 ;
        RECT 184.950 502.950 187.050 505.050 ;
        RECT 193.950 502.950 196.050 505.050 ;
        RECT 181.950 493.950 184.050 496.050 ;
        RECT 151.950 487.800 154.050 489.900 ;
        RECT 160.950 487.800 163.050 489.900 ;
        RECT 172.950 487.800 175.050 489.900 ;
        RECT 178.950 487.950 181.050 490.050 ;
        RECT 175.950 469.950 178.050 472.050 ;
        RECT 145.950 457.950 148.050 460.050 ;
        RECT 140.400 448.050 141.600 450.600 ;
        RECT 142.950 449.100 145.050 451.200 ;
        RECT 139.500 447.150 141.600 448.050 ;
        RECT 139.500 445.950 142.050 447.150 ;
        RECT 129.750 443.100 138.300 444.300 ;
        RECT 112.950 436.950 115.050 439.050 ;
        RECT 127.500 438.600 129.600 440.700 ;
        RECT 130.800 440.100 132.900 442.200 ;
        RECT 134.700 441.300 136.800 443.100 ;
        RECT 139.950 442.800 142.050 445.950 ;
        RECT 131.400 438.900 132.600 440.100 ;
        RECT 130.950 436.800 133.050 438.900 ;
        RECT 146.400 433.050 147.600 457.950 ;
        RECT 154.950 454.950 157.050 457.050 ;
        RECT 155.400 451.200 156.600 454.950 ;
        RECT 154.950 449.100 157.050 451.200 ;
        RECT 155.400 448.050 156.600 449.100 ;
        RECT 176.400 448.050 177.600 469.950 ;
        RECT 154.950 445.950 157.050 448.050 ;
        RECT 157.950 445.950 160.050 448.050 ;
        RECT 169.950 445.950 172.050 448.050 ;
        RECT 175.950 445.950 178.050 448.050 ;
        RECT 151.950 442.950 154.050 445.050 ;
        RECT 158.400 444.900 159.600 445.950 ;
        RECT 145.950 430.950 148.050 433.050 ;
        RECT 100.950 424.950 103.050 427.050 ;
        RECT 109.950 424.950 112.050 427.050 ;
        RECT 88.950 418.950 91.050 421.050 ;
        RECT 89.400 409.050 90.600 418.950 ;
        RECT 91.950 415.950 94.050 421.050 ;
        RECT 97.950 416.100 100.050 418.200 ;
        RECT 103.950 417.000 106.050 421.050 ;
        RECT 106.950 418.950 109.050 424.050 ;
        RECT 98.400 415.050 99.600 416.100 ;
        RECT 104.400 415.050 105.600 417.000 ;
        RECT 94.950 412.950 97.050 415.050 ;
        RECT 97.950 412.950 100.050 415.050 ;
        RECT 100.950 412.950 103.050 415.050 ;
        RECT 103.950 412.950 106.050 415.050 ;
        RECT 95.400 411.600 96.600 412.950 ;
        RECT 101.400 411.900 102.600 412.950 ;
        RECT 110.400 411.900 111.600 424.950 ;
        RECT 136.950 422.400 139.050 424.500 ;
        RECT 118.950 420.600 123.000 421.050 ;
        RECT 118.950 418.950 123.600 420.600 ;
        RECT 122.400 415.050 123.600 418.950 ;
        RECT 112.950 412.950 115.050 415.050 ;
        RECT 118.950 412.950 121.050 415.050 ;
        RECT 121.950 412.950 124.050 415.050 ;
        RECT 124.950 412.950 127.050 415.050 ;
        RECT 133.950 412.950 136.050 415.050 ;
        RECT 92.400 410.400 96.600 411.600 ;
        RECT 88.950 406.950 91.050 409.050 ;
        RECT 92.400 406.050 93.600 410.400 ;
        RECT 100.950 409.800 103.050 411.900 ;
        RECT 109.950 409.800 112.050 411.900 ;
        RECT 113.400 409.050 114.600 412.950 ;
        RECT 119.400 411.000 120.600 412.950 ;
        RECT 94.950 406.950 97.050 409.050 ;
        RECT 112.950 406.950 115.050 409.050 ;
        RECT 118.950 406.950 121.050 411.000 ;
        RECT 88.950 403.800 91.050 405.900 ;
        RECT 91.950 403.950 94.050 406.050 ;
        RECT 89.400 391.050 90.600 403.800 ;
        RECT 88.950 388.950 91.050 391.050 ;
        RECT 70.950 385.950 73.050 388.050 ;
        RECT 85.950 385.950 88.050 388.050 ;
        RECT 67.950 376.950 70.050 379.050 ;
        RECT 68.400 367.050 69.600 376.950 ;
        RECT 71.400 373.050 72.600 385.950 ;
        RECT 88.950 381.300 91.050 383.400 ;
        RECT 79.950 376.950 82.050 379.050 ;
        RECT 89.850 377.700 91.050 381.300 ;
        RECT 70.950 370.950 73.050 373.050 ;
        RECT 73.950 371.100 76.050 373.200 ;
        RECT 74.400 370.050 75.600 371.100 ;
        RECT 80.400 370.050 81.600 376.950 ;
        RECT 88.950 375.600 91.050 377.700 ;
        RECT 73.950 367.950 76.050 370.050 ;
        RECT 76.950 367.950 79.050 370.050 ;
        RECT 79.950 367.950 82.050 370.050 ;
        RECT 85.950 367.950 88.050 370.050 ;
        RECT 67.950 364.950 70.050 367.050 ;
        RECT 67.950 361.800 70.050 363.900 ;
        RECT 64.950 355.950 67.050 358.050 ;
        RECT 52.950 331.800 55.050 333.900 ;
        RECT 58.950 331.800 61.050 333.900 ;
        RECT 46.950 328.950 49.050 331.050 ;
        RECT 41.400 320.400 45.600 321.600 ;
        RECT 40.950 316.950 43.050 319.050 ;
        RECT 1.950 304.950 4.050 307.050 ;
        RECT 13.950 304.950 16.050 307.050 ;
        RECT 14.400 292.050 15.600 304.950 ;
        RECT 13.950 289.950 16.050 292.050 ;
        RECT 13.950 256.950 16.050 259.050 ;
        RECT 14.400 229.050 15.600 256.950 ;
        RECT 22.950 229.950 25.050 232.050 ;
        RECT 13.950 226.950 16.050 229.050 ;
        RECT 7.950 224.400 10.050 226.500 ;
        RECT 4.950 220.950 7.050 223.050 ;
        RECT 5.400 214.050 6.600 220.950 ;
        RECT 4.950 211.950 7.050 214.050 ;
        RECT 8.700 204.600 9.900 224.400 ;
        RECT 14.400 223.050 15.600 226.950 ;
        RECT 13.950 220.950 16.050 223.050 ;
        RECT 13.950 215.400 16.050 217.500 ;
        RECT 14.400 214.050 15.600 215.400 ;
        RECT 13.950 211.950 16.050 214.050 ;
        RECT 16.950 208.950 19.050 211.050 ;
        RECT 7.950 202.500 10.050 204.600 ;
        RECT 17.400 181.050 18.600 208.950 ;
        RECT 23.400 193.050 24.600 229.950 ;
        RECT 28.950 225.300 31.050 227.400 ;
        RECT 28.950 221.700 30.150 225.300 ;
        RECT 28.950 219.600 31.050 221.700 ;
        RECT 28.950 204.600 30.150 219.600 ;
        RECT 31.950 211.950 34.050 214.050 ;
        RECT 32.400 210.600 33.600 211.950 ;
        RECT 31.950 208.500 34.050 210.600 ;
        RECT 28.950 202.500 31.050 204.600 ;
        RECT 34.950 202.950 37.050 205.050 ;
        RECT 35.400 196.050 36.600 202.950 ;
        RECT 41.400 199.050 42.600 316.950 ;
        RECT 44.400 286.050 45.600 320.400 ;
        RECT 47.400 292.050 48.600 328.950 ;
        RECT 64.950 322.950 67.050 325.050 ;
        RECT 50.400 297.000 60.600 297.600 ;
        RECT 49.950 296.400 60.600 297.000 ;
        RECT 49.950 292.950 52.050 296.400 ;
        RECT 52.950 293.100 55.050 295.200 ;
        RECT 53.400 292.050 54.600 293.100 ;
        RECT 59.400 292.050 60.600 296.400 ;
        RECT 65.400 292.050 66.600 322.950 ;
        RECT 68.400 294.600 69.600 361.800 ;
        RECT 77.400 358.050 78.600 367.950 ;
        RECT 82.950 364.950 85.050 367.050 ;
        RECT 86.400 366.600 87.600 367.950 ;
        RECT 76.950 355.950 79.050 358.050 ;
        RECT 76.950 339.000 79.050 343.050 ;
        RECT 77.400 337.050 78.600 339.000 ;
        RECT 83.400 337.050 84.600 364.950 ;
        RECT 85.950 364.500 88.050 366.600 ;
        RECT 89.850 360.600 91.050 375.600 ;
        RECT 95.400 373.050 96.600 406.950 ;
        RECT 103.950 388.950 106.050 391.050 ;
        RECT 97.950 379.950 100.050 382.050 ;
        RECT 94.950 370.950 97.050 373.050 ;
        RECT 88.950 358.500 91.050 360.600 ;
        RECT 98.400 339.600 99.600 379.950 ;
        RECT 104.400 370.050 105.600 388.950 ;
        RECT 109.950 380.400 112.050 382.500 ;
        RECT 103.950 367.950 106.050 370.050 ;
        RECT 110.100 360.600 111.300 380.400 ;
        RECT 112.950 372.000 115.050 376.050 ;
        RECT 113.400 370.050 114.600 372.000 ;
        RECT 112.950 367.950 115.050 370.050 ;
        RECT 109.950 358.500 112.050 360.600 ;
        RECT 95.400 338.400 99.600 339.600 ;
        RECT 73.950 334.950 76.050 337.050 ;
        RECT 76.950 334.950 79.050 337.050 ;
        RECT 79.950 334.950 82.050 337.050 ;
        RECT 82.950 334.950 85.050 337.050 ;
        RECT 85.950 334.950 88.050 337.050 ;
        RECT 74.400 333.900 75.600 334.950 ;
        RECT 73.950 331.800 76.050 333.900 ;
        RECT 74.400 328.050 75.600 331.800 ;
        RECT 80.400 330.600 81.600 334.950 ;
        RECT 77.400 329.400 81.600 330.600 ;
        RECT 73.950 325.950 76.050 328.050 ;
        RECT 77.400 322.050 78.600 329.400 ;
        RECT 79.950 325.950 82.050 328.050 ;
        RECT 76.950 319.950 79.050 322.050 ;
        RECT 73.950 313.950 76.050 316.050 ;
        RECT 70.950 295.950 73.050 301.050 ;
        RECT 68.400 293.400 72.600 294.600 ;
        RECT 46.950 289.950 49.050 292.050 ;
        RECT 52.950 289.950 55.050 292.050 ;
        RECT 55.950 289.950 58.050 292.050 ;
        RECT 58.950 289.950 61.050 292.050 ;
        RECT 61.950 289.950 64.050 292.050 ;
        RECT 64.950 289.950 67.050 292.050 ;
        RECT 56.400 288.900 57.600 289.950 ;
        RECT 46.950 286.800 49.050 288.900 ;
        RECT 55.950 286.800 58.050 288.900 ;
        RECT 62.400 288.000 63.600 289.950 ;
        RECT 43.950 283.950 46.050 286.050 ;
        RECT 43.950 250.950 46.050 253.050 ;
        RECT 44.400 210.600 45.600 250.950 ;
        RECT 47.400 216.600 48.600 286.800 ;
        RECT 61.950 283.950 64.050 288.000 ;
        RECT 71.400 286.050 72.600 293.400 ;
        RECT 70.950 283.950 73.050 286.050 ;
        RECT 67.950 280.950 70.050 283.050 ;
        RECT 61.950 268.950 64.050 271.050 ;
        RECT 55.950 260.100 58.050 262.200 ;
        RECT 56.400 259.050 57.600 260.100 ;
        RECT 62.400 259.050 63.600 268.950 ;
        RECT 52.950 256.950 55.050 259.050 ;
        RECT 55.950 256.950 58.050 259.050 ;
        RECT 58.950 256.950 61.050 259.050 ;
        RECT 61.950 256.950 64.050 259.050 ;
        RECT 49.950 253.950 52.050 256.050 ;
        RECT 50.400 220.050 51.600 253.950 ;
        RECT 53.400 238.050 54.600 256.950 ;
        RECT 59.400 255.000 60.600 256.950 ;
        RECT 58.950 250.950 61.050 255.000 ;
        RECT 52.950 235.950 55.050 238.050 ;
        RECT 64.950 235.950 67.050 238.050 ;
        RECT 49.950 217.950 52.050 220.050 ;
        RECT 47.400 215.400 51.600 216.600 ;
        RECT 55.950 216.000 58.050 220.050 ;
        RECT 50.400 214.050 51.600 215.400 ;
        RECT 56.400 214.050 57.600 216.000 ;
        RECT 49.950 211.950 52.050 214.050 ;
        RECT 52.950 211.950 55.050 214.050 ;
        RECT 55.950 211.950 58.050 214.050 ;
        RECT 58.950 211.950 61.050 214.050 ;
        RECT 43.950 208.500 46.050 210.600 ;
        RECT 40.950 196.950 43.050 199.050 ;
        RECT 28.950 193.950 31.050 196.050 ;
        RECT 34.950 193.950 37.050 196.050 ;
        RECT 22.950 190.950 25.050 193.050 ;
        RECT 23.400 181.050 24.600 190.950 ;
        RECT 13.950 178.950 16.050 181.050 ;
        RECT 16.950 178.950 19.050 181.050 ;
        RECT 19.950 178.950 22.050 181.050 ;
        RECT 22.950 178.950 25.050 181.050 ;
        RECT 14.400 177.900 15.600 178.950 ;
        RECT 13.950 175.800 16.050 177.900 ;
        RECT 20.400 142.050 21.600 178.950 ;
        RECT 19.950 139.950 22.050 142.050 ;
        RECT 19.950 133.950 22.050 136.050 ;
        RECT 20.400 133.050 21.600 133.950 ;
        RECT 29.400 133.050 30.600 193.950 ;
        RECT 37.950 182.100 40.050 184.200 ;
        RECT 44.400 184.050 45.600 208.500 ;
        RECT 53.400 205.050 54.600 211.950 ;
        RECT 59.400 210.900 60.600 211.950 ;
        RECT 58.950 208.800 61.050 210.900 ;
        RECT 65.400 208.050 66.600 235.950 ;
        RECT 68.400 223.050 69.600 280.950 ;
        RECT 74.400 262.200 75.600 313.950 ;
        RECT 76.950 307.950 79.050 310.050 ;
        RECT 77.400 295.050 78.600 307.950 ;
        RECT 80.400 295.200 81.600 325.950 ;
        RECT 86.400 325.050 87.600 334.950 ;
        RECT 95.400 333.900 96.600 338.400 ;
        RECT 103.950 338.100 106.050 340.200 ;
        RECT 104.400 337.050 105.600 338.100 ;
        RECT 112.950 337.950 115.050 340.050 ;
        RECT 115.950 337.950 118.050 340.050 ;
        RECT 100.950 334.950 103.050 337.050 ;
        RECT 103.950 334.950 106.050 337.050 ;
        RECT 106.950 334.950 109.050 337.050 ;
        RECT 94.950 331.800 97.050 333.900 ;
        RECT 85.950 322.950 88.050 325.050 ;
        RECT 91.950 322.950 94.050 325.050 ;
        RECT 85.950 298.950 88.050 301.050 ;
        RECT 76.950 292.950 79.050 295.050 ;
        RECT 79.950 293.100 82.050 295.200 ;
        RECT 80.400 292.050 81.600 293.100 ;
        RECT 86.400 292.050 87.600 298.950 ;
        RECT 92.400 292.050 93.600 322.950 ;
        RECT 101.400 310.050 102.600 334.950 ;
        RECT 107.400 333.900 108.600 334.950 ;
        RECT 106.950 331.800 109.050 333.900 ;
        RECT 100.950 307.950 103.050 310.050 ;
        RECT 109.950 307.950 112.050 310.050 ;
        RECT 100.950 303.300 103.050 305.400 ;
        RECT 101.850 299.700 103.050 303.300 ;
        RECT 100.950 297.600 103.050 299.700 ;
        RECT 79.950 289.950 82.050 292.050 ;
        RECT 82.950 289.950 85.050 292.050 ;
        RECT 85.950 289.950 88.050 292.050 ;
        RECT 88.950 289.950 91.050 292.050 ;
        RECT 91.950 289.950 94.050 292.050 ;
        RECT 97.950 289.950 100.050 292.050 ;
        RECT 76.950 283.950 79.050 289.050 ;
        RECT 83.400 288.000 84.600 289.950 ;
        RECT 89.400 288.900 90.600 289.950 ;
        RECT 82.950 283.950 85.050 288.000 ;
        RECT 88.950 286.800 91.050 288.900 ;
        RECT 98.400 288.600 99.600 289.950 ;
        RECT 97.950 286.500 100.050 288.600 ;
        RECT 101.850 282.600 103.050 297.600 ;
        RECT 106.950 292.950 109.050 295.050 ;
        RECT 100.950 280.500 103.050 282.600 ;
        RECT 100.950 268.950 103.050 271.050 ;
        RECT 73.950 260.100 76.050 262.200 ;
        RECT 85.950 260.100 88.050 262.200 ;
        RECT 86.400 259.050 87.600 260.100 ;
        RECT 101.400 259.050 102.600 268.950 ;
        RECT 107.400 262.050 108.600 292.950 ;
        RECT 110.400 262.200 111.600 307.950 ;
        RECT 113.400 294.600 114.600 337.950 ;
        RECT 116.400 333.900 117.600 337.950 ;
        RECT 115.950 331.800 118.050 333.900 ;
        RECT 119.400 310.050 120.600 406.950 ;
        RECT 125.400 403.050 126.600 412.950 ;
        RECT 134.400 411.000 135.600 412.950 ;
        RECT 127.950 406.950 130.050 409.050 ;
        RECT 133.950 406.950 136.050 411.000 ;
        RECT 124.950 400.950 127.050 403.050 ;
        RECT 124.950 397.800 127.050 399.900 ;
        RECT 121.950 370.950 124.050 373.050 ;
        RECT 122.400 349.050 123.600 370.950 ;
        RECT 125.400 361.050 126.600 397.800 ;
        RECT 128.400 376.050 129.600 406.950 ;
        RECT 137.700 402.600 138.900 422.400 ;
        RECT 148.950 421.950 151.050 424.050 ;
        RECT 142.950 412.950 145.050 415.050 ;
        RECT 143.400 411.600 144.600 412.950 ;
        RECT 149.400 412.050 150.600 421.950 ;
        RECT 152.400 418.500 153.600 442.950 ;
        RECT 157.950 442.800 160.050 444.900 ;
        RECT 170.400 442.050 171.600 445.950 ;
        RECT 169.950 439.950 172.050 442.050 ;
        RECT 157.950 422.400 160.050 424.500 ;
        RECT 151.950 416.400 154.050 418.500 ;
        RECT 142.950 409.500 145.050 411.600 ;
        RECT 148.950 409.950 151.050 412.050 ;
        RECT 157.950 407.400 159.150 422.400 ;
        RECT 160.950 416.400 163.050 418.500 ;
        RECT 161.400 415.050 162.600 416.400 ;
        RECT 160.950 412.950 163.050 415.050 ;
        RECT 163.950 409.800 166.050 411.900 ;
        RECT 157.950 405.300 160.050 407.400 ;
        RECT 136.950 400.500 139.050 402.600 ;
        RECT 157.950 401.700 159.150 405.300 ;
        RECT 157.950 399.600 160.050 401.700 ;
        RECT 142.950 376.950 145.050 379.050 ;
        RECT 127.950 373.950 130.050 376.050 ;
        RECT 130.950 371.100 133.050 373.200 ;
        RECT 131.400 370.050 132.600 371.100 ;
        RECT 130.950 367.950 133.050 370.050 ;
        RECT 136.950 367.950 139.050 370.050 ;
        RECT 137.400 366.600 138.600 367.950 ;
        RECT 137.400 365.400 141.600 366.600 ;
        RECT 140.400 361.050 141.600 365.400 ;
        RECT 124.950 358.950 127.050 361.050 ;
        RECT 139.950 358.950 142.050 361.050 ;
        RECT 121.950 346.950 124.050 349.050 ;
        RECT 133.950 346.950 136.050 349.050 ;
        RECT 121.950 337.950 124.050 343.050 ;
        RECT 127.950 338.100 130.050 340.200 ;
        RECT 128.400 337.050 129.600 338.100 ;
        RECT 134.400 337.050 135.600 346.950 ;
        RECT 124.950 334.950 127.050 337.050 ;
        RECT 127.950 334.950 130.050 337.050 ;
        RECT 130.950 334.950 133.050 337.050 ;
        RECT 133.950 334.950 136.050 337.050 ;
        RECT 125.400 333.900 126.600 334.950 ;
        RECT 131.400 333.900 132.600 334.950 ;
        RECT 124.950 331.800 127.050 333.900 ;
        RECT 130.950 331.800 133.050 333.900 ;
        RECT 140.400 316.050 141.600 358.950 ;
        RECT 139.950 313.950 142.050 316.050 ;
        RECT 118.950 307.950 121.050 310.050 ;
        RECT 121.950 302.400 124.050 304.500 ;
        RECT 113.400 293.400 117.600 294.600 ;
        RECT 116.400 292.050 117.600 293.400 ;
        RECT 115.950 289.950 118.050 292.050 ;
        RECT 122.100 282.600 123.300 302.400 ;
        RECT 127.950 301.950 130.050 304.050 ;
        RECT 136.950 302.400 139.050 304.500 ;
        RECT 143.400 304.050 144.600 376.950 ;
        RECT 145.950 370.950 148.050 373.050 ;
        RECT 154.950 371.100 157.050 373.200 ;
        RECT 146.400 343.050 147.600 370.950 ;
        RECT 155.400 370.050 156.600 371.100 ;
        RECT 151.950 367.950 154.050 370.050 ;
        RECT 154.950 367.950 157.050 370.050 ;
        RECT 157.950 367.950 160.050 370.050 ;
        RECT 152.400 358.050 153.600 367.950 ;
        RECT 158.400 366.000 159.600 367.950 ;
        RECT 157.950 361.950 160.050 366.000 ;
        RECT 151.950 355.950 154.050 358.050 ;
        RECT 145.950 340.950 148.050 343.050 ;
        RECT 160.950 340.950 163.050 343.050 ;
        RECT 151.950 338.100 154.050 340.200 ;
        RECT 152.400 337.050 153.600 338.100 ;
        RECT 148.950 334.950 151.050 337.050 ;
        RECT 151.950 334.950 154.050 337.050 ;
        RECT 154.950 334.950 157.050 337.050 ;
        RECT 149.400 333.000 150.600 334.950 ;
        RECT 148.950 328.950 151.050 333.000 ;
        RECT 148.950 322.950 151.050 325.050 ;
        RECT 128.400 294.600 129.600 301.950 ;
        RECT 125.400 293.400 129.600 294.600 ;
        RECT 133.950 294.000 136.050 298.050 ;
        RECT 125.400 292.050 126.600 293.400 ;
        RECT 134.400 292.050 135.600 294.000 ;
        RECT 124.950 289.950 127.050 292.050 ;
        RECT 133.950 289.950 136.050 292.050 ;
        RECT 137.700 282.600 138.900 302.400 ;
        RECT 142.950 301.950 145.050 304.050 ;
        RECT 142.950 293.400 145.050 295.500 ;
        RECT 143.400 292.050 144.600 293.400 ;
        RECT 142.950 289.950 145.050 292.050 ;
        RECT 121.950 280.500 124.050 282.600 ;
        RECT 136.950 280.500 139.050 282.600 ;
        RECT 149.400 280.050 150.600 322.950 ;
        RECT 155.400 322.050 156.600 334.950 ;
        RECT 161.400 331.050 162.600 340.950 ;
        RECT 164.400 340.050 165.600 409.800 ;
        RECT 170.400 400.050 171.600 439.950 ;
        RECT 182.400 439.050 183.600 493.950 ;
        RECT 185.400 484.050 186.600 502.950 ;
        RECT 194.400 493.050 195.600 502.950 ;
        RECT 199.950 493.950 202.050 499.050 ;
        RECT 190.950 490.950 193.050 493.050 ;
        RECT 193.950 490.950 196.050 493.050 ;
        RECT 196.950 490.950 199.050 493.050 ;
        RECT 187.950 487.950 190.050 490.050 ;
        RECT 191.400 489.900 192.600 490.950 ;
        RECT 184.950 481.950 187.050 484.050 ;
        RECT 184.950 449.100 187.050 451.200 ;
        RECT 172.950 436.950 175.050 439.050 ;
        RECT 181.950 436.950 184.050 439.050 ;
        RECT 169.950 397.950 172.050 400.050 ;
        RECT 173.400 382.050 174.600 436.950 ;
        RECT 185.400 436.050 186.600 449.100 ;
        RECT 188.400 439.050 189.600 487.950 ;
        RECT 190.950 487.800 193.050 489.900 ;
        RECT 197.400 478.050 198.600 490.950 ;
        RECT 203.400 487.050 204.600 514.950 ;
        RECT 215.400 502.050 216.600 586.950 ;
        RECT 226.950 578.400 229.050 580.500 ;
        RECT 220.950 568.950 223.050 571.050 ;
        RECT 221.400 532.050 222.600 568.950 ;
        RECT 227.100 558.600 228.300 578.400 ;
        RECT 233.400 573.600 234.600 619.950 ;
        RECT 236.400 610.050 237.600 650.400 ;
        RECT 239.400 640.050 240.600 652.950 ;
        RECT 244.950 650.100 247.050 652.200 ;
        RECT 250.950 651.000 253.050 655.050 ;
        RECT 268.950 651.000 271.050 655.050 ;
        RECT 245.400 649.050 246.600 650.100 ;
        RECT 251.400 649.050 252.600 651.000 ;
        RECT 269.400 649.050 270.600 651.000 ;
        RECT 275.400 649.050 276.600 658.950 ;
        RECT 244.950 646.950 247.050 649.050 ;
        RECT 247.950 646.950 250.050 649.050 ;
        RECT 250.950 646.950 253.050 649.050 ;
        RECT 253.950 646.950 256.050 649.050 ;
        RECT 265.950 646.950 268.050 649.050 ;
        RECT 268.950 646.950 271.050 649.050 ;
        RECT 271.950 646.950 274.050 649.050 ;
        RECT 274.950 646.950 277.050 649.050 ;
        RECT 238.950 637.950 241.050 640.050 ;
        RECT 248.400 634.050 249.600 646.950 ;
        RECT 254.400 645.900 255.600 646.950 ;
        RECT 253.950 643.800 256.050 645.900 ;
        RECT 266.400 634.050 267.600 646.950 ;
        RECT 272.400 645.900 273.600 646.950 ;
        RECT 271.950 643.800 274.050 645.900 ;
        RECT 247.950 631.950 250.050 634.050 ;
        RECT 265.950 631.950 268.050 634.050 ;
        RECT 284.400 622.050 285.600 683.100 ;
        RECT 296.400 682.050 297.600 683.100 ;
        RECT 292.950 679.950 295.050 682.050 ;
        RECT 295.950 679.950 298.050 682.050 ;
        RECT 289.950 673.950 292.050 676.050 ;
        RECT 286.950 652.950 289.050 655.050 ;
        RECT 287.400 645.900 288.600 652.950 ;
        RECT 286.950 643.800 289.050 645.900 ;
        RECT 283.950 619.950 286.050 622.050 ;
        RECT 290.400 616.050 291.600 673.950 ;
        RECT 293.400 670.050 294.600 679.950 ;
        RECT 302.400 676.050 303.600 683.100 ;
        RECT 305.400 679.050 306.600 689.400 ;
        RECT 311.400 682.050 312.600 691.950 ;
        RECT 316.950 683.100 319.050 685.200 ;
        RECT 317.400 682.050 318.600 683.100 ;
        RECT 310.950 679.950 313.050 682.050 ;
        RECT 313.950 679.950 316.050 682.050 ;
        RECT 316.950 679.950 319.050 682.050 ;
        RECT 304.950 676.950 307.050 679.050 ;
        RECT 314.400 678.900 315.600 679.950 ;
        RECT 313.950 676.800 316.050 678.900 ;
        RECT 301.950 673.950 304.050 676.050 ;
        RECT 292.950 667.950 295.050 670.050 ;
        RECT 313.950 667.950 316.050 670.050 ;
        RECT 293.400 652.050 294.600 667.950 ;
        RECT 304.950 664.950 307.050 667.050 ;
        RECT 292.950 649.950 295.050 652.050 ;
        RECT 298.950 651.000 301.050 655.050 ;
        RECT 299.400 649.050 300.600 651.000 ;
        RECT 305.400 649.050 306.600 664.950 ;
        RECT 314.400 661.050 315.600 667.950 ;
        RECT 323.400 667.050 324.600 694.950 ;
        RECT 325.950 691.950 328.050 694.050 ;
        RECT 322.950 664.950 325.050 667.050 ;
        RECT 326.400 664.050 327.600 691.950 ;
        RECT 329.400 688.050 330.600 697.950 ;
        RECT 331.950 691.950 334.050 694.050 ;
        RECT 328.950 685.950 331.050 688.050 ;
        RECT 332.400 682.050 333.600 691.950 ;
        RECT 356.400 685.200 357.600 700.950 ;
        RECT 359.400 690.600 360.600 728.100 ;
        RECT 362.400 694.050 363.600 784.950 ;
        RECT 365.400 763.050 366.600 817.950 ;
        RECT 371.400 805.050 372.600 829.950 ;
        RECT 374.400 820.050 375.600 841.950 ;
        RECT 377.400 841.050 378.600 865.950 ;
        RECT 385.950 844.950 388.050 847.050 ;
        RECT 394.950 844.950 397.050 847.050 ;
        RECT 376.950 838.950 379.050 841.050 ;
        RECT 379.950 840.000 382.050 844.050 ;
        RECT 380.400 838.050 381.600 840.000 ;
        RECT 386.400 838.050 387.600 844.950 ;
        RECT 379.950 835.950 382.050 838.050 ;
        RECT 382.950 835.950 385.050 838.050 ;
        RECT 385.950 835.950 388.050 838.050 ;
        RECT 388.950 835.950 391.050 838.050 ;
        RECT 383.400 834.900 384.600 835.950 ;
        RECT 389.400 834.900 390.600 835.950 ;
        RECT 382.950 832.800 385.050 834.900 ;
        RECT 388.950 832.800 391.050 834.900 ;
        RECT 395.400 829.050 396.600 844.950 ;
        RECT 397.950 841.950 400.050 844.050 ;
        RECT 398.400 832.050 399.600 841.950 ;
        RECT 406.950 839.100 409.050 841.200 ;
        RECT 412.950 840.000 415.050 844.050 ;
        RECT 407.400 838.050 408.600 839.100 ;
        RECT 413.400 838.050 414.600 840.000 ;
        RECT 403.950 835.950 406.050 838.050 ;
        RECT 406.950 835.950 409.050 838.050 ;
        RECT 409.950 835.950 412.050 838.050 ;
        RECT 412.950 835.950 415.050 838.050 ;
        RECT 400.950 832.950 403.050 835.050 ;
        RECT 397.950 829.950 400.050 832.050 ;
        RECT 394.950 826.950 397.050 829.050 ;
        RECT 397.950 820.950 400.050 823.050 ;
        RECT 373.950 817.950 376.050 820.050 ;
        RECT 388.950 817.950 391.050 820.050 ;
        RECT 376.950 814.950 379.050 817.050 ;
        RECT 377.400 805.050 378.600 814.950 ;
        RECT 385.950 806.100 388.050 808.200 ;
        RECT 370.950 802.950 373.050 805.050 ;
        RECT 373.950 802.950 376.050 805.050 ;
        RECT 376.950 802.950 379.050 805.050 ;
        RECT 379.950 802.950 382.050 805.050 ;
        RECT 374.400 796.050 375.600 802.950 ;
        RECT 380.400 801.000 381.600 802.950 ;
        RECT 379.950 796.950 382.050 801.000 ;
        RECT 373.950 793.950 376.050 796.050 ;
        RECT 374.400 778.050 375.600 793.950 ;
        RECT 373.950 775.950 376.050 778.050 ;
        RECT 382.950 775.950 385.050 778.050 ;
        RECT 373.950 769.950 376.050 772.050 ;
        RECT 364.950 760.950 367.050 763.050 ;
        RECT 367.950 762.000 370.050 766.050 ;
        RECT 368.400 760.050 369.600 762.000 ;
        RECT 374.400 760.050 375.600 769.950 ;
        RECT 367.950 757.950 370.050 760.050 ;
        RECT 370.950 757.950 373.050 760.050 ;
        RECT 373.950 757.950 376.050 760.050 ;
        RECT 376.950 757.950 379.050 760.050 ;
        RECT 371.400 756.900 372.600 757.950 ;
        RECT 370.950 754.800 373.050 756.900 ;
        RECT 373.950 748.950 376.050 751.050 ;
        RECT 367.950 728.100 370.050 730.200 ;
        RECT 368.400 727.050 369.600 728.100 ;
        RECT 374.400 727.050 375.600 748.950 ;
        RECT 377.400 736.050 378.600 757.950 ;
        RECT 376.950 733.950 379.050 736.050 ;
        RECT 367.950 724.950 370.050 727.050 ;
        RECT 370.950 724.950 373.050 727.050 ;
        RECT 373.950 724.950 376.050 727.050 ;
        RECT 376.950 724.950 379.050 727.050 ;
        RECT 371.400 723.900 372.600 724.950 ;
        RECT 370.950 721.800 373.050 723.900 ;
        RECT 371.400 712.050 372.600 721.800 ;
        RECT 377.400 718.050 378.600 724.950 ;
        RECT 376.950 715.950 379.050 718.050 ;
        RECT 383.400 715.050 384.600 775.950 ;
        RECT 386.400 772.050 387.600 806.100 ;
        RECT 389.400 802.050 390.600 817.950 ;
        RECT 398.400 805.050 399.600 820.950 ;
        RECT 401.400 820.050 402.600 832.950 ;
        RECT 400.950 817.950 403.050 820.050 ;
        RECT 404.400 808.200 405.600 835.950 ;
        RECT 406.950 829.950 409.050 832.050 ;
        RECT 407.400 825.600 408.600 829.950 ;
        RECT 410.400 829.050 411.600 835.950 ;
        RECT 409.950 826.950 412.050 829.050 ;
        RECT 407.400 824.400 411.600 825.600 ;
        RECT 403.950 806.100 406.050 808.200 ;
        RECT 404.400 805.050 405.600 806.100 ;
        RECT 394.950 802.950 397.050 805.050 ;
        RECT 397.950 802.950 400.050 805.050 ;
        RECT 400.950 802.950 403.050 805.050 ;
        RECT 403.950 802.950 406.050 805.050 ;
        RECT 388.950 799.950 391.050 802.050 ;
        RECT 395.400 799.050 396.600 802.950 ;
        RECT 401.400 801.900 402.600 802.950 ;
        RECT 400.950 799.800 403.050 801.900 ;
        RECT 394.950 796.950 397.050 799.050 ;
        RECT 388.950 790.950 391.050 793.050 ;
        RECT 385.950 769.950 388.050 772.050 ;
        RECT 389.400 736.050 390.600 790.950 ;
        RECT 395.400 760.050 396.600 796.950 ;
        RECT 401.400 778.050 402.600 799.800 ;
        RECT 410.400 781.050 411.600 824.400 ;
        RECT 415.950 811.950 418.050 814.050 ;
        RECT 416.400 808.050 417.600 811.950 ;
        RECT 415.950 805.950 418.050 808.050 ;
        RECT 422.400 805.050 423.600 868.950 ;
        RECT 431.400 856.050 432.600 877.950 ;
        RECT 442.950 874.950 445.050 879.900 ;
        RECT 448.950 877.800 451.050 879.900 ;
        RECT 455.400 874.050 456.600 884.100 ;
        RECT 464.400 883.050 465.600 884.100 ;
        RECT 470.400 883.050 471.600 884.100 ;
        RECT 475.800 883.950 477.900 886.050 ;
        RECT 478.950 884.100 481.050 886.200 ;
        RECT 484.950 884.100 487.050 886.200 ;
        RECT 460.950 880.950 463.050 883.050 ;
        RECT 463.950 880.950 466.050 883.050 ;
        RECT 466.950 880.950 469.050 883.050 ;
        RECT 469.950 880.950 472.050 883.050 ;
        RECT 461.400 879.900 462.600 880.950 ;
        RECT 460.950 877.800 463.050 879.900 ;
        RECT 467.400 879.000 468.600 880.950 ;
        RECT 476.400 879.900 477.600 883.950 ;
        RECT 448.950 871.950 451.050 874.050 ;
        RECT 454.950 871.950 457.050 874.050 ;
        RECT 427.800 853.950 429.900 856.050 ;
        RECT 430.950 853.950 433.050 856.050 ;
        RECT 439.950 853.950 442.050 856.050 ;
        RECT 428.400 841.050 429.600 853.950 ;
        RECT 433.950 844.950 436.050 847.050 ;
        RECT 427.950 838.950 430.050 841.050 ;
        RECT 434.400 838.050 435.600 844.950 ;
        RECT 440.400 838.050 441.600 853.950 ;
        RECT 445.950 839.100 448.050 841.200 ;
        RECT 430.950 835.950 433.050 838.050 ;
        RECT 433.950 835.950 436.050 838.050 ;
        RECT 436.950 835.950 439.050 838.050 ;
        RECT 439.950 835.950 442.050 838.050 ;
        RECT 431.400 834.900 432.600 835.950 ;
        RECT 437.400 834.900 438.600 835.950 ;
        RECT 430.950 832.800 433.050 834.900 ;
        RECT 436.950 832.800 439.050 834.900 ;
        RECT 442.950 829.950 445.050 834.900 ;
        RECT 439.950 826.950 442.050 829.050 ;
        RECT 430.950 817.950 433.050 820.050 ;
        RECT 418.950 802.950 421.050 805.050 ;
        RECT 421.950 802.950 424.050 805.050 ;
        RECT 424.950 802.950 427.050 805.050 ;
        RECT 419.400 801.900 420.600 802.950 ;
        RECT 418.950 799.800 421.050 801.900 ;
        RECT 425.400 781.050 426.600 802.950 ;
        RECT 403.950 778.950 406.050 781.050 ;
        RECT 409.950 778.950 412.050 781.050 ;
        RECT 424.950 778.950 427.050 781.050 ;
        RECT 400.950 775.950 403.050 778.050 ;
        RECT 394.950 757.950 397.050 760.050 ;
        RECT 397.950 757.950 400.050 760.050 ;
        RECT 398.400 756.900 399.600 757.950 ;
        RECT 404.400 757.050 405.600 778.950 ;
        RECT 424.950 769.950 427.050 772.050 ;
        RECT 425.400 763.200 426.600 769.950 ;
        RECT 406.950 762.600 411.000 763.050 ;
        RECT 406.950 760.950 411.600 762.600 ;
        RECT 424.950 761.100 427.050 763.200 ;
        RECT 431.400 762.600 432.600 817.950 ;
        RECT 433.950 806.100 436.050 808.200 ;
        RECT 434.400 790.050 435.600 806.100 ;
        RECT 440.400 805.050 441.600 826.950 ;
        RECT 446.400 826.050 447.600 839.100 ;
        RECT 449.400 832.050 450.600 871.950 ;
        RECT 461.400 852.600 462.600 877.800 ;
        RECT 466.950 874.950 469.050 879.000 ;
        RECT 475.950 877.800 478.050 879.900 ;
        RECT 463.950 852.600 466.050 853.050 ;
        RECT 461.400 851.400 466.050 852.600 ;
        RECT 463.950 850.950 466.050 851.400 ;
        RECT 457.950 839.100 460.050 841.200 ;
        RECT 458.400 838.050 459.600 839.100 ;
        RECT 464.400 838.050 465.600 850.950 ;
        RECT 467.400 841.200 468.600 874.950 ;
        RECT 479.400 871.050 480.600 884.100 ;
        RECT 485.400 883.050 486.600 884.100 ;
        RECT 491.400 883.050 492.600 889.950 ;
        RECT 499.950 883.950 502.050 886.050 ;
        RECT 508.950 884.100 511.050 886.200 ;
        RECT 484.950 880.950 487.050 883.050 ;
        RECT 487.950 880.950 490.050 883.050 ;
        RECT 490.950 880.950 493.050 883.050 ;
        RECT 493.950 880.950 496.050 883.050 ;
        RECT 488.400 879.900 489.600 880.950 ;
        RECT 487.950 877.800 490.050 879.900 ;
        RECT 494.400 879.000 495.600 880.950 ;
        RECT 493.950 874.950 496.050 879.000 ;
        RECT 500.400 877.050 501.600 883.950 ;
        RECT 509.400 883.050 510.600 884.100 ;
        RECT 520.950 883.950 523.050 886.050 ;
        RECT 529.950 884.100 532.050 886.200 ;
        RECT 535.950 884.100 538.050 886.200 ;
        RECT 508.950 880.950 511.050 883.050 ;
        RECT 511.950 880.950 514.050 883.050 ;
        RECT 512.400 879.900 513.600 880.950 ;
        RECT 511.950 877.800 514.050 879.900 ;
        RECT 499.950 874.950 502.050 877.050 ;
        RECT 478.950 868.950 481.050 871.050 ;
        RECT 521.400 868.050 522.600 883.950 ;
        RECT 530.400 883.050 531.600 884.100 ;
        RECT 536.400 883.050 537.600 884.100 ;
        RECT 542.400 883.050 543.600 889.950 ;
        RECT 556.200 887.100 558.300 889.200 ;
        RECT 560.400 888.900 561.600 891.450 ;
        RECT 544.950 883.950 547.050 886.050 ;
        RECT 526.950 880.950 529.050 883.050 ;
        RECT 529.950 880.950 532.050 883.050 ;
        RECT 532.950 880.950 535.050 883.050 ;
        RECT 535.950 880.950 538.050 883.050 ;
        RECT 541.950 880.950 544.050 883.050 ;
        RECT 520.950 865.950 523.050 868.050 ;
        RECT 469.950 844.950 472.050 847.050 ;
        RECT 484.950 844.950 487.050 847.050 ;
        RECT 502.950 844.950 505.050 847.050 ;
        RECT 514.950 844.950 517.050 847.050 ;
        RECT 466.950 839.100 469.050 841.200 ;
        RECT 454.950 835.950 457.050 838.050 ;
        RECT 457.950 835.950 460.050 838.050 ;
        RECT 460.950 835.950 463.050 838.050 ;
        RECT 463.950 835.950 466.050 838.050 ;
        RECT 455.400 835.050 456.600 835.950 ;
        RECT 451.950 833.400 456.600 835.050 ;
        RECT 461.400 834.000 462.600 835.950 ;
        RECT 470.400 835.050 471.600 844.950 ;
        RECT 478.950 839.100 481.050 841.200 ;
        RECT 479.400 838.050 480.600 839.100 ;
        RECT 485.400 838.050 486.600 844.950 ;
        RECT 493.950 839.100 496.050 841.200 ;
        RECT 478.950 835.950 481.050 838.050 ;
        RECT 481.950 835.950 484.050 838.050 ;
        RECT 484.950 835.950 487.050 838.050 ;
        RECT 487.950 835.950 490.050 838.050 ;
        RECT 451.950 832.950 456.000 833.400 ;
        RECT 448.950 829.950 451.050 832.050 ;
        RECT 460.950 829.950 463.050 834.000 ;
        RECT 469.950 832.950 472.050 835.050 ;
        RECT 482.400 834.900 483.600 835.950 ;
        RECT 481.950 832.800 484.050 834.900 ;
        RECT 488.400 829.050 489.600 835.950 ;
        RECT 463.950 826.950 466.050 829.050 ;
        RECT 487.950 826.950 490.050 829.050 ;
        RECT 445.950 823.950 448.050 826.050 ;
        RECT 454.950 808.950 457.050 811.050 ;
        RECT 445.950 806.100 448.050 808.200 ;
        RECT 446.400 805.050 447.600 806.100 ;
        RECT 439.950 802.950 442.050 805.050 ;
        RECT 442.950 802.950 445.050 805.050 ;
        RECT 445.950 802.950 448.050 805.050 ;
        RECT 448.950 802.950 451.050 805.050 ;
        RECT 443.400 796.050 444.600 802.950 ;
        RECT 449.400 801.900 450.600 802.950 ;
        RECT 455.400 801.900 456.600 808.950 ;
        RECT 464.400 805.050 465.600 826.950 ;
        RECT 494.400 823.050 495.600 839.100 ;
        RECT 503.400 838.050 504.600 844.950 ;
        RECT 508.950 839.100 511.050 841.200 ;
        RECT 509.400 838.050 510.600 839.100 ;
        RECT 499.950 835.950 502.050 838.050 ;
        RECT 502.950 835.950 505.050 838.050 ;
        RECT 505.950 835.950 508.050 838.050 ;
        RECT 508.950 835.950 511.050 838.050 ;
        RECT 500.400 829.050 501.600 835.950 ;
        RECT 506.400 834.000 507.600 835.950 ;
        RECT 515.400 835.050 516.600 844.950 ;
        RECT 505.950 829.950 508.050 834.000 ;
        RECT 511.950 829.950 514.050 835.050 ;
        RECT 514.950 832.950 517.050 835.050 ;
        RECT 521.400 832.050 522.600 865.950 ;
        RECT 527.400 856.050 528.600 880.950 ;
        RECT 533.400 879.900 534.600 880.950 ;
        RECT 532.950 877.800 535.050 879.900 ;
        RECT 545.400 877.050 546.600 883.950 ;
        RECT 554.400 883.200 555.600 885.600 ;
        RECT 553.950 883.050 556.050 883.200 ;
        RECT 551.400 881.100 556.050 883.050 ;
        RECT 556.950 882.000 557.850 887.100 ;
        RECT 559.500 886.800 561.600 888.900 ;
        RECT 563.400 885.900 564.600 892.950 ;
        RECT 601.950 889.950 604.050 892.050 ;
        RECT 613.950 889.950 616.050 892.050 ;
        RECT 640.950 889.950 643.050 892.050 ;
        RECT 667.950 889.950 670.050 892.050 ;
        RECT 566.250 887.400 568.350 889.500 ;
        RECT 563.400 885.000 565.800 885.900 ;
        RECT 558.750 883.800 565.800 885.000 ;
        RECT 558.750 882.900 560.850 883.800 ;
        RECT 563.700 882.000 565.800 882.900 ;
        RECT 556.950 881.100 565.800 882.000 ;
        RECT 551.400 880.950 553.950 881.100 ;
        RECT 544.950 874.950 547.050 877.050 ;
        RECT 551.400 868.050 552.600 880.950 ;
        RECT 556.950 874.500 557.850 881.100 ;
        RECT 563.700 880.800 565.800 881.100 ;
        RECT 559.500 878.100 561.600 880.200 ;
        RECT 556.800 872.400 558.900 874.500 ;
        RECT 550.950 865.950 553.050 868.050 ;
        RECT 560.400 862.050 561.600 878.100 ;
        RECT 566.700 874.800 567.600 887.400 ;
        RECT 574.950 884.100 577.050 886.200 ;
        RECT 580.950 884.100 583.050 886.200 ;
        RECT 586.950 884.100 589.050 886.200 ;
        RECT 568.500 881.100 570.600 883.200 ;
        RECT 569.400 879.900 570.600 881.100 ;
        RECT 568.950 877.800 571.050 879.900 ;
        RECT 575.400 877.050 576.600 884.100 ;
        RECT 581.400 883.050 582.600 884.100 ;
        RECT 587.400 883.050 588.600 884.100 ;
        RECT 592.950 883.950 595.050 889.050 ;
        RECT 595.950 883.950 598.050 886.050 ;
        RECT 580.950 880.950 583.050 883.050 ;
        RECT 583.950 880.950 586.050 883.050 ;
        RECT 586.950 880.950 589.050 883.050 ;
        RECT 589.950 880.950 592.050 883.050 ;
        RECT 584.400 879.900 585.600 880.950 ;
        RECT 590.400 879.900 591.600 880.950 ;
        RECT 583.950 877.800 586.050 879.900 ;
        RECT 589.950 877.800 592.050 879.900 ;
        RECT 592.950 877.950 595.050 880.050 ;
        RECT 596.400 879.900 597.600 883.950 ;
        RECT 574.950 874.950 577.050 877.050 ;
        RECT 565.800 872.700 567.900 874.800 ;
        RECT 575.400 862.050 576.600 874.950 ;
        RECT 559.950 859.950 562.050 862.050 ;
        RECT 574.950 859.950 577.050 862.050 ;
        RECT 526.950 853.950 529.050 856.050 ;
        RECT 560.400 853.050 561.600 859.950 ;
        RECT 544.950 850.950 547.050 853.050 ;
        RECT 559.950 850.950 562.050 853.050 ;
        RECT 541.950 844.950 544.050 847.050 ;
        RECT 542.400 841.200 543.600 844.950 ;
        RECT 529.950 839.100 532.050 841.200 ;
        RECT 535.950 839.100 538.050 841.200 ;
        RECT 541.950 839.100 544.050 841.200 ;
        RECT 530.400 838.050 531.600 839.100 ;
        RECT 536.400 838.050 537.600 839.100 ;
        RECT 526.950 835.950 529.050 838.050 ;
        RECT 529.950 835.950 532.050 838.050 ;
        RECT 532.950 835.950 535.050 838.050 ;
        RECT 535.950 835.950 538.050 838.050 ;
        RECT 527.400 834.900 528.600 835.950 ;
        RECT 526.950 832.800 529.050 834.900 ;
        RECT 520.950 829.950 523.050 832.050 ;
        RECT 533.400 829.050 534.600 835.950 ;
        RECT 538.950 832.950 541.050 835.050 ;
        RECT 499.950 826.950 502.050 829.050 ;
        RECT 532.950 826.950 535.050 829.050 ;
        RECT 535.950 823.950 538.050 826.050 ;
        RECT 493.950 820.950 496.050 823.050 ;
        RECT 514.950 820.950 517.050 823.050 ;
        RECT 478.950 811.950 481.050 814.050 ;
        RECT 469.950 807.000 472.050 811.050 ;
        RECT 470.400 805.050 471.600 807.000 ;
        RECT 463.950 802.950 466.050 805.050 ;
        RECT 466.950 802.950 469.050 805.050 ;
        RECT 469.950 802.950 472.050 805.050 ;
        RECT 472.950 802.950 475.050 805.050 ;
        RECT 448.950 799.800 451.050 801.900 ;
        RECT 454.950 799.800 457.050 801.900 ;
        RECT 442.950 793.950 445.050 796.050 ;
        RECT 467.400 790.050 468.600 802.950 ;
        RECT 473.400 801.900 474.600 802.950 ;
        RECT 479.400 801.900 480.600 811.950 ;
        RECT 490.950 806.100 493.050 808.200 ;
        RECT 491.400 805.050 492.600 806.100 ;
        RECT 515.400 805.050 516.600 820.950 ;
        RECT 536.400 820.050 537.600 823.950 ;
        RECT 539.400 823.050 540.600 832.950 ;
        RECT 542.400 825.600 543.600 839.100 ;
        RECT 545.400 835.050 546.600 850.950 ;
        RECT 553.950 844.950 556.050 847.050 ;
        RECT 554.400 838.050 555.600 844.950 ;
        RECT 577.500 844.500 579.600 846.600 ;
        RECT 559.950 839.100 562.050 841.200 ;
        RECT 560.400 838.050 561.600 839.100 ;
        RECT 550.950 835.950 553.050 838.050 ;
        RECT 553.950 835.950 556.050 838.050 ;
        RECT 556.950 835.950 559.050 838.050 ;
        RECT 559.950 835.950 562.050 838.050 ;
        RECT 544.950 832.950 547.050 835.050 ;
        RECT 551.400 834.900 552.600 835.950 ;
        RECT 550.950 832.800 553.050 834.900 ;
        RECT 557.400 829.050 558.600 835.950 ;
        RECT 562.800 832.950 564.900 835.050 ;
        RECT 565.950 832.950 568.050 838.050 ;
        RECT 574.950 835.950 577.050 838.050 ;
        RECT 577.950 837.300 579.000 844.500 ;
        RECT 581.400 840.900 582.600 843.450 ;
        RECT 587.100 843.300 589.200 845.400 ;
        RECT 580.800 838.800 582.900 840.900 ;
        RECT 583.800 839.700 585.900 841.800 ;
        RECT 583.800 837.300 584.700 839.700 ;
        RECT 577.950 836.100 584.700 837.300 ;
        RECT 575.400 833.400 576.600 835.950 ;
        RECT 556.950 826.950 559.050 829.050 ;
        RECT 542.400 824.400 546.600 825.600 ;
        RECT 538.950 820.950 541.050 823.050 ;
        RECT 545.400 820.050 546.600 824.400 ;
        RECT 563.400 823.050 564.600 832.950 ;
        RECT 565.950 829.800 568.050 831.900 ;
        RECT 577.950 830.700 578.850 836.100 ;
        RECT 579.750 834.300 581.850 835.200 ;
        RECT 587.400 834.300 588.300 843.300 ;
        RECT 590.400 838.050 591.600 840.600 ;
        RECT 593.400 838.050 594.600 877.950 ;
        RECT 595.950 877.800 598.050 879.900 ;
        RECT 596.400 850.050 597.600 877.800 ;
        RECT 602.400 874.050 603.600 889.950 ;
        RECT 607.950 884.100 610.050 886.200 ;
        RECT 608.400 883.050 609.600 884.100 ;
        RECT 614.400 883.050 615.600 889.950 ;
        RECT 622.950 883.950 625.050 886.050 ;
        RECT 634.950 884.100 637.050 886.200 ;
        RECT 607.950 880.950 610.050 883.050 ;
        RECT 610.950 880.950 613.050 883.050 ;
        RECT 613.950 880.950 616.050 883.050 ;
        RECT 616.950 880.950 619.050 883.050 ;
        RECT 611.400 879.000 612.600 880.950 ;
        RECT 617.400 879.900 618.600 880.950 ;
        RECT 610.950 874.950 613.050 879.000 ;
        RECT 616.950 877.800 619.050 879.900 ;
        RECT 623.400 877.050 624.600 883.950 ;
        RECT 635.400 883.050 636.600 884.100 ;
        RECT 641.400 883.050 642.600 889.950 ;
        RECT 649.950 883.950 652.050 886.050 ;
        RECT 655.950 884.100 658.050 886.200 ;
        RECT 661.950 884.100 664.050 886.200 ;
        RECT 668.400 886.050 669.600 889.950 ;
        RECT 670.950 886.950 673.050 889.050 ;
        RECT 631.950 880.950 634.050 883.050 ;
        RECT 634.950 880.950 637.050 883.050 ;
        RECT 637.950 880.950 640.050 883.050 ;
        RECT 640.950 880.950 643.050 883.050 ;
        RECT 622.950 874.950 625.050 877.050 ;
        RECT 601.950 871.950 604.050 874.050 ;
        RECT 595.950 847.950 598.050 850.050 ;
        RECT 596.400 841.200 597.600 847.950 ;
        RECT 595.950 839.100 598.050 841.200 ;
        RECT 602.400 838.050 603.600 871.950 ;
        RECT 632.400 862.050 633.600 880.950 ;
        RECT 634.950 874.950 637.050 877.050 ;
        RECT 635.400 868.050 636.600 874.950 ;
        RECT 638.400 871.050 639.600 880.950 ;
        RECT 650.400 879.900 651.600 883.950 ;
        RECT 656.400 883.050 657.600 884.100 ;
        RECT 662.400 883.050 663.600 884.100 ;
        RECT 667.950 883.950 670.050 886.050 ;
        RECT 655.950 880.950 658.050 883.050 ;
        RECT 658.950 880.950 661.050 883.050 ;
        RECT 661.950 880.950 664.050 883.050 ;
        RECT 664.950 880.950 667.050 883.050 ;
        RECT 649.950 877.800 652.050 879.900 ;
        RECT 659.400 879.000 660.600 880.950 ;
        RECT 665.400 879.900 666.600 880.950 ;
        RECT 671.400 879.900 672.600 886.950 ;
        RECT 680.400 883.050 681.600 892.950 ;
        RECT 676.950 880.950 679.050 883.050 ;
        RECT 679.950 880.950 682.050 883.050 ;
        RECT 682.950 880.950 685.050 883.050 ;
        RECT 677.400 879.900 678.600 880.950 ;
        RECT 683.400 879.900 684.600 880.950 ;
        RECT 637.950 868.950 640.050 871.050 ;
        RECT 634.950 865.950 637.050 868.050 ;
        RECT 631.950 859.950 634.050 862.050 ;
        RECT 616.950 853.950 619.050 856.050 ;
        RECT 607.950 850.950 610.050 853.050 ;
        RECT 608.400 838.050 609.600 850.950 ;
        RECT 589.500 835.950 591.600 838.050 ;
        RECT 592.950 835.950 595.050 838.050 ;
        RECT 601.950 835.950 604.050 838.050 ;
        RECT 604.950 835.950 607.050 838.050 ;
        RECT 607.950 835.950 610.050 838.050 ;
        RECT 610.950 835.950 613.050 838.050 ;
        RECT 579.750 833.100 588.300 834.300 ;
        RECT 605.400 834.000 606.600 835.950 ;
        RECT 580.800 832.050 582.900 832.200 ;
        RECT 566.400 826.050 567.600 829.800 ;
        RECT 577.500 828.600 579.600 830.700 ;
        RECT 580.800 830.100 583.050 832.050 ;
        RECT 584.700 831.300 586.800 833.100 ;
        RECT 580.950 829.950 583.050 830.100 ;
        RECT 604.950 829.950 607.050 834.000 ;
        RECT 581.400 827.550 582.600 829.950 ;
        RECT 611.400 826.050 612.600 835.950 ;
        RECT 617.400 832.050 618.600 853.950 ;
        RECT 628.950 839.100 631.050 841.200 ;
        RECT 634.950 840.000 637.050 844.050 ;
        RECT 640.950 841.950 643.050 844.050 ;
        RECT 629.400 838.050 630.600 839.100 ;
        RECT 635.400 838.050 636.600 840.000 ;
        RECT 625.950 835.950 628.050 838.050 ;
        RECT 628.950 835.950 631.050 838.050 ;
        RECT 631.950 835.950 634.050 838.050 ;
        RECT 634.950 835.950 637.050 838.050 ;
        RECT 626.400 835.050 627.600 835.950 ;
        RECT 622.950 832.950 627.600 835.050 ;
        RECT 616.950 829.950 619.050 832.050 ;
        RECT 626.400 826.050 627.600 832.950 ;
        RECT 628.950 826.950 631.050 829.050 ;
        RECT 565.950 823.950 568.050 826.050 ;
        RECT 571.950 823.950 574.050 826.050 ;
        RECT 610.950 823.950 613.050 826.050 ;
        RECT 625.950 823.950 628.050 826.050 ;
        RECT 562.950 820.950 565.050 823.050 ;
        RECT 535.950 817.950 538.050 820.050 ;
        RECT 544.950 817.950 547.050 820.050 ;
        RECT 553.950 814.950 556.050 817.050 ;
        RECT 526.950 811.950 529.050 814.050 ;
        RECT 538.950 811.950 541.050 814.050 ;
        RECT 527.400 808.050 528.600 811.950 ;
        RECT 526.950 805.950 529.050 808.050 ;
        RECT 539.400 805.050 540.600 811.950 ;
        RECT 554.400 808.200 555.600 814.950 ;
        RECT 553.950 806.100 556.050 808.200 ;
        RECT 560.400 806.400 567.600 807.600 ;
        RECT 554.400 805.050 555.600 806.100 ;
        RECT 560.400 805.050 561.600 806.400 ;
        RECT 487.950 802.950 490.050 805.050 ;
        RECT 490.950 802.950 493.050 805.050 ;
        RECT 496.950 802.950 499.050 805.050 ;
        RECT 511.950 802.950 514.050 805.050 ;
        RECT 514.950 802.950 517.050 805.050 ;
        RECT 517.950 802.950 520.050 805.050 ;
        RECT 535.950 802.950 538.050 805.050 ;
        RECT 538.950 802.950 541.050 805.050 ;
        RECT 550.950 802.950 553.050 805.050 ;
        RECT 553.950 802.950 556.050 805.050 ;
        RECT 556.950 802.950 559.050 805.050 ;
        RECT 559.950 802.950 562.050 805.050 ;
        RECT 472.950 799.800 475.050 801.900 ;
        RECT 478.950 799.800 481.050 801.900 ;
        RECT 479.400 796.050 480.600 799.800 ;
        RECT 478.950 793.950 481.050 796.050 ;
        RECT 488.400 790.050 489.600 802.950 ;
        RECT 433.950 787.950 436.050 790.050 ;
        RECT 466.950 787.950 469.050 790.050 ;
        RECT 487.950 787.950 490.050 790.050 ;
        RECT 497.400 787.050 498.600 802.950 ;
        RECT 512.400 787.050 513.600 802.950 ;
        RECT 518.400 801.900 519.600 802.950 ;
        RECT 536.400 801.900 537.600 802.950 ;
        RECT 517.950 799.800 520.050 801.900 ;
        RECT 535.950 799.800 538.050 801.900 ;
        RECT 518.400 795.600 519.600 799.800 ;
        RECT 518.400 794.400 522.600 795.600 ;
        RECT 496.950 784.950 499.050 787.050 ;
        RECT 511.950 784.950 514.050 787.050 ;
        RECT 460.950 775.950 463.050 778.050 ;
        RECT 472.950 775.950 475.050 778.050 ;
        RECT 428.400 761.400 432.600 762.600 ;
        RECT 410.400 760.050 411.600 760.950 ;
        RECT 409.950 757.950 412.050 760.050 ;
        RECT 412.950 757.950 415.050 760.050 ;
        RECT 397.950 754.800 400.050 756.900 ;
        RECT 403.950 754.950 406.050 757.050 ;
        RECT 406.950 754.950 409.050 757.050 ;
        RECT 413.400 756.900 414.600 757.950 ;
        RECT 388.950 733.950 391.050 736.050 ;
        RECT 385.950 728.100 388.050 730.200 ;
        RECT 391.950 728.100 394.050 730.200 ;
        RECT 397.950 728.100 400.050 730.200 ;
        RECT 386.400 718.050 387.600 728.100 ;
        RECT 392.400 727.050 393.600 728.100 ;
        RECT 398.400 727.050 399.600 728.100 ;
        RECT 391.950 724.950 394.050 727.050 ;
        RECT 394.950 724.950 397.050 727.050 ;
        RECT 397.950 724.950 400.050 727.050 ;
        RECT 395.400 720.600 396.600 724.950 ;
        RECT 392.400 719.400 396.600 720.600 ;
        RECT 385.950 715.950 388.050 718.050 ;
        RECT 382.950 712.950 385.050 715.050 ;
        RECT 392.400 712.050 393.600 719.400 ;
        RECT 394.950 715.950 397.050 718.050 ;
        RECT 370.950 709.950 373.050 712.050 ;
        RECT 391.950 709.950 394.050 712.050 ;
        RECT 373.950 694.950 376.050 697.050 ;
        RECT 388.950 694.950 391.050 697.050 ;
        RECT 361.950 691.950 364.050 694.050 ;
        RECT 359.400 689.400 363.600 690.600 ;
        RECT 340.950 683.100 343.050 685.200 ;
        RECT 341.400 682.050 342.600 683.100 ;
        RECT 349.950 682.950 352.050 685.050 ;
        RECT 355.950 683.100 358.050 685.200 ;
        RECT 331.950 679.950 334.050 682.050 ;
        RECT 334.950 679.950 337.050 682.050 ;
        RECT 340.950 679.950 343.050 682.050 ;
        RECT 346.950 679.950 349.050 682.050 ;
        RECT 335.400 678.900 336.600 679.950 ;
        RECT 334.950 676.800 337.050 678.900 ;
        RECT 347.400 670.050 348.600 679.950 ;
        RECT 346.950 667.950 349.050 670.050 ;
        RECT 328.950 664.950 331.050 667.050 ;
        RECT 325.950 661.950 328.050 664.050 ;
        RECT 307.950 655.950 310.050 661.050 ;
        RECT 313.950 658.950 316.050 661.050 ;
        RECT 310.950 655.950 313.050 658.050 ;
        RECT 316.950 655.950 322.050 658.050 ;
        RECT 295.950 646.950 298.050 649.050 ;
        RECT 298.950 646.950 301.050 649.050 ;
        RECT 301.950 646.950 304.050 649.050 ;
        RECT 304.950 646.950 307.050 649.050 ;
        RECT 296.400 645.900 297.600 646.950 ;
        RECT 295.950 643.800 298.050 645.900 ;
        RECT 302.400 637.050 303.600 646.950 ;
        RECT 307.950 643.950 310.050 646.050 ;
        RECT 301.950 634.950 304.050 637.050 ;
        RECT 295.950 631.950 298.050 634.050 ;
        RECT 289.950 613.950 292.050 616.050 ;
        RECT 266.100 610.200 268.200 612.300 ;
        RECT 275.100 610.500 277.200 612.600 ;
        RECT 235.950 607.950 238.050 610.050 ;
        RECT 236.400 605.400 243.600 606.600 ;
        RECT 247.950 606.000 250.050 610.050 ;
        RECT 236.400 589.050 237.600 605.400 ;
        RECT 242.400 604.050 243.600 605.400 ;
        RECT 248.400 604.050 249.600 606.000 ;
        RECT 241.950 601.950 244.050 604.050 ;
        RECT 244.950 601.950 247.050 604.050 ;
        RECT 247.950 601.950 250.050 604.050 ;
        RECT 250.950 601.950 253.050 604.050 ;
        RECT 263.400 603.900 264.600 606.450 ;
        RECT 245.400 600.900 246.600 601.950 ;
        RECT 244.950 598.800 247.050 600.900 ;
        RECT 251.400 600.000 252.600 601.950 ;
        RECT 263.400 601.800 265.500 603.900 ;
        RECT 250.950 595.950 253.050 600.000 ;
        RECT 256.950 595.950 259.050 598.050 ;
        RECT 266.400 597.600 267.300 610.200 ;
        RECT 272.400 606.900 273.600 609.450 ;
        RECT 272.400 604.800 274.500 606.900 ;
        RECT 268.200 603.900 270.300 604.200 ;
        RECT 276.150 603.900 277.050 610.500 ;
        RECT 286.950 604.950 289.050 607.050 ;
        RECT 268.200 603.000 277.050 603.900 ;
        RECT 268.200 602.100 270.300 603.000 ;
        RECT 273.150 601.200 275.250 602.100 ;
        RECT 268.200 600.000 275.250 601.200 ;
        RECT 268.200 599.100 270.600 600.000 ;
        RECT 238.950 592.950 241.050 595.050 ;
        RECT 235.950 586.950 238.050 589.050 ;
        RECT 233.400 572.400 237.600 573.600 ;
        RECT 229.950 568.950 232.050 571.050 ;
        RECT 230.400 562.050 231.600 568.950 ;
        RECT 236.400 565.050 237.600 572.400 ;
        RECT 239.400 568.050 240.600 592.950 ;
        RECT 247.950 586.950 250.050 589.050 ;
        RECT 248.400 571.050 249.600 586.950 ;
        RECT 244.950 568.950 247.050 571.050 ;
        RECT 247.950 568.950 250.050 571.050 ;
        RECT 250.950 568.950 253.050 571.050 ;
        RECT 238.950 565.950 241.050 568.050 ;
        RECT 245.400 567.900 246.600 568.950 ;
        RECT 244.950 565.800 247.050 567.900 ;
        RECT 235.950 562.950 238.050 565.050 ;
        RECT 229.950 559.950 232.050 562.050 ;
        RECT 226.950 556.500 229.050 558.600 ;
        RECT 236.400 541.050 237.600 562.950 ;
        RECT 241.950 553.950 244.050 556.050 ;
        RECT 235.950 538.950 238.050 541.050 ;
        RECT 223.950 532.950 226.050 535.050 ;
        RECT 220.950 529.950 223.050 532.050 ;
        RECT 224.400 526.050 225.600 532.950 ;
        RECT 229.950 528.000 232.050 532.050 ;
        RECT 235.950 529.950 238.050 532.050 ;
        RECT 230.400 526.050 231.600 528.000 ;
        RECT 220.950 523.950 223.050 526.050 ;
        RECT 223.950 523.950 226.050 526.050 ;
        RECT 226.950 523.950 229.050 526.050 ;
        RECT 229.950 523.950 232.050 526.050 ;
        RECT 221.400 517.050 222.600 523.950 ;
        RECT 227.400 522.900 228.600 523.950 ;
        RECT 226.950 520.800 229.050 522.900 ;
        RECT 220.950 514.950 223.050 517.050 ;
        RECT 229.950 511.950 232.050 514.050 ;
        RECT 217.950 502.950 220.050 505.050 ;
        RECT 226.950 502.950 229.050 505.050 ;
        RECT 208.950 499.950 211.050 502.050 ;
        RECT 214.950 499.950 217.050 502.050 ;
        RECT 205.950 496.950 208.050 499.050 ;
        RECT 202.950 484.950 205.050 487.050 ;
        RECT 206.400 478.050 207.600 496.950 ;
        RECT 209.400 489.900 210.600 499.950 ;
        RECT 211.950 493.950 214.050 499.050 ;
        RECT 218.400 493.050 219.600 502.950 ;
        RECT 227.400 496.050 228.600 502.950 ;
        RECT 226.950 493.950 229.050 496.050 ;
        RECT 214.950 490.950 217.050 493.050 ;
        RECT 217.950 490.950 220.050 493.050 ;
        RECT 223.950 490.950 226.050 493.050 ;
        RECT 208.950 487.800 211.050 489.900 ;
        RECT 215.400 484.050 216.600 490.950 ;
        RECT 224.400 489.900 225.600 490.950 ;
        RECT 223.800 487.800 225.900 489.900 ;
        RECT 226.950 487.800 229.050 489.900 ;
        RECT 214.950 481.950 217.050 484.050 ;
        RECT 196.950 475.950 199.050 478.050 ;
        RECT 205.950 475.950 208.050 478.050 ;
        RECT 197.400 472.050 198.600 475.950 ;
        RECT 196.950 469.950 199.050 472.050 ;
        RECT 208.950 457.950 211.050 460.050 ;
        RECT 220.950 457.950 223.050 460.050 ;
        RECT 199.950 454.950 202.050 457.050 ;
        RECT 193.950 449.100 196.050 451.200 ;
        RECT 194.400 448.050 195.600 449.100 ;
        RECT 200.400 448.050 201.600 454.950 ;
        RECT 193.950 445.950 196.050 448.050 ;
        RECT 196.950 445.950 199.050 448.050 ;
        RECT 199.950 445.950 202.050 448.050 ;
        RECT 202.950 445.950 205.050 448.050 ;
        RECT 187.950 436.950 190.050 439.050 ;
        RECT 184.950 433.950 187.050 436.050 ;
        RECT 181.950 430.950 184.050 433.050 ;
        RECT 182.400 415.050 183.600 430.950 ;
        RECT 197.400 424.050 198.600 445.950 ;
        RECT 203.400 444.900 204.600 445.950 ;
        RECT 202.950 442.800 205.050 444.900 ;
        RECT 209.400 430.050 210.600 457.950 ;
        RECT 214.950 449.100 217.050 454.050 ;
        RECT 215.400 448.050 216.600 449.100 ;
        RECT 221.400 448.050 222.600 457.950 ;
        RECT 227.400 451.050 228.600 487.800 ;
        RECT 230.400 466.050 231.600 511.950 ;
        RECT 236.400 511.050 237.600 529.950 ;
        RECT 238.950 526.950 241.050 529.050 ;
        RECT 239.400 517.050 240.600 526.950 ;
        RECT 242.400 520.050 243.600 553.950 ;
        RECT 251.400 550.050 252.600 568.950 ;
        RECT 250.950 547.950 253.050 550.050 ;
        RECT 257.400 549.600 258.600 595.950 ;
        RECT 265.650 595.500 267.750 597.600 ;
        RECT 269.400 595.050 270.600 599.100 ;
        RECT 272.400 596.100 274.500 598.200 ;
        RECT 276.150 597.900 277.050 603.000 ;
        RECT 277.950 601.800 280.050 603.900 ;
        RECT 278.400 599.400 279.600 601.800 ;
        RECT 268.950 592.950 271.050 595.050 ;
        RECT 268.950 583.950 271.050 586.050 ;
        RECT 269.400 571.050 270.600 583.950 ;
        RECT 272.400 577.050 273.600 596.100 ;
        RECT 275.700 595.800 277.800 597.900 ;
        RECT 287.400 589.050 288.600 604.950 ;
        RECT 296.400 604.050 297.600 631.950 ;
        RECT 292.950 601.950 295.050 604.050 ;
        RECT 295.950 601.950 298.050 604.050 ;
        RECT 298.950 601.950 301.050 604.050 ;
        RECT 293.400 595.050 294.600 601.950 ;
        RECT 292.950 592.950 295.050 595.050 ;
        RECT 299.400 589.050 300.600 601.950 ;
        RECT 308.400 589.050 309.600 643.950 ;
        RECT 311.400 637.050 312.600 655.950 ;
        RECT 316.950 650.100 319.050 652.200 ;
        RECT 322.950 650.100 325.050 652.200 ;
        RECT 317.400 649.050 318.600 650.100 ;
        RECT 323.400 649.050 324.600 650.100 ;
        RECT 316.950 646.950 319.050 649.050 ;
        RECT 319.950 646.950 322.050 649.050 ;
        RECT 322.950 646.950 325.050 649.050 ;
        RECT 320.400 637.050 321.600 646.950 ;
        RECT 310.950 634.950 313.050 637.050 ;
        RECT 319.950 634.950 322.050 637.050 ;
        RECT 329.400 634.050 330.600 664.950 ;
        RECT 340.950 658.950 343.050 661.050 ;
        RECT 341.400 649.050 342.600 658.950 ;
        RECT 337.950 646.950 340.050 649.050 ;
        RECT 340.950 646.950 343.050 649.050 ;
        RECT 343.950 646.950 346.050 649.050 ;
        RECT 328.950 631.950 331.050 634.050 ;
        RECT 316.950 605.100 319.050 607.200 ;
        RECT 322.950 606.000 325.050 610.050 ;
        RECT 317.400 604.050 318.600 605.100 ;
        RECT 323.400 604.050 324.600 606.000 ;
        RECT 338.400 604.050 339.600 646.950 ;
        RECT 344.400 645.000 345.600 646.950 ;
        RECT 343.950 640.950 346.050 645.000 ;
        RECT 350.400 625.050 351.600 682.950 ;
        RECT 356.400 682.050 357.600 683.100 ;
        RECT 362.400 682.050 363.600 689.400 ;
        RECT 374.400 688.050 375.600 694.950 ;
        RECT 376.950 688.950 379.050 691.050 ;
        RECT 382.950 688.950 385.050 691.050 ;
        RECT 367.950 684.000 370.050 688.050 ;
        RECT 373.950 685.950 376.050 688.050 ;
        RECT 368.400 682.050 369.600 684.000 ;
        RECT 355.950 679.950 358.050 682.050 ;
        RECT 358.950 679.950 361.050 682.050 ;
        RECT 361.950 679.950 364.050 682.050 ;
        RECT 364.950 679.950 367.050 682.050 ;
        RECT 367.950 679.950 370.050 682.050 ;
        RECT 359.400 678.900 360.600 679.950 ;
        RECT 358.950 676.800 361.050 678.900 ;
        RECT 358.950 670.950 361.050 673.050 ;
        RECT 352.950 667.950 355.050 670.050 ;
        RECT 355.950 667.950 358.050 670.050 ;
        RECT 353.400 646.050 354.600 667.950 ;
        RECT 352.950 643.950 355.050 646.050 ;
        RECT 356.400 628.050 357.600 667.950 ;
        RECT 359.400 652.200 360.600 670.950 ;
        RECT 365.400 670.050 366.600 679.950 ;
        RECT 364.950 667.950 367.050 670.050 ;
        RECT 374.400 660.600 375.600 685.950 ;
        RECT 377.400 678.900 378.600 688.950 ;
        RECT 383.400 682.050 384.600 688.950 ;
        RECT 389.400 682.050 390.600 694.950 ;
        RECT 382.950 679.950 385.050 682.050 ;
        RECT 385.950 679.950 388.050 682.050 ;
        RECT 388.950 679.950 391.050 682.050 ;
        RECT 386.400 678.900 387.600 679.950 ;
        RECT 376.950 676.800 379.050 678.900 ;
        RECT 385.950 676.800 388.050 678.900 ;
        RECT 395.400 673.050 396.600 715.950 ;
        RECT 397.950 697.950 400.050 700.050 ;
        RECT 398.400 679.050 399.600 697.950 ;
        RECT 407.400 697.050 408.600 754.950 ;
        RECT 412.950 754.800 415.050 756.900 ;
        RECT 415.950 745.950 418.050 748.050 ;
        RECT 416.400 730.200 417.600 745.950 ;
        RECT 415.950 728.100 418.050 730.200 ;
        RECT 416.400 727.050 417.600 728.100 ;
        RECT 412.950 724.950 415.050 727.050 ;
        RECT 415.950 724.950 418.050 727.050 ;
        RECT 418.950 724.950 421.050 727.050 ;
        RECT 413.400 700.050 414.600 724.950 ;
        RECT 419.400 723.600 420.600 724.950 ;
        RECT 419.400 722.400 423.600 723.600 ;
        RECT 418.950 712.950 421.050 715.050 ;
        RECT 412.950 697.950 415.050 700.050 ;
        RECT 406.950 694.950 409.050 697.050 ;
        RECT 415.950 694.950 418.050 697.050 ;
        RECT 416.400 691.050 417.600 694.950 ;
        RECT 415.950 688.950 418.050 691.050 ;
        RECT 403.950 683.100 406.050 685.200 ;
        RECT 409.950 683.100 412.050 685.200 ;
        RECT 416.400 685.050 417.600 688.950 ;
        RECT 404.400 682.050 405.600 683.100 ;
        RECT 410.400 682.050 411.600 683.100 ;
        RECT 415.950 682.950 418.050 685.050 ;
        RECT 403.950 679.950 406.050 682.050 ;
        RECT 406.950 679.950 409.050 682.050 ;
        RECT 409.950 679.950 412.050 682.050 ;
        RECT 412.950 679.950 415.050 682.050 ;
        RECT 397.950 676.950 400.050 679.050 ;
        RECT 407.400 678.900 408.600 679.950 ;
        RECT 406.950 676.800 409.050 678.900 ;
        RECT 413.400 673.050 414.600 679.950 ;
        RECT 415.950 676.950 418.050 679.050 ;
        RECT 394.950 670.950 397.050 673.050 ;
        RECT 409.800 670.950 411.900 673.050 ;
        RECT 412.950 670.950 415.050 673.050 ;
        RECT 385.950 667.950 388.050 670.050 ;
        RECT 379.950 664.950 382.050 667.050 ;
        RECT 374.400 659.400 378.600 660.600 ;
        RECT 358.950 650.100 361.050 652.200 ;
        RECT 367.950 651.600 370.050 655.050 ;
        RECT 365.400 651.000 370.050 651.600 ;
        RECT 365.400 650.400 369.600 651.000 ;
        RECT 365.400 649.050 366.600 650.400 ;
        RECT 361.950 646.950 364.050 649.050 ;
        RECT 364.950 646.950 367.050 649.050 ;
        RECT 370.950 646.950 373.050 649.050 ;
        RECT 362.400 645.900 363.600 646.950 ;
        RECT 361.950 643.800 364.050 645.900 ;
        RECT 371.400 640.050 372.600 646.950 ;
        RECT 377.400 640.050 378.600 659.400 ;
        RECT 370.950 637.950 373.050 640.050 ;
        RECT 376.950 637.950 379.050 640.050 ;
        RECT 355.950 625.950 358.050 628.050 ;
        RECT 349.950 622.950 352.050 625.050 ;
        RECT 370.950 622.950 373.050 625.050 ;
        RECT 358.950 613.950 361.050 616.050 ;
        RECT 346.950 606.000 349.050 610.050 ;
        RECT 359.400 607.200 360.600 613.950 ;
        RECT 347.400 604.050 348.600 606.000 ;
        RECT 358.950 605.100 361.050 607.200 ;
        RECT 364.950 606.000 367.050 610.050 ;
        RECT 359.400 604.050 360.600 605.100 ;
        RECT 365.400 604.050 366.600 606.000 ;
        RECT 316.950 601.950 319.050 604.050 ;
        RECT 319.950 601.950 322.050 604.050 ;
        RECT 322.950 601.950 325.050 604.050 ;
        RECT 337.950 601.950 340.050 604.050 ;
        RECT 340.950 601.950 343.050 604.050 ;
        RECT 346.950 601.950 349.050 604.050 ;
        RECT 358.950 601.950 361.050 604.050 ;
        RECT 361.950 601.950 364.050 604.050 ;
        RECT 364.950 601.950 367.050 604.050 ;
        RECT 320.400 589.050 321.600 601.950 ;
        RECT 325.950 598.950 328.050 601.050 ;
        RECT 322.950 592.950 325.050 598.050 ;
        RECT 326.400 591.600 327.600 598.950 ;
        RECT 328.950 595.950 334.050 598.050 ;
        RECT 341.400 592.050 342.600 601.950 ;
        RECT 358.950 595.950 361.050 598.050 ;
        RECT 328.950 591.600 331.050 592.050 ;
        RECT 326.400 590.400 331.050 591.600 ;
        RECT 328.950 589.950 331.050 590.400 ;
        RECT 340.950 589.950 343.050 592.050 ;
        RECT 286.950 586.950 289.050 589.050 ;
        RECT 298.950 586.950 301.050 589.050 ;
        RECT 307.950 586.950 310.050 589.050 ;
        RECT 319.950 586.950 322.050 589.050 ;
        RECT 271.950 574.950 274.050 577.050 ;
        RECT 277.950 574.950 280.050 577.050 ;
        RECT 265.950 568.950 268.050 571.050 ;
        RECT 268.950 568.950 271.050 571.050 ;
        RECT 271.950 568.950 274.050 571.050 ;
        RECT 266.400 567.000 267.600 568.950 ;
        RECT 272.400 567.900 273.600 568.950 ;
        RECT 265.950 562.950 268.050 567.000 ;
        RECT 271.950 565.800 274.050 567.900 ;
        RECT 259.950 549.600 262.050 550.050 ;
        RECT 257.400 548.400 262.050 549.600 ;
        RECT 259.950 547.950 262.050 548.400 ;
        RECT 253.950 527.100 256.050 529.200 ;
        RECT 254.400 526.050 255.600 527.100 ;
        RECT 247.950 523.950 250.050 526.050 ;
        RECT 253.950 523.950 256.050 526.050 ;
        RECT 248.400 523.050 249.600 523.950 ;
        RECT 248.400 522.000 253.050 523.050 ;
        RECT 247.950 520.950 253.050 522.000 ;
        RECT 241.950 517.950 244.050 520.050 ;
        RECT 247.950 517.950 250.050 520.950 ;
        RECT 238.950 514.950 241.050 517.050 ;
        RECT 250.950 514.950 253.050 517.050 ;
        RECT 235.950 508.950 238.050 511.050 ;
        RECT 239.400 502.050 240.600 514.950 ;
        RECT 251.400 505.050 252.600 514.950 ;
        RECT 253.950 511.950 256.050 514.050 ;
        RECT 250.950 502.950 253.050 505.050 ;
        RECT 238.950 499.950 241.050 502.050 ;
        RECT 247.800 499.950 249.900 502.050 ;
        RECT 238.950 494.100 241.050 496.200 ;
        RECT 239.400 493.050 240.600 494.100 ;
        RECT 235.950 490.950 238.050 493.050 ;
        RECT 238.950 490.950 241.050 493.050 ;
        RECT 241.950 490.950 244.050 493.050 ;
        RECT 236.400 489.900 237.600 490.950 ;
        RECT 235.950 487.800 238.050 489.900 ;
        RECT 242.400 478.050 243.600 490.950 ;
        RECT 244.950 487.950 247.050 490.050 ;
        RECT 241.950 475.950 244.050 478.050 ;
        RECT 229.950 463.950 232.050 466.050 ;
        RECT 238.950 463.950 241.050 466.050 ;
        RECT 232.950 459.300 235.050 461.400 ;
        RECT 233.850 455.700 235.050 459.300 ;
        RECT 232.950 453.600 235.050 455.700 ;
        RECT 226.950 448.950 229.050 451.050 ;
        RECT 214.950 445.950 217.050 448.050 ;
        RECT 217.950 445.950 220.050 448.050 ;
        RECT 220.950 445.950 223.050 448.050 ;
        RECT 229.950 445.950 232.050 448.050 ;
        RECT 218.400 439.050 219.600 445.950 ;
        RECT 226.950 444.600 229.050 445.050 ;
        RECT 230.400 444.600 231.600 445.950 ;
        RECT 226.950 443.400 231.600 444.600 ;
        RECT 226.950 442.950 229.050 443.400 ;
        RECT 217.950 436.950 220.050 439.050 ;
        RECT 208.950 427.950 211.050 430.050 ;
        RECT 196.950 421.950 199.050 424.050 ;
        RECT 227.400 418.200 228.600 442.950 ;
        RECT 233.850 438.600 235.050 453.600 ;
        RECT 239.400 445.050 240.600 463.950 ;
        RECT 241.950 451.950 244.050 454.050 ;
        RECT 238.950 442.950 241.050 445.050 ;
        RECT 232.950 436.500 235.050 438.600 ;
        RECT 235.950 427.950 238.050 430.050 ;
        RECT 188.400 416.400 195.600 417.600 ;
        RECT 188.400 415.050 189.600 416.400 ;
        RECT 178.950 412.950 181.050 415.050 ;
        RECT 181.950 412.950 184.050 415.050 ;
        RECT 184.950 412.950 187.050 415.050 ;
        RECT 187.950 412.950 190.050 415.050 ;
        RECT 179.400 411.900 180.600 412.950 ;
        RECT 185.400 411.900 186.600 412.950 ;
        RECT 178.950 409.800 181.050 411.900 ;
        RECT 184.950 409.800 187.050 411.900 ;
        RECT 194.400 406.050 195.600 416.400 ;
        RECT 196.950 416.100 199.050 418.200 ;
        RECT 202.950 416.100 205.050 418.200 ;
        RECT 208.950 416.100 211.050 418.200 ;
        RECT 197.400 412.050 198.600 416.100 ;
        RECT 203.400 415.050 204.600 416.100 ;
        RECT 209.400 415.050 210.600 416.100 ;
        RECT 214.800 415.950 216.900 418.050 ;
        RECT 217.950 415.950 220.050 418.050 ;
        RECT 226.950 416.100 229.050 418.200 ;
        RECT 232.950 416.100 235.050 418.200 ;
        RECT 202.950 412.950 205.050 415.050 ;
        RECT 205.950 412.950 208.050 415.050 ;
        RECT 208.950 412.950 211.050 415.050 ;
        RECT 196.950 409.950 199.050 412.050 ;
        RECT 193.950 403.950 196.050 406.050 ;
        RECT 190.950 394.950 193.050 397.050 ;
        RECT 187.950 391.950 190.050 394.050 ;
        RECT 172.950 379.950 175.050 382.050 ;
        RECT 172.950 371.100 175.050 373.200 ;
        RECT 178.950 371.100 181.050 373.200 ;
        RECT 173.400 370.050 174.600 371.100 ;
        RECT 179.400 370.050 180.600 371.100 ;
        RECT 184.950 370.950 187.050 373.050 ;
        RECT 169.950 367.950 172.050 370.050 ;
        RECT 172.950 367.950 175.050 370.050 ;
        RECT 175.950 367.950 178.050 370.050 ;
        RECT 178.950 367.950 181.050 370.050 ;
        RECT 170.400 358.050 171.600 367.950 ;
        RECT 169.950 355.950 172.050 358.050 ;
        RECT 176.400 343.050 177.600 367.950 ;
        RECT 181.950 364.950 184.050 367.050 ;
        RECT 182.400 352.050 183.600 364.950 ;
        RECT 185.400 364.050 186.600 370.950 ;
        RECT 184.950 361.950 187.050 364.050 ;
        RECT 188.400 358.050 189.600 391.950 ;
        RECT 191.400 367.050 192.600 394.950 ;
        RECT 206.400 394.050 207.600 412.950 ;
        RECT 215.400 406.050 216.600 415.950 ;
        RECT 214.950 403.950 217.050 406.050 ;
        RECT 205.950 391.950 208.050 394.050 ;
        RECT 211.950 381.300 214.050 383.400 ;
        RECT 212.850 377.700 214.050 381.300 ;
        RECT 211.950 375.600 214.050 377.700 ;
        RECT 199.950 371.100 202.050 373.200 ;
        RECT 200.400 370.050 201.600 371.100 ;
        RECT 196.950 367.950 199.050 370.050 ;
        RECT 199.950 367.950 202.050 370.050 ;
        RECT 202.950 367.950 205.050 370.050 ;
        RECT 208.950 367.950 211.050 370.050 ;
        RECT 190.950 364.950 193.050 367.050 ;
        RECT 197.400 361.050 198.600 367.950 ;
        RECT 203.400 366.000 204.600 367.950 ;
        RECT 202.950 361.950 205.050 366.000 ;
        RECT 205.950 364.950 208.050 367.050 ;
        RECT 209.400 366.000 210.600 367.950 ;
        RECT 196.950 358.950 199.050 361.050 ;
        RECT 187.950 355.950 190.050 358.050 ;
        RECT 181.950 349.950 184.050 352.050 ;
        RECT 196.950 349.950 199.050 352.050 ;
        RECT 187.950 343.950 190.050 346.050 ;
        RECT 175.950 340.950 178.050 343.050 ;
        RECT 181.950 340.950 184.050 343.050 ;
        RECT 163.950 337.950 166.050 340.050 ;
        RECT 172.950 338.100 175.050 340.200 ;
        RECT 164.400 331.050 165.600 337.950 ;
        RECT 173.400 337.050 174.600 338.100 ;
        RECT 169.950 334.950 172.050 337.050 ;
        RECT 172.950 334.950 175.050 337.050 ;
        RECT 175.950 334.950 178.050 337.050 ;
        RECT 170.400 333.000 171.600 334.950 ;
        RECT 160.950 328.950 163.050 331.050 ;
        RECT 163.950 328.950 166.050 331.050 ;
        RECT 169.950 328.950 172.050 333.000 ;
        RECT 176.400 328.050 177.600 334.950 ;
        RECT 175.950 325.950 178.050 328.050 ;
        RECT 182.400 322.050 183.600 340.950 ;
        RECT 188.400 337.050 189.600 343.950 ;
        RECT 187.950 334.950 190.050 337.050 ;
        RECT 190.950 334.950 193.050 337.050 ;
        RECT 154.950 319.950 157.050 322.050 ;
        RECT 181.950 319.950 184.050 322.050 ;
        RECT 191.400 310.050 192.600 334.950 ;
        RECT 197.400 310.050 198.600 349.950 ;
        RECT 199.950 343.950 202.050 346.050 ;
        RECT 200.400 328.050 201.600 343.950 ;
        RECT 206.400 337.050 207.600 364.950 ;
        RECT 208.950 361.950 211.050 366.000 ;
        RECT 212.850 360.600 214.050 375.600 ;
        RECT 218.400 361.050 219.600 415.950 ;
        RECT 227.400 415.050 228.600 416.100 ;
        RECT 223.950 412.950 226.050 415.050 ;
        RECT 226.950 412.950 229.050 415.050 ;
        RECT 224.400 411.900 225.600 412.950 ;
        RECT 223.950 409.800 226.050 411.900 ;
        RECT 233.400 400.050 234.600 416.100 ;
        RECT 236.400 411.600 237.600 427.950 ;
        RECT 242.400 427.050 243.600 451.950 ;
        RECT 245.400 450.600 246.600 487.950 ;
        RECT 248.400 454.050 249.600 499.950 ;
        RECT 250.950 499.800 253.050 501.900 ;
        RECT 251.400 490.050 252.600 499.800 ;
        RECT 250.950 487.950 253.050 490.050 ;
        RECT 254.400 478.050 255.600 511.950 ;
        RECT 260.400 499.050 261.600 547.950 ;
        RECT 278.400 538.050 279.600 574.950 ;
        RECT 329.400 571.050 330.600 589.950 ;
        RECT 334.950 572.100 337.050 574.200 ;
        RECT 335.400 571.050 336.600 572.100 ;
        RECT 340.950 571.950 343.050 574.050 ;
        RECT 310.950 568.950 313.050 571.050 ;
        RECT 325.950 568.950 328.050 571.050 ;
        RECT 328.950 568.950 331.050 571.050 ;
        RECT 331.950 568.950 334.050 571.050 ;
        RECT 334.950 568.950 337.050 571.050 ;
        RECT 298.950 565.800 301.050 567.900 ;
        RECT 280.950 538.950 283.050 541.050 ;
        RECT 262.950 535.950 265.050 538.050 ;
        RECT 277.950 535.950 280.050 538.050 ;
        RECT 263.400 514.050 264.600 535.950 ;
        RECT 274.950 532.950 277.050 535.050 ;
        RECT 268.950 527.100 271.050 529.200 ;
        RECT 269.400 526.050 270.600 527.100 ;
        RECT 275.400 526.050 276.600 532.950 ;
        RECT 268.950 523.950 271.050 526.050 ;
        RECT 271.950 523.950 274.050 526.050 ;
        RECT 274.950 523.950 277.050 526.050 ;
        RECT 262.950 511.950 265.050 514.050 ;
        RECT 272.400 511.050 273.600 523.950 ;
        RECT 281.400 520.050 282.600 538.950 ;
        RECT 292.950 527.100 295.050 529.200 ;
        RECT 293.400 526.050 294.600 527.100 ;
        RECT 289.950 523.950 292.050 526.050 ;
        RECT 292.950 523.950 295.050 526.050 ;
        RECT 283.950 520.950 286.050 523.050 ;
        RECT 290.400 522.000 291.600 523.950 ;
        RECT 280.950 514.950 283.050 520.050 ;
        RECT 271.950 508.950 274.050 511.050 ;
        RECT 262.950 499.950 265.050 502.050 ;
        RECT 277.950 500.400 280.050 502.500 ;
        RECT 259.950 496.950 262.050 499.050 ;
        RECT 263.400 493.050 264.600 499.950 ;
        RECT 268.950 495.000 271.050 499.050 ;
        RECT 269.400 493.050 270.600 495.000 ;
        RECT 274.950 494.400 277.050 496.500 ;
        RECT 275.400 493.050 276.600 494.400 ;
        RECT 259.950 490.950 262.050 493.050 ;
        RECT 262.950 490.950 265.050 493.050 ;
        RECT 265.950 490.950 268.050 493.050 ;
        RECT 268.950 490.950 271.050 493.050 ;
        RECT 274.950 490.950 277.050 493.050 ;
        RECT 260.400 489.900 261.600 490.950 ;
        RECT 259.950 487.800 262.050 489.900 ;
        RECT 262.950 481.950 265.050 484.050 ;
        RECT 253.950 475.950 256.050 478.050 ;
        RECT 263.400 474.600 264.600 481.950 ;
        RECT 266.400 478.050 267.600 490.950 ;
        RECT 278.850 485.400 280.050 500.400 ;
        RECT 277.950 483.300 280.050 485.400 ;
        RECT 278.850 479.700 280.050 483.300 ;
        RECT 265.950 475.950 268.050 478.050 ;
        RECT 277.950 477.600 280.050 479.700 ;
        RECT 263.400 473.400 267.600 474.600 ;
        RECT 259.950 463.950 262.050 466.050 ;
        RECT 253.950 458.400 256.050 460.500 ;
        RECT 247.950 451.950 250.050 454.050 ;
        RECT 245.400 449.400 249.600 450.600 ;
        RECT 248.400 448.050 249.600 449.400 ;
        RECT 247.950 445.950 250.050 448.050 ;
        RECT 254.100 438.600 255.300 458.400 ;
        RECT 260.400 450.600 261.600 463.950 ;
        RECT 257.400 449.400 264.600 450.600 ;
        RECT 257.400 448.050 258.600 449.400 ;
        RECT 256.950 445.950 259.050 448.050 ;
        RECT 253.950 436.500 256.050 438.600 ;
        RECT 241.950 424.950 244.050 427.050 ;
        RECT 259.950 424.950 262.050 427.050 ;
        RECT 253.950 422.400 256.050 424.500 ;
        RECT 244.950 416.100 247.050 418.200 ;
        RECT 250.950 416.400 253.050 418.500 ;
        RECT 245.400 415.050 246.600 416.100 ;
        RECT 251.400 415.050 252.600 416.400 ;
        RECT 241.950 412.950 244.050 415.050 ;
        RECT 244.950 412.950 247.050 415.050 ;
        RECT 250.950 412.950 253.050 415.050 ;
        RECT 238.950 411.600 241.050 412.050 ;
        RECT 236.400 410.400 241.050 411.600 ;
        RECT 238.950 409.950 241.050 410.400 ;
        RECT 239.400 402.600 240.600 409.950 ;
        RECT 242.400 406.050 243.600 412.950 ;
        RECT 254.850 407.400 256.050 422.400 ;
        RECT 241.950 403.950 244.050 406.050 ;
        RECT 247.950 403.950 250.050 406.050 ;
        RECT 253.950 405.300 256.050 407.400 ;
        RECT 239.400 401.400 243.600 402.600 ;
        RECT 220.950 397.950 223.050 400.050 ;
        RECT 232.950 397.950 235.050 400.050 ;
        RECT 221.400 364.050 222.600 397.950 ;
        RECT 232.950 380.400 235.050 382.500 ;
        RECT 226.950 371.400 229.050 373.500 ;
        RECT 227.400 370.050 228.600 371.400 ;
        RECT 226.950 367.950 229.050 370.050 ;
        RECT 220.950 361.950 223.050 364.050 ;
        RECT 211.950 358.500 214.050 360.600 ;
        RECT 217.950 358.950 220.050 361.050 ;
        RECT 233.100 360.600 234.300 380.400 ;
        RECT 238.950 379.950 241.050 382.050 ;
        RECT 239.400 372.600 240.600 379.950 ;
        RECT 236.400 371.400 240.600 372.600 ;
        RECT 236.400 370.050 237.600 371.400 ;
        RECT 235.950 367.950 238.050 370.050 ;
        RECT 238.950 364.950 241.050 367.050 ;
        RECT 239.400 361.050 240.600 364.950 ;
        RECT 232.950 358.500 235.050 360.600 ;
        RECT 238.950 358.950 241.050 361.050 ;
        RECT 242.400 355.050 243.600 401.400 ;
        RECT 244.950 382.950 247.050 385.050 ;
        RECT 245.400 366.900 246.600 382.950 ;
        RECT 248.400 373.200 249.600 403.950 ;
        RECT 254.850 401.700 256.050 405.300 ;
        RECT 253.950 399.600 256.050 401.700 ;
        RECT 260.400 385.050 261.600 424.950 ;
        RECT 263.400 411.600 264.600 449.400 ;
        RECT 266.400 430.050 267.600 473.400 ;
        RECT 284.400 463.050 285.600 520.950 ;
        RECT 289.950 517.950 292.050 522.000 ;
        RECT 299.400 517.050 300.600 565.800 ;
        RECT 311.400 562.050 312.600 568.950 ;
        RECT 326.400 562.050 327.600 568.950 ;
        RECT 332.400 565.050 333.600 568.950 ;
        RECT 328.950 563.400 333.600 565.050 ;
        RECT 328.950 562.950 333.000 563.400 ;
        RECT 310.950 559.950 313.050 562.050 ;
        RECT 325.950 559.950 328.050 562.050 ;
        RECT 311.400 535.050 312.600 559.950 ;
        RECT 313.950 538.950 316.050 541.050 ;
        RECT 304.950 532.950 307.050 535.050 ;
        RECT 301.950 529.950 304.050 532.050 ;
        RECT 302.400 519.600 303.600 529.950 ;
        RECT 305.400 522.600 306.600 532.950 ;
        RECT 310.950 529.950 313.050 535.050 ;
        RECT 314.400 526.050 315.600 538.950 ;
        RECT 325.950 537.300 328.050 539.400 ;
        RECT 341.400 538.050 342.600 571.950 ;
        RECT 355.950 561.600 358.050 562.050 ;
        RECT 359.400 561.600 360.600 595.950 ;
        RECT 362.400 595.050 363.600 601.950 ;
        RECT 361.950 592.950 364.050 595.050 ;
        RECT 371.400 573.600 372.600 622.950 ;
        RECT 380.400 610.050 381.600 664.950 ;
        RECT 386.400 661.050 387.600 667.950 ;
        RECT 385.950 658.950 388.050 661.050 ;
        RECT 400.950 658.950 403.050 661.050 ;
        RECT 388.950 655.950 391.050 658.050 ;
        RECT 389.400 649.050 390.600 655.950 ;
        RECT 401.400 652.200 402.600 658.950 ;
        RECT 394.950 650.100 397.050 652.200 ;
        RECT 400.950 650.100 403.050 652.200 ;
        RECT 395.400 649.050 396.600 650.100 ;
        RECT 385.950 646.950 388.050 649.050 ;
        RECT 388.950 646.950 391.050 649.050 ;
        RECT 391.950 646.950 394.050 649.050 ;
        RECT 394.950 646.950 397.050 649.050 ;
        RECT 386.400 645.900 387.600 646.950 ;
        RECT 392.400 645.900 393.600 646.950 ;
        RECT 385.950 643.800 388.050 645.900 ;
        RECT 391.950 643.800 394.050 645.900 ;
        RECT 385.950 631.950 388.050 634.050 ;
        RECT 373.950 607.950 376.050 610.050 ;
        RECT 379.950 607.950 382.050 610.050 ;
        RECT 382.950 607.950 385.050 613.050 ;
        RECT 374.400 600.900 375.600 607.950 ;
        RECT 380.400 604.050 381.600 607.950 ;
        RECT 386.400 604.050 387.600 631.950 ;
        RECT 397.950 625.950 400.050 628.050 ;
        RECT 391.950 619.950 394.050 622.050 ;
        RECT 392.400 604.050 393.600 619.950 ;
        RECT 379.950 601.950 382.050 604.050 ;
        RECT 382.950 601.950 385.050 604.050 ;
        RECT 385.950 601.950 388.050 604.050 ;
        RECT 388.950 601.950 391.050 604.050 ;
        RECT 391.950 601.950 394.050 604.050 ;
        RECT 383.400 600.900 384.600 601.950 ;
        RECT 373.950 598.800 376.050 600.900 ;
        RECT 382.950 598.800 385.050 600.900 ;
        RECT 389.400 592.050 390.600 601.950 ;
        RECT 398.400 601.050 399.600 625.950 ;
        RECT 397.950 598.950 400.050 601.050 ;
        RECT 388.950 589.950 391.050 592.050 ;
        RECT 385.950 583.950 388.050 586.050 ;
        RECT 355.950 560.400 360.600 561.600 ;
        RECT 368.400 572.400 372.600 573.600 ;
        RECT 355.950 559.950 358.050 560.400 ;
        RECT 326.850 533.700 328.050 537.300 ;
        RECT 334.950 535.950 337.050 538.050 ;
        RECT 340.950 535.950 343.050 538.050 ;
        RECT 346.950 536.400 349.050 538.500 ;
        RECT 325.950 531.600 328.050 533.700 ;
        RECT 310.950 523.950 313.050 526.050 ;
        RECT 313.950 523.950 316.050 526.050 ;
        RECT 316.950 523.950 319.050 526.050 ;
        RECT 322.950 523.950 325.050 526.050 ;
        RECT 305.400 521.400 309.600 522.600 ;
        RECT 302.400 518.400 306.600 519.600 ;
        RECT 286.950 514.950 289.050 517.050 ;
        RECT 298.950 514.950 301.050 517.050 ;
        RECT 287.400 496.500 288.600 514.950 ;
        RECT 298.950 500.400 301.050 502.500 ;
        RECT 286.950 494.400 289.050 496.500 ;
        RECT 287.400 469.050 288.600 494.400 ;
        RECT 292.950 490.950 295.050 493.050 ;
        RECT 293.400 481.050 294.600 490.950 ;
        RECT 292.950 478.950 295.050 481.050 ;
        RECT 299.100 480.600 300.300 500.400 ;
        RECT 305.400 496.050 306.600 518.400 ;
        RECT 304.950 493.950 307.050 496.050 ;
        RECT 301.950 490.950 304.050 493.050 ;
        RECT 302.400 489.600 303.600 490.950 ;
        RECT 301.950 487.500 304.050 489.600 ;
        RECT 298.950 478.500 301.050 480.600 ;
        RECT 304.950 478.950 307.050 481.050 ;
        RECT 298.950 472.950 301.050 475.050 ;
        RECT 286.950 466.950 289.050 469.050 ;
        RECT 283.950 460.950 286.050 463.050 ;
        RECT 289.950 459.300 292.050 461.400 ;
        RECT 290.850 455.700 292.050 459.300 ;
        RECT 271.950 450.000 274.050 454.050 ;
        RECT 289.950 453.600 292.050 455.700 ;
        RECT 272.400 448.050 273.600 450.000 ;
        RECT 277.950 449.100 280.050 451.200 ;
        RECT 278.400 448.050 279.600 449.100 ;
        RECT 271.950 445.950 274.050 448.050 ;
        RECT 274.950 445.950 277.050 448.050 ;
        RECT 277.950 445.950 280.050 448.050 ;
        RECT 286.950 445.950 289.050 448.050 ;
        RECT 275.400 436.050 276.600 445.950 ;
        RECT 283.950 442.950 286.050 445.050 ;
        RECT 287.400 444.000 288.600 445.950 ;
        RECT 274.950 433.950 277.050 436.050 ;
        RECT 265.950 427.950 268.050 430.050 ;
        RECT 274.950 422.400 277.050 424.500 ;
        RECT 268.950 412.950 271.050 415.050 ;
        RECT 262.950 409.500 265.050 411.600 ;
        RECT 259.950 382.950 262.050 385.050 ;
        RECT 260.400 379.050 261.600 382.950 ;
        RECT 263.400 382.050 264.600 409.500 ;
        RECT 262.950 379.950 265.050 382.050 ;
        RECT 259.950 376.950 262.050 379.050 ;
        RECT 265.950 373.950 268.050 376.050 ;
        RECT 247.950 371.100 250.050 373.200 ;
        RECT 253.950 371.100 256.050 373.200 ;
        RECT 259.950 371.100 262.050 373.200 ;
        RECT 254.400 370.050 255.600 371.100 ;
        RECT 260.400 370.050 261.600 371.100 ;
        RECT 250.950 367.950 253.050 370.050 ;
        RECT 253.950 367.950 256.050 370.050 ;
        RECT 256.950 367.950 259.050 370.050 ;
        RECT 259.950 367.950 262.050 370.050 ;
        RECT 251.400 366.900 252.600 367.950 ;
        RECT 244.950 364.800 247.050 366.900 ;
        RECT 250.950 364.800 253.050 366.900 ;
        RECT 257.400 361.050 258.600 367.950 ;
        RECT 256.950 358.950 259.050 361.050 ;
        RECT 256.950 355.800 259.050 357.900 ;
        RECT 229.950 352.950 232.050 355.050 ;
        RECT 241.950 352.950 244.050 355.050 ;
        RECT 217.950 343.950 220.050 346.050 ;
        RECT 205.950 334.950 208.050 337.050 ;
        RECT 211.950 334.950 214.050 337.050 ;
        RECT 212.400 333.000 213.600 334.950 ;
        RECT 211.950 328.950 214.050 333.000 ;
        RECT 199.950 325.950 202.050 328.050 ;
        RECT 212.400 325.050 213.600 328.950 ;
        RECT 218.400 325.050 219.600 343.950 ;
        RECT 223.950 338.100 226.050 340.200 ;
        RECT 224.400 331.050 225.600 338.100 ;
        RECT 230.400 337.050 231.600 352.950 ;
        RECT 241.950 346.950 244.050 349.050 ;
        RECT 235.950 338.100 238.050 340.200 ;
        RECT 236.400 337.050 237.600 338.100 ;
        RECT 229.950 334.950 232.050 337.050 ;
        RECT 232.950 334.950 235.050 337.050 ;
        RECT 235.950 334.950 238.050 337.050 ;
        RECT 233.400 333.900 234.600 334.950 ;
        RECT 232.950 331.800 235.050 333.900 ;
        RECT 223.950 328.950 226.050 331.050 ;
        RECT 229.950 328.950 232.050 331.050 ;
        RECT 211.950 322.950 214.050 325.050 ;
        RECT 217.950 322.950 220.050 325.050 ;
        RECT 190.950 307.950 193.050 310.050 ;
        RECT 196.950 307.950 199.050 310.050 ;
        RECT 214.950 307.950 217.050 310.050 ;
        RECT 157.950 303.300 160.050 305.400 ;
        RECT 157.950 299.700 159.150 303.300 ;
        RECT 172.950 302.400 175.050 304.500 ;
        RECT 193.950 303.300 196.050 305.400 ;
        RECT 157.950 297.600 160.050 299.700 ;
        RECT 151.950 293.400 154.050 295.500 ;
        RECT 142.950 277.950 145.050 280.050 ;
        RECT 148.950 277.950 151.050 280.050 ;
        RECT 139.950 274.950 142.050 277.050 ;
        RECT 106.950 259.950 109.050 262.050 ;
        RECT 109.950 260.100 112.050 262.200 ;
        RECT 112.950 259.950 115.050 262.050 ;
        RECT 121.950 260.100 124.050 262.200 ;
        RECT 127.950 260.100 130.050 262.200 ;
        RECT 136.950 260.100 139.050 262.200 ;
        RECT 79.950 256.950 82.050 259.050 ;
        RECT 85.950 256.950 88.050 259.050 ;
        RECT 100.950 256.950 103.050 259.050 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 80.400 250.050 81.600 256.950 ;
        RECT 79.950 247.950 82.050 250.050 ;
        RECT 80.400 232.050 81.600 247.950 ;
        RECT 104.400 244.050 105.600 256.950 ;
        RECT 113.400 255.900 114.600 259.950 ;
        RECT 122.400 259.050 123.600 260.100 ;
        RECT 128.400 259.050 129.600 260.100 ;
        RECT 118.950 256.950 121.050 259.050 ;
        RECT 121.950 256.950 124.050 259.050 ;
        RECT 124.950 256.950 127.050 259.050 ;
        RECT 127.950 256.950 130.050 259.050 ;
        RECT 130.950 256.950 133.050 259.050 ;
        RECT 119.400 255.900 120.600 256.950 ;
        RECT 112.950 253.800 115.050 255.900 ;
        RECT 118.950 253.800 121.050 255.900 ;
        RECT 103.950 243.600 106.050 244.050 ;
        RECT 103.950 242.400 108.600 243.600 ;
        RECT 103.950 241.950 106.050 242.400 ;
        RECT 79.950 229.950 82.050 232.050 ;
        RECT 67.950 220.950 70.050 223.050 ;
        RECT 91.950 220.950 94.050 223.050 ;
        RECT 73.950 215.100 76.050 217.200 ;
        RECT 79.800 215.100 81.900 217.200 ;
        RECT 74.400 214.050 75.600 215.100 ;
        RECT 70.950 211.950 73.050 214.050 ;
        RECT 73.950 211.950 76.050 214.050 ;
        RECT 71.400 210.000 72.600 211.950 ;
        RECT 64.950 205.950 67.050 208.050 ;
        RECT 70.950 205.950 73.050 210.000 ;
        RECT 80.400 205.050 81.600 215.100 ;
        RECT 82.950 214.950 85.050 217.050 ;
        RECT 83.400 210.900 84.600 214.950 ;
        RECT 92.400 214.050 93.600 220.950 ;
        RECT 97.950 216.000 100.050 220.050 ;
        RECT 98.400 214.050 99.600 216.000 ;
        RECT 91.950 211.950 94.050 214.050 ;
        RECT 94.950 211.950 97.050 214.050 ;
        RECT 97.950 211.950 100.050 214.050 ;
        RECT 100.950 211.950 103.050 214.050 ;
        RECT 82.950 208.800 85.050 210.900 ;
        RECT 52.950 202.950 55.050 205.050 ;
        RECT 67.950 202.950 70.050 205.050 ;
        RECT 79.950 202.950 82.050 205.050 ;
        RECT 52.950 196.950 55.050 199.050 ;
        RECT 46.950 190.950 49.050 193.050 ;
        RECT 38.400 181.050 39.600 182.100 ;
        RECT 43.950 181.950 46.050 184.050 ;
        RECT 34.950 178.950 37.050 181.050 ;
        RECT 37.950 178.950 40.050 181.050 ;
        RECT 40.950 178.950 43.050 181.050 ;
        RECT 35.400 177.900 36.600 178.950 ;
        RECT 34.950 175.800 37.050 177.900 ;
        RECT 41.400 177.000 42.600 178.950 ;
        RECT 40.950 172.950 43.050 177.000 ;
        RECT 47.400 175.050 48.600 190.950 ;
        RECT 49.950 182.100 52.050 184.200 ;
        RECT 46.950 172.950 49.050 175.050 ;
        RECT 47.400 145.050 48.600 172.950 ;
        RECT 46.950 142.950 49.050 145.050 ;
        RECT 20.400 131.400 25.050 133.050 ;
        RECT 21.000 130.950 25.050 131.400 ;
        RECT 28.950 130.950 31.050 133.050 ;
        RECT 50.400 130.050 51.600 182.100 ;
        RECT 53.400 177.900 54.600 196.950 ;
        RECT 61.950 182.100 64.050 184.200 ;
        RECT 62.400 181.050 63.600 182.100 ;
        RECT 68.400 181.050 69.600 202.950 ;
        RECT 79.950 199.800 82.050 201.900 ;
        RECT 73.950 196.950 76.050 199.050 ;
        RECT 58.950 178.950 61.050 181.050 ;
        RECT 61.950 178.950 64.050 181.050 ;
        RECT 64.950 178.950 67.050 181.050 ;
        RECT 67.950 178.950 70.050 181.050 ;
        RECT 59.400 177.900 60.600 178.950 ;
        RECT 65.400 177.900 66.600 178.950 ;
        RECT 52.950 175.800 55.050 177.900 ;
        RECT 58.950 175.800 61.050 177.900 ;
        RECT 64.950 175.800 67.050 177.900 ;
        RECT 74.400 175.050 75.600 196.950 ;
        RECT 80.400 181.050 81.600 199.800 ;
        RECT 95.400 199.050 96.600 211.950 ;
        RECT 101.400 205.050 102.600 211.950 ;
        RECT 107.400 210.900 108.600 242.400 ;
        RECT 125.400 223.050 126.600 256.950 ;
        RECT 131.400 255.900 132.600 256.950 ;
        RECT 137.400 256.050 138.600 260.100 ;
        RECT 130.950 253.800 133.050 255.900 ;
        RECT 136.950 253.950 139.050 256.050 ;
        RECT 140.400 244.050 141.600 274.950 ;
        RECT 143.400 262.050 144.600 277.950 ;
        RECT 152.400 277.050 153.600 293.400 ;
        RECT 157.950 282.600 159.150 297.600 ;
        RECT 169.950 293.400 172.050 298.050 ;
        RECT 170.400 292.050 171.600 293.400 ;
        RECT 160.950 289.950 163.050 292.050 ;
        RECT 169.950 289.950 172.050 292.050 ;
        RECT 161.400 288.600 162.600 289.950 ;
        RECT 161.400 287.400 165.600 288.600 ;
        RECT 164.400 283.050 165.600 287.400 ;
        RECT 166.950 286.950 169.050 289.050 ;
        RECT 157.950 280.500 160.050 282.600 ;
        RECT 163.950 280.950 166.050 283.050 ;
        RECT 151.950 274.950 154.050 277.050 ;
        RECT 148.950 265.950 151.050 268.050 ;
        RECT 160.950 266.400 163.050 268.500 ;
        RECT 142.950 259.950 145.050 262.050 ;
        RECT 149.400 259.050 150.600 265.950 ;
        RECT 157.950 260.400 160.050 262.500 ;
        RECT 158.400 259.050 159.600 260.400 ;
        RECT 145.950 256.950 148.050 259.050 ;
        RECT 148.950 256.950 151.050 259.050 ;
        RECT 151.950 256.950 154.050 259.050 ;
        RECT 157.950 256.950 160.050 259.050 ;
        RECT 146.400 250.050 147.600 256.950 ;
        RECT 152.400 255.900 153.600 256.950 ;
        RECT 151.950 253.800 154.050 255.900 ;
        RECT 161.850 251.400 163.050 266.400 ;
        RECT 145.950 247.950 148.050 250.050 ;
        RECT 160.950 249.300 163.050 251.400 ;
        RECT 161.850 245.700 163.050 249.300 ;
        RECT 139.950 241.950 142.050 244.050 ;
        RECT 160.950 243.600 163.050 245.700 ;
        RECT 167.400 229.050 168.600 286.950 ;
        RECT 173.700 282.600 174.900 302.400 ;
        RECT 193.950 299.700 195.150 303.300 ;
        RECT 193.950 297.600 196.050 299.700 ;
        RECT 179.400 293.400 186.600 294.600 ;
        RECT 179.400 292.050 180.600 293.400 ;
        RECT 178.950 289.950 181.050 292.050 ;
        RECT 185.400 283.050 186.600 293.400 ;
        RECT 172.950 280.500 175.050 282.600 ;
        RECT 184.950 280.950 187.050 283.050 ;
        RECT 193.950 282.600 195.150 297.600 ;
        RECT 215.400 292.050 216.600 307.950 ;
        RECT 221.400 293.400 228.600 294.600 ;
        RECT 221.400 292.050 222.600 293.400 ;
        RECT 196.950 289.950 199.050 292.050 ;
        RECT 214.950 289.950 217.050 292.050 ;
        RECT 217.950 289.950 220.050 292.050 ;
        RECT 220.950 289.950 223.050 292.050 ;
        RECT 197.400 288.600 198.600 289.950 ;
        RECT 197.400 287.400 201.600 288.600 ;
        RECT 193.950 280.500 196.050 282.600 ;
        RECT 169.950 274.950 172.050 277.050 ;
        RECT 127.950 226.950 130.050 229.050 ;
        RECT 166.950 226.950 169.050 229.050 ;
        RECT 124.950 220.950 127.050 223.050 ;
        RECT 124.950 217.800 127.050 219.900 ;
        RECT 115.950 215.100 118.050 217.200 ;
        RECT 116.400 214.050 117.600 215.100 ;
        RECT 112.950 211.950 115.050 214.050 ;
        RECT 115.950 211.950 118.050 214.050 ;
        RECT 118.950 211.950 121.050 214.050 ;
        RECT 113.400 210.900 114.600 211.950 ;
        RECT 119.400 210.900 120.600 211.950 ;
        RECT 106.950 208.800 109.050 210.900 ;
        RECT 112.950 208.800 115.050 210.900 ;
        RECT 118.950 208.800 121.050 210.900 ;
        RECT 100.950 202.950 103.050 205.050 ;
        RECT 97.950 199.950 100.050 202.050 ;
        RECT 94.950 196.950 97.050 199.050 ;
        RECT 98.400 196.050 99.600 199.950 ;
        RECT 125.400 199.050 126.600 217.800 ;
        RECT 124.950 196.950 127.050 199.050 ;
        RECT 97.950 193.950 100.050 196.050 ;
        RECT 100.950 188.400 103.050 190.500 ;
        RECT 121.950 188.400 124.050 190.500 ;
        RECT 85.950 182.100 88.050 184.200 ;
        RECT 97.950 182.400 100.050 184.500 ;
        RECT 86.400 181.050 87.600 182.100 ;
        RECT 98.400 181.050 99.600 182.400 ;
        RECT 79.950 178.950 82.050 181.050 ;
        RECT 82.950 178.950 85.050 181.050 ;
        RECT 85.950 178.950 88.050 181.050 ;
        RECT 88.950 178.950 91.050 181.050 ;
        RECT 97.950 178.950 100.050 181.050 ;
        RECT 83.400 177.900 84.600 178.950 ;
        RECT 82.950 175.800 85.050 177.900 ;
        RECT 73.950 172.950 76.050 175.050 ;
        RECT 79.950 172.950 82.050 175.050 ;
        RECT 80.400 145.050 81.600 172.950 ;
        RECT 73.950 142.950 76.050 145.050 ;
        RECT 79.950 142.950 82.050 145.050 ;
        RECT 55.950 137.100 58.050 139.200 ;
        RECT 56.400 136.050 57.600 137.100 ;
        RECT 61.950 136.950 64.050 139.050 ;
        RECT 55.950 133.950 58.050 136.050 ;
        RECT 19.950 127.950 22.050 130.050 ;
        RECT 49.950 127.950 52.050 130.050 ;
        RECT 55.950 127.950 58.050 130.050 ;
        RECT 16.500 108.300 18.600 110.400 ;
        RECT 20.400 108.900 21.600 127.950 ;
        RECT 43.950 109.950 46.050 112.050 ;
        RECT 14.400 103.050 15.600 105.600 ;
        RECT 4.950 100.950 7.050 103.050 ;
        RECT 13.950 100.950 16.050 103.050 ;
        RECT 16.950 102.900 17.850 108.300 ;
        RECT 19.800 106.800 21.900 108.900 ;
        RECT 23.700 105.900 25.800 107.700 ;
        RECT 18.750 104.700 27.300 105.900 ;
        RECT 18.750 103.800 20.850 104.700 ;
        RECT 16.950 101.700 23.700 102.900 ;
        RECT 5.400 91.050 6.600 100.950 ;
        RECT 16.950 94.500 18.000 101.700 ;
        RECT 19.800 98.100 21.900 100.200 ;
        RECT 22.800 99.300 23.700 101.700 ;
        RECT 20.400 95.550 21.600 98.100 ;
        RECT 22.800 97.200 24.900 99.300 ;
        RECT 26.400 95.700 27.300 104.700 ;
        RECT 44.400 103.050 45.600 109.950 ;
        RECT 49.950 104.100 52.050 106.200 ;
        RECT 50.400 103.050 51.600 104.100 ;
        RECT 28.500 100.950 30.600 103.050 ;
        RECT 29.400 98.400 30.600 100.950 ;
        RECT 31.950 97.950 34.050 103.050 ;
        RECT 43.950 100.950 46.050 103.050 ;
        RECT 46.950 100.950 49.050 103.050 ;
        RECT 49.950 100.950 52.050 103.050 ;
        RECT 47.400 99.900 48.600 100.950 ;
        RECT 46.950 97.800 49.050 99.900 ;
        RECT 16.500 92.400 18.600 94.500 ;
        RECT 26.100 93.600 28.200 95.700 ;
        RECT 4.950 88.950 7.050 91.050 ;
        RECT 16.950 88.950 19.050 91.050 ;
        RECT 17.400 73.050 18.600 88.950 ;
        RECT 16.950 70.950 19.050 73.050 ;
        RECT 52.950 70.950 55.050 73.050 ;
        RECT 17.400 58.050 18.600 70.950 ;
        RECT 25.950 58.950 28.050 61.050 ;
        RECT 34.950 59.100 37.050 61.200 ;
        RECT 13.950 55.950 16.050 58.050 ;
        RECT 16.950 55.950 19.050 58.050 ;
        RECT 19.950 55.950 22.050 58.050 ;
        RECT 14.400 40.050 15.600 55.950 ;
        RECT 20.400 54.600 21.600 55.950 ;
        RECT 26.400 54.600 27.600 58.950 ;
        RECT 35.400 58.050 36.600 59.100 ;
        RECT 53.400 58.050 54.600 70.950 ;
        RECT 56.400 67.050 57.600 127.950 ;
        RECT 62.400 105.600 63.600 136.950 ;
        RECT 74.400 136.050 75.600 142.950 ;
        RECT 83.400 141.600 84.600 175.800 ;
        RECT 89.400 172.050 90.600 178.950 ;
        RECT 101.850 173.400 103.050 188.400 ;
        RECT 115.950 178.950 118.050 181.050 ;
        RECT 88.950 169.950 91.050 172.050 ;
        RECT 100.950 171.300 103.050 173.400 ;
        RECT 101.850 167.700 103.050 171.300 ;
        RECT 100.950 165.600 103.050 167.700 ;
        RECT 112.950 142.950 115.050 145.050 ;
        RECT 80.400 140.400 84.600 141.600 ;
        RECT 80.400 136.050 81.600 140.400 ;
        RECT 85.950 139.950 88.050 142.050 ;
        RECT 91.950 141.600 94.050 142.200 ;
        RECT 103.950 141.600 106.050 142.050 ;
        RECT 91.950 140.400 106.050 141.600 ;
        RECT 91.950 140.100 94.050 140.400 ;
        RECT 103.950 139.950 106.050 140.400 ;
        RECT 106.950 139.950 109.050 142.050 ;
        RECT 73.950 133.950 76.050 136.050 ;
        RECT 76.950 133.950 79.050 136.050 ;
        RECT 79.950 133.950 82.050 136.050 ;
        RECT 77.400 132.900 78.600 133.950 ;
        RECT 86.400 133.050 87.600 139.950 ;
        RECT 91.950 136.950 94.050 139.050 ;
        RECT 100.950 137.100 103.050 139.200 ;
        RECT 92.400 136.050 93.600 136.950 ;
        RECT 101.400 136.050 102.600 137.100 ;
        RECT 91.950 133.950 94.050 136.050 ;
        RECT 97.950 133.950 100.050 136.050 ;
        RECT 100.950 133.950 103.050 136.050 ;
        RECT 76.950 130.800 79.050 132.900 ;
        RECT 85.950 130.950 88.050 133.050 ;
        RECT 98.400 132.000 99.600 133.950 ;
        RECT 79.950 127.950 82.050 130.050 ;
        RECT 91.950 127.950 94.050 130.050 ;
        RECT 97.950 127.950 100.050 132.000 ;
        RECT 76.950 109.950 79.050 112.050 ;
        RECT 59.400 104.400 63.600 105.600 ;
        RECT 59.400 82.050 60.600 104.400 ;
        RECT 67.950 104.100 70.050 106.200 ;
        RECT 68.400 103.050 69.600 104.100 ;
        RECT 64.950 100.950 67.050 103.050 ;
        RECT 67.950 100.950 70.050 103.050 ;
        RECT 70.950 100.950 73.050 103.050 ;
        RECT 61.950 97.950 64.050 100.050 ;
        RECT 62.400 94.050 63.600 97.950 ;
        RECT 61.950 91.950 64.050 94.050 ;
        RECT 58.950 79.950 61.050 82.050 ;
        RECT 55.950 64.950 58.050 67.050 ;
        RECT 62.400 64.050 63.600 91.950 ;
        RECT 65.400 88.050 66.600 100.950 ;
        RECT 64.950 85.950 67.050 88.050 ;
        RECT 71.400 73.050 72.600 100.950 ;
        RECT 73.950 97.950 76.050 100.050 ;
        RECT 70.950 70.950 73.050 73.050 ;
        RECT 70.950 64.950 73.050 67.050 ;
        RECT 61.950 61.950 64.050 64.050 ;
        RECT 58.950 59.100 61.050 61.200 ;
        RECT 67.950 59.100 70.050 61.200 ;
        RECT 59.400 58.050 60.600 59.100 ;
        RECT 31.950 55.950 34.050 58.050 ;
        RECT 34.950 55.950 37.050 58.050 ;
        RECT 37.950 55.950 40.050 58.050 ;
        RECT 52.950 55.950 55.050 58.050 ;
        RECT 55.950 55.950 58.050 58.050 ;
        RECT 58.950 55.950 61.050 58.050 ;
        RECT 61.950 55.950 64.050 58.050 ;
        RECT 20.400 53.400 27.600 54.600 ;
        RECT 32.400 49.050 33.600 55.950 ;
        RECT 31.950 46.950 34.050 49.050 ;
        RECT 13.950 37.950 16.050 40.050 ;
        RECT 14.400 31.050 15.600 37.950 ;
        RECT 32.400 34.050 33.600 46.950 ;
        RECT 22.950 31.950 25.050 34.050 ;
        RECT 31.950 31.950 34.050 34.050 ;
        RECT 13.950 28.950 16.050 31.050 ;
        RECT 16.950 26.100 19.050 28.200 ;
        RECT 17.400 25.050 18.600 26.100 ;
        RECT 13.950 22.950 16.050 25.050 ;
        RECT 16.950 22.950 19.050 25.050 ;
        RECT 14.400 21.900 15.600 22.950 ;
        RECT 23.400 21.900 24.600 31.950 ;
        RECT 31.950 26.100 34.050 28.200 ;
        RECT 38.400 28.050 39.600 55.950 ;
        RECT 56.400 54.900 57.600 55.950 ;
        RECT 55.950 52.800 58.050 54.900 ;
        RECT 46.950 43.950 49.050 46.050 ;
        RECT 47.400 40.050 48.600 43.950 ;
        RECT 58.950 40.950 61.050 43.050 ;
        RECT 62.400 42.600 63.600 55.950 ;
        RECT 64.950 52.950 67.050 55.050 ;
        RECT 65.400 46.050 66.600 52.950 ;
        RECT 64.950 43.950 67.050 46.050 ;
        RECT 68.400 42.600 69.600 59.100 ;
        RECT 71.400 43.050 72.600 64.950 ;
        RECT 74.400 48.600 75.600 97.950 ;
        RECT 77.400 97.050 78.600 109.950 ;
        RECT 76.950 94.950 79.050 97.050 ;
        RECT 80.400 85.050 81.600 127.950 ;
        RECT 85.950 112.950 88.050 115.050 ;
        RECT 86.400 103.050 87.600 112.950 ;
        RECT 92.400 106.200 93.600 127.950 ;
        RECT 98.400 124.050 99.600 127.950 ;
        RECT 97.950 121.950 100.050 124.050 ;
        RECT 107.400 115.050 108.600 139.950 ;
        RECT 97.950 112.950 100.050 115.050 ;
        RECT 106.950 112.950 109.050 115.050 ;
        RECT 91.950 104.100 94.050 106.200 ;
        RECT 92.400 103.050 93.600 104.100 ;
        RECT 85.950 100.950 88.050 103.050 ;
        RECT 88.950 100.950 91.050 103.050 ;
        RECT 91.950 100.950 94.050 103.050 ;
        RECT 89.400 99.000 90.600 100.950 ;
        RECT 88.950 94.950 91.050 99.000 ;
        RECT 79.950 82.950 82.050 85.050 ;
        RECT 91.950 82.950 94.050 85.050 ;
        RECT 79.950 59.100 82.050 61.200 ;
        RECT 85.950 60.000 88.050 64.050 ;
        RECT 92.400 61.050 93.600 82.950 ;
        RECT 94.950 73.950 97.050 76.050 ;
        RECT 80.400 58.050 81.600 59.100 ;
        RECT 86.400 58.050 87.600 60.000 ;
        RECT 91.950 58.950 94.050 61.050 ;
        RECT 79.950 55.950 82.050 58.050 ;
        RECT 82.950 55.950 85.050 58.050 ;
        RECT 85.950 55.950 88.050 58.050 ;
        RECT 88.950 55.950 91.050 58.050 ;
        RECT 83.400 54.000 84.600 55.950 ;
        RECT 82.950 49.950 85.050 54.000 ;
        RECT 89.400 51.600 90.600 55.950 ;
        RECT 91.950 52.950 94.050 55.050 ;
        RECT 86.400 50.400 90.600 51.600 ;
        RECT 86.400 48.600 87.600 50.400 ;
        RECT 74.400 47.400 87.600 48.600 ;
        RECT 92.400 46.050 93.600 52.950 ;
        RECT 95.400 52.050 96.600 73.950 ;
        RECT 98.400 64.050 99.600 112.950 ;
        RECT 103.950 104.100 106.050 106.200 ;
        RECT 104.400 103.050 105.600 104.100 ;
        RECT 103.950 100.950 106.050 103.050 ;
        RECT 106.950 100.950 109.050 103.050 ;
        RECT 107.400 99.900 108.600 100.950 ;
        RECT 106.950 97.800 109.050 99.900 ;
        RECT 97.950 61.950 100.050 64.050 ;
        RECT 113.400 61.200 114.600 142.950 ;
        RECT 116.400 133.050 117.600 178.950 ;
        RECT 122.100 168.600 123.300 188.400 ;
        RECT 128.400 184.050 129.600 226.950 ;
        RECT 157.950 220.950 160.050 223.050 ;
        RECT 170.400 222.600 171.600 274.950 ;
        RECT 200.400 271.050 201.600 287.400 ;
        RECT 199.950 268.950 202.050 271.050 ;
        RECT 181.950 266.400 184.050 268.500 ;
        RECT 175.950 256.950 178.050 259.050 ;
        RECT 176.400 255.600 177.600 256.950 ;
        RECT 175.950 253.500 178.050 255.600 ;
        RECT 182.100 246.600 183.300 266.400 ;
        RECT 196.950 265.950 199.050 268.050 ;
        RECT 190.950 259.950 193.050 262.050 ;
        RECT 184.950 256.950 187.050 259.050 ;
        RECT 185.400 255.600 186.600 256.950 ;
        RECT 191.400 255.600 192.600 259.950 ;
        RECT 193.950 256.950 196.050 259.050 ;
        RECT 185.400 254.400 189.600 255.600 ;
        RECT 181.950 244.500 184.050 246.600 ;
        RECT 188.400 229.050 189.600 254.400 ;
        RECT 190.950 253.500 193.050 255.600 ;
        RECT 194.400 250.050 195.600 256.950 ;
        RECT 197.400 255.900 198.600 265.950 ;
        RECT 205.950 260.100 208.050 262.200 ;
        RECT 211.950 260.100 214.050 262.200 ;
        RECT 206.400 259.050 207.600 260.100 ;
        RECT 212.400 259.050 213.600 260.100 ;
        RECT 202.950 256.950 205.050 259.050 ;
        RECT 205.950 256.950 208.050 259.050 ;
        RECT 208.950 256.950 211.050 259.050 ;
        RECT 211.950 256.950 214.050 259.050 ;
        RECT 203.400 255.900 204.600 256.950 ;
        RECT 209.400 255.900 210.600 256.950 ;
        RECT 218.400 255.900 219.600 289.950 ;
        RECT 227.400 289.050 228.600 293.400 ;
        RECT 226.950 286.950 229.050 289.050 ;
        RECT 220.950 280.950 223.050 283.050 ;
        RECT 221.400 262.050 222.600 280.950 ;
        RECT 230.400 280.050 231.600 328.950 ;
        RECT 242.400 313.050 243.600 346.950 ;
        RECT 250.950 338.100 253.050 340.200 ;
        RECT 251.400 337.050 252.600 338.100 ;
        RECT 257.400 337.050 258.600 355.800 ;
        RECT 262.950 349.950 265.050 352.050 ;
        RECT 263.400 340.200 264.600 349.950 ;
        RECT 262.950 338.100 265.050 340.200 ;
        RECT 247.950 334.950 250.050 337.050 ;
        RECT 250.950 334.950 253.050 337.050 ;
        RECT 253.950 334.950 256.050 337.050 ;
        RECT 256.950 334.950 259.050 337.050 ;
        RECT 248.400 333.000 249.600 334.950 ;
        RECT 254.400 333.900 255.600 334.950 ;
        RECT 247.950 328.950 250.050 333.000 ;
        RECT 253.950 331.800 256.050 333.900 ;
        RECT 263.400 333.600 264.600 338.100 ;
        RECT 260.400 332.400 264.600 333.600 ;
        RECT 256.950 328.950 259.050 331.050 ;
        RECT 235.950 310.950 238.050 313.050 ;
        RECT 241.950 310.950 244.050 313.050 ;
        RECT 236.400 292.050 237.600 310.950 ;
        RECT 241.950 304.950 244.050 307.050 ;
        RECT 242.400 292.050 243.600 304.950 ;
        RECT 250.950 303.300 253.050 305.400 ;
        RECT 251.850 299.700 253.050 303.300 ;
        RECT 250.950 297.600 253.050 299.700 ;
        RECT 235.950 289.950 238.050 292.050 ;
        RECT 238.950 289.950 241.050 292.050 ;
        RECT 241.950 289.950 244.050 292.050 ;
        RECT 247.950 289.950 250.050 292.050 ;
        RECT 239.400 288.900 240.600 289.950 ;
        RECT 238.950 286.800 241.050 288.900 ;
        RECT 248.400 288.600 249.600 289.950 ;
        RECT 247.950 286.500 250.050 288.600 ;
        RECT 244.950 280.950 247.050 283.050 ;
        RECT 251.850 282.600 253.050 297.600 ;
        RECT 257.400 289.050 258.600 328.950 ;
        RECT 256.950 286.950 259.050 289.050 ;
        RECT 229.950 277.950 232.050 280.050 ;
        RECT 226.950 274.950 229.050 277.050 ;
        RECT 220.950 259.950 223.050 262.050 ;
        RECT 227.400 259.050 228.600 274.950 ;
        RECT 232.950 271.950 235.050 274.050 ;
        RECT 233.400 259.050 234.600 271.950 ;
        RECT 238.950 268.950 241.050 271.050 ;
        RECT 223.950 256.950 226.050 259.050 ;
        RECT 226.950 256.950 229.050 259.050 ;
        RECT 229.950 256.950 232.050 259.050 ;
        RECT 232.950 256.950 235.050 259.050 ;
        RECT 224.400 255.900 225.600 256.950 ;
        RECT 196.950 253.800 199.050 255.900 ;
        RECT 202.950 253.800 205.050 255.900 ;
        RECT 208.950 253.800 211.050 255.900 ;
        RECT 217.950 253.800 220.050 255.900 ;
        RECT 223.950 253.800 226.050 255.900 ;
        RECT 230.400 250.050 231.600 256.950 ;
        RECT 193.950 247.950 196.050 250.050 ;
        RECT 199.950 247.950 202.050 250.050 ;
        RECT 205.950 247.950 208.050 250.050 ;
        RECT 229.950 247.950 232.050 250.050 ;
        RECT 190.950 241.950 193.050 244.050 ;
        RECT 187.950 226.950 190.050 229.050 ;
        RECT 170.400 221.400 174.600 222.600 ;
        RECT 130.950 214.950 133.050 217.050 ;
        RECT 139.950 215.100 142.050 217.200 ;
        RECT 127.950 181.950 130.050 184.050 ;
        RECT 124.950 178.950 127.050 181.050 ;
        RECT 125.400 177.600 126.600 178.950 ;
        RECT 124.950 175.500 127.050 177.600 ;
        RECT 131.400 175.050 132.600 214.950 ;
        RECT 140.400 214.050 141.600 215.100 ;
        RECT 158.400 214.050 159.600 220.950 ;
        RECT 163.950 215.100 166.050 217.200 ;
        RECT 169.950 215.100 172.050 220.050 ;
        RECT 164.400 214.050 165.600 215.100 ;
        RECT 136.950 211.950 139.050 214.050 ;
        RECT 139.950 211.950 142.050 214.050 ;
        RECT 142.950 211.950 145.050 214.050 ;
        RECT 157.950 211.950 160.050 214.050 ;
        RECT 160.950 211.950 163.050 214.050 ;
        RECT 163.950 211.950 166.050 214.050 ;
        RECT 166.950 211.950 169.050 214.050 ;
        RECT 137.400 205.050 138.600 211.950 ;
        RECT 143.400 205.050 144.600 211.950 ;
        RECT 154.950 208.800 157.050 210.900 ;
        RECT 136.950 202.950 139.050 205.050 ;
        RECT 142.950 202.950 145.050 205.050 ;
        RECT 151.950 202.950 154.050 205.050 ;
        RECT 143.400 196.050 144.600 202.950 ;
        RECT 142.950 193.950 145.050 196.050 ;
        RECT 133.950 181.950 136.050 184.050 ;
        RECT 142.950 182.100 145.050 184.200 ;
        RECT 130.950 172.950 133.050 175.050 ;
        RECT 134.400 172.050 135.600 181.950 ;
        RECT 143.400 181.050 144.600 182.100 ;
        RECT 139.950 178.950 142.050 181.050 ;
        RECT 142.950 178.950 145.050 181.050 ;
        RECT 145.950 178.950 148.050 181.050 ;
        RECT 140.400 177.900 141.600 178.950 ;
        RECT 139.950 175.800 142.050 177.900 ;
        RECT 136.950 172.950 139.050 175.050 ;
        RECT 133.950 169.950 136.050 172.050 ;
        RECT 121.950 166.500 124.050 168.600 ;
        RECT 121.950 138.000 124.050 142.050 ;
        RECT 122.400 136.050 123.600 138.000 ;
        RECT 127.950 137.100 130.050 139.200 ;
        RECT 128.400 136.050 129.600 137.100 ;
        RECT 121.950 133.950 124.050 136.050 ;
        RECT 124.950 133.950 127.050 136.050 ;
        RECT 127.950 133.950 130.050 136.050 ;
        RECT 130.950 133.950 133.050 136.050 ;
        RECT 115.950 130.950 118.050 133.050 ;
        RECT 125.400 132.900 126.600 133.950 ;
        RECT 131.400 132.900 132.600 133.950 ;
        RECT 124.950 130.800 127.050 132.900 ;
        RECT 130.950 130.800 133.050 132.900 ;
        RECT 115.800 104.100 117.900 106.200 ;
        RECT 118.950 104.100 121.050 106.200 ;
        RECT 124.950 104.100 127.050 106.200 ;
        RECT 130.950 104.100 133.050 106.200 ;
        RECT 116.400 100.050 117.600 104.100 ;
        RECT 115.950 97.950 118.050 100.050 ;
        RECT 116.400 88.050 117.600 97.950 ;
        RECT 119.400 97.050 120.600 104.100 ;
        RECT 125.400 103.050 126.600 104.100 ;
        RECT 131.400 103.050 132.600 104.100 ;
        RECT 124.950 100.950 127.050 103.050 ;
        RECT 127.950 100.950 130.050 103.050 ;
        RECT 130.950 100.950 133.050 103.050 ;
        RECT 128.400 99.900 129.600 100.950 ;
        RECT 127.950 97.800 130.050 99.900 ;
        RECT 118.950 94.950 121.050 97.050 ;
        RECT 115.950 85.950 118.050 88.050 ;
        RECT 137.400 85.050 138.600 172.950 ;
        RECT 146.400 154.050 147.600 178.950 ;
        RECT 152.400 177.900 153.600 202.950 ;
        RECT 151.950 175.800 154.050 177.900 ;
        RECT 148.950 169.950 151.050 172.050 ;
        RECT 145.950 151.950 148.050 154.050 ;
        RECT 145.950 141.600 148.050 142.050 ;
        RECT 149.400 141.600 150.600 169.950 ;
        RECT 155.400 157.050 156.600 208.800 ;
        RECT 161.400 207.600 162.600 211.950 ;
        RECT 167.400 210.900 168.600 211.950 ;
        RECT 166.950 208.800 169.050 210.900 ;
        RECT 158.400 206.400 162.600 207.600 ;
        RECT 154.950 154.950 157.050 157.050 ;
        RECT 145.950 140.400 150.600 141.600 ;
        RECT 145.950 139.950 148.050 140.400 ;
        RECT 146.400 136.050 147.600 139.950 ;
        RECT 151.950 137.100 154.050 139.200 ;
        RECT 152.400 136.050 153.600 137.100 ;
        RECT 142.950 133.950 145.050 136.050 ;
        RECT 145.950 133.950 148.050 136.050 ;
        RECT 148.950 133.950 151.050 136.050 ;
        RECT 151.950 133.950 154.050 136.050 ;
        RECT 143.400 124.050 144.600 133.950 ;
        RECT 149.400 132.900 150.600 133.950 ;
        RECT 148.950 130.800 151.050 132.900 ;
        RECT 142.950 121.950 145.050 124.050 ;
        RECT 158.400 112.050 159.600 206.400 ;
        RECT 173.400 205.050 174.600 221.400 ;
        RECT 181.950 215.100 184.050 217.200 ;
        RECT 182.400 214.050 183.600 215.100 ;
        RECT 191.400 214.050 192.600 241.950 ;
        RECT 178.950 211.950 181.050 214.050 ;
        RECT 181.950 211.950 184.050 214.050 ;
        RECT 184.950 211.950 187.050 214.050 ;
        RECT 190.950 211.950 193.050 214.050 ;
        RECT 179.400 210.900 180.600 211.950 ;
        RECT 178.950 208.800 181.050 210.900 ;
        RECT 180.000 207.750 183.000 208.050 ;
        RECT 178.950 205.950 184.050 207.750 ;
        RECT 178.950 205.650 181.050 205.950 ;
        RECT 181.950 205.650 184.050 205.950 ;
        RECT 172.950 202.950 175.050 205.050 ;
        RECT 166.950 196.950 169.050 199.050 ;
        RECT 167.400 181.050 168.600 196.950 ;
        RECT 173.400 196.050 174.600 202.950 ;
        RECT 185.400 202.050 186.600 211.950 ;
        RECT 196.950 202.950 199.050 205.050 ;
        RECT 178.950 199.950 181.050 202.050 ;
        RECT 184.950 199.950 187.050 202.050 ;
        RECT 172.950 193.950 175.050 196.050 ;
        RECT 173.400 181.050 174.600 193.950 ;
        RECT 163.950 178.950 166.050 181.050 ;
        RECT 166.950 178.950 169.050 181.050 ;
        RECT 169.950 178.950 172.050 181.050 ;
        RECT 172.950 178.950 175.050 181.050 ;
        RECT 164.400 177.900 165.600 178.950 ;
        RECT 163.950 175.800 166.050 177.900 ;
        RECT 170.400 169.050 171.600 178.950 ;
        RECT 175.950 172.950 178.050 177.900 ;
        RECT 169.950 166.950 172.050 169.050 ;
        RECT 179.400 160.050 180.600 199.950 ;
        RECT 181.950 181.950 184.050 187.050 ;
        RECT 187.950 182.100 190.050 184.200 ;
        RECT 188.400 181.050 189.600 182.100 ;
        RECT 184.950 178.950 187.050 181.050 ;
        RECT 187.950 178.950 190.050 181.050 ;
        RECT 190.950 178.950 193.050 181.050 ;
        RECT 185.400 177.900 186.600 178.950 ;
        RECT 184.950 175.800 187.050 177.900 ;
        RECT 191.400 177.000 192.600 178.950 ;
        RECT 190.950 172.950 193.050 177.000 ;
        RECT 197.400 175.050 198.600 202.950 ;
        RECT 200.400 175.050 201.600 247.950 ;
        RECT 206.400 238.050 207.600 247.950 ;
        RECT 205.950 235.950 208.050 238.050 ;
        RECT 206.400 214.050 207.600 235.950 ;
        RECT 223.950 225.300 226.050 227.400 ;
        RECT 239.400 226.050 240.600 268.950 ;
        RECT 241.950 256.950 244.050 259.050 ;
        RECT 242.400 244.050 243.600 256.950 ;
        RECT 241.950 241.950 244.050 244.050 ;
        RECT 245.400 241.050 246.600 280.950 ;
        RECT 250.950 280.500 253.050 282.600 ;
        RECT 250.950 274.950 253.050 277.050 ;
        RECT 251.400 259.050 252.600 274.950 ;
        RECT 257.400 268.050 258.600 286.950 ;
        RECT 260.400 283.050 261.600 332.400 ;
        RECT 266.400 331.050 267.600 373.950 ;
        RECT 269.400 358.050 270.600 412.950 ;
        RECT 275.100 402.600 276.300 422.400 ;
        RECT 277.950 412.950 280.050 415.050 ;
        RECT 278.400 411.600 279.600 412.950 ;
        RECT 277.950 409.500 280.050 411.600 ;
        RECT 274.950 400.500 277.050 402.600 ;
        RECT 277.950 391.950 280.050 394.050 ;
        RECT 278.400 379.050 279.600 391.950 ;
        RECT 284.400 385.050 285.600 442.950 ;
        RECT 286.950 439.950 289.050 444.000 ;
        RECT 290.850 438.600 292.050 453.600 ;
        RECT 295.950 449.100 298.050 451.200 ;
        RECT 289.950 436.500 292.050 438.600 ;
        RECT 296.400 433.050 297.600 449.100 ;
        RECT 299.400 439.050 300.600 472.950 ;
        RECT 305.400 472.050 306.600 478.950 ;
        RECT 308.400 475.050 309.600 521.400 ;
        RECT 311.400 478.050 312.600 523.950 ;
        RECT 317.400 517.050 318.600 523.950 ;
        RECT 323.400 522.600 324.600 523.950 ;
        RECT 320.400 521.400 324.600 522.600 ;
        RECT 316.950 514.950 319.050 517.050 ;
        RECT 317.400 493.050 318.600 514.950 ;
        RECT 320.400 508.050 321.600 521.400 ;
        RECT 326.850 516.600 328.050 531.600 ;
        RECT 331.950 523.950 334.050 526.050 ;
        RECT 325.950 514.500 328.050 516.600 ;
        RECT 319.950 505.950 322.050 508.050 ;
        RECT 328.950 505.950 331.050 508.050 ;
        RECT 322.950 495.000 325.050 499.050 ;
        RECT 329.400 496.050 330.600 505.950 ;
        RECT 332.400 502.050 333.600 523.950 ;
        RECT 331.950 499.950 334.050 502.050 ;
        RECT 331.950 496.800 334.050 498.900 ;
        RECT 323.400 493.050 324.600 495.000 ;
        RECT 328.950 493.950 331.050 496.050 ;
        RECT 316.950 490.950 319.050 493.050 ;
        RECT 319.950 490.950 322.050 493.050 ;
        RECT 322.950 490.950 325.050 493.050 ;
        RECT 325.950 490.950 328.050 493.050 ;
        RECT 316.950 484.950 319.050 487.050 ;
        RECT 310.950 475.950 313.050 478.050 ;
        RECT 307.950 472.950 310.050 475.050 ;
        RECT 304.950 469.950 307.050 472.050 ;
        RECT 301.950 466.950 304.050 469.050 ;
        RECT 302.400 457.050 303.600 466.950 ;
        RECT 317.400 466.050 318.600 484.950 ;
        RECT 320.400 478.050 321.600 490.950 ;
        RECT 326.400 490.050 327.600 490.950 ;
        RECT 326.400 488.400 331.050 490.050 ;
        RECT 327.000 487.950 331.050 488.400 ;
        RECT 332.400 487.050 333.600 496.800 ;
        RECT 331.950 484.950 334.050 487.050 ;
        RECT 319.950 475.950 322.050 478.050 ;
        RECT 325.950 475.950 328.050 478.050 ;
        RECT 316.950 463.950 319.050 466.050 ;
        RECT 310.950 458.400 313.050 460.500 ;
        RECT 301.950 454.950 304.050 457.050 ;
        RECT 304.950 449.400 307.050 451.500 ;
        RECT 305.400 448.050 306.600 449.400 ;
        RECT 304.950 445.950 307.050 448.050 ;
        RECT 298.950 436.950 301.050 439.050 ;
        RECT 311.100 438.600 312.300 458.400 ;
        RECT 317.400 450.600 318.600 463.950 ;
        RECT 319.950 460.950 322.050 463.050 ;
        RECT 314.400 449.400 318.600 450.600 ;
        RECT 314.400 448.050 315.600 449.400 ;
        RECT 313.950 445.950 316.050 448.050 ;
        RECT 316.950 442.950 319.050 445.050 ;
        RECT 310.950 436.500 313.050 438.600 ;
        RECT 295.950 430.950 298.050 433.050 ;
        RECT 317.400 432.600 318.600 442.950 ;
        RECT 320.400 436.050 321.600 460.950 ;
        RECT 319.950 433.950 322.050 436.050 ;
        RECT 317.400 431.400 321.600 432.600 ;
        RECT 295.950 427.800 298.050 429.900 ;
        RECT 296.400 415.050 297.600 427.800 ;
        RECT 304.950 421.950 307.050 424.050 ;
        RECT 292.950 412.950 295.050 415.050 ;
        RECT 295.950 412.950 298.050 415.050 ;
        RECT 298.950 412.950 301.050 415.050 ;
        RECT 293.400 394.050 294.600 412.950 ;
        RECT 299.400 403.050 300.600 412.950 ;
        RECT 305.400 411.900 306.600 421.950 ;
        RECT 307.950 416.100 310.050 418.200 ;
        RECT 313.950 416.100 316.050 418.200 ;
        RECT 304.950 409.800 307.050 411.900 ;
        RECT 298.950 400.950 301.050 403.050 ;
        RECT 292.950 391.950 295.050 394.050 ;
        RECT 283.950 382.950 286.050 385.050 ;
        RECT 277.950 376.950 280.050 379.050 ;
        RECT 271.950 371.100 274.050 373.200 ;
        RECT 272.400 367.050 273.600 371.100 ;
        RECT 278.400 370.050 279.600 376.950 ;
        RECT 284.400 371.400 291.600 372.600 ;
        RECT 298.950 372.000 301.050 376.050 ;
        RECT 284.400 370.050 285.600 371.400 ;
        RECT 277.950 367.950 280.050 370.050 ;
        RECT 280.950 367.950 283.050 370.050 ;
        RECT 283.950 367.950 286.050 370.050 ;
        RECT 271.950 364.950 274.050 367.050 ;
        RECT 281.400 366.900 282.600 367.950 ;
        RECT 280.950 364.800 283.050 366.900 ;
        RECT 290.400 358.050 291.600 371.400 ;
        RECT 299.400 370.050 300.600 372.000 ;
        RECT 298.950 367.950 301.050 370.050 ;
        RECT 301.950 367.950 304.050 370.050 ;
        RECT 302.400 366.000 303.600 367.950 ;
        RECT 301.950 361.950 304.050 366.000 ;
        RECT 268.950 355.950 271.050 358.050 ;
        RECT 289.950 355.950 292.050 358.050 ;
        RECT 308.400 352.050 309.600 416.100 ;
        RECT 314.400 415.050 315.600 416.100 ;
        RECT 320.400 415.050 321.600 431.400 ;
        RECT 326.400 417.600 327.600 475.950 ;
        RECT 331.950 457.950 334.050 460.050 ;
        RECT 332.400 448.050 333.600 457.950 ;
        RECT 335.400 454.050 336.600 535.950 ;
        RECT 340.950 527.400 343.050 529.500 ;
        RECT 341.400 526.050 342.600 527.400 ;
        RECT 340.950 523.950 343.050 526.050 ;
        RECT 337.950 520.950 340.050 523.050 ;
        RECT 338.400 511.050 339.600 520.950 ;
        RECT 347.100 516.600 348.300 536.400 ;
        RECT 349.950 532.950 352.050 535.050 ;
        RECT 350.400 526.050 351.600 532.950 ;
        RECT 349.950 523.950 352.050 526.050 ;
        RECT 346.950 514.500 349.050 516.600 ;
        RECT 352.950 514.950 355.050 517.050 ;
        RECT 337.950 508.950 340.050 511.050 ;
        RECT 346.950 508.950 349.050 511.050 ;
        RECT 337.950 499.950 340.050 502.050 ;
        RECT 338.400 493.050 339.600 499.950 ;
        RECT 347.400 493.050 348.600 508.950 ;
        RECT 353.400 502.050 354.600 514.950 ;
        RECT 352.950 499.950 355.050 502.050 ;
        RECT 356.400 498.600 357.600 559.950 ;
        RECT 368.400 556.050 369.600 572.400 ;
        RECT 373.950 568.950 376.050 571.050 ;
        RECT 367.950 553.950 370.050 556.050 ;
        RECT 374.400 538.050 375.600 568.950 ;
        RECT 386.400 562.050 387.600 583.950 ;
        RECT 389.400 574.050 390.600 589.950 ;
        RECT 388.950 571.950 391.050 574.050 ;
        RECT 394.950 572.100 397.050 574.200 ;
        RECT 395.400 571.050 396.600 572.100 ;
        RECT 391.950 568.950 394.050 571.050 ;
        RECT 394.950 568.950 397.050 571.050 ;
        RECT 392.400 562.050 393.600 568.950 ;
        RECT 401.400 567.600 402.600 650.100 ;
        RECT 410.400 649.050 411.600 670.950 ;
        RECT 416.400 652.050 417.600 676.950 ;
        RECT 419.400 676.050 420.600 712.950 ;
        RECT 422.400 712.050 423.600 722.400 ;
        RECT 425.400 721.050 426.600 761.100 ;
        RECT 428.400 742.050 429.600 761.400 ;
        RECT 436.950 761.100 439.050 763.200 ;
        RECT 442.950 761.100 445.050 763.200 ;
        RECT 437.400 760.050 438.600 761.100 ;
        RECT 443.400 760.050 444.600 761.100 ;
        RECT 461.400 760.050 462.600 775.950 ;
        RECT 469.950 766.950 472.050 769.050 ;
        RECT 433.950 757.950 436.050 760.050 ;
        RECT 436.950 757.950 439.050 760.050 ;
        RECT 439.950 757.950 442.050 760.050 ;
        RECT 442.950 757.950 445.050 760.050 ;
        RECT 445.950 757.950 448.050 760.050 ;
        RECT 457.950 757.950 460.050 760.050 ;
        RECT 460.950 757.950 463.050 760.050 ;
        RECT 463.950 757.950 466.050 760.050 ;
        RECT 434.400 756.900 435.600 757.950 ;
        RECT 433.950 754.800 436.050 756.900 ;
        RECT 440.400 742.050 441.600 757.950 ;
        RECT 446.400 748.050 447.600 757.950 ;
        RECT 451.950 754.800 454.050 756.900 ;
        RECT 445.950 745.950 448.050 748.050 ;
        RECT 427.950 739.950 430.050 742.050 ;
        RECT 439.950 739.950 442.050 742.050 ;
        RECT 436.950 724.950 439.050 727.050 ;
        RECT 424.950 718.950 427.050 721.050 ;
        RECT 433.950 718.950 436.050 721.050 ;
        RECT 421.950 709.950 424.050 712.050 ;
        RECT 422.400 697.050 423.600 709.950 ;
        RECT 427.950 697.950 430.050 700.050 ;
        RECT 421.950 694.950 424.050 697.050 ;
        RECT 421.950 691.800 424.050 693.900 ;
        RECT 418.950 673.950 421.050 676.050 ;
        RECT 422.400 667.050 423.600 691.800 ;
        RECT 428.400 682.050 429.600 697.950 ;
        RECT 434.400 682.050 435.600 718.950 ;
        RECT 437.400 712.050 438.600 724.950 ;
        RECT 436.950 709.950 439.050 712.050 ;
        RECT 452.400 709.050 453.600 754.800 ;
        RECT 458.400 748.050 459.600 757.950 ;
        RECT 464.400 756.900 465.600 757.950 ;
        RECT 463.950 754.800 466.050 756.900 ;
        RECT 457.950 745.950 460.050 748.050 ;
        RECT 460.950 733.950 463.050 736.050 ;
        RECT 461.400 727.050 462.600 733.950 ;
        RECT 466.950 729.600 469.050 730.200 ;
        RECT 470.400 729.600 471.600 766.950 ;
        RECT 473.400 742.050 474.600 775.950 ;
        RECT 493.950 766.950 496.050 769.050 ;
        RECT 505.950 766.950 508.050 769.050 ;
        RECT 481.950 762.000 484.050 766.050 ;
        RECT 482.400 760.050 483.600 762.000 ;
        RECT 487.950 761.100 490.050 763.200 ;
        RECT 488.400 760.050 489.600 761.100 ;
        RECT 478.950 757.950 481.050 760.050 ;
        RECT 481.950 757.950 484.050 760.050 ;
        RECT 484.950 757.950 487.050 760.050 ;
        RECT 487.950 757.950 490.050 760.050 ;
        RECT 479.400 751.050 480.600 757.950 ;
        RECT 485.400 756.900 486.600 757.950 ;
        RECT 494.400 757.050 495.600 766.950 ;
        RECT 499.950 763.950 502.050 766.050 ;
        RECT 496.950 761.100 499.050 763.200 ;
        RECT 484.950 754.800 487.050 756.900 ;
        RECT 490.950 755.400 495.600 757.050 ;
        RECT 490.950 754.950 495.000 755.400 ;
        RECT 478.950 748.950 481.050 751.050 ;
        RECT 493.950 748.950 496.050 751.050 ;
        RECT 475.950 742.950 478.050 745.050 ;
        RECT 472.950 739.950 475.050 742.050 ;
        RECT 472.950 733.950 475.050 736.050 ;
        RECT 466.950 728.400 471.600 729.600 ;
        RECT 466.950 728.100 469.050 728.400 ;
        RECT 467.400 727.050 468.600 728.100 ;
        RECT 457.950 724.950 460.050 727.050 ;
        RECT 460.950 724.950 463.050 727.050 ;
        RECT 463.950 724.950 466.050 727.050 ;
        RECT 466.950 724.950 469.050 727.050 ;
        RECT 451.950 706.950 454.050 709.050 ;
        RECT 458.400 697.050 459.600 724.950 ;
        RECT 464.400 715.050 465.600 724.950 ;
        RECT 469.950 721.800 472.050 723.900 ;
        RECT 463.950 712.950 466.050 715.050 ;
        RECT 448.950 694.950 451.050 697.050 ;
        RECT 457.950 694.950 460.050 697.050 ;
        RECT 439.950 683.100 442.050 685.200 ;
        RECT 445.950 683.100 448.050 685.200 ;
        RECT 440.400 682.050 441.600 683.100 ;
        RECT 427.950 679.950 430.050 682.050 ;
        RECT 430.950 679.950 433.050 682.050 ;
        RECT 433.950 679.950 436.050 682.050 ;
        RECT 436.950 679.950 439.050 682.050 ;
        RECT 439.950 679.950 442.050 682.050 ;
        RECT 427.950 672.600 430.050 676.050 ;
        RECT 431.400 675.600 432.600 679.950 ;
        RECT 437.400 678.900 438.600 679.950 ;
        RECT 436.950 676.800 439.050 678.900 ;
        RECT 446.400 678.600 447.600 683.100 ;
        RECT 449.400 679.050 450.600 694.950 ;
        RECT 457.950 684.000 460.050 688.050 ;
        RECT 458.400 682.050 459.600 684.000 ;
        RECT 463.950 683.100 466.050 685.200 ;
        RECT 464.400 682.050 465.600 683.100 ;
        RECT 454.950 679.950 457.050 682.050 ;
        RECT 457.950 679.950 460.050 682.050 ;
        RECT 460.950 679.950 463.050 682.050 ;
        RECT 463.950 679.950 466.050 682.050 ;
        RECT 443.400 677.400 447.600 678.600 ;
        RECT 431.400 674.400 435.600 675.600 ;
        RECT 427.950 672.000 432.600 672.600 ;
        RECT 428.400 671.400 432.600 672.000 ;
        RECT 424.950 667.800 427.050 669.900 ;
        RECT 421.950 664.950 424.050 667.050 ;
        RECT 421.950 652.950 424.050 655.050 ;
        RECT 415.950 649.950 418.050 652.050 ;
        RECT 406.950 646.950 409.050 649.050 ;
        RECT 409.950 646.950 412.050 649.050 ;
        RECT 412.950 646.950 415.050 649.050 ;
        RECT 403.950 643.800 406.050 645.900 ;
        RECT 404.400 586.050 405.600 643.800 ;
        RECT 407.400 640.050 408.600 646.950 ;
        RECT 413.400 645.900 414.600 646.950 ;
        RECT 412.950 643.800 415.050 645.900 ;
        RECT 415.950 643.950 418.050 646.050 ;
        RECT 422.400 645.900 423.600 652.950 ;
        RECT 425.400 652.050 426.600 667.800 ;
        RECT 424.950 649.950 427.050 652.050 ;
        RECT 431.400 649.050 432.600 671.400 ;
        RECT 434.400 655.050 435.600 674.400 ;
        RECT 439.950 673.950 442.050 676.050 ;
        RECT 433.950 652.950 436.050 655.050 ;
        RECT 427.950 646.950 430.050 649.050 ;
        RECT 430.950 646.950 433.050 649.050 ;
        RECT 433.950 646.950 436.050 649.050 ;
        RECT 428.400 645.900 429.600 646.950 ;
        RECT 406.950 637.950 409.050 640.050 ;
        RECT 407.400 622.050 408.600 637.950 ;
        RECT 416.400 637.050 417.600 643.950 ;
        RECT 421.950 643.800 424.050 645.900 ;
        RECT 427.950 643.800 430.050 645.900 ;
        RECT 434.400 645.000 435.600 646.950 ;
        RECT 409.950 634.950 412.050 637.050 ;
        RECT 412.950 634.950 415.050 637.050 ;
        RECT 415.950 634.950 418.050 637.050 ;
        RECT 406.950 619.950 409.050 622.050 ;
        RECT 410.400 604.050 411.600 634.950 ;
        RECT 413.400 625.050 414.600 634.950 ;
        RECT 412.950 622.950 415.050 625.050 ;
        RECT 422.400 613.050 423.600 643.800 ;
        RECT 433.950 640.950 436.050 645.000 ;
        RECT 440.400 639.600 441.600 673.950 ;
        RECT 443.400 643.050 444.600 677.400 ;
        RECT 448.950 676.950 451.050 679.050 ;
        RECT 455.400 678.000 456.600 679.950 ;
        RECT 461.400 678.900 462.600 679.950 ;
        RECT 454.950 673.950 457.050 678.000 ;
        RECT 460.950 676.800 463.050 678.900 ;
        RECT 466.950 678.600 469.050 679.050 ;
        RECT 470.400 678.600 471.600 721.800 ;
        RECT 473.400 715.050 474.600 733.950 ;
        RECT 476.400 718.050 477.600 742.950 ;
        RECT 478.950 739.950 481.050 742.050 ;
        RECT 479.400 730.200 480.600 739.950 ;
        RECT 478.950 728.100 481.050 730.200 ;
        RECT 484.950 728.100 487.050 730.200 ;
        RECT 490.950 728.100 493.050 730.200 ;
        RECT 485.400 727.050 486.600 728.100 ;
        RECT 481.950 724.950 484.050 727.050 ;
        RECT 484.950 724.950 487.050 727.050 ;
        RECT 482.400 723.900 483.600 724.950 ;
        RECT 481.950 721.800 484.050 723.900 ;
        RECT 475.950 715.950 478.050 718.050 ;
        RECT 472.950 712.950 475.050 715.050 ;
        RECT 472.950 706.950 475.050 709.050 ;
        RECT 473.400 697.050 474.600 706.950 ;
        RECT 491.400 706.050 492.600 728.100 ;
        RECT 494.400 723.600 495.600 748.950 ;
        RECT 497.400 733.050 498.600 761.100 ;
        RECT 500.400 756.600 501.600 763.950 ;
        RECT 506.400 760.050 507.600 766.950 ;
        RECT 511.950 762.000 514.050 766.050 ;
        RECT 512.400 760.050 513.600 762.000 ;
        RECT 505.950 757.950 508.050 760.050 ;
        RECT 508.950 757.950 511.050 760.050 ;
        RECT 511.950 757.950 514.050 760.050 ;
        RECT 514.950 757.950 517.050 760.050 ;
        RECT 500.400 755.400 504.600 756.600 ;
        RECT 496.950 730.950 499.050 733.050 ;
        RECT 503.400 727.050 504.600 755.400 ;
        RECT 509.400 751.050 510.600 757.950 ;
        RECT 515.400 756.900 516.600 757.950 ;
        RECT 521.400 757.050 522.600 794.400 ;
        RECT 551.400 790.050 552.600 802.950 ;
        RECT 557.400 801.900 558.600 802.950 ;
        RECT 556.950 799.800 559.050 801.900 ;
        RECT 550.950 787.950 553.050 790.050 ;
        RECT 556.950 787.950 559.050 790.050 ;
        RECT 557.400 784.050 558.600 787.950 ;
        RECT 566.400 787.050 567.600 806.400 ;
        RECT 572.400 790.050 573.600 823.950 ;
        RECT 580.950 817.950 583.050 820.050 ;
        RECT 581.400 805.050 582.600 817.950 ;
        RECT 604.950 814.950 607.050 817.050 ;
        RECT 586.950 806.100 589.050 808.200 ;
        RECT 598.950 806.100 601.050 808.200 ;
        RECT 587.400 805.050 588.600 806.100 ;
        RECT 599.400 805.050 600.600 806.100 ;
        RECT 605.400 805.050 606.600 814.950 ;
        RECT 622.950 808.950 625.050 811.050 ;
        RECT 613.950 806.100 616.050 808.200 ;
        RECT 577.950 802.950 580.050 805.050 ;
        RECT 580.950 802.950 583.050 805.050 ;
        RECT 583.950 802.950 586.050 805.050 ;
        RECT 586.950 802.950 589.050 805.050 ;
        RECT 598.950 802.950 601.050 805.050 ;
        RECT 601.950 802.950 604.050 805.050 ;
        RECT 604.950 802.950 607.050 805.050 ;
        RECT 607.950 802.950 610.050 805.050 ;
        RECT 578.400 790.050 579.600 802.950 ;
        RECT 584.400 801.900 585.600 802.950 ;
        RECT 602.400 801.900 603.600 802.950 ;
        RECT 608.400 801.900 609.600 802.950 ;
        RECT 583.950 799.800 586.050 801.900 ;
        RECT 601.950 799.800 604.050 801.900 ;
        RECT 607.950 799.800 610.050 801.900 ;
        RECT 571.950 787.950 574.050 790.050 ;
        RECT 577.950 787.950 580.050 790.050 ;
        RECT 559.950 784.950 562.050 787.050 ;
        RECT 565.950 784.950 568.050 787.050 ;
        RECT 526.950 781.950 529.050 784.050 ;
        RECT 556.950 781.950 559.050 784.050 ;
        RECT 523.950 760.950 526.050 763.050 ;
        RECT 514.950 754.800 517.050 756.900 ;
        RECT 520.950 754.950 523.050 757.050 ;
        RECT 524.400 751.050 525.600 760.950 ;
        RECT 508.950 748.950 511.050 751.050 ;
        RECT 523.950 748.950 526.050 751.050 ;
        RECT 520.950 739.950 523.050 742.050 ;
        RECT 511.950 727.950 514.050 730.050 ;
        RECT 499.950 724.950 502.050 727.050 ;
        RECT 502.950 724.950 505.050 727.050 ;
        RECT 505.950 724.950 508.050 727.050 ;
        RECT 494.400 722.400 498.600 723.600 ;
        RECT 493.950 715.950 496.050 718.050 ;
        RECT 490.950 703.950 493.050 706.050 ;
        RECT 472.950 694.950 475.050 697.050 ;
        RECT 466.950 677.400 471.600 678.600 ;
        RECT 466.950 676.950 469.050 677.400 ;
        RECT 467.400 673.050 468.600 676.950 ;
        RECT 473.400 676.050 474.600 694.950 ;
        RECT 481.950 684.000 484.050 688.050 ;
        RECT 482.400 682.050 483.600 684.000 ;
        RECT 487.950 683.100 490.050 685.200 ;
        RECT 488.400 682.050 489.600 683.100 ;
        RECT 490.950 682.950 493.050 688.050 ;
        RECT 478.950 679.950 481.050 682.050 ;
        RECT 481.950 679.950 484.050 682.050 ;
        RECT 484.950 679.950 487.050 682.050 ;
        RECT 487.950 679.950 490.050 682.050 ;
        RECT 479.400 679.050 480.600 679.950 ;
        RECT 475.950 677.400 480.600 679.050 ;
        RECT 485.400 678.900 486.600 679.950 ;
        RECT 494.400 679.050 495.600 715.950 ;
        RECT 475.950 676.950 480.000 677.400 ;
        RECT 484.950 676.800 487.050 678.900 ;
        RECT 493.950 676.950 496.050 679.050 ;
        RECT 469.800 673.800 471.900 675.900 ;
        RECT 472.950 673.950 475.050 676.050 ;
        RECT 478.950 673.950 481.050 676.050 ;
        RECT 466.950 670.950 469.050 673.050 ;
        RECT 457.950 667.950 460.050 670.050 ;
        RECT 454.950 661.950 457.050 664.050 ;
        RECT 445.950 655.950 448.050 658.050 ;
        RECT 446.400 643.050 447.600 655.950 ;
        RECT 455.400 649.050 456.600 661.950 ;
        RECT 458.400 655.050 459.600 667.950 ;
        RECT 463.950 661.950 466.050 664.050 ;
        RECT 457.800 652.950 459.900 655.050 ;
        RECT 460.950 651.000 463.050 655.050 ;
        RECT 464.400 652.050 465.600 661.950 ;
        RECT 461.400 649.050 462.600 651.000 ;
        RECT 463.950 649.950 466.050 652.050 ;
        RECT 451.950 646.950 454.050 649.050 ;
        RECT 454.950 646.950 457.050 649.050 ;
        RECT 457.950 646.950 460.050 649.050 ;
        RECT 460.950 646.950 463.050 649.050 ;
        RECT 452.400 645.900 453.600 646.950 ;
        RECT 458.400 645.900 459.600 646.950 ;
        RECT 451.950 643.800 454.050 645.900 ;
        RECT 457.950 643.800 460.050 645.900 ;
        RECT 463.950 643.800 466.050 645.900 ;
        RECT 442.950 640.950 445.050 643.050 ;
        RECT 445.950 640.950 448.050 643.050 ;
        RECT 440.400 638.400 444.600 639.600 ;
        RECT 427.950 634.950 430.050 637.050 ;
        RECT 424.950 628.950 427.050 631.050 ;
        RECT 425.400 622.050 426.600 628.950 ;
        RECT 428.400 628.050 429.600 634.950 ;
        RECT 436.950 628.950 439.050 631.050 ;
        RECT 427.950 625.950 430.050 628.050 ;
        RECT 437.400 625.050 438.600 628.950 ;
        RECT 436.950 622.950 439.050 625.050 ;
        RECT 424.950 619.950 427.050 622.050 ;
        RECT 433.950 619.950 436.050 622.050 ;
        RECT 434.400 616.050 435.600 619.950 ;
        RECT 424.950 613.950 427.050 616.050 ;
        RECT 433.950 613.950 436.050 616.050 ;
        RECT 421.950 610.950 424.050 613.050 ;
        RECT 409.950 601.950 412.050 604.050 ;
        RECT 412.950 601.950 415.050 604.050 ;
        RECT 413.400 600.900 414.600 601.950 ;
        RECT 412.950 598.800 415.050 600.900 ;
        RECT 403.950 583.950 406.050 586.050 ;
        RECT 425.400 574.200 426.600 613.950 ;
        RECT 430.950 610.950 433.050 613.050 ;
        RECT 431.400 604.050 432.600 610.950 ;
        RECT 430.950 601.950 433.050 604.050 ;
        RECT 443.400 600.600 444.600 638.400 ;
        RECT 464.400 637.050 465.600 643.800 ;
        RECT 467.400 640.050 468.600 670.950 ;
        RECT 470.400 664.050 471.600 673.800 ;
        RECT 469.950 661.950 472.050 664.050 ;
        RECT 469.950 649.950 472.050 652.050 ;
        RECT 466.950 637.950 469.050 640.050 ;
        RECT 463.950 634.950 466.050 637.050 ;
        RECT 451.950 616.950 454.050 619.050 ;
        RECT 452.400 607.200 453.600 616.950 ;
        RECT 451.950 605.100 454.050 607.200 ;
        RECT 452.400 604.050 453.600 605.100 ;
        RECT 451.950 601.950 454.050 604.050 ;
        RECT 464.400 600.600 465.600 634.950 ;
        RECT 470.400 628.050 471.600 649.950 ;
        RECT 479.400 649.050 480.600 673.950 ;
        RECT 487.950 670.950 490.050 673.050 ;
        RECT 484.950 667.950 487.050 670.050 ;
        RECT 485.400 652.050 486.600 667.950 ;
        RECT 484.950 649.950 487.050 652.050 ;
        RECT 475.950 646.950 478.050 649.050 ;
        RECT 478.950 646.950 481.050 649.050 ;
        RECT 481.950 646.950 484.050 649.050 ;
        RECT 476.400 645.900 477.600 646.950 ;
        RECT 475.950 643.800 478.050 645.900 ;
        RECT 469.950 625.950 472.050 628.050 ;
        RECT 476.400 619.050 477.600 643.800 ;
        RECT 482.400 643.050 483.600 646.950 ;
        RECT 481.950 640.950 484.050 643.050 ;
        RECT 478.950 637.950 481.050 640.050 ;
        RECT 475.950 616.950 478.050 619.050 ;
        RECT 472.950 605.100 475.050 607.200 ;
        RECT 473.400 604.050 474.600 605.100 ;
        RECT 479.400 604.050 480.600 637.950 ;
        RECT 482.400 634.050 483.600 640.950 ;
        RECT 481.950 631.950 484.050 634.050 ;
        RECT 488.400 631.050 489.600 670.950 ;
        RECT 497.400 655.050 498.600 722.400 ;
        RECT 500.400 685.050 501.600 724.950 ;
        RECT 506.400 703.050 507.600 724.950 ;
        RECT 505.950 700.950 508.050 703.050 ;
        RECT 499.950 682.950 502.050 685.050 ;
        RECT 505.950 683.100 508.050 685.200 ;
        RECT 512.400 685.050 513.600 727.950 ;
        RECT 521.400 727.050 522.600 739.950 ;
        RECT 527.400 730.050 528.600 781.950 ;
        RECT 550.950 775.950 553.050 778.050 ;
        RECT 551.400 771.600 552.600 775.950 ;
        RECT 556.950 771.600 559.050 772.050 ;
        RECT 551.400 770.400 559.050 771.600 ;
        RECT 556.950 769.950 559.050 770.400 ;
        RECT 553.950 766.950 556.050 769.050 ;
        RECT 532.950 761.100 535.050 763.200 ;
        RECT 541.950 761.100 544.050 763.200 ;
        RECT 547.950 761.100 550.050 763.200 ;
        RECT 533.400 760.050 534.600 761.100 ;
        RECT 532.950 757.950 535.050 760.050 ;
        RECT 535.950 757.950 538.050 760.050 ;
        RECT 529.950 754.950 532.050 757.050 ;
        RECT 526.950 727.950 529.050 730.050 ;
        RECT 517.950 724.950 520.050 727.050 ;
        RECT 520.950 724.950 523.050 727.050 ;
        RECT 518.400 715.050 519.600 724.950 ;
        RECT 517.950 712.950 520.050 715.050 ;
        RECT 520.950 709.950 523.050 712.050 ;
        RECT 514.950 691.950 517.050 694.050 ;
        RECT 506.400 682.050 507.600 683.100 ;
        RECT 511.950 682.950 514.050 685.050 ;
        RECT 515.400 682.050 516.600 691.950 ;
        RECT 499.950 679.800 502.050 681.900 ;
        RECT 505.950 679.950 508.050 682.050 ;
        RECT 514.950 679.950 517.050 682.050 ;
        RECT 500.400 673.050 501.600 679.800 ;
        RECT 521.400 678.600 522.600 709.950 ;
        RECT 530.400 687.600 531.600 754.950 ;
        RECT 536.400 751.050 537.600 757.950 ;
        RECT 542.400 751.050 543.600 761.100 ;
        RECT 548.400 760.050 549.600 761.100 ;
        RECT 554.400 760.050 555.600 766.950 ;
        RECT 560.400 763.050 561.600 784.950 ;
        RECT 571.950 778.950 574.050 781.050 ;
        RECT 562.950 766.950 565.050 769.050 ;
        RECT 559.950 760.950 562.050 763.050 ;
        RECT 547.950 757.950 550.050 760.050 ;
        RECT 550.950 757.950 553.050 760.050 ;
        RECT 553.950 757.950 556.050 760.050 ;
        RECT 556.950 757.950 559.050 760.050 ;
        RECT 535.950 748.950 538.050 751.050 ;
        RECT 541.950 748.950 544.050 751.050 ;
        RECT 551.400 745.050 552.600 757.950 ;
        RECT 557.400 756.900 558.600 757.950 ;
        RECT 563.400 757.050 564.600 766.950 ;
        RECT 565.950 761.100 568.050 763.200 ;
        RECT 572.400 763.050 573.600 778.950 ;
        RECT 578.400 772.050 579.600 787.950 ;
        RECT 602.400 784.050 603.600 799.800 ;
        RECT 601.950 781.950 604.050 784.050 ;
        RECT 614.400 781.050 615.600 806.100 ;
        RECT 623.400 793.050 624.600 808.950 ;
        RECT 629.400 805.050 630.600 826.950 ;
        RECT 632.400 811.050 633.600 835.950 ;
        RECT 631.950 808.950 634.050 811.050 ;
        RECT 634.950 806.100 637.050 808.200 ;
        RECT 641.400 808.050 642.600 841.950 ;
        RECT 650.400 840.600 651.600 877.800 ;
        RECT 658.950 874.950 661.050 879.000 ;
        RECT 664.950 877.800 667.050 879.900 ;
        RECT 670.950 877.800 673.050 879.900 ;
        RECT 676.950 877.800 679.050 879.900 ;
        RECT 682.950 877.800 685.050 879.900 ;
        RECT 683.400 874.050 684.600 877.800 ;
        RECT 682.950 871.950 685.050 874.050 ;
        RECT 689.400 871.050 690.600 892.950 ;
        RECT 706.950 889.050 709.050 889.200 ;
        RECT 703.950 887.100 709.050 889.050 ;
        RECT 721.950 888.600 726.000 889.050 ;
        RECT 703.950 886.950 708.000 887.100 ;
        RECT 721.950 886.950 726.600 888.600 ;
        RECT 700.950 884.100 703.050 886.200 ;
        RECT 701.400 883.050 702.600 884.100 ;
        RECT 706.950 883.950 709.050 886.050 ;
        RECT 707.400 883.050 708.600 883.950 ;
        RECT 725.400 883.050 726.600 886.950 ;
        RECT 730.950 884.100 733.050 886.200 ;
        RECT 731.400 883.050 732.600 884.100 ;
        RECT 739.950 883.950 742.050 886.050 ;
        RECT 748.950 884.100 751.050 886.200 ;
        RECT 754.950 884.100 757.050 886.200 ;
        RECT 763.950 884.100 766.050 886.200 ;
        RECT 772.950 884.100 775.050 886.200 ;
        RECT 700.950 880.950 703.050 883.050 ;
        RECT 703.950 880.950 706.050 883.050 ;
        RECT 706.950 880.950 709.050 883.050 ;
        RECT 709.950 880.950 712.050 883.050 ;
        RECT 724.950 880.950 727.050 883.050 ;
        RECT 727.950 880.950 730.050 883.050 ;
        RECT 730.950 880.950 733.050 883.050 ;
        RECT 733.950 880.950 736.050 883.050 ;
        RECT 704.400 879.000 705.600 880.950 ;
        RECT 710.400 879.900 711.600 880.950 ;
        RECT 728.400 879.900 729.600 880.950 ;
        RECT 703.950 874.950 706.050 879.000 ;
        RECT 709.950 877.800 712.050 879.900 ;
        RECT 727.950 877.800 730.050 879.900 ;
        RECT 734.400 879.000 735.600 880.950 ;
        RECT 688.950 868.950 691.050 871.050 ;
        RECT 658.950 859.950 661.050 862.050 ;
        RECT 685.950 859.950 688.050 862.050 ;
        RECT 650.400 839.400 654.600 840.600 ;
        RECT 653.400 838.050 654.600 839.400 ;
        RECT 659.400 838.050 660.600 859.950 ;
        RECT 686.400 844.050 687.600 859.950 ;
        RECT 664.950 841.950 667.050 844.050 ;
        RECT 667.950 841.950 670.050 844.050 ;
        RECT 665.400 838.050 666.600 841.950 ;
        RECT 652.950 835.950 655.050 838.050 ;
        RECT 655.950 835.950 658.050 838.050 ;
        RECT 658.950 835.950 661.050 838.050 ;
        RECT 664.950 835.950 667.050 838.050 ;
        RECT 656.400 834.900 657.600 835.950 ;
        RECT 668.400 835.050 669.600 841.950 ;
        RECT 673.950 840.000 676.050 844.050 ;
        RECT 685.950 841.950 688.050 844.050 ;
        RECT 674.400 838.050 675.600 840.000 ;
        RECT 679.950 839.100 682.050 841.200 ;
        RECT 680.400 838.050 681.600 839.100 ;
        RECT 673.950 835.950 676.050 838.050 ;
        RECT 676.950 835.950 679.050 838.050 ;
        RECT 679.950 835.950 682.050 838.050 ;
        RECT 655.950 832.800 658.050 834.900 ;
        RECT 667.950 832.950 670.050 835.050 ;
        RECT 677.400 834.900 678.600 835.950 ;
        RECT 686.400 835.050 687.600 841.950 ;
        RECT 691.950 840.000 694.050 844.050 ;
        RECT 692.400 838.050 693.600 840.000 ;
        RECT 697.950 839.100 700.050 841.200 ;
        RECT 698.400 838.050 699.600 839.100 ;
        RECT 691.950 835.950 694.050 838.050 ;
        RECT 694.950 835.950 697.050 838.050 ;
        RECT 697.950 835.950 700.050 838.050 ;
        RECT 676.950 832.800 679.050 834.900 ;
        RECT 685.950 832.950 688.050 835.050 ;
        RECT 695.400 826.050 696.600 835.950 ;
        RECT 694.950 823.950 697.050 826.050 ;
        RECT 697.950 820.950 700.050 823.050 ;
        RECT 652.950 811.950 655.050 814.050 ;
        RECT 653.400 808.200 654.600 811.950 ;
        RECT 635.400 805.050 636.600 806.100 ;
        RECT 640.950 805.950 643.050 808.050 ;
        RECT 643.950 806.100 646.050 808.200 ;
        RECT 652.950 806.100 655.050 808.200 ;
        RECT 658.950 806.100 661.050 808.200 ;
        RECT 628.950 802.950 631.050 805.050 ;
        RECT 631.950 802.950 634.050 805.050 ;
        RECT 634.950 802.950 637.050 805.050 ;
        RECT 637.950 802.950 640.050 805.050 ;
        RECT 632.400 801.900 633.600 802.950 ;
        RECT 631.950 796.950 634.050 801.900 ;
        RECT 638.400 796.050 639.600 802.950 ;
        RECT 644.400 802.050 645.600 806.100 ;
        RECT 653.400 805.050 654.600 806.100 ;
        RECT 659.400 805.050 660.600 806.100 ;
        RECT 667.950 805.950 670.050 808.050 ;
        RECT 676.950 806.100 679.050 808.200 ;
        RECT 682.950 806.100 685.050 808.200 ;
        RECT 652.950 802.950 655.050 805.050 ;
        RECT 655.950 802.950 658.050 805.050 ;
        RECT 658.950 802.950 661.050 805.050 ;
        RECT 661.950 802.950 664.050 805.050 ;
        RECT 643.950 799.950 646.050 802.050 ;
        RECT 649.950 799.950 652.050 802.050 ;
        RECT 656.400 801.900 657.600 802.950 ;
        RECT 643.950 796.800 646.050 798.900 ;
        RECT 637.950 793.950 640.050 796.050 ;
        RECT 622.950 790.950 625.050 793.050 ;
        RECT 637.950 790.800 640.050 792.900 ;
        RECT 613.950 778.950 616.050 781.050 ;
        RECT 589.950 772.950 592.050 775.050 ;
        RECT 577.950 769.950 580.050 772.050 ;
        RECT 571.950 762.600 576.000 763.050 ;
        RECT 556.950 754.800 559.050 756.900 ;
        RECT 559.950 754.950 562.050 757.050 ;
        RECT 562.950 754.950 565.050 757.050 ;
        RECT 550.950 742.950 553.050 745.050 ;
        RECT 553.950 739.950 556.050 742.050 ;
        RECT 532.950 736.950 535.050 739.050 ;
        RECT 533.400 712.050 534.600 736.950 ;
        RECT 550.950 733.950 553.050 736.050 ;
        RECT 541.950 729.000 544.050 733.050 ;
        RECT 542.400 727.050 543.600 729.000 ;
        RECT 538.950 724.950 541.050 727.050 ;
        RECT 541.950 724.950 544.050 727.050 ;
        RECT 532.950 709.950 535.050 712.050 ;
        RECT 539.400 709.050 540.600 724.950 ;
        RECT 538.950 706.950 541.050 709.050 ;
        RECT 551.400 706.050 552.600 733.950 ;
        RECT 544.950 703.950 547.050 706.050 ;
        RECT 550.950 703.950 553.050 706.050 ;
        RECT 538.800 702.000 540.900 702.900 ;
        RECT 538.800 700.800 541.050 702.000 ;
        RECT 541.950 700.950 544.050 703.050 ;
        RECT 538.950 697.950 541.050 700.800 ;
        RECT 530.400 686.400 537.600 687.600 ;
        RECT 529.950 683.100 532.050 685.200 ;
        RECT 530.400 682.050 531.600 683.100 ;
        RECT 536.400 682.050 537.600 686.400 ;
        RECT 526.950 679.950 529.050 682.050 ;
        RECT 529.950 679.950 532.050 682.050 ;
        RECT 532.950 679.950 535.050 682.050 ;
        RECT 535.950 679.950 538.050 682.050 ;
        RECT 521.400 677.400 525.600 678.600 ;
        RECT 527.400 678.000 528.600 679.950 ;
        RECT 533.400 678.900 534.600 679.950 ;
        RECT 542.400 678.900 543.600 700.950 ;
        RECT 545.400 700.050 546.600 703.950 ;
        RECT 554.400 703.050 555.600 739.950 ;
        RECT 560.400 736.050 561.600 754.950 ;
        RECT 562.950 748.950 565.050 751.050 ;
        RECT 559.950 733.950 562.050 736.050 ;
        RECT 563.400 727.050 564.600 748.950 ;
        RECT 566.400 748.050 567.600 761.100 ;
        RECT 571.950 760.950 576.600 762.600 ;
        RECT 580.950 761.100 583.050 763.200 ;
        RECT 575.400 760.050 576.600 760.950 ;
        RECT 581.400 760.050 582.600 761.100 ;
        RECT 574.950 757.950 577.050 760.050 ;
        RECT 577.950 757.950 580.050 760.050 ;
        RECT 580.950 757.950 583.050 760.050 ;
        RECT 583.950 757.950 586.050 760.050 ;
        RECT 578.400 756.900 579.600 757.950 ;
        RECT 577.950 754.800 580.050 756.900 ;
        RECT 584.400 751.050 585.600 757.950 ;
        RECT 583.950 748.950 586.050 751.050 ;
        RECT 565.950 745.950 568.050 748.050 ;
        RECT 571.800 745.950 573.900 748.050 ;
        RECT 574.950 745.950 577.050 748.050 ;
        RECT 559.950 724.950 562.050 727.050 ;
        RECT 562.950 724.950 565.050 727.050 ;
        RECT 560.400 715.050 561.600 724.950 ;
        RECT 572.400 721.050 573.600 745.950 ;
        RECT 562.950 718.950 565.050 721.050 ;
        RECT 571.950 718.950 574.050 721.050 ;
        RECT 559.950 712.950 562.050 715.050 ;
        RECT 553.950 700.950 556.050 703.050 ;
        RECT 544.950 697.950 547.050 700.050 ;
        RECT 544.950 691.950 547.050 694.050 ;
        RECT 545.400 685.200 546.600 691.950 ;
        RECT 563.400 685.200 564.600 718.950 ;
        RECT 565.950 712.950 568.050 715.050 ;
        RECT 571.950 712.950 574.050 715.050 ;
        RECT 544.950 683.100 547.050 685.200 ;
        RECT 550.950 683.100 553.050 685.200 ;
        RECT 562.950 683.100 565.050 685.200 ;
        RECT 508.950 673.950 511.050 676.050 ;
        RECT 520.950 673.950 523.050 676.050 ;
        RECT 499.950 670.950 502.050 673.050 ;
        RECT 505.950 655.950 508.050 658.050 ;
        RECT 496.950 652.950 499.050 655.050 ;
        RECT 499.950 650.100 502.050 652.200 ;
        RECT 506.400 652.050 507.600 655.950 ;
        RECT 500.400 649.050 501.600 650.100 ;
        RECT 505.950 649.950 508.050 652.050 ;
        RECT 493.950 646.950 496.050 649.050 ;
        RECT 499.950 646.950 502.050 649.050 ;
        RECT 502.950 646.950 505.050 649.050 ;
        RECT 494.400 634.050 495.600 646.950 ;
        RECT 503.400 645.900 504.600 646.950 ;
        RECT 502.950 643.800 505.050 645.900 ;
        RECT 503.400 637.050 504.600 643.800 ;
        RECT 509.400 640.050 510.600 673.950 ;
        RECT 511.950 664.950 514.050 667.050 ;
        RECT 512.400 646.050 513.600 664.950 ;
        RECT 521.400 664.050 522.600 673.950 ;
        RECT 520.950 661.950 523.050 664.050 ;
        RECT 521.400 649.050 522.600 661.950 ;
        RECT 524.400 661.050 525.600 677.400 ;
        RECT 526.950 676.050 529.050 678.000 ;
        RECT 532.950 676.800 535.050 678.900 ;
        RECT 541.950 676.800 544.050 678.900 ;
        RECT 545.400 676.050 546.600 683.100 ;
        RECT 551.400 682.050 552.600 683.100 ;
        RECT 550.950 679.950 553.050 682.050 ;
        RECT 553.950 679.950 556.050 682.050 ;
        RECT 554.400 678.900 555.600 679.950 ;
        RECT 553.950 676.800 556.050 678.900 ;
        RECT 526.800 675.000 529.050 676.050 ;
        RECT 526.800 673.950 528.900 675.000 ;
        RECT 529.950 673.950 532.050 676.050 ;
        RECT 544.950 673.950 547.050 676.050 ;
        RECT 550.950 673.950 553.050 676.050 ;
        RECT 530.400 670.050 531.600 673.950 ;
        RECT 529.950 667.950 532.050 670.050 ;
        RECT 523.950 658.950 526.050 661.050 ;
        RECT 529.950 650.100 532.050 652.200 ;
        RECT 541.950 651.600 544.050 652.200 ;
        RECT 544.950 651.600 547.050 655.050 ;
        RECT 547.950 652.950 550.050 655.050 ;
        RECT 541.950 651.000 547.050 651.600 ;
        RECT 541.950 650.400 546.600 651.000 ;
        RECT 541.950 650.100 544.050 650.400 ;
        RECT 517.950 646.950 520.050 649.050 ;
        RECT 520.950 646.950 523.050 649.050 ;
        RECT 511.950 643.950 514.050 646.050 ;
        RECT 518.400 645.900 519.600 646.950 ;
        RECT 517.950 643.800 520.050 645.900 ;
        RECT 508.950 637.950 511.050 640.050 ;
        RECT 502.950 634.950 505.050 637.050 ;
        RECT 493.950 631.950 496.050 634.050 ;
        RECT 505.950 631.950 508.050 634.050 ;
        RECT 487.950 628.950 490.050 631.050 ;
        RECT 484.950 616.950 487.050 619.050 ;
        RECT 485.400 606.600 486.600 616.950 ;
        RECT 490.950 614.400 493.050 616.500 ;
        RECT 485.400 605.400 489.600 606.600 ;
        RECT 488.400 604.050 489.600 605.400 ;
        RECT 472.950 601.950 475.050 604.050 ;
        RECT 475.950 601.950 478.050 604.050 ;
        RECT 478.950 601.950 481.050 604.050 ;
        RECT 481.950 601.950 484.050 604.050 ;
        RECT 487.950 601.950 490.050 604.050 ;
        RECT 476.400 600.900 477.600 601.950 ;
        RECT 440.400 599.400 444.600 600.600 ;
        RECT 461.400 599.400 465.600 600.600 ;
        RECT 424.950 572.100 427.050 574.200 ;
        RECT 433.950 572.100 436.050 574.200 ;
        RECT 409.950 568.950 412.050 571.050 ;
        RECT 410.400 567.900 411.600 568.950 ;
        RECT 398.400 566.400 402.600 567.600 ;
        RECT 385.950 559.950 388.050 562.050 ;
        RECT 391.950 559.950 394.050 562.050 ;
        RECT 391.950 553.950 394.050 556.050 ;
        RECT 388.950 547.950 391.050 550.050 ;
        RECT 389.400 541.050 390.600 547.950 ;
        RECT 392.400 544.050 393.600 553.950 ;
        RECT 391.950 541.950 394.050 544.050 ;
        RECT 388.950 538.950 391.050 541.050 ;
        RECT 358.950 535.950 361.050 538.050 ;
        RECT 373.950 535.950 376.050 538.050 ;
        RECT 359.400 508.050 360.600 535.950 ;
        RECT 382.950 529.950 385.050 532.050 ;
        RECT 373.950 527.100 376.050 529.200 ;
        RECT 379.950 527.100 382.050 529.200 ;
        RECT 374.400 526.050 375.600 527.100 ;
        RECT 370.950 523.950 373.050 526.050 ;
        RECT 373.950 523.950 376.050 526.050 ;
        RECT 371.400 520.050 372.600 523.950 ;
        RECT 380.400 520.050 381.600 527.100 ;
        RECT 383.400 520.050 384.600 529.950 ;
        RECT 392.400 526.050 393.600 541.950 ;
        RECT 398.400 526.050 399.600 566.400 ;
        RECT 409.950 565.800 412.050 567.900 ;
        RECT 425.400 556.050 426.600 572.100 ;
        RECT 434.400 571.050 435.600 572.100 ;
        RECT 430.950 568.950 433.050 571.050 ;
        RECT 433.950 568.950 436.050 571.050 ;
        RECT 431.400 567.900 432.600 568.950 ;
        RECT 430.950 565.800 433.050 567.900 ;
        RECT 436.950 567.600 439.050 567.900 ;
        RECT 440.400 567.600 441.600 599.400 ;
        RECT 448.950 572.100 451.050 574.200 ;
        RECT 449.400 571.050 450.600 572.100 ;
        RECT 448.950 568.950 451.050 571.050 ;
        RECT 451.950 568.950 454.050 571.050 ;
        RECT 452.400 567.900 453.600 568.950 ;
        RECT 436.950 566.400 441.600 567.600 ;
        RECT 436.950 565.800 439.050 566.400 ;
        RECT 451.950 565.800 454.050 567.900 ;
        RECT 424.950 553.950 427.050 556.050 ;
        RECT 400.950 535.950 403.050 538.050 ;
        RECT 424.950 536.400 427.050 538.500 ;
        RECT 388.950 523.950 391.050 526.050 ;
        RECT 391.950 523.950 394.050 526.050 ;
        RECT 397.950 523.950 400.050 526.050 ;
        RECT 371.400 518.400 376.050 520.050 ;
        RECT 372.000 517.950 376.050 518.400 ;
        RECT 379.950 517.950 382.050 520.050 ;
        RECT 382.950 517.950 385.050 520.050 ;
        RECT 389.400 511.050 390.600 523.950 ;
        RECT 401.400 523.050 402.600 535.950 ;
        RECT 421.950 532.950 424.050 535.050 ;
        RECT 406.950 528.000 409.050 532.050 ;
        RECT 407.400 526.050 408.600 528.000 ;
        RECT 412.950 527.100 415.050 529.200 ;
        RECT 413.400 526.050 414.600 527.100 ;
        RECT 422.400 526.050 423.600 532.950 ;
        RECT 406.950 523.950 409.050 526.050 ;
        RECT 409.950 523.950 412.050 526.050 ;
        RECT 412.950 523.950 415.050 526.050 ;
        RECT 415.950 523.950 418.050 526.050 ;
        RECT 421.950 523.950 424.050 526.050 ;
        RECT 400.950 520.950 403.050 523.050 ;
        RECT 410.400 522.900 411.600 523.950 ;
        RECT 409.950 520.800 412.050 522.900 ;
        RECT 397.950 517.950 400.050 520.050 ;
        RECT 388.950 508.950 391.050 511.050 ;
        RECT 358.950 505.950 361.050 508.050 ;
        RECT 370.950 505.950 373.050 508.050 ;
        RECT 361.950 500.400 364.050 502.500 ;
        RECT 356.400 497.400 360.600 498.600 ;
        RECT 352.950 494.100 355.050 496.200 ;
        RECT 353.400 493.050 354.600 494.100 ;
        RECT 359.400 493.050 360.600 497.400 ;
        RECT 337.950 490.950 340.050 493.050 ;
        RECT 343.950 490.950 346.050 493.050 ;
        RECT 346.950 490.950 349.050 493.050 ;
        RECT 349.950 490.950 352.050 493.050 ;
        RECT 352.950 490.950 355.050 493.050 ;
        RECT 358.950 490.950 361.050 493.050 ;
        RECT 344.400 489.000 345.600 490.950 ;
        RECT 350.400 489.900 351.600 490.950 ;
        RECT 343.950 484.950 346.050 489.000 ;
        RECT 349.950 487.800 352.050 489.900 ;
        RECT 355.950 487.950 358.050 490.050 ;
        RECT 337.950 475.950 340.050 478.050 ;
        RECT 334.950 451.950 337.050 454.050 ;
        RECT 338.400 448.050 339.600 475.950 ;
        RECT 346.950 469.950 349.050 472.050 ;
        RECT 331.950 445.950 334.050 448.050 ;
        RECT 334.950 445.950 337.050 448.050 ;
        RECT 337.950 445.950 340.050 448.050 ;
        RECT 340.950 445.950 343.050 448.050 ;
        RECT 328.950 442.950 331.050 445.050 ;
        RECT 335.400 444.900 336.600 445.950 ;
        RECT 329.400 421.050 330.600 442.950 ;
        RECT 334.950 442.800 337.050 444.900 ;
        RECT 341.400 444.000 342.600 445.950 ;
        RECT 347.400 445.050 348.600 469.950 ;
        RECT 350.400 457.050 351.600 487.800 ;
        RECT 356.400 466.050 357.600 487.950 ;
        RECT 362.850 485.400 364.050 500.400 ;
        RECT 371.400 489.600 372.600 505.950 ;
        RECT 391.950 502.950 394.050 505.050 ;
        RECT 382.950 500.400 385.050 502.500 ;
        RECT 376.950 490.950 379.050 493.050 ;
        RECT 370.950 487.500 373.050 489.600 ;
        RECT 361.950 483.300 364.050 485.400 ;
        RECT 362.850 479.700 364.050 483.300 ;
        RECT 361.950 477.600 364.050 479.700 ;
        RECT 371.400 475.050 372.600 487.500 ;
        RECT 377.400 484.050 378.600 490.950 ;
        RECT 376.950 481.950 379.050 484.050 ;
        RECT 383.100 480.600 384.300 500.400 ;
        RECT 385.950 490.950 388.050 493.050 ;
        RECT 386.400 489.600 387.600 490.950 ;
        RECT 385.950 487.500 388.050 489.600 ;
        RECT 392.400 484.050 393.600 502.950 ;
        RECT 398.400 502.050 399.600 517.950 ;
        RECT 409.950 502.950 412.050 505.050 ;
        RECT 397.950 499.950 400.050 502.050 ;
        RECT 391.950 481.950 394.050 484.050 ;
        RECT 398.400 481.050 399.600 499.950 ;
        RECT 410.400 499.050 411.600 502.950 ;
        RECT 416.400 502.050 417.600 523.950 ;
        RECT 418.950 520.950 421.050 523.050 ;
        RECT 419.400 511.050 420.600 520.950 ;
        RECT 425.700 516.600 426.900 536.400 ;
        RECT 430.950 535.950 433.050 538.050 ;
        RECT 431.400 526.050 432.600 535.950 ;
        RECT 430.950 523.950 433.050 526.050 ;
        RECT 437.400 519.600 438.600 565.800 ;
        RECT 442.950 562.950 445.050 565.050 ;
        RECT 443.400 550.050 444.600 562.950 ;
        RECT 442.950 547.950 445.050 550.050 ;
        RECT 461.400 547.050 462.600 599.400 ;
        RECT 475.950 598.800 478.050 600.900 ;
        RECT 472.950 595.950 475.050 598.050 ;
        RECT 463.950 571.950 466.050 574.050 ;
        RECT 460.950 544.950 463.050 547.050 ;
        RECT 464.400 544.050 465.600 571.950 ;
        RECT 473.400 571.050 474.600 595.950 ;
        RECT 472.950 568.950 475.050 571.050 ;
        RECT 475.950 568.950 478.050 571.050 ;
        RECT 476.400 567.900 477.600 568.950 ;
        RECT 482.400 568.050 483.600 601.950 ;
        RECT 484.950 592.950 487.050 595.050 ;
        RECT 491.700 594.600 492.900 614.400 ;
        RECT 502.950 607.950 505.050 610.050 ;
        RECT 496.950 605.400 499.050 607.500 ;
        RECT 497.400 604.050 498.600 605.400 ;
        RECT 496.950 601.950 499.050 604.050 ;
        RECT 503.400 600.600 504.600 607.950 ;
        RECT 500.400 599.400 504.600 600.600 ;
        RECT 475.950 565.800 478.050 567.900 ;
        RECT 481.950 565.950 484.050 568.050 ;
        RECT 472.950 562.950 475.050 565.050 ;
        RECT 466.950 553.950 469.050 556.050 ;
        RECT 439.950 541.950 442.050 544.050 ;
        RECT 463.950 541.950 466.050 544.050 ;
        RECT 440.400 522.600 441.600 541.950 ;
        RECT 467.400 541.050 468.600 553.950 ;
        RECT 469.950 541.950 472.050 544.050 ;
        RECT 445.950 537.300 448.050 539.400 ;
        RECT 466.950 538.950 469.050 541.050 ;
        RECT 445.950 533.700 447.150 537.300 ;
        RECT 457.950 535.950 460.050 538.050 ;
        RECT 445.950 531.600 448.050 533.700 ;
        RECT 439.950 520.500 442.050 522.600 ;
        RECT 437.400 518.400 441.600 519.600 ;
        RECT 424.950 514.500 427.050 516.600 ;
        RECT 418.950 508.950 421.050 511.050 ;
        RECT 433.950 508.950 436.050 511.050 ;
        RECT 415.950 499.950 418.050 502.050 ;
        RECT 409.950 496.950 412.050 499.050 ;
        RECT 406.950 494.100 409.050 496.200 ;
        RECT 407.400 493.050 408.600 494.100 ;
        RECT 406.950 490.950 409.050 493.050 ;
        RECT 409.950 490.950 412.050 493.050 ;
        RECT 410.400 484.050 411.600 490.950 ;
        RECT 382.950 478.500 385.050 480.600 ;
        RECT 397.950 478.950 400.050 481.050 ;
        RECT 409.950 478.950 412.050 484.050 ;
        RECT 370.950 472.950 373.050 475.050 ;
        RECT 361.950 469.950 364.050 472.050 ;
        RECT 355.950 463.950 358.050 466.050 ;
        RECT 362.400 457.050 363.600 469.950 ;
        RECT 416.400 466.050 417.600 499.950 ;
        RECT 419.400 478.050 420.600 508.950 ;
        RECT 434.400 502.050 435.600 508.950 ;
        RECT 433.950 499.950 436.050 502.050 ;
        RECT 427.950 495.000 430.050 499.050 ;
        RECT 428.400 493.050 429.600 495.000 ;
        RECT 434.400 493.050 435.600 499.950 ;
        RECT 424.950 490.950 427.050 493.050 ;
        RECT 427.950 490.950 430.050 493.050 ;
        RECT 430.950 490.950 433.050 493.050 ;
        RECT 433.950 490.950 436.050 493.050 ;
        RECT 425.400 489.900 426.600 490.950 ;
        RECT 431.400 489.900 432.600 490.950 ;
        RECT 440.400 490.050 441.600 518.400 ;
        RECT 445.950 516.600 447.150 531.600 ;
        RECT 454.950 529.800 457.050 531.900 ;
        RECT 448.950 523.950 451.050 526.050 ;
        RECT 449.400 522.600 450.600 523.950 ;
        RECT 448.950 520.500 451.050 522.600 ;
        RECT 445.950 514.500 448.050 516.600 ;
        RECT 442.950 499.950 445.050 502.050 ;
        RECT 451.950 499.950 454.050 502.050 ;
        RECT 424.950 487.800 427.050 489.900 ;
        RECT 430.950 487.800 433.050 489.900 ;
        RECT 439.950 487.950 442.050 490.050 ;
        RECT 443.400 484.050 444.600 499.950 ;
        RECT 452.400 493.050 453.600 499.950 ;
        RECT 455.400 499.050 456.600 529.800 ;
        RECT 458.400 523.050 459.600 535.950 ;
        RECT 470.400 532.050 471.600 541.950 ;
        RECT 469.950 529.950 472.050 532.050 ;
        RECT 473.400 529.050 474.600 562.950 ;
        RECT 478.950 553.950 481.050 556.050 ;
        RECT 475.950 532.950 478.050 535.050 ;
        RECT 472.950 528.600 475.050 529.050 ;
        RECT 470.400 527.400 475.050 528.600 ;
        RECT 470.400 526.050 471.600 527.400 ;
        RECT 472.950 526.950 475.050 527.400 ;
        RECT 466.950 523.950 469.050 526.050 ;
        RECT 469.950 523.950 472.050 526.050 ;
        RECT 457.950 520.950 460.050 523.050 ;
        RECT 467.400 522.900 468.600 523.950 ;
        RECT 466.950 520.800 469.050 522.900 ;
        RECT 472.950 520.950 475.050 523.050 ;
        RECT 457.950 502.950 460.050 505.050 ;
        RECT 454.950 496.950 457.050 499.050 ;
        RECT 458.400 493.050 459.600 502.950 ;
        RECT 466.950 500.400 469.050 502.500 ;
        RECT 448.950 490.950 451.050 493.050 ;
        RECT 451.950 490.950 454.050 493.050 ;
        RECT 454.950 490.950 457.050 493.050 ;
        RECT 457.950 490.950 460.050 493.050 ;
        RECT 463.950 490.950 466.050 493.050 ;
        RECT 449.400 489.900 450.600 490.950 ;
        RECT 455.400 489.900 456.600 490.950 ;
        RECT 448.950 487.800 451.050 489.900 ;
        RECT 454.950 487.800 457.050 489.900 ;
        RECT 424.950 481.950 427.050 484.050 ;
        RECT 442.950 481.950 445.050 484.050 ;
        RECT 418.950 475.950 421.050 478.050 ;
        RECT 421.950 472.950 424.050 475.050 ;
        RECT 370.950 463.950 373.050 466.050 ;
        RECT 415.950 463.950 418.050 466.050 ;
        RECT 349.950 454.950 352.050 457.050 ;
        RECT 361.950 454.950 364.050 457.050 ;
        RECT 340.950 439.950 343.050 444.000 ;
        RECT 346.950 442.950 349.050 445.050 ;
        RECT 337.950 436.950 340.050 439.050 ;
        RECT 328.950 418.950 331.050 421.050 ;
        RECT 334.950 418.950 337.050 421.050 ;
        RECT 326.400 416.400 330.600 417.600 ;
        RECT 313.950 412.950 316.050 415.050 ;
        RECT 316.950 412.950 319.050 415.050 ;
        RECT 319.950 412.950 322.050 415.050 ;
        RECT 322.950 412.950 325.050 415.050 ;
        RECT 317.400 411.900 318.600 412.950 ;
        RECT 323.400 411.900 324.600 412.950 ;
        RECT 316.950 409.800 319.050 411.900 ;
        RECT 322.950 409.800 325.050 411.900 ;
        RECT 329.400 409.050 330.600 416.400 ;
        RECT 328.950 408.600 331.050 409.050 ;
        RECT 328.950 407.400 333.600 408.600 ;
        RECT 328.950 406.950 331.050 407.400 ;
        RECT 316.950 382.950 319.050 385.050 ;
        RECT 307.950 349.950 310.050 352.050 ;
        RECT 277.950 346.950 280.050 349.050 ;
        RECT 271.950 338.100 274.050 340.200 ;
        RECT 272.400 337.050 273.600 338.100 ;
        RECT 278.400 337.050 279.600 346.950 ;
        RECT 289.950 344.400 292.050 346.500 ;
        RECT 310.950 344.400 313.050 346.500 ;
        RECT 271.950 334.950 274.050 337.050 ;
        RECT 274.950 334.950 277.050 337.050 ;
        RECT 277.950 334.950 280.050 337.050 ;
        RECT 286.950 334.950 289.050 337.050 ;
        RECT 265.950 328.950 268.050 331.050 ;
        RECT 275.400 325.050 276.600 334.950 ;
        RECT 287.400 333.600 288.600 334.950 ;
        RECT 280.950 331.500 283.050 333.600 ;
        RECT 286.950 331.500 289.050 333.600 ;
        RECT 274.950 322.950 277.050 325.050 ;
        RECT 271.950 302.400 274.050 304.500 ;
        RECT 265.950 298.950 268.050 301.050 ;
        RECT 266.400 292.050 267.600 298.950 ;
        RECT 265.950 289.950 268.050 292.050 ;
        RECT 259.950 280.950 262.050 283.050 ;
        RECT 272.100 282.600 273.300 302.400 ;
        RECT 281.400 295.500 282.600 331.500 ;
        RECT 290.700 324.600 291.900 344.400 ;
        RECT 304.950 337.950 307.050 340.050 ;
        RECT 295.950 334.950 298.050 337.050 ;
        RECT 289.950 322.500 292.050 324.600 ;
        RECT 292.950 304.950 295.050 307.050 ;
        RECT 293.400 301.050 294.600 304.950 ;
        RECT 283.950 298.950 286.050 301.050 ;
        RECT 292.950 298.950 295.050 301.050 ;
        RECT 274.950 293.400 277.050 295.500 ;
        RECT 280.950 293.400 283.050 295.500 ;
        RECT 275.400 292.050 276.600 293.400 ;
        RECT 274.950 289.950 277.050 292.050 ;
        RECT 271.950 280.500 274.050 282.600 ;
        RECT 281.400 277.050 282.600 293.400 ;
        RECT 284.400 280.050 285.600 298.950 ;
        RECT 293.400 292.050 294.600 298.950 ;
        RECT 296.400 298.050 297.600 334.950 ;
        RECT 298.950 331.950 301.050 334.050 ;
        RECT 305.400 333.900 306.600 337.950 ;
        RECT 299.400 301.050 300.600 331.950 ;
        RECT 304.950 331.800 307.050 333.900 ;
        RECT 310.950 329.400 312.150 344.400 ;
        RECT 313.950 338.400 316.050 340.500 ;
        RECT 317.400 339.600 318.600 382.950 ;
        RECT 322.950 371.100 325.050 373.200 ;
        RECT 323.400 370.050 324.600 371.100 ;
        RECT 322.950 367.950 325.050 370.050 ;
        RECT 325.950 367.950 328.050 370.050 ;
        RECT 326.400 361.050 327.600 367.950 ;
        RECT 332.400 364.050 333.600 407.400 ;
        RECT 335.400 376.050 336.600 418.950 ;
        RECT 338.400 412.050 339.600 436.950 ;
        RECT 350.400 424.050 351.600 454.950 ;
        RECT 355.950 449.100 358.050 451.200 ;
        RECT 356.400 448.050 357.600 449.100 ;
        RECT 362.400 448.050 363.600 454.950 ;
        RECT 355.950 445.950 358.050 448.050 ;
        RECT 358.950 445.950 361.050 448.050 ;
        RECT 361.950 445.950 364.050 448.050 ;
        RECT 364.950 445.950 367.050 448.050 ;
        RECT 359.400 444.900 360.600 445.950 ;
        RECT 358.950 442.800 361.050 444.900 ;
        RECT 365.400 444.600 366.600 445.950 ;
        RECT 365.400 443.400 369.600 444.600 ;
        RECT 364.950 439.950 367.050 442.050 ;
        RECT 358.950 433.950 361.050 436.050 ;
        RECT 349.950 421.950 352.050 424.050 ;
        RECT 346.950 416.100 349.050 418.200 ;
        RECT 352.950 416.100 355.050 418.200 ;
        RECT 347.400 415.050 348.600 416.100 ;
        RECT 353.400 415.050 354.600 416.100 ;
        RECT 343.950 412.950 346.050 415.050 ;
        RECT 346.950 412.950 349.050 415.050 ;
        RECT 349.950 412.950 352.050 415.050 ;
        RECT 352.950 412.950 355.050 415.050 ;
        RECT 337.950 409.950 340.050 412.050 ;
        RECT 344.400 411.900 345.600 412.950 ;
        RECT 343.950 409.800 346.050 411.900 ;
        RECT 350.400 411.000 351.600 412.950 ;
        RECT 349.950 406.950 352.050 411.000 ;
        RECT 359.400 400.050 360.600 433.950 ;
        RECT 365.400 424.050 366.600 439.950 ;
        RECT 368.400 439.050 369.600 443.400 ;
        RECT 371.400 442.050 372.600 463.950 ;
        RECT 394.950 459.300 397.050 461.400 ;
        RECT 395.850 455.700 397.050 459.300 ;
        RECT 415.950 458.400 418.050 460.500 ;
        RECT 394.950 453.600 397.050 455.700 ;
        RECT 382.950 449.100 385.050 451.200 ;
        RECT 383.400 448.050 384.600 449.100 ;
        RECT 379.950 445.950 382.050 448.050 ;
        RECT 382.950 445.950 385.050 448.050 ;
        RECT 385.950 445.950 388.050 448.050 ;
        RECT 391.950 445.950 394.050 448.050 ;
        RECT 373.950 442.950 376.050 445.050 ;
        RECT 380.400 444.900 381.600 445.950 ;
        RECT 370.950 439.950 373.050 442.050 ;
        RECT 367.950 436.950 370.050 439.050 ;
        RECT 374.400 433.050 375.600 442.950 ;
        RECT 379.950 442.800 382.050 444.900 ;
        RECT 379.950 439.650 382.050 441.750 ;
        RECT 373.950 430.950 376.050 433.050 ;
        RECT 364.950 421.950 367.050 424.050 ;
        RECT 365.400 415.050 366.600 421.950 ;
        RECT 380.400 421.050 381.600 439.650 ;
        RECT 386.400 430.050 387.600 445.950 ;
        RECT 392.400 444.600 393.600 445.950 ;
        RECT 391.950 442.500 394.050 444.600 ;
        RECT 395.850 438.600 397.050 453.600 ;
        RECT 400.950 451.950 403.050 454.050 ;
        RECT 394.950 436.500 397.050 438.600 ;
        RECT 401.400 432.600 402.600 451.950 ;
        RECT 409.950 450.000 412.050 454.050 ;
        RECT 410.400 448.050 411.600 450.000 ;
        RECT 409.950 445.950 412.050 448.050 ;
        RECT 406.950 442.950 409.050 445.050 ;
        RECT 398.400 431.400 402.600 432.600 ;
        RECT 385.950 427.950 388.050 430.050 ;
        RECT 386.400 424.050 387.600 427.950 ;
        RECT 385.950 421.950 388.050 424.050 ;
        RECT 379.950 418.950 382.050 421.050 ;
        RECT 370.950 416.100 373.050 418.200 ;
        RECT 371.400 415.050 372.600 416.100 ;
        RECT 364.950 412.950 367.050 415.050 ;
        RECT 367.950 412.950 370.050 415.050 ;
        RECT 370.950 412.950 373.050 415.050 ;
        RECT 373.950 412.950 376.050 415.050 ;
        RECT 368.400 411.000 369.600 412.950 ;
        RECT 367.950 406.950 370.050 411.000 ;
        RECT 374.400 403.050 375.600 412.950 ;
        RECT 380.400 412.050 381.600 418.950 ;
        RECT 382.950 415.950 385.050 418.050 ;
        RECT 391.950 417.000 394.050 421.050 ;
        RECT 379.950 409.950 382.050 412.050 ;
        RECT 383.400 406.050 384.600 415.950 ;
        RECT 392.400 415.050 393.600 417.000 ;
        RECT 398.400 415.050 399.600 431.400 ;
        RECT 388.950 412.950 391.050 415.050 ;
        RECT 391.950 412.950 394.050 415.050 ;
        RECT 394.950 412.950 397.050 415.050 ;
        RECT 397.950 412.950 400.050 415.050 ;
        RECT 385.950 409.950 388.050 412.050 ;
        RECT 389.400 411.900 390.600 412.950 ;
        RECT 395.400 411.900 396.600 412.950 ;
        RECT 407.400 411.900 408.600 442.950 ;
        RECT 416.100 438.600 417.300 458.400 ;
        RECT 422.400 457.050 423.600 472.950 ;
        RECT 421.950 454.950 424.050 457.050 ;
        RECT 422.400 450.600 423.600 454.950 ;
        RECT 419.400 449.400 423.600 450.600 ;
        RECT 419.400 448.050 420.600 449.400 ;
        RECT 418.950 445.950 421.050 448.050 ;
        RECT 415.950 436.500 418.050 438.600 ;
        RECT 425.400 430.050 426.600 481.950 ;
        RECT 427.950 469.950 430.050 472.050 ;
        RECT 424.950 427.950 427.050 430.050 ;
        RECT 424.950 424.800 427.050 426.900 ;
        RECT 409.950 415.950 412.050 418.050 ;
        RECT 418.950 416.100 421.050 418.200 ;
        RECT 382.950 403.950 385.050 406.050 ;
        RECT 361.950 402.600 364.050 403.050 ;
        RECT 367.950 402.600 370.050 403.050 ;
        RECT 361.950 401.400 370.050 402.600 ;
        RECT 361.950 400.950 364.050 401.400 ;
        RECT 367.950 400.950 370.050 401.400 ;
        RECT 373.950 400.950 376.050 403.050 ;
        RECT 358.950 397.950 361.050 400.050 ;
        RECT 364.950 397.950 367.050 400.050 ;
        RECT 340.950 382.950 343.050 385.050 ;
        RECT 334.950 373.950 337.050 376.050 ;
        RECT 341.400 370.050 342.600 382.950 ;
        RECT 358.950 381.300 361.050 383.400 ;
        RECT 359.850 377.700 361.050 381.300 ;
        RECT 346.950 372.000 349.050 376.050 ;
        RECT 358.950 375.600 361.050 377.700 ;
        RECT 347.400 370.050 348.600 372.000 ;
        RECT 337.950 367.950 340.050 370.050 ;
        RECT 340.950 367.950 343.050 370.050 ;
        RECT 343.950 367.950 346.050 370.050 ;
        RECT 346.950 367.950 349.050 370.050 ;
        RECT 355.950 367.950 358.050 370.050 ;
        RECT 338.400 366.900 339.600 367.950 ;
        RECT 344.400 366.900 345.600 367.950 ;
        RECT 337.950 364.800 340.050 366.900 ;
        RECT 343.950 364.800 346.050 366.900 ;
        RECT 356.400 366.000 357.600 367.950 ;
        RECT 331.950 361.950 334.050 364.050 ;
        RECT 325.950 358.950 328.050 361.050 ;
        RECT 338.400 349.050 339.600 364.800 ;
        RECT 355.950 361.950 358.050 366.000 ;
        RECT 359.850 360.600 361.050 375.600 ;
        RECT 358.950 358.500 361.050 360.600 ;
        RECT 361.950 352.950 364.050 355.050 ;
        RECT 337.950 346.950 340.050 349.050 ;
        RECT 317.400 338.400 321.600 339.600 ;
        RECT 314.400 337.050 315.600 338.400 ;
        RECT 313.950 334.950 316.050 337.050 ;
        RECT 310.950 327.300 313.050 329.400 ;
        RECT 310.950 323.700 312.150 327.300 ;
        RECT 310.950 321.600 313.050 323.700 ;
        RECT 304.950 313.950 307.050 316.050 ;
        RECT 298.950 298.950 301.050 301.050 ;
        RECT 295.950 295.950 298.050 298.050 ;
        RECT 300.000 294.600 304.050 295.050 ;
        RECT 299.400 292.950 304.050 294.600 ;
        RECT 299.400 292.050 300.600 292.950 ;
        RECT 289.950 289.950 292.050 292.050 ;
        RECT 292.950 289.950 295.050 292.050 ;
        RECT 295.950 289.950 298.050 292.050 ;
        RECT 298.950 289.950 301.050 292.050 ;
        RECT 290.400 288.000 291.600 289.950 ;
        RECT 296.400 288.900 297.600 289.950 ;
        RECT 289.950 283.950 292.050 288.000 ;
        RECT 295.950 286.800 298.050 288.900 ;
        RECT 301.950 283.950 304.050 286.050 ;
        RECT 283.950 277.950 286.050 280.050 ;
        RECT 274.950 274.950 277.050 277.050 ;
        RECT 280.950 274.950 283.050 277.050 ;
        RECT 271.950 271.950 274.050 274.050 ;
        RECT 256.950 265.950 259.050 268.050 ;
        RECT 265.950 266.400 268.050 268.500 ;
        RECT 257.400 259.050 258.600 265.950 ;
        RECT 262.950 260.400 265.050 262.500 ;
        RECT 263.400 259.050 264.600 260.400 ;
        RECT 250.950 256.950 253.050 259.050 ;
        RECT 253.950 256.950 256.050 259.050 ;
        RECT 256.950 256.950 259.050 259.050 ;
        RECT 262.950 256.950 265.050 259.050 ;
        RECT 254.400 250.050 255.600 256.950 ;
        RECT 266.850 251.400 268.050 266.400 ;
        RECT 253.950 247.950 256.050 250.050 ;
        RECT 265.950 249.300 268.050 251.400 ;
        RECT 266.850 245.700 268.050 249.300 ;
        RECT 265.950 243.600 268.050 245.700 ;
        RECT 272.400 244.050 273.600 271.950 ;
        RECT 271.950 241.950 274.050 244.050 ;
        RECT 244.950 238.950 247.050 241.050 ;
        RECT 256.950 238.950 259.050 241.050 ;
        RECT 250.950 226.950 253.050 229.050 ;
        RECT 224.850 221.700 226.050 225.300 ;
        RECT 232.950 223.950 235.050 226.050 ;
        RECT 238.950 223.950 241.050 226.050 ;
        RECT 244.950 224.400 247.050 226.500 ;
        RECT 223.950 219.600 226.050 221.700 ;
        RECT 211.950 215.100 214.050 217.200 ;
        RECT 212.400 214.050 213.600 215.100 ;
        RECT 205.950 211.950 208.050 214.050 ;
        RECT 208.950 211.950 211.050 214.050 ;
        RECT 211.950 211.950 214.050 214.050 ;
        RECT 214.950 211.950 217.050 214.050 ;
        RECT 220.950 211.950 223.050 214.050 ;
        RECT 209.400 210.000 210.600 211.950 ;
        RECT 208.950 205.950 211.050 210.000 ;
        RECT 215.400 196.050 216.600 211.950 ;
        RECT 221.400 210.600 222.600 211.950 ;
        RECT 220.950 208.500 223.050 210.600 ;
        RECT 224.850 204.600 226.050 219.600 ;
        RECT 229.950 214.950 232.050 217.050 ;
        RECT 230.400 210.600 231.600 214.950 ;
        RECT 229.950 208.500 232.050 210.600 ;
        RECT 223.950 202.500 226.050 204.600 ;
        RECT 214.950 193.950 217.050 196.050 ;
        RECT 211.950 187.950 214.050 190.050 ;
        RECT 223.950 188.400 226.050 190.500 ;
        RECT 212.400 181.050 213.600 187.950 ;
        RECT 220.950 182.400 223.050 184.500 ;
        RECT 221.400 181.050 222.600 182.400 ;
        RECT 208.950 178.950 211.050 181.050 ;
        RECT 211.950 178.950 214.050 181.050 ;
        RECT 214.950 178.950 217.050 181.050 ;
        RECT 220.950 178.950 223.050 181.050 ;
        RECT 209.400 177.000 210.600 178.950 ;
        RECT 215.400 177.900 216.600 178.950 ;
        RECT 196.950 172.950 199.050 175.050 ;
        RECT 199.950 172.950 202.050 175.050 ;
        RECT 208.950 172.950 211.050 177.000 ;
        RECT 214.950 175.800 217.050 177.900 ;
        RECT 215.400 169.050 216.600 175.800 ;
        RECT 224.850 173.400 226.050 188.400 ;
        RECT 223.950 171.300 226.050 173.400 ;
        RECT 214.950 166.950 217.050 169.050 ;
        RECT 224.850 167.700 226.050 171.300 ;
        RECT 223.950 165.600 226.050 167.700 ;
        RECT 178.950 157.950 181.050 160.050 ;
        RECT 202.950 147.300 205.050 149.400 ;
        RECT 203.850 143.700 205.050 147.300 ;
        RECT 223.950 146.400 226.050 148.500 ;
        RECT 202.950 141.600 205.050 143.700 ;
        RECT 217.950 142.950 220.050 145.050 ;
        RECT 160.950 136.950 163.050 139.050 ;
        RECT 169.950 137.100 172.050 139.200 ;
        RECT 184.950 137.100 187.050 139.200 ;
        RECT 190.950 137.100 193.050 139.200 ;
        RECT 142.950 109.950 145.050 112.050 ;
        RECT 157.950 109.950 160.050 112.050 ;
        RECT 143.400 103.050 144.600 109.950 ;
        RECT 142.950 100.950 145.050 103.050 ;
        RECT 136.950 82.950 139.050 85.050 ;
        RECT 115.950 79.950 118.050 82.050 ;
        RECT 100.950 59.100 103.050 61.200 ;
        RECT 106.950 59.100 109.050 61.200 ;
        RECT 112.950 59.100 115.050 61.200 ;
        RECT 101.400 58.050 102.600 59.100 ;
        RECT 107.400 58.050 108.600 59.100 ;
        RECT 100.950 55.950 103.050 58.050 ;
        RECT 103.950 55.950 106.050 58.050 ;
        RECT 106.950 55.950 109.050 58.050 ;
        RECT 97.950 52.950 100.050 55.050 ;
        RECT 104.400 54.900 105.600 55.950 ;
        RECT 94.950 49.950 97.050 52.050 ;
        RECT 79.950 43.950 82.050 46.050 ;
        RECT 91.950 43.950 94.050 46.050 ;
        RECT 62.400 41.400 69.600 42.600 ;
        RECT 70.950 40.950 73.050 43.050 ;
        RECT 46.950 37.950 49.050 40.050 ;
        RECT 32.400 25.050 33.600 26.100 ;
        RECT 37.950 25.950 40.050 28.050 ;
        RECT 59.400 25.050 60.600 40.950 ;
        RECT 80.400 25.050 81.600 43.950 ;
        RECT 88.950 32.400 91.050 34.500 ;
        RECT 85.950 26.400 88.050 28.500 ;
        RECT 86.400 25.050 87.600 26.400 ;
        RECT 28.950 22.950 31.050 25.050 ;
        RECT 31.950 22.950 34.050 25.050 ;
        RECT 34.950 22.950 37.050 25.050 ;
        RECT 58.950 22.950 61.050 25.050 ;
        RECT 79.950 22.950 82.050 25.050 ;
        RECT 85.950 22.950 88.050 25.050 ;
        RECT 29.400 21.900 30.600 22.950 ;
        RECT 35.400 21.900 36.600 22.950 ;
        RECT 13.950 19.800 16.050 21.900 ;
        RECT 22.950 19.800 25.050 21.900 ;
        RECT 28.950 19.800 31.050 21.900 ;
        RECT 34.950 19.800 37.050 21.900 ;
        RECT 89.850 17.400 91.050 32.400 ;
        RECT 98.400 28.500 99.600 52.950 ;
        RECT 103.950 52.800 106.050 54.900 ;
        RECT 109.950 32.400 112.050 34.500 ;
        RECT 97.950 26.400 100.050 28.500 ;
        RECT 103.950 22.950 106.050 25.050 ;
        RECT 104.400 21.600 105.600 22.950 ;
        RECT 103.950 19.500 106.050 21.600 ;
        RECT 88.950 15.300 91.050 17.400 ;
        RECT 89.850 11.700 91.050 15.300 ;
        RECT 110.100 12.600 111.300 32.400 ;
        RECT 116.400 27.600 117.600 79.950 ;
        RECT 161.400 79.050 162.600 136.950 ;
        RECT 170.400 136.050 171.600 137.100 ;
        RECT 169.950 133.950 172.050 136.050 ;
        RECT 175.950 133.950 178.050 136.050 ;
        RECT 172.950 130.950 175.050 133.050 ;
        RECT 173.400 121.050 174.600 130.950 ;
        RECT 176.400 127.050 177.600 133.950 ;
        RECT 185.400 133.050 186.600 137.100 ;
        RECT 191.400 136.050 192.600 137.100 ;
        RECT 190.950 133.950 193.050 136.050 ;
        RECT 193.950 133.950 196.050 136.050 ;
        RECT 199.950 133.950 202.050 136.050 ;
        RECT 184.950 130.950 187.050 133.050 ;
        RECT 194.400 132.900 195.600 133.950 ;
        RECT 193.950 130.800 196.050 132.900 ;
        RECT 200.400 132.600 201.600 133.950 ;
        RECT 175.950 124.950 178.050 127.050 ;
        RECT 172.950 118.950 175.050 121.050 ;
        RECT 166.950 104.100 169.050 106.200 ;
        RECT 167.400 103.050 168.600 104.100 ;
        RECT 173.400 103.050 174.600 118.950 ;
        RECT 187.950 104.100 190.050 106.200 ;
        RECT 188.400 103.050 189.600 104.100 ;
        RECT 194.400 103.050 195.600 130.800 ;
        RECT 199.950 130.500 202.050 132.600 ;
        RECT 203.850 126.600 205.050 141.600 ;
        RECT 218.400 136.050 219.600 142.950 ;
        RECT 217.950 133.950 220.050 136.050 ;
        RECT 224.100 126.600 225.300 146.400 ;
        RECT 226.950 137.400 229.050 139.500 ;
        RECT 227.400 136.050 228.600 137.400 ;
        RECT 226.950 133.950 229.050 136.050 ;
        RECT 229.950 130.950 232.050 133.050 ;
        RECT 202.950 124.500 205.050 126.600 ;
        RECT 223.950 124.500 226.050 126.600 ;
        RECT 223.950 110.400 226.050 112.500 ;
        RECT 214.950 104.100 217.050 106.200 ;
        RECT 220.950 104.400 223.050 106.500 ;
        RECT 215.400 103.050 216.600 104.100 ;
        RECT 221.400 103.050 222.600 104.400 ;
        RECT 166.950 100.950 169.050 103.050 ;
        RECT 169.950 100.950 172.050 103.050 ;
        RECT 172.950 100.950 175.050 103.050 ;
        RECT 187.950 100.950 190.050 103.050 ;
        RECT 190.950 100.950 193.050 103.050 ;
        RECT 193.950 100.950 196.050 103.050 ;
        RECT 211.950 100.950 214.050 103.050 ;
        RECT 214.950 100.950 217.050 103.050 ;
        RECT 220.950 100.950 223.050 103.050 ;
        RECT 170.400 99.000 171.600 100.950 ;
        RECT 191.400 99.900 192.600 100.950 ;
        RECT 212.400 99.900 213.600 100.950 ;
        RECT 169.950 94.950 172.050 99.000 ;
        RECT 190.950 97.800 193.050 99.900 ;
        RECT 211.950 97.800 214.050 99.900 ;
        RECT 224.850 95.400 226.050 110.400 ;
        RECT 196.950 91.950 199.050 94.050 ;
        RECT 223.950 93.300 226.050 95.400 ;
        RECT 172.950 82.950 175.050 85.050 ;
        RECT 166.950 79.950 169.050 82.050 ;
        RECT 151.950 76.950 154.050 79.050 ;
        RECT 160.950 76.950 163.050 79.050 ;
        RECT 139.950 69.300 142.050 71.400 ;
        RECT 140.850 65.700 142.050 69.300 ;
        RECT 139.950 63.600 142.050 65.700 ;
        RECT 152.400 63.600 153.600 76.950 ;
        RECT 160.950 68.400 163.050 70.500 ;
        RECT 121.950 59.100 124.050 61.200 ;
        RECT 127.950 59.100 130.050 61.200 ;
        RECT 122.400 58.050 123.600 59.100 ;
        RECT 128.400 58.050 129.600 59.100 ;
        RECT 121.950 55.950 124.050 58.050 ;
        RECT 124.950 55.950 127.050 58.050 ;
        RECT 127.950 55.950 130.050 58.050 ;
        RECT 136.950 55.950 139.050 58.050 ;
        RECT 116.400 26.400 120.600 27.600 ;
        RECT 112.950 22.950 115.050 25.050 ;
        RECT 113.400 21.600 114.600 22.950 ;
        RECT 119.400 21.600 120.600 26.400 ;
        RECT 125.400 25.050 126.600 55.950 ;
        RECT 137.400 54.000 138.600 55.950 ;
        RECT 136.950 49.950 139.050 54.000 ;
        RECT 130.950 46.950 133.050 49.050 ;
        RECT 140.850 48.600 142.050 63.600 ;
        RECT 149.400 62.400 153.600 63.600 ;
        RECT 145.950 59.100 148.050 61.200 ;
        RECT 131.400 25.050 132.600 46.950 ;
        RECT 139.950 46.500 142.050 48.600 ;
        RECT 146.400 37.050 147.600 59.100 ;
        RECT 149.400 49.050 150.600 62.400 ;
        RECT 151.950 60.600 156.000 61.050 ;
        RECT 151.950 58.950 156.600 60.600 ;
        RECT 155.400 58.050 156.600 58.950 ;
        RECT 154.950 55.950 157.050 58.050 ;
        RECT 151.950 52.950 154.050 55.050 ;
        RECT 148.950 46.950 151.050 49.050 ;
        RECT 145.950 34.950 148.050 37.050 ;
        RECT 149.400 28.200 150.600 46.950 ;
        RECT 152.400 30.600 153.600 52.950 ;
        RECT 161.100 48.600 162.300 68.400 ;
        RECT 167.400 60.600 168.600 79.950 ;
        RECT 173.400 67.050 174.600 82.950 ;
        RECT 172.950 64.950 175.050 67.050 ;
        RECT 164.400 59.400 168.600 60.600 ;
        RECT 164.400 58.050 165.600 59.400 ;
        RECT 163.950 55.950 166.050 58.050 ;
        RECT 173.400 54.900 174.600 64.950 ;
        RECT 181.950 59.100 184.050 61.200 ;
        RECT 182.400 58.050 183.600 59.100 ;
        RECT 178.950 55.950 181.050 58.050 ;
        RECT 181.950 55.950 184.050 58.050 ;
        RECT 184.950 55.950 187.050 58.050 ;
        RECT 172.950 52.800 175.050 54.900 ;
        RECT 160.950 46.500 163.050 48.600 ;
        RECT 179.400 31.050 180.600 55.950 ;
        RECT 185.400 54.900 186.600 55.950 ;
        RECT 184.950 52.800 187.050 54.900 ;
        RECT 197.400 43.050 198.600 91.950 ;
        RECT 224.850 89.700 226.050 93.300 ;
        RECT 214.950 85.950 217.050 88.050 ;
        RECT 223.950 87.600 226.050 89.700 ;
        RECT 215.400 76.050 216.600 85.950 ;
        RECT 230.400 82.050 231.600 130.950 ;
        RECT 233.400 127.050 234.600 223.950 ;
        RECT 241.950 220.950 244.050 223.050 ;
        RECT 242.400 216.600 243.600 220.950 ;
        RECT 239.400 215.400 243.600 216.600 ;
        RECT 239.400 214.050 240.600 215.400 ;
        RECT 238.950 211.950 241.050 214.050 ;
        RECT 245.100 204.600 246.300 224.400 ;
        RECT 251.400 216.600 252.600 226.950 ;
        RECT 248.400 215.400 255.600 216.600 ;
        RECT 248.400 214.050 249.600 215.400 ;
        RECT 247.950 211.950 250.050 214.050 ;
        RECT 244.950 202.500 247.050 204.600 ;
        RECT 244.950 188.400 247.050 190.500 ;
        RECT 238.950 178.950 241.050 181.050 ;
        RECT 239.400 177.600 240.600 178.950 ;
        RECT 238.950 175.500 241.050 177.600 ;
        RECT 245.100 168.600 246.300 188.400 ;
        RECT 247.950 178.950 250.050 181.050 ;
        RECT 248.400 177.600 249.600 178.950 ;
        RECT 254.400 177.600 255.600 215.400 ;
        RECT 247.950 175.500 250.050 177.600 ;
        RECT 253.950 175.500 256.050 177.600 ;
        RECT 244.950 166.500 247.050 168.600 ;
        RECT 250.950 148.950 253.050 151.050 ;
        RECT 244.950 137.100 247.050 139.200 ;
        RECT 245.400 136.050 246.600 137.100 ;
        RECT 251.400 136.050 252.600 148.950 ;
        RECT 241.950 133.950 244.050 136.050 ;
        RECT 244.950 133.950 247.050 136.050 ;
        RECT 247.950 133.950 250.050 136.050 ;
        RECT 250.950 133.950 253.050 136.050 ;
        RECT 238.950 130.950 241.050 133.050 ;
        RECT 242.400 132.000 243.600 133.950 ;
        RECT 248.400 132.900 249.600 133.950 ;
        RECT 232.950 124.950 235.050 127.050 ;
        RECT 239.400 121.050 240.600 130.950 ;
        RECT 241.950 127.950 244.050 132.000 ;
        RECT 247.950 130.800 250.050 132.900 ;
        RECT 253.950 127.950 256.050 130.050 ;
        RECT 238.950 118.950 241.050 121.050 ;
        RECT 244.950 110.400 247.050 112.500 ;
        RECT 232.950 104.100 235.050 106.200 ;
        RECT 233.400 100.050 234.600 104.100 ;
        RECT 238.950 100.950 241.050 103.050 ;
        RECT 232.950 97.950 235.050 100.050 ;
        RECT 239.400 94.050 240.600 100.950 ;
        RECT 238.950 91.950 241.050 94.050 ;
        RECT 245.100 90.600 246.300 110.400 ;
        RECT 247.950 100.950 250.050 103.050 ;
        RECT 248.400 99.600 249.600 100.950 ;
        RECT 254.400 99.900 255.600 127.950 ;
        RECT 248.400 98.400 252.600 99.600 ;
        RECT 244.950 88.500 247.050 90.600 ;
        RECT 251.400 82.050 252.600 98.400 ;
        RECT 253.950 97.800 256.050 99.900 ;
        RECT 217.950 79.950 220.050 82.050 ;
        RECT 229.950 79.950 232.050 82.050 ;
        RECT 250.950 79.950 253.050 82.050 ;
        RECT 214.950 73.950 217.050 76.050 ;
        RECT 205.950 59.100 208.050 61.200 ;
        RECT 211.950 59.100 214.050 61.200 ;
        RECT 206.400 58.050 207.600 59.100 ;
        RECT 212.400 58.050 213.600 59.100 ;
        RECT 202.950 55.950 205.050 58.050 ;
        RECT 205.950 55.950 208.050 58.050 ;
        RECT 208.950 55.950 211.050 58.050 ;
        RECT 211.950 55.950 214.050 58.050 ;
        RECT 196.950 40.950 199.050 43.050 ;
        RECT 190.950 32.400 193.050 34.500 ;
        RECT 152.400 29.400 156.600 30.600 ;
        RECT 148.950 26.100 151.050 28.200 ;
        RECT 149.400 25.050 150.600 26.100 ;
        RECT 155.400 25.050 156.600 29.400 ;
        RECT 163.950 28.950 166.050 31.050 ;
        RECT 172.950 30.600 177.000 31.050 ;
        RECT 172.950 28.950 177.600 30.600 ;
        RECT 178.950 28.950 181.050 31.050 ;
        RECT 124.950 22.950 127.050 25.050 ;
        RECT 130.950 22.950 133.050 25.050 ;
        RECT 133.950 22.950 136.050 25.050 ;
        RECT 148.950 22.950 151.050 25.050 ;
        RECT 151.950 22.950 154.050 25.050 ;
        RECT 154.950 22.950 157.050 25.050 ;
        RECT 157.950 22.950 160.050 25.050 ;
        RECT 134.400 21.900 135.600 22.950 ;
        RECT 152.400 21.900 153.600 22.950 ;
        RECT 113.400 20.400 120.600 21.600 ;
        RECT 133.950 19.800 136.050 21.900 ;
        RECT 151.950 19.800 154.050 21.900 ;
        RECT 158.400 21.600 159.600 22.950 ;
        RECT 164.400 21.600 165.600 28.950 ;
        RECT 166.950 25.950 169.050 28.050 ;
        RECT 167.400 21.900 168.600 25.950 ;
        RECT 176.400 25.050 177.600 28.950 ;
        RECT 187.950 26.400 190.050 31.050 ;
        RECT 188.400 25.050 189.600 26.400 ;
        RECT 172.950 22.950 175.050 25.050 ;
        RECT 175.950 22.950 178.050 25.050 ;
        RECT 178.950 22.950 181.050 25.050 ;
        RECT 187.950 22.950 190.050 25.050 ;
        RECT 173.400 21.900 174.600 22.950 ;
        RECT 179.400 21.900 180.600 22.950 ;
        RECT 158.400 20.400 165.600 21.600 ;
        RECT 166.950 19.800 169.050 21.900 ;
        RECT 172.950 19.800 175.050 21.900 ;
        RECT 178.950 19.800 181.050 21.900 ;
        RECT 191.850 17.400 193.050 32.400 ;
        RECT 203.400 27.600 204.600 55.950 ;
        RECT 209.400 54.900 210.600 55.950 ;
        RECT 208.950 52.800 211.050 54.900 ;
        RECT 211.950 32.400 214.050 34.500 ;
        RECT 200.400 26.400 204.600 27.600 ;
        RECT 200.400 21.600 201.600 26.400 ;
        RECT 205.950 22.950 208.050 25.050 ;
        RECT 206.400 21.600 207.600 22.950 ;
        RECT 199.950 19.500 202.050 21.600 ;
        RECT 205.950 19.500 208.050 21.600 ;
        RECT 190.950 15.300 193.050 17.400 ;
        RECT 88.950 9.600 91.050 11.700 ;
        RECT 109.950 10.500 112.050 12.600 ;
        RECT 191.850 11.700 193.050 15.300 ;
        RECT 212.100 12.600 213.300 32.400 ;
        RECT 218.400 27.600 219.600 79.950 ;
        RECT 229.950 70.950 232.050 73.050 ;
        RECT 230.400 67.050 231.600 70.950 ;
        RECT 244.950 69.300 247.050 71.400 ;
        RECT 229.950 64.950 232.050 67.050 ;
        RECT 245.850 65.700 247.050 69.300 ;
        RECT 253.950 67.950 256.050 70.050 ;
        RECT 244.950 63.600 247.050 65.700 ;
        RECT 226.950 59.100 229.050 61.200 ;
        RECT 232.950 59.100 235.050 61.200 ;
        RECT 227.400 58.050 228.600 59.100 ;
        RECT 233.400 58.050 234.600 59.100 ;
        RECT 223.950 55.950 226.050 58.050 ;
        RECT 226.950 55.950 229.050 58.050 ;
        RECT 229.950 55.950 232.050 58.050 ;
        RECT 232.950 55.950 235.050 58.050 ;
        RECT 241.950 55.950 244.050 58.050 ;
        RECT 224.400 54.900 225.600 55.950 ;
        RECT 223.950 52.800 226.050 54.900 ;
        RECT 224.400 46.050 225.600 52.800 ;
        RECT 226.950 49.950 229.050 52.050 ;
        RECT 223.950 43.950 226.050 46.050 ;
        RECT 218.400 26.400 222.600 27.600 ;
        RECT 214.950 22.950 217.050 25.050 ;
        RECT 215.400 21.600 216.600 22.950 ;
        RECT 221.400 21.600 222.600 26.400 ;
        RECT 214.950 19.500 217.050 21.600 ;
        RECT 220.950 19.500 223.050 21.600 ;
        RECT 190.950 9.600 193.050 11.700 ;
        RECT 211.950 10.500 214.050 12.600 ;
        RECT 227.400 7.050 228.600 49.950 ;
        RECT 230.400 43.050 231.600 55.950 ;
        RECT 235.950 52.950 238.050 55.050 ;
        RECT 242.400 54.600 243.600 55.950 ;
        RECT 239.400 53.400 243.600 54.600 ;
        RECT 229.950 40.950 232.050 43.050 ;
        RECT 236.400 25.050 237.600 52.950 ;
        RECT 239.400 43.050 240.600 53.400 ;
        RECT 245.850 48.600 247.050 63.600 ;
        RECT 250.950 58.950 253.050 61.050 ;
        RECT 244.950 46.500 247.050 48.600 ;
        RECT 251.400 46.050 252.600 58.950 ;
        RECT 250.950 43.950 253.050 46.050 ;
        RECT 238.950 40.950 241.050 43.050 ;
        RECT 244.950 40.950 247.050 43.050 ;
        RECT 232.950 22.950 235.050 25.050 ;
        RECT 235.950 22.950 238.050 25.050 ;
        RECT 238.950 22.950 241.050 25.050 ;
        RECT 233.400 7.050 234.600 22.950 ;
        RECT 239.400 21.900 240.600 22.950 ;
        RECT 245.400 22.050 246.600 40.950 ;
        RECT 254.400 37.050 255.600 67.950 ;
        RECT 257.400 61.050 258.600 238.950 ;
        RECT 268.950 235.950 271.050 238.050 ;
        RECT 269.400 217.200 270.600 235.950 ;
        RECT 275.400 229.050 276.600 274.950 ;
        RECT 286.950 266.400 289.050 268.500 ;
        RECT 280.950 256.950 283.050 259.050 ;
        RECT 281.400 255.600 282.600 256.950 ;
        RECT 280.950 253.500 283.050 255.600 ;
        RECT 287.100 246.600 288.300 266.400 ;
        RECT 295.950 265.950 298.050 268.050 ;
        RECT 289.950 256.950 292.050 259.050 ;
        RECT 290.400 255.600 291.600 256.950 ;
        RECT 296.400 255.600 297.600 265.950 ;
        RECT 302.400 262.200 303.600 283.950 ;
        RECT 305.400 268.050 306.600 313.950 ;
        RECT 320.400 301.050 321.600 338.400 ;
        RECT 328.950 338.100 331.050 340.200 ;
        RECT 329.400 337.050 330.600 338.100 ;
        RECT 328.950 334.950 331.050 337.050 ;
        RECT 331.950 334.950 334.050 337.050 ;
        RECT 332.400 333.900 333.600 334.950 ;
        RECT 331.950 331.800 334.050 333.900 ;
        RECT 340.950 301.950 343.050 304.050 ;
        RECT 352.950 303.300 355.050 305.400 ;
        RECT 319.950 298.950 322.050 301.050 ;
        RECT 331.950 298.950 334.050 301.050 ;
        RECT 307.950 293.100 310.050 295.200 ;
        RECT 304.950 265.950 307.050 268.050 ;
        RECT 308.400 262.200 309.600 293.100 ;
        RECT 310.950 292.950 313.050 295.050 ;
        RECT 316.950 293.100 319.050 295.200 ;
        RECT 322.950 293.100 325.050 295.200 ;
        RECT 311.400 289.050 312.600 292.950 ;
        RECT 317.400 292.050 318.600 293.100 ;
        RECT 323.400 292.050 324.600 293.100 ;
        RECT 316.950 289.950 319.050 292.050 ;
        RECT 319.950 289.950 322.050 292.050 ;
        RECT 322.950 289.950 325.050 292.050 ;
        RECT 310.950 286.950 313.050 289.050 ;
        RECT 320.400 288.900 321.600 289.950 ;
        RECT 319.950 286.800 322.050 288.900 ;
        RECT 319.950 265.950 322.050 268.050 ;
        RECT 301.950 260.100 304.050 262.200 ;
        RECT 307.950 260.100 310.050 262.200 ;
        RECT 302.400 255.600 303.600 260.100 ;
        RECT 308.400 259.050 309.600 260.100 ;
        RECT 307.950 256.950 310.050 259.050 ;
        RECT 313.950 256.950 316.050 259.050 ;
        RECT 314.400 255.900 315.600 256.950 ;
        RECT 320.400 255.900 321.600 265.950 ;
        RECT 332.400 262.200 333.600 298.950 ;
        RECT 341.400 292.050 342.600 301.950 ;
        RECT 353.850 299.700 355.050 303.300 ;
        RECT 352.950 297.600 355.050 299.700 ;
        RECT 337.950 289.950 340.050 292.050 ;
        RECT 340.950 289.950 343.050 292.050 ;
        RECT 343.950 289.950 346.050 292.050 ;
        RECT 349.950 289.950 352.050 292.050 ;
        RECT 338.400 288.900 339.600 289.950 ;
        RECT 337.950 286.800 340.050 288.900 ;
        RECT 344.400 280.050 345.600 289.950 ;
        RECT 350.400 288.600 351.600 289.950 ;
        RECT 349.950 286.500 352.050 288.600 ;
        RECT 353.850 282.600 355.050 297.600 ;
        RECT 362.400 286.050 363.600 352.950 ;
        RECT 365.400 343.050 366.600 397.950 ;
        RECT 367.950 391.950 370.050 394.050 ;
        RECT 364.950 340.950 367.050 343.050 ;
        RECT 368.400 340.050 369.600 391.950 ;
        RECT 379.950 380.400 382.050 382.500 ;
        RECT 373.950 371.400 376.050 373.500 ;
        RECT 374.400 370.050 375.600 371.400 ;
        RECT 373.950 367.950 376.050 370.050 ;
        RECT 370.950 364.950 373.050 367.050 ;
        RECT 371.400 355.050 372.600 364.950 ;
        RECT 380.100 360.600 381.300 380.400 ;
        RECT 382.950 376.950 385.050 379.050 ;
        RECT 383.400 370.050 384.600 376.950 ;
        RECT 386.400 373.050 387.600 409.950 ;
        RECT 388.950 409.800 391.050 411.900 ;
        RECT 394.950 409.800 397.050 411.900 ;
        RECT 406.950 409.800 409.050 411.900 ;
        RECT 389.400 394.050 390.600 409.800 ;
        RECT 410.400 400.050 411.600 415.950 ;
        RECT 419.400 415.050 420.600 416.100 ;
        RECT 425.400 415.050 426.600 424.800 ;
        RECT 428.400 418.050 429.600 469.950 ;
        RECT 436.950 463.950 439.050 466.050 ;
        RECT 455.400 465.600 456.600 487.800 ;
        RECT 464.400 486.600 465.600 490.950 ;
        RECT 461.400 485.400 465.600 486.600 ;
        RECT 455.400 464.400 459.600 465.600 ;
        RECT 437.400 448.050 438.600 463.950 ;
        RECT 451.950 459.300 454.050 461.400 ;
        RECT 452.850 455.700 454.050 459.300 ;
        RECT 451.950 453.600 454.050 455.700 ;
        RECT 436.950 445.950 439.050 448.050 ;
        RECT 442.950 445.950 445.050 448.050 ;
        RECT 448.950 445.950 451.050 448.050 ;
        RECT 443.400 444.600 444.600 445.950 ;
        RECT 449.400 444.600 450.600 445.950 ;
        RECT 439.950 442.500 442.050 444.600 ;
        RECT 443.400 443.400 447.600 444.600 ;
        RECT 433.950 422.400 436.050 424.500 ;
        RECT 440.400 424.050 441.600 442.500 ;
        RECT 442.950 424.950 445.050 427.050 ;
        RECT 427.950 415.950 430.050 418.050 ;
        RECT 415.950 412.950 418.050 415.050 ;
        RECT 418.950 412.950 421.050 415.050 ;
        RECT 421.950 412.950 424.050 415.050 ;
        RECT 424.950 412.950 427.050 415.050 ;
        RECT 430.950 412.950 433.050 415.050 ;
        RECT 416.400 406.050 417.600 412.950 ;
        RECT 422.400 411.900 423.600 412.950 ;
        RECT 421.950 409.800 424.050 411.900 ;
        RECT 431.400 411.000 432.600 412.950 ;
        RECT 424.950 406.950 427.050 409.050 ;
        RECT 430.950 406.950 433.050 411.000 ;
        RECT 415.950 403.950 418.050 406.050 ;
        RECT 409.950 397.950 412.050 400.050 ;
        RECT 388.950 391.950 391.050 394.050 ;
        RECT 394.950 381.300 397.050 383.400 ;
        RECT 400.950 382.950 403.050 385.050 ;
        RECT 395.850 377.700 397.050 381.300 ;
        RECT 394.950 375.600 397.050 377.700 ;
        RECT 385.950 370.950 388.050 373.050 ;
        RECT 382.950 367.950 385.050 370.050 ;
        RECT 391.950 367.950 394.050 370.050 ;
        RECT 392.400 366.600 393.600 367.950 ;
        RECT 389.400 365.400 393.600 366.600 ;
        RECT 379.950 358.500 382.050 360.600 ;
        RECT 389.400 358.050 390.600 365.400 ;
        RECT 395.850 360.600 397.050 375.600 ;
        RECT 394.950 358.500 397.050 360.600 ;
        RECT 388.950 355.950 391.050 358.050 ;
        RECT 370.950 352.950 373.050 355.050 ;
        RECT 379.950 346.950 382.050 349.050 ;
        RECT 367.950 337.950 370.050 340.050 ;
        RECT 370.950 334.950 373.050 337.050 ;
        RECT 371.400 310.050 372.600 334.950 ;
        RECT 380.400 310.050 381.600 346.950 ;
        RECT 389.400 337.050 390.600 355.950 ;
        RECT 394.950 338.100 397.050 340.200 ;
        RECT 395.400 337.050 396.600 338.100 ;
        RECT 388.950 334.950 391.050 337.050 ;
        RECT 391.950 334.950 394.050 337.050 ;
        RECT 394.950 334.950 397.050 337.050 ;
        RECT 392.400 333.900 393.600 334.950 ;
        RECT 391.950 331.800 394.050 333.900 ;
        RECT 401.400 322.050 402.600 382.950 ;
        RECT 415.950 380.400 418.050 382.500 ;
        RECT 425.400 382.050 426.600 406.950 ;
        RECT 434.700 402.600 435.900 422.400 ;
        RECT 439.950 421.950 442.050 424.050 ;
        RECT 443.400 418.050 444.600 424.950 ;
        RECT 446.400 421.050 447.600 443.400 ;
        RECT 448.950 442.500 451.050 444.600 ;
        RECT 452.850 438.600 454.050 453.600 ;
        RECT 451.950 436.500 454.050 438.600 ;
        RECT 458.400 430.050 459.600 464.400 ;
        RECT 461.400 457.050 462.600 485.400 ;
        RECT 467.700 480.600 468.900 500.400 ;
        RECT 473.400 499.050 474.600 520.950 ;
        RECT 476.400 517.050 477.600 532.950 ;
        RECT 475.950 514.950 478.050 517.050 ;
        RECT 472.950 496.950 475.050 499.050 ;
        RECT 479.400 496.500 480.600 553.950 ;
        RECT 485.400 544.050 486.600 592.950 ;
        RECT 490.950 592.500 493.050 594.600 ;
        RECT 500.400 577.050 501.600 599.400 ;
        RECT 506.400 597.600 507.600 631.950 ;
        RECT 503.400 596.400 507.600 597.600 ;
        RECT 511.950 615.300 514.050 617.400 ;
        RECT 511.950 611.700 513.150 615.300 ;
        RECT 511.950 609.600 514.050 611.700 ;
        RECT 493.950 573.000 496.050 577.050 ;
        RECT 499.950 574.950 502.050 577.050 ;
        RECT 494.400 571.050 495.600 573.000 ;
        RECT 493.950 568.950 496.050 571.050 ;
        RECT 496.950 568.950 499.050 571.050 ;
        RECT 497.400 567.900 498.600 568.950 ;
        RECT 496.950 565.800 499.050 567.900 ;
        RECT 497.400 564.600 498.600 565.800 ;
        RECT 497.400 563.400 501.600 564.600 ;
        RECT 484.950 541.950 487.050 544.050 ;
        RECT 496.950 541.950 499.050 544.050 ;
        RECT 481.950 538.950 484.050 541.050 ;
        RECT 482.400 529.200 483.600 538.950 ;
        RECT 493.950 535.950 496.050 538.050 ;
        RECT 494.400 532.200 495.600 535.950 ;
        RECT 493.950 530.100 496.050 532.200 ;
        RECT 481.950 527.100 484.050 529.200 ;
        RECT 487.950 527.100 490.050 529.200 ;
        RECT 497.400 529.050 498.600 541.950 ;
        RECT 500.400 529.050 501.600 563.400 ;
        RECT 503.400 559.050 504.600 596.400 ;
        RECT 511.950 594.600 513.150 609.600 ;
        RECT 518.400 607.050 519.600 643.800 ;
        RECT 530.400 640.050 531.600 650.100 ;
        RECT 542.400 649.050 543.600 650.100 ;
        RECT 541.950 646.950 544.050 649.050 ;
        RECT 548.400 643.050 549.600 652.950 ;
        RECT 551.400 646.050 552.600 673.950 ;
        RECT 554.400 670.050 555.600 676.800 ;
        RECT 563.400 676.050 564.600 683.100 ;
        RECT 556.950 673.950 559.050 676.050 ;
        RECT 562.950 673.950 565.050 676.050 ;
        RECT 553.950 667.950 556.050 670.050 ;
        RECT 553.950 658.950 556.050 661.050 ;
        RECT 550.950 643.950 553.050 646.050 ;
        RECT 541.950 640.950 544.050 643.050 ;
        RECT 547.950 640.950 550.050 643.050 ;
        RECT 520.950 637.950 523.050 640.050 ;
        RECT 529.950 637.950 532.050 640.050 ;
        RECT 517.950 604.950 520.050 607.050 ;
        RECT 514.950 601.950 517.050 604.050 ;
        RECT 515.400 600.600 516.600 601.950 ;
        RECT 521.400 601.050 522.600 637.950 ;
        RECT 529.950 634.800 532.050 636.900 ;
        RECT 526.950 628.950 529.050 631.050 ;
        RECT 514.950 598.500 517.050 600.600 ;
        RECT 520.950 598.950 523.050 601.050 ;
        RECT 527.400 598.050 528.600 628.950 ;
        RECT 520.950 595.800 523.050 597.900 ;
        RECT 526.950 595.950 529.050 598.050 ;
        RECT 511.950 592.500 514.050 594.600 ;
        RECT 511.950 572.100 514.050 574.200 ;
        RECT 512.400 571.050 513.600 572.100 ;
        RECT 511.950 568.950 514.050 571.050 ;
        RECT 514.950 568.950 517.050 571.050 ;
        RECT 515.400 567.000 516.600 568.950 ;
        RECT 514.950 562.950 517.050 567.000 ;
        RECT 502.950 556.950 505.050 559.050 ;
        RECT 502.950 550.950 505.050 553.050 ;
        RECT 488.400 526.050 489.600 527.100 ;
        RECT 493.950 526.950 496.050 529.050 ;
        RECT 496.950 526.950 499.050 529.050 ;
        RECT 499.950 526.950 502.050 529.050 ;
        RECT 494.400 526.050 495.600 526.950 ;
        RECT 487.950 523.950 490.050 526.050 ;
        RECT 490.950 523.950 493.050 526.050 ;
        RECT 493.950 523.950 496.050 526.050 ;
        RECT 481.950 511.950 484.050 514.050 ;
        RECT 478.950 494.400 481.050 496.500 ;
        RECT 472.950 490.950 475.050 493.050 ;
        RECT 473.400 484.050 474.600 490.950 ;
        RECT 472.950 481.950 475.050 484.050 ;
        RECT 466.950 478.500 469.050 480.600 ;
        RECT 472.950 458.400 475.050 460.500 ;
        RECT 460.950 454.950 463.050 457.050 ;
        RECT 466.950 449.400 469.050 451.500 ;
        RECT 467.400 448.050 468.600 449.400 ;
        RECT 466.950 445.950 469.050 448.050 ;
        RECT 473.100 438.600 474.300 458.400 ;
        RECT 482.400 457.050 483.600 511.950 ;
        RECT 491.400 508.050 492.600 523.950 ;
        RECT 496.950 520.950 499.050 523.050 ;
        RECT 490.950 505.950 493.050 508.050 ;
        RECT 487.950 500.400 490.050 502.500 ;
        RECT 487.950 485.400 489.150 500.400 ;
        RECT 490.950 494.400 493.050 496.500 ;
        RECT 491.400 493.050 492.600 494.400 ;
        RECT 490.950 490.950 493.050 493.050 ;
        RECT 487.950 483.300 490.050 485.400 ;
        RECT 487.950 479.700 489.150 483.300 ;
        RECT 487.950 477.600 490.050 479.700 ;
        RECT 493.950 475.950 496.050 478.050 ;
        RECT 494.400 469.050 495.600 475.950 ;
        RECT 493.950 466.950 496.050 469.050 ;
        RECT 497.400 463.050 498.600 520.950 ;
        RECT 500.400 514.050 501.600 526.950 ;
        RECT 499.950 511.950 502.050 514.050 ;
        RECT 499.950 505.950 502.050 508.050 ;
        RECT 500.400 484.050 501.600 505.950 ;
        RECT 503.400 496.050 504.600 550.950 ;
        RECT 505.950 535.950 508.050 538.050 ;
        RECT 506.400 529.050 507.600 535.950 ;
        RECT 505.950 526.950 508.050 529.050 ;
        RECT 508.950 528.000 511.050 532.050 ;
        RECT 509.400 526.050 510.600 528.000 ;
        RECT 515.400 526.050 516.600 562.950 ;
        RECT 521.400 553.050 522.600 595.800 ;
        RECT 530.400 595.050 531.600 634.800 ;
        RECT 535.950 606.000 538.050 610.050 ;
        RECT 536.400 604.050 537.600 606.000 ;
        RECT 542.400 604.050 543.600 640.950 ;
        RECT 551.400 625.050 552.600 643.950 ;
        RECT 550.950 622.950 553.050 625.050 ;
        RECT 554.400 622.050 555.600 658.950 ;
        RECT 557.400 655.050 558.600 673.950 ;
        RECT 566.400 661.050 567.600 712.950 ;
        RECT 572.400 700.050 573.600 712.950 ;
        RECT 571.950 697.950 574.050 700.050 ;
        RECT 575.400 694.050 576.600 745.950 ;
        RECT 590.400 742.050 591.600 772.950 ;
        RECT 607.950 769.950 610.050 772.050 ;
        RECT 595.950 762.000 598.050 766.050 ;
        RECT 596.400 760.050 597.600 762.000 ;
        RECT 595.950 757.950 598.050 760.050 ;
        RECT 598.950 757.950 601.050 760.050 ;
        RECT 599.400 756.900 600.600 757.950 ;
        RECT 598.950 754.800 601.050 756.900 ;
        RECT 598.950 748.950 601.050 751.050 ;
        RECT 589.950 739.950 592.050 742.050 ;
        RECT 583.950 724.950 586.050 727.050 ;
        RECT 592.950 724.950 595.050 727.050 ;
        RECT 584.400 706.050 585.600 724.950 ;
        RECT 593.400 723.600 594.600 724.950 ;
        RECT 590.400 722.400 594.600 723.600 ;
        RECT 590.400 709.050 591.600 722.400 ;
        RECT 599.400 709.050 600.600 748.950 ;
        RECT 608.400 748.050 609.600 769.950 ;
        RECT 610.950 763.950 613.050 766.050 ;
        RECT 611.400 751.050 612.600 763.950 ;
        RECT 616.950 761.100 619.050 763.200 ;
        RECT 622.950 761.100 625.050 763.200 ;
        RECT 631.950 761.100 634.050 763.200 ;
        RECT 617.400 760.050 618.600 761.100 ;
        RECT 623.400 760.050 624.600 761.100 ;
        RECT 616.950 757.950 619.050 760.050 ;
        RECT 619.950 757.950 622.050 760.050 ;
        RECT 622.950 757.950 625.050 760.050 ;
        RECT 625.950 757.950 628.050 760.050 ;
        RECT 610.950 748.950 613.050 751.050 ;
        RECT 607.950 745.950 610.050 748.050 ;
        RECT 604.950 736.950 607.050 739.050 ;
        RECT 610.950 736.950 613.050 739.050 ;
        RECT 605.400 727.050 606.600 736.950 ;
        RECT 611.400 727.050 612.600 736.950 ;
        RECT 604.950 724.950 607.050 727.050 ;
        RECT 607.950 724.950 610.050 727.050 ;
        RECT 610.950 724.950 613.050 727.050 ;
        RECT 613.950 724.950 616.050 727.050 ;
        RECT 608.400 723.900 609.600 724.950 ;
        RECT 614.400 723.900 615.600 724.950 ;
        RECT 607.950 721.800 610.050 723.900 ;
        RECT 613.950 721.800 616.050 723.900 ;
        RECT 620.400 723.600 621.600 757.950 ;
        RECT 626.400 751.050 627.600 757.950 ;
        RECT 625.950 748.950 628.050 751.050 ;
        RECT 622.950 739.950 625.050 742.050 ;
        RECT 617.400 722.400 621.600 723.600 ;
        RECT 607.950 712.950 610.050 715.050 ;
        RECT 589.950 706.950 592.050 709.050 ;
        RECT 598.950 706.950 601.050 709.050 ;
        RECT 583.950 703.950 586.050 706.050 ;
        RECT 586.950 700.950 589.050 703.050 ;
        RECT 574.950 691.950 577.050 694.050 ;
        RECT 583.950 691.950 586.050 694.050 ;
        RECT 574.950 683.100 577.050 685.200 ;
        RECT 580.950 683.100 583.050 685.200 ;
        RECT 584.400 685.050 585.600 691.950 ;
        RECT 575.400 682.050 576.600 683.100 ;
        RECT 581.400 682.050 582.600 683.100 ;
        RECT 583.950 682.950 586.050 685.050 ;
        RECT 571.950 679.950 574.050 682.050 ;
        RECT 574.950 679.950 577.050 682.050 ;
        RECT 577.950 679.950 580.050 682.050 ;
        RECT 580.950 679.950 583.050 682.050 ;
        RECT 572.400 664.050 573.600 679.950 ;
        RECT 578.400 673.050 579.600 679.950 ;
        RECT 583.950 676.950 586.050 679.050 ;
        RECT 580.950 673.950 583.050 676.050 ;
        RECT 577.950 670.950 580.050 673.050 ;
        RECT 571.950 661.950 574.050 664.050 ;
        RECT 565.950 658.950 568.050 661.050 ;
        RECT 556.950 652.950 559.050 655.050 ;
        RECT 559.950 651.000 562.050 655.050 ;
        RECT 571.950 652.950 574.050 655.050 ;
        RECT 560.400 649.050 561.600 651.000 ;
        RECT 559.950 646.950 562.050 649.050 ;
        RECT 562.950 646.950 565.050 649.050 ;
        RECT 563.400 645.900 564.600 646.950 ;
        RECT 572.400 645.900 573.600 652.950 ;
        RECT 581.400 649.050 582.600 673.950 ;
        RECT 584.400 673.050 585.600 676.950 ;
        RECT 587.400 676.050 588.600 700.950 ;
        RECT 586.950 673.950 589.050 676.050 ;
        RECT 583.950 670.950 586.050 673.050 ;
        RECT 590.400 667.050 591.600 706.950 ;
        RECT 608.400 694.050 609.600 712.950 ;
        RECT 610.950 706.950 613.050 709.050 ;
        RECT 607.950 691.950 610.050 694.050 ;
        RECT 595.950 687.600 598.050 691.050 ;
        RECT 595.950 687.000 600.600 687.600 ;
        RECT 596.400 686.400 600.600 687.000 ;
        RECT 599.400 682.050 600.600 686.400 ;
        RECT 604.950 683.100 607.050 685.200 ;
        RECT 605.400 682.050 606.600 683.100 ;
        RECT 595.950 679.950 598.050 682.050 ;
        RECT 598.950 679.950 601.050 682.050 ;
        RECT 601.950 679.950 604.050 682.050 ;
        RECT 604.950 679.950 607.050 682.050 ;
        RECT 589.950 666.600 592.050 667.050 ;
        RECT 589.950 665.400 594.600 666.600 ;
        RECT 589.950 664.950 592.050 665.400 ;
        RECT 586.950 650.100 589.050 652.200 ;
        RECT 587.400 649.050 588.600 650.100 ;
        RECT 577.950 646.950 580.050 649.050 ;
        RECT 580.950 646.950 583.050 649.050 ;
        RECT 583.950 646.950 586.050 649.050 ;
        RECT 586.950 646.950 589.050 649.050 ;
        RECT 578.400 645.900 579.600 646.950 ;
        RECT 562.950 643.800 565.050 645.900 ;
        RECT 571.950 643.800 574.050 645.900 ;
        RECT 577.950 643.800 580.050 645.900 ;
        RECT 563.400 630.600 564.600 643.800 ;
        RECT 584.400 637.050 585.600 646.950 ;
        RECT 583.950 634.950 586.050 637.050 ;
        RECT 589.950 634.950 592.050 637.050 ;
        RECT 563.400 629.400 567.600 630.600 ;
        RECT 553.950 619.950 556.050 622.050 ;
        RECT 547.950 616.950 550.050 619.050 ;
        RECT 548.400 606.600 549.600 616.950 ;
        RECT 553.950 614.400 556.050 616.500 ;
        RECT 550.950 606.600 553.050 607.500 ;
        RECT 548.400 605.400 553.050 606.600 ;
        RECT 551.400 604.050 552.600 605.400 ;
        RECT 535.950 601.950 538.050 604.050 ;
        RECT 538.950 601.950 541.050 604.050 ;
        RECT 541.950 601.950 544.050 604.050 ;
        RECT 544.950 601.950 547.050 604.050 ;
        RECT 550.950 601.950 553.050 604.050 ;
        RECT 532.950 598.950 535.050 601.050 ;
        RECT 539.400 600.900 540.600 601.950 ;
        RECT 529.950 592.950 532.050 595.050 ;
        RECT 533.400 586.050 534.600 598.950 ;
        RECT 538.950 598.800 541.050 600.900 ;
        RECT 545.400 589.050 546.600 601.950 ;
        RECT 554.700 594.600 555.900 614.400 ;
        RECT 559.950 610.950 562.050 613.050 ;
        RECT 560.400 604.050 561.600 610.950 ;
        RECT 566.400 604.050 567.600 629.400 ;
        RECT 574.950 615.300 577.050 617.400 ;
        RECT 586.950 616.950 589.050 619.050 ;
        RECT 574.950 611.700 576.150 615.300 ;
        RECT 574.950 609.600 577.050 611.700 ;
        RECT 568.950 604.950 571.050 607.050 ;
        RECT 559.950 601.950 562.050 604.050 ;
        RECT 565.950 601.950 568.050 604.050 ;
        RECT 559.950 595.950 562.050 598.050 ;
        RECT 553.950 592.500 556.050 594.600 ;
        RECT 544.950 586.950 547.050 589.050 ;
        RECT 532.950 583.950 535.050 586.050 ;
        RECT 541.950 577.950 544.050 580.050 ;
        RECT 550.950 578.400 553.050 580.500 ;
        RECT 526.950 571.950 529.050 574.050 ;
        RECT 535.950 572.100 538.050 574.200 ;
        RECT 527.400 567.900 528.600 571.950 ;
        RECT 536.400 571.050 537.600 572.100 ;
        RECT 542.400 571.050 543.600 577.950 ;
        RECT 532.950 568.950 535.050 571.050 ;
        RECT 535.950 568.950 538.050 571.050 ;
        RECT 538.950 568.950 541.050 571.050 ;
        RECT 541.950 568.950 544.050 571.050 ;
        RECT 547.950 568.950 550.050 571.050 ;
        RECT 533.400 567.900 534.600 568.950 ;
        RECT 526.950 565.800 529.050 567.900 ;
        RECT 532.950 565.800 535.050 567.900 ;
        RECT 539.400 562.050 540.600 568.950 ;
        RECT 548.400 562.050 549.600 568.950 ;
        RECT 538.950 559.950 541.050 562.050 ;
        RECT 547.950 559.950 550.050 562.050 ;
        RECT 532.950 556.950 535.050 559.050 ;
        RECT 520.800 550.950 522.900 553.050 ;
        RECT 533.400 541.050 534.600 556.950 ;
        RECT 538.950 556.800 541.050 558.900 ;
        RECT 551.700 558.600 552.900 578.400 ;
        RECT 560.400 574.050 561.600 595.950 ;
        RECT 562.950 583.950 565.050 586.050 ;
        RECT 559.950 571.950 562.050 574.050 ;
        RECT 556.950 568.950 559.050 571.050 ;
        RECT 557.400 568.050 558.600 568.950 ;
        RECT 553.950 566.400 558.600 568.050 ;
        RECT 553.950 565.950 558.000 566.400 ;
        RECT 559.950 565.950 562.050 568.050 ;
        RECT 560.400 562.050 561.600 565.950 ;
        RECT 559.950 559.950 562.050 562.050 ;
        RECT 532.950 538.950 535.050 541.050 ;
        RECT 520.950 535.050 523.050 538.050 ;
        RECT 526.950 536.400 529.050 538.500 ;
        RECT 517.950 531.600 520.050 535.050 ;
        RECT 520.950 534.000 526.050 535.050 ;
        RECT 521.400 533.400 526.050 534.000 ;
        RECT 522.000 532.950 526.050 533.400 ;
        RECT 517.950 531.000 522.600 531.600 ;
        RECT 518.400 530.400 522.600 531.000 ;
        RECT 521.400 528.600 522.600 530.400 ;
        RECT 523.950 528.600 526.050 529.500 ;
        RECT 521.400 527.400 526.050 528.600 ;
        RECT 524.400 526.050 525.600 527.400 ;
        RECT 508.950 523.950 511.050 526.050 ;
        RECT 511.950 523.950 514.050 526.050 ;
        RECT 514.950 523.950 517.050 526.050 ;
        RECT 517.950 523.950 520.050 526.050 ;
        RECT 523.950 523.950 526.050 526.050 ;
        RECT 512.400 522.900 513.600 523.950 ;
        RECT 518.400 522.900 519.600 523.950 ;
        RECT 511.950 520.800 514.050 522.900 ;
        RECT 517.950 520.800 520.050 522.900 ;
        RECT 527.700 516.600 528.900 536.400 ;
        RECT 532.950 532.950 535.050 535.050 ;
        RECT 533.400 526.050 534.600 532.950 ;
        RECT 539.400 526.050 540.600 556.800 ;
        RECT 550.950 556.500 553.050 558.600 ;
        RECT 547.950 537.300 550.050 539.400 ;
        RECT 547.950 533.700 549.150 537.300 ;
        RECT 547.950 531.600 550.050 533.700 ;
        RECT 532.950 523.950 535.050 526.050 ;
        RECT 538.950 523.950 541.050 526.050 ;
        RECT 538.950 520.800 541.050 522.900 ;
        RECT 526.950 514.500 529.050 516.600 ;
        RECT 505.950 511.950 508.050 514.050 ;
        RECT 502.950 493.950 505.050 496.050 ;
        RECT 506.400 493.050 507.600 511.950 ;
        RECT 511.950 505.950 514.050 508.050 ;
        RECT 523.950 505.950 526.050 508.050 ;
        RECT 532.950 505.950 535.050 508.050 ;
        RECT 512.400 493.050 513.600 505.950 ;
        RECT 520.950 502.950 523.050 505.050 ;
        RECT 505.950 490.950 508.050 493.050 ;
        RECT 508.950 490.950 511.050 493.050 ;
        RECT 511.950 490.950 514.050 493.050 ;
        RECT 514.950 490.950 517.050 493.050 ;
        RECT 502.950 487.950 505.050 490.050 ;
        RECT 509.400 489.900 510.600 490.950 ;
        RECT 499.950 481.950 502.050 484.050 ;
        RECT 503.400 475.050 504.600 487.950 ;
        RECT 508.950 487.800 511.050 489.900 ;
        RECT 515.400 484.050 516.600 490.950 ;
        RECT 514.950 481.950 517.050 484.050 ;
        RECT 502.950 472.950 505.050 475.050 ;
        RECT 496.950 460.950 499.050 463.050 ;
        RECT 505.950 460.950 508.050 463.050 ;
        RECT 502.950 457.950 505.050 460.050 ;
        RECT 475.950 454.950 478.050 457.050 ;
        RECT 481.950 454.950 484.050 457.050 ;
        RECT 496.950 454.950 499.050 457.050 ;
        RECT 476.400 448.050 477.600 454.950 ;
        RECT 481.950 448.950 484.050 451.050 ;
        RECT 475.950 445.950 478.050 448.050 ;
        RECT 472.950 436.500 475.050 438.600 ;
        RECT 457.950 427.950 460.050 430.050 ;
        RECT 482.400 427.050 483.600 448.950 ;
        RECT 497.400 448.050 498.600 454.950 ;
        RECT 490.950 445.950 493.050 448.050 ;
        RECT 496.950 445.950 499.050 448.050 ;
        RECT 487.950 436.950 490.050 439.050 ;
        RECT 469.950 424.950 472.050 427.050 ;
        RECT 481.950 424.950 484.050 427.050 ;
        RECT 454.950 422.400 457.050 424.500 ;
        RECT 445.950 418.950 448.050 421.050 ;
        RECT 442.950 415.950 445.050 418.050 ;
        RECT 439.950 412.950 442.050 415.050 ;
        RECT 433.950 400.500 436.050 402.600 ;
        RECT 440.400 400.050 441.600 412.950 ;
        RECT 439.950 397.950 442.050 400.050 ;
        RECT 446.400 397.050 447.600 418.950 ;
        RECT 448.950 415.950 451.050 418.050 ;
        RECT 445.950 396.600 448.050 397.050 ;
        RECT 443.400 395.400 448.050 396.600 ;
        RECT 409.950 371.400 412.050 373.500 ;
        RECT 410.400 370.050 411.600 371.400 ;
        RECT 409.950 367.950 412.050 370.050 ;
        RECT 409.950 361.950 412.050 364.050 ;
        RECT 403.950 338.100 406.050 340.200 ;
        RECT 400.950 319.950 403.050 322.050 ;
        RECT 404.400 319.050 405.600 338.100 ;
        RECT 410.400 337.050 411.600 361.950 ;
        RECT 416.100 360.600 417.300 380.400 ;
        RECT 424.950 379.950 427.050 382.050 ;
        RECT 430.950 380.400 433.050 382.500 ;
        RECT 418.950 371.400 421.050 373.500 ;
        RECT 427.950 371.400 430.050 373.500 ;
        RECT 419.400 370.050 420.600 371.400 ;
        RECT 428.400 370.050 429.600 371.400 ;
        RECT 418.950 367.950 421.050 370.050 ;
        RECT 427.950 367.950 430.050 370.050 ;
        RECT 421.950 364.950 424.050 367.050 ;
        RECT 415.950 358.500 418.050 360.600 ;
        RECT 422.400 349.050 423.600 364.950 ;
        RECT 431.700 360.600 432.900 380.400 ;
        RECT 436.950 371.400 439.050 373.500 ;
        RECT 437.400 370.050 438.600 371.400 ;
        RECT 436.950 367.950 439.050 370.050 ;
        RECT 430.950 358.500 433.050 360.600 ;
        RECT 421.950 346.950 424.050 349.050 ;
        RECT 415.950 338.100 418.050 340.200 ;
        RECT 424.950 338.100 427.050 340.200 ;
        RECT 443.400 339.600 444.600 395.400 ;
        RECT 445.950 394.950 448.050 395.400 ;
        RECT 449.400 393.600 450.600 415.950 ;
        RECT 454.950 407.400 456.150 422.400 ;
        RECT 457.950 416.400 460.050 418.500 ;
        RECT 463.950 416.400 466.050 418.500 ;
        RECT 458.400 415.050 459.600 416.400 ;
        RECT 457.950 412.950 460.050 415.050 ;
        RECT 454.950 405.300 457.050 407.400 ;
        RECT 454.950 401.700 456.150 405.300 ;
        RECT 464.400 403.050 465.600 416.400 ;
        RECT 470.400 412.050 471.600 424.950 ;
        RECT 481.950 417.000 484.050 421.050 ;
        RECT 482.400 415.050 483.600 417.000 ;
        RECT 475.950 412.950 478.050 415.050 ;
        RECT 481.950 412.950 484.050 415.050 ;
        RECT 469.950 409.950 472.050 412.050 ;
        RECT 476.400 411.900 477.600 412.950 ;
        RECT 475.950 409.800 478.050 411.900 ;
        RECT 454.950 399.600 457.050 401.700 ;
        RECT 463.950 400.950 466.050 403.050 ;
        RECT 440.400 338.400 444.600 339.600 ;
        RECT 446.400 392.400 450.600 393.600 ;
        RECT 416.400 337.050 417.600 338.100 ;
        RECT 409.950 334.950 412.050 337.050 ;
        RECT 412.950 334.950 415.050 337.050 ;
        RECT 415.950 334.950 418.050 337.050 ;
        RECT 418.950 334.950 421.050 337.050 ;
        RECT 413.400 333.900 414.600 334.950 ;
        RECT 412.950 331.800 415.050 333.900 ;
        RECT 419.400 319.050 420.600 334.950 ;
        RECT 425.400 325.050 426.600 338.100 ;
        RECT 440.400 337.050 441.600 338.400 ;
        RECT 433.950 334.950 436.050 337.050 ;
        RECT 439.950 334.950 442.050 337.050 ;
        RECT 424.950 322.950 427.050 325.050 ;
        RECT 434.400 319.050 435.600 334.950 ;
        RECT 446.400 325.050 447.600 392.400 ;
        RECT 451.950 381.300 454.050 383.400 ;
        RECT 488.400 382.050 489.600 436.950 ;
        RECT 491.400 421.050 492.600 445.950 ;
        RECT 503.400 424.050 504.600 457.950 ;
        RECT 502.950 421.950 505.050 424.050 ;
        RECT 490.950 418.950 493.050 421.050 ;
        RECT 496.950 416.100 499.050 418.200 ;
        RECT 497.400 415.050 498.600 416.100 ;
        RECT 502.950 415.950 505.050 420.900 ;
        RECT 496.950 412.950 499.050 415.050 ;
        RECT 499.950 412.950 502.050 415.050 ;
        RECT 500.400 411.000 501.600 412.950 ;
        RECT 499.950 406.950 502.050 411.000 ;
        RECT 451.950 377.700 453.150 381.300 ;
        RECT 487.950 379.950 490.050 382.050 ;
        RECT 493.950 379.950 496.050 382.050 ;
        RECT 451.950 375.600 454.050 377.700 ;
        RECT 451.950 360.600 453.150 375.600 ;
        RECT 460.950 371.400 463.050 373.500 ;
        RECT 454.950 367.950 457.050 370.050 ;
        RECT 455.400 366.600 456.600 367.950 ;
        RECT 454.950 364.500 457.050 366.600 ;
        RECT 461.400 361.050 462.600 371.400 ;
        RECT 472.950 371.100 475.050 373.200 ;
        RECT 473.400 370.050 474.600 371.100 ;
        RECT 494.400 370.050 495.600 379.950 ;
        RECT 499.950 371.100 502.050 373.200 ;
        RECT 506.400 373.050 507.600 460.950 ;
        RECT 514.950 445.950 517.050 448.050 ;
        RECT 515.400 444.000 516.600 445.950 ;
        RECT 514.950 441.600 517.050 444.000 ;
        RECT 512.400 440.400 517.050 441.600 ;
        RECT 508.950 427.950 511.050 430.050 ;
        RECT 509.400 411.900 510.600 427.950 ;
        RECT 508.950 409.800 511.050 411.900 ;
        RECT 508.950 397.950 511.050 400.050 ;
        RECT 500.400 370.050 501.600 371.100 ;
        RECT 505.950 370.950 508.050 373.050 ;
        RECT 469.950 367.950 472.050 370.050 ;
        RECT 472.950 367.950 475.050 370.050 ;
        RECT 475.950 367.950 478.050 370.050 ;
        RECT 493.950 367.950 496.050 370.050 ;
        RECT 496.950 367.950 499.050 370.050 ;
        RECT 499.950 367.950 502.050 370.050 ;
        RECT 502.950 367.950 505.050 370.050 ;
        RECT 470.400 367.050 471.600 367.950 ;
        RECT 468.000 366.600 471.600 367.050 ;
        RECT 476.400 366.900 477.600 367.950 ;
        RECT 497.400 366.900 498.600 367.950 ;
        RECT 466.950 364.950 471.600 366.600 ;
        RECT 466.950 364.500 469.050 364.950 ;
        RECT 451.950 358.500 454.050 360.600 ;
        RECT 460.950 358.950 463.050 361.050 ;
        RECT 463.950 349.950 466.050 352.050 ;
        RECT 451.950 339.000 454.050 343.050 ;
        RECT 452.400 337.050 453.600 339.000 ;
        RECT 451.950 334.950 454.050 337.050 ;
        RECT 457.950 334.950 460.050 337.050 ;
        RECT 448.950 331.950 451.050 334.050 ;
        RECT 445.950 322.950 448.050 325.050 ;
        RECT 436.950 319.950 439.050 322.050 ;
        RECT 403.950 316.950 406.050 319.050 ;
        RECT 418.950 316.950 421.050 319.050 ;
        RECT 433.950 316.950 436.050 319.050 ;
        RECT 370.950 307.950 373.050 310.050 ;
        RECT 379.950 307.950 382.050 310.050 ;
        RECT 373.950 302.400 376.050 304.500 ;
        RECT 367.950 293.400 370.050 295.500 ;
        RECT 368.400 292.050 369.600 293.400 ;
        RECT 367.950 289.950 370.050 292.050 ;
        RECT 361.950 283.950 364.050 286.050 ;
        RECT 374.100 282.600 375.300 302.400 ;
        RECT 380.400 298.050 381.600 307.950 ;
        RECT 397.950 301.950 400.050 304.050 ;
        RECT 379.950 295.950 382.050 298.050 ;
        RECT 380.400 294.600 381.600 295.950 ;
        RECT 377.400 293.400 381.600 294.600 ;
        RECT 377.400 292.050 378.600 293.400 ;
        RECT 385.950 292.950 388.050 295.050 ;
        RECT 376.950 289.950 379.050 292.050 ;
        RECT 379.950 283.950 382.050 286.050 ;
        RECT 352.950 280.500 355.050 282.600 ;
        RECT 373.950 280.500 376.050 282.600 ;
        RECT 343.950 277.950 346.050 280.050 ;
        RECT 349.950 265.950 352.050 268.050 ;
        RECT 367.950 266.400 370.050 268.500 ;
        RECT 325.950 259.950 328.050 262.050 ;
        RECT 331.950 260.100 334.050 262.200 ;
        RECT 290.400 254.400 294.600 255.600 ;
        RECT 286.950 244.500 289.050 246.600 ;
        RECT 293.400 229.050 294.600 254.400 ;
        RECT 295.950 253.500 298.050 255.600 ;
        RECT 302.400 254.400 306.600 255.600 ;
        RECT 274.950 226.950 277.050 229.050 ;
        RECT 292.950 226.950 295.050 229.050 ;
        RECT 277.950 220.950 280.050 223.050 ;
        RECT 262.950 215.100 265.050 217.200 ;
        RECT 268.950 215.100 271.050 217.200 ;
        RECT 263.400 214.050 264.600 215.100 ;
        RECT 269.400 214.050 270.600 215.100 ;
        RECT 274.950 214.950 277.050 217.050 ;
        RECT 262.950 211.950 265.050 214.050 ;
        RECT 265.950 211.950 268.050 214.050 ;
        RECT 268.950 211.950 271.050 214.050 ;
        RECT 266.400 210.900 267.600 211.950 ;
        RECT 265.950 208.800 268.050 210.900 ;
        RECT 259.950 187.950 262.050 190.050 ;
        RECT 260.400 177.900 261.600 187.950 ;
        RECT 275.400 184.200 276.600 214.950 ;
        RECT 278.400 202.050 279.600 220.950 ;
        RECT 305.400 217.200 306.600 254.400 ;
        RECT 313.950 253.800 316.050 255.900 ;
        RECT 319.950 253.800 322.050 255.900 ;
        RECT 280.950 215.100 283.050 217.200 ;
        RECT 286.950 215.100 289.050 217.200 ;
        RECT 292.950 215.100 295.050 217.200 ;
        RECT 301.800 215.100 303.900 217.200 ;
        RECT 304.950 215.100 307.050 217.200 ;
        RECT 310.950 215.100 313.050 217.200 ;
        RECT 316.950 216.000 319.050 220.050 ;
        RECT 281.400 211.050 282.600 215.100 ;
        RECT 287.400 214.050 288.600 215.100 ;
        RECT 293.400 214.050 294.600 215.100 ;
        RECT 286.950 211.950 289.050 214.050 ;
        RECT 289.950 211.950 292.050 214.050 ;
        RECT 292.950 211.950 295.050 214.050 ;
        RECT 295.950 211.950 298.050 214.050 ;
        RECT 280.950 208.950 283.050 211.050 ;
        RECT 280.950 205.800 283.050 207.900 ;
        RECT 277.950 199.950 280.050 202.050 ;
        RECT 268.950 182.100 271.050 184.200 ;
        RECT 274.950 182.100 277.050 184.200 ;
        RECT 269.400 181.050 270.600 182.100 ;
        RECT 275.400 181.050 276.600 182.100 ;
        RECT 265.950 178.950 268.050 181.050 ;
        RECT 268.950 178.950 271.050 181.050 ;
        RECT 271.950 178.950 274.050 181.050 ;
        RECT 274.950 178.950 277.050 181.050 ;
        RECT 266.400 177.900 267.600 178.950 ;
        RECT 259.950 175.800 262.050 177.900 ;
        RECT 265.950 175.800 268.050 177.900 ;
        RECT 268.950 172.950 271.050 175.050 ;
        RECT 269.400 166.050 270.600 172.950 ;
        RECT 268.950 163.950 271.050 166.050 ;
        RECT 259.950 142.950 262.050 145.050 ;
        RECT 260.400 132.900 261.600 142.950 ;
        RECT 269.400 139.200 270.600 163.950 ;
        RECT 272.400 163.050 273.600 178.950 ;
        RECT 281.400 175.050 282.600 205.800 ;
        RECT 290.400 202.050 291.600 211.950 ;
        RECT 296.400 210.900 297.600 211.950 ;
        RECT 302.400 211.050 303.600 215.100 ;
        RECT 295.950 208.800 298.050 210.900 ;
        RECT 301.950 208.950 304.050 211.050 ;
        RECT 289.950 199.950 292.050 202.050 ;
        RECT 283.950 181.950 286.050 184.050 ;
        RECT 289.950 182.100 292.050 184.200 ;
        RECT 295.950 182.100 298.050 184.200 ;
        RECT 284.400 175.050 285.600 181.950 ;
        RECT 290.400 181.050 291.600 182.100 ;
        RECT 296.400 181.050 297.600 182.100 ;
        RECT 289.950 178.950 292.050 181.050 ;
        RECT 292.950 178.950 295.050 181.050 ;
        RECT 295.950 178.950 298.050 181.050 ;
        RECT 298.950 178.950 301.050 181.050 ;
        RECT 293.400 177.000 294.600 178.950 ;
        RECT 299.400 177.000 300.600 178.950 ;
        RECT 274.950 169.950 277.050 175.050 ;
        RECT 280.950 172.950 283.050 175.050 ;
        RECT 283.950 172.950 286.050 175.050 ;
        RECT 292.950 172.950 295.050 177.000 ;
        RECT 298.950 172.950 301.050 177.000 ;
        RECT 305.400 172.050 306.600 215.100 ;
        RECT 311.400 214.050 312.600 215.100 ;
        RECT 317.400 214.050 318.600 216.000 ;
        RECT 310.950 211.950 313.050 214.050 ;
        RECT 313.950 211.950 316.050 214.050 ;
        RECT 316.950 211.950 319.050 214.050 ;
        RECT 319.950 211.950 322.050 214.050 ;
        RECT 314.400 210.900 315.600 211.950 ;
        RECT 313.950 208.800 316.050 210.900 ;
        RECT 320.400 196.050 321.600 211.950 ;
        RECT 326.400 210.900 327.600 259.950 ;
        RECT 332.400 259.050 333.600 260.100 ;
        RECT 350.400 259.050 351.600 265.950 ;
        RECT 331.950 256.950 334.050 259.050 ;
        RECT 334.950 256.950 337.050 259.050 ;
        RECT 349.950 256.950 352.050 259.050 ;
        RECT 355.950 256.950 358.050 259.050 ;
        RECT 364.950 256.950 367.050 259.050 ;
        RECT 335.400 220.050 336.600 256.950 ;
        RECT 356.400 238.050 357.600 256.950 ;
        RECT 365.400 255.600 366.600 256.950 ;
        RECT 364.950 253.500 367.050 255.600 ;
        RECT 368.700 246.600 369.900 266.400 ;
        RECT 373.950 256.950 376.050 259.050 ;
        RECT 374.400 250.050 375.600 256.950 ;
        RECT 373.950 247.950 376.050 250.050 ;
        RECT 367.950 244.500 370.050 246.600 ;
        RECT 380.400 241.050 381.600 283.950 ;
        RECT 386.400 280.050 387.600 292.950 ;
        RECT 398.400 292.050 399.600 301.950 ;
        RECT 404.400 295.200 405.600 316.950 ;
        RECT 437.400 298.050 438.600 319.950 ;
        RECT 442.950 301.950 445.050 304.050 ;
        RECT 427.950 295.950 430.050 298.050 ;
        RECT 436.950 295.950 439.050 298.050 ;
        RECT 403.950 293.100 406.050 295.200 ;
        RECT 421.950 293.100 424.050 295.200 ;
        RECT 404.400 292.050 405.600 293.100 ;
        RECT 422.400 292.050 423.600 293.100 ;
        RECT 394.950 289.950 397.050 292.050 ;
        RECT 397.950 289.950 400.050 292.050 ;
        RECT 400.950 289.950 403.050 292.050 ;
        RECT 403.950 289.950 406.050 292.050 ;
        RECT 415.950 289.950 418.050 292.050 ;
        RECT 421.950 289.950 424.050 292.050 ;
        RECT 395.400 288.900 396.600 289.950 ;
        RECT 394.950 286.800 397.050 288.900 ;
        RECT 385.950 277.950 388.050 280.050 ;
        RECT 388.950 266.400 391.050 268.500 ;
        RECT 388.950 251.400 390.150 266.400 ;
        RECT 391.950 260.400 394.050 262.500 ;
        RECT 392.400 259.050 393.600 260.400 ;
        RECT 391.950 256.950 394.050 259.050 ;
        RECT 388.950 249.300 391.050 251.400 ;
        RECT 388.950 245.700 390.150 249.300 ;
        RECT 388.950 243.600 391.050 245.700 ;
        RECT 401.400 241.050 402.600 289.950 ;
        RECT 416.400 268.050 417.600 289.950 ;
        RECT 428.400 274.050 429.600 295.950 ;
        RECT 437.400 292.050 438.600 295.950 ;
        RECT 443.400 292.050 444.600 301.950 ;
        RECT 436.950 289.950 439.050 292.050 ;
        RECT 439.950 289.950 442.050 292.050 ;
        RECT 442.950 289.950 445.050 292.050 ;
        RECT 427.950 271.950 430.050 274.050 ;
        RECT 418.950 268.950 421.050 271.050 ;
        RECT 415.950 265.950 418.050 268.050 ;
        RECT 419.400 265.050 420.600 268.950 ;
        RECT 418.950 262.950 421.050 265.050 ;
        RECT 428.400 264.600 429.600 271.950 ;
        RECT 425.400 263.400 429.600 264.600 ;
        RECT 440.400 264.600 441.600 289.950 ;
        RECT 445.950 283.950 448.050 286.050 ;
        RECT 440.400 263.400 444.600 264.600 ;
        RECT 406.950 260.100 409.050 262.200 ;
        RECT 415.950 260.100 418.050 262.200 ;
        RECT 407.400 259.050 408.600 260.100 ;
        RECT 406.950 256.950 409.050 259.050 ;
        RECT 409.950 256.950 412.050 259.050 ;
        RECT 410.400 255.900 411.600 256.950 ;
        RECT 409.950 253.800 412.050 255.900 ;
        RECT 367.950 238.950 370.050 241.050 ;
        RECT 379.950 238.950 382.050 241.050 ;
        RECT 400.950 238.950 403.050 241.050 ;
        RECT 355.950 235.950 358.050 238.050 ;
        RECT 328.950 217.950 331.050 220.050 ;
        RECT 334.950 217.950 337.050 220.050 ;
        RECT 325.950 208.800 328.050 210.900 ;
        RECT 313.950 193.950 316.050 196.050 ;
        RECT 319.950 193.950 322.050 196.050 ;
        RECT 307.950 190.950 310.050 193.050 ;
        RECT 308.400 175.050 309.600 190.950 ;
        RECT 314.400 181.050 315.600 193.950 ;
        RECT 329.400 187.050 330.600 217.950 ;
        RECT 337.950 215.100 340.050 217.200 ;
        RECT 338.400 214.050 339.600 215.100 ;
        RECT 349.950 214.950 352.050 217.050 ;
        RECT 355.950 215.100 358.050 217.200 ;
        RECT 334.950 211.950 337.050 214.050 ;
        RECT 337.950 211.950 340.050 214.050 ;
        RECT 340.950 211.950 343.050 214.050 ;
        RECT 335.400 210.900 336.600 211.950 ;
        RECT 341.400 210.900 342.600 211.950 ;
        RECT 334.950 208.800 337.050 210.900 ;
        RECT 340.950 208.800 343.050 210.900 ;
        RECT 350.400 196.050 351.600 214.950 ;
        RECT 356.400 214.050 357.600 215.100 ;
        RECT 364.950 214.950 367.050 217.050 ;
        RECT 355.950 211.950 358.050 214.050 ;
        RECT 358.950 211.950 361.050 214.050 ;
        RECT 359.400 210.900 360.600 211.950 ;
        RECT 365.400 210.900 366.600 214.950 ;
        RECT 368.400 211.050 369.600 238.950 ;
        RECT 412.950 217.950 415.050 220.050 ;
        RECT 373.950 215.100 376.050 217.200 ;
        RECT 382.950 215.100 385.050 217.200 ;
        RECT 397.950 215.100 400.050 217.200 ;
        RECT 406.950 215.100 409.050 217.200 ;
        RECT 374.400 214.050 375.600 215.100 ;
        RECT 383.400 214.050 384.600 215.100 ;
        RECT 398.400 214.050 399.600 215.100 ;
        RECT 407.400 214.050 408.600 215.100 ;
        RECT 373.950 211.950 376.050 214.050 ;
        RECT 376.950 211.950 379.050 214.050 ;
        RECT 382.950 211.950 385.050 214.050 ;
        RECT 397.950 211.950 400.050 214.050 ;
        RECT 403.950 211.950 406.050 214.050 ;
        RECT 406.950 211.950 409.050 214.050 ;
        RECT 358.950 208.800 361.050 210.900 ;
        RECT 364.800 208.800 366.900 210.900 ;
        RECT 367.950 208.950 370.050 211.050 ;
        RECT 377.400 202.050 378.600 211.950 ;
        RECT 379.950 208.950 382.050 211.050 ;
        RECT 404.400 210.900 405.600 211.950 ;
        RECT 376.950 199.950 379.050 202.050 ;
        RECT 359.400 197.400 366.600 198.600 ;
        RECT 349.950 193.950 352.050 196.050 ;
        RECT 359.400 193.050 360.600 197.400 ;
        RECT 361.950 193.950 364.050 196.050 ;
        RECT 358.950 190.950 361.050 193.050 ;
        RECT 328.950 184.950 331.050 187.050 ;
        RECT 337.500 186.300 339.600 188.400 ;
        RECT 341.400 186.900 342.600 189.450 ;
        RECT 319.950 182.100 322.050 184.200 ;
        RECT 325.950 182.100 328.050 184.200 ;
        RECT 320.400 181.050 321.600 182.100 ;
        RECT 326.400 181.050 327.600 182.100 ;
        RECT 335.400 181.050 336.600 183.600 ;
        RECT 313.950 178.950 316.050 181.050 ;
        RECT 316.950 178.950 319.050 181.050 ;
        RECT 319.950 178.950 322.050 181.050 ;
        RECT 325.950 178.950 328.050 181.050 ;
        RECT 334.950 178.950 337.050 181.050 ;
        RECT 337.950 180.900 338.850 186.300 ;
        RECT 340.800 184.800 342.900 186.900 ;
        RECT 344.700 183.900 346.800 185.700 ;
        RECT 352.950 184.950 355.050 187.050 ;
        RECT 339.750 182.700 348.300 183.900 ;
        RECT 339.750 181.800 341.850 182.700 ;
        RECT 337.950 179.700 344.700 180.900 ;
        RECT 317.400 177.900 318.600 178.950 ;
        RECT 316.950 175.800 319.050 177.900 ;
        RECT 307.950 172.950 310.050 175.050 ;
        RECT 326.400 172.050 327.600 178.950 ;
        RECT 337.950 172.500 339.000 179.700 ;
        RECT 340.800 176.100 342.900 178.200 ;
        RECT 343.800 177.300 344.700 179.700 ;
        RECT 341.400 173.550 342.600 176.100 ;
        RECT 343.800 175.200 345.900 177.300 ;
        RECT 347.400 173.700 348.300 182.700 ;
        RECT 349.500 178.950 351.600 181.050 ;
        RECT 350.400 176.400 351.600 178.950 ;
        RECT 353.400 177.900 354.600 184.950 ;
        RECT 355.950 181.950 361.050 184.050 ;
        RECT 362.400 181.050 363.600 193.950 ;
        RECT 365.400 193.050 366.600 197.400 ;
        RECT 364.950 190.950 367.050 193.050 ;
        RECT 367.950 182.100 370.050 184.200 ;
        RECT 368.400 181.050 369.600 182.100 ;
        RECT 361.950 178.950 364.050 181.050 ;
        RECT 364.950 178.950 367.050 181.050 ;
        RECT 367.950 178.950 370.050 181.050 ;
        RECT 370.950 178.950 373.050 181.050 ;
        RECT 365.400 177.900 366.600 178.950 ;
        RECT 371.400 177.900 372.600 178.950 ;
        RECT 377.400 177.900 378.600 199.950 ;
        RECT 352.950 175.800 355.050 177.900 ;
        RECT 364.950 175.800 367.050 177.900 ;
        RECT 370.950 175.800 373.050 177.900 ;
        RECT 376.950 175.800 379.050 177.900 ;
        RECT 304.950 169.950 307.050 172.050 ;
        RECT 316.950 169.950 319.050 172.050 ;
        RECT 325.950 169.950 328.050 172.050 ;
        RECT 337.500 170.400 339.600 172.500 ;
        RECT 347.100 171.600 349.200 173.700 ;
        RECT 271.950 160.950 274.050 163.050 ;
        RECT 274.950 154.950 277.050 157.050 ;
        RECT 275.400 142.050 276.600 154.950 ;
        RECT 313.950 151.950 316.050 154.050 ;
        RECT 307.950 147.300 310.050 149.400 ;
        RECT 295.950 142.950 298.050 145.050 ;
        RECT 308.850 143.700 310.050 147.300 ;
        RECT 268.950 137.100 271.050 139.200 ;
        RECT 274.950 138.000 277.050 142.050 ;
        RECT 280.950 139.950 283.050 142.050 ;
        RECT 269.400 136.050 270.600 137.100 ;
        RECT 275.400 136.050 276.600 138.000 ;
        RECT 268.950 133.950 271.050 136.050 ;
        RECT 271.950 133.950 274.050 136.050 ;
        RECT 274.950 133.950 277.050 136.050 ;
        RECT 272.400 132.900 273.600 133.950 ;
        RECT 259.950 130.800 262.050 132.900 ;
        RECT 271.950 130.800 274.050 132.900 ;
        RECT 281.400 121.050 282.600 139.950 ;
        RECT 283.950 136.950 286.050 139.050 ;
        RECT 289.950 137.100 292.050 139.200 ;
        RECT 284.400 127.050 285.600 136.950 ;
        RECT 290.400 136.050 291.600 137.100 ;
        RECT 296.400 136.050 297.600 142.950 ;
        RECT 307.950 141.600 310.050 143.700 ;
        RECT 289.950 133.950 292.050 136.050 ;
        RECT 292.950 133.950 295.050 136.050 ;
        RECT 295.950 133.950 298.050 136.050 ;
        RECT 298.950 133.950 301.050 136.050 ;
        RECT 304.950 133.950 307.050 136.050 ;
        RECT 293.400 132.900 294.600 133.950 ;
        RECT 292.950 130.800 295.050 132.900 ;
        RECT 286.950 127.950 289.050 130.050 ;
        RECT 283.950 124.950 286.050 127.050 ;
        RECT 280.950 118.950 283.050 121.050 ;
        RECT 287.400 118.050 288.600 127.950 ;
        RECT 299.400 127.050 300.600 133.950 ;
        RECT 305.400 132.600 306.600 133.950 ;
        RECT 302.400 131.400 306.600 132.600 ;
        RECT 298.950 124.950 301.050 127.050 ;
        RECT 302.400 121.050 303.600 131.400 ;
        RECT 308.850 126.600 310.050 141.600 ;
        RECT 307.950 124.500 310.050 126.600 ;
        RECT 314.400 121.050 315.600 151.950 ;
        RECT 301.950 118.950 304.050 121.050 ;
        RECT 307.950 118.950 310.050 121.050 ;
        RECT 313.950 118.950 316.050 121.050 ;
        RECT 286.950 115.950 289.050 118.050 ;
        RECT 277.950 112.950 280.050 115.050 ;
        RECT 262.950 104.100 265.050 106.200 ;
        RECT 268.950 104.100 271.050 106.200 ;
        RECT 263.400 103.050 264.600 104.100 ;
        RECT 269.400 103.050 270.600 104.100 ;
        RECT 262.950 100.950 265.050 103.050 ;
        RECT 265.950 100.950 268.050 103.050 ;
        RECT 268.950 100.950 271.050 103.050 ;
        RECT 271.950 100.950 274.050 103.050 ;
        RECT 266.400 99.900 267.600 100.950 ;
        RECT 265.950 97.800 268.050 99.900 ;
        RECT 272.400 99.000 273.600 100.950 ;
        RECT 271.950 94.950 274.050 99.000 ;
        RECT 274.950 97.950 277.050 100.050 ;
        RECT 268.950 93.600 271.050 94.050 ;
        RECT 275.400 93.600 276.600 97.950 ;
        RECT 278.400 97.050 279.600 112.950 ;
        RECT 301.950 110.400 304.050 112.500 ;
        RECT 293.400 104.400 300.600 105.600 ;
        RECT 293.400 103.050 294.600 104.400 ;
        RECT 299.400 103.050 300.600 104.400 ;
        RECT 289.950 100.950 292.050 103.050 ;
        RECT 292.950 100.950 295.050 103.050 ;
        RECT 298.950 100.950 301.050 103.050 ;
        RECT 290.400 99.900 291.600 100.950 ;
        RECT 289.950 97.800 292.050 99.900 ;
        RECT 277.950 94.950 280.050 97.050 ;
        RECT 302.850 95.400 304.050 110.400 ;
        RECT 308.400 99.900 309.600 118.950 ;
        RECT 317.400 118.050 318.600 169.950 ;
        RECT 380.400 163.050 381.600 208.950 ;
        RECT 403.950 208.800 406.050 210.900 ;
        RECT 409.950 190.950 412.050 193.050 ;
        RECT 400.950 184.950 403.050 187.050 ;
        RECT 391.950 182.100 394.050 184.200 ;
        RECT 397.950 182.100 400.050 184.200 ;
        RECT 392.400 181.050 393.600 182.100 ;
        RECT 388.950 178.950 391.050 181.050 ;
        RECT 391.950 178.950 394.050 181.050 ;
        RECT 389.400 172.050 390.600 178.950 ;
        RECT 398.400 172.050 399.600 182.100 ;
        RECT 388.950 169.950 391.050 172.050 ;
        RECT 397.950 169.950 400.050 172.050 ;
        RECT 340.950 160.950 346.050 163.050 ;
        RECT 379.950 160.950 382.050 163.050 ;
        RECT 367.950 157.950 370.050 160.050 ;
        RECT 368.400 151.050 369.600 157.950 ;
        RECT 367.950 148.950 370.050 151.050 ;
        RECT 328.950 146.400 331.050 148.500 ;
        RECT 322.950 137.400 325.050 139.500 ;
        RECT 323.400 136.050 324.600 137.400 ;
        RECT 322.950 133.950 325.050 136.050 ;
        RECT 329.100 126.600 330.300 146.400 ;
        RECT 340.950 145.950 343.050 148.050 ;
        RECT 331.950 137.400 334.050 139.500 ;
        RECT 332.400 136.050 333.600 137.400 ;
        RECT 331.950 133.950 334.050 136.050 ;
        RECT 341.400 133.050 342.600 145.950 ;
        RECT 361.950 142.950 364.050 145.050 ;
        RECT 343.950 136.950 346.050 139.050 ;
        RECT 349.950 137.100 352.050 139.200 ;
        RECT 334.950 130.950 337.050 133.050 ;
        RECT 340.950 130.950 343.050 133.050 ;
        RECT 328.950 124.500 331.050 126.600 ;
        RECT 316.950 115.950 319.050 118.050 ;
        RECT 322.950 110.400 325.050 112.500 ;
        RECT 316.950 100.950 319.050 103.050 ;
        RECT 307.950 97.800 310.050 99.900 ;
        RECT 317.400 99.600 318.600 100.950 ;
        RECT 316.950 97.500 319.050 99.600 ;
        RECT 268.950 92.400 276.600 93.600 ;
        RECT 301.950 93.300 304.050 95.400 ;
        RECT 268.950 91.950 271.050 92.400 ;
        RECT 259.950 88.950 262.050 91.050 ;
        RECT 302.850 89.700 304.050 93.300 ;
        RECT 316.950 91.950 319.050 94.050 ;
        RECT 256.950 58.950 259.050 61.050 ;
        RECT 260.400 58.050 261.600 88.950 ;
        RECT 301.950 87.600 304.050 89.700 ;
        RECT 271.950 79.950 274.050 82.050 ;
        RECT 298.950 79.950 301.050 82.050 ;
        RECT 265.950 68.400 268.050 70.500 ;
        RECT 259.950 55.950 262.050 58.050 ;
        RECT 266.100 48.600 267.300 68.400 ;
        RECT 272.400 60.600 273.600 79.950 ;
        RECT 269.400 59.400 273.600 60.600 ;
        RECT 269.400 58.050 270.600 59.400 ;
        RECT 286.950 59.100 289.050 61.200 ;
        RECT 287.400 58.050 288.600 59.100 ;
        RECT 268.950 55.950 271.050 58.050 ;
        RECT 286.950 55.950 289.050 58.050 ;
        RECT 265.950 46.500 268.050 48.600 ;
        RECT 283.950 46.800 286.050 48.900 ;
        RECT 284.400 40.050 285.600 46.800 ;
        RECT 265.950 37.950 268.050 40.050 ;
        RECT 283.800 37.950 285.900 40.050 ;
        RECT 286.950 37.950 289.050 40.050 ;
        RECT 253.950 34.950 256.050 37.050 ;
        RECT 256.950 26.100 259.050 28.200 ;
        RECT 257.400 25.050 258.600 26.100 ;
        RECT 253.950 22.950 256.050 25.050 ;
        RECT 256.950 22.950 259.050 25.050 ;
        RECT 259.950 22.950 262.050 25.050 ;
        RECT 238.950 19.800 241.050 21.900 ;
        RECT 244.950 19.950 247.050 22.050 ;
        RECT 254.400 21.900 255.600 22.950 ;
        RECT 260.400 21.900 261.600 22.950 ;
        RECT 266.400 21.900 267.600 37.950 ;
        RECT 277.950 31.950 280.050 34.050 ;
        RECT 268.950 25.950 271.050 28.050 ;
        RECT 253.950 19.800 256.050 21.900 ;
        RECT 259.950 19.800 262.050 21.900 ;
        RECT 265.950 19.800 268.050 21.900 ;
        RECT 269.400 19.050 270.600 25.950 ;
        RECT 278.400 25.050 279.600 31.950 ;
        RECT 284.400 25.050 285.600 37.950 ;
        RECT 287.400 28.050 288.600 37.950 ;
        RECT 292.950 32.400 295.050 34.500 ;
        RECT 286.950 25.950 289.050 28.050 ;
        RECT 274.950 22.950 277.050 25.050 ;
        RECT 277.950 22.950 280.050 25.050 ;
        RECT 280.950 22.950 283.050 25.050 ;
        RECT 283.950 22.950 286.050 25.050 ;
        RECT 289.950 22.950 292.050 25.050 ;
        RECT 275.400 21.000 276.600 22.950 ;
        RECT 281.400 21.900 282.600 22.950 ;
        RECT 268.950 16.950 271.050 19.050 ;
        RECT 274.950 16.950 277.050 21.000 ;
        RECT 280.950 19.800 283.050 21.900 ;
        RECT 290.400 21.600 291.600 22.950 ;
        RECT 289.950 19.500 292.050 21.600 ;
        RECT 293.700 12.600 294.900 32.400 ;
        RECT 299.400 31.050 300.600 79.950 ;
        RECT 310.950 64.950 313.050 67.050 ;
        RECT 304.950 59.100 307.050 61.200 ;
        RECT 305.400 58.050 306.600 59.100 ;
        RECT 311.400 58.050 312.600 64.950 ;
        RECT 304.950 55.950 307.050 58.050 ;
        RECT 307.950 55.950 310.050 58.050 ;
        RECT 310.950 55.950 313.050 58.050 ;
        RECT 308.400 54.000 309.600 55.950 ;
        RECT 307.950 49.950 310.050 54.000 ;
        RECT 317.400 52.050 318.600 91.950 ;
        RECT 323.100 90.600 324.300 110.400 ;
        RECT 331.950 109.950 334.050 112.050 ;
        RECT 332.400 106.050 333.600 109.950 ;
        RECT 331.950 103.950 334.050 106.050 ;
        RECT 325.950 100.950 328.050 103.050 ;
        RECT 326.400 99.600 327.600 100.950 ;
        RECT 335.400 100.050 336.600 130.950 ;
        RECT 340.950 118.950 343.050 121.050 ;
        RECT 341.400 103.050 342.600 118.950 ;
        RECT 344.400 118.050 345.600 136.950 ;
        RECT 350.400 136.050 351.600 137.100 ;
        RECT 349.950 133.950 352.050 136.050 ;
        RECT 355.950 133.950 358.050 136.050 ;
        RECT 356.400 127.050 357.600 133.950 ;
        RECT 355.950 124.950 358.050 127.050 ;
        RECT 343.950 115.950 346.050 118.050 ;
        RECT 344.400 109.050 345.600 115.950 ;
        RECT 346.950 109.950 349.050 112.050 ;
        RECT 343.950 106.950 346.050 109.050 ;
        RECT 347.400 103.050 348.600 109.950 ;
        RECT 352.950 104.100 355.050 106.200 ;
        RECT 358.950 104.100 361.050 106.200 ;
        RECT 353.400 103.050 354.600 104.100 ;
        RECT 340.950 100.950 343.050 103.050 ;
        RECT 343.950 100.950 346.050 103.050 ;
        RECT 346.950 100.950 349.050 103.050 ;
        RECT 349.950 100.950 352.050 103.050 ;
        RECT 352.950 100.950 355.050 103.050 ;
        RECT 328.950 99.600 331.050 100.050 ;
        RECT 326.400 98.400 331.050 99.600 ;
        RECT 328.950 97.950 331.050 98.400 ;
        RECT 334.950 97.950 337.050 100.050 ;
        RECT 344.400 99.900 345.600 100.950 ;
        RECT 322.950 88.500 325.050 90.600 ;
        RECT 329.400 82.050 330.600 97.950 ;
        RECT 343.950 97.800 346.050 99.900 ;
        RECT 328.950 79.950 331.050 82.050 ;
        RECT 328.950 59.100 331.050 61.200 ;
        RECT 334.950 59.100 337.050 61.200 ;
        RECT 329.400 58.050 330.600 59.100 ;
        RECT 335.400 58.050 336.600 59.100 ;
        RECT 350.400 58.050 351.600 100.950 ;
        RECT 359.400 85.050 360.600 104.100 ;
        RECT 362.400 94.050 363.600 142.950 ;
        RECT 367.950 137.100 370.050 139.200 ;
        RECT 373.950 137.100 376.050 139.200 ;
        RECT 379.950 137.100 382.050 139.200 ;
        RECT 368.400 136.050 369.600 137.100 ;
        RECT 374.400 136.050 375.600 137.100 ;
        RECT 367.950 133.950 370.050 136.050 ;
        RECT 370.950 133.950 373.050 136.050 ;
        RECT 373.950 133.950 376.050 136.050 ;
        RECT 371.400 132.900 372.600 133.950 ;
        RECT 370.950 130.800 373.050 132.900 ;
        RECT 364.950 104.100 367.050 106.200 ;
        RECT 370.950 104.100 373.050 109.050 ;
        RECT 376.950 105.600 379.050 106.200 ;
        RECT 380.400 105.600 381.600 137.100 ;
        RECT 401.400 127.050 402.600 184.950 ;
        RECT 410.400 181.050 411.600 190.950 ;
        RECT 413.400 187.050 414.600 217.950 ;
        RECT 416.400 216.600 417.600 260.100 ;
        RECT 419.400 220.200 420.600 262.950 ;
        RECT 425.400 259.050 426.600 263.400 ;
        RECT 430.950 260.100 433.050 262.200 ;
        RECT 439.950 260.100 442.050 262.200 ;
        RECT 431.400 259.050 432.600 260.100 ;
        RECT 424.950 256.950 427.050 259.050 ;
        RECT 427.950 256.950 430.050 259.050 ;
        RECT 430.950 256.950 433.050 259.050 ;
        RECT 433.950 256.950 436.050 259.050 ;
        RECT 428.400 255.900 429.600 256.950 ;
        RECT 434.400 255.900 435.600 256.950 ;
        RECT 427.950 253.800 430.050 255.900 ;
        RECT 433.950 253.800 436.050 255.900 ;
        RECT 440.400 250.050 441.600 260.100 ;
        RECT 443.400 255.900 444.600 263.400 ;
        RECT 446.400 262.050 447.600 283.950 ;
        RECT 449.400 265.050 450.600 331.950 ;
        RECT 458.400 322.050 459.600 334.950 ;
        RECT 457.950 319.950 460.050 322.050 ;
        RECT 464.400 301.050 465.600 349.950 ;
        RECT 466.950 340.950 469.050 343.050 ;
        RECT 467.400 334.050 468.600 340.950 ;
        RECT 466.950 331.950 469.050 334.050 ;
        RECT 470.400 304.050 471.600 364.950 ;
        RECT 475.950 364.800 478.050 366.900 ;
        RECT 496.950 364.800 499.050 366.900 ;
        RECT 476.400 352.050 477.600 364.800 ;
        RECT 503.400 361.050 504.600 367.950 ;
        RECT 505.950 364.950 508.050 367.050 ;
        RECT 502.950 358.950 505.050 361.050 ;
        RECT 478.950 352.950 481.050 355.050 ;
        RECT 475.950 349.950 478.050 352.050 ;
        RECT 479.400 342.600 480.600 352.950 ;
        RECT 496.950 346.950 499.050 349.050 ;
        RECT 476.400 341.400 480.600 342.600 ;
        RECT 476.400 337.050 477.600 341.400 ;
        RECT 481.950 339.000 484.050 343.050 ;
        RECT 490.950 340.950 493.050 346.050 ;
        RECT 482.400 337.050 483.600 339.000 ;
        RECT 497.400 337.050 498.600 346.950 ;
        RECT 502.950 338.100 505.050 340.200 ;
        RECT 506.400 339.600 507.600 364.950 ;
        RECT 509.400 349.050 510.600 397.950 ;
        RECT 512.400 391.050 513.600 440.400 ;
        RECT 514.950 439.950 517.050 440.400 ;
        RECT 521.400 436.050 522.600 502.950 ;
        RECT 524.400 502.050 525.600 505.950 ;
        RECT 523.950 499.950 526.050 502.050 ;
        RECT 523.950 496.800 526.050 498.900 ;
        RECT 524.400 469.050 525.600 496.800 ;
        RECT 533.400 496.200 534.600 505.950 ;
        RECT 532.950 494.100 535.050 496.200 ;
        RECT 533.400 493.050 534.600 494.100 ;
        RECT 529.950 490.950 532.050 493.050 ;
        RECT 532.950 490.950 535.050 493.050 ;
        RECT 526.950 487.950 529.050 490.050 ;
        RECT 530.400 489.000 531.600 490.950 ;
        RECT 523.950 466.950 526.050 469.050 ;
        RECT 520.950 433.950 523.050 436.050 ;
        RECT 520.950 424.950 523.050 427.050 ;
        RECT 521.400 415.050 522.600 424.950 ;
        RECT 524.400 424.050 525.600 466.950 ;
        RECT 523.950 421.950 526.050 424.050 ;
        RECT 527.400 418.200 528.600 487.950 ;
        RECT 529.950 484.950 532.050 489.000 ;
        RECT 530.400 460.050 531.600 484.950 ;
        RECT 539.400 463.050 540.600 520.800 ;
        RECT 547.950 516.600 549.150 531.600 ;
        RECT 559.950 528.600 562.050 529.050 ;
        RECT 563.400 528.600 564.600 583.950 ;
        RECT 566.400 562.050 567.600 601.950 ;
        RECT 569.400 589.050 570.600 604.950 ;
        RECT 574.950 594.600 576.150 609.600 ;
        RECT 577.950 601.950 580.050 604.050 ;
        RECT 578.400 600.600 579.600 601.950 ;
        RECT 577.950 598.500 580.050 600.600 ;
        RECT 574.950 592.500 577.050 594.600 ;
        RECT 568.950 586.950 571.050 589.050 ;
        RECT 571.950 578.400 574.050 580.500 ;
        RECT 571.950 563.400 573.150 578.400 ;
        RECT 583.950 576.600 586.050 577.050 ;
        RECT 587.400 576.600 588.600 616.950 ;
        RECT 590.400 600.600 591.600 634.950 ;
        RECT 593.400 606.600 594.600 665.400 ;
        RECT 596.400 640.050 597.600 679.950 ;
        RECT 602.400 678.900 603.600 679.950 ;
        RECT 601.950 676.800 604.050 678.900 ;
        RECT 611.400 652.050 612.600 706.950 ;
        RECT 617.400 679.050 618.600 722.400 ;
        RECT 623.400 709.050 624.600 739.950 ;
        RECT 632.400 739.050 633.600 761.100 ;
        RECT 638.400 742.050 639.600 790.800 ;
        RECT 644.400 760.050 645.600 796.800 ;
        RECT 650.400 792.600 651.600 799.950 ;
        RECT 655.950 796.950 658.050 801.900 ;
        RECT 662.400 801.000 663.600 802.950 ;
        RECT 661.950 796.950 664.050 801.000 ;
        RECT 650.400 791.400 654.600 792.600 ;
        RECT 649.950 787.950 652.050 790.050 ;
        RECT 650.400 763.050 651.600 787.950 ;
        RECT 649.950 760.950 652.050 763.050 ;
        RECT 643.950 757.950 646.050 760.050 ;
        RECT 646.950 757.950 649.050 760.050 ;
        RECT 640.950 754.950 643.050 757.050 ;
        RECT 647.400 756.900 648.600 757.950 ;
        RECT 641.400 745.050 642.600 754.950 ;
        RECT 646.950 754.800 649.050 756.900 ;
        RECT 640.950 742.950 643.050 745.050 ;
        RECT 637.950 739.950 640.050 742.050 ;
        RECT 631.950 736.950 634.050 739.050 ;
        RECT 653.400 733.050 654.600 791.400 ;
        RECT 662.400 790.050 663.600 796.950 ;
        RECT 668.400 796.050 669.600 805.950 ;
        RECT 677.400 805.050 678.600 806.100 ;
        RECT 683.400 805.050 684.600 806.100 ;
        RECT 688.950 805.950 691.050 808.050 ;
        RECT 673.950 802.950 676.050 805.050 ;
        RECT 676.950 802.950 679.050 805.050 ;
        RECT 679.950 802.950 682.050 805.050 ;
        RECT 682.950 802.950 685.050 805.050 ;
        RECT 674.400 801.000 675.600 802.950 ;
        RECT 680.400 801.000 681.600 802.950 ;
        RECT 689.400 801.900 690.600 805.950 ;
        RECT 698.400 805.050 699.600 820.950 ;
        RECT 704.400 820.050 705.600 874.950 ;
        RECT 728.400 868.050 729.600 877.800 ;
        RECT 730.950 874.050 733.050 877.050 ;
        RECT 733.950 874.950 736.050 879.000 ;
        RECT 736.950 877.950 739.050 880.050 ;
        RECT 730.800 873.000 733.050 874.050 ;
        RECT 730.800 871.950 732.900 873.000 ;
        RECT 727.950 865.950 730.050 868.050 ;
        RECT 728.400 858.600 729.600 865.950 ;
        RECT 728.400 857.400 732.600 858.600 ;
        RECT 715.950 853.950 718.050 856.050 ;
        RECT 716.400 838.050 717.600 853.950 ;
        RECT 724.950 844.950 727.050 847.050 ;
        RECT 725.400 841.200 726.600 844.950 ;
        RECT 724.950 839.100 727.050 841.200 ;
        RECT 725.400 838.050 726.600 839.100 ;
        RECT 715.950 835.950 718.050 838.050 ;
        RECT 718.950 835.950 721.050 838.050 ;
        RECT 724.950 835.950 727.050 838.050 ;
        RECT 706.950 829.800 709.050 831.900 ;
        RECT 703.950 817.950 706.050 820.050 ;
        RECT 707.400 817.050 708.600 829.800 ;
        RECT 712.950 817.950 715.050 820.050 ;
        RECT 706.950 814.950 709.050 817.050 ;
        RECT 703.950 811.950 706.050 814.050 ;
        RECT 704.400 805.050 705.600 811.950 ;
        RECT 697.950 802.950 700.050 805.050 ;
        RECT 700.950 802.950 703.050 805.050 ;
        RECT 703.950 802.950 706.050 805.050 ;
        RECT 706.950 802.950 709.050 805.050 ;
        RECT 701.400 801.900 702.600 802.950 ;
        RECT 707.400 801.900 708.600 802.950 ;
        RECT 673.950 798.600 676.050 801.000 ;
        RECT 671.400 797.400 676.050 798.600 ;
        RECT 667.950 793.950 670.050 796.050 ;
        RECT 661.950 787.950 664.050 790.050 ;
        RECT 667.950 781.950 670.050 784.050 ;
        RECT 655.950 760.950 658.050 763.050 ;
        RECT 661.950 761.100 664.050 763.200 ;
        RECT 668.400 763.050 669.600 781.950 ;
        RECT 656.400 751.050 657.600 760.950 ;
        RECT 662.400 760.050 663.600 761.100 ;
        RECT 667.950 760.950 670.050 763.050 ;
        RECT 661.950 757.950 664.050 760.050 ;
        RECT 664.950 757.950 667.050 760.050 ;
        RECT 658.950 754.950 661.050 757.050 ;
        RECT 655.950 748.950 658.050 751.050 ;
        RECT 646.950 730.950 649.050 733.050 ;
        RECT 652.950 730.950 655.050 733.050 ;
        RECT 659.400 732.600 660.600 754.950 ;
        RECT 665.400 745.050 666.600 757.950 ;
        RECT 664.950 742.950 667.050 745.050 ;
        RECT 671.400 733.050 672.600 797.400 ;
        RECT 673.950 796.950 676.050 797.400 ;
        RECT 679.950 796.950 682.050 801.000 ;
        RECT 688.950 799.800 691.050 801.900 ;
        RECT 700.950 799.800 703.050 801.900 ;
        RECT 706.950 799.800 709.050 801.900 ;
        RECT 694.950 793.950 697.050 796.050 ;
        RECT 676.950 769.950 679.050 772.050 ;
        RECT 677.400 760.050 678.600 769.950 ;
        RECT 682.950 766.950 685.050 769.050 ;
        RECT 683.400 763.200 684.600 766.950 ;
        RECT 682.950 761.100 685.050 763.200 ;
        RECT 683.400 760.050 684.600 761.100 ;
        RECT 676.950 757.950 679.050 760.050 ;
        RECT 679.950 757.950 682.050 760.050 ;
        RECT 682.950 757.950 685.050 760.050 ;
        RECT 685.950 757.950 688.050 760.050 ;
        RECT 673.950 753.600 676.050 757.050 ;
        RECT 673.950 753.000 678.600 753.600 ;
        RECT 674.400 752.400 678.600 753.000 ;
        RECT 656.400 731.400 660.600 732.600 ;
        RECT 631.950 724.950 634.050 727.050 ;
        RECT 640.950 724.950 643.050 727.050 ;
        RECT 632.400 723.900 633.600 724.950 ;
        RECT 631.950 721.800 634.050 723.900 ;
        RECT 641.400 718.050 642.600 724.950 ;
        RECT 640.950 715.950 643.050 718.050 ;
        RECT 622.950 706.950 625.050 709.050 ;
        RECT 631.950 706.950 634.050 709.050 ;
        RECT 622.950 703.800 625.050 705.900 ;
        RECT 623.400 685.200 624.600 703.800 ;
        RECT 632.400 694.050 633.600 706.950 ;
        RECT 640.950 694.950 643.050 697.050 ;
        RECT 631.950 691.950 634.050 694.050 ;
        RECT 622.950 683.100 625.050 685.200 ;
        RECT 623.400 682.050 624.600 683.100 ;
        RECT 632.400 682.050 633.600 691.950 ;
        RECT 641.400 685.050 642.600 694.950 ;
        RECT 647.400 691.050 648.600 730.950 ;
        RECT 656.400 727.050 657.600 731.400 ;
        RECT 670.950 730.950 673.050 733.050 ;
        RECT 677.400 727.050 678.600 752.400 ;
        RECT 680.400 751.050 681.600 757.950 ;
        RECT 679.950 748.950 682.050 751.050 ;
        RECT 686.400 748.050 687.600 757.950 ;
        RECT 695.400 756.900 696.600 793.950 ;
        RECT 713.400 775.050 714.600 817.950 ;
        RECT 719.400 817.050 720.600 835.950 ;
        RECT 731.400 834.600 732.600 857.400 ;
        RECT 733.950 855.600 736.050 856.050 ;
        RECT 737.400 855.600 738.600 877.950 ;
        RECT 740.400 874.050 741.600 883.950 ;
        RECT 749.400 883.050 750.600 884.100 ;
        RECT 755.400 883.050 756.600 884.100 ;
        RECT 748.950 880.950 751.050 883.050 ;
        RECT 751.950 880.950 754.050 883.050 ;
        RECT 754.950 880.950 757.050 883.050 ;
        RECT 757.950 880.950 760.050 883.050 ;
        RECT 752.400 879.900 753.600 880.950 ;
        RECT 751.950 877.800 754.050 879.900 ;
        RECT 758.400 879.000 759.600 880.950 ;
        RECT 739.950 871.950 742.050 874.050 ;
        RECT 733.950 854.400 738.600 855.600 ;
        RECT 733.950 853.950 736.050 854.400 ;
        RECT 734.400 835.050 735.600 853.950 ;
        RECT 742.950 840.000 745.050 844.050 ;
        RECT 743.400 838.050 744.600 840.000 ;
        RECT 748.950 839.100 751.050 841.200 ;
        RECT 752.400 841.050 753.600 877.800 ;
        RECT 757.950 874.950 760.050 879.000 ;
        RECT 764.400 871.050 765.600 884.100 ;
        RECT 773.400 883.050 774.600 884.100 ;
        RECT 779.400 883.050 780.600 892.950 ;
        RECT 820.950 889.950 823.050 892.050 ;
        RECT 886.950 889.950 889.050 892.050 ;
        RECT 790.950 884.100 793.050 886.200 ;
        RECT 799.950 884.100 802.050 886.200 ;
        RECT 805.950 884.100 808.050 886.200 ;
        RECT 811.950 884.100 814.050 886.200 ;
        RECT 769.950 880.950 772.050 883.050 ;
        RECT 772.950 880.950 775.050 883.050 ;
        RECT 775.950 880.950 778.050 883.050 ;
        RECT 778.950 880.950 781.050 883.050 ;
        RECT 770.400 879.900 771.600 880.950 ;
        RECT 776.400 879.900 777.600 880.950 ;
        RECT 769.950 877.800 772.050 879.900 ;
        RECT 775.950 874.950 778.050 879.900 ;
        RECT 763.950 868.950 766.050 871.050 ;
        RECT 772.950 868.950 775.050 871.050 ;
        RECT 749.400 838.050 750.600 839.100 ;
        RECT 751.950 838.950 754.050 841.050 ;
        RECT 754.950 839.100 757.050 844.050 ;
        RECT 760.950 839.100 763.050 841.200 ;
        RECT 766.950 839.100 769.050 841.200 ;
        RECT 773.400 841.050 774.600 868.950 ;
        RECT 739.950 835.950 742.050 838.050 ;
        RECT 742.950 835.950 745.050 838.050 ;
        RECT 745.950 835.950 748.050 838.050 ;
        RECT 748.950 835.950 751.050 838.050 ;
        RECT 728.400 833.400 732.600 834.600 ;
        RECT 718.950 814.950 721.050 817.050 ;
        RECT 728.400 805.050 729.600 833.400 ;
        RECT 733.950 832.950 736.050 835.050 ;
        RECT 740.400 834.900 741.600 835.950 ;
        RECT 739.950 832.800 742.050 834.900 ;
        RECT 746.400 814.050 747.600 835.950 ;
        RECT 751.950 832.950 754.050 835.050 ;
        RECT 748.950 826.950 751.050 829.050 ;
        RECT 749.400 820.050 750.600 826.950 ;
        RECT 752.400 825.600 753.600 832.950 ;
        RECT 755.400 829.050 756.600 839.100 ;
        RECT 761.400 838.050 762.600 839.100 ;
        RECT 767.400 838.050 768.600 839.100 ;
        RECT 772.950 838.950 775.050 841.050 ;
        RECT 760.950 835.950 763.050 838.050 ;
        RECT 763.950 835.950 766.050 838.050 ;
        RECT 766.950 835.950 769.050 838.050 ;
        RECT 769.950 835.950 772.050 838.050 ;
        RECT 764.400 834.900 765.600 835.950 ;
        RECT 770.400 834.900 771.600 835.950 ;
        RECT 776.400 835.050 777.600 874.950 ;
        RECT 791.400 874.050 792.600 884.100 ;
        RECT 800.400 883.050 801.600 884.100 ;
        RECT 796.950 880.950 799.050 883.050 ;
        RECT 799.950 880.950 802.050 883.050 ;
        RECT 797.400 879.900 798.600 880.950 ;
        RECT 796.950 877.800 799.050 879.900 ;
        RECT 790.950 871.950 793.050 874.050 ;
        RECT 806.400 856.050 807.600 884.100 ;
        RECT 812.400 883.050 813.600 884.100 ;
        RECT 811.950 880.950 814.050 883.050 ;
        RECT 814.950 880.950 817.050 883.050 ;
        RECT 815.400 879.900 816.600 880.950 ;
        RECT 814.950 877.800 817.050 879.900 ;
        RECT 793.950 853.950 796.050 856.050 ;
        RECT 805.950 853.950 808.050 856.050 ;
        RECT 787.950 839.100 790.050 841.200 ;
        RECT 788.400 838.050 789.600 839.100 ;
        RECT 794.400 838.050 795.600 853.950 ;
        RECT 799.950 844.950 802.050 847.050 ;
        RECT 784.950 835.950 787.050 838.050 ;
        RECT 787.950 835.950 790.050 838.050 ;
        RECT 790.950 835.950 793.050 838.050 ;
        RECT 793.950 835.950 796.050 838.050 ;
        RECT 763.950 832.800 766.050 834.900 ;
        RECT 769.950 832.800 772.050 834.900 ;
        RECT 775.950 832.950 778.050 835.050 ;
        RECT 785.400 834.900 786.600 835.950 ;
        RECT 791.400 834.900 792.600 835.950 ;
        RECT 800.400 835.050 801.600 844.950 ;
        RECT 821.400 841.200 822.600 889.950 ;
        RECT 847.950 886.950 850.050 889.050 ;
        RECT 823.950 884.100 826.050 886.200 ;
        RECT 832.950 884.100 835.050 886.200 ;
        RECT 838.950 884.100 841.050 886.200 ;
        RECT 824.400 868.050 825.600 884.100 ;
        RECT 833.400 883.050 834.600 884.100 ;
        RECT 839.400 883.050 840.600 884.100 ;
        RECT 844.950 883.950 847.050 886.050 ;
        RECT 829.950 880.950 832.050 883.050 ;
        RECT 832.950 880.950 835.050 883.050 ;
        RECT 835.950 880.950 838.050 883.050 ;
        RECT 838.950 880.950 841.050 883.050 ;
        RECT 830.400 874.050 831.600 880.950 ;
        RECT 836.400 879.900 837.600 880.950 ;
        RECT 835.950 877.800 838.050 879.900 ;
        RECT 829.950 871.950 832.050 874.050 ;
        RECT 823.950 865.950 826.050 868.050 ;
        RECT 845.400 850.050 846.600 883.950 ;
        RECT 848.400 879.600 849.600 886.950 ;
        RECT 853.950 885.000 856.050 889.050 ;
        RECT 854.400 883.050 855.600 885.000 ;
        RECT 859.950 884.100 862.050 886.200 ;
        RECT 860.400 883.050 861.600 884.100 ;
        RECT 871.950 883.950 874.050 886.050 ;
        RECT 880.950 884.100 883.050 886.200 ;
        RECT 853.950 880.950 856.050 883.050 ;
        RECT 856.950 880.950 859.050 883.050 ;
        RECT 859.950 880.950 862.050 883.050 ;
        RECT 862.950 880.950 865.050 883.050 ;
        RECT 848.400 878.400 852.600 879.600 ;
        RECT 835.950 847.950 838.050 850.050 ;
        RECT 844.950 847.950 847.050 850.050 ;
        RECT 808.950 839.100 811.050 841.200 ;
        RECT 814.950 839.100 817.050 841.200 ;
        RECT 820.950 839.100 823.050 841.200 ;
        RECT 809.400 838.050 810.600 839.100 ;
        RECT 815.400 838.050 816.600 839.100 ;
        RECT 836.400 838.050 837.600 847.950 ;
        RECT 841.950 839.100 844.050 841.200 ;
        RECT 842.400 838.050 843.600 839.100 ;
        RECT 808.950 835.950 811.050 838.050 ;
        RECT 811.950 835.950 814.050 838.050 ;
        RECT 814.950 835.950 817.050 838.050 ;
        RECT 817.950 835.950 820.050 838.050 ;
        RECT 835.950 835.950 838.050 838.050 ;
        RECT 838.950 835.950 841.050 838.050 ;
        RECT 841.950 835.950 844.050 838.050 ;
        RECT 844.950 835.950 847.050 838.050 ;
        RECT 784.950 832.800 787.050 834.900 ;
        RECT 790.950 832.800 793.050 834.900 ;
        RECT 799.950 832.950 802.050 835.050 ;
        RECT 764.400 831.600 765.600 832.800 ;
        RECT 761.400 830.400 765.600 831.600 ;
        RECT 754.950 826.950 757.050 829.050 ;
        RECT 752.400 824.400 756.600 825.600 ;
        RECT 748.950 817.950 751.050 820.050 ;
        RECT 745.950 811.950 748.050 814.050 ;
        RECT 733.950 806.100 736.050 808.200 ;
        RECT 734.400 805.050 735.600 806.100 ;
        RECT 749.400 805.050 750.600 817.950 ;
        RECT 755.400 805.050 756.600 824.400 ;
        RECT 724.950 802.950 727.050 805.050 ;
        RECT 727.950 802.950 730.050 805.050 ;
        RECT 730.950 802.950 733.050 805.050 ;
        RECT 733.950 802.950 736.050 805.050 ;
        RECT 745.950 802.950 748.050 805.050 ;
        RECT 748.950 802.950 751.050 805.050 ;
        RECT 751.950 802.950 754.050 805.050 ;
        RECT 754.950 802.950 757.050 805.050 ;
        RECT 725.400 796.050 726.600 802.950 ;
        RECT 724.950 793.950 727.050 796.050 ;
        RECT 725.400 787.050 726.600 793.950 ;
        RECT 731.400 787.050 732.600 802.950 ;
        RECT 746.400 801.900 747.600 802.950 ;
        RECT 745.950 799.800 748.050 801.900 ;
        RECT 752.400 796.050 753.600 802.950 ;
        RECT 761.400 801.900 762.600 830.400 ;
        RECT 766.950 829.950 769.050 832.050 ;
        RECT 767.400 814.050 768.600 829.950 ;
        RECT 775.950 829.800 778.050 831.900 ;
        RECT 766.950 811.950 769.050 814.050 ;
        RECT 760.950 799.800 763.050 801.900 ;
        RECT 767.400 801.600 768.600 811.950 ;
        RECT 776.400 805.050 777.600 829.800 ;
        RECT 812.400 823.050 813.600 835.950 ;
        RECT 811.950 820.950 814.050 823.050 ;
        RECT 796.950 817.950 799.050 820.050 ;
        RECT 781.950 806.100 784.050 808.200 ;
        RECT 790.950 806.100 793.050 808.200 ;
        RECT 782.400 805.050 783.600 806.100 ;
        RECT 772.950 802.950 775.050 805.050 ;
        RECT 775.950 802.950 778.050 805.050 ;
        RECT 778.950 802.950 781.050 805.050 ;
        RECT 781.950 802.950 784.050 805.050 ;
        RECT 773.400 801.600 774.600 802.950 ;
        RECT 767.400 800.400 774.600 801.600 ;
        RECT 751.950 793.950 754.050 796.050 ;
        RECT 724.950 784.950 727.050 787.050 ;
        RECT 730.950 784.950 733.050 787.050 ;
        RECT 718.950 775.950 721.050 778.050 ;
        RECT 712.950 772.950 715.050 775.050 ;
        RECT 706.950 766.950 712.050 769.050 ;
        RECT 715.950 766.950 718.050 772.050 ;
        RECT 697.950 761.100 700.050 763.200 ;
        RECT 706.950 761.100 709.050 763.200 ;
        RECT 712.950 762.000 715.050 766.050 ;
        RECT 694.950 754.800 697.050 756.900 ;
        RECT 688.950 751.950 691.050 754.050 ;
        RECT 685.950 745.950 688.050 748.050 ;
        RECT 689.400 745.050 690.600 751.950 ;
        RECT 698.400 751.050 699.600 761.100 ;
        RECT 707.400 760.050 708.600 761.100 ;
        RECT 713.400 760.050 714.600 762.000 ;
        RECT 703.950 757.950 706.050 760.050 ;
        RECT 706.950 757.950 709.050 760.050 ;
        RECT 709.950 757.950 712.050 760.050 ;
        RECT 712.950 757.950 715.050 760.050 ;
        RECT 704.400 756.900 705.600 757.950 ;
        RECT 710.400 756.900 711.600 757.950 ;
        RECT 703.950 754.800 706.050 756.900 ;
        RECT 709.950 754.800 712.050 756.900 ;
        RECT 697.950 748.950 700.050 751.050 ;
        RECT 688.950 742.950 691.050 745.050 ;
        RECT 710.400 742.050 711.600 754.800 ;
        RECT 719.400 754.050 720.600 775.950 ;
        RECT 748.950 769.950 751.050 772.050 ;
        RECT 724.950 761.100 727.050 763.200 ;
        RECT 730.950 761.100 733.050 766.050 ;
        RECT 742.950 761.100 745.050 763.200 ;
        RECT 725.400 760.050 726.600 761.100 ;
        RECT 731.400 760.050 732.600 761.100 ;
        RECT 724.950 757.950 727.050 760.050 ;
        RECT 727.950 757.950 730.050 760.050 ;
        RECT 730.950 757.950 733.050 760.050 ;
        RECT 733.950 757.950 736.050 760.050 ;
        RECT 739.950 757.950 742.050 760.050 ;
        RECT 728.400 756.000 729.600 757.950 ;
        RECT 712.950 751.950 715.050 754.050 ;
        RECT 718.950 751.950 721.050 754.050 ;
        RECT 727.950 751.950 730.050 756.000 ;
        RECT 734.400 754.050 735.600 757.950 ;
        RECT 730.950 752.400 735.600 754.050 ;
        RECT 730.950 751.950 735.000 752.400 ;
        RECT 736.950 751.950 739.050 754.050 ;
        RECT 709.950 739.950 712.050 742.050 ;
        RECT 682.950 728.100 685.050 730.200 ;
        RECT 691.950 728.100 694.050 730.200 ;
        RECT 700.950 728.100 703.050 730.200 ;
        RECT 706.950 729.000 709.050 733.050 ;
        RECT 683.400 727.050 684.600 728.100 ;
        RECT 652.950 724.950 655.050 727.050 ;
        RECT 655.950 724.950 658.050 727.050 ;
        RECT 658.950 724.950 661.050 727.050 ;
        RECT 676.950 724.950 679.050 727.050 ;
        RECT 679.950 724.950 682.050 727.050 ;
        RECT 682.950 724.950 685.050 727.050 ;
        RECT 685.950 724.950 688.050 727.050 ;
        RECT 653.400 723.900 654.600 724.950 ;
        RECT 652.950 721.800 655.050 723.900 ;
        RECT 652.950 715.950 655.050 718.050 ;
        RECT 653.400 699.600 654.600 715.950 ;
        RECT 655.950 706.950 658.050 709.050 ;
        RECT 656.400 702.600 657.600 706.950 ;
        RECT 659.400 706.050 660.600 724.950 ;
        RECT 680.400 718.050 681.600 724.950 ;
        RECT 686.400 723.000 687.600 724.950 ;
        RECT 685.950 720.600 688.050 723.000 ;
        RECT 685.950 719.400 690.600 720.600 ;
        RECT 685.950 718.950 688.050 719.400 ;
        RECT 679.950 715.950 682.050 718.050 ;
        RECT 658.800 703.950 660.900 706.050 ;
        RECT 661.950 702.600 664.050 706.050 ;
        RECT 656.400 702.000 664.050 702.600 ;
        RECT 656.400 701.400 663.600 702.000 ;
        RECT 653.400 698.400 657.600 699.600 ;
        RECT 646.950 688.950 649.050 691.050 ;
        RECT 652.950 688.950 655.050 691.050 ;
        RECT 648.000 687.600 652.050 688.050 ;
        RECT 647.400 685.950 652.050 687.600 ;
        RECT 640.950 682.950 643.050 685.050 ;
        RECT 647.400 682.050 648.600 685.950 ;
        RECT 653.400 685.050 654.600 688.950 ;
        RECT 652.950 682.950 655.050 685.050 ;
        RECT 622.950 679.950 625.050 682.050 ;
        RECT 631.950 679.950 634.050 682.050 ;
        RECT 643.950 679.950 646.050 682.050 ;
        RECT 646.950 679.950 649.050 682.050 ;
        RECT 649.950 679.950 652.050 682.050 ;
        RECT 616.950 676.950 619.050 679.050 ;
        RECT 634.950 676.950 637.050 679.050 ;
        RECT 644.400 678.900 645.600 679.950 ;
        RECT 622.950 661.950 625.050 664.050 ;
        RECT 616.950 652.950 619.050 655.050 ;
        RECT 610.950 649.950 613.050 652.050 ;
        RECT 617.400 649.050 618.600 652.950 ;
        RECT 623.400 649.050 624.600 661.950 ;
        RECT 628.950 651.000 631.050 655.050 ;
        RECT 635.400 652.050 636.600 676.950 ;
        RECT 643.950 676.800 646.050 678.900 ;
        RECT 650.400 673.050 651.600 679.950 ;
        RECT 652.950 676.950 655.050 679.050 ;
        RECT 649.950 670.950 652.050 673.050 ;
        RECT 637.950 652.950 640.050 655.050 ;
        RECT 629.400 649.050 630.600 651.000 ;
        RECT 634.950 649.950 637.050 652.050 ;
        RECT 638.400 649.050 639.600 652.950 ;
        RECT 650.400 649.050 651.600 670.950 ;
        RECT 653.400 661.050 654.600 676.950 ;
        RECT 652.950 658.950 655.050 661.050 ;
        RECT 656.400 652.050 657.600 698.400 ;
        RECT 655.950 649.950 658.050 652.050 ;
        RECT 601.950 646.950 604.050 649.050 ;
        RECT 616.950 646.950 619.050 649.050 ;
        RECT 622.950 646.950 625.050 649.050 ;
        RECT 625.950 646.950 628.050 649.050 ;
        RECT 628.950 646.950 631.050 649.050 ;
        RECT 631.950 646.950 634.050 649.050 ;
        RECT 637.950 646.950 640.050 649.050 ;
        RECT 646.950 646.950 649.050 649.050 ;
        RECT 649.950 646.950 652.050 649.050 ;
        RECT 652.950 646.950 655.050 649.050 ;
        RECT 598.950 643.950 601.050 646.050 ;
        RECT 595.950 637.950 598.050 640.050 ;
        RECT 599.400 619.050 600.600 643.950 ;
        RECT 602.400 640.050 603.600 646.950 ;
        RECT 610.950 643.950 613.050 646.050 ;
        RECT 626.400 645.900 627.600 646.950 ;
        RECT 601.950 637.950 604.050 640.050 ;
        RECT 607.950 625.950 610.050 628.050 ;
        RECT 598.950 616.950 601.050 619.050 ;
        RECT 593.400 605.400 597.600 606.600 ;
        RECT 596.400 604.050 597.600 605.400 ;
        RECT 601.950 605.100 604.050 607.200 ;
        RECT 602.400 604.050 603.600 605.100 ;
        RECT 595.950 601.950 598.050 604.050 ;
        RECT 598.950 601.950 601.050 604.050 ;
        RECT 601.950 601.950 604.050 604.050 ;
        RECT 599.400 600.900 600.600 601.950 ;
        RECT 590.400 599.400 594.600 600.600 ;
        RECT 590.400 592.050 591.600 599.400 ;
        RECT 589.950 589.950 592.050 592.050 ;
        RECT 593.400 589.050 594.600 599.400 ;
        RECT 598.950 598.800 601.050 600.900 ;
        RECT 604.950 598.950 607.050 601.050 ;
        RECT 592.950 586.950 595.050 589.050 ;
        RECT 583.950 575.400 588.600 576.600 ;
        RECT 583.950 574.950 586.050 575.400 ;
        RECT 574.950 572.400 577.050 574.500 ;
        RECT 575.400 571.050 576.600 572.400 ;
        RECT 574.950 568.950 577.050 571.050 ;
        RECT 584.400 567.900 585.600 574.950 ;
        RECT 589.950 572.100 592.050 574.200 ;
        RECT 605.400 573.600 606.600 598.950 ;
        RECT 608.400 577.050 609.600 625.950 ;
        RECT 611.400 612.600 612.600 643.950 ;
        RECT 625.950 643.800 628.050 645.900 ;
        RECT 632.400 645.000 633.600 646.950 ;
        RECT 631.950 640.950 634.050 645.000 ;
        RECT 632.400 628.050 633.600 640.950 ;
        RECT 638.400 640.050 639.600 646.950 ;
        RECT 643.950 640.950 646.050 646.050 ;
        RECT 647.400 640.050 648.600 646.950 ;
        RECT 653.400 645.900 654.600 646.950 ;
        RECT 652.950 643.800 655.050 645.900 ;
        RECT 655.950 643.950 658.050 646.050 ;
        RECT 637.950 637.950 640.050 640.050 ;
        RECT 646.950 637.950 649.050 640.050 ;
        RECT 631.950 625.950 634.050 628.050 ;
        RECT 647.400 625.050 648.600 637.950 ;
        RECT 646.950 622.950 649.050 625.050 ;
        RECT 634.950 619.950 637.050 622.050 ;
        RECT 622.950 616.950 625.050 619.050 ;
        RECT 631.950 616.950 634.050 619.050 ;
        RECT 611.400 611.400 615.600 612.600 ;
        RECT 610.950 607.950 613.050 610.050 ;
        RECT 611.400 601.050 612.600 607.950 ;
        RECT 614.400 607.050 615.600 611.400 ;
        RECT 613.950 604.950 616.050 607.050 ;
        RECT 616.950 606.000 619.050 610.050 ;
        RECT 617.400 604.050 618.600 606.000 ;
        RECT 623.400 604.050 624.600 616.950 ;
        RECT 628.950 605.100 631.050 610.050 ;
        RECT 616.950 601.950 619.050 604.050 ;
        RECT 619.950 601.950 622.050 604.050 ;
        RECT 622.950 601.950 625.050 604.050 ;
        RECT 625.950 601.950 628.050 604.050 ;
        RECT 610.950 598.950 613.050 601.050 ;
        RECT 616.950 592.950 619.050 595.050 ;
        RECT 607.950 574.950 610.050 577.050 ;
        RECT 602.400 572.400 606.600 573.600 ;
        RECT 590.400 571.050 591.600 572.100 ;
        RECT 589.950 568.950 592.050 571.050 ;
        RECT 592.950 568.950 595.050 571.050 ;
        RECT 593.400 567.900 594.600 568.950 ;
        RECT 583.950 565.800 586.050 567.900 ;
        RECT 592.950 565.800 595.050 567.900 ;
        RECT 565.950 559.950 568.050 562.050 ;
        RECT 571.950 561.300 574.050 563.400 ;
        RECT 577.950 562.950 580.050 565.050 ;
        RECT 571.950 557.700 573.150 561.300 ;
        RECT 571.950 555.600 574.050 557.700 ;
        RECT 578.400 541.050 579.600 562.950 ;
        RECT 577.950 538.950 580.050 541.050 ;
        RECT 578.400 531.600 579.600 538.950 ;
        RECT 578.400 530.400 582.600 531.600 ;
        RECT 559.950 527.400 564.600 528.600 ;
        RECT 559.950 526.950 562.050 527.400 ;
        RECT 568.950 527.100 571.050 529.200 ;
        RECT 576.000 528.600 580.050 529.050 ;
        RECT 550.950 523.950 553.050 526.050 ;
        RECT 551.400 522.600 552.600 523.950 ;
        RECT 550.950 520.500 553.050 522.600 ;
        RECT 556.950 520.500 559.050 522.600 ;
        RECT 547.950 514.500 550.050 516.600 ;
        RECT 547.950 499.950 550.050 502.050 ;
        RECT 548.400 493.050 549.600 499.950 ;
        RECT 557.400 496.050 558.600 520.500 ;
        RECT 556.950 493.950 559.050 496.050 ;
        RECT 547.950 490.950 550.050 493.050 ;
        RECT 544.950 472.950 547.050 475.050 ;
        RECT 538.950 460.950 541.050 463.050 ;
        RECT 529.950 457.950 532.050 460.050 ;
        RECT 541.950 457.950 544.050 460.050 ;
        RECT 542.400 450.600 543.600 457.950 ;
        RECT 545.400 454.050 546.600 472.950 ;
        RECT 556.950 469.950 559.050 472.050 ;
        RECT 550.950 463.950 553.050 466.050 ;
        RECT 544.950 451.950 547.050 454.050 ;
        RECT 539.400 449.400 543.600 450.600 ;
        RECT 539.400 448.050 540.600 449.400 ;
        RECT 535.950 445.950 538.050 448.050 ;
        RECT 538.950 445.950 541.050 448.050 ;
        RECT 526.950 416.100 529.050 418.200 ;
        RECT 536.400 418.050 537.600 445.950 ;
        RECT 545.400 442.050 546.600 451.950 ;
        RECT 544.950 439.950 547.050 442.050 ;
        RECT 538.950 433.950 541.050 436.050 ;
        RECT 539.400 418.200 540.600 433.950 ;
        RECT 544.950 424.950 547.050 427.050 ;
        RECT 527.400 415.050 528.600 416.100 ;
        RECT 532.950 415.950 535.050 418.050 ;
        RECT 535.950 415.950 538.050 418.050 ;
        RECT 538.950 416.100 541.050 418.200 ;
        RECT 517.950 412.950 520.050 415.050 ;
        RECT 520.950 412.950 523.050 415.050 ;
        RECT 523.950 412.950 526.050 415.050 ;
        RECT 526.950 412.950 529.050 415.050 ;
        RECT 518.400 412.050 519.600 412.950 ;
        RECT 514.950 410.400 519.600 412.050 ;
        RECT 524.400 411.900 525.600 412.950 ;
        RECT 514.950 409.950 519.000 410.400 ;
        RECT 523.950 409.800 526.050 411.900 ;
        RECT 533.400 408.600 534.600 415.950 ;
        RECT 539.400 415.050 540.600 416.100 ;
        RECT 545.400 415.050 546.600 424.950 ;
        RECT 551.400 421.050 552.600 463.950 ;
        RECT 557.400 460.050 558.600 469.950 ;
        RECT 560.400 466.050 561.600 526.950 ;
        RECT 569.400 526.050 570.600 527.100 ;
        RECT 575.400 526.950 580.050 528.600 ;
        RECT 575.400 526.050 576.600 526.950 ;
        RECT 565.950 523.950 568.050 526.050 ;
        RECT 568.950 523.950 571.050 526.050 ;
        RECT 571.950 523.950 574.050 526.050 ;
        RECT 574.950 523.950 577.050 526.050 ;
        RECT 562.950 511.950 565.050 514.050 ;
        RECT 563.400 487.050 564.600 511.950 ;
        RECT 566.400 508.050 567.600 523.950 ;
        RECT 572.400 522.900 573.600 523.950 ;
        RECT 571.950 520.800 574.050 522.900 ;
        RECT 581.400 514.050 582.600 530.400 ;
        RECT 580.950 511.950 583.050 514.050 ;
        RECT 565.950 505.950 568.050 508.050 ;
        RECT 574.950 494.100 577.050 496.200 ;
        RECT 575.400 493.050 576.600 494.100 ;
        RECT 580.950 493.950 583.050 499.050 ;
        RECT 584.400 498.600 585.600 565.800 ;
        RECT 602.400 535.050 603.600 572.400 ;
        RECT 610.950 572.100 613.050 574.200 ;
        RECT 611.400 571.050 612.600 572.100 ;
        RECT 607.950 568.950 610.050 571.050 ;
        RECT 610.950 568.950 613.050 571.050 ;
        RECT 608.400 564.600 609.600 568.950 ;
        RECT 608.400 563.400 612.600 564.600 ;
        RECT 607.950 556.950 610.050 559.050 ;
        RECT 601.950 532.950 604.050 535.050 ;
        RECT 589.950 528.600 594.000 529.050 ;
        RECT 589.950 526.950 594.600 528.600 ;
        RECT 601.950 528.000 604.050 531.900 ;
        RECT 593.400 526.050 594.600 526.950 ;
        RECT 602.400 526.050 603.600 528.000 ;
        RECT 592.950 523.950 595.050 526.050 ;
        RECT 601.950 523.950 604.050 526.050 ;
        RECT 589.950 520.950 592.050 523.050 ;
        RECT 590.400 508.050 591.600 520.950 ;
        RECT 589.950 505.950 592.050 508.050 ;
        RECT 591.000 504.900 594.000 505.050 ;
        RECT 589.950 504.450 594.000 504.900 ;
        RECT 589.950 504.000 594.600 504.450 ;
        RECT 589.950 502.950 595.050 504.000 ;
        RECT 595.950 502.950 598.050 505.050 ;
        RECT 604.950 502.950 607.050 505.050 ;
        RECT 589.950 502.800 592.050 502.950 ;
        RECT 592.950 499.950 595.050 502.950 ;
        RECT 584.400 497.400 588.600 498.600 ;
        RECT 574.950 490.950 577.050 493.050 ;
        RECT 577.950 490.950 580.050 493.050 ;
        RECT 583.950 490.950 586.050 493.050 ;
        RECT 578.400 489.000 579.600 490.950 ;
        RECT 562.950 484.950 565.050 487.050 ;
        RECT 577.950 484.950 580.050 489.000 ;
        RECT 584.400 484.050 585.600 490.950 ;
        RECT 587.400 487.050 588.600 497.400 ;
        RECT 596.400 493.050 597.600 502.950 ;
        RECT 601.950 494.100 604.050 496.200 ;
        RECT 605.400 496.050 606.600 502.950 ;
        RECT 602.400 493.050 603.600 494.100 ;
        RECT 604.950 493.950 607.050 496.050 ;
        RECT 592.950 490.950 595.050 493.050 ;
        RECT 595.950 490.950 598.050 493.050 ;
        RECT 598.950 490.950 601.050 493.050 ;
        RECT 601.950 490.950 604.050 493.050 ;
        RECT 593.400 490.050 594.600 490.950 ;
        RECT 589.950 488.400 594.600 490.050 ;
        RECT 589.950 487.950 594.000 488.400 ;
        RECT 586.950 484.950 589.050 487.050 ;
        RECT 592.950 486.600 597.000 487.050 ;
        RECT 592.950 484.950 597.600 486.600 ;
        RECT 583.950 481.950 586.050 484.050 ;
        RECT 586.950 481.800 589.050 483.900 ;
        RECT 589.950 481.950 592.050 484.050 ;
        RECT 559.950 463.950 562.050 466.050 ;
        RECT 568.950 460.950 571.050 463.050 ;
        RECT 556.950 457.950 559.050 460.050 ;
        RECT 559.950 449.100 562.050 451.200 ;
        RECT 560.400 448.050 561.600 449.100 ;
        RECT 556.950 445.950 559.050 448.050 ;
        RECT 559.950 445.950 562.050 448.050 ;
        RECT 557.400 444.000 558.600 445.950 ;
        RECT 556.950 439.950 559.050 444.000 ;
        RECT 569.400 442.050 570.600 460.950 ;
        RECT 587.400 454.050 588.600 481.800 ;
        RECT 590.400 469.050 591.600 481.950 ;
        RECT 589.950 466.950 592.050 469.050 ;
        RECT 586.950 451.950 589.050 454.050 ;
        RECT 590.400 451.200 591.600 466.950 ;
        RECT 596.400 454.200 597.600 484.950 ;
        RECT 599.400 484.050 600.600 490.950 ;
        RECT 604.950 487.950 607.050 490.050 ;
        RECT 598.950 481.950 601.050 484.050 ;
        RECT 595.950 452.100 598.050 454.200 ;
        RECT 589.950 449.100 592.050 451.200 ;
        RECT 590.400 448.050 591.600 449.100 ;
        RECT 601.950 448.950 604.050 451.050 ;
        RECT 574.950 445.950 577.050 448.050 ;
        RECT 589.950 445.950 592.050 448.050 ;
        RECT 592.950 445.950 595.050 448.050 ;
        RECT 562.950 439.950 565.050 442.050 ;
        RECT 568.950 439.950 571.050 442.050 ;
        RECT 550.950 418.950 553.050 421.050 ;
        RECT 556.950 418.950 559.050 421.050 ;
        RECT 553.950 415.950 556.050 418.050 ;
        RECT 538.950 412.950 541.050 415.050 ;
        RECT 541.950 412.950 544.050 415.050 ;
        RECT 544.950 412.950 547.050 415.050 ;
        RECT 547.950 412.950 550.050 415.050 ;
        RECT 535.950 409.950 538.050 412.050 ;
        RECT 542.400 411.900 543.600 412.950 ;
        RECT 530.400 407.400 534.600 408.600 ;
        RECT 511.950 388.950 514.050 391.050 ;
        RECT 511.950 379.950 514.050 382.050 ;
        RECT 508.950 346.950 511.050 349.050 ;
        RECT 506.400 338.400 510.600 339.600 ;
        RECT 503.400 337.050 504.600 338.100 ;
        RECT 475.950 334.950 478.050 337.050 ;
        RECT 478.950 334.950 481.050 337.050 ;
        RECT 481.950 334.950 484.050 337.050 ;
        RECT 493.950 334.950 496.050 337.050 ;
        RECT 496.950 334.950 499.050 337.050 ;
        RECT 499.950 334.950 502.050 337.050 ;
        RECT 502.950 334.950 505.050 337.050 ;
        RECT 479.400 333.000 480.600 334.950 ;
        RECT 494.400 333.000 495.600 334.950 ;
        RECT 500.400 333.900 501.600 334.950 ;
        RECT 509.400 333.900 510.600 338.400 ;
        RECT 478.950 328.950 481.050 333.000 ;
        RECT 493.950 328.950 496.050 333.000 ;
        RECT 499.950 331.800 502.050 333.900 ;
        RECT 508.950 331.800 511.050 333.900 ;
        RECT 478.950 322.950 481.050 325.050 ;
        RECT 469.950 301.950 472.050 304.050 ;
        RECT 463.950 298.950 466.050 301.050 ;
        RECT 472.950 298.950 475.050 301.050 ;
        RECT 451.950 295.950 454.050 298.050 ;
        RECT 465.000 297.600 469.050 298.050 ;
        RECT 464.400 295.950 469.050 297.600 ;
        RECT 448.950 262.950 451.050 265.050 ;
        RECT 445.950 259.950 448.050 262.050 ;
        RECT 449.400 259.050 450.600 262.950 ;
        RECT 452.400 262.050 453.600 295.950 ;
        RECT 454.950 292.950 457.050 295.050 ;
        RECT 455.400 268.050 456.600 292.950 ;
        RECT 464.400 292.050 465.600 295.950 ;
        RECT 460.950 289.950 463.050 292.050 ;
        RECT 463.950 289.950 466.050 292.050 ;
        RECT 466.950 289.950 469.050 292.050 ;
        RECT 461.400 288.000 462.600 289.950 ;
        RECT 467.400 288.000 468.600 289.950 ;
        RECT 460.950 280.950 463.050 288.000 ;
        RECT 466.950 283.950 469.050 288.000 ;
        RECT 473.400 283.050 474.600 298.950 ;
        RECT 479.400 295.200 480.600 322.950 ;
        RECT 499.950 302.400 502.050 304.500 ;
        RECT 478.950 293.100 481.050 295.200 ;
        RECT 484.950 294.000 487.050 298.050 ;
        RECT 496.950 294.000 499.050 298.050 ;
        RECT 479.400 292.050 480.600 293.100 ;
        RECT 485.400 292.050 486.600 294.000 ;
        RECT 497.400 292.050 498.600 294.000 ;
        RECT 478.950 289.950 481.050 292.050 ;
        RECT 481.950 289.950 484.050 292.050 ;
        RECT 484.950 289.950 487.050 292.050 ;
        RECT 487.950 289.950 490.050 292.050 ;
        RECT 496.950 289.950 499.050 292.050 ;
        RECT 475.950 286.950 478.050 289.050 ;
        RECT 472.950 280.950 475.050 283.050 ;
        RECT 454.950 265.950 457.050 268.050 ;
        RECT 466.950 266.400 469.050 268.500 ;
        RECT 451.950 259.950 454.050 262.050 ;
        RECT 448.950 256.950 451.050 259.050 ;
        RECT 454.950 256.950 457.050 259.050 ;
        RECT 463.950 256.950 466.050 259.050 ;
        RECT 442.800 253.800 444.900 255.900 ;
        RECT 445.950 250.950 448.050 256.050 ;
        RECT 451.950 253.950 454.050 256.050 ;
        RECT 439.950 247.950 442.050 250.050 ;
        RECT 448.950 247.950 451.050 250.050 ;
        RECT 433.950 241.950 436.050 244.050 ;
        RECT 434.400 235.050 435.600 241.950 ;
        RECT 445.950 238.950 448.050 241.050 ;
        RECT 433.950 232.950 436.050 235.050 ;
        RECT 436.950 224.400 439.050 226.500 ;
        RECT 418.950 218.100 421.050 220.200 ;
        RECT 418.950 216.600 421.050 217.050 ;
        RECT 416.400 215.400 421.050 216.600 ;
        RECT 418.950 214.950 421.050 215.400 ;
        RECT 424.950 215.100 427.050 217.200 ;
        RECT 433.950 216.000 436.050 220.050 ;
        RECT 419.400 214.050 420.600 214.950 ;
        RECT 425.400 214.050 426.600 215.100 ;
        RECT 434.400 214.050 435.600 216.000 ;
        RECT 418.950 211.950 421.050 214.050 ;
        RECT 421.950 211.950 424.050 214.050 ;
        RECT 424.950 211.950 427.050 214.050 ;
        RECT 433.950 211.950 436.050 214.050 ;
        RECT 422.400 202.050 423.600 211.950 ;
        RECT 437.700 204.600 438.900 224.400 ;
        RECT 442.950 223.950 445.050 226.050 ;
        RECT 443.400 214.050 444.600 223.950 ;
        RECT 446.400 216.600 447.600 238.950 ;
        RECT 449.400 220.050 450.600 247.950 ;
        RECT 448.950 217.950 451.050 220.050 ;
        RECT 446.400 215.400 450.600 216.600 ;
        RECT 442.950 211.950 445.050 214.050 ;
        RECT 449.400 210.600 450.600 215.400 ;
        RECT 446.400 209.400 450.600 210.600 ;
        RECT 436.950 202.500 439.050 204.600 ;
        RECT 415.950 199.950 418.050 202.050 ;
        RECT 421.950 199.950 424.050 202.050 ;
        RECT 412.950 184.950 415.050 187.050 ;
        RECT 416.400 181.050 417.600 199.950 ;
        RECT 421.950 190.950 424.050 193.050 ;
        RECT 406.950 178.950 409.050 181.050 ;
        RECT 409.950 178.950 412.050 181.050 ;
        RECT 412.950 178.950 415.050 181.050 ;
        RECT 415.950 178.950 418.050 181.050 ;
        RECT 407.400 160.050 408.600 178.950 ;
        RECT 413.400 177.900 414.600 178.950 ;
        RECT 412.950 175.800 415.050 177.900 ;
        RECT 418.950 160.950 421.050 163.050 ;
        RECT 406.950 157.950 409.050 160.050 ;
        RECT 406.950 136.950 409.050 139.050 ;
        RECT 412.950 137.100 415.050 139.200 ;
        RECT 400.950 124.950 403.050 127.050 ;
        RECT 407.400 118.050 408.600 136.950 ;
        RECT 413.400 136.050 414.600 137.100 ;
        RECT 412.950 133.950 415.050 136.050 ;
        RECT 406.950 115.950 409.050 118.050 ;
        RECT 415.950 115.950 418.050 118.050 ;
        RECT 385.950 110.400 388.050 112.500 ;
        RECT 376.950 104.400 381.600 105.600 ;
        RECT 382.950 104.400 385.050 106.500 ;
        RECT 376.950 104.100 379.050 104.400 ;
        RECT 361.950 91.950 364.050 94.050 ;
        RECT 358.950 82.950 361.050 85.050 ;
        RECT 365.400 73.050 366.600 104.100 ;
        RECT 371.400 103.050 372.600 104.100 ;
        RECT 377.400 103.050 378.600 104.100 ;
        RECT 383.400 103.050 384.600 104.400 ;
        RECT 370.950 100.950 373.050 103.050 ;
        RECT 373.950 100.950 376.050 103.050 ;
        RECT 376.950 100.950 379.050 103.050 ;
        RECT 382.950 100.950 385.050 103.050 ;
        RECT 374.400 99.900 375.600 100.950 ;
        RECT 373.950 97.800 376.050 99.900 ;
        RECT 386.850 95.400 388.050 110.400 ;
        RECT 391.950 109.950 394.050 112.050 ;
        RECT 406.950 110.400 409.050 112.500 ;
        RECT 392.400 97.050 393.600 109.950 ;
        RECT 394.950 103.950 397.050 106.050 ;
        RECT 395.400 100.050 396.600 103.950 ;
        RECT 400.950 100.950 403.050 103.050 ;
        RECT 394.950 97.950 397.050 100.050 ;
        RECT 401.400 99.000 402.600 100.950 ;
        RECT 385.950 93.300 388.050 95.400 ;
        RECT 391.950 94.950 394.050 97.050 ;
        RECT 400.950 94.950 403.050 99.000 ;
        RECT 386.850 89.700 388.050 93.300 ;
        RECT 407.100 90.600 408.300 110.400 ;
        RECT 409.950 100.950 412.050 103.050 ;
        RECT 410.400 99.600 411.600 100.950 ;
        RECT 416.400 99.600 417.600 115.950 ;
        RECT 409.950 97.500 412.050 99.600 ;
        RECT 415.950 97.500 418.050 99.600 ;
        RECT 385.950 87.600 388.050 89.700 ;
        RECT 406.950 88.500 409.050 90.600 ;
        RECT 403.950 82.950 406.050 85.050 ;
        RECT 364.950 70.950 367.050 73.050 ;
        RECT 361.950 64.950 364.050 67.050 ;
        RECT 358.950 58.950 361.050 61.050 ;
        RECT 325.950 55.950 328.050 58.050 ;
        RECT 328.950 55.950 331.050 58.050 ;
        RECT 331.950 55.950 334.050 58.050 ;
        RECT 334.950 55.950 337.050 58.050 ;
        RECT 340.950 55.950 343.050 58.050 ;
        RECT 346.950 55.950 349.050 58.050 ;
        RECT 349.950 55.950 352.050 58.050 ;
        RECT 352.950 55.950 355.050 58.050 ;
        RECT 326.400 54.900 327.600 55.950 ;
        RECT 325.950 52.800 328.050 54.900 ;
        RECT 316.950 49.950 319.050 52.050 ;
        RECT 304.950 31.950 307.050 34.050 ;
        RECT 313.950 32.400 316.050 34.500 ;
        RECT 298.950 28.950 301.050 31.050 ;
        RECT 298.950 22.950 301.050 25.050 ;
        RECT 299.400 21.600 300.600 22.950 ;
        RECT 305.400 22.050 306.600 31.950 ;
        RECT 298.950 19.500 301.050 21.600 ;
        RECT 304.950 19.950 307.050 22.050 ;
        RECT 313.950 17.400 315.150 32.400 ;
        RECT 316.950 26.400 319.050 28.500 ;
        RECT 332.400 28.200 333.600 55.950 ;
        RECT 341.400 52.050 342.600 55.950 ;
        RECT 347.400 54.900 348.600 55.950 ;
        RECT 353.400 54.900 354.600 55.950 ;
        RECT 346.950 52.800 349.050 54.900 ;
        RECT 340.950 49.950 343.050 52.050 ;
        RECT 340.950 37.950 343.050 40.050 ;
        RECT 341.400 34.050 342.600 37.950 ;
        RECT 340.950 31.950 343.050 34.050 ;
        RECT 317.400 25.050 318.600 26.400 ;
        RECT 331.950 26.100 334.050 28.200 ;
        RECT 332.400 25.050 333.600 26.100 ;
        RECT 316.950 22.950 319.050 25.050 ;
        RECT 331.950 22.950 334.050 25.050 ;
        RECT 334.950 22.950 337.050 25.050 ;
        RECT 335.400 21.600 336.600 22.950 ;
        RECT 341.400 21.600 342.600 31.950 ;
        RECT 347.400 28.200 348.600 52.800 ;
        RECT 352.950 49.950 355.050 54.900 ;
        RECT 359.400 34.050 360.600 58.950 ;
        RECT 362.400 55.050 363.600 64.950 ;
        RECT 388.950 61.950 391.050 64.050 ;
        RECT 370.950 59.100 373.050 61.200 ;
        RECT 376.950 59.100 379.050 61.200 ;
        RECT 371.400 58.050 372.600 59.100 ;
        RECT 377.400 58.050 378.600 59.100 ;
        RECT 385.950 58.950 388.050 61.050 ;
        RECT 370.950 55.950 373.050 58.050 ;
        RECT 373.950 55.950 376.050 58.050 ;
        RECT 376.950 55.950 379.050 58.050 ;
        RECT 379.950 55.950 382.050 58.050 ;
        RECT 361.950 52.950 364.050 55.050 ;
        RECT 374.400 54.900 375.600 55.950 ;
        RECT 373.950 52.800 376.050 54.900 ;
        RECT 380.400 37.050 381.600 55.950 ;
        RECT 386.400 52.050 387.600 58.950 ;
        RECT 385.950 49.950 388.050 52.050 ;
        RECT 389.400 40.050 390.600 61.950 ;
        RECT 391.950 60.600 396.000 61.050 ;
        RECT 391.950 58.950 396.600 60.600 ;
        RECT 395.400 58.050 396.600 58.950 ;
        RECT 394.950 55.950 397.050 58.050 ;
        RECT 397.950 55.950 400.050 58.050 ;
        RECT 398.400 54.900 399.600 55.950 ;
        RECT 397.950 52.800 400.050 54.900 ;
        RECT 398.400 43.050 399.600 52.800 ;
        RECT 404.400 52.050 405.600 82.950 ;
        RECT 416.400 64.050 417.600 97.500 ;
        RECT 419.400 97.050 420.600 160.950 ;
        RECT 422.400 109.050 423.600 190.950 ;
        RECT 442.950 187.950 445.050 190.050 ;
        RECT 424.950 184.950 427.050 187.050 ;
        RECT 425.400 177.900 426.600 184.950 ;
        RECT 430.950 183.000 433.050 187.050 ;
        RECT 431.400 181.050 432.600 183.000 ;
        RECT 436.950 182.100 439.050 184.200 ;
        RECT 437.400 181.050 438.600 182.100 ;
        RECT 430.950 178.950 433.050 181.050 ;
        RECT 433.950 178.950 436.050 181.050 ;
        RECT 436.950 178.950 439.050 181.050 ;
        RECT 424.950 175.800 427.050 177.900 ;
        RECT 434.400 172.050 435.600 178.950 ;
        RECT 433.950 169.950 436.050 172.050 ;
        RECT 430.950 163.950 433.050 166.050 ;
        RECT 431.400 136.050 432.600 163.950 ;
        RECT 443.400 160.050 444.600 187.950 ;
        RECT 442.950 157.950 445.050 160.050 ;
        RECT 436.950 145.950 439.050 148.050 ;
        RECT 437.400 136.050 438.600 145.950 ;
        RECT 442.950 139.950 445.050 142.050 ;
        RECT 430.950 133.950 433.050 136.050 ;
        RECT 433.950 133.950 436.050 136.050 ;
        RECT 436.950 133.950 439.050 136.050 ;
        RECT 434.400 132.900 435.600 133.950 ;
        RECT 433.950 130.800 436.050 132.900 ;
        RECT 443.400 124.050 444.600 139.950 ;
        RECT 442.950 121.950 445.050 124.050 ;
        RECT 427.950 109.950 430.050 112.050 ;
        RECT 421.950 106.950 424.050 109.050 ;
        RECT 421.950 103.800 424.050 105.900 ;
        RECT 422.400 99.900 423.600 103.800 ;
        RECT 428.400 103.050 429.600 109.950 ;
        RECT 433.950 105.000 436.050 109.050 ;
        RECT 434.400 103.050 435.600 105.000 ;
        RECT 442.950 104.100 445.050 106.200 ;
        RECT 427.950 100.950 430.050 103.050 ;
        RECT 430.950 100.950 433.050 103.050 ;
        RECT 433.950 100.950 436.050 103.050 ;
        RECT 436.950 100.950 439.050 103.050 ;
        RECT 431.400 99.900 432.600 100.950 ;
        RECT 421.950 97.800 424.050 99.900 ;
        RECT 430.950 97.800 433.050 99.900 ;
        RECT 437.400 97.050 438.600 100.950 ;
        RECT 418.950 94.950 421.050 97.050 ;
        RECT 436.950 94.950 439.050 97.050 ;
        RECT 427.950 67.950 430.050 70.050 ;
        RECT 415.950 61.950 418.050 64.050 ;
        RECT 412.950 59.100 415.050 61.200 ;
        RECT 418.950 59.100 421.050 61.200 ;
        RECT 424.950 59.100 427.050 61.200 ;
        RECT 413.400 58.050 414.600 59.100 ;
        RECT 419.400 58.050 420.600 59.100 ;
        RECT 409.950 55.950 412.050 58.050 ;
        RECT 412.950 55.950 415.050 58.050 ;
        RECT 415.950 55.950 418.050 58.050 ;
        RECT 418.950 55.950 421.050 58.050 ;
        RECT 403.950 49.950 406.050 52.050 ;
        RECT 403.950 46.800 406.050 48.900 ;
        RECT 397.950 40.950 400.050 43.050 ;
        RECT 388.950 37.950 391.050 40.050 ;
        RECT 394.950 37.950 397.050 40.050 ;
        RECT 370.950 34.950 373.050 37.050 ;
        RECT 379.950 34.950 382.050 37.050 ;
        RECT 358.950 31.950 361.050 34.050 ;
        RECT 364.950 32.400 367.050 34.500 ;
        RECT 346.950 26.100 349.050 28.200 ;
        RECT 355.950 26.100 358.050 28.200 ;
        RECT 361.950 26.400 364.050 28.500 ;
        RECT 356.400 25.050 357.600 26.100 ;
        RECT 362.400 25.050 363.600 26.400 ;
        RECT 352.950 22.950 355.050 25.050 ;
        RECT 355.950 22.950 358.050 25.050 ;
        RECT 361.950 22.950 364.050 25.050 ;
        RECT 353.400 21.900 354.600 22.950 ;
        RECT 335.400 20.400 342.600 21.600 ;
        RECT 352.950 19.800 355.050 21.900 ;
        RECT 365.850 17.400 367.050 32.400 ;
        RECT 371.400 21.900 372.600 34.950 ;
        RECT 385.950 32.400 388.050 34.500 ;
        RECT 379.950 22.950 382.050 25.050 ;
        RECT 370.950 19.800 373.050 21.900 ;
        RECT 380.400 21.600 381.600 22.950 ;
        RECT 379.950 19.500 382.050 21.600 ;
        RECT 313.950 15.300 316.050 17.400 ;
        RECT 364.950 15.300 367.050 17.400 ;
        RECT 292.950 10.500 295.050 12.600 ;
        RECT 313.950 11.700 315.150 15.300 ;
        RECT 365.850 11.700 367.050 15.300 ;
        RECT 386.100 12.600 387.300 32.400 ;
        RECT 388.950 22.950 391.050 25.050 ;
        RECT 389.400 21.600 390.600 22.950 ;
        RECT 395.400 21.600 396.600 37.950 ;
        RECT 397.950 34.950 400.050 37.050 ;
        RECT 398.400 21.900 399.600 34.950 ;
        RECT 404.400 25.050 405.600 46.800 ;
        RECT 410.400 37.050 411.600 55.950 ;
        RECT 416.400 54.000 417.600 55.950 ;
        RECT 415.950 49.950 418.050 54.000 ;
        RECT 425.400 49.050 426.600 59.100 ;
        RECT 424.950 46.950 427.050 49.050 ;
        RECT 409.950 34.950 412.050 37.050 ;
        RECT 418.950 31.950 421.050 34.050 ;
        RECT 409.950 26.100 412.050 28.200 ;
        RECT 410.400 25.050 411.600 26.100 ;
        RECT 403.950 22.950 406.050 25.050 ;
        RECT 406.950 22.950 409.050 25.050 ;
        RECT 409.950 22.950 412.050 25.050 ;
        RECT 412.950 22.950 415.050 25.050 ;
        RECT 407.400 21.900 408.600 22.950 ;
        RECT 413.400 21.900 414.600 22.950 ;
        RECT 419.400 21.900 420.600 31.950 ;
        RECT 425.400 28.050 426.600 46.950 ;
        RECT 428.400 40.050 429.600 67.950 ;
        RECT 437.400 61.200 438.600 94.950 ;
        RECT 443.400 88.050 444.600 104.100 ;
        RECT 442.950 85.950 445.050 88.050 ;
        RECT 443.400 70.050 444.600 85.950 ;
        RECT 446.400 85.050 447.600 209.400 ;
        RECT 452.400 193.050 453.600 253.950 ;
        RECT 455.400 232.050 456.600 256.950 ;
        RECT 464.400 255.600 465.600 256.950 ;
        RECT 463.950 253.500 466.050 255.600 ;
        RECT 464.400 250.050 465.600 253.500 ;
        RECT 463.950 247.950 466.050 250.050 ;
        RECT 467.700 246.600 468.900 266.400 ;
        RECT 476.400 262.050 477.600 286.950 ;
        RECT 482.400 283.050 483.600 289.950 ;
        RECT 488.400 288.900 489.600 289.950 ;
        RECT 487.950 286.800 490.050 288.900 ;
        RECT 481.950 280.950 484.050 283.050 ;
        RECT 500.700 282.600 501.900 302.400 ;
        RECT 505.950 293.400 508.050 295.500 ;
        RECT 506.400 292.050 507.600 293.400 ;
        RECT 505.950 289.950 508.050 292.050 ;
        RECT 512.400 283.050 513.600 379.950 ;
        RECT 530.400 376.050 531.600 407.400 ;
        RECT 536.400 406.050 537.600 409.950 ;
        RECT 541.950 409.800 544.050 411.900 ;
        RECT 548.400 406.050 549.600 412.950 ;
        RECT 535.950 405.600 538.050 406.050 ;
        RECT 533.400 404.400 538.050 405.600 ;
        RECT 517.950 373.950 520.050 376.050 ;
        RECT 529.950 373.950 532.050 376.050 ;
        RECT 514.950 370.950 517.050 373.050 ;
        RECT 515.400 358.050 516.600 370.950 ;
        RECT 514.950 355.950 517.050 358.050 ;
        RECT 518.400 349.050 519.600 373.950 ;
        RECT 523.950 371.100 526.050 373.200 ;
        RECT 524.400 370.050 525.600 371.100 ;
        RECT 533.400 370.050 534.600 404.400 ;
        RECT 535.950 403.950 538.050 404.400 ;
        RECT 547.950 403.950 550.050 406.050 ;
        RECT 550.950 388.950 553.050 391.050 ;
        RECT 538.950 382.950 541.050 385.050 ;
        RECT 523.950 367.950 526.050 370.050 ;
        RECT 529.950 367.950 532.050 370.050 ;
        RECT 532.950 367.950 535.050 370.050 ;
        RECT 530.400 366.900 531.600 367.950 ;
        RECT 529.950 364.800 532.050 366.900 ;
        RECT 532.950 361.950 535.050 364.050 ;
        RECT 517.950 346.950 520.050 349.050 ;
        RECT 518.400 346.050 519.600 346.950 ;
        RECT 514.950 344.400 519.600 346.050 ;
        RECT 514.950 343.950 519.000 344.400 ;
        RECT 515.400 342.000 525.600 342.600 ;
        RECT 514.950 341.400 525.600 342.000 ;
        RECT 514.950 337.950 517.050 341.400 ;
        RECT 517.950 338.100 520.050 340.200 ;
        RECT 518.400 337.050 519.600 338.100 ;
        RECT 524.400 337.050 525.600 341.400 ;
        RECT 533.400 340.050 534.600 361.950 ;
        RECT 539.400 355.050 540.600 382.950 ;
        RECT 541.950 373.950 544.050 376.050 ;
        RECT 542.400 364.050 543.600 373.950 ;
        RECT 551.400 370.050 552.600 388.950 ;
        RECT 554.400 376.050 555.600 415.950 ;
        RECT 557.400 411.900 558.600 418.950 ;
        RECT 563.400 415.050 564.600 439.950 ;
        RECT 575.400 430.050 576.600 445.950 ;
        RECT 574.950 427.950 577.050 430.050 ;
        RECT 571.950 424.950 574.050 427.050 ;
        RECT 568.950 416.100 571.050 418.200 ;
        RECT 572.400 418.050 573.600 424.950 ;
        RECT 575.400 418.200 576.600 427.950 ;
        RECT 593.400 421.050 594.600 445.950 ;
        RECT 595.950 439.950 598.050 442.050 ;
        RECT 592.950 418.950 595.050 421.050 ;
        RECT 569.400 415.050 570.600 416.100 ;
        RECT 571.950 415.950 574.050 418.050 ;
        RECT 574.950 416.100 577.050 418.200 ;
        RECT 562.950 412.950 565.050 415.050 ;
        RECT 565.950 412.950 568.050 415.050 ;
        RECT 568.950 412.950 571.050 415.050 ;
        RECT 556.950 409.800 559.050 411.900 ;
        RECT 566.400 376.050 567.600 412.950 ;
        RECT 575.400 385.050 576.600 416.100 ;
        RECT 577.950 415.950 580.050 418.050 ;
        RECT 580.950 415.950 583.050 418.050 ;
        RECT 589.950 416.100 592.050 418.200 ;
        RECT 578.400 400.050 579.600 415.950 ;
        RECT 577.950 397.950 580.050 400.050 ;
        RECT 574.950 382.950 577.050 385.050 ;
        RECT 553.950 373.950 556.050 376.050 ;
        RECT 556.950 372.000 559.050 376.050 ;
        RECT 565.950 375.600 568.050 376.050 ;
        RECT 563.400 374.400 568.050 375.600 ;
        RECT 557.400 370.050 558.600 372.000 ;
        RECT 547.950 367.950 550.050 370.050 ;
        RECT 550.950 367.950 553.050 370.050 ;
        RECT 553.950 367.950 556.050 370.050 ;
        RECT 556.950 367.950 559.050 370.050 ;
        RECT 548.400 366.000 549.600 367.950 ;
        RECT 541.950 361.950 544.050 364.050 ;
        RECT 547.950 361.950 550.050 366.000 ;
        RECT 538.950 352.950 541.050 355.050 ;
        RECT 532.950 337.950 535.050 340.050 ;
        RECT 539.400 339.600 540.600 352.950 ;
        RECT 541.950 346.950 544.050 349.050 ;
        RECT 536.400 338.400 540.600 339.600 ;
        RECT 517.950 334.950 520.050 337.050 ;
        RECT 520.950 334.950 523.050 337.050 ;
        RECT 523.950 334.950 526.050 337.050 ;
        RECT 526.950 334.950 529.050 337.050 ;
        RECT 514.950 331.950 517.050 334.050 ;
        RECT 521.400 333.000 522.600 334.950 ;
        RECT 527.400 333.000 528.600 334.950 ;
        RECT 532.950 334.800 535.050 336.900 ;
        RECT 499.950 280.500 502.050 282.600 ;
        RECT 505.950 280.950 508.050 283.050 ;
        RECT 511.950 280.950 514.050 283.050 ;
        RECT 481.950 271.950 484.050 274.050 ;
        RECT 478.950 268.950 481.050 271.050 ;
        RECT 475.950 259.950 478.050 262.050 ;
        RECT 472.950 256.950 475.050 259.050 ;
        RECT 473.400 250.050 474.600 256.950 ;
        RECT 475.950 253.950 478.050 256.050 ;
        RECT 472.950 247.950 475.050 250.050 ;
        RECT 466.950 244.500 469.050 246.600 ;
        RECT 476.400 241.050 477.600 253.950 ;
        RECT 479.400 250.050 480.600 268.950 ;
        RECT 478.950 247.950 481.050 250.050 ;
        RECT 466.950 238.950 469.050 241.050 ;
        RECT 475.950 238.950 478.050 241.050 ;
        RECT 454.950 229.950 457.050 232.050 ;
        RECT 457.950 225.300 460.050 227.400 ;
        RECT 457.950 221.700 459.150 225.300 ;
        RECT 457.950 219.600 460.050 221.700 ;
        RECT 457.950 204.600 459.150 219.600 ;
        RECT 460.950 211.950 463.050 214.050 ;
        RECT 461.400 210.600 462.600 211.950 ;
        RECT 460.950 208.500 463.050 210.600 ;
        RECT 457.950 202.500 460.050 204.600 ;
        RECT 463.950 202.950 466.050 205.050 ;
        RECT 451.950 190.950 454.050 193.050 ;
        RECT 451.950 187.800 454.050 189.900 ;
        RECT 452.400 181.050 453.600 187.800 ;
        RECT 451.950 178.950 454.050 181.050 ;
        RECT 454.950 178.950 457.050 181.050 ;
        RECT 455.400 177.900 456.600 178.950 ;
        RECT 464.400 178.050 465.600 202.950 ;
        RECT 454.950 175.800 457.050 177.900 ;
        RECT 463.950 175.950 466.050 178.050 ;
        RECT 467.400 175.050 468.600 238.950 ;
        RECT 469.950 229.950 472.050 232.050 ;
        RECT 470.400 193.050 471.600 229.950 ;
        RECT 482.400 223.050 483.600 271.950 ;
        RECT 487.950 266.400 490.050 268.500 ;
        RECT 487.950 251.400 489.150 266.400 ;
        RECT 490.950 261.000 493.050 265.050 ;
        RECT 496.950 262.950 499.050 265.050 ;
        RECT 491.400 259.050 492.600 261.000 ;
        RECT 490.950 256.950 493.050 259.050 ;
        RECT 487.950 249.300 490.050 251.400 ;
        RECT 487.950 245.700 489.150 249.300 ;
        RECT 497.400 247.050 498.600 262.950 ;
        RECT 506.400 262.200 507.600 280.950 ;
        RECT 515.400 280.050 516.600 331.950 ;
        RECT 520.950 328.950 523.050 333.000 ;
        RECT 526.950 328.950 529.050 333.000 ;
        RECT 533.400 328.050 534.600 334.800 ;
        RECT 536.400 333.900 537.600 338.400 ;
        RECT 542.400 337.050 543.600 346.950 ;
        RECT 547.950 338.100 550.050 340.200 ;
        RECT 554.400 340.050 555.600 367.950 ;
        RECT 556.950 352.950 559.050 355.050 ;
        RECT 548.400 337.050 549.600 338.100 ;
        RECT 553.950 337.950 556.050 340.050 ;
        RECT 541.950 334.950 544.050 337.050 ;
        RECT 544.950 334.950 547.050 337.050 ;
        RECT 547.950 334.950 550.050 337.050 ;
        RECT 550.950 334.950 553.050 337.050 ;
        RECT 545.400 333.900 546.600 334.950 ;
        RECT 551.400 333.900 552.600 334.950 ;
        RECT 557.400 334.050 558.600 352.950 ;
        RECT 563.400 342.600 564.600 374.400 ;
        RECT 565.950 373.950 568.050 374.400 ;
        RECT 565.950 370.800 568.050 372.900 ;
        RECT 574.950 371.100 577.050 373.200 ;
        RECT 560.400 341.400 564.600 342.600 ;
        RECT 535.950 331.800 538.050 333.900 ;
        RECT 544.950 331.800 547.050 333.900 ;
        RECT 550.950 331.800 553.050 333.900 ;
        RECT 556.950 331.950 559.050 334.050 ;
        RECT 541.950 330.600 544.050 331.050 ;
        RECT 547.950 330.600 550.050 331.050 ;
        RECT 541.950 329.400 550.050 330.600 ;
        RECT 541.950 328.950 544.050 329.400 ;
        RECT 547.950 328.950 550.050 329.400 ;
        RECT 556.950 328.800 559.050 330.900 ;
        RECT 532.950 325.950 535.050 328.050 ;
        RECT 537.000 327.900 541.050 328.050 ;
        RECT 535.950 325.950 541.050 327.900 ;
        RECT 535.950 325.800 538.050 325.950 ;
        RECT 520.950 303.300 523.050 305.400 ;
        RECT 520.950 299.700 522.150 303.300 ;
        RECT 520.950 297.600 523.050 299.700 ;
        RECT 550.950 298.950 553.050 301.050 ;
        RECT 520.950 282.600 522.150 297.600 ;
        RECT 541.950 293.100 544.050 295.200 ;
        RECT 542.400 292.050 543.600 293.100 ;
        RECT 551.400 292.050 552.600 298.950 ;
        RECT 523.950 289.950 526.050 292.050 ;
        RECT 541.950 289.950 544.050 292.050 ;
        RECT 544.950 289.950 547.050 292.050 ;
        RECT 550.950 289.950 553.050 292.050 ;
        RECT 524.400 288.000 525.600 289.950 ;
        RECT 523.950 285.600 526.050 288.000 ;
        RECT 523.950 284.400 528.600 285.600 ;
        RECT 523.950 283.950 526.050 284.400 ;
        RECT 520.950 280.500 523.050 282.600 ;
        RECT 514.950 277.950 517.050 280.050 ;
        RECT 511.950 268.950 514.050 271.050 ;
        RECT 499.950 260.100 502.050 262.200 ;
        RECT 505.950 260.100 508.050 262.200 ;
        RECT 487.950 243.600 490.050 245.700 ;
        RECT 496.950 244.950 499.050 247.050 ;
        RECT 500.400 238.050 501.600 260.100 ;
        RECT 506.400 259.050 507.600 260.100 ;
        RECT 512.400 259.050 513.600 268.950 ;
        RECT 520.950 259.950 523.050 262.050 ;
        RECT 527.400 261.600 528.600 284.400 ;
        RECT 545.400 280.050 546.600 289.950 ;
        RECT 553.950 286.950 556.050 289.050 ;
        RECT 544.950 277.950 547.050 280.050 ;
        RECT 554.400 268.050 555.600 286.950 ;
        RECT 557.400 271.050 558.600 328.800 ;
        RECT 560.400 288.900 561.600 341.400 ;
        RECT 566.400 339.600 567.600 370.800 ;
        RECT 575.400 370.050 576.600 371.100 ;
        RECT 581.400 370.050 582.600 415.950 ;
        RECT 590.400 415.050 591.600 416.100 ;
        RECT 596.400 415.050 597.600 439.950 ;
        RECT 586.950 412.950 589.050 415.050 ;
        RECT 589.950 412.950 592.050 415.050 ;
        RECT 592.950 412.950 595.050 415.050 ;
        RECT 595.950 412.950 598.050 415.050 ;
        RECT 587.400 388.050 588.600 412.950 ;
        RECT 593.400 411.000 594.600 412.950 ;
        RECT 592.950 406.950 595.050 411.000 ;
        RECT 598.950 409.950 601.050 412.050 ;
        RECT 586.950 385.950 589.050 388.050 ;
        RECT 589.950 379.950 592.050 382.050 ;
        RECT 571.950 367.950 574.050 370.050 ;
        RECT 574.950 367.950 577.050 370.050 ;
        RECT 577.950 367.950 580.050 370.050 ;
        RECT 580.950 367.950 583.050 370.050 ;
        RECT 572.400 366.900 573.600 367.950 ;
        RECT 571.950 364.800 574.050 366.900 ;
        RECT 571.950 349.950 574.050 352.050 ;
        RECT 563.400 338.400 567.600 339.600 ;
        RECT 563.400 331.050 564.600 338.400 ;
        RECT 572.400 337.050 573.600 349.950 ;
        RECT 578.400 340.050 579.600 367.950 ;
        RECT 583.950 358.950 586.050 361.050 ;
        RECT 577.950 337.950 580.050 340.050 ;
        RECT 568.950 334.950 571.050 337.050 ;
        RECT 571.950 334.950 574.050 337.050 ;
        RECT 574.950 334.950 577.050 337.050 ;
        RECT 569.400 333.900 570.600 334.950 ;
        RECT 568.950 331.800 571.050 333.900 ;
        RECT 562.950 328.950 565.050 331.050 ;
        RECT 569.400 325.050 570.600 331.800 ;
        RECT 575.400 328.050 576.600 334.950 ;
        RECT 574.950 325.950 577.050 328.050 ;
        RECT 568.950 322.950 571.050 325.050 ;
        RECT 584.400 313.050 585.600 358.950 ;
        RECT 586.950 346.950 589.050 349.050 ;
        RECT 587.400 316.050 588.600 346.950 ;
        RECT 590.400 337.050 591.600 379.950 ;
        RECT 599.400 373.200 600.600 409.950 ;
        RECT 602.400 376.050 603.600 448.950 ;
        RECT 605.400 418.050 606.600 487.950 ;
        RECT 608.400 457.050 609.600 556.950 ;
        RECT 611.400 553.050 612.600 563.400 ;
        RECT 617.400 559.050 618.600 592.950 ;
        RECT 620.400 592.050 621.600 601.950 ;
        RECT 626.400 600.900 627.600 601.950 ;
        RECT 625.950 598.800 628.050 600.900 ;
        RECT 626.400 595.050 627.600 598.800 ;
        RECT 628.950 595.950 631.050 601.050 ;
        RECT 625.950 592.950 628.050 595.050 ;
        RECT 632.400 592.050 633.600 616.950 ;
        RECT 635.400 610.050 636.600 619.950 ;
        RECT 656.400 613.050 657.600 643.950 ;
        RECT 659.400 640.050 660.600 701.400 ;
        RECT 664.950 688.950 667.050 691.050 ;
        RECT 665.400 678.900 666.600 688.950 ;
        RECT 667.950 683.100 670.050 688.050 ;
        RECT 673.950 683.100 676.050 685.200 ;
        RECT 674.400 682.050 675.600 683.100 ;
        RECT 680.400 682.050 681.600 715.950 ;
        RECT 685.950 700.950 688.050 703.050 ;
        RECT 670.950 679.950 673.050 682.050 ;
        RECT 673.950 679.950 676.050 682.050 ;
        RECT 676.950 679.950 679.050 682.050 ;
        RECT 679.950 679.950 682.050 682.050 ;
        RECT 671.400 678.900 672.600 679.950 ;
        RECT 677.400 678.900 678.600 679.950 ;
        RECT 664.950 676.800 667.050 678.900 ;
        RECT 670.950 676.800 673.050 678.900 ;
        RECT 676.950 676.800 679.050 678.900 ;
        RECT 682.950 676.950 685.050 679.050 ;
        RECT 686.400 678.900 687.600 700.950 ;
        RECT 683.400 664.050 684.600 676.950 ;
        RECT 685.950 676.800 688.050 678.900 ;
        RECT 682.800 661.950 684.900 664.050 ;
        RECT 685.950 661.950 688.050 664.050 ;
        RECT 676.950 658.950 679.050 661.050 ;
        RECT 667.950 651.000 670.050 655.050 ;
        RECT 668.400 649.050 669.600 651.000 ;
        RECT 677.400 649.050 678.600 658.950 ;
        RECT 679.950 652.950 682.050 655.050 ;
        RECT 664.950 646.950 667.050 649.050 ;
        RECT 667.950 646.950 670.050 649.050 ;
        RECT 670.950 646.950 673.050 649.050 ;
        RECT 676.950 646.950 679.050 649.050 ;
        RECT 661.950 640.950 664.050 643.050 ;
        RECT 658.950 637.950 661.050 640.050 ;
        RECT 640.950 610.950 643.050 613.050 ;
        RECT 655.950 610.950 658.050 613.050 ;
        RECT 634.950 607.950 637.050 610.050 ;
        RECT 641.400 607.200 642.600 610.950 ;
        RECT 662.400 609.600 663.600 640.950 ;
        RECT 665.400 634.050 666.600 646.950 ;
        RECT 671.400 645.000 672.600 646.950 ;
        RECT 670.950 640.950 673.050 645.000 ;
        RECT 673.950 640.950 676.050 646.050 ;
        RECT 676.950 640.950 679.050 643.050 ;
        RECT 673.950 637.800 676.050 639.900 ;
        RECT 664.950 631.950 667.050 634.050 ;
        RECT 667.950 619.950 670.050 622.050 ;
        RECT 656.400 608.400 663.600 609.600 ;
        RECT 640.950 605.100 643.050 607.200 ;
        RECT 646.950 605.100 649.050 607.200 ;
        RECT 656.400 606.600 657.600 608.400 ;
        RECT 653.400 605.400 657.600 606.600 ;
        RECT 641.400 604.050 642.600 605.100 ;
        RECT 647.400 604.050 648.600 605.100 ;
        RECT 640.950 601.950 643.050 604.050 ;
        RECT 643.950 601.950 646.050 604.050 ;
        RECT 646.950 601.950 649.050 604.050 ;
        RECT 634.950 592.950 637.050 598.050 ;
        RECT 644.400 595.050 645.600 601.950 ;
        RECT 643.950 592.950 646.050 595.050 ;
        RECT 619.950 589.950 622.050 592.050 ;
        RECT 631.950 589.950 634.050 592.050 ;
        RECT 619.950 577.950 622.050 580.050 ;
        RECT 620.400 559.050 621.600 577.950 ;
        RECT 653.400 577.050 654.600 605.400 ;
        RECT 661.950 605.100 664.050 607.200 ;
        RECT 662.400 604.050 663.600 605.100 ;
        RECT 668.400 604.050 669.600 619.950 ;
        RECT 658.950 601.950 661.050 604.050 ;
        RECT 661.950 601.950 664.050 604.050 ;
        RECT 664.950 601.950 667.050 604.050 ;
        RECT 667.950 601.950 670.050 604.050 ;
        RECT 659.400 601.050 660.600 601.950 ;
        RECT 655.950 598.950 660.600 601.050 ;
        RECT 665.400 600.000 666.600 601.950 ;
        RECT 659.400 585.600 660.600 598.950 ;
        RECT 664.950 595.950 667.050 600.000 ;
        RECT 670.950 598.950 673.050 601.050 ;
        RECT 671.400 595.050 672.600 598.950 ;
        RECT 670.950 592.950 673.050 595.050 ;
        RECT 667.950 589.950 670.050 592.050 ;
        RECT 659.400 584.400 663.600 585.600 ;
        RECT 658.950 580.950 661.050 583.050 ;
        RECT 652.950 574.950 655.050 577.050 ;
        RECT 622.950 572.100 625.050 574.200 ;
        RECT 631.950 572.100 634.050 574.200 ;
        RECT 616.800 556.950 618.900 559.050 ;
        RECT 619.950 556.950 622.050 559.050 ;
        RECT 610.950 550.950 613.050 553.050 ;
        RECT 623.400 550.050 624.600 572.100 ;
        RECT 632.400 571.050 633.600 572.100 ;
        RECT 640.950 571.950 643.050 574.050 ;
        RECT 631.950 568.950 634.050 571.050 ;
        RECT 634.950 568.950 637.050 571.050 ;
        RECT 635.400 562.050 636.600 568.950 ;
        RECT 634.950 559.950 637.050 562.050 ;
        RECT 631.950 550.950 634.050 553.050 ;
        RECT 622.950 547.950 625.050 550.050 ;
        RECT 610.950 532.950 613.050 535.050 ;
        RECT 625.950 532.950 628.050 535.050 ;
        RECT 611.400 505.050 612.600 532.950 ;
        RECT 626.400 529.200 627.600 532.950 ;
        RECT 619.950 527.100 622.050 529.200 ;
        RECT 625.950 527.100 628.050 529.200 ;
        RECT 620.400 526.050 621.600 527.100 ;
        RECT 626.400 526.050 627.600 527.100 ;
        RECT 616.950 523.950 619.050 526.050 ;
        RECT 619.950 523.950 622.050 526.050 ;
        RECT 622.950 523.950 625.050 526.050 ;
        RECT 625.950 523.950 628.050 526.050 ;
        RECT 617.400 517.050 618.600 523.950 ;
        RECT 623.400 519.600 624.600 523.950 ;
        RECT 620.400 518.400 624.600 519.600 ;
        RECT 616.950 514.950 619.050 517.050 ;
        RECT 610.950 502.950 613.050 505.050 ;
        RECT 613.950 494.100 616.050 496.200 ;
        RECT 614.400 493.050 615.600 494.100 ;
        RECT 620.400 493.050 621.600 518.400 ;
        RECT 628.950 502.950 631.050 505.050 ;
        RECT 613.950 490.950 616.050 493.050 ;
        RECT 616.950 490.950 619.050 493.050 ;
        RECT 619.950 490.950 622.050 493.050 ;
        RECT 622.950 490.950 625.050 493.050 ;
        RECT 610.950 487.950 613.050 490.050 ;
        RECT 611.400 460.050 612.600 487.950 ;
        RECT 617.400 484.050 618.600 490.950 ;
        RECT 623.400 489.000 624.600 490.950 ;
        RECT 622.950 484.950 625.050 489.000 ;
        RECT 616.950 481.950 619.050 484.050 ;
        RECT 610.950 457.950 613.050 460.050 ;
        RECT 607.950 454.950 610.050 457.050 ;
        RECT 607.950 451.800 610.050 453.900 ;
        RECT 608.400 442.050 609.600 451.800 ;
        RECT 616.950 449.100 619.050 451.200 ;
        RECT 629.400 450.600 630.600 502.950 ;
        RECT 632.400 478.050 633.600 550.950 ;
        RECT 641.400 535.050 642.600 571.950 ;
        RECT 652.950 568.950 655.050 571.050 ;
        RECT 653.400 562.050 654.600 568.950 ;
        RECT 655.950 565.950 658.050 568.050 ;
        RECT 652.950 559.950 655.050 562.050 ;
        RECT 652.950 553.950 655.050 556.050 ;
        RECT 640.950 532.950 643.050 535.050 ;
        RECT 640.950 527.100 643.050 529.200 ;
        RECT 641.400 526.050 642.600 527.100 ;
        RECT 646.950 526.950 649.050 529.050 ;
        RECT 637.950 523.950 640.050 526.050 ;
        RECT 640.950 523.950 643.050 526.050 ;
        RECT 638.400 522.900 639.600 523.950 ;
        RECT 637.950 520.800 640.050 522.900 ;
        RECT 643.950 520.950 646.050 523.050 ;
        RECT 634.950 505.950 637.050 508.050 ;
        RECT 635.400 496.050 636.600 505.950 ;
        RECT 640.950 502.950 643.050 505.050 ;
        RECT 634.950 493.950 637.050 496.050 ;
        RECT 641.400 493.050 642.600 502.950 ;
        RECT 644.400 499.050 645.600 520.950 ;
        RECT 643.950 496.950 646.050 499.050 ;
        RECT 647.400 496.200 648.600 526.950 ;
        RECT 649.950 502.950 652.050 505.050 ;
        RECT 646.950 494.100 649.050 496.200 ;
        RECT 637.950 490.950 640.050 493.050 ;
        RECT 640.950 490.950 643.050 493.050 ;
        RECT 643.950 490.950 646.050 493.050 ;
        RECT 638.400 489.900 639.600 490.950 ;
        RECT 637.950 487.800 640.050 489.900 ;
        RECT 634.950 484.950 637.050 487.050 ;
        RECT 639.000 486.750 642.000 487.050 ;
        RECT 637.950 486.600 642.000 486.750 ;
        RECT 644.400 486.600 645.600 490.950 ;
        RECT 650.400 489.900 651.600 502.950 ;
        RECT 649.950 487.800 652.050 489.900 ;
        RECT 653.400 489.600 654.600 553.950 ;
        RECT 656.400 529.050 657.600 565.950 ;
        RECT 659.400 532.050 660.600 580.950 ;
        RECT 655.950 526.950 658.050 529.050 ;
        RECT 658.950 528.000 661.050 532.050 ;
        RECT 662.400 531.600 663.600 584.400 ;
        RECT 664.950 583.950 667.050 586.050 ;
        RECT 665.400 550.050 666.600 583.950 ;
        RECT 668.400 574.050 669.600 589.950 ;
        RECT 671.400 586.050 672.600 592.950 ;
        RECT 670.950 583.950 673.050 586.050 ;
        RECT 674.400 583.050 675.600 637.800 ;
        RECT 677.400 592.050 678.600 640.950 ;
        RECT 680.400 637.050 681.600 652.950 ;
        RECT 686.400 651.600 687.600 661.950 ;
        RECT 689.400 655.050 690.600 719.400 ;
        RECT 692.400 703.050 693.600 728.100 ;
        RECT 701.400 727.050 702.600 728.100 ;
        RECT 707.400 727.050 708.600 729.000 ;
        RECT 697.950 724.950 700.050 727.050 ;
        RECT 700.950 724.950 703.050 727.050 ;
        RECT 703.950 724.950 706.050 727.050 ;
        RECT 706.950 724.950 709.050 727.050 ;
        RECT 698.400 718.050 699.600 724.950 ;
        RECT 704.400 723.900 705.600 724.950 ;
        RECT 703.950 718.950 706.050 723.900 ;
        RECT 697.950 715.950 700.050 718.050 ;
        RECT 691.950 700.950 694.050 703.050 ;
        RECT 709.950 697.950 712.050 700.050 ;
        RECT 691.950 694.950 694.050 697.050 ;
        RECT 692.400 685.050 693.600 694.950 ;
        RECT 691.950 682.950 694.050 685.050 ;
        RECT 697.950 683.100 700.050 685.200 ;
        RECT 703.950 683.100 706.050 685.200 ;
        RECT 698.400 682.050 699.600 683.100 ;
        RECT 704.400 682.050 705.600 683.100 ;
        RECT 694.950 679.950 697.050 682.050 ;
        RECT 697.950 679.950 700.050 682.050 ;
        RECT 700.950 679.950 703.050 682.050 ;
        RECT 703.950 679.950 706.050 682.050 ;
        RECT 691.950 676.950 694.050 679.050 ;
        RECT 692.400 673.050 693.600 676.950 ;
        RECT 691.950 670.950 694.050 673.050 ;
        RECT 695.400 669.600 696.600 679.950 ;
        RECT 701.400 673.050 702.600 679.950 ;
        RECT 706.950 676.950 709.050 679.050 ;
        RECT 700.950 670.950 703.050 673.050 ;
        RECT 703.950 669.600 706.050 670.050 ;
        RECT 695.400 668.400 706.050 669.600 ;
        RECT 703.950 667.950 706.050 668.400 ;
        RECT 703.950 664.800 706.050 666.900 ;
        RECT 691.950 658.950 694.050 661.050 ;
        RECT 692.400 655.200 693.600 658.950 ;
        RECT 688.950 652.950 691.050 655.050 ;
        RECT 691.950 653.100 694.050 655.200 ;
        RECT 704.400 655.050 705.600 664.800 ;
        RECT 683.400 650.400 687.600 651.600 ;
        RECT 679.950 634.950 682.050 637.050 ;
        RECT 679.950 628.950 682.050 631.050 ;
        RECT 680.400 607.050 681.600 628.950 ;
        RECT 683.400 610.050 684.600 650.400 ;
        RECT 691.950 649.950 694.050 652.050 ;
        RECT 697.950 650.100 700.050 652.200 ;
        RECT 703.950 650.100 706.050 655.050 ;
        RECT 692.400 649.050 693.600 649.950 ;
        RECT 698.400 649.050 699.600 650.100 ;
        RECT 688.950 646.950 691.050 649.050 ;
        RECT 691.950 646.950 694.050 649.050 ;
        RECT 694.950 646.950 697.050 649.050 ;
        RECT 697.950 646.950 700.050 649.050 ;
        RECT 700.950 646.950 703.050 649.050 ;
        RECT 689.400 645.900 690.600 646.950 ;
        RECT 688.950 643.800 691.050 645.900 ;
        RECT 689.400 640.050 690.600 643.800 ;
        RECT 688.950 637.950 691.050 640.050 ;
        RECT 695.400 637.050 696.600 646.950 ;
        RECT 701.400 645.900 702.600 646.950 ;
        RECT 707.400 646.050 708.600 676.950 ;
        RECT 710.400 661.050 711.600 697.950 ;
        RECT 713.400 670.050 714.600 751.950 ;
        RECT 737.400 745.050 738.600 751.950 ;
        RECT 740.400 748.050 741.600 757.950 ;
        RECT 739.950 745.950 742.050 748.050 ;
        RECT 736.950 742.950 739.050 745.050 ;
        RECT 715.950 739.950 718.050 742.050 ;
        RECT 716.400 697.050 717.600 739.950 ;
        RECT 727.950 728.100 730.050 730.200 ;
        RECT 733.950 728.100 736.050 730.200 ;
        RECT 743.400 730.050 744.600 761.100 ;
        RECT 749.400 760.050 750.600 769.950 ;
        RECT 754.950 761.100 757.050 763.200 ;
        RECT 755.400 760.050 756.600 761.100 ;
        RECT 748.950 757.950 751.050 760.050 ;
        RECT 751.950 757.950 754.050 760.050 ;
        RECT 754.950 757.950 757.050 760.050 ;
        RECT 752.400 756.900 753.600 757.950 ;
        RECT 751.950 754.800 754.050 756.900 ;
        RECT 757.950 748.950 760.050 751.050 ;
        RECT 728.400 727.050 729.600 728.100 ;
        RECT 734.400 727.050 735.600 728.100 ;
        RECT 742.950 727.950 745.050 730.050 ;
        RECT 748.950 728.100 751.050 730.200 ;
        RECT 749.400 727.050 750.600 728.100 ;
        RECT 724.950 724.950 727.050 727.050 ;
        RECT 727.950 724.950 730.050 727.050 ;
        RECT 730.950 724.950 733.050 727.050 ;
        RECT 733.950 724.950 736.050 727.050 ;
        RECT 745.950 724.950 748.050 727.050 ;
        RECT 748.950 724.950 751.050 727.050 ;
        RECT 725.400 723.900 726.600 724.950 ;
        RECT 724.950 721.800 727.050 723.900 ;
        RECT 721.950 712.950 724.050 715.050 ;
        RECT 715.800 694.950 717.900 697.050 ;
        RECT 718.950 694.950 721.050 697.050 ;
        RECT 719.400 682.050 720.600 694.950 ;
        RECT 722.400 688.050 723.600 712.950 ;
        RECT 724.950 700.950 727.050 703.050 ;
        RECT 725.400 694.050 726.600 700.950 ;
        RECT 731.400 700.050 732.600 724.950 ;
        RECT 736.950 721.950 739.050 724.050 ;
        RECT 737.400 703.050 738.600 721.950 ;
        RECT 736.950 700.950 739.050 703.050 ;
        RECT 730.950 697.950 733.050 700.050 ;
        RECT 737.400 697.050 738.600 700.950 ;
        RECT 736.950 694.950 739.050 697.050 ;
        RECT 746.400 694.050 747.600 724.950 ;
        RECT 724.950 691.950 727.050 694.050 ;
        RECT 745.950 691.950 748.050 694.050 ;
        RECT 748.950 688.950 751.050 691.050 ;
        RECT 721.950 685.950 724.050 688.050 ;
        RECT 749.400 685.200 750.600 688.950 ;
        RECT 724.950 683.100 727.050 685.200 ;
        RECT 733.950 683.100 736.050 685.200 ;
        RECT 742.950 683.100 745.050 685.200 ;
        RECT 748.950 683.100 751.050 685.200 ;
        RECT 725.400 682.050 726.600 683.100 ;
        RECT 718.950 679.950 721.050 682.050 ;
        RECT 721.950 679.950 724.050 682.050 ;
        RECT 724.950 679.950 727.050 682.050 ;
        RECT 727.950 679.950 730.050 682.050 ;
        RECT 722.400 678.900 723.600 679.950 ;
        RECT 728.400 678.900 729.600 679.950 ;
        RECT 721.950 676.800 724.050 678.900 ;
        RECT 727.950 676.800 730.050 678.900 ;
        RECT 712.950 667.950 715.050 670.050 ;
        RECT 730.950 667.950 733.050 670.050 ;
        RECT 709.950 658.950 712.050 661.050 ;
        RECT 721.950 651.000 724.050 655.050 ;
        RECT 722.400 649.050 723.600 651.000 ;
        RECT 727.950 649.950 730.050 655.050 ;
        RECT 712.950 646.950 715.050 649.050 ;
        RECT 718.950 646.950 721.050 649.050 ;
        RECT 721.950 646.950 724.050 649.050 ;
        RECT 724.950 646.950 727.050 649.050 ;
        RECT 700.950 643.800 703.050 645.900 ;
        RECT 706.950 643.950 709.050 646.050 ;
        RECT 709.950 643.950 712.050 646.050 ;
        RECT 713.400 645.900 714.600 646.950 ;
        RECT 719.400 645.900 720.600 646.950 ;
        RECT 694.950 634.950 697.050 637.050 ;
        RECT 694.950 616.950 697.050 619.050 ;
        RECT 682.950 607.950 685.050 610.050 ;
        RECT 679.950 604.950 682.050 607.050 ;
        RECT 682.950 601.950 685.050 604.050 ;
        RECT 683.400 600.000 684.600 601.950 ;
        RECT 682.950 595.950 685.050 600.000 ;
        RECT 691.950 598.950 694.050 601.050 ;
        RECT 679.950 592.950 682.050 595.050 ;
        RECT 676.950 589.950 679.050 592.050 ;
        RECT 680.400 586.050 681.600 592.950 ;
        RECT 679.950 583.950 682.050 586.050 ;
        RECT 673.950 580.950 676.050 583.050 ;
        RECT 667.950 571.950 670.050 574.050 ;
        RECT 673.950 572.100 676.050 574.200 ;
        RECT 685.950 572.100 688.050 574.200 ;
        RECT 692.400 574.050 693.600 598.950 ;
        RECT 695.400 598.050 696.600 616.950 ;
        RECT 701.400 607.050 702.600 643.800 ;
        RECT 703.950 637.950 706.050 640.050 ;
        RECT 704.400 619.050 705.600 637.950 ;
        RECT 706.950 634.950 709.050 637.050 ;
        RECT 707.400 625.050 708.600 634.950 ;
        RECT 706.950 622.950 709.050 625.050 ;
        RECT 703.950 616.950 706.050 619.050 ;
        RECT 710.400 607.200 711.600 643.950 ;
        RECT 712.950 643.800 715.050 645.900 ;
        RECT 718.950 643.800 721.050 645.900 ;
        RECT 713.400 622.050 714.600 643.800 ;
        RECT 721.950 637.950 724.050 640.050 ;
        RECT 712.950 619.950 715.050 622.050 ;
        RECT 718.950 619.950 721.050 622.050 ;
        RECT 719.400 610.050 720.600 619.950 ;
        RECT 718.950 607.950 721.050 610.050 ;
        RECT 700.950 604.950 703.050 607.050 ;
        RECT 709.950 605.100 712.050 607.200 ;
        RECT 722.400 606.600 723.600 637.950 ;
        RECT 725.400 622.050 726.600 646.950 ;
        RECT 727.950 643.950 730.050 646.050 ;
        RECT 728.400 640.050 729.600 643.950 ;
        RECT 727.950 637.950 730.050 640.050 ;
        RECT 731.400 633.600 732.600 667.950 ;
        RECT 734.400 646.050 735.600 683.100 ;
        RECT 743.400 682.050 744.600 683.100 ;
        RECT 749.400 682.050 750.600 683.100 ;
        RECT 739.950 679.950 742.050 682.050 ;
        RECT 742.950 679.950 745.050 682.050 ;
        RECT 745.950 679.950 748.050 682.050 ;
        RECT 748.950 679.950 751.050 682.050 ;
        RECT 740.400 678.900 741.600 679.950 ;
        RECT 746.400 678.900 747.600 679.950 ;
        RECT 758.400 679.050 759.600 748.950 ;
        RECT 761.400 727.050 762.600 799.800 ;
        RECT 779.400 793.050 780.600 802.950 ;
        RECT 791.400 799.050 792.600 806.100 ;
        RECT 797.400 805.050 798.600 817.950 ;
        RECT 818.400 817.050 819.600 835.950 ;
        RECT 839.400 834.900 840.600 835.950 ;
        RECT 838.950 832.800 841.050 834.900 ;
        RECT 817.950 814.950 820.050 817.050 ;
        RECT 811.950 808.950 814.050 811.050 ;
        RECT 802.950 806.100 805.050 808.200 ;
        RECT 803.400 805.050 804.600 806.100 ;
        RECT 796.950 802.950 799.050 805.050 ;
        RECT 799.950 802.950 802.050 805.050 ;
        RECT 802.950 802.950 805.050 805.050 ;
        RECT 805.950 802.950 808.050 805.050 ;
        RECT 800.400 801.900 801.600 802.950 ;
        RECT 799.950 799.800 802.050 801.900 ;
        RECT 790.950 796.950 793.050 799.050 ;
        RECT 778.950 790.950 781.050 793.050 ;
        RECT 779.400 787.050 780.600 790.950 ;
        RECT 778.950 784.950 781.050 787.050 ;
        RECT 763.950 772.950 766.050 775.050 ;
        RECT 764.400 757.050 765.600 772.950 ;
        RECT 800.400 763.200 801.600 799.800 ;
        RECT 806.400 787.050 807.600 802.950 ;
        RECT 808.950 796.950 811.050 799.050 ;
        RECT 805.950 784.950 808.050 787.050 ;
        RECT 805.950 772.950 808.050 775.050 ;
        RECT 766.950 761.100 769.050 763.200 ;
        RECT 772.950 761.100 775.050 763.200 ;
        RECT 778.950 761.100 781.050 763.200 ;
        RECT 763.950 754.950 766.050 757.050 ;
        RECT 767.400 754.050 768.600 761.100 ;
        RECT 773.400 760.050 774.600 761.100 ;
        RECT 779.400 760.050 780.600 761.100 ;
        RECT 784.950 760.950 787.050 763.050 ;
        RECT 790.950 761.100 793.050 763.200 ;
        RECT 799.950 761.100 802.050 763.200 ;
        RECT 772.950 757.950 775.050 760.050 ;
        RECT 775.950 757.950 778.050 760.050 ;
        RECT 778.950 757.950 781.050 760.050 ;
        RECT 766.950 751.950 769.050 754.050 ;
        RECT 772.950 739.950 775.050 742.050 ;
        RECT 766.950 728.100 769.050 730.200 ;
        RECT 773.400 729.600 774.600 739.950 ;
        RECT 776.400 739.050 777.600 757.950 ;
        RECT 785.400 754.050 786.600 760.950 ;
        RECT 791.400 760.050 792.600 761.100 ;
        RECT 800.400 760.050 801.600 761.100 ;
        RECT 790.950 757.950 793.050 760.050 ;
        RECT 796.950 757.950 799.050 760.050 ;
        RECT 799.950 757.950 802.050 760.050 ;
        RECT 797.400 756.900 798.600 757.950 ;
        RECT 796.950 754.800 799.050 756.900 ;
        RECT 784.950 751.950 787.050 754.050 ;
        RECT 806.400 745.050 807.600 772.950 ;
        RECT 809.400 756.600 810.600 796.950 ;
        RECT 812.400 787.050 813.600 808.950 ;
        RECT 820.950 807.000 823.050 811.050 ;
        RECT 821.400 805.050 822.600 807.000 ;
        RECT 826.950 806.100 829.050 808.200 ;
        RECT 827.400 805.050 828.600 806.100 ;
        RECT 845.400 805.050 846.600 835.950 ;
        RECT 851.400 814.050 852.600 878.400 ;
        RECT 857.400 876.600 858.600 880.950 ;
        RECT 854.400 875.400 858.600 876.600 ;
        RECT 854.400 826.050 855.600 875.400 ;
        RECT 863.400 874.050 864.600 880.950 ;
        RECT 856.950 871.950 859.050 874.050 ;
        RECT 862.950 871.950 865.050 874.050 ;
        RECT 853.950 823.950 856.050 826.050 ;
        RECT 850.950 811.950 853.050 814.050 ;
        RECT 857.400 813.600 858.600 871.950 ;
        RECT 872.400 844.200 873.600 883.950 ;
        RECT 881.400 883.050 882.600 884.100 ;
        RECT 887.400 883.050 888.600 889.950 ;
        RECT 877.950 880.950 880.050 883.050 ;
        RECT 880.950 880.950 883.050 883.050 ;
        RECT 883.950 880.950 886.050 883.050 ;
        RECT 886.950 880.950 889.050 883.050 ;
        RECT 865.950 840.000 868.050 844.050 ;
        RECT 871.950 842.100 874.050 844.200 ;
        RECT 878.400 844.050 879.600 880.950 ;
        RECT 877.950 841.950 880.050 844.050 ;
        RECT 884.400 841.050 885.600 880.950 ;
        RECT 886.950 841.950 889.050 844.050 ;
        RECT 866.400 838.050 867.600 840.000 ;
        RECT 871.950 838.950 874.050 841.050 ;
        RECT 883.950 838.950 886.050 841.050 ;
        RECT 872.400 838.050 873.600 838.950 ;
        RECT 862.950 835.950 865.050 838.050 ;
        RECT 865.950 835.950 868.050 838.050 ;
        RECT 868.950 835.950 871.050 838.050 ;
        RECT 871.950 835.950 874.050 838.050 ;
        RECT 863.400 834.900 864.600 835.950 ;
        RECT 869.400 834.900 870.600 835.950 ;
        RECT 862.950 832.800 865.050 834.900 ;
        RECT 868.950 832.800 871.050 834.900 ;
        RECT 868.950 820.950 871.050 823.050 ;
        RECT 857.400 812.400 861.600 813.600 ;
        RECT 850.950 806.100 853.050 808.200 ;
        RECT 851.400 805.050 852.600 806.100 ;
        RECT 817.950 802.950 820.050 805.050 ;
        RECT 820.950 802.950 823.050 805.050 ;
        RECT 823.950 802.950 826.050 805.050 ;
        RECT 826.950 802.950 829.050 805.050 ;
        RECT 844.950 802.950 847.050 805.050 ;
        RECT 847.950 802.950 850.050 805.050 ;
        RECT 850.950 802.950 853.050 805.050 ;
        RECT 853.950 802.950 856.050 805.050 ;
        RECT 818.400 801.000 819.600 802.950 ;
        RECT 824.400 801.900 825.600 802.950 ;
        RECT 817.950 796.950 820.050 801.000 ;
        RECT 823.950 799.800 826.050 801.900 ;
        RECT 848.400 799.050 849.600 802.950 ;
        RECT 854.400 801.900 855.600 802.950 ;
        RECT 853.950 799.800 856.050 801.900 ;
        RECT 860.400 801.600 861.600 812.400 ;
        RECT 869.400 805.050 870.600 820.950 ;
        RECT 874.950 806.100 877.050 808.200 ;
        RECT 883.950 806.100 886.050 808.200 ;
        RECT 875.400 805.050 876.600 806.100 ;
        RECT 868.950 802.950 871.050 805.050 ;
        RECT 871.950 802.950 874.050 805.050 ;
        RECT 874.950 802.950 877.050 805.050 ;
        RECT 877.950 802.950 880.050 805.050 ;
        RECT 872.400 801.900 873.600 802.950 ;
        RECT 857.400 800.400 861.600 801.600 ;
        RECT 847.950 796.950 850.050 799.050 ;
        RECT 835.950 790.950 838.050 793.050 ;
        RECT 811.950 784.950 814.050 787.050 ;
        RECT 814.950 761.100 817.050 763.200 ;
        RECT 820.950 761.100 823.050 763.200 ;
        RECT 826.950 763.050 829.050 763.200 ;
        RECT 826.950 761.100 832.050 763.050 ;
        RECT 815.400 760.050 816.600 761.100 ;
        RECT 821.400 760.050 822.600 761.100 ;
        RECT 828.000 760.950 832.050 761.100 ;
        RECT 832.950 760.950 835.050 763.050 ;
        RECT 814.950 757.950 817.050 760.050 ;
        RECT 817.950 757.950 820.050 760.050 ;
        RECT 820.950 757.950 823.050 760.050 ;
        RECT 823.950 757.950 826.050 760.050 ;
        RECT 818.400 756.900 819.600 757.950 ;
        RECT 824.400 756.900 825.600 757.950 ;
        RECT 833.400 757.050 834.600 760.950 ;
        RECT 811.950 756.600 814.050 756.900 ;
        RECT 809.400 755.400 814.050 756.600 ;
        RECT 811.950 754.800 814.050 755.400 ;
        RECT 817.950 754.800 820.050 756.900 ;
        RECT 823.950 754.800 826.050 756.900 ;
        RECT 832.950 754.950 835.050 757.050 ;
        RECT 812.400 751.050 813.600 754.800 ;
        RECT 811.950 748.950 814.050 751.050 ;
        RECT 817.950 748.950 820.050 751.050 ;
        RECT 805.950 742.950 808.050 745.050 ;
        RECT 775.950 736.950 778.050 739.050 ;
        RECT 781.950 733.950 784.050 736.050 ;
        RECT 793.950 733.950 796.050 736.050 ;
        RECT 811.950 733.950 814.050 736.050 ;
        RECT 773.400 728.400 777.600 729.600 ;
        RECT 767.400 727.050 768.600 728.100 ;
        RECT 760.950 724.950 763.050 727.050 ;
        RECT 766.950 724.950 769.050 727.050 ;
        RECT 769.950 724.950 772.050 727.050 ;
        RECT 770.400 718.050 771.600 724.950 ;
        RECT 769.950 715.950 772.050 718.050 ;
        RECT 776.400 700.050 777.600 728.400 ;
        RECT 760.950 697.950 763.050 700.050 ;
        RECT 775.950 697.950 778.050 700.050 ;
        RECT 739.950 676.800 742.050 678.900 ;
        RECT 745.950 676.800 748.050 678.900 ;
        RECT 757.950 676.950 760.050 679.050 ;
        RECT 740.400 654.600 741.600 676.800 ;
        RECT 761.400 672.600 762.600 697.950 ;
        RECT 775.950 691.950 778.050 694.050 ;
        RECT 776.400 685.200 777.600 691.950 ;
        RECT 769.950 683.100 772.050 685.200 ;
        RECT 775.950 683.100 778.050 685.200 ;
        RECT 770.400 682.050 771.600 683.100 ;
        RECT 776.400 682.050 777.600 683.100 ;
        RECT 766.950 679.950 769.050 682.050 ;
        RECT 769.950 679.950 772.050 682.050 ;
        RECT 772.950 679.950 775.050 682.050 ;
        RECT 775.950 679.950 778.050 682.050 ;
        RECT 758.400 671.400 762.600 672.600 ;
        RECT 748.950 655.050 751.050 655.200 ;
        RECT 740.400 653.400 744.600 654.600 ;
        RECT 743.400 649.050 744.600 653.400 ;
        RECT 745.950 653.100 751.050 655.050 ;
        RECT 745.950 652.950 750.000 653.100 ;
        RECT 748.950 649.950 751.050 652.050 ;
        RECT 749.400 649.050 750.600 649.950 ;
        RECT 742.950 646.950 745.050 649.050 ;
        RECT 745.950 646.950 748.050 649.050 ;
        RECT 748.950 646.950 751.050 649.050 ;
        RECT 751.950 646.950 754.050 649.050 ;
        RECT 733.950 643.950 736.050 646.050 ;
        RECT 746.400 645.000 747.600 646.950 ;
        RECT 752.400 645.900 753.600 646.950 ;
        RECT 745.950 640.950 748.050 645.000 ;
        RECT 751.950 643.800 754.050 645.900 ;
        RECT 748.950 640.950 751.050 643.050 ;
        RECT 745.950 637.800 748.050 639.900 ;
        RECT 728.400 633.000 732.600 633.600 ;
        RECT 727.950 632.400 732.600 633.000 ;
        RECT 727.950 628.950 730.050 632.400 ;
        RECT 742.950 631.950 745.050 634.050 ;
        RECT 739.950 627.600 742.050 631.050 ;
        RECT 737.400 627.000 742.050 627.600 ;
        RECT 737.400 626.400 741.600 627.000 ;
        RECT 724.950 619.950 727.050 622.050 ;
        RECT 733.950 613.950 736.050 616.050 ;
        RECT 719.400 605.400 723.600 606.600 ;
        RECT 724.950 606.000 727.050 610.050 ;
        RECT 734.400 607.050 735.600 613.950 ;
        RECT 710.400 604.050 711.600 605.100 ;
        RECT 709.950 601.950 712.050 604.050 ;
        RECT 700.950 598.950 703.050 601.050 ;
        RECT 706.950 598.950 709.050 601.050 ;
        RECT 694.950 595.950 697.050 598.050 ;
        RECT 701.400 580.050 702.600 598.950 ;
        RECT 707.400 595.050 708.600 598.950 ;
        RECT 706.950 592.950 709.050 595.050 ;
        RECT 700.950 577.950 703.050 580.050 ;
        RECT 674.400 571.050 675.600 572.100 ;
        RECT 670.950 568.950 673.050 571.050 ;
        RECT 673.950 568.950 676.050 571.050 ;
        RECT 679.950 568.950 682.050 571.050 ;
        RECT 671.400 568.050 672.600 568.950 ;
        RECT 667.950 566.400 672.600 568.050 ;
        RECT 667.950 565.950 672.000 566.400 ;
        RECT 680.400 559.050 681.600 568.950 ;
        RECT 682.950 565.950 685.050 568.050 ;
        RECT 673.950 556.950 676.050 559.050 ;
        RECT 679.950 556.950 682.050 559.050 ;
        RECT 664.950 547.950 667.050 550.050 ;
        RECT 670.950 547.950 673.050 550.050 ;
        RECT 662.400 530.400 666.600 531.600 ;
        RECT 665.400 529.200 666.600 530.400 ;
        RECT 659.400 526.050 660.600 528.000 ;
        RECT 664.950 527.100 667.050 529.200 ;
        RECT 665.400 526.050 666.600 527.100 ;
        RECT 658.950 523.950 661.050 526.050 ;
        RECT 661.950 523.950 664.050 526.050 ;
        RECT 664.950 523.950 667.050 526.050 ;
        RECT 662.400 514.050 663.600 523.950 ;
        RECT 664.950 517.950 667.050 520.050 ;
        RECT 661.950 511.950 664.050 514.050 ;
        RECT 665.400 505.050 666.600 517.950 ;
        RECT 664.950 502.950 667.050 505.050 ;
        RECT 671.400 502.050 672.600 547.950 ;
        RECT 674.400 529.050 675.600 556.950 ;
        RECT 679.950 547.950 682.050 550.050 ;
        RECT 673.950 526.950 676.050 529.050 ;
        RECT 680.400 526.050 681.600 547.950 ;
        RECT 683.400 532.050 684.600 565.950 ;
        RECT 686.400 562.050 687.600 572.100 ;
        RECT 691.950 571.950 694.050 574.050 ;
        RECT 697.950 572.100 700.050 574.200 ;
        RECT 707.400 574.050 708.600 592.950 ;
        RECT 712.950 583.950 715.050 586.050 ;
        RECT 698.400 571.050 699.600 572.100 ;
        RECT 706.950 571.950 709.050 574.050 ;
        RECT 713.400 571.050 714.600 583.950 ;
        RECT 719.400 571.050 720.600 605.400 ;
        RECT 725.400 604.050 726.600 606.000 ;
        RECT 733.950 604.950 736.050 607.050 ;
        RECT 724.950 601.950 727.050 604.050 ;
        RECT 727.950 601.950 730.050 604.050 ;
        RECT 728.400 600.900 729.600 601.950 ;
        RECT 727.950 598.800 730.050 600.900 ;
        RECT 733.950 595.950 736.050 600.900 ;
        RECT 724.950 592.950 727.050 595.050 ;
        RECT 721.950 589.950 724.050 592.050 ;
        RECT 722.400 583.050 723.600 589.950 ;
        RECT 721.950 580.950 724.050 583.050 ;
        RECT 725.400 577.050 726.600 592.950 ;
        RECT 733.950 592.800 736.050 594.900 ;
        RECT 727.950 586.950 730.050 589.050 ;
        RECT 724.950 574.950 727.050 577.050 ;
        RECT 694.950 568.950 697.050 571.050 ;
        RECT 697.950 568.950 700.050 571.050 ;
        RECT 700.950 568.950 703.050 571.050 ;
        RECT 712.950 568.950 715.050 571.050 ;
        RECT 715.950 568.950 718.050 571.050 ;
        RECT 718.950 568.950 721.050 571.050 ;
        RECT 721.950 568.950 724.050 571.050 ;
        RECT 695.400 567.900 696.600 568.950 ;
        RECT 694.950 565.800 697.050 567.900 ;
        RECT 685.950 559.950 688.050 562.050 ;
        RECT 686.400 541.050 687.600 559.950 ;
        RECT 701.400 559.050 702.600 568.950 ;
        RECT 705.000 567.900 709.050 568.050 ;
        RECT 703.950 565.950 709.050 567.900 ;
        RECT 703.950 565.800 706.050 565.950 ;
        RECT 716.400 562.050 717.600 568.950 ;
        RECT 722.400 567.900 723.600 568.950 ;
        RECT 721.950 565.800 724.050 567.900 ;
        RECT 715.950 559.950 718.050 562.050 ;
        RECT 724.950 561.600 727.050 562.050 ;
        RECT 728.400 561.600 729.600 586.950 ;
        RECT 734.400 574.050 735.600 592.800 ;
        RECT 737.400 586.050 738.600 626.400 ;
        RECT 743.400 622.050 744.600 631.950 ;
        RECT 746.400 628.050 747.600 637.800 ;
        RECT 749.400 637.050 750.600 640.950 ;
        RECT 754.950 637.950 757.050 640.050 ;
        RECT 748.950 634.950 751.050 637.050 ;
        RECT 745.950 625.950 748.050 628.050 ;
        RECT 742.950 619.950 745.050 622.050 ;
        RECT 749.400 610.050 750.600 634.950 ;
        RECT 755.400 634.050 756.600 637.950 ;
        RECT 754.950 631.950 757.050 634.050 ;
        RECT 758.400 631.050 759.600 671.400 ;
        RECT 767.400 670.050 768.600 679.950 ;
        RECT 773.400 678.000 774.600 679.950 ;
        RECT 772.950 673.950 775.050 678.000 ;
        RECT 782.400 670.050 783.600 733.950 ;
        RECT 787.950 728.100 790.050 730.200 ;
        RECT 788.400 727.050 789.600 728.100 ;
        RECT 794.400 727.050 795.600 733.950 ;
        RECT 812.400 727.050 813.600 733.950 ;
        RECT 818.400 727.050 819.600 748.950 ;
        RECT 829.950 742.950 832.050 745.050 ;
        RECT 823.950 733.950 826.050 736.050 ;
        RECT 787.950 724.950 790.050 727.050 ;
        RECT 790.950 724.950 793.050 727.050 ;
        RECT 793.950 724.950 796.050 727.050 ;
        RECT 796.950 724.950 799.050 727.050 ;
        RECT 808.950 724.950 811.050 727.050 ;
        RECT 811.950 724.950 814.050 727.050 ;
        RECT 814.950 724.950 817.050 727.050 ;
        RECT 817.950 724.950 820.050 727.050 ;
        RECT 791.400 715.050 792.600 724.950 ;
        RECT 797.400 723.000 798.600 724.950 ;
        RECT 796.950 718.950 799.050 723.000 ;
        RECT 802.950 718.950 805.050 721.050 ;
        RECT 790.950 712.950 793.050 715.050 ;
        RECT 793.950 700.950 796.050 703.050 ;
        RECT 787.950 684.000 790.050 688.050 ;
        RECT 788.400 682.050 789.600 684.000 ;
        RECT 794.400 682.050 795.600 700.950 ;
        RECT 803.400 688.050 804.600 718.950 ;
        RECT 805.950 715.950 808.050 718.050 ;
        RECT 802.950 685.950 805.050 688.050 ;
        RECT 787.950 679.950 790.050 682.050 ;
        RECT 790.950 679.950 793.050 682.050 ;
        RECT 793.950 679.950 796.050 682.050 ;
        RECT 796.950 679.950 799.050 682.050 ;
        RECT 791.400 678.900 792.600 679.950 ;
        RECT 797.400 679.050 798.600 679.950 ;
        RECT 790.950 676.800 793.050 678.900 ;
        RECT 797.400 677.400 802.050 679.050 ;
        RECT 798.000 676.950 802.050 677.400 ;
        RECT 760.950 667.950 763.050 670.050 ;
        RECT 766.950 667.950 769.050 670.050 ;
        RECT 781.950 667.950 784.050 670.050 ;
        RECT 761.400 661.050 762.600 667.950 ;
        RECT 791.400 667.050 792.600 676.800 ;
        RECT 803.400 676.050 804.600 685.950 ;
        RECT 806.400 679.050 807.600 715.950 ;
        RECT 809.400 712.050 810.600 724.950 ;
        RECT 815.400 723.900 816.600 724.950 ;
        RECT 824.400 724.050 825.600 733.950 ;
        RECT 826.950 728.100 829.050 730.200 ;
        RECT 814.950 718.950 817.050 723.900 ;
        RECT 823.950 721.950 826.050 724.050 ;
        RECT 808.950 709.950 811.050 712.050 ;
        RECT 827.400 703.050 828.600 728.100 ;
        RECT 826.950 700.950 829.050 703.050 ;
        RECT 814.950 683.100 817.050 685.200 ;
        RECT 820.950 683.100 823.050 685.200 ;
        RECT 826.950 683.100 829.050 685.200 ;
        RECT 815.400 682.050 816.600 683.100 ;
        RECT 821.400 682.050 822.600 683.100 ;
        RECT 811.950 679.950 814.050 682.050 ;
        RECT 814.950 679.950 817.050 682.050 ;
        RECT 817.950 679.950 820.050 682.050 ;
        RECT 820.950 679.950 823.050 682.050 ;
        RECT 805.950 676.950 808.050 679.050 ;
        RECT 812.400 678.000 813.600 679.950 ;
        RECT 796.950 673.950 799.050 676.050 ;
        RECT 802.950 673.950 805.050 676.050 ;
        RECT 811.950 673.950 814.050 678.000 ;
        RECT 772.950 664.950 775.050 667.050 ;
        RECT 790.950 664.950 793.050 667.050 ;
        RECT 760.950 658.950 763.050 661.050 ;
        RECT 763.950 655.050 766.050 658.050 ;
        RECT 760.950 654.000 766.050 655.050 ;
        RECT 760.950 653.400 765.600 654.000 ;
        RECT 760.950 652.950 765.000 653.400 ;
        RECT 766.950 650.100 769.050 652.200 ;
        RECT 767.400 649.050 768.600 650.100 ;
        RECT 773.400 649.050 774.600 664.950 ;
        RECT 781.950 655.950 784.050 658.050 ;
        RECT 763.950 646.950 766.050 649.050 ;
        RECT 766.950 646.950 769.050 649.050 ;
        RECT 769.950 646.950 772.050 649.050 ;
        RECT 772.950 646.950 775.050 649.050 ;
        RECT 760.950 643.950 763.050 646.050 ;
        RECT 764.400 645.000 765.600 646.950 ;
        RECT 757.950 628.950 760.050 631.050 ;
        RECT 757.950 625.800 760.050 627.900 ;
        RECT 758.400 615.600 759.600 625.800 ;
        RECT 761.400 619.050 762.600 643.950 ;
        RECT 763.950 640.950 766.050 645.000 ;
        RECT 760.950 616.950 763.050 619.050 ;
        RECT 764.400 616.050 765.600 640.950 ;
        RECT 766.950 637.950 769.050 640.050 ;
        RECT 767.400 631.050 768.600 637.950 ;
        RECT 770.400 637.050 771.600 646.950 ;
        RECT 782.400 646.050 783.600 655.950 ;
        RECT 790.950 650.100 793.050 652.200 ;
        RECT 791.400 649.050 792.600 650.100 ;
        RECT 797.400 649.050 798.600 673.950 ;
        RECT 805.950 664.950 808.050 667.050 ;
        RECT 802.950 649.950 805.050 652.050 ;
        RECT 787.950 646.950 790.050 649.050 ;
        RECT 790.950 646.950 793.050 649.050 ;
        RECT 793.950 646.950 796.050 649.050 ;
        RECT 796.950 646.950 799.050 649.050 ;
        RECT 781.950 643.950 784.050 646.050 ;
        RECT 788.400 645.900 789.600 646.950 ;
        RECT 787.950 645.600 790.050 645.900 ;
        RECT 785.400 644.400 790.050 645.600 ;
        RECT 769.950 634.950 772.050 637.050 ;
        RECT 766.950 628.950 769.050 631.050 ;
        RECT 769.950 619.950 772.050 622.050 ;
        RECT 766.950 616.950 769.050 619.050 ;
        RECT 758.400 614.400 762.600 615.600 ;
        RECT 739.950 607.950 742.050 610.050 ;
        RECT 748.950 607.950 751.050 610.050 ;
        RECT 740.400 595.050 741.600 607.950 ;
        RECT 742.950 606.600 747.000 607.050 ;
        RECT 742.950 604.950 747.600 606.600 ;
        RECT 751.950 606.000 754.050 610.050 ;
        RECT 746.400 604.050 747.600 604.950 ;
        RECT 752.400 604.050 753.600 606.000 ;
        RECT 757.950 604.950 760.050 610.050 ;
        RECT 745.950 601.950 748.050 604.050 ;
        RECT 748.950 601.950 751.050 604.050 ;
        RECT 751.950 601.950 754.050 604.050 ;
        RECT 754.950 601.950 757.050 604.050 ;
        RECT 742.950 595.950 745.050 601.050 ;
        RECT 739.950 592.950 742.050 595.050 ;
        RECT 749.400 592.050 750.600 601.950 ;
        RECT 755.400 600.900 756.600 601.950 ;
        RECT 754.950 598.800 757.050 600.900 ;
        RECT 761.400 592.050 762.600 614.400 ;
        RECT 763.950 613.950 766.050 616.050 ;
        RECT 767.400 607.050 768.600 616.950 ;
        RECT 766.950 604.950 769.050 607.050 ;
        RECT 770.400 604.050 771.600 619.950 ;
        RECT 775.950 610.950 778.050 613.050 ;
        RECT 776.400 604.050 777.600 610.950 ;
        RECT 781.950 605.100 784.050 607.200 ;
        RECT 785.400 607.050 786.600 644.400 ;
        RECT 787.950 643.800 790.050 644.400 ;
        RECT 794.400 631.050 795.600 646.950 ;
        RECT 793.950 628.950 796.050 631.050 ;
        RECT 787.950 619.950 790.050 622.050 ;
        RECT 782.400 604.050 783.600 605.100 ;
        RECT 784.950 604.950 787.050 607.050 ;
        RECT 769.950 601.950 772.050 604.050 ;
        RECT 772.950 601.950 775.050 604.050 ;
        RECT 775.950 601.950 778.050 604.050 ;
        RECT 778.950 601.950 781.050 604.050 ;
        RECT 781.950 601.950 784.050 604.050 ;
        RECT 766.950 598.950 769.050 601.050 ;
        RECT 748.950 589.950 751.050 592.050 ;
        RECT 760.950 589.950 763.050 592.050 ;
        RECT 736.950 583.950 739.050 586.050 ;
        RECT 751.950 583.950 754.050 586.050 ;
        RECT 736.950 574.950 739.050 580.050 ;
        RECT 733.950 571.950 736.050 574.050 ;
        RECT 742.950 572.100 745.050 574.200 ;
        RECT 743.400 571.050 744.600 572.100 ;
        RECT 739.950 568.950 742.050 571.050 ;
        RECT 742.950 568.950 745.050 571.050 ;
        RECT 745.950 568.950 748.050 571.050 ;
        RECT 740.400 562.050 741.600 568.950 ;
        RECT 746.400 568.050 747.600 568.950 ;
        RECT 746.400 566.400 751.050 568.050 ;
        RECT 747.000 565.950 751.050 566.400 ;
        RECT 745.950 562.950 748.050 565.050 ;
        RECT 724.950 560.400 729.600 561.600 ;
        RECT 724.950 559.950 727.050 560.400 ;
        RECT 739.950 559.950 742.050 562.050 ;
        RECT 700.950 556.950 703.050 559.050 ;
        RECT 685.950 538.950 688.050 541.050 ;
        RECT 701.400 538.050 702.600 556.950 ;
        RECT 715.950 547.950 718.050 550.050 ;
        RECT 712.950 544.950 715.050 547.050 ;
        RECT 700.950 535.950 703.050 538.050 ;
        RECT 682.950 529.950 685.050 532.050 ;
        RECT 685.950 528.000 688.050 532.050 ;
        RECT 691.950 529.950 694.050 532.050 ;
        RECT 686.400 526.050 687.600 528.000 ;
        RECT 676.950 523.950 679.050 526.050 ;
        RECT 679.950 523.950 682.050 526.050 ;
        RECT 682.950 523.950 685.050 526.050 ;
        RECT 685.950 523.950 688.050 526.050 ;
        RECT 673.950 520.950 676.050 523.050 ;
        RECT 670.950 499.950 673.050 502.050 ;
        RECT 661.950 494.100 664.050 496.200 ;
        RECT 667.950 494.100 670.050 496.200 ;
        RECT 662.400 493.050 663.600 494.100 ;
        RECT 668.400 493.050 669.600 494.100 ;
        RECT 658.950 490.950 661.050 493.050 ;
        RECT 661.950 490.950 664.050 493.050 ;
        RECT 664.950 490.950 667.050 493.050 ;
        RECT 667.950 490.950 670.050 493.050 ;
        RECT 653.400 488.400 657.600 489.600 ;
        RECT 637.950 485.400 645.600 486.600 ;
        RECT 637.950 484.950 642.600 485.400 ;
        RECT 635.400 481.050 636.600 484.950 ;
        RECT 637.950 484.650 640.050 484.950 ;
        RECT 634.950 478.950 637.050 481.050 ;
        RECT 631.950 475.950 634.050 478.050 ;
        RECT 635.400 450.600 636.600 478.950 ;
        RECT 641.400 451.200 642.600 484.950 ;
        RECT 649.950 475.950 652.050 478.050 ;
        RECT 626.400 449.400 630.600 450.600 ;
        RECT 632.400 449.400 636.600 450.600 ;
        RECT 617.400 448.050 618.600 449.100 ;
        RECT 613.950 445.950 616.050 448.050 ;
        RECT 616.950 445.950 619.050 448.050 ;
        RECT 619.950 445.950 622.050 448.050 ;
        RECT 607.950 439.950 610.050 442.050 ;
        RECT 614.400 430.050 615.600 445.950 ;
        RECT 620.400 444.000 621.600 445.950 ;
        RECT 619.950 439.950 622.050 444.000 ;
        RECT 613.950 427.950 616.050 430.050 ;
        RECT 619.800 427.950 621.900 430.050 ;
        RECT 622.950 427.950 625.050 430.050 ;
        RECT 604.950 415.950 607.050 418.050 ;
        RECT 610.950 417.000 613.050 421.050 ;
        RECT 611.400 415.050 612.600 417.000 ;
        RECT 616.950 415.950 619.050 421.050 ;
        RECT 620.400 418.050 621.600 427.950 ;
        RECT 619.950 415.950 622.050 418.050 ;
        RECT 607.950 412.950 610.050 415.050 ;
        RECT 610.950 412.950 613.050 415.050 ;
        RECT 604.950 409.950 607.050 412.050 ;
        RECT 605.400 397.050 606.600 409.950 ;
        RECT 608.400 406.050 609.600 412.950 ;
        RECT 619.950 412.800 622.050 414.900 ;
        RECT 607.950 403.950 610.050 406.050 ;
        RECT 616.950 400.950 619.050 403.050 ;
        RECT 617.400 397.050 618.600 400.950 ;
        RECT 604.950 394.950 607.050 397.050 ;
        RECT 616.950 394.950 619.050 397.050 ;
        RECT 604.950 379.950 607.050 382.050 ;
        RECT 601.950 373.950 604.050 376.050 ;
        RECT 598.950 371.100 601.050 373.200 ;
        RECT 599.400 370.050 600.600 371.100 ;
        RECT 605.400 370.050 606.600 379.950 ;
        RECT 620.400 379.050 621.600 412.800 ;
        RECT 623.400 388.050 624.600 427.950 ;
        RECT 626.400 418.050 627.600 449.400 ;
        RECT 632.400 448.050 633.600 449.400 ;
        RECT 640.950 449.100 643.050 451.200 ;
        RECT 641.400 448.050 642.600 449.100 ;
        RECT 631.950 445.950 634.050 448.050 ;
        RECT 640.950 445.950 643.050 448.050 ;
        RECT 634.800 442.950 636.900 445.050 ;
        RECT 635.400 424.050 636.600 442.950 ;
        RECT 628.950 421.950 631.050 424.050 ;
        RECT 634.950 421.950 637.050 424.050 ;
        RECT 625.950 415.950 628.050 418.050 ;
        RECT 629.400 415.050 630.600 421.950 ;
        RECT 650.400 421.050 651.600 475.950 ;
        RECT 656.400 451.050 657.600 488.400 ;
        RECT 659.400 460.050 660.600 490.950 ;
        RECT 665.400 489.900 666.600 490.950 ;
        RECT 664.950 487.800 667.050 489.900 ;
        RECT 670.950 478.950 673.050 481.050 ;
        RECT 658.950 457.950 661.050 460.050 ;
        RECT 664.950 454.950 667.050 457.050 ;
        RECT 652.800 448.950 654.900 451.050 ;
        RECT 655.800 448.950 657.900 451.050 ;
        RECT 658.950 449.100 661.050 451.200 ;
        RECT 653.400 424.050 654.600 448.950 ;
        RECT 659.400 448.050 660.600 449.100 ;
        RECT 665.400 448.050 666.600 454.950 ;
        RECT 671.400 448.050 672.600 478.950 ;
        RECT 674.400 472.050 675.600 520.950 ;
        RECT 677.400 505.050 678.600 523.950 ;
        RECT 683.400 522.900 684.600 523.950 ;
        RECT 682.950 520.800 685.050 522.900 ;
        RECT 692.400 511.050 693.600 529.950 ;
        RECT 706.950 527.100 709.050 529.200 ;
        RECT 707.400 526.050 708.600 527.100 ;
        RECT 706.950 523.950 709.050 526.050 ;
        RECT 713.400 514.050 714.600 544.950 ;
        RECT 694.950 511.950 697.050 514.050 ;
        RECT 700.950 511.950 703.050 514.050 ;
        RECT 712.950 511.950 715.050 514.050 ;
        RECT 716.400 513.600 717.600 547.950 ;
        RECT 725.400 526.050 726.600 559.950 ;
        RECT 746.400 556.050 747.600 562.950 ;
        RECT 748.950 556.950 751.050 559.050 ;
        RECT 745.950 553.950 748.050 556.050 ;
        RECT 749.400 553.050 750.600 556.950 ;
        RECT 748.950 550.950 751.050 553.050 ;
        RECT 742.950 547.950 745.050 550.050 ;
        RECT 730.950 541.950 733.050 544.050 ;
        RECT 736.950 541.950 739.050 544.050 ;
        RECT 731.400 526.050 732.600 541.950 ;
        RECT 721.950 523.950 724.050 526.050 ;
        RECT 724.950 523.950 727.050 526.050 ;
        RECT 727.950 523.950 730.050 526.050 ;
        RECT 730.950 523.950 733.050 526.050 ;
        RECT 718.950 520.950 721.050 523.050 ;
        RECT 719.400 517.050 720.600 520.950 ;
        RECT 718.950 514.950 721.050 517.050 ;
        RECT 722.400 513.600 723.600 523.950 ;
        RECT 716.400 512.400 723.600 513.600 ;
        RECT 691.950 508.950 694.050 511.050 ;
        RECT 682.950 505.950 685.050 508.050 ;
        RECT 676.950 502.950 679.050 505.050 ;
        RECT 683.400 499.050 684.600 505.950 ;
        RECT 695.400 505.050 696.600 511.950 ;
        RECT 685.950 502.950 688.050 505.050 ;
        RECT 694.950 502.950 697.050 505.050 ;
        RECT 697.950 502.950 700.050 505.050 ;
        RECT 676.950 496.950 679.050 499.050 ;
        RECT 682.950 496.950 685.050 499.050 ;
        RECT 673.950 469.950 676.050 472.050 ;
        RECT 674.400 451.200 675.600 469.950 ;
        RECT 677.400 463.050 678.600 496.950 ;
        RECT 686.400 493.050 687.600 502.950 ;
        RECT 694.950 493.950 697.050 496.050 ;
        RECT 682.950 490.950 685.050 493.050 ;
        RECT 685.950 490.950 688.050 493.050 ;
        RECT 688.950 490.950 691.050 493.050 ;
        RECT 683.400 489.900 684.600 490.950 ;
        RECT 689.400 489.900 690.600 490.950 ;
        RECT 695.400 489.900 696.600 493.950 ;
        RECT 682.950 487.800 685.050 489.900 ;
        RECT 688.950 487.800 691.050 489.900 ;
        RECT 694.950 484.950 697.050 489.900 ;
        RECT 698.400 481.050 699.600 502.950 ;
        RECT 701.400 490.050 702.600 511.950 ;
        RECT 716.400 508.050 717.600 512.400 ;
        RECT 715.950 505.950 718.050 508.050 ;
        RECT 703.950 499.950 706.050 505.050 ;
        RECT 706.950 499.950 709.050 502.050 ;
        RECT 721.950 499.950 724.050 502.050 ;
        RECT 707.400 493.050 708.600 499.950 ;
        RECT 712.950 494.100 715.050 496.200 ;
        RECT 713.400 493.050 714.600 494.100 ;
        RECT 706.950 490.950 709.050 493.050 ;
        RECT 709.950 490.950 712.050 493.050 ;
        RECT 712.950 490.950 715.050 493.050 ;
        RECT 715.950 490.950 718.050 493.050 ;
        RECT 700.950 487.950 703.050 490.050 ;
        RECT 710.400 489.900 711.600 490.950 ;
        RECT 709.950 487.800 712.050 489.900 ;
        RECT 706.950 484.950 709.050 487.050 ;
        RECT 697.950 478.950 700.050 481.050 ;
        RECT 707.400 478.050 708.600 484.950 ;
        RECT 691.950 475.950 694.050 478.050 ;
        RECT 706.950 475.950 709.050 478.050 ;
        RECT 676.950 460.950 679.050 463.050 ;
        RECT 676.950 454.950 679.050 457.050 ;
        RECT 673.950 449.100 676.050 451.200 ;
        RECT 658.950 445.950 661.050 448.050 ;
        RECT 664.950 445.950 667.050 448.050 ;
        RECT 670.950 445.950 673.050 448.050 ;
        RECT 655.950 427.950 658.050 430.050 ;
        RECT 652.950 421.950 655.050 424.050 ;
        RECT 640.950 418.950 643.050 421.050 ;
        RECT 649.950 418.950 652.050 421.050 ;
        RECT 656.400 420.600 657.600 427.950 ;
        RECT 661.950 421.950 664.050 424.050 ;
        RECT 673.950 421.950 676.050 424.050 ;
        RECT 653.400 419.400 657.600 420.600 ;
        RECT 634.950 416.100 637.050 418.200 ;
        RECT 635.400 415.050 636.600 416.100 ;
        RECT 628.950 412.950 631.050 415.050 ;
        RECT 631.950 412.950 634.050 415.050 ;
        RECT 634.950 412.950 637.050 415.050 ;
        RECT 625.950 409.950 628.050 412.050 ;
        RECT 626.400 391.050 627.600 409.950 ;
        RECT 625.950 388.950 628.050 391.050 ;
        RECT 622.950 385.950 625.050 388.050 ;
        RECT 623.400 379.050 624.600 385.950 ;
        RECT 632.400 385.050 633.600 412.950 ;
        RECT 641.400 409.050 642.600 418.950 ;
        RECT 653.400 415.050 654.600 419.400 ;
        RECT 649.950 412.950 652.050 415.050 ;
        RECT 652.950 412.950 655.050 415.050 ;
        RECT 650.400 411.000 651.600 412.950 ;
        RECT 637.950 403.950 640.050 406.050 ;
        RECT 640.950 403.950 643.050 409.050 ;
        RECT 649.950 406.950 652.050 411.000 ;
        RECT 662.400 409.050 663.600 421.950 ;
        RECT 674.400 415.050 675.600 421.950 ;
        RECT 677.400 421.050 678.600 454.950 ;
        RECT 679.950 448.950 682.050 451.050 ;
        RECT 680.400 427.050 681.600 448.950 ;
        RECT 692.400 448.050 693.600 475.950 ;
        RECT 700.950 466.950 703.050 469.050 ;
        RECT 701.400 463.050 702.600 466.950 ;
        RECT 697.800 460.950 699.900 463.050 ;
        RECT 700.950 460.950 703.050 463.050 ;
        RECT 688.950 445.950 691.050 448.050 ;
        RECT 691.950 445.950 694.050 448.050 ;
        RECT 689.400 444.900 690.600 445.950 ;
        RECT 698.400 444.900 699.600 460.950 ;
        RECT 710.400 453.600 711.600 487.800 ;
        RECT 716.400 484.050 717.600 490.950 ;
        RECT 715.950 481.950 718.050 484.050 ;
        RECT 707.400 452.400 711.600 453.600 ;
        RECT 707.400 448.050 708.600 452.400 ;
        RECT 712.950 449.100 715.050 451.200 ;
        RECT 713.400 448.050 714.600 449.100 ;
        RECT 703.950 445.950 706.050 448.050 ;
        RECT 706.950 445.950 709.050 448.050 ;
        RECT 709.950 445.950 712.050 448.050 ;
        RECT 712.950 445.950 715.050 448.050 ;
        RECT 704.400 444.900 705.600 445.950 ;
        RECT 688.950 442.800 691.050 444.900 ;
        RECT 697.950 442.800 700.050 444.900 ;
        RECT 703.950 442.800 706.050 444.900 ;
        RECT 689.400 436.050 690.600 442.800 ;
        RECT 710.400 439.050 711.600 445.950 ;
        RECT 709.950 436.950 712.050 439.050 ;
        RECT 688.950 433.950 691.050 436.050 ;
        RECT 715.950 427.950 718.050 430.050 ;
        RECT 679.950 424.950 682.050 427.050 ;
        RECT 688.950 421.950 691.050 424.050 ;
        RECT 676.950 418.950 679.050 421.050 ;
        RECT 689.400 418.200 690.600 421.950 ;
        RECT 679.950 416.100 682.050 418.200 ;
        RECT 680.400 415.050 681.600 416.100 ;
        RECT 685.800 415.950 687.900 418.050 ;
        RECT 688.950 416.100 691.050 418.200 ;
        RECT 697.950 416.100 700.050 418.200 ;
        RECT 703.950 416.100 706.050 418.200 ;
        RECT 712.950 416.100 715.050 418.200 ;
        RECT 670.950 412.950 673.050 415.050 ;
        RECT 673.950 412.950 676.050 415.050 ;
        RECT 676.950 412.950 679.050 415.050 ;
        RECT 679.950 412.950 682.050 415.050 ;
        RECT 667.950 409.950 670.050 412.050 ;
        RECT 671.400 411.900 672.600 412.950 ;
        RECT 661.950 406.950 664.050 409.050 ;
        RECT 634.950 400.950 637.050 403.050 ;
        RECT 631.950 382.950 634.050 385.050 ;
        RECT 613.950 376.950 616.050 379.050 ;
        RECT 616.950 376.950 619.050 379.050 ;
        RECT 619.950 376.950 622.050 379.050 ;
        RECT 622.950 376.950 625.050 379.050 ;
        RECT 614.400 370.050 615.600 376.950 ;
        RECT 595.950 367.950 598.050 370.050 ;
        RECT 598.950 367.950 601.050 370.050 ;
        RECT 601.950 367.950 604.050 370.050 ;
        RECT 604.950 367.950 607.050 370.050 ;
        RECT 607.950 367.950 610.050 370.050 ;
        RECT 613.950 367.950 616.050 370.050 ;
        RECT 596.400 366.900 597.600 367.950 ;
        RECT 595.950 364.800 598.050 366.900 ;
        RECT 602.400 349.050 603.600 367.950 ;
        RECT 608.400 367.050 609.600 367.950 ;
        RECT 608.400 365.400 613.050 367.050 ;
        RECT 609.000 364.950 613.050 365.400 ;
        RECT 613.950 355.950 616.050 358.050 ;
        RECT 601.950 346.950 604.050 349.050 ;
        RECT 599.400 342.900 600.600 345.450 ;
        RECT 595.200 339.900 597.300 341.700 ;
        RECT 599.100 340.800 601.200 342.900 ;
        RECT 602.400 342.300 604.500 344.400 ;
        RECT 593.700 338.700 602.250 339.900 ;
        RECT 590.400 334.950 592.500 337.050 ;
        RECT 590.400 332.400 591.600 334.950 ;
        RECT 593.700 329.700 594.600 338.700 ;
        RECT 600.150 337.800 602.250 338.700 ;
        RECT 603.150 336.900 604.050 342.300 ;
        RECT 610.950 340.950 613.050 343.050 ;
        RECT 605.400 337.050 606.600 339.600 ;
        RECT 611.400 337.050 612.600 340.950 ;
        RECT 597.300 335.700 604.050 336.900 ;
        RECT 597.300 333.300 598.200 335.700 ;
        RECT 596.100 331.200 598.200 333.300 ;
        RECT 599.100 332.100 601.200 334.200 ;
        RECT 592.800 327.600 594.900 329.700 ;
        RECT 599.400 329.550 600.600 332.100 ;
        RECT 603.000 328.500 604.050 335.700 ;
        RECT 604.950 334.950 607.050 337.050 ;
        RECT 610.950 334.950 613.050 337.050 ;
        RECT 602.400 326.400 604.500 328.500 ;
        RECT 598.950 316.950 601.050 319.050 ;
        RECT 586.950 313.950 589.050 316.050 ;
        RECT 583.950 310.950 586.050 313.050 ;
        RECT 595.950 307.950 598.050 310.050 ;
        RECT 589.950 298.950 592.050 301.050 ;
        RECT 590.400 295.200 591.600 298.950 ;
        RECT 565.950 293.100 568.050 295.200 ;
        RECT 566.400 292.050 567.600 293.100 ;
        RECT 574.950 292.950 577.050 295.050 ;
        RECT 580.950 293.100 583.050 295.200 ;
        RECT 589.950 293.100 592.050 295.200 ;
        RECT 565.950 289.950 568.050 292.050 ;
        RECT 568.950 289.950 571.050 292.050 ;
        RECT 569.400 288.900 570.600 289.950 ;
        RECT 559.950 286.800 562.050 288.900 ;
        RECT 568.950 286.800 571.050 288.900 ;
        RECT 575.400 277.050 576.600 292.950 ;
        RECT 581.400 292.050 582.600 293.100 ;
        RECT 590.400 292.050 591.600 293.100 ;
        RECT 580.950 289.950 583.050 292.050 ;
        RECT 583.950 289.950 586.050 292.050 ;
        RECT 589.950 289.950 592.050 292.050 ;
        RECT 584.400 288.000 585.600 289.950 ;
        RECT 583.950 283.950 586.050 288.000 ;
        RECT 574.950 274.950 577.050 277.050 ;
        RECT 596.400 271.050 597.600 307.950 ;
        RECT 599.400 274.050 600.600 316.950 ;
        RECT 607.950 293.100 610.050 295.200 ;
        RECT 608.400 292.050 609.600 293.100 ;
        RECT 604.950 289.950 607.050 292.050 ;
        RECT 607.950 289.950 610.050 292.050 ;
        RECT 605.400 288.900 606.600 289.950 ;
        RECT 604.950 286.800 607.050 288.900 ;
        RECT 614.400 286.050 615.600 355.950 ;
        RECT 617.400 333.900 618.600 376.950 ;
        RECT 619.950 370.950 622.050 375.900 ;
        RECT 631.950 373.950 634.050 376.050 ;
        RECT 625.950 371.100 628.050 373.200 ;
        RECT 626.400 370.050 627.600 371.100 ;
        RECT 622.950 367.950 625.050 370.050 ;
        RECT 625.950 367.950 628.050 370.050 ;
        RECT 623.400 366.900 624.600 367.950 ;
        RECT 632.400 366.900 633.600 373.950 ;
        RECT 622.950 364.800 625.050 366.900 ;
        RECT 631.950 364.800 634.050 366.900 ;
        RECT 623.400 343.050 624.600 364.800 ;
        RECT 631.950 358.950 634.050 361.050 ;
        RECT 622.950 340.950 625.050 343.050 ;
        RECT 625.950 338.100 628.050 340.200 ;
        RECT 626.400 337.050 627.600 338.100 ;
        RECT 632.400 337.050 633.600 358.950 ;
        RECT 635.400 358.050 636.600 400.950 ;
        RECT 638.400 366.600 639.600 403.950 ;
        RECT 643.950 397.950 646.050 400.050 ;
        RECT 644.400 370.050 645.600 397.950 ;
        RECT 650.400 382.050 651.600 406.950 ;
        RECT 668.400 406.050 669.600 409.950 ;
        RECT 670.950 406.950 673.050 411.900 ;
        RECT 677.400 406.050 678.600 412.950 ;
        RECT 682.950 406.950 685.050 409.050 ;
        RECT 667.950 403.950 670.050 406.050 ;
        RECT 676.950 403.950 679.050 406.050 ;
        RECT 679.950 391.950 682.050 394.050 ;
        RECT 658.950 388.950 661.050 391.050 ;
        RECT 649.950 379.950 652.050 382.050 ;
        RECT 649.950 376.800 652.050 378.900 ;
        RECT 650.400 370.050 651.600 376.800 ;
        RECT 643.950 367.950 646.050 370.050 ;
        RECT 646.950 367.950 649.050 370.050 ;
        RECT 649.950 367.950 652.050 370.050 ;
        RECT 652.950 367.950 655.050 370.050 ;
        RECT 638.400 365.400 642.600 366.600 ;
        RECT 634.950 355.950 637.050 358.050 ;
        RECT 637.950 337.950 640.050 340.050 ;
        RECT 622.950 334.950 625.050 337.050 ;
        RECT 625.950 334.950 628.050 337.050 ;
        RECT 628.950 334.950 631.050 337.050 ;
        RECT 631.950 334.950 634.050 337.050 ;
        RECT 616.950 331.800 619.050 333.900 ;
        RECT 617.400 286.050 618.600 331.800 ;
        RECT 623.400 328.050 624.600 334.950 ;
        RECT 629.400 333.900 630.600 334.950 ;
        RECT 628.950 331.800 631.050 333.900 ;
        RECT 622.950 325.950 625.050 328.050 ;
        RECT 638.400 316.050 639.600 337.950 ;
        RECT 641.400 333.600 642.600 365.400 ;
        RECT 643.950 361.950 646.050 364.050 ;
        RECT 644.400 352.050 645.600 361.950 ;
        RECT 647.400 355.050 648.600 367.950 ;
        RECT 653.400 361.050 654.600 367.950 ;
        RECT 652.950 358.950 655.050 361.050 ;
        RECT 646.950 352.950 649.050 355.050 ;
        RECT 652.950 352.950 655.050 355.050 ;
        RECT 643.950 349.950 646.050 352.050 ;
        RECT 646.950 338.100 649.050 340.200 ;
        RECT 647.400 337.050 648.600 338.100 ;
        RECT 653.400 337.050 654.600 352.950 ;
        RECT 659.400 340.050 660.600 388.950 ;
        RECT 664.950 376.950 667.050 379.050 ;
        RECT 665.400 370.050 666.600 376.950 ;
        RECT 680.400 370.050 681.600 391.950 ;
        RECT 664.950 367.950 667.050 370.050 ;
        RECT 667.950 367.950 670.050 370.050 ;
        RECT 679.950 367.950 682.050 370.050 ;
        RECT 668.400 361.050 669.600 367.950 ;
        RECT 667.950 358.950 670.050 361.050 ;
        RECT 683.400 354.600 684.600 406.950 ;
        RECT 686.400 394.050 687.600 415.950 ;
        RECT 689.400 406.050 690.600 416.100 ;
        RECT 698.400 415.050 699.600 416.100 ;
        RECT 704.400 415.050 705.600 416.100 ;
        RECT 694.950 412.950 697.050 415.050 ;
        RECT 697.950 412.950 700.050 415.050 ;
        RECT 700.950 412.950 703.050 415.050 ;
        RECT 703.950 412.950 706.050 415.050 ;
        RECT 706.950 412.950 709.050 415.050 ;
        RECT 695.400 411.900 696.600 412.950 ;
        RECT 694.950 409.800 697.050 411.900 ;
        RECT 688.950 403.950 691.050 406.050 ;
        RECT 701.400 397.050 702.600 412.950 ;
        RECT 700.950 394.950 703.050 397.050 ;
        RECT 707.400 394.050 708.600 412.950 ;
        RECT 713.400 411.600 714.600 416.100 ;
        RECT 710.400 410.400 714.600 411.600 ;
        RECT 685.950 391.950 688.050 394.050 ;
        RECT 706.950 391.950 709.050 394.050 ;
        RECT 706.950 384.600 709.050 385.050 ;
        RECT 710.400 384.600 711.600 410.400 ;
        RECT 716.400 409.050 717.600 427.950 ;
        RECT 718.950 424.950 721.050 427.050 ;
        RECT 719.400 411.900 720.600 424.950 ;
        RECT 722.400 418.050 723.600 499.950 ;
        RECT 724.950 496.950 727.050 499.050 ;
        RECT 725.400 472.050 726.600 496.950 ;
        RECT 728.400 496.200 729.600 523.950 ;
        RECT 737.400 499.050 738.600 541.950 ;
        RECT 739.950 529.950 742.050 532.050 ;
        RECT 740.400 514.050 741.600 529.950 ;
        RECT 743.400 529.050 744.600 547.950 ;
        RECT 742.950 526.950 745.050 529.050 ;
        RECT 749.400 528.600 750.600 550.950 ;
        RECT 752.400 532.050 753.600 583.950 ;
        RECT 754.950 580.950 757.050 583.050 ;
        RECT 755.400 574.050 756.600 580.950 ;
        RECT 754.950 571.950 757.050 574.050 ;
        RECT 760.950 572.100 763.050 574.200 ;
        RECT 761.400 571.050 762.600 572.100 ;
        RECT 767.400 571.050 768.600 598.950 ;
        RECT 773.400 597.600 774.600 601.950 ;
        RECT 770.400 596.400 774.600 597.600 ;
        RECT 770.400 574.050 771.600 596.400 ;
        RECT 772.950 592.950 775.050 595.050 ;
        RECT 769.950 571.950 772.050 574.050 ;
        RECT 757.950 568.950 760.050 571.050 ;
        RECT 760.950 568.950 763.050 571.050 ;
        RECT 763.950 568.950 766.050 571.050 ;
        RECT 766.950 568.950 769.050 571.050 ;
        RECT 754.950 559.950 757.050 562.050 ;
        RECT 755.400 553.050 756.600 559.950 ;
        RECT 754.950 550.950 757.050 553.050 ;
        RECT 755.400 544.050 756.600 550.950 ;
        RECT 754.950 541.950 757.050 544.050 ;
        RECT 751.950 529.950 754.050 532.050 ;
        RECT 746.400 527.400 750.600 528.600 ;
        RECT 746.400 526.050 747.600 527.400 ;
        RECT 755.400 526.050 756.600 541.950 ;
        RECT 758.400 538.050 759.600 568.950 ;
        RECT 764.400 562.050 765.600 568.950 ;
        RECT 766.950 562.950 769.050 565.050 ;
        RECT 769.950 562.950 772.050 568.050 ;
        RECT 763.950 559.950 766.050 562.050 ;
        RECT 767.400 553.050 768.600 562.950 ;
        RECT 766.950 550.950 769.050 553.050 ;
        RECT 766.950 547.800 769.050 549.900 ;
        RECT 763.950 544.950 766.050 547.050 ;
        RECT 760.950 538.950 763.050 541.050 ;
        RECT 757.950 535.950 760.050 538.050 ;
        RECT 745.950 523.950 748.050 526.050 ;
        RECT 751.950 523.950 754.050 526.050 ;
        RECT 754.950 523.950 757.050 526.050 ;
        RECT 742.950 520.950 745.050 523.050 ;
        RECT 739.950 511.950 742.050 514.050 ;
        RECT 739.950 505.950 742.050 508.050 ;
        RECT 736.950 496.950 739.050 499.050 ;
        RECT 727.950 494.100 730.050 496.200 ;
        RECT 733.950 494.100 736.050 496.200 ;
        RECT 734.400 493.050 735.600 494.100 ;
        RECT 740.400 493.050 741.600 505.950 ;
        RECT 743.400 495.600 744.600 520.950 ;
        RECT 752.400 517.050 753.600 523.950 ;
        RECT 751.950 516.600 754.050 517.050 ;
        RECT 751.950 515.400 756.600 516.600 ;
        RECT 751.950 514.950 754.050 515.400 ;
        RECT 748.950 511.950 751.050 514.050 ;
        RECT 743.400 494.400 747.600 495.600 ;
        RECT 730.950 490.950 733.050 493.050 ;
        RECT 733.950 490.950 736.050 493.050 ;
        RECT 736.950 490.950 739.050 493.050 ;
        RECT 739.950 490.950 742.050 493.050 ;
        RECT 731.400 489.900 732.600 490.950 ;
        RECT 730.950 487.800 733.050 489.900 ;
        RECT 737.400 487.050 738.600 490.950 ;
        RECT 736.950 484.950 739.050 487.050 ;
        RECT 724.950 469.950 727.050 472.050 ;
        RECT 727.950 460.950 730.050 463.050 ;
        RECT 728.400 448.050 729.600 460.950 ;
        RECT 737.400 460.050 738.600 484.950 ;
        RECT 746.400 474.600 747.600 494.400 ;
        RECT 743.400 473.400 747.600 474.600 ;
        RECT 743.400 462.600 744.600 473.400 ;
        RECT 745.950 469.950 748.050 472.050 ;
        RECT 740.400 461.400 744.600 462.600 ;
        RECT 736.950 457.950 739.050 460.050 ;
        RECT 727.950 445.950 730.050 448.050 ;
        RECT 730.950 445.950 733.050 448.050 ;
        RECT 724.950 442.950 727.050 445.050 ;
        RECT 725.400 427.050 726.600 442.950 ;
        RECT 724.950 424.950 727.050 427.050 ;
        RECT 731.400 421.050 732.600 445.950 ;
        RECT 736.950 436.950 739.050 439.050 ;
        RECT 730.950 418.950 733.050 421.050 ;
        RECT 737.400 418.050 738.600 436.950 ;
        RECT 740.400 430.050 741.600 461.400 ;
        RECT 742.950 457.950 745.050 460.050 ;
        RECT 743.400 445.050 744.600 457.950 ;
        RECT 742.950 442.950 745.050 445.050 ;
        RECT 746.400 430.050 747.600 469.950 ;
        RECT 749.400 466.050 750.600 511.950 ;
        RECT 755.400 496.050 756.600 515.400 ;
        RECT 754.950 493.950 757.050 496.050 ;
        RECT 761.400 493.050 762.600 538.950 ;
        RECT 764.400 502.050 765.600 544.950 ;
        RECT 767.400 538.050 768.600 547.800 ;
        RECT 773.400 547.050 774.600 592.950 ;
        RECT 779.400 592.050 780.600 601.950 ;
        RECT 784.950 598.950 787.050 601.050 ;
        RECT 785.400 595.050 786.600 598.950 ;
        RECT 788.400 595.050 789.600 619.950 ;
        RECT 794.400 619.050 795.600 628.950 ;
        RECT 793.950 616.950 796.050 619.050 ;
        RECT 793.950 613.800 796.050 615.900 ;
        RECT 790.950 607.950 793.050 613.050 ;
        RECT 794.400 607.050 795.600 613.800 ;
        RECT 796.950 607.950 799.050 613.050 ;
        RECT 803.400 607.050 804.600 649.950 ;
        RECT 806.400 634.050 807.600 664.950 ;
        RECT 811.950 658.950 814.050 661.050 ;
        RECT 812.400 649.050 813.600 658.950 ;
        RECT 818.400 655.050 819.600 679.950 ;
        RECT 823.950 673.950 826.050 676.050 ;
        RECT 817.950 652.950 820.050 655.050 ;
        RECT 811.950 646.950 814.050 649.050 ;
        RECT 824.400 640.050 825.600 673.950 ;
        RECT 827.400 673.050 828.600 683.100 ;
        RECT 826.950 670.950 829.050 673.050 ;
        RECT 830.400 667.050 831.600 742.950 ;
        RECT 833.400 742.050 834.600 754.950 ;
        RECT 836.400 751.050 837.600 790.950 ;
        RECT 848.400 775.050 849.600 796.950 ;
        RECT 847.950 772.950 850.050 775.050 ;
        RECT 841.950 762.600 846.000 763.050 ;
        RECT 841.950 760.950 846.600 762.600 ;
        RECT 850.950 760.950 853.050 766.050 ;
        RECT 857.400 763.050 858.600 800.400 ;
        RECT 871.950 796.950 874.050 801.900 ;
        RECT 878.400 801.000 879.600 802.950 ;
        RECT 877.950 796.950 880.050 801.000 ;
        RECT 880.950 796.950 883.050 799.050 ;
        RECT 874.950 784.950 877.050 787.050 ;
        RECT 856.950 760.950 859.050 763.050 ;
        RECT 859.950 761.100 862.050 763.200 ;
        RECT 865.950 762.000 868.050 766.050 ;
        RECT 845.400 760.050 846.600 760.950 ;
        RECT 860.400 760.050 861.600 761.100 ;
        RECT 866.400 760.050 867.600 762.000 ;
        RECT 844.950 757.950 847.050 760.050 ;
        RECT 847.950 757.950 850.050 760.050 ;
        RECT 853.950 757.950 856.050 760.050 ;
        RECT 859.950 757.950 862.050 760.050 ;
        RECT 862.950 757.950 865.050 760.050 ;
        RECT 865.950 757.950 868.050 760.050 ;
        RECT 868.950 757.950 871.050 760.050 ;
        RECT 848.400 753.600 849.600 757.950 ;
        RECT 850.950 754.950 853.050 757.050 ;
        RECT 845.400 752.400 849.600 753.600 ;
        RECT 835.950 748.950 838.050 751.050 ;
        RECT 832.950 739.950 835.050 742.050 ;
        RECT 845.400 730.200 846.600 752.400 ;
        RECT 847.950 741.600 850.050 742.050 ;
        RECT 851.400 741.600 852.600 754.950 ;
        RECT 847.950 740.400 852.600 741.600 ;
        RECT 847.950 739.950 850.050 740.400 ;
        RECT 838.950 728.100 841.050 730.200 ;
        RECT 844.950 728.100 847.050 730.200 ;
        RECT 848.400 730.050 849.600 739.950 ;
        RECT 850.950 730.950 853.050 733.050 ;
        RECT 839.400 727.050 840.600 728.100 ;
        RECT 845.400 727.050 846.600 728.100 ;
        RECT 847.950 727.950 850.050 730.050 ;
        RECT 835.950 724.950 838.050 727.050 ;
        RECT 838.950 724.950 841.050 727.050 ;
        RECT 841.950 724.950 844.050 727.050 ;
        RECT 844.950 724.950 847.050 727.050 ;
        RECT 832.950 706.950 835.050 709.050 ;
        RECT 833.400 676.050 834.600 706.950 ;
        RECT 836.400 694.050 837.600 724.950 ;
        RECT 842.400 723.000 843.600 724.950 ;
        RECT 841.950 718.950 844.050 723.000 ;
        RECT 835.950 691.950 838.050 694.050 ;
        RECT 841.950 684.000 844.050 688.050 ;
        RECT 847.950 684.000 850.050 688.050 ;
        RECT 851.400 685.050 852.600 730.950 ;
        RECT 842.400 682.050 843.600 684.000 ;
        RECT 848.400 682.050 849.600 684.000 ;
        RECT 850.950 682.950 853.050 685.050 ;
        RECT 838.950 679.950 841.050 682.050 ;
        RECT 841.950 679.950 844.050 682.050 ;
        RECT 844.950 679.950 847.050 682.050 ;
        RECT 847.950 679.950 850.050 682.050 ;
        RECT 839.400 678.900 840.600 679.950 ;
        RECT 838.950 676.800 841.050 678.900 ;
        RECT 832.950 673.950 835.050 676.050 ;
        RECT 841.950 670.950 844.050 673.050 ;
        RECT 842.400 667.050 843.600 670.950 ;
        RECT 845.400 670.050 846.600 679.950 ;
        RECT 850.950 676.950 853.050 679.050 ;
        RECT 844.950 667.950 847.050 670.050 ;
        RECT 829.950 664.950 832.050 667.050 ;
        RECT 841.950 664.950 844.050 667.050 ;
        RECT 832.950 661.950 835.050 664.050 ;
        RECT 833.400 658.050 834.600 661.950 ;
        RECT 851.400 661.050 852.600 676.950 ;
        RECT 854.400 670.050 855.600 757.950 ;
        RECT 863.400 756.000 864.600 757.950 ;
        RECT 869.400 756.900 870.600 757.950 ;
        RECT 856.950 751.950 859.050 754.050 ;
        RECT 862.950 751.950 865.050 756.000 ;
        RECT 868.950 754.800 871.050 756.900 ;
        RECT 857.400 730.050 858.600 751.950 ;
        RECT 865.950 739.950 868.050 742.050 ;
        RECT 859.950 733.950 862.050 736.050 ;
        RECT 856.950 727.950 859.050 730.050 ;
        RECT 860.400 727.050 861.600 733.950 ;
        RECT 866.400 727.050 867.600 739.950 ;
        RECT 875.400 730.050 876.600 784.950 ;
        RECT 877.950 781.950 880.050 784.050 ;
        RECT 874.950 727.950 877.050 730.050 ;
        RECT 859.950 724.950 862.050 727.050 ;
        RECT 862.950 724.950 865.050 727.050 ;
        RECT 865.950 724.950 868.050 727.050 ;
        RECT 868.950 724.950 871.050 727.050 ;
        RECT 856.950 721.950 859.050 724.050 ;
        RECT 857.400 688.050 858.600 721.950 ;
        RECT 859.950 718.950 862.050 721.050 ;
        RECT 860.400 688.050 861.600 718.950 ;
        RECT 863.400 718.050 864.600 724.950 ;
        RECT 869.400 723.900 870.600 724.950 ;
        RECT 868.950 721.800 871.050 723.900 ;
        RECT 871.950 721.950 874.050 724.050 ;
        RECT 862.950 715.950 865.050 718.050 ;
        RECT 856.950 685.950 859.050 688.050 ;
        RECT 859.950 685.950 862.050 688.050 ;
        RECT 860.400 682.050 861.600 685.950 ;
        RECT 865.950 683.100 868.050 688.050 ;
        RECT 872.400 685.050 873.600 721.950 ;
        RECT 866.400 682.050 867.600 683.100 ;
        RECT 871.950 682.950 874.050 685.050 ;
        RECT 874.950 683.100 877.050 685.200 ;
        RECT 859.950 679.950 862.050 682.050 ;
        RECT 862.950 679.950 865.050 682.050 ;
        RECT 865.950 679.950 868.050 682.050 ;
        RECT 868.950 679.950 871.050 682.050 ;
        RECT 859.950 673.950 862.050 676.050 ;
        RECT 853.950 667.950 856.050 670.050 ;
        RECT 843.000 660.600 847.050 661.050 ;
        RECT 842.400 658.950 847.050 660.600 ;
        RECT 850.950 658.950 853.050 661.050 ;
        RECT 832.950 655.950 835.050 658.050 ;
        RECT 829.950 649.950 832.050 655.050 ;
        RECT 835.950 650.100 838.050 652.200 ;
        RECT 836.400 649.050 837.600 650.100 ;
        RECT 842.400 649.050 843.600 658.950 ;
        RECT 832.950 646.950 835.050 649.050 ;
        RECT 835.950 646.950 838.050 649.050 ;
        RECT 838.950 646.950 841.050 649.050 ;
        RECT 841.950 646.950 844.050 649.050 ;
        RECT 829.950 643.950 832.050 646.050 ;
        RECT 814.950 637.950 817.050 640.050 ;
        RECT 823.950 637.950 826.050 640.050 ;
        RECT 805.950 631.950 808.050 634.050 ;
        RECT 805.950 616.950 808.050 619.050 ;
        RECT 790.950 604.800 793.050 606.900 ;
        RECT 793.950 604.950 796.050 607.050 ;
        RECT 802.950 606.600 805.050 607.050 ;
        RECT 800.400 605.400 805.050 606.600 ;
        RECT 784.950 592.950 787.050 595.050 ;
        RECT 787.950 592.950 790.050 595.050 ;
        RECT 778.950 589.950 781.050 592.050 ;
        RECT 784.950 583.950 787.050 586.050 ;
        RECT 781.950 580.950 784.050 583.050 ;
        RECT 775.950 574.950 778.050 577.050 ;
        RECT 776.400 571.050 777.600 574.950 ;
        RECT 782.400 574.050 783.600 580.950 ;
        RECT 785.400 577.050 786.600 583.950 ;
        RECT 791.400 580.050 792.600 604.800 ;
        RECT 800.400 604.050 801.600 605.400 ;
        RECT 802.950 604.950 805.050 605.400 ;
        RECT 796.950 601.950 799.050 604.050 ;
        RECT 799.950 601.950 802.050 604.050 ;
        RECT 797.400 600.900 798.600 601.950 ;
        RECT 796.950 598.800 799.050 600.900 ;
        RECT 802.950 598.950 805.050 601.050 ;
        RECT 796.950 592.950 799.050 595.050 ;
        RECT 790.950 577.950 793.050 580.050 ;
        RECT 797.400 577.050 798.600 592.950 ;
        RECT 799.950 577.950 802.050 580.050 ;
        RECT 784.950 574.950 787.050 577.050 ;
        RECT 796.950 574.950 799.050 577.050 ;
        RECT 781.950 571.950 784.050 574.050 ;
        RECT 787.950 572.100 790.050 574.200 ;
        RECT 793.950 572.100 796.050 574.200 ;
        RECT 800.400 574.050 801.600 577.950 ;
        RECT 803.400 577.050 804.600 598.950 ;
        RECT 806.400 586.050 807.600 616.950 ;
        RECT 811.950 613.950 814.050 616.050 ;
        RECT 808.950 604.950 811.050 607.050 ;
        RECT 805.950 583.950 808.050 586.050 ;
        RECT 802.950 574.950 805.050 577.050 ;
        RECT 788.400 571.050 789.600 572.100 ;
        RECT 794.400 571.050 795.600 572.100 ;
        RECT 799.950 571.950 802.050 574.050 ;
        RECT 805.950 573.600 808.050 577.050 ;
        RECT 809.400 574.050 810.600 604.950 ;
        RECT 812.400 598.050 813.600 613.950 ;
        RECT 815.400 607.050 816.600 637.950 ;
        RECT 817.950 616.950 820.050 619.050 ;
        RECT 814.950 604.950 817.050 607.050 ;
        RECT 818.400 604.050 819.600 616.950 ;
        RECT 823.950 606.000 826.050 610.050 ;
        RECT 830.400 606.600 831.600 643.950 ;
        RECT 833.400 640.050 834.600 646.950 ;
        RECT 835.950 640.950 838.050 643.050 ;
        RECT 832.950 637.950 835.050 640.050 ;
        RECT 836.400 607.050 837.600 640.950 ;
        RECT 839.400 607.200 840.600 646.950 ;
        RECT 844.950 637.950 847.050 640.050 ;
        RECT 845.400 607.200 846.600 637.950 ;
        RECT 824.400 604.050 825.600 606.000 ;
        RECT 830.400 605.400 834.600 606.600 ;
        RECT 817.950 601.950 820.050 604.050 ;
        RECT 820.950 601.950 823.050 604.050 ;
        RECT 823.950 601.950 826.050 604.050 ;
        RECT 826.950 601.950 829.050 604.050 ;
        RECT 811.950 595.950 814.050 598.050 ;
        RECT 821.400 592.050 822.600 601.950 ;
        RECT 827.400 600.900 828.600 601.950 ;
        RECT 826.950 598.800 829.050 600.900 ;
        RECT 829.950 598.950 832.050 601.050 ;
        RECT 830.400 592.050 831.600 598.950 ;
        RECT 820.950 589.950 823.050 592.050 ;
        RECT 826.800 591.000 828.900 592.050 ;
        RECT 826.800 589.950 829.050 591.000 ;
        RECT 829.950 589.950 832.050 592.050 ;
        RECT 826.950 588.600 829.050 589.950 ;
        RECT 833.400 589.050 834.600 605.400 ;
        RECT 835.950 604.950 838.050 607.050 ;
        RECT 838.950 605.100 841.050 607.200 ;
        RECT 844.950 605.100 847.050 607.200 ;
        RECT 851.400 607.050 852.600 658.950 ;
        RECT 839.400 604.050 840.600 605.100 ;
        RECT 845.400 604.050 846.600 605.100 ;
        RECT 850.950 604.950 853.050 607.050 ;
        RECT 838.950 601.950 841.050 604.050 ;
        RECT 841.950 601.950 844.050 604.050 ;
        RECT 844.950 601.950 847.050 604.050 ;
        RECT 847.950 601.950 850.050 604.050 ;
        RECT 835.950 598.950 838.050 601.050 ;
        RECT 826.950 588.000 831.600 588.600 ;
        RECT 827.400 587.400 831.600 588.000 ;
        RECT 826.950 583.950 829.050 586.050 ;
        RECT 817.950 580.950 820.050 583.050 ;
        RECT 803.400 573.000 808.050 573.600 ;
        RECT 803.400 572.400 807.600 573.000 ;
        RECT 775.950 568.950 778.050 571.050 ;
        RECT 784.950 568.950 787.050 571.050 ;
        RECT 787.950 568.950 790.050 571.050 ;
        RECT 790.950 568.950 793.050 571.050 ;
        RECT 793.950 568.950 796.050 571.050 ;
        RECT 796.950 568.950 799.050 571.050 ;
        RECT 785.400 568.050 786.600 568.950 ;
        RECT 781.950 566.400 786.600 568.050 ;
        RECT 791.400 567.900 792.600 568.950 ;
        RECT 797.400 568.050 798.600 568.950 ;
        RECT 781.950 565.950 786.000 566.400 ;
        RECT 790.950 565.800 793.050 567.900 ;
        RECT 797.400 566.400 802.050 568.050 ;
        RECT 798.000 565.950 802.050 566.400 ;
        RECT 781.950 562.800 784.050 564.900 ;
        RECT 787.950 562.950 790.050 565.050 ;
        RECT 775.950 556.950 778.050 559.050 ;
        RECT 776.400 552.600 777.600 556.950 ;
        RECT 776.400 551.400 780.600 552.600 ;
        RECT 772.950 544.950 775.050 547.050 ;
        RECT 772.950 538.950 775.050 541.050 ;
        RECT 766.950 535.950 769.050 538.050 ;
        RECT 766.950 527.100 769.050 529.200 ;
        RECT 767.400 505.050 768.600 527.100 ;
        RECT 773.400 526.050 774.600 538.950 ;
        RECT 779.400 529.050 780.600 551.400 ;
        RECT 782.400 547.050 783.600 562.800 ;
        RECT 784.950 559.950 787.050 562.050 ;
        RECT 781.950 544.950 784.050 547.050 ;
        RECT 779.400 526.950 784.050 529.050 ;
        RECT 779.400 526.050 780.600 526.950 ;
        RECT 772.950 523.950 775.050 526.050 ;
        RECT 775.950 523.950 778.050 526.050 ;
        RECT 778.950 523.950 781.050 526.050 ;
        RECT 776.400 522.900 777.600 523.950 ;
        RECT 785.400 523.050 786.600 559.950 ;
        RECT 788.400 553.050 789.600 562.950 ;
        RECT 803.400 559.050 804.600 572.400 ;
        RECT 808.950 571.950 811.050 574.050 ;
        RECT 818.400 571.050 819.600 580.950 ;
        RECT 823.950 577.950 826.050 580.050 ;
        RECT 824.400 571.050 825.600 577.950 ;
        RECT 827.400 574.050 828.600 583.950 ;
        RECT 830.400 583.050 831.600 587.400 ;
        RECT 832.950 586.950 835.050 589.050 ;
        RECT 829.950 580.950 832.050 583.050 ;
        RECT 829.950 579.600 832.050 579.900 ;
        RECT 829.950 578.400 834.600 579.600 ;
        RECT 829.950 577.800 832.050 578.400 ;
        RECT 826.950 571.950 829.050 574.050 ;
        RECT 808.950 568.800 811.050 570.900 ;
        RECT 814.950 568.950 817.050 571.050 ;
        RECT 817.950 568.950 820.050 571.050 ;
        RECT 820.950 568.950 823.050 571.050 ;
        RECT 823.950 568.950 826.050 571.050 ;
        RECT 805.950 562.950 808.050 565.050 ;
        RECT 802.950 556.950 805.050 559.050 ;
        RECT 787.950 550.950 790.050 553.050 ;
        RECT 790.950 541.950 793.050 544.050 ;
        RECT 787.950 538.950 790.050 541.050 ;
        RECT 775.950 520.800 778.050 522.900 ;
        RECT 781.950 520.950 784.050 523.050 ;
        RECT 784.950 520.950 787.050 523.050 ;
        RECT 778.950 514.950 781.050 517.050 ;
        RECT 775.950 511.950 778.050 514.050 ;
        RECT 769.950 508.950 772.050 511.050 ;
        RECT 766.950 502.950 769.050 505.050 ;
        RECT 763.950 499.950 766.050 502.050 ;
        RECT 770.400 496.050 771.600 508.950 ;
        RECT 772.950 496.950 775.050 499.050 ;
        RECT 769.950 493.950 772.050 496.050 ;
        RECT 757.950 490.950 760.050 493.050 ;
        RECT 760.950 490.950 763.050 493.050 ;
        RECT 766.950 490.950 769.050 493.050 ;
        RECT 754.950 487.950 757.050 490.050 ;
        RECT 755.400 475.050 756.600 487.950 ;
        RECT 758.400 484.050 759.600 490.950 ;
        RECT 767.400 489.600 768.600 490.950 ;
        RECT 764.400 488.400 768.600 489.600 ;
        RECT 764.400 484.050 765.600 488.400 ;
        RECT 766.950 484.950 772.050 487.050 ;
        RECT 773.400 484.050 774.600 496.950 ;
        RECT 776.400 496.050 777.600 511.950 ;
        RECT 779.400 498.600 780.600 514.950 ;
        RECT 782.400 514.050 783.600 520.950 ;
        RECT 781.950 511.950 784.050 514.050 ;
        RECT 779.400 497.400 783.600 498.600 ;
        RECT 775.950 493.950 778.050 496.050 ;
        RECT 782.400 493.050 783.600 497.400 ;
        RECT 788.400 493.050 789.600 538.950 ;
        RECT 791.400 538.050 792.600 541.950 ;
        RECT 790.950 535.950 793.050 538.050 ;
        RECT 793.950 532.950 796.050 535.050 ;
        RECT 794.400 529.200 795.600 532.950 ;
        RECT 793.950 527.100 796.050 529.200 ;
        RECT 799.950 527.100 802.050 529.200 ;
        RECT 794.400 526.050 795.600 527.100 ;
        RECT 800.400 526.050 801.600 527.100 ;
        RECT 793.950 523.950 796.050 526.050 ;
        RECT 796.950 523.950 799.050 526.050 ;
        RECT 799.950 523.950 802.050 526.050 ;
        RECT 790.950 520.800 793.050 522.900 ;
        RECT 791.400 499.050 792.600 520.800 ;
        RECT 797.400 520.050 798.600 523.950 ;
        RECT 802.950 520.950 805.050 523.050 ;
        RECT 797.400 518.400 802.050 520.050 ;
        RECT 798.000 517.950 802.050 518.400 ;
        RECT 803.400 511.050 804.600 520.950 ;
        RECT 802.950 508.950 805.050 511.050 ;
        RECT 806.400 508.050 807.600 562.950 ;
        RECT 809.400 553.050 810.600 568.800 ;
        RECT 815.400 567.900 816.600 568.950 ;
        RECT 814.950 565.800 817.050 567.900 ;
        RECT 821.400 567.000 822.600 568.950 ;
        RECT 820.950 562.950 823.050 567.000 ;
        RECT 830.400 564.600 831.600 577.800 ;
        RECT 833.400 573.600 834.600 578.400 ;
        RECT 836.400 577.050 837.600 598.950 ;
        RECT 842.400 597.600 843.600 601.950 ;
        RECT 848.400 600.900 849.600 601.950 ;
        RECT 854.400 601.050 855.600 667.950 ;
        RECT 856.950 661.950 859.050 664.050 ;
        RECT 857.400 658.050 858.600 661.950 ;
        RECT 856.950 655.950 859.050 658.050 ;
        RECT 860.400 649.050 861.600 673.950 ;
        RECT 863.400 670.050 864.600 679.950 ;
        RECT 862.950 667.950 865.050 670.050 ;
        RECT 869.400 667.050 870.600 679.950 ;
        RECT 871.950 676.950 874.050 679.050 ;
        RECT 868.950 664.950 871.050 667.050 ;
        RECT 865.950 650.100 868.050 652.200 ;
        RECT 872.400 652.050 873.600 676.950 ;
        RECT 875.400 676.050 876.600 683.100 ;
        RECT 874.950 673.950 877.050 676.050 ;
        RECT 878.400 667.050 879.600 781.950 ;
        RECT 881.400 685.050 882.600 796.950 ;
        RECT 884.400 784.050 885.600 806.100 ;
        RECT 883.950 781.950 886.050 784.050 ;
        RECT 887.400 709.050 888.600 841.950 ;
        RECT 892.950 838.950 895.050 841.050 ;
        RECT 889.950 811.950 892.050 814.050 ;
        RECT 890.400 724.050 891.600 811.950 ;
        RECT 893.400 757.050 894.600 838.950 ;
        RECT 895.950 823.950 898.050 826.050 ;
        RECT 892.950 754.950 895.050 757.050 ;
        RECT 896.400 733.050 897.600 823.950 ;
        RECT 895.950 730.950 898.050 733.050 ;
        RECT 889.950 721.950 892.050 724.050 ;
        RECT 886.950 706.950 889.050 709.050 ;
        RECT 880.950 682.950 883.050 685.050 ;
        RECT 883.950 679.950 886.050 682.050 ;
        RECT 880.950 673.950 883.050 679.050 ;
        RECT 877.950 664.950 880.050 667.050 ;
        RECT 884.400 664.050 885.600 679.950 ;
        RECT 892.950 676.950 895.050 679.050 ;
        RECT 889.950 673.950 892.050 676.050 ;
        RECT 883.950 661.950 886.050 664.050 ;
        RECT 866.400 649.050 867.600 650.100 ;
        RECT 871.950 649.950 874.050 652.050 ;
        RECT 874.950 650.100 877.050 652.200 ;
        RECT 883.950 650.100 886.050 652.200 ;
        RECT 859.950 646.950 862.050 649.050 ;
        RECT 862.950 646.950 865.050 649.050 ;
        RECT 865.950 646.950 868.050 649.050 ;
        RECT 868.950 646.950 871.050 649.050 ;
        RECT 863.400 643.050 864.600 646.950 ;
        RECT 862.950 640.950 865.050 643.050 ;
        RECT 859.950 613.950 862.050 616.050 ;
        RECT 856.950 604.950 859.050 607.050 ;
        RECT 847.950 598.800 850.050 600.900 ;
        RECT 853.950 598.950 856.050 601.050 ;
        RECT 842.400 596.400 846.600 597.600 ;
        RECT 841.950 592.950 844.050 595.050 ;
        RECT 838.950 586.950 841.050 589.050 ;
        RECT 839.400 580.050 840.600 586.950 ;
        RECT 838.950 577.950 841.050 580.050 ;
        RECT 835.950 574.950 838.050 577.050 ;
        RECT 833.400 572.400 837.600 573.600 ;
        RECT 836.400 571.050 837.600 572.400 ;
        RECT 842.400 571.050 843.600 592.950 ;
        RECT 845.400 592.050 846.600 596.400 ;
        RECT 853.950 595.800 856.050 597.900 ;
        RECT 844.950 589.950 847.050 592.050 ;
        RECT 845.400 577.050 846.600 589.950 ;
        RECT 850.950 577.950 853.050 580.050 ;
        RECT 844.950 574.950 847.050 577.050 ;
        RECT 835.950 568.950 838.050 571.050 ;
        RECT 838.950 568.950 841.050 571.050 ;
        RECT 841.950 568.950 844.050 571.050 ;
        RECT 844.950 568.950 847.050 571.050 ;
        RECT 832.950 565.950 835.050 568.050 ;
        RECT 839.400 567.000 840.600 568.950 ;
        RECT 827.400 563.400 831.600 564.600 ;
        RECT 811.950 556.950 814.050 559.050 ;
        RECT 808.950 550.950 811.050 553.050 ;
        RECT 808.950 544.950 811.050 547.050 ;
        RECT 809.400 529.050 810.600 544.950 ;
        RECT 812.400 544.050 813.600 556.950 ;
        RECT 820.950 544.950 823.050 547.050 ;
        RECT 811.950 541.950 814.050 544.050 ;
        RECT 811.950 532.950 814.050 535.050 ;
        RECT 808.950 526.950 811.050 529.050 ;
        RECT 812.400 526.050 813.600 532.950 ;
        RECT 821.400 526.050 822.600 544.950 ;
        RECT 823.950 538.950 826.050 541.050 ;
        RECT 824.400 529.050 825.600 538.950 ;
        RECT 823.950 526.950 826.050 529.050 ;
        RECT 811.950 523.950 814.050 526.050 ;
        RECT 817.950 523.950 820.050 526.050 ;
        RECT 820.950 523.950 823.050 526.050 ;
        RECT 808.950 517.950 811.050 523.050 ;
        RECT 814.950 520.950 817.050 523.050 ;
        RECT 799.950 505.950 802.050 508.050 ;
        RECT 805.950 505.950 808.050 508.050 ;
        RECT 796.950 499.950 799.050 502.050 ;
        RECT 790.950 496.950 793.050 499.050 ;
        RECT 778.950 490.950 781.050 493.050 ;
        RECT 781.950 490.950 784.050 493.050 ;
        RECT 784.950 490.950 787.050 493.050 ;
        RECT 787.950 490.950 790.050 493.050 ;
        RECT 790.950 490.950 793.050 493.050 ;
        RECT 779.400 490.050 780.600 490.950 ;
        RECT 775.950 488.400 780.600 490.050 ;
        RECT 785.400 489.900 786.600 490.950 ;
        RECT 775.950 487.950 780.000 488.400 ;
        RECT 784.950 487.800 787.050 489.900 ;
        RECT 775.950 484.800 778.050 486.900 ;
        RECT 781.950 484.950 784.050 487.050 ;
        RECT 787.950 484.950 790.050 487.050 ;
        RECT 757.950 481.950 760.050 484.050 ;
        RECT 763.950 481.950 766.050 484.050 ;
        RECT 754.950 472.950 757.050 475.050 ;
        RECT 748.950 463.950 751.050 466.050 ;
        RECT 758.400 460.050 759.600 481.950 ;
        RECT 766.950 481.800 769.050 483.900 ;
        RECT 772.950 481.950 775.050 484.050 ;
        RECT 763.950 472.950 766.050 475.050 ;
        RECT 757.950 457.950 760.050 460.050 ;
        RECT 757.950 449.100 760.050 451.200 ;
        RECT 758.400 448.050 759.600 449.100 ;
        RECT 754.950 445.950 757.050 448.050 ;
        RECT 757.950 445.950 760.050 448.050 ;
        RECT 755.400 444.900 756.600 445.950 ;
        RECT 754.950 442.800 757.050 444.900 ;
        RECT 760.950 430.950 763.050 433.050 ;
        RECT 764.400 432.600 765.600 472.950 ;
        RECT 767.400 442.050 768.600 481.800 ;
        RECT 776.400 478.050 777.600 484.800 ;
        RECT 778.950 481.950 781.050 484.050 ;
        RECT 775.950 475.950 778.050 478.050 ;
        RECT 779.400 475.050 780.600 481.950 ;
        RECT 782.400 478.050 783.600 484.950 ;
        RECT 784.950 478.950 787.050 481.050 ;
        RECT 781.950 475.950 784.050 478.050 ;
        RECT 772.950 472.950 775.050 475.050 ;
        RECT 778.950 472.950 781.050 475.050 ;
        RECT 773.400 448.050 774.600 472.950 ;
        RECT 779.400 463.050 780.600 472.950 ;
        RECT 781.950 463.950 784.050 466.050 ;
        RECT 778.950 460.950 781.050 463.050 ;
        RECT 779.400 448.050 780.600 460.950 ;
        RECT 782.400 451.050 783.600 463.950 ;
        RECT 781.950 448.950 784.050 451.050 ;
        RECT 772.950 445.950 775.050 448.050 ;
        RECT 775.950 445.950 778.050 448.050 ;
        RECT 778.950 445.950 781.050 448.050 ;
        RECT 769.950 442.950 772.050 445.050 ;
        RECT 776.400 444.000 777.600 445.950 ;
        RECT 766.950 439.950 769.050 442.050 ;
        RECT 764.400 431.400 768.600 432.600 ;
        RECT 739.950 427.950 742.050 430.050 ;
        RECT 745.950 427.950 748.050 430.050 ;
        RECT 751.950 421.950 754.050 424.050 ;
        RECT 739.950 418.950 742.050 421.050 ;
        RECT 721.950 415.950 724.050 418.050 ;
        RECT 736.950 415.950 739.050 418.050 ;
        RECT 724.950 412.950 727.050 415.050 ;
        RECT 733.950 412.950 736.050 415.050 ;
        RECT 718.950 409.800 721.050 411.900 ;
        RECT 715.950 406.950 718.050 409.050 ;
        RECT 712.950 394.950 715.050 397.050 ;
        RECT 706.950 383.400 711.600 384.600 ;
        RECT 706.950 382.950 709.050 383.400 ;
        RECT 692.100 376.200 694.200 378.300 ;
        RECT 701.100 376.500 703.200 378.600 ;
        RECT 689.400 369.900 690.600 372.450 ;
        RECT 689.400 367.800 691.500 369.900 ;
        RECT 692.400 363.600 693.300 376.200 ;
        RECT 698.400 372.900 699.600 375.450 ;
        RECT 698.400 370.800 700.500 372.900 ;
        RECT 694.200 369.900 696.300 370.200 ;
        RECT 702.150 369.900 703.050 376.500 ;
        RECT 707.400 373.050 708.600 382.950 ;
        RECT 706.950 370.950 709.050 373.050 ;
        RECT 709.950 371.100 712.050 373.200 ;
        RECT 694.200 369.000 703.050 369.900 ;
        RECT 694.200 368.100 696.300 369.000 ;
        RECT 699.150 367.200 701.250 368.100 ;
        RECT 694.200 366.000 701.250 367.200 ;
        RECT 694.200 365.100 696.300 366.000 ;
        RECT 691.650 361.500 693.750 363.600 ;
        RECT 698.400 362.100 700.500 364.200 ;
        RECT 702.150 363.900 703.050 369.000 ;
        RECT 703.950 367.800 706.050 369.900 ;
        RECT 704.400 365.400 705.600 367.800 ;
        RECT 710.400 364.050 711.600 371.100 ;
        RECT 698.400 360.000 699.600 362.100 ;
        RECT 701.700 361.800 703.800 363.900 ;
        RECT 709.950 361.950 712.050 364.050 ;
        RECT 697.950 355.950 700.050 360.000 ;
        RECT 683.400 353.400 687.600 354.600 ;
        RECT 658.950 337.950 661.050 340.050 ;
        RECT 670.950 338.100 673.050 340.200 ;
        RECT 676.950 339.000 679.050 343.050 ;
        RECT 671.400 337.050 672.600 338.100 ;
        RECT 677.400 337.050 678.600 339.000 ;
        RECT 682.950 337.950 685.050 340.050 ;
        RECT 646.950 334.950 649.050 337.050 ;
        RECT 649.950 334.950 652.050 337.050 ;
        RECT 652.950 334.950 655.050 337.050 ;
        RECT 655.950 334.950 658.050 337.050 ;
        RECT 661.950 334.950 664.050 337.050 ;
        RECT 667.950 334.950 670.050 337.050 ;
        RECT 670.950 334.950 673.050 337.050 ;
        RECT 673.950 334.950 676.050 337.050 ;
        RECT 676.950 334.950 679.050 337.050 ;
        RECT 641.400 332.400 645.600 333.600 ;
        RECT 619.950 313.950 622.050 316.050 ;
        RECT 637.950 313.950 640.050 316.050 ;
        RECT 613.950 283.950 616.050 286.050 ;
        RECT 616.950 283.950 619.050 286.050 ;
        RECT 616.950 274.950 619.050 277.050 ;
        RECT 598.950 271.950 601.050 274.050 ;
        RECT 556.950 268.950 559.050 271.050 ;
        RECT 580.950 268.950 583.050 271.050 ;
        RECT 589.950 268.950 592.050 271.050 ;
        RECT 595.950 268.950 598.050 271.050 ;
        RECT 547.950 265.950 550.050 268.050 ;
        RECT 553.950 265.950 556.050 268.050 ;
        RECT 524.400 260.400 528.600 261.600 ;
        RECT 505.950 256.950 508.050 259.050 ;
        RECT 508.950 256.950 511.050 259.050 ;
        RECT 511.950 256.950 514.050 259.050 ;
        RECT 514.950 256.950 517.050 259.050 ;
        RECT 509.400 253.050 510.600 256.950 ;
        RECT 515.400 255.900 516.600 256.950 ;
        RECT 521.400 255.900 522.600 259.950 ;
        RECT 514.950 253.800 517.050 255.900 ;
        RECT 520.950 253.800 523.050 255.900 ;
        RECT 508.950 250.950 511.050 253.050 ;
        RECT 499.950 235.950 502.050 238.050 ;
        RECT 509.400 235.050 510.600 250.950 ;
        RECT 517.950 238.950 520.050 241.050 ;
        RECT 508.950 232.950 511.050 235.050 ;
        RECT 487.950 223.950 490.050 226.050 ;
        RECT 481.950 222.600 484.050 223.050 ;
        RECT 481.950 221.400 486.600 222.600 ;
        RECT 481.950 220.950 484.050 221.400 ;
        RECT 478.950 215.100 481.050 217.200 ;
        RECT 479.400 214.050 480.600 215.100 ;
        RECT 475.950 211.950 478.050 214.050 ;
        RECT 478.950 211.950 481.050 214.050 ;
        RECT 476.400 210.900 477.600 211.950 ;
        RECT 485.400 211.050 486.600 221.400 ;
        RECT 475.950 208.800 478.050 210.900 ;
        RECT 484.950 208.950 487.050 211.050 ;
        RECT 476.400 199.050 477.600 208.800 ;
        RECT 481.950 207.900 486.000 208.050 ;
        RECT 481.950 205.950 487.050 207.900 ;
        RECT 484.950 205.800 487.050 205.950 ;
        RECT 488.400 202.050 489.600 223.950 ;
        RECT 496.950 215.100 499.050 217.200 ;
        RECT 504.000 216.600 508.050 217.050 ;
        RECT 497.400 214.050 498.600 215.100 ;
        RECT 503.400 214.950 508.050 216.600 ;
        RECT 503.400 214.050 504.600 214.950 ;
        RECT 493.950 211.950 496.050 214.050 ;
        RECT 496.950 211.950 499.050 214.050 ;
        RECT 499.950 211.950 502.050 214.050 ;
        RECT 502.950 211.950 505.050 214.050 ;
        RECT 494.400 210.900 495.600 211.950 ;
        RECT 493.950 208.800 496.050 210.900 ;
        RECT 490.950 202.950 493.050 208.050 ;
        RECT 500.400 202.050 501.600 211.950 ;
        RECT 505.950 208.950 508.050 211.050 ;
        RECT 506.400 205.050 507.600 208.950 ;
        RECT 505.950 202.950 508.050 205.050 ;
        RECT 509.400 202.050 510.600 232.950 ;
        RECT 518.400 223.050 519.600 238.950 ;
        RECT 517.950 220.950 520.050 223.050 ;
        RECT 511.950 217.950 514.050 220.050 ;
        RECT 487.950 199.950 490.050 202.050 ;
        RECT 499.950 199.950 502.050 202.050 ;
        RECT 508.950 199.950 511.050 202.050 ;
        RECT 475.950 196.950 478.050 199.050 ;
        RECT 469.950 190.950 472.050 193.050 ;
        RECT 484.950 188.400 487.050 190.500 ;
        RECT 505.950 188.400 508.050 190.500 ;
        RECT 476.400 182.400 483.600 183.600 ;
        RECT 476.400 181.050 477.600 182.400 ;
        RECT 482.400 181.050 483.600 182.400 ;
        RECT 472.950 178.950 475.050 181.050 ;
        RECT 475.950 178.950 478.050 181.050 ;
        RECT 481.950 178.950 484.050 181.050 ;
        RECT 473.400 177.900 474.600 178.950 ;
        RECT 472.950 175.800 475.050 177.900 ;
        RECT 466.950 172.950 469.050 175.050 ;
        RECT 473.400 157.050 474.600 175.800 ;
        RECT 475.950 172.950 478.050 175.050 ;
        RECT 485.850 173.400 487.050 188.400 ;
        RECT 499.950 178.950 502.050 181.050 ;
        RECT 472.950 154.950 475.050 157.050 ;
        RECT 463.950 145.950 466.050 148.050 ;
        RECT 469.950 147.300 472.050 149.400 ;
        RECT 451.950 137.100 454.050 139.200 ;
        RECT 457.950 138.000 460.050 142.050 ;
        RECT 464.400 139.050 465.600 145.950 ;
        RECT 470.850 143.700 472.050 147.300 ;
        RECT 469.950 141.600 472.050 143.700 ;
        RECT 452.400 136.050 453.600 137.100 ;
        RECT 458.400 136.050 459.600 138.000 ;
        RECT 463.950 136.950 466.050 139.050 ;
        RECT 451.950 133.950 454.050 136.050 ;
        RECT 454.950 133.950 457.050 136.050 ;
        RECT 457.950 133.950 460.050 136.050 ;
        RECT 460.950 133.950 463.050 136.050 ;
        RECT 466.950 133.950 469.050 136.050 ;
        RECT 455.400 127.050 456.600 133.950 ;
        RECT 454.950 124.950 457.050 127.050 ;
        RECT 461.400 123.600 462.600 133.950 ;
        RECT 467.400 132.600 468.600 133.950 ;
        RECT 466.950 130.500 469.050 132.600 ;
        RECT 470.850 126.600 472.050 141.600 ;
        RECT 476.400 133.050 477.600 172.950 ;
        RECT 484.950 171.300 487.050 173.400 ;
        RECT 485.850 167.700 487.050 171.300 ;
        RECT 484.950 165.600 487.050 167.700 ;
        RECT 490.950 146.400 493.050 148.500 ;
        RECT 500.400 148.050 501.600 178.950 ;
        RECT 506.100 168.600 507.300 188.400 ;
        RECT 512.400 184.050 513.600 217.950 ;
        RECT 518.400 214.050 519.600 220.950 ;
        RECT 524.400 214.050 525.600 260.400 ;
        RECT 532.950 260.100 535.050 262.200 ;
        RECT 533.400 259.050 534.600 260.100 ;
        RECT 529.950 256.950 532.050 259.050 ;
        RECT 532.950 256.950 535.050 259.050 ;
        RECT 535.950 256.950 538.050 259.050 ;
        RECT 530.400 250.050 531.600 256.950 ;
        RECT 536.400 255.000 537.600 256.950 ;
        RECT 535.950 250.950 538.050 255.000 ;
        RECT 529.950 247.950 532.050 250.050 ;
        RECT 548.400 229.050 549.600 265.950 ;
        RECT 556.950 260.100 559.050 262.200 ;
        RECT 557.400 259.050 558.600 260.100 ;
        RECT 565.950 259.950 568.050 262.050 ;
        RECT 553.950 256.950 556.050 259.050 ;
        RECT 556.950 256.950 559.050 259.050 ;
        RECT 559.950 256.950 562.050 259.050 ;
        RECT 554.400 250.050 555.600 256.950 ;
        RECT 553.950 247.950 556.050 250.050 ;
        RECT 560.400 241.050 561.600 256.950 ;
        RECT 559.950 238.950 562.050 241.050 ;
        RECT 547.950 228.600 550.050 229.050 ;
        RECT 545.400 227.400 550.050 228.600 ;
        RECT 535.950 225.300 538.050 227.400 ;
        RECT 536.850 221.700 538.050 225.300 ;
        RECT 535.950 219.600 538.050 221.700 ;
        RECT 517.950 211.950 520.050 214.050 ;
        RECT 520.950 211.950 523.050 214.050 ;
        RECT 523.950 211.950 526.050 214.050 ;
        RECT 532.950 211.950 535.050 214.050 ;
        RECT 514.950 205.950 517.050 211.050 ;
        RECT 521.400 210.000 522.600 211.950 ;
        RECT 533.400 210.600 534.600 211.950 ;
        RECT 520.950 205.950 523.050 210.000 ;
        RECT 532.950 208.500 535.050 210.600 ;
        RECT 536.850 204.600 538.050 219.600 ;
        RECT 535.950 202.500 538.050 204.600 ;
        RECT 514.950 199.950 517.050 202.050 ;
        RECT 511.950 181.950 514.050 184.050 ;
        RECT 508.950 178.950 511.050 181.050 ;
        RECT 509.400 177.600 510.600 178.950 ;
        RECT 508.950 172.950 511.050 177.600 ;
        RECT 505.950 166.500 508.050 168.600 ;
        RECT 511.950 163.950 514.050 166.050 ;
        RECT 502.950 157.950 505.050 160.050 ;
        RECT 478.950 137.400 481.050 139.500 ;
        RECT 484.950 137.400 487.050 139.500 ;
        RECT 475.950 130.950 478.050 133.050 ;
        RECT 479.400 127.050 480.600 137.400 ;
        RECT 485.400 136.050 486.600 137.400 ;
        RECT 484.950 133.950 487.050 136.050 ;
        RECT 469.950 124.500 472.050 126.600 ;
        RECT 478.950 124.950 481.050 127.050 ;
        RECT 491.100 126.600 492.300 146.400 ;
        RECT 499.950 145.950 502.050 148.050 ;
        RECT 493.950 137.400 496.050 139.500 ;
        RECT 499.950 137.400 502.050 139.500 ;
        RECT 494.400 136.050 495.600 137.400 ;
        RECT 493.950 133.950 496.050 136.050 ;
        RECT 490.950 124.500 493.050 126.600 ;
        RECT 461.400 122.400 465.600 123.600 ;
        RECT 457.950 109.950 460.050 112.050 ;
        RECT 451.950 104.100 454.050 106.200 ;
        RECT 452.400 103.050 453.600 104.100 ;
        RECT 458.400 103.050 459.600 109.950 ;
        RECT 451.950 100.950 454.050 103.050 ;
        RECT 454.950 100.950 457.050 103.050 ;
        RECT 457.950 100.950 460.050 103.050 ;
        RECT 455.400 99.900 456.600 100.950 ;
        RECT 464.400 100.050 465.600 122.400 ;
        RECT 475.950 121.950 478.050 124.050 ;
        RECT 476.400 103.050 477.600 121.950 ;
        RECT 500.400 121.050 501.600 137.400 ;
        RECT 487.950 118.950 490.050 121.050 ;
        RECT 499.950 118.950 502.050 121.050 ;
        RECT 481.950 104.100 484.050 106.200 ;
        RECT 482.400 103.050 483.600 104.100 ;
        RECT 472.950 100.950 475.050 103.050 ;
        RECT 475.950 100.950 478.050 103.050 ;
        RECT 478.950 100.950 481.050 103.050 ;
        RECT 481.950 100.950 484.050 103.050 ;
        RECT 454.950 97.800 457.050 99.900 ;
        RECT 463.950 97.950 466.050 100.050 ;
        RECT 473.400 94.050 474.600 100.950 ;
        RECT 472.950 91.950 475.050 94.050 ;
        RECT 479.400 91.050 480.600 100.950 ;
        RECT 478.950 88.950 481.050 91.050 ;
        RECT 445.950 82.950 448.050 85.050 ;
        RECT 454.950 70.950 457.050 73.050 ;
        RECT 442.950 67.950 445.050 70.050 ;
        RECT 436.950 59.100 439.050 61.200 ;
        RECT 437.400 58.050 438.600 59.100 ;
        RECT 445.950 58.950 448.050 61.050 ;
        RECT 436.950 55.950 439.050 58.050 ;
        RECT 446.400 54.900 447.600 58.950 ;
        RECT 455.400 58.050 456.600 70.950 ;
        RECT 472.950 67.950 475.050 70.050 ;
        RECT 469.950 61.950 472.050 64.050 ;
        RECT 460.950 59.100 463.050 61.200 ;
        RECT 461.400 58.050 462.600 59.100 ;
        RECT 451.950 55.950 454.050 58.050 ;
        RECT 454.950 55.950 457.050 58.050 ;
        RECT 457.950 55.950 460.050 58.050 ;
        RECT 460.950 55.950 463.050 58.050 ;
        RECT 452.400 54.900 453.600 55.950 ;
        RECT 445.950 52.800 448.050 54.900 ;
        RECT 451.950 52.800 454.050 54.900 ;
        RECT 451.950 46.950 454.050 49.050 ;
        RECT 427.950 37.950 430.050 40.050 ;
        RECT 430.950 31.950 433.050 34.050 ;
        RECT 424.950 25.950 427.050 28.050 ;
        RECT 431.400 25.050 432.600 31.950 ;
        RECT 442.950 26.400 445.050 28.500 ;
        RECT 427.950 22.950 430.050 25.050 ;
        RECT 430.950 22.950 433.050 25.050 ;
        RECT 433.950 22.950 436.050 25.050 ;
        RECT 428.400 21.900 429.600 22.950 ;
        RECT 434.400 21.900 435.600 22.950 ;
        RECT 443.400 22.050 444.600 26.400 ;
        RECT 452.400 25.050 453.600 46.950 ;
        RECT 458.400 34.050 459.600 55.950 ;
        RECT 463.950 52.950 466.050 55.050 ;
        RECT 464.400 49.050 465.600 52.950 ;
        RECT 463.950 46.950 466.050 49.050 ;
        RECT 470.400 39.600 471.600 61.950 ;
        RECT 473.400 54.900 474.600 67.950 ;
        RECT 479.400 58.050 480.600 88.950 ;
        RECT 488.400 64.050 489.600 118.950 ;
        RECT 490.950 114.600 493.050 115.050 ;
        RECT 496.950 114.600 499.050 115.050 ;
        RECT 490.950 113.400 499.050 114.600 ;
        RECT 490.950 112.950 493.050 113.400 ;
        RECT 496.950 112.950 499.050 113.400 ;
        RECT 493.950 109.950 496.050 112.050 ;
        RECT 494.400 103.050 495.600 109.950 ;
        RECT 493.950 100.950 496.050 103.050 ;
        RECT 496.950 100.950 499.050 103.050 ;
        RECT 497.400 99.900 498.600 100.950 ;
        RECT 496.950 97.800 499.050 99.900 ;
        RECT 503.400 73.050 504.600 157.950 ;
        RECT 508.950 154.950 511.050 157.050 ;
        RECT 509.400 136.050 510.600 154.950 ;
        RECT 512.400 142.050 513.600 163.950 ;
        RECT 515.400 160.050 516.600 199.950 ;
        RECT 523.950 196.950 526.050 199.050 ;
        RECT 538.950 196.950 541.050 199.050 ;
        RECT 517.950 184.950 520.050 187.050 ;
        RECT 518.400 178.050 519.600 184.950 ;
        RECT 524.400 181.050 525.600 196.950 ;
        RECT 535.950 190.950 538.050 193.050 ;
        RECT 529.950 182.100 532.050 184.200 ;
        RECT 530.400 181.050 531.600 182.100 ;
        RECT 523.950 178.950 526.050 181.050 ;
        RECT 526.950 178.950 529.050 181.050 ;
        RECT 529.950 178.950 532.050 181.050 ;
        RECT 517.950 175.950 520.050 178.050 ;
        RECT 527.400 177.900 528.600 178.950 ;
        RECT 526.950 175.800 529.050 177.900 ;
        RECT 514.950 157.950 517.050 160.050 ;
        RECT 536.400 154.050 537.600 190.950 ;
        RECT 539.400 177.900 540.600 196.950 ;
        RECT 545.400 193.050 546.600 227.400 ;
        RECT 547.950 226.950 550.050 227.400 ;
        RECT 556.950 224.400 559.050 226.500 ;
        RECT 550.950 220.950 553.050 223.050 ;
        RECT 551.400 214.050 552.600 220.950 ;
        RECT 550.950 211.950 553.050 214.050 ;
        RECT 557.100 204.600 558.300 224.400 ;
        RECT 559.950 216.000 562.050 220.050 ;
        RECT 560.400 214.050 561.600 216.000 ;
        RECT 559.950 211.950 562.050 214.050 ;
        RECT 556.950 202.500 559.050 204.600 ;
        RECT 566.400 196.050 567.600 259.950 ;
        RECT 581.400 259.050 582.600 268.950 ;
        RECT 574.950 256.950 577.050 259.050 ;
        RECT 580.950 256.950 583.050 259.050 ;
        RECT 583.950 256.950 586.050 259.050 ;
        RECT 575.400 226.050 576.600 256.950 ;
        RECT 584.400 255.900 585.600 256.950 ;
        RECT 583.950 253.800 586.050 255.900 ;
        RECT 583.950 226.950 586.050 229.050 ;
        RECT 574.950 223.950 577.050 226.050 ;
        RECT 571.950 220.950 574.050 223.050 ;
        RECT 568.950 214.950 571.050 217.050 ;
        RECT 569.400 210.600 570.600 214.950 ;
        RECT 572.400 211.050 573.600 220.950 ;
        RECT 577.950 215.100 580.050 217.200 ;
        RECT 578.400 214.050 579.600 215.100 ;
        RECT 584.400 214.050 585.600 226.950 ;
        RECT 590.400 219.600 591.600 268.950 ;
        RECT 592.950 265.950 595.050 268.050 ;
        RECT 593.400 255.900 594.600 265.950 ;
        RECT 610.950 262.950 613.050 265.050 ;
        RECT 601.950 260.100 604.050 262.200 ;
        RECT 602.400 259.050 603.600 260.100 ;
        RECT 598.950 256.950 601.050 259.050 ;
        RECT 601.950 256.950 604.050 259.050 ;
        RECT 604.950 256.950 607.050 259.050 ;
        RECT 599.400 255.900 600.600 256.950 ;
        RECT 592.950 253.800 595.050 255.900 ;
        RECT 598.950 253.800 601.050 255.900 ;
        RECT 605.400 247.050 606.600 256.950 ;
        RECT 604.950 244.950 607.050 247.050 ;
        RECT 595.950 238.950 598.050 241.050 ;
        RECT 590.400 218.400 594.600 219.600 ;
        RECT 589.950 215.100 592.050 217.200 ;
        RECT 577.950 211.950 580.050 214.050 ;
        RECT 580.950 211.950 583.050 214.050 ;
        RECT 583.950 211.950 586.050 214.050 ;
        RECT 568.800 208.500 570.900 210.600 ;
        RECT 571.950 208.950 574.050 211.050 ;
        RECT 581.400 205.050 582.600 211.950 ;
        RECT 590.400 205.050 591.600 215.100 ;
        RECT 580.950 202.950 583.050 205.050 ;
        RECT 589.950 202.950 592.050 205.050 ;
        RECT 565.950 193.950 568.050 196.050 ;
        RECT 577.950 193.950 580.050 196.050 ;
        RECT 544.950 190.950 547.050 193.050 ;
        RECT 574.950 190.950 577.050 193.050 ;
        RECT 547.950 187.950 550.050 190.050 ;
        RECT 562.950 188.400 565.050 190.500 ;
        RECT 548.400 181.050 549.600 187.950 ;
        RECT 544.950 178.950 547.050 181.050 ;
        RECT 547.950 178.950 550.050 181.050 ;
        RECT 550.950 178.950 553.050 181.050 ;
        RECT 559.950 178.950 562.050 181.050 ;
        RECT 545.400 177.900 546.600 178.950 ;
        RECT 551.400 177.900 552.600 178.950 ;
        RECT 538.950 175.800 541.050 177.900 ;
        RECT 544.950 175.800 547.050 177.900 ;
        RECT 550.950 175.800 553.050 177.900 ;
        RECT 560.400 177.000 561.600 178.950 ;
        RECT 559.950 172.950 562.050 177.000 ;
        RECT 563.700 168.600 564.900 188.400 ;
        RECT 568.950 178.950 571.050 181.050 ;
        RECT 569.400 172.050 570.600 178.950 ;
        RECT 568.950 169.950 571.050 172.050 ;
        RECT 562.950 166.500 565.050 168.600 ;
        RECT 575.400 157.050 576.600 190.950 ;
        RECT 578.400 177.900 579.600 193.950 ;
        RECT 583.950 188.400 586.050 190.500 ;
        RECT 577.950 175.800 580.050 177.900 ;
        RECT 583.950 173.400 585.150 188.400 ;
        RECT 586.950 182.400 589.050 184.500 ;
        RECT 587.400 181.050 588.600 182.400 ;
        RECT 586.950 178.950 589.050 181.050 ;
        RECT 583.950 171.300 586.050 173.400 ;
        RECT 583.950 167.700 585.150 171.300 ;
        RECT 583.950 165.600 586.050 167.700 ;
        RECT 574.950 154.950 577.050 157.050 ;
        RECT 526.950 151.950 529.050 154.050 ;
        RECT 535.950 151.950 538.050 154.050 ;
        RECT 514.950 145.950 517.050 148.050 ;
        RECT 511.950 139.950 514.050 142.050 ;
        RECT 515.400 136.050 516.600 145.950 ;
        RECT 520.950 137.100 523.050 139.200 ;
        RECT 521.400 136.050 522.600 137.100 ;
        RECT 508.950 133.950 511.050 136.050 ;
        RECT 511.950 133.950 514.050 136.050 ;
        RECT 514.950 133.950 517.050 136.050 ;
        RECT 517.950 133.950 520.050 136.050 ;
        RECT 520.950 133.950 523.050 136.050 ;
        RECT 505.950 130.950 508.050 133.050 ;
        RECT 512.400 132.900 513.600 133.950 ;
        RECT 506.400 100.050 507.600 130.950 ;
        RECT 511.950 130.800 514.050 132.900 ;
        RECT 518.400 132.000 519.600 133.950 ;
        RECT 517.950 127.950 520.050 132.000 ;
        RECT 520.950 127.950 523.050 130.050 ;
        RECT 514.950 104.100 517.050 106.200 ;
        RECT 515.400 103.050 516.600 104.100 ;
        RECT 521.400 103.050 522.600 127.950 ;
        RECT 523.950 124.950 526.050 130.050 ;
        RECT 514.950 100.950 517.050 103.050 ;
        RECT 517.950 100.950 520.050 103.050 ;
        RECT 520.950 100.950 523.050 103.050 ;
        RECT 505.950 97.950 508.050 100.050 ;
        RECT 511.950 97.950 514.050 100.050 ;
        RECT 502.950 70.950 505.050 73.050 ;
        RECT 505.950 67.950 508.050 70.050 ;
        RECT 487.950 61.950 490.050 64.050 ;
        RECT 499.950 59.100 502.050 61.200 ;
        RECT 500.400 58.050 501.600 59.100 ;
        RECT 506.400 58.050 507.600 67.950 ;
        RECT 478.950 55.950 481.050 58.050 ;
        RECT 481.950 55.950 484.050 58.050 ;
        RECT 496.950 55.950 499.050 58.050 ;
        RECT 499.950 55.950 502.050 58.050 ;
        RECT 502.950 55.950 505.050 58.050 ;
        RECT 505.950 55.950 508.050 58.050 ;
        RECT 482.400 54.900 483.600 55.950 ;
        RECT 472.950 52.800 475.050 54.900 ;
        RECT 481.950 52.800 484.050 54.900 ;
        RECT 497.400 43.050 498.600 55.950 ;
        RECT 503.400 54.900 504.600 55.950 ;
        RECT 502.950 52.800 505.050 54.900 ;
        RECT 496.950 40.950 499.050 43.050 ;
        RECT 470.400 38.400 474.600 39.600 ;
        RECT 457.950 31.950 460.050 34.050 ;
        RECT 466.950 32.400 469.050 34.500 ;
        RECT 463.950 26.400 466.050 28.500 ;
        RECT 464.400 25.050 465.600 26.400 ;
        RECT 448.950 22.950 451.050 25.050 ;
        RECT 451.950 22.950 454.050 25.050 ;
        RECT 454.950 22.950 457.050 25.050 ;
        RECT 463.950 22.950 466.050 25.050 ;
        RECT 389.400 20.400 396.600 21.600 ;
        RECT 397.950 19.800 400.050 21.900 ;
        RECT 406.950 19.800 409.050 21.900 ;
        RECT 412.950 19.800 415.050 21.900 ;
        RECT 418.950 19.800 421.050 21.900 ;
        RECT 427.950 19.800 430.050 21.900 ;
        RECT 433.950 19.800 436.050 21.900 ;
        RECT 442.950 19.950 445.050 22.050 ;
        RECT 449.400 21.900 450.600 22.950 ;
        RECT 448.950 19.800 451.050 21.900 ;
        RECT 455.400 16.050 456.600 22.950 ;
        RECT 467.850 17.400 469.050 32.400 ;
        RECT 473.400 28.050 474.600 38.400 ;
        RECT 475.950 31.950 478.050 34.050 ;
        RECT 487.950 32.400 490.050 34.500 ;
        RECT 472.950 25.950 475.050 28.050 ;
        RECT 476.400 21.600 477.600 31.950 ;
        RECT 481.950 22.950 484.050 25.050 ;
        RECT 482.400 21.600 483.600 22.950 ;
        RECT 475.950 19.500 478.050 21.600 ;
        RECT 481.950 19.500 484.050 21.600 ;
        RECT 454.950 13.950 457.050 16.050 ;
        RECT 466.950 15.300 469.050 17.400 ;
        RECT 313.950 9.600 316.050 11.700 ;
        RECT 364.950 9.600 367.050 11.700 ;
        RECT 385.950 10.500 388.050 12.600 ;
        RECT 455.400 7.050 456.600 13.950 ;
        RECT 467.850 11.700 469.050 15.300 ;
        RECT 488.100 12.600 489.300 32.400 ;
        RECT 512.400 28.050 513.600 97.950 ;
        RECT 514.950 70.950 517.050 73.050 ;
        RECT 511.950 25.950 514.050 28.050 ;
        RECT 490.950 22.950 493.050 25.050 ;
        RECT 508.950 22.950 511.050 25.050 ;
        RECT 491.400 21.600 492.600 22.950 ;
        RECT 509.400 21.900 510.600 22.950 ;
        RECT 490.950 19.500 493.050 21.600 ;
        RECT 508.950 19.800 511.050 21.900 ;
        RECT 515.400 19.050 516.600 70.950 ;
        RECT 518.400 54.900 519.600 100.950 ;
        RECT 527.400 94.050 528.600 151.950 ;
        RECT 575.400 139.200 576.600 154.950 ;
        RECT 538.950 137.100 541.050 139.200 ;
        RECT 547.950 137.100 550.050 139.200 ;
        RECT 553.950 137.100 556.050 139.200 ;
        RECT 562.950 137.100 565.050 139.200 ;
        RECT 568.950 137.100 571.050 139.200 ;
        RECT 574.950 137.100 577.050 139.200 ;
        RECT 539.400 136.050 540.600 137.100 ;
        RECT 548.400 136.050 549.600 137.100 ;
        RECT 538.950 133.950 541.050 136.050 ;
        RECT 544.950 133.950 547.050 136.050 ;
        RECT 547.950 133.950 550.050 136.050 ;
        RECT 545.400 132.000 546.600 133.950 ;
        RECT 544.950 127.950 547.050 132.000 ;
        RECT 541.950 126.600 544.050 127.050 ;
        RECT 547.950 126.600 550.050 130.050 ;
        RECT 541.950 126.000 550.050 126.600 ;
        RECT 541.950 125.400 549.600 126.000 ;
        RECT 541.950 124.950 544.050 125.400 ;
        RECT 532.950 104.100 535.050 106.200 ;
        RECT 538.950 104.100 541.050 106.200 ;
        RECT 554.400 106.050 555.600 137.100 ;
        RECT 563.400 136.050 564.600 137.100 ;
        RECT 569.400 136.050 570.600 137.100 ;
        RECT 580.950 136.950 583.050 139.050 ;
        RECT 589.950 137.100 592.050 139.200 ;
        RECT 593.400 139.050 594.600 218.400 ;
        RECT 596.400 187.050 597.600 238.950 ;
        RECT 611.400 220.050 612.600 262.950 ;
        RECT 617.400 259.050 618.600 274.950 ;
        RECT 620.400 271.050 621.600 313.950 ;
        RECT 625.950 310.950 628.050 313.050 ;
        RECT 626.400 292.050 627.600 310.950 ;
        RECT 631.950 293.100 634.050 295.200 ;
        RECT 638.400 295.050 639.600 313.950 ;
        RECT 632.400 292.050 633.600 293.100 ;
        RECT 637.950 292.950 640.050 295.050 ;
        RECT 640.950 293.100 643.050 295.200 ;
        RECT 625.950 289.950 628.050 292.050 ;
        RECT 628.950 289.950 631.050 292.050 ;
        RECT 631.950 289.950 634.050 292.050 ;
        RECT 634.950 289.950 637.050 292.050 ;
        RECT 629.400 288.000 630.600 289.950 ;
        RECT 628.950 283.950 631.050 288.000 ;
        RECT 619.950 268.950 622.050 271.050 ;
        RECT 631.950 268.950 634.050 271.050 ;
        RECT 622.950 261.000 625.050 265.050 ;
        RECT 623.400 259.050 624.600 261.000 ;
        RECT 616.950 256.950 619.050 259.050 ;
        RECT 619.950 256.950 622.050 259.050 ;
        RECT 622.950 256.950 625.050 259.050 ;
        RECT 625.950 256.950 628.050 259.050 ;
        RECT 620.400 250.050 621.600 256.950 ;
        RECT 626.400 255.900 627.600 256.950 ;
        RECT 632.400 256.050 633.600 268.950 ;
        RECT 625.950 253.800 628.050 255.900 ;
        RECT 631.950 253.950 634.050 256.050 ;
        RECT 619.950 247.950 622.050 250.050 ;
        RECT 632.400 247.050 633.600 253.950 ;
        RECT 631.950 244.950 634.050 247.050 ;
        RECT 622.950 223.950 625.050 226.050 ;
        RECT 610.950 217.950 613.050 220.050 ;
        RECT 616.950 217.950 619.050 220.050 ;
        RECT 601.950 215.100 604.050 217.200 ;
        RECT 607.950 215.100 610.050 217.200 ;
        RECT 602.400 214.050 603.600 215.100 ;
        RECT 608.400 214.050 609.600 215.100 ;
        RECT 601.950 211.950 604.050 214.050 ;
        RECT 604.950 211.950 607.050 214.050 ;
        RECT 607.950 211.950 610.050 214.050 ;
        RECT 610.950 211.950 613.050 214.050 ;
        RECT 605.400 210.900 606.600 211.950 ;
        RECT 604.950 208.800 607.050 210.900 ;
        RECT 611.400 199.050 612.600 211.950 ;
        RECT 613.950 208.950 616.050 211.050 ;
        RECT 610.950 196.950 613.050 199.050 ;
        RECT 611.400 193.050 612.600 196.950 ;
        RECT 614.400 196.050 615.600 208.950 ;
        RECT 617.400 208.050 618.600 217.950 ;
        RECT 623.400 214.050 624.600 223.950 ;
        RECT 631.950 215.100 634.050 217.200 ;
        RECT 635.400 216.600 636.600 289.950 ;
        RECT 637.950 286.950 640.050 289.050 ;
        RECT 638.400 256.050 639.600 286.950 ;
        RECT 641.400 277.050 642.600 293.100 ;
        RECT 644.400 280.050 645.600 332.400 ;
        RECT 650.400 325.050 651.600 334.950 ;
        RECT 656.400 331.050 657.600 334.950 ;
        RECT 662.400 331.050 663.600 334.950 ;
        RECT 652.950 328.950 655.050 331.050 ;
        RECT 649.950 322.950 652.050 325.050 ;
        RECT 653.400 310.050 654.600 328.950 ;
        RECT 655.950 325.950 658.050 331.050 ;
        RECT 661.950 328.950 664.050 331.050 ;
        RECT 661.950 325.800 664.050 327.900 ;
        RECT 652.950 307.950 655.050 310.050 ;
        RECT 652.950 301.950 655.050 304.050 ;
        RECT 646.950 292.950 649.050 295.050 ;
        RECT 647.400 288.900 648.600 292.950 ;
        RECT 653.400 292.050 654.600 301.950 ;
        RECT 652.950 289.950 655.050 292.050 ;
        RECT 655.950 289.950 658.050 292.050 ;
        RECT 656.400 288.900 657.600 289.950 ;
        RECT 646.950 286.800 649.050 288.900 ;
        RECT 655.950 286.800 658.050 288.900 ;
        RECT 656.400 283.050 657.600 286.800 ;
        RECT 662.400 286.050 663.600 325.800 ;
        RECT 668.400 325.050 669.600 334.950 ;
        RECT 674.400 333.900 675.600 334.950 ;
        RECT 673.950 331.800 676.050 333.900 ;
        RECT 676.950 325.950 679.050 328.050 ;
        RECT 667.950 322.950 670.050 325.050 ;
        RECT 670.950 293.100 673.050 295.200 ;
        RECT 671.400 292.050 672.600 293.100 ;
        RECT 667.950 289.950 670.050 292.050 ;
        RECT 670.950 289.950 673.050 292.050 ;
        RECT 661.950 283.950 664.050 286.050 ;
        RECT 655.950 280.950 658.050 283.050 ;
        RECT 668.400 280.050 669.600 289.950 ;
        RECT 643.950 277.950 646.050 280.050 ;
        RECT 664.800 277.950 666.900 280.050 ;
        RECT 667.950 277.950 670.050 280.050 ;
        RECT 640.950 274.950 643.050 277.050 ;
        RECT 649.200 263.100 651.300 265.200 ;
        RECT 653.400 264.900 654.600 267.450 ;
        RECT 655.950 265.950 658.050 268.050 ;
        RECT 647.400 259.200 648.600 261.600 ;
        RECT 646.950 257.100 649.050 259.200 ;
        RECT 649.950 258.000 650.850 263.100 ;
        RECT 652.500 262.800 654.600 264.900 ;
        RECT 656.400 261.900 657.600 265.950 ;
        RECT 659.250 263.400 661.350 265.500 ;
        RECT 656.400 261.000 658.800 261.900 ;
        RECT 651.750 259.800 658.800 261.000 ;
        RECT 651.750 258.900 653.850 259.800 ;
        RECT 656.700 258.000 658.800 258.900 ;
        RECT 649.950 257.100 658.800 258.000 ;
        RECT 637.950 253.950 640.050 256.050 ;
        RECT 638.400 250.050 639.600 253.950 ;
        RECT 649.950 250.500 650.850 257.100 ;
        RECT 656.700 256.800 658.800 257.100 ;
        RECT 652.500 254.100 654.600 256.200 ;
        RECT 637.950 247.950 640.050 250.050 ;
        RECT 649.800 248.400 651.900 250.500 ;
        RECT 653.400 232.050 654.600 254.100 ;
        RECT 659.700 250.800 660.600 263.400 ;
        RECT 661.500 257.100 663.600 259.200 ;
        RECT 662.400 254.550 663.600 257.100 ;
        RECT 658.800 248.700 660.900 250.800 ;
        RECT 665.400 235.050 666.600 277.950 ;
        RECT 677.400 277.050 678.600 325.950 ;
        RECT 683.400 294.600 684.600 337.950 ;
        RECT 686.400 313.050 687.600 353.400 ;
        RECT 688.950 352.950 691.050 355.050 ;
        RECT 689.400 333.900 690.600 352.950 ;
        RECT 706.950 343.950 709.050 346.050 ;
        RECT 691.950 339.600 696.000 340.050 ;
        RECT 691.950 337.950 696.600 339.600 ;
        RECT 700.950 338.100 703.050 340.200 ;
        RECT 707.400 340.050 708.600 343.950 ;
        RECT 695.400 337.050 696.600 337.950 ;
        RECT 701.400 337.050 702.600 338.100 ;
        RECT 706.950 337.950 709.050 340.050 ;
        RECT 713.400 339.600 714.600 394.950 ;
        RECT 715.950 385.950 718.050 388.050 ;
        RECT 716.400 346.050 717.600 385.950 ;
        RECT 719.400 379.050 720.600 409.800 ;
        RECT 725.400 406.050 726.600 412.950 ;
        RECT 734.400 411.900 735.600 412.950 ;
        RECT 733.950 409.800 736.050 411.900 ;
        RECT 740.400 409.050 741.600 418.950 ;
        RECT 742.950 415.950 745.050 418.050 ;
        RECT 739.950 406.950 742.050 409.050 ;
        RECT 724.950 403.950 727.050 406.050 ;
        RECT 736.950 400.950 739.050 403.050 ;
        RECT 733.950 394.950 736.050 397.050 ;
        RECT 718.950 376.950 721.050 379.050 ;
        RECT 721.950 371.100 724.050 373.200 ;
        RECT 727.950 371.100 730.050 373.200 ;
        RECT 734.400 373.050 735.600 394.950 ;
        RECT 737.400 382.050 738.600 400.950 ;
        RECT 736.950 379.950 739.050 382.050 ;
        RECT 740.400 373.200 741.600 406.950 ;
        RECT 743.400 376.050 744.600 415.950 ;
        RECT 752.400 415.050 753.600 421.950 ;
        RECT 757.950 417.000 760.050 421.050 ;
        RECT 761.400 418.050 762.600 430.950 ;
        RECT 763.950 427.950 766.050 430.050 ;
        RECT 758.400 415.050 759.600 417.000 ;
        RECT 760.950 415.950 763.050 418.050 ;
        RECT 748.950 412.950 751.050 415.050 ;
        RECT 751.950 412.950 754.050 415.050 ;
        RECT 754.950 412.950 757.050 415.050 ;
        RECT 757.950 412.950 760.050 415.050 ;
        RECT 749.400 412.050 750.600 412.950 ;
        RECT 745.950 410.400 750.600 412.050 ;
        RECT 755.400 411.000 756.600 412.950 ;
        RECT 745.950 409.950 750.000 410.400 ;
        RECT 754.950 406.950 757.050 411.000 ;
        RECT 760.950 409.950 763.050 412.050 ;
        RECT 748.800 391.950 750.900 394.050 ;
        RECT 751.950 391.950 754.050 394.050 ;
        RECT 749.400 376.050 750.600 391.950 ;
        RECT 742.950 373.950 745.050 376.050 ;
        RECT 748.950 373.950 751.050 376.050 ;
        RECT 722.400 370.050 723.600 371.100 ;
        RECT 728.400 370.050 729.600 371.100 ;
        RECT 733.950 370.950 736.050 373.050 ;
        RECT 739.950 372.600 742.050 373.200 ;
        RECT 737.400 371.400 742.050 372.600 ;
        RECT 721.950 367.950 724.050 370.050 ;
        RECT 724.950 367.950 727.050 370.050 ;
        RECT 727.950 367.950 730.050 370.050 ;
        RECT 730.950 367.950 733.050 370.050 ;
        RECT 725.400 349.050 726.600 367.950 ;
        RECT 731.400 366.000 732.600 367.950 ;
        RECT 730.950 361.950 733.050 366.000 ;
        RECT 733.950 364.950 736.050 367.050 ;
        RECT 737.400 366.900 738.600 371.400 ;
        RECT 739.950 371.100 742.050 371.400 ;
        RECT 745.950 371.100 748.050 373.200 ;
        RECT 752.400 373.050 753.600 391.950 ;
        RECT 757.950 373.950 760.050 376.050 ;
        RECT 746.400 370.050 747.600 371.100 ;
        RECT 751.950 370.950 754.050 373.050 ;
        RECT 754.950 370.950 757.050 373.050 ;
        RECT 742.950 367.950 745.050 370.050 ;
        RECT 745.950 367.950 748.050 370.050 ;
        RECT 748.950 367.950 751.050 370.050 ;
        RECT 743.400 366.900 744.600 367.950 ;
        RECT 749.400 367.050 750.600 367.950 ;
        RECT 718.950 346.950 721.050 349.050 ;
        RECT 724.950 346.950 727.050 349.050 ;
        RECT 715.950 343.950 718.050 346.050 ;
        RECT 719.400 340.200 720.600 346.950 ;
        RECT 727.950 343.950 730.050 346.050 ;
        RECT 710.400 338.400 714.600 339.600 ;
        RECT 694.950 334.950 697.050 337.050 ;
        RECT 697.950 334.950 700.050 337.050 ;
        RECT 700.950 334.950 703.050 337.050 ;
        RECT 703.950 334.950 706.050 337.050 ;
        RECT 688.950 331.800 691.050 333.900 ;
        RECT 698.400 325.050 699.600 334.950 ;
        RECT 704.400 333.900 705.600 334.950 ;
        RECT 703.950 331.800 706.050 333.900 ;
        RECT 706.950 331.950 709.050 334.050 ;
        RECT 697.950 322.950 700.050 325.050 ;
        RECT 704.400 316.050 705.600 331.800 ;
        RECT 703.950 313.950 706.050 316.050 ;
        RECT 685.950 310.950 688.050 313.050 ;
        RECT 703.950 295.950 706.050 298.050 ;
        RECT 680.400 293.400 684.600 294.600 ;
        RECT 680.400 288.900 681.600 293.400 ;
        RECT 685.950 293.100 688.050 295.200 ;
        RECT 691.950 293.100 694.050 295.200 ;
        RECT 700.950 293.100 703.050 295.200 ;
        RECT 686.400 292.050 687.600 293.100 ;
        RECT 692.400 292.050 693.600 293.100 ;
        RECT 685.950 289.950 688.050 292.050 ;
        RECT 688.950 289.950 691.050 292.050 ;
        RECT 691.950 289.950 694.050 292.050 ;
        RECT 694.950 289.950 697.050 292.050 ;
        RECT 689.400 288.900 690.600 289.950 ;
        RECT 679.950 286.800 682.050 288.900 ;
        RECT 688.950 286.800 691.050 288.900 ;
        RECT 685.950 283.950 688.050 286.050 ;
        RECT 667.950 274.800 670.050 276.900 ;
        RECT 676.950 274.950 679.050 277.050 ;
        RECT 664.950 232.950 667.050 235.050 ;
        RECT 652.950 229.950 655.050 232.050 ;
        RECT 646.950 223.950 649.050 226.050 ;
        RECT 635.400 215.400 639.600 216.600 ;
        RECT 632.400 214.050 633.600 215.100 ;
        RECT 622.950 211.950 625.050 214.050 ;
        RECT 628.950 211.950 631.050 214.050 ;
        RECT 631.950 211.950 634.050 214.050 ;
        RECT 629.400 210.000 630.600 211.950 ;
        RECT 616.950 205.950 619.050 208.050 ;
        RECT 628.950 205.950 631.050 210.000 ;
        RECT 631.950 202.950 634.050 205.050 ;
        RECT 632.400 199.050 633.600 202.950 ;
        RECT 634.950 199.950 637.050 202.050 ;
        RECT 631.950 196.950 634.050 199.050 ;
        RECT 635.400 196.050 636.600 199.950 ;
        RECT 613.950 193.950 616.050 196.050 ;
        RECT 634.950 193.950 637.050 196.050 ;
        RECT 638.400 193.050 639.600 215.400 ;
        RECT 640.950 214.950 643.050 217.050 ;
        RECT 641.400 202.050 642.600 214.950 ;
        RECT 647.400 214.050 648.600 223.950 ;
        RECT 655.950 215.100 658.050 217.200 ;
        RECT 656.400 214.050 657.600 215.100 ;
        RECT 664.950 214.950 667.050 217.050 ;
        RECT 646.950 211.950 649.050 214.050 ;
        RECT 652.950 211.950 655.050 214.050 ;
        RECT 655.950 211.950 658.050 214.050 ;
        RECT 653.400 210.600 654.600 211.950 ;
        RECT 650.400 209.400 654.600 210.600 ;
        RECT 640.950 199.950 643.050 202.050 ;
        RECT 643.950 196.950 646.050 202.050 ;
        RECT 610.950 190.950 613.050 193.050 ;
        RECT 637.950 190.950 640.050 193.050 ;
        RECT 619.950 187.950 622.050 190.050 ;
        RECT 595.950 184.950 598.050 187.050 ;
        RECT 598.950 182.100 601.050 184.200 ;
        RECT 607.950 182.100 610.050 184.200 ;
        RECT 613.950 183.000 616.050 187.050 ;
        RECT 599.400 163.050 600.600 182.100 ;
        RECT 608.400 181.050 609.600 182.100 ;
        RECT 614.400 181.050 615.600 183.000 ;
        RECT 604.950 178.950 607.050 181.050 ;
        RECT 607.950 178.950 610.050 181.050 ;
        RECT 610.950 178.950 613.050 181.050 ;
        RECT 613.950 178.950 616.050 181.050 ;
        RECT 605.400 177.900 606.600 178.950 ;
        RECT 604.950 175.800 607.050 177.900 ;
        RECT 611.400 174.600 612.600 178.950 ;
        RECT 608.400 173.400 612.600 174.600 ;
        RECT 598.950 160.950 601.050 163.050 ;
        RECT 608.400 139.200 609.600 173.400 ;
        RECT 620.400 172.050 621.600 187.950 ;
        RECT 650.400 187.050 651.600 209.400 ;
        RECT 658.800 202.950 660.900 205.050 ;
        RECT 661.950 202.950 664.050 205.050 ;
        RECT 652.950 187.950 655.050 190.050 ;
        RECT 649.950 184.950 652.050 187.050 ;
        RECT 628.950 182.100 631.050 184.200 ;
        RECT 629.400 181.050 630.600 182.100 ;
        RECT 643.950 181.950 646.050 184.050 ;
        RECT 625.950 178.950 628.050 181.050 ;
        RECT 628.950 178.950 631.050 181.050 ;
        RECT 631.950 178.950 634.050 181.050 ;
        RECT 626.400 177.900 627.600 178.950 ;
        RECT 625.950 175.800 628.050 177.900 ;
        RECT 619.950 169.950 622.050 172.050 ;
        RECT 632.400 157.050 633.600 178.950 ;
        RECT 644.400 175.050 645.600 181.950 ;
        RECT 653.400 181.050 654.600 187.950 ;
        RECT 659.400 187.050 660.600 202.950 ;
        RECT 658.950 184.950 661.050 187.050 ;
        RECT 659.400 181.050 660.600 184.950 ;
        RECT 662.400 183.600 663.600 202.950 ;
        RECT 665.400 196.050 666.600 214.950 ;
        RECT 664.950 193.950 667.050 196.050 ;
        RECT 662.400 182.400 666.600 183.600 ;
        RECT 649.950 178.950 652.050 181.050 ;
        RECT 652.950 178.950 655.050 181.050 ;
        RECT 655.950 178.950 658.050 181.050 ;
        RECT 658.950 178.950 661.050 181.050 ;
        RECT 650.400 177.000 651.600 178.950 ;
        RECT 656.400 177.900 657.600 178.950 ;
        RECT 665.400 177.900 666.600 182.400 ;
        RECT 643.950 172.950 646.050 175.050 ;
        RECT 649.950 172.950 652.050 177.000 ;
        RECT 655.950 175.800 658.050 177.900 ;
        RECT 664.950 175.800 667.050 177.900 ;
        RECT 652.950 172.950 655.050 175.050 ;
        RECT 634.950 160.950 637.050 163.050 ;
        RECT 631.950 154.950 634.050 157.050 ;
        RECT 619.950 147.300 622.050 149.400 ;
        RECT 620.850 143.700 622.050 147.300 ;
        RECT 619.950 141.600 622.050 143.700 ;
        RECT 562.950 133.950 565.050 136.050 ;
        RECT 565.950 133.950 568.050 136.050 ;
        RECT 568.950 133.950 571.050 136.050 ;
        RECT 571.950 133.950 574.050 136.050 ;
        RECT 566.400 132.000 567.600 133.950 ;
        RECT 565.950 127.950 568.050 132.000 ;
        RECT 572.400 130.050 573.600 133.950 ;
        RECT 577.950 130.800 580.050 132.900 ;
        RECT 568.950 128.400 573.600 130.050 ;
        RECT 568.950 127.950 573.000 128.400 ;
        RECT 578.400 106.050 579.600 130.800 ;
        RECT 581.400 130.050 582.600 136.950 ;
        RECT 590.400 136.050 591.600 137.100 ;
        RECT 592.950 136.950 595.050 139.050 ;
        RECT 598.950 136.950 601.050 139.050 ;
        RECT 607.950 137.100 610.050 139.200 ;
        RECT 586.950 133.950 589.050 136.050 ;
        RECT 589.950 133.950 592.050 136.050 ;
        RECT 587.400 132.900 588.600 133.950 ;
        RECT 586.950 130.800 589.050 132.900 ;
        RECT 580.950 127.950 583.050 130.050 ;
        RECT 586.950 112.950 592.050 115.050 ;
        RECT 592.950 112.950 598.050 115.050 ;
        RECT 589.950 109.800 592.050 111.900 ;
        RECT 599.400 111.600 600.600 136.950 ;
        RECT 608.400 136.050 609.600 137.100 ;
        RECT 607.950 133.950 610.050 136.050 ;
        RECT 610.950 133.950 613.050 136.050 ;
        RECT 616.950 133.950 619.050 136.050 ;
        RECT 611.400 132.000 612.600 133.950 ;
        RECT 610.950 127.950 613.050 132.000 ;
        RECT 613.950 130.950 616.050 133.050 ;
        RECT 617.400 132.000 618.600 133.950 ;
        RECT 596.400 110.400 600.600 111.600 ;
        RECT 533.400 103.050 534.600 104.100 ;
        RECT 539.400 103.050 540.600 104.100 ;
        RECT 553.950 103.950 556.050 106.050 ;
        RECT 563.400 104.400 570.600 105.600 ;
        RECT 563.400 103.050 564.600 104.400 ;
        RECT 532.950 100.950 535.050 103.050 ;
        RECT 535.950 100.950 538.050 103.050 ;
        RECT 538.950 100.950 541.050 103.050 ;
        RECT 541.950 100.950 544.050 103.050 ;
        RECT 559.950 100.950 562.050 103.050 ;
        RECT 562.950 100.950 565.050 103.050 ;
        RECT 526.950 91.950 529.050 94.050 ;
        RECT 536.400 91.050 537.600 100.950 ;
        RECT 542.400 99.900 543.600 100.950 ;
        RECT 560.400 99.900 561.600 100.950 ;
        RECT 541.950 97.800 544.050 99.900 ;
        RECT 559.950 97.800 562.050 99.900 ;
        RECT 569.400 91.050 570.600 104.400 ;
        RECT 577.950 103.950 580.050 106.050 ;
        RECT 580.950 105.000 583.050 109.050 ;
        RECT 581.400 103.050 582.600 105.000 ;
        RECT 574.950 100.950 577.050 103.050 ;
        RECT 580.950 100.950 583.050 103.050 ;
        RECT 583.950 100.950 586.050 103.050 ;
        RECT 575.400 99.900 576.600 100.950 ;
        RECT 574.800 97.800 576.900 99.900 ;
        RECT 577.950 97.950 580.050 100.050 ;
        RECT 584.400 99.900 585.600 100.950 ;
        RECT 590.400 100.050 591.600 109.800 ;
        RECT 535.950 88.950 538.050 91.050 ;
        RECT 568.950 90.600 571.050 91.050 ;
        RECT 568.950 89.400 573.600 90.600 ;
        RECT 568.950 88.950 571.050 89.400 ;
        RECT 523.950 82.950 526.050 85.050 ;
        RECT 524.400 58.050 525.600 82.950 ;
        RECT 541.950 59.100 544.050 61.200 ;
        RECT 562.950 60.000 565.050 64.050 ;
        RECT 568.950 60.000 571.050 64.050 ;
        RECT 572.400 61.050 573.600 89.400 ;
        RECT 578.400 64.050 579.600 97.950 ;
        RECT 583.950 97.800 586.050 99.900 ;
        RECT 589.950 97.950 592.050 100.050 ;
        RECT 596.400 69.600 597.600 110.400 ;
        RECT 599.400 108.000 606.600 108.600 ;
        RECT 598.950 107.400 606.600 108.000 ;
        RECT 598.950 103.950 601.050 107.400 ;
        RECT 605.400 103.050 606.600 107.400 ;
        RECT 614.400 105.600 615.600 130.950 ;
        RECT 616.950 127.950 619.050 132.000 ;
        RECT 620.850 126.600 622.050 141.600 ;
        RECT 635.400 136.050 636.600 160.950 ;
        RECT 640.950 146.400 643.050 148.500 ;
        RECT 628.950 133.950 631.050 136.050 ;
        RECT 634.950 133.950 637.050 136.050 ;
        RECT 619.950 124.500 622.050 126.600 ;
        RECT 629.400 121.050 630.600 133.950 ;
        RECT 634.950 127.950 637.050 130.050 ;
        RECT 628.950 118.950 631.050 121.050 ;
        RECT 631.950 115.950 634.050 118.050 ;
        RECT 616.950 105.600 619.050 106.200 ;
        RECT 614.400 104.400 619.050 105.600 ;
        RECT 616.950 104.100 619.050 104.400 ;
        RECT 622.950 104.100 625.050 106.200 ;
        RECT 628.950 105.600 631.050 109.050 ;
        RECT 632.400 105.600 633.600 115.950 ;
        RECT 628.950 105.000 633.600 105.600 ;
        RECT 629.400 104.400 633.600 105.000 ;
        RECT 601.950 100.950 604.050 103.050 ;
        RECT 604.950 100.950 607.050 103.050 ;
        RECT 607.950 100.950 610.050 103.050 ;
        RECT 602.400 99.900 603.600 100.950 ;
        RECT 608.400 99.900 609.600 100.950 ;
        RECT 617.400 100.050 618.600 104.100 ;
        RECT 623.400 103.050 624.600 104.100 ;
        RECT 629.400 103.050 630.600 104.400 ;
        RECT 622.950 100.950 625.050 103.050 ;
        RECT 625.950 100.950 628.050 103.050 ;
        RECT 628.950 100.950 631.050 103.050 ;
        RECT 601.950 97.800 604.050 99.900 ;
        RECT 607.950 97.800 610.050 99.900 ;
        RECT 616.950 97.950 619.050 100.050 ;
        RECT 616.950 91.950 619.050 94.050 ;
        RECT 596.400 68.400 600.600 69.600 ;
        RECT 595.950 64.950 598.050 67.050 ;
        RECT 577.950 61.950 580.050 64.050 ;
        RECT 542.400 58.050 543.600 59.100 ;
        RECT 563.400 58.050 564.600 60.000 ;
        RECT 569.400 58.050 570.600 60.000 ;
        RECT 571.950 58.950 574.050 61.050 ;
        RECT 577.950 60.600 580.050 60.900 ;
        RECT 580.950 60.600 583.050 64.050 ;
        RECT 577.950 60.000 583.050 60.600 ;
        RECT 586.950 60.000 589.050 64.050 ;
        RECT 577.950 59.400 582.600 60.000 ;
        RECT 577.950 58.800 580.050 59.400 ;
        RECT 523.950 55.950 526.050 58.050 ;
        RECT 541.950 55.950 544.050 58.050 ;
        RECT 544.950 55.950 547.050 58.050 ;
        RECT 559.950 55.950 562.050 58.050 ;
        RECT 562.950 55.950 565.050 58.050 ;
        RECT 565.950 55.950 568.050 58.050 ;
        RECT 568.950 55.950 571.050 58.050 ;
        RECT 545.400 54.900 546.600 55.950 ;
        RECT 560.400 54.900 561.600 55.950 ;
        RECT 566.400 54.900 567.600 55.950 ;
        RECT 578.400 54.900 579.600 58.800 ;
        RECT 587.400 58.050 588.600 60.000 ;
        RECT 583.950 55.950 586.050 58.050 ;
        RECT 586.950 55.950 589.050 58.050 ;
        RECT 589.950 55.950 592.050 58.050 ;
        RECT 584.400 54.900 585.600 55.950 ;
        RECT 590.400 54.900 591.600 55.950 ;
        RECT 596.400 54.900 597.600 64.950 ;
        RECT 517.950 52.800 520.050 54.900 ;
        RECT 544.950 52.800 547.050 54.900 ;
        RECT 559.950 52.800 562.050 54.900 ;
        RECT 565.950 52.800 568.050 54.900 ;
        RECT 577.950 52.800 580.050 54.900 ;
        RECT 583.950 52.800 586.050 54.900 ;
        RECT 589.950 52.800 592.050 54.900 ;
        RECT 595.950 52.800 598.050 54.900 ;
        RECT 538.950 31.950 541.050 34.050 ;
        RECT 553.950 31.950 556.050 34.050 ;
        RECT 565.950 32.400 568.050 34.500 ;
        RECT 523.950 26.100 526.050 28.200 ;
        RECT 529.950 26.100 532.050 28.200 ;
        RECT 524.400 25.050 525.600 26.100 ;
        RECT 530.400 25.050 531.600 26.100 ;
        RECT 523.950 22.950 526.050 25.050 ;
        RECT 526.950 22.950 529.050 25.050 ;
        RECT 529.950 22.950 532.050 25.050 ;
        RECT 532.950 22.950 535.050 25.050 ;
        RECT 527.400 21.000 528.600 22.950 ;
        RECT 533.400 21.900 534.600 22.950 ;
        RECT 539.400 21.900 540.600 31.950 ;
        RECT 544.950 25.950 547.050 28.050 ;
        RECT 514.950 16.950 517.050 19.050 ;
        RECT 526.950 16.950 529.050 21.000 ;
        RECT 532.950 19.800 535.050 21.900 ;
        RECT 538.950 19.800 541.050 21.900 ;
        RECT 545.400 13.050 546.600 25.950 ;
        RECT 554.400 25.050 555.600 31.950 ;
        RECT 550.950 22.950 553.050 25.050 ;
        RECT 553.950 22.950 556.050 25.050 ;
        RECT 556.950 22.950 559.050 25.050 ;
        RECT 562.950 22.950 565.050 25.050 ;
        RECT 551.400 21.000 552.600 22.950 ;
        RECT 550.950 16.950 553.050 21.000 ;
        RECT 557.400 16.050 558.600 22.950 ;
        RECT 563.400 21.600 564.600 22.950 ;
        RECT 562.950 19.500 565.050 21.600 ;
        RECT 556.950 13.950 559.050 16.050 ;
        RECT 466.950 9.600 469.050 11.700 ;
        RECT 487.950 10.500 490.050 12.600 ;
        RECT 544.950 10.950 547.050 13.050 ;
        RECT 553.950 12.600 556.050 13.050 ;
        RECT 559.950 12.600 562.050 13.050 ;
        RECT 566.700 12.600 567.900 32.400 ;
        RECT 577.950 31.950 580.050 34.050 ;
        RECT 586.950 32.400 589.050 34.500 ;
        RECT 578.400 25.050 579.600 31.950 ;
        RECT 580.950 26.400 583.050 28.500 ;
        RECT 571.950 22.950 574.050 25.050 ;
        RECT 577.950 22.950 580.050 25.050 ;
        RECT 572.400 13.050 573.600 22.950 ;
        RECT 581.400 16.050 582.600 26.400 ;
        RECT 586.950 17.400 588.150 32.400 ;
        RECT 589.950 26.400 592.050 28.500 ;
        RECT 590.400 25.050 591.600 26.400 ;
        RECT 589.950 22.950 592.050 25.050 ;
        RECT 580.950 13.950 583.050 16.050 ;
        RECT 586.950 15.300 589.050 17.400 ;
        RECT 553.950 11.400 562.050 12.600 ;
        RECT 553.950 10.950 556.050 11.400 ;
        RECT 559.950 10.950 562.050 11.400 ;
        RECT 565.950 10.500 568.050 12.600 ;
        RECT 571.950 10.950 574.050 13.050 ;
        RECT 586.950 11.700 588.150 15.300 ;
        RECT 586.950 9.600 589.050 11.700 ;
        RECT 599.400 7.050 600.600 68.400 ;
        RECT 607.950 59.100 610.050 61.200 ;
        RECT 608.400 58.050 609.600 59.100 ;
        RECT 604.950 55.950 607.050 58.050 ;
        RECT 607.950 55.950 610.050 58.050 ;
        RECT 610.950 55.950 613.050 58.050 ;
        RECT 605.400 54.900 606.600 55.950 ;
        RECT 611.400 54.900 612.600 55.950 ;
        RECT 604.950 52.800 607.050 54.900 ;
        RECT 610.950 52.800 613.050 54.900 ;
        RECT 612.000 30.600 616.050 31.050 ;
        RECT 611.400 28.950 616.050 30.600 ;
        RECT 611.400 25.050 612.600 28.950 ;
        RECT 617.400 28.200 618.600 91.950 ;
        RECT 626.400 91.050 627.600 100.950 ;
        RECT 625.950 88.950 628.050 91.050 ;
        RECT 635.400 64.050 636.600 127.950 ;
        RECT 641.100 126.600 642.300 146.400 ;
        RECT 643.950 137.400 646.050 139.500 ;
        RECT 644.400 136.050 645.600 137.400 ;
        RECT 649.950 136.950 652.050 139.050 ;
        RECT 643.950 133.950 646.050 136.050 ;
        RECT 640.950 124.500 643.050 126.600 ;
        RECT 650.400 112.050 651.600 136.950 ;
        RECT 653.400 130.050 654.600 172.950 ;
        RECT 668.400 157.050 669.600 274.800 ;
        RECT 670.950 259.950 673.050 262.050 ;
        RECT 679.950 260.100 682.050 262.200 ;
        RECT 686.400 262.050 687.600 283.950 ;
        RECT 671.400 241.050 672.600 259.950 ;
        RECT 680.400 259.050 681.600 260.100 ;
        RECT 685.950 259.950 688.050 262.050 ;
        RECT 676.950 256.950 679.050 259.050 ;
        RECT 679.950 256.950 682.050 259.050 ;
        RECT 682.950 256.950 685.050 259.050 ;
        RECT 673.950 253.950 676.050 256.050 ;
        RECT 677.400 255.000 678.600 256.950 ;
        RECT 683.400 255.900 684.600 256.950 ;
        RECT 670.950 238.950 673.050 241.050 ;
        RECT 674.400 219.600 675.600 253.950 ;
        RECT 676.950 250.950 679.050 255.000 ;
        RECT 682.950 253.800 685.050 255.900 ;
        RECT 685.950 253.950 688.050 256.050 ;
        RECT 689.400 255.900 690.600 286.800 ;
        RECT 695.400 261.600 696.600 289.950 ;
        RECT 701.400 289.050 702.600 293.100 ;
        RECT 700.950 286.950 703.050 289.050 ;
        RECT 700.950 280.950 703.050 283.050 ;
        RECT 697.950 271.950 700.050 274.050 ;
        RECT 692.400 260.400 696.600 261.600 ;
        RECT 674.400 218.400 678.600 219.600 ;
        RECT 677.400 214.050 678.600 218.400 ;
        RECT 682.950 215.100 685.050 217.200 ;
        RECT 686.400 217.050 687.600 253.950 ;
        RECT 688.950 253.800 691.050 255.900 ;
        RECT 692.400 253.050 693.600 260.400 ;
        RECT 698.400 259.050 699.600 271.950 ;
        RECT 701.400 270.600 702.600 280.950 ;
        RECT 704.400 280.050 705.600 295.950 ;
        RECT 707.400 288.900 708.600 331.950 ;
        RECT 710.400 298.050 711.600 338.400 ;
        RECT 718.950 338.100 721.050 340.200 ;
        RECT 724.950 339.000 727.050 343.050 ;
        RECT 728.400 340.050 729.600 343.950 ;
        RECT 719.400 337.050 720.600 338.100 ;
        RECT 725.400 337.050 726.600 339.000 ;
        RECT 727.950 337.950 730.050 340.050 ;
        RECT 730.950 337.950 733.050 340.050 ;
        RECT 715.950 334.950 718.050 337.050 ;
        RECT 718.950 334.950 721.050 337.050 ;
        RECT 721.950 334.950 724.050 337.050 ;
        RECT 724.950 334.950 727.050 337.050 ;
        RECT 716.400 333.900 717.600 334.950 ;
        RECT 722.400 333.900 723.600 334.950 ;
        RECT 715.950 331.800 718.050 333.900 ;
        RECT 721.950 331.800 724.050 333.900 ;
        RECT 727.950 331.950 730.050 334.050 ;
        RECT 731.400 333.900 732.600 337.950 ;
        RECT 715.950 301.950 718.050 304.050 ;
        RECT 709.950 295.950 712.050 298.050 ;
        RECT 716.400 295.200 717.600 301.950 ;
        RECT 715.950 293.100 718.050 295.200 ;
        RECT 716.400 292.050 717.600 293.100 ;
        RECT 722.400 292.050 723.600 331.800 ;
        RECT 728.400 300.600 729.600 331.950 ;
        RECT 730.950 331.800 733.050 333.900 ;
        RECT 725.400 299.400 729.600 300.600 ;
        RECT 725.400 295.050 726.600 299.400 ;
        RECT 734.400 298.050 735.600 364.950 ;
        RECT 736.950 364.800 739.050 366.900 ;
        RECT 742.950 364.800 745.050 366.900 ;
        RECT 749.400 366.000 754.050 367.050 ;
        RECT 748.950 364.950 754.050 366.000 ;
        RECT 748.950 361.950 751.050 364.950 ;
        RECT 755.400 355.050 756.600 370.950 ;
        RECT 754.950 352.950 757.050 355.050 ;
        RECT 748.950 346.950 751.050 349.050 ;
        RECT 736.950 340.950 739.050 343.050 ;
        RECT 737.400 301.050 738.600 340.950 ;
        RECT 742.950 338.100 745.050 340.200 ;
        RECT 743.400 337.050 744.600 338.100 ;
        RECT 749.400 337.050 750.600 346.950 ;
        RECT 742.950 334.950 745.050 337.050 ;
        RECT 745.950 334.950 748.050 337.050 ;
        RECT 748.950 334.950 751.050 337.050 ;
        RECT 751.950 334.950 754.050 337.050 ;
        RECT 746.400 328.050 747.600 334.950 ;
        RECT 752.400 333.900 753.600 334.950 ;
        RECT 751.950 331.800 754.050 333.900 ;
        RECT 745.950 325.950 748.050 328.050 ;
        RECT 745.950 322.800 748.050 324.900 ;
        RECT 736.950 298.950 739.050 301.050 ;
        RECT 727.950 295.950 730.050 298.050 ;
        RECT 733.950 295.950 736.050 298.050 ;
        RECT 724.950 292.950 727.050 295.050 ;
        RECT 712.950 289.950 715.050 292.050 ;
        RECT 715.950 289.950 718.050 292.050 ;
        RECT 718.950 289.950 721.050 292.050 ;
        RECT 721.950 289.950 724.050 292.050 ;
        RECT 706.950 286.800 709.050 288.900 ;
        RECT 709.950 286.950 712.050 289.050 ;
        RECT 713.400 288.900 714.600 289.950 ;
        RECT 710.400 283.050 711.600 286.950 ;
        RECT 712.950 286.800 715.050 288.900 ;
        RECT 719.400 283.050 720.600 289.950 ;
        RECT 709.950 280.950 712.050 283.050 ;
        RECT 718.950 280.950 721.050 283.050 ;
        RECT 703.950 277.950 706.050 280.050 ;
        RECT 701.400 269.400 705.600 270.600 ;
        RECT 704.400 262.200 705.600 269.400 ;
        RECT 712.950 268.950 715.050 271.050 ;
        RECT 703.950 260.100 706.050 262.200 ;
        RECT 704.400 259.050 705.600 260.100 ;
        RECT 697.950 256.950 700.050 259.050 ;
        RECT 700.950 256.950 703.050 259.050 ;
        RECT 703.950 256.950 706.050 259.050 ;
        RECT 706.950 256.950 709.050 259.050 ;
        RECT 701.400 255.000 702.600 256.950 ;
        RECT 707.400 255.900 708.600 256.950 ;
        RECT 691.950 250.950 694.050 253.050 ;
        RECT 700.950 250.950 703.050 255.000 ;
        RECT 706.950 253.800 709.050 255.900 ;
        RECT 713.400 253.050 714.600 268.950 ;
        RECT 728.400 268.050 729.600 295.950 ;
        RECT 730.950 292.950 733.050 295.050 ;
        RECT 739.950 293.100 742.050 295.200 ;
        RECT 727.950 265.950 730.050 268.050 ;
        RECT 721.950 260.100 724.050 262.200 ;
        RECT 727.950 260.100 730.050 262.200 ;
        RECT 731.400 262.050 732.600 292.950 ;
        RECT 740.400 292.050 741.600 293.100 ;
        RECT 746.400 292.050 747.600 322.800 ;
        RECT 751.950 307.950 754.050 310.050 ;
        RECT 736.950 289.950 739.050 292.050 ;
        RECT 739.950 289.950 742.050 292.050 ;
        RECT 742.950 289.950 745.050 292.050 ;
        RECT 745.950 289.950 748.050 292.050 ;
        RECT 737.400 288.900 738.600 289.950 ;
        RECT 743.400 288.900 744.600 289.950 ;
        RECT 736.950 286.800 739.050 288.900 ;
        RECT 742.950 286.800 745.050 288.900 ;
        RECT 745.950 274.950 748.050 277.050 ;
        RECT 733.950 265.950 736.050 268.050 ;
        RECT 742.950 265.950 745.050 268.050 ;
        RECT 722.400 259.050 723.600 260.100 ;
        RECT 728.400 259.050 729.600 260.100 ;
        RECT 730.950 259.950 733.050 262.050 ;
        RECT 718.950 256.950 721.050 259.050 ;
        RECT 721.950 256.950 724.050 259.050 ;
        RECT 724.950 256.950 727.050 259.050 ;
        RECT 727.950 256.950 730.050 259.050 ;
        RECT 719.400 255.900 720.600 256.950 ;
        RECT 718.950 253.800 721.050 255.900 ;
        RECT 725.400 255.000 726.600 256.950 ;
        RECT 734.400 255.900 735.600 265.950 ;
        RECT 743.400 262.050 744.600 265.950 ;
        RECT 736.950 259.950 739.050 262.050 ;
        RECT 739.950 259.950 742.050 262.050 ;
        RECT 742.950 259.950 745.050 262.050 ;
        RECT 712.950 250.950 715.050 253.050 ;
        RECT 724.950 250.950 727.050 255.000 ;
        RECT 733.950 253.800 736.050 255.900 ;
        RECT 721.950 238.950 724.050 241.050 ;
        RECT 688.950 232.950 691.050 235.050 ;
        RECT 718.950 232.950 721.050 235.050 ;
        RECT 683.400 214.050 684.600 215.100 ;
        RECT 685.950 214.950 688.050 217.050 ;
        RECT 673.950 211.950 676.050 214.050 ;
        RECT 676.950 211.950 679.050 214.050 ;
        RECT 679.950 211.950 682.050 214.050 ;
        RECT 682.950 211.950 685.050 214.050 ;
        RECT 674.400 186.600 675.600 211.950 ;
        RECT 680.400 202.050 681.600 211.950 ;
        RECT 679.950 199.950 682.050 202.050 ;
        RECT 682.950 193.950 685.050 196.050 ;
        RECT 671.400 186.000 675.600 186.600 ;
        RECT 670.950 185.400 675.600 186.000 ;
        RECT 670.950 181.950 673.050 185.400 ;
        RECT 676.950 183.000 679.050 187.050 ;
        RECT 677.400 181.050 678.600 183.000 ;
        RECT 683.400 181.050 684.600 193.950 ;
        RECT 689.400 183.600 690.600 232.950 ;
        RECT 691.950 229.950 694.050 232.050 ;
        RECT 692.400 186.600 693.600 229.950 ;
        RECT 697.800 219.300 699.900 221.400 ;
        RECT 707.400 220.500 709.500 222.600 ;
        RECT 694.950 214.050 697.050 217.050 ;
        RECT 695.400 211.950 697.500 214.050 ;
        RECT 695.400 190.050 696.600 211.950 ;
        RECT 698.700 210.300 699.600 219.300 ;
        RECT 701.100 215.700 703.200 217.800 ;
        RECT 704.400 216.900 705.600 219.450 ;
        RECT 702.300 213.300 703.200 215.700 ;
        RECT 704.100 214.800 706.200 216.900 ;
        RECT 708.000 213.300 709.050 220.500 ;
        RECT 719.400 214.050 720.600 232.950 ;
        RECT 702.300 212.100 709.050 213.300 ;
        RECT 705.150 210.300 707.250 211.200 ;
        RECT 698.700 209.100 707.250 210.300 ;
        RECT 700.200 207.300 702.300 209.100 ;
        RECT 704.100 206.100 706.200 208.200 ;
        RECT 708.150 206.700 709.050 212.100 ;
        RECT 709.950 211.950 712.050 214.050 ;
        RECT 715.800 211.950 717.900 214.050 ;
        RECT 718.950 211.950 721.050 214.050 ;
        RECT 710.400 209.400 711.600 211.950 ;
        RECT 700.950 199.950 703.050 202.050 ;
        RECT 694.950 187.950 697.050 190.050 ;
        RECT 692.400 185.400 696.600 186.600 ;
        RECT 689.400 182.400 693.600 183.600 ;
        RECT 673.950 178.950 676.050 181.050 ;
        RECT 676.950 178.950 679.050 181.050 ;
        RECT 679.950 178.950 682.050 181.050 ;
        RECT 682.950 178.950 685.050 181.050 ;
        RECT 685.950 178.950 688.050 181.050 ;
        RECT 674.400 177.000 675.600 178.950 ;
        RECT 673.950 172.950 676.050 177.000 ;
        RECT 680.400 171.600 681.600 178.950 ;
        RECT 686.400 177.900 687.600 178.950 ;
        RECT 685.950 175.800 688.050 177.900 ;
        RECT 680.400 170.400 684.600 171.600 ;
        RECT 679.950 166.950 682.050 169.050 ;
        RECT 667.950 154.950 670.050 157.050 ;
        RECT 673.950 147.300 676.050 149.400 ;
        RECT 674.850 143.700 676.050 147.300 ;
        RECT 673.950 141.600 676.050 143.700 ;
        RECT 655.950 136.950 658.050 139.050 ;
        RECT 661.950 137.100 664.050 139.200 ;
        RECT 652.950 127.950 655.050 130.050 ;
        RECT 656.400 118.050 657.600 136.950 ;
        RECT 662.400 136.050 663.600 137.100 ;
        RECT 661.950 133.950 664.050 136.050 ;
        RECT 664.950 133.950 667.050 136.050 ;
        RECT 670.950 133.950 673.050 136.050 ;
        RECT 665.400 132.600 666.600 133.950 ;
        RECT 671.400 132.600 672.600 133.950 ;
        RECT 665.400 131.400 672.600 132.600 ;
        RECT 674.850 126.600 676.050 141.600 ;
        RECT 680.400 130.050 681.600 166.950 ;
        RECT 679.950 127.950 682.050 130.050 ;
        RECT 673.950 124.500 676.050 126.600 ;
        RECT 683.400 118.050 684.600 170.400 ;
        RECT 692.400 169.050 693.600 182.400 ;
        RECT 691.950 166.950 694.050 169.050 ;
        RECT 695.400 163.050 696.600 185.400 ;
        RECT 701.400 181.050 702.600 199.950 ;
        RECT 704.400 199.050 705.600 206.100 ;
        RECT 707.400 204.600 709.500 206.700 ;
        RECT 703.800 196.950 705.900 199.050 ;
        RECT 706.950 196.950 709.050 199.050 ;
        RECT 707.400 181.050 708.600 196.950 ;
        RECT 716.400 196.050 717.600 211.950 ;
        RECT 722.400 204.600 723.600 238.950 ;
        RECT 737.400 229.050 738.600 259.950 ;
        RECT 740.400 238.050 741.600 259.950 ;
        RECT 746.400 259.050 747.600 274.950 ;
        RECT 752.400 268.050 753.600 307.950 ;
        RECT 758.400 304.050 759.600 373.950 ;
        RECT 761.400 351.600 762.600 409.950 ;
        RECT 764.400 394.050 765.600 427.950 ;
        RECT 767.400 418.050 768.600 431.400 ;
        RECT 770.400 421.050 771.600 442.950 ;
        RECT 775.950 439.950 778.050 444.000 ;
        RECT 781.950 442.950 784.050 445.050 ;
        RECT 778.950 439.950 781.050 442.050 ;
        RECT 776.400 421.050 777.600 439.950 ;
        RECT 779.400 433.050 780.600 439.950 ;
        RECT 778.950 430.950 781.050 433.050 ;
        RECT 769.950 418.950 772.050 421.050 ;
        RECT 772.800 420.000 774.900 421.050 ;
        RECT 772.800 418.950 775.050 420.000 ;
        RECT 775.950 418.950 778.050 421.050 ;
        RECT 766.950 415.950 769.050 418.050 ;
        RECT 772.950 417.000 775.050 418.950 ;
        RECT 773.400 415.050 774.600 417.000 ;
        RECT 769.950 412.950 772.050 415.050 ;
        RECT 772.950 412.950 775.050 415.050 ;
        RECT 775.950 412.950 778.050 415.050 ;
        RECT 766.950 409.950 769.050 412.050 ;
        RECT 763.950 391.950 766.050 394.050 ;
        RECT 767.400 388.050 768.600 409.950 ;
        RECT 770.400 403.050 771.600 412.950 ;
        RECT 776.400 411.900 777.600 412.950 ;
        RECT 775.950 409.800 778.050 411.900 ;
        RECT 769.950 400.950 772.050 403.050 ;
        RECT 782.400 388.050 783.600 442.950 ;
        RECT 766.950 385.950 769.050 388.050 ;
        RECT 781.950 385.950 784.050 388.050 ;
        RECT 766.800 375.300 768.900 377.400 ;
        RECT 776.400 376.500 778.500 378.600 ;
        RECT 764.400 370.050 765.600 372.600 ;
        RECT 764.400 367.950 766.500 370.050 ;
        RECT 767.700 366.300 768.600 375.300 ;
        RECT 770.100 371.700 772.200 373.800 ;
        RECT 773.400 372.900 774.600 375.450 ;
        RECT 771.300 369.300 772.200 371.700 ;
        RECT 773.100 370.800 775.200 372.900 ;
        RECT 777.000 369.300 778.050 376.500 ;
        RECT 771.300 368.100 778.050 369.300 ;
        RECT 774.150 366.300 776.250 367.200 ;
        RECT 767.700 365.100 776.250 366.300 ;
        RECT 763.950 361.800 766.050 363.900 ;
        RECT 769.200 363.300 771.300 365.100 ;
        RECT 773.100 362.100 775.200 364.200 ;
        RECT 777.150 362.700 778.050 368.100 ;
        RECT 778.950 367.950 781.050 370.050 ;
        RECT 779.400 365.400 780.600 367.950 ;
        RECT 764.400 358.050 765.600 361.800 ;
        RECT 763.950 355.950 766.050 358.050 ;
        RECT 761.400 350.400 765.600 351.600 ;
        RECT 760.950 346.950 763.050 349.050 ;
        RECT 761.400 333.900 762.600 346.950 ;
        RECT 764.400 340.050 765.600 350.400 ;
        RECT 773.400 343.050 774.600 362.100 ;
        RECT 776.400 360.600 778.500 362.700 ;
        RECT 778.950 355.950 781.050 358.050 ;
        RECT 775.950 352.950 778.050 355.050 ;
        RECT 772.950 342.600 775.050 343.050 ;
        RECT 770.400 341.400 775.050 342.600 ;
        RECT 770.400 340.200 771.600 341.400 ;
        RECT 772.950 340.950 775.050 341.400 ;
        RECT 763.950 337.950 766.050 340.050 ;
        RECT 769.950 338.100 772.050 340.200 ;
        RECT 770.400 337.050 771.600 338.100 ;
        RECT 776.400 337.050 777.600 352.950 ;
        RECT 779.400 340.050 780.600 355.950 ;
        RECT 781.950 340.950 784.050 343.050 ;
        RECT 778.950 337.950 781.050 340.050 ;
        RECT 766.950 334.950 769.050 337.050 ;
        RECT 769.950 334.950 772.050 337.050 ;
        RECT 772.950 334.950 775.050 337.050 ;
        RECT 775.950 334.950 778.050 337.050 ;
        RECT 760.950 331.800 763.050 333.900 ;
        RECT 763.950 331.950 766.050 334.050 ;
        RECT 767.400 333.900 768.600 334.950 ;
        RECT 773.400 333.900 774.600 334.950 ;
        RECT 764.400 322.050 765.600 331.950 ;
        RECT 766.950 331.800 769.050 333.900 ;
        RECT 772.950 331.800 775.050 333.900 ;
        RECT 778.950 331.950 781.050 334.050 ;
        RECT 782.400 333.900 783.600 340.950 ;
        RECT 779.400 328.050 780.600 331.950 ;
        RECT 781.950 331.800 784.050 333.900 ;
        RECT 778.950 325.950 781.050 328.050 ;
        RECT 763.950 319.950 766.050 322.050 ;
        RECT 778.950 313.950 781.050 316.050 ;
        RECT 757.950 301.950 760.050 304.050 ;
        RECT 775.950 301.950 778.050 304.050 ;
        RECT 754.950 298.950 757.050 301.050 ;
        RECT 755.400 288.900 756.600 298.950 ;
        RECT 757.950 292.950 760.050 298.050 ;
        RECT 760.950 294.000 763.050 298.050 ;
        RECT 766.950 294.000 769.050 298.050 ;
        RECT 761.400 292.050 762.600 294.000 ;
        RECT 767.400 292.050 768.600 294.000 ;
        RECT 760.950 289.950 763.050 292.050 ;
        RECT 763.950 289.950 766.050 292.050 ;
        RECT 766.950 289.950 769.050 292.050 ;
        RECT 769.950 289.950 772.050 292.050 ;
        RECT 764.400 288.900 765.600 289.950 ;
        RECT 754.950 286.800 757.050 288.900 ;
        RECT 763.950 286.800 766.050 288.900 ;
        RECT 770.400 280.050 771.600 289.950 ;
        RECT 769.950 277.950 772.050 280.050 ;
        RECT 760.950 271.950 763.050 274.050 ;
        RECT 751.950 265.950 754.050 268.050 ;
        RECT 751.950 260.100 754.050 262.200 ;
        RECT 752.400 259.050 753.600 260.100 ;
        RECT 745.950 256.950 748.050 259.050 ;
        RECT 748.950 256.950 751.050 259.050 ;
        RECT 751.950 256.950 754.050 259.050 ;
        RECT 754.950 256.950 757.050 259.050 ;
        RECT 739.950 235.950 742.050 238.050 ;
        RECT 749.400 235.050 750.600 256.950 ;
        RECT 751.950 250.950 754.050 253.050 ;
        RECT 748.950 232.950 751.050 235.050 ;
        RECT 736.950 226.950 739.050 229.050 ;
        RECT 748.950 226.950 751.050 229.050 ;
        RECT 730.500 220.500 732.600 222.600 ;
        RECT 727.950 211.950 730.050 214.050 ;
        RECT 730.950 213.300 732.000 220.500 ;
        RECT 734.400 216.900 735.600 219.450 ;
        RECT 740.100 219.300 742.200 221.400 ;
        RECT 733.800 214.800 735.900 216.900 ;
        RECT 736.800 215.700 738.900 217.800 ;
        RECT 736.800 213.300 737.700 215.700 ;
        RECT 730.950 212.100 737.700 213.300 ;
        RECT 728.400 209.400 729.600 211.950 ;
        RECT 730.950 206.700 731.850 212.100 ;
        RECT 732.750 210.300 734.850 211.200 ;
        RECT 740.400 210.300 741.300 219.300 ;
        RECT 743.400 214.050 744.600 216.600 ;
        RECT 742.500 211.950 744.600 214.050 ;
        RECT 745.950 211.950 748.050 214.050 ;
        RECT 732.750 209.100 741.300 210.300 ;
        RECT 730.500 204.600 732.600 206.700 ;
        RECT 733.800 206.100 735.900 208.200 ;
        RECT 737.700 207.300 739.800 209.100 ;
        RECT 734.400 204.900 735.600 206.100 ;
        RECT 722.400 203.400 726.600 204.600 ;
        RECT 721.950 199.950 724.050 202.050 ;
        RECT 715.950 193.950 718.050 196.050 ;
        RECT 715.950 187.950 718.050 190.050 ;
        RECT 700.950 178.950 703.050 181.050 ;
        RECT 703.950 178.950 706.050 181.050 ;
        RECT 706.950 178.950 709.050 181.050 ;
        RECT 694.950 160.950 697.050 163.050 ;
        RECT 694.950 146.400 697.050 148.500 ;
        RECT 688.950 142.950 691.050 145.050 ;
        RECT 689.400 136.050 690.600 142.950 ;
        RECT 688.950 133.950 691.050 136.050 ;
        RECT 688.950 127.950 691.050 130.050 ;
        RECT 655.950 115.950 658.050 118.050 ;
        RECT 670.950 115.950 673.050 118.050 ;
        RECT 682.950 115.950 685.050 118.050 ;
        RECT 649.950 109.950 652.050 112.050 ;
        RECT 658.950 110.400 661.050 112.500 ;
        RECT 649.950 104.100 652.050 106.200 ;
        RECT 655.950 104.400 658.050 106.500 ;
        RECT 650.400 103.050 651.600 104.100 ;
        RECT 656.400 103.050 657.600 104.400 ;
        RECT 646.950 100.950 649.050 103.050 ;
        RECT 649.950 100.950 652.050 103.050 ;
        RECT 655.950 100.950 658.050 103.050 ;
        RECT 643.950 64.950 646.050 67.050 ;
        RECT 634.950 61.950 637.050 64.050 ;
        RECT 619.950 59.100 622.050 61.200 ;
        RECT 625.950 59.100 628.050 61.200 ;
        RECT 620.400 55.050 621.600 59.100 ;
        RECT 626.400 58.050 627.600 59.100 ;
        RECT 635.400 58.050 636.600 61.950 ;
        RECT 644.400 58.050 645.600 64.950 ;
        RECT 647.400 64.050 648.600 100.950 ;
        RECT 652.950 97.950 655.050 100.050 ;
        RECT 646.950 61.950 649.050 64.050 ;
        RECT 625.950 55.950 628.050 58.050 ;
        RECT 628.950 55.950 631.050 58.050 ;
        RECT 634.950 55.950 637.050 58.050 ;
        RECT 640.950 55.950 643.050 58.050 ;
        RECT 643.950 55.950 646.050 58.050 ;
        RECT 646.950 55.950 649.050 58.050 ;
        RECT 619.950 52.950 622.050 55.050 ;
        RECT 629.400 54.900 630.600 55.950 ;
        RECT 641.400 54.900 642.600 55.950 ;
        RECT 647.400 54.900 648.600 55.950 ;
        RECT 653.400 54.900 654.600 97.950 ;
        RECT 659.850 95.400 661.050 110.400 ;
        RECT 671.400 106.050 672.600 115.950 ;
        RECT 679.950 110.400 682.050 112.500 ;
        RECT 670.950 103.950 673.050 106.050 ;
        RECT 673.950 100.950 676.050 103.050 ;
        RECT 674.400 99.600 675.600 100.950 ;
        RECT 673.950 97.500 676.050 99.600 ;
        RECT 658.950 93.300 661.050 95.400 ;
        RECT 659.850 89.700 661.050 93.300 ;
        RECT 673.950 91.950 676.050 94.050 ;
        RECT 658.950 87.600 661.050 89.700 ;
        RECT 667.950 59.100 670.050 61.200 ;
        RECT 668.400 58.050 669.600 59.100 ;
        RECT 674.400 58.050 675.600 91.950 ;
        RECT 680.100 90.600 681.300 110.400 ;
        RECT 682.950 100.950 685.050 103.050 ;
        RECT 683.400 99.600 684.600 100.950 ;
        RECT 682.950 98.400 687.600 99.600 ;
        RECT 682.950 97.500 685.050 98.400 ;
        RECT 679.950 88.500 682.050 90.600 ;
        RECT 679.950 59.100 682.050 61.200 ;
        RECT 686.400 60.600 687.600 98.400 ;
        RECT 689.400 79.050 690.600 127.950 ;
        RECT 695.100 126.600 696.300 146.400 ;
        RECT 697.950 138.000 700.050 142.050 ;
        RECT 698.400 136.050 699.600 138.000 ;
        RECT 697.950 133.950 700.050 136.050 ;
        RECT 694.950 124.500 697.050 126.600 ;
        RECT 704.400 124.050 705.600 178.950 ;
        RECT 716.400 172.050 717.600 187.950 ;
        RECT 722.400 181.050 723.600 199.950 ;
        RECT 725.400 187.050 726.600 203.400 ;
        RECT 733.950 202.800 736.050 204.900 ;
        RECT 746.400 199.050 747.600 211.950 ;
        RECT 749.400 202.050 750.600 226.950 ;
        RECT 748.950 199.950 751.050 202.050 ;
        RECT 745.950 196.950 748.050 199.050 ;
        RECT 724.950 184.950 727.050 187.050 ;
        RECT 730.950 184.950 733.050 187.050 ;
        RECT 721.950 178.950 724.050 181.050 ;
        RECT 724.950 178.950 727.050 181.050 ;
        RECT 715.950 169.950 718.050 172.050 ;
        RECT 706.950 142.950 709.050 145.050 ;
        RECT 707.400 127.050 708.600 142.950 ;
        RECT 725.400 142.050 726.600 178.950 ;
        RECT 715.950 137.100 718.050 142.050 ;
        RECT 724.950 139.950 727.050 142.050 ;
        RECT 721.950 137.100 724.050 139.200 ;
        RECT 716.400 136.050 717.600 137.100 ;
        RECT 722.400 136.050 723.600 137.100 ;
        RECT 712.950 133.950 715.050 136.050 ;
        RECT 715.950 133.950 718.050 136.050 ;
        RECT 718.950 133.950 721.050 136.050 ;
        RECT 721.950 133.950 724.050 136.050 ;
        RECT 724.950 133.950 727.050 136.050 ;
        RECT 713.400 132.900 714.600 133.950 ;
        RECT 712.950 130.800 715.050 132.900 ;
        RECT 715.950 127.950 718.050 130.050 ;
        RECT 706.950 124.950 709.050 127.050 ;
        RECT 703.950 121.950 706.050 124.050 ;
        RECT 700.950 112.950 703.050 115.050 ;
        RECT 691.950 109.950 694.050 112.050 ;
        RECT 692.400 99.600 693.600 109.950 ;
        RECT 701.400 103.050 702.600 112.950 ;
        RECT 706.950 104.100 709.050 106.200 ;
        RECT 707.400 103.050 708.600 104.100 ;
        RECT 700.950 100.950 703.050 103.050 ;
        RECT 703.950 100.950 706.050 103.050 ;
        RECT 706.950 100.950 709.050 103.050 ;
        RECT 709.950 100.950 712.050 103.050 ;
        RECT 691.950 97.500 694.050 99.600 ;
        RECT 704.400 88.050 705.600 100.950 ;
        RECT 710.400 94.050 711.600 100.950 ;
        RECT 716.400 94.050 717.600 127.950 ;
        RECT 719.400 127.050 720.600 133.950 ;
        RECT 718.950 124.950 721.050 127.050 ;
        RECT 725.400 124.050 726.600 133.950 ;
        RECT 727.950 130.950 730.050 133.050 ;
        RECT 728.400 124.050 729.600 130.950 ;
        RECT 724.800 121.950 726.900 124.050 ;
        RECT 727.950 121.950 730.050 124.050 ;
        RECT 724.950 104.100 727.050 106.200 ;
        RECT 731.400 106.050 732.600 184.950 ;
        RECT 739.950 183.000 742.050 187.050 ;
        RECT 740.400 181.050 741.600 183.000 ;
        RECT 746.400 181.050 747.600 196.950 ;
        RECT 752.400 183.600 753.600 250.950 ;
        RECT 755.400 232.050 756.600 256.950 ;
        RECT 757.950 250.950 760.050 256.050 ;
        RECT 754.950 229.950 757.050 232.050 ;
        RECT 761.400 220.200 762.600 271.950 ;
        RECT 770.400 268.050 771.600 277.950 ;
        RECT 776.400 274.050 777.600 301.950 ;
        RECT 775.950 271.950 778.050 274.050 ;
        RECT 763.950 265.950 766.050 268.050 ;
        RECT 769.950 265.950 772.050 268.050 ;
        RECT 764.400 255.900 765.600 265.950 ;
        RECT 772.950 261.000 775.050 265.050 ;
        RECT 779.400 262.050 780.600 313.950 ;
        RECT 785.400 298.050 786.600 478.950 ;
        RECT 788.400 454.050 789.600 484.950 ;
        RECT 791.400 475.050 792.600 490.950 ;
        RECT 797.400 487.050 798.600 499.950 ;
        RECT 796.950 484.950 799.050 487.050 ;
        RECT 790.950 472.950 793.050 475.050 ;
        RECT 800.400 469.050 801.600 505.950 ;
        RECT 811.950 502.050 814.050 505.050 ;
        RECT 808.950 501.000 814.050 502.050 ;
        RECT 808.950 500.400 813.600 501.000 ;
        RECT 808.950 499.950 813.000 500.400 ;
        RECT 805.950 495.000 808.050 499.050 ;
        RECT 806.400 493.050 807.600 495.000 ;
        RECT 811.950 494.100 814.050 496.200 ;
        RECT 815.400 495.600 816.600 520.950 ;
        RECT 818.400 511.050 819.600 523.950 ;
        RECT 823.950 520.950 826.050 523.050 ;
        RECT 817.950 508.950 820.050 511.050 ;
        RECT 820.950 505.950 823.050 508.050 ;
        RECT 815.400 494.400 819.600 495.600 ;
        RECT 812.400 493.050 813.600 494.100 ;
        RECT 805.950 490.950 808.050 493.050 ;
        RECT 808.950 490.950 811.050 493.050 ;
        RECT 811.950 490.950 814.050 493.050 ;
        RECT 805.950 481.950 808.050 484.050 ;
        RECT 799.950 466.950 802.050 469.050 ;
        RECT 806.400 460.050 807.600 481.950 ;
        RECT 809.400 463.050 810.600 490.950 ;
        RECT 814.950 487.950 817.050 490.050 ;
        RECT 811.950 466.950 814.050 469.050 ;
        RECT 808.950 460.950 811.050 463.050 ;
        RECT 805.950 457.950 808.050 460.050 ;
        RECT 796.500 454.500 798.600 456.600 ;
        RECT 787.950 451.950 790.050 454.050 ;
        RECT 787.950 445.950 790.050 448.050 ;
        RECT 793.950 445.950 796.050 448.050 ;
        RECT 796.950 447.300 798.000 454.500 ;
        RECT 800.400 450.900 801.600 453.450 ;
        RECT 806.100 453.300 808.200 455.400 ;
        RECT 799.800 448.800 801.900 450.900 ;
        RECT 802.800 449.700 804.900 451.800 ;
        RECT 802.800 447.300 803.700 449.700 ;
        RECT 796.950 446.100 803.700 447.300 ;
        RECT 788.400 435.600 789.600 445.950 ;
        RECT 794.400 443.400 795.600 445.950 ;
        RECT 796.950 440.700 797.850 446.100 ;
        RECT 798.750 444.300 800.850 445.200 ;
        RECT 806.400 444.300 807.300 453.300 ;
        RECT 809.400 448.050 810.600 450.600 ;
        RECT 808.500 445.950 810.600 448.050 ;
        RECT 798.750 443.100 807.300 444.300 ;
        RECT 796.500 438.600 798.600 440.700 ;
        RECT 799.800 440.100 801.900 442.200 ;
        RECT 803.700 441.300 805.800 443.100 ;
        RECT 790.950 435.600 793.050 436.050 ;
        RECT 788.400 434.400 793.050 435.600 ;
        RECT 790.950 433.950 793.050 434.400 ;
        RECT 791.400 420.600 792.600 433.950 ;
        RECT 800.400 430.050 801.600 440.100 ;
        RECT 799.950 427.950 802.050 430.050 ;
        RECT 805.950 427.950 808.050 430.050 ;
        RECT 791.400 419.400 795.600 420.600 ;
        RECT 794.400 415.050 795.600 419.400 ;
        RECT 790.950 412.950 793.050 415.050 ;
        RECT 793.950 412.950 796.050 415.050 ;
        RECT 799.950 412.950 802.050 415.050 ;
        RECT 791.400 411.900 792.600 412.950 ;
        RECT 790.950 409.800 793.050 411.900 ;
        RECT 796.950 409.950 799.050 412.050 ;
        RECT 787.950 382.950 790.050 385.050 ;
        RECT 788.400 370.050 789.600 382.950 ;
        RECT 797.400 373.200 798.600 409.950 ;
        RECT 800.400 397.050 801.600 412.950 ;
        RECT 806.400 409.050 807.600 427.950 ;
        RECT 808.950 421.950 811.050 424.050 ;
        RECT 805.950 406.950 808.050 409.050 ;
        RECT 799.950 394.950 802.050 397.050 ;
        RECT 809.400 391.050 810.600 421.950 ;
        RECT 812.400 409.050 813.600 466.950 ;
        RECT 815.400 451.200 816.600 487.950 ;
        RECT 818.400 487.050 819.600 494.400 ;
        RECT 817.950 484.950 820.050 487.050 ;
        RECT 817.950 460.950 820.050 463.050 ;
        RECT 818.400 454.050 819.600 460.950 ;
        RECT 821.400 457.050 822.600 505.950 ;
        RECT 824.400 496.050 825.600 520.950 ;
        RECT 827.400 517.050 828.600 563.400 ;
        RECT 829.950 532.950 832.050 535.050 ;
        RECT 826.950 514.950 829.050 517.050 ;
        RECT 830.400 496.200 831.600 532.950 ;
        RECT 833.400 520.050 834.600 565.950 ;
        RECT 835.950 562.950 838.050 565.050 ;
        RECT 838.950 562.950 841.050 567.000 ;
        RECT 836.400 556.050 837.600 562.950 ;
        RECT 845.400 556.050 846.600 568.950 ;
        RECT 847.950 565.950 850.050 568.050 ;
        RECT 848.400 559.050 849.600 565.950 ;
        RECT 847.950 556.950 850.050 559.050 ;
        RECT 835.950 553.950 838.050 556.050 ;
        RECT 844.950 553.950 847.050 556.050 ;
        RECT 836.400 529.050 837.600 553.950 ;
        RECT 851.400 550.050 852.600 577.950 ;
        RECT 850.950 547.950 853.050 550.050 ;
        RECT 854.400 547.050 855.600 595.800 ;
        RECT 857.400 574.050 858.600 604.950 ;
        RECT 860.400 598.050 861.600 613.950 ;
        RECT 863.400 607.050 864.600 640.950 ;
        RECT 869.400 631.050 870.600 646.950 ;
        RECT 871.950 643.950 874.050 646.050 ;
        RECT 868.950 628.950 871.050 631.050 ;
        RECT 872.400 622.050 873.600 643.950 ;
        RECT 875.400 631.050 876.600 650.100 ;
        RECT 884.400 649.050 885.600 650.100 ;
        RECT 890.400 649.050 891.600 673.950 ;
        RECT 893.400 652.050 894.600 676.950 ;
        RECT 892.950 649.950 895.050 652.050 ;
        RECT 880.950 646.950 883.050 649.050 ;
        RECT 883.950 646.950 886.050 649.050 ;
        RECT 886.950 646.950 889.050 649.050 ;
        RECT 889.950 646.950 892.050 649.050 ;
        RECT 881.400 645.000 882.600 646.950 ;
        RECT 887.400 645.900 888.600 646.950 ;
        RECT 880.950 640.950 883.050 645.000 ;
        RECT 886.950 643.800 889.050 645.900 ;
        RECT 892.950 643.950 895.050 646.050 ;
        RECT 883.950 637.950 886.050 640.050 ;
        RECT 877.950 631.950 880.050 634.050 ;
        RECT 874.950 628.950 877.050 631.050 ;
        RECT 871.950 619.950 874.050 622.050 ;
        RECT 874.950 613.950 877.050 616.050 ;
        RECT 862.950 604.950 865.050 607.050 ;
        RECT 868.950 606.000 871.050 610.050 ;
        RECT 869.400 604.050 870.600 606.000 ;
        RECT 875.400 604.050 876.600 613.950 ;
        RECT 878.400 607.050 879.600 631.950 ;
        RECT 880.950 628.950 883.050 631.050 ;
        RECT 877.950 604.950 880.050 607.050 ;
        RECT 865.950 601.950 868.050 604.050 ;
        RECT 868.950 601.950 871.050 604.050 ;
        RECT 871.950 601.950 874.050 604.050 ;
        RECT 874.950 601.950 877.050 604.050 ;
        RECT 859.950 595.950 862.050 598.050 ;
        RECT 866.400 597.600 867.600 601.950 ;
        RECT 872.400 600.900 873.600 601.950 ;
        RECT 871.950 598.800 874.050 600.900 ;
        RECT 877.950 598.950 880.050 601.050 ;
        RECT 866.400 596.400 870.600 597.600 ;
        RECT 865.950 592.950 868.050 595.050 ;
        RECT 862.950 583.950 865.050 586.050 ;
        RECT 856.950 571.950 859.050 574.050 ;
        RECT 863.400 571.050 864.600 583.950 ;
        RECT 866.400 583.050 867.600 592.950 ;
        RECT 869.400 586.050 870.600 596.400 ;
        RECT 872.400 595.050 873.600 598.800 ;
        RECT 871.950 592.950 874.050 595.050 ;
        RECT 868.950 583.950 871.050 586.050 ;
        RECT 865.950 580.950 868.050 583.050 ;
        RECT 868.950 573.000 871.050 577.050 ;
        RECT 869.400 571.050 870.600 573.000 ;
        RECT 859.950 568.950 862.050 571.050 ;
        RECT 862.950 568.950 865.050 571.050 ;
        RECT 865.950 568.950 868.050 571.050 ;
        RECT 868.950 568.950 871.050 571.050 ;
        RECT 860.400 567.000 861.600 568.950 ;
        RECT 859.950 562.950 862.050 567.000 ;
        RECT 866.400 559.050 867.600 568.950 ;
        RECT 865.950 556.950 868.050 559.050 ;
        RECT 874.950 556.950 877.050 559.050 ;
        RECT 853.950 544.950 856.050 547.050 ;
        RECT 847.950 532.950 850.050 535.050 ;
        RECT 862.950 532.950 865.050 535.050 ;
        RECT 835.950 526.950 838.050 529.050 ;
        RECT 841.950 527.100 844.050 529.200 ;
        RECT 842.400 526.050 843.600 527.100 ;
        RECT 848.400 526.050 849.600 532.950 ;
        RECT 853.950 527.100 856.050 529.200 ;
        RECT 838.950 523.950 841.050 526.050 ;
        RECT 841.950 523.950 844.050 526.050 ;
        RECT 844.950 523.950 847.050 526.050 ;
        RECT 847.950 523.950 850.050 526.050 ;
        RECT 835.950 520.950 838.050 523.050 ;
        RECT 832.950 517.950 835.050 520.050 ;
        RECT 836.400 508.050 837.600 520.950 ;
        RECT 839.400 517.050 840.600 523.950 ;
        RECT 841.950 517.950 844.050 520.050 ;
        RECT 838.950 514.950 841.050 517.050 ;
        RECT 835.950 505.950 838.050 508.050 ;
        RECT 832.950 502.950 835.050 505.050 ;
        RECT 833.400 499.050 834.600 502.950 ;
        RECT 832.950 496.950 835.050 499.050 ;
        RECT 823.950 493.950 826.050 496.050 ;
        RECT 829.950 494.100 832.050 496.200 ;
        RECT 830.400 493.050 831.600 494.100 ;
        RECT 838.950 493.950 841.050 496.050 ;
        RECT 826.950 490.950 829.050 493.050 ;
        RECT 829.950 490.950 832.050 493.050 ;
        RECT 832.950 490.950 835.050 493.050 ;
        RECT 823.950 487.950 826.050 490.050 ;
        RECT 827.400 489.000 828.600 490.950 ;
        RECT 824.400 460.050 825.600 487.950 ;
        RECT 826.950 484.950 829.050 489.000 ;
        RECT 833.400 484.050 834.600 490.950 ;
        RECT 835.950 487.950 838.050 490.050 ;
        RECT 832.950 481.950 835.050 484.050 ;
        RECT 829.950 475.950 832.050 478.050 ;
        RECT 830.400 466.050 831.600 475.950 ;
        RECT 829.950 463.950 832.050 466.050 ;
        RECT 823.950 457.950 826.050 460.050 ;
        RECT 832.950 457.950 835.050 460.050 ;
        RECT 820.800 454.950 822.900 457.050 ;
        RECT 823.950 454.800 826.050 456.900 ;
        RECT 817.950 451.950 820.050 454.050 ;
        RECT 824.400 451.200 825.600 454.800 ;
        RECT 814.950 449.100 817.050 451.200 ;
        RECT 823.950 449.100 826.050 451.200 ;
        RECT 829.950 449.100 832.050 451.200 ;
        RECT 833.400 451.050 834.600 457.950 ;
        RECT 824.400 448.050 825.600 449.100 ;
        RECT 830.400 448.050 831.600 449.100 ;
        RECT 832.950 448.950 835.050 451.050 ;
        RECT 820.950 445.950 823.050 448.050 ;
        RECT 823.950 445.950 826.050 448.050 ;
        RECT 826.950 445.950 829.050 448.050 ;
        RECT 829.950 445.950 832.050 448.050 ;
        RECT 814.950 439.950 817.050 445.050 ;
        RECT 821.400 436.050 822.600 445.950 ;
        RECT 820.950 433.950 823.050 436.050 ;
        RECT 827.400 427.050 828.600 445.950 ;
        RECT 832.950 442.950 835.050 445.050 ;
        RECT 833.400 436.050 834.600 442.950 ;
        RECT 836.400 436.050 837.600 487.950 ;
        RECT 839.400 478.050 840.600 493.950 ;
        RECT 838.950 475.950 841.050 478.050 ;
        RECT 839.400 451.200 840.600 475.950 ;
        RECT 842.400 472.050 843.600 517.950 ;
        RECT 845.400 484.050 846.600 523.950 ;
        RECT 854.400 520.050 855.600 527.100 ;
        RECT 863.400 526.050 864.600 532.950 ;
        RECT 868.950 527.100 871.050 529.200 ;
        RECT 869.400 526.050 870.600 527.100 ;
        RECT 859.950 523.950 862.050 526.050 ;
        RECT 862.950 523.950 865.050 526.050 ;
        RECT 865.950 523.950 868.050 526.050 ;
        RECT 868.950 523.950 871.050 526.050 ;
        RECT 860.400 522.000 861.600 523.950 ;
        RECT 859.950 520.050 862.050 522.000 ;
        RECT 853.950 517.950 856.050 520.050 ;
        RECT 859.800 519.000 862.050 520.050 ;
        RECT 859.800 517.950 861.900 519.000 ;
        RECT 862.950 517.950 865.050 520.050 ;
        RECT 847.950 505.950 850.050 508.050 ;
        RECT 848.400 496.050 849.600 505.950 ;
        RECT 853.950 502.950 856.050 505.050 ;
        RECT 854.400 499.050 855.600 502.950 ;
        RECT 853.950 496.950 856.050 499.050 ;
        RECT 847.950 493.950 850.050 496.050 ;
        RECT 854.400 493.050 855.600 496.950 ;
        RECT 859.800 494.100 861.900 496.200 ;
        RECT 863.400 496.050 864.600 517.950 ;
        RECT 866.400 501.600 867.600 523.950 ;
        RECT 875.400 522.600 876.600 556.950 ;
        RECT 878.400 541.050 879.600 598.950 ;
        RECT 881.400 598.050 882.600 628.950 ;
        RECT 880.950 595.950 883.050 598.050 ;
        RECT 884.400 592.050 885.600 637.950 ;
        RECT 887.400 616.050 888.600 643.800 ;
        RECT 893.400 640.050 894.600 643.950 ;
        RECT 892.950 637.950 895.050 640.050 ;
        RECT 886.950 613.950 889.050 616.050 ;
        RECT 886.950 609.600 891.000 610.050 ;
        RECT 886.950 607.950 891.600 609.600 ;
        RECT 890.400 604.050 891.600 607.950 ;
        RECT 889.950 601.950 892.050 604.050 ;
        RECT 892.950 601.950 895.050 604.050 ;
        RECT 893.400 600.600 894.600 601.950 ;
        RECT 893.400 599.400 897.600 600.600 ;
        RECT 896.400 598.050 897.600 599.400 ;
        RECT 895.950 595.950 898.050 598.050 ;
        RECT 883.950 589.950 886.050 592.050 ;
        RECT 892.950 589.950 895.050 592.050 ;
        RECT 889.950 583.950 892.050 586.050 ;
        RECT 880.950 562.950 883.050 565.050 ;
        RECT 877.950 538.950 880.050 541.050 ;
        RECT 877.950 532.950 880.050 535.050 ;
        RECT 872.400 521.400 876.600 522.600 ;
        RECT 872.400 505.050 873.600 521.400 ;
        RECT 878.400 508.050 879.600 532.950 ;
        RECT 877.950 505.950 880.050 508.050 ;
        RECT 871.950 502.950 874.050 505.050 ;
        RECT 866.400 500.400 870.600 501.600 ;
        RECT 865.950 496.950 868.050 499.050 ;
        RECT 860.400 493.050 861.600 494.100 ;
        RECT 862.950 493.950 865.050 496.050 ;
        RECT 850.950 490.950 853.050 493.050 ;
        RECT 853.950 490.950 856.050 493.050 ;
        RECT 856.950 490.950 859.050 493.050 ;
        RECT 859.950 490.950 862.050 493.050 ;
        RECT 844.950 481.950 847.050 484.050 ;
        RECT 841.950 469.950 844.050 472.050 ;
        RECT 851.400 466.050 852.600 490.950 ;
        RECT 853.950 484.950 856.050 487.050 ;
        RECT 844.950 463.950 847.050 466.050 ;
        RECT 850.950 463.950 853.050 466.050 ;
        RECT 838.950 449.100 841.050 451.200 ;
        RECT 845.400 451.050 846.600 463.950 ;
        RECT 847.950 460.950 850.050 463.050 ;
        RECT 841.950 448.950 844.050 451.050 ;
        RECT 844.950 448.950 847.050 451.050 ;
        RECT 832.800 433.950 834.900 436.050 ;
        RECT 835.950 433.950 838.050 436.050 ;
        RECT 826.950 424.950 829.050 427.050 ;
        RECT 838.950 424.950 841.050 427.050 ;
        RECT 814.950 421.950 817.050 424.050 ;
        RECT 815.400 418.050 816.600 421.950 ;
        RECT 814.950 415.950 817.050 418.050 ;
        RECT 820.950 416.100 823.050 418.200 ;
        RECT 826.950 417.000 829.050 421.050 ;
        RECT 821.400 415.050 822.600 416.100 ;
        RECT 827.400 415.050 828.600 417.000 ;
        RECT 832.950 415.950 835.050 418.050 ;
        RECT 817.950 412.950 820.050 415.050 ;
        RECT 820.950 412.950 823.050 415.050 ;
        RECT 823.950 412.950 826.050 415.050 ;
        RECT 826.950 412.950 829.050 415.050 ;
        RECT 814.950 409.950 817.050 412.050 ;
        RECT 818.400 411.000 819.600 412.950 ;
        RECT 824.400 411.000 825.600 412.950 ;
        RECT 811.950 406.950 814.050 409.050 ;
        RECT 811.950 400.950 814.050 403.050 ;
        RECT 808.950 388.950 811.050 391.050 ;
        RECT 809.400 376.050 810.600 388.950 ;
        RECT 808.950 373.950 811.050 376.050 ;
        RECT 796.950 371.100 799.050 373.200 ;
        RECT 802.950 371.100 805.050 373.200 ;
        RECT 797.400 370.050 798.600 371.100 ;
        RECT 803.400 370.050 804.600 371.100 ;
        RECT 787.950 367.950 790.050 370.050 ;
        RECT 796.950 367.950 799.050 370.050 ;
        RECT 799.950 367.950 802.050 370.050 ;
        RECT 802.950 367.950 805.050 370.050 ;
        RECT 805.950 367.950 808.050 370.050 ;
        RECT 793.950 364.950 796.050 367.050 ;
        RECT 787.950 346.950 790.050 349.050 ;
        RECT 788.400 340.050 789.600 346.950 ;
        RECT 794.400 343.200 795.600 364.950 ;
        RECT 800.400 345.600 801.600 367.950 ;
        RECT 806.400 366.000 807.600 367.950 ;
        RECT 805.950 361.950 808.050 366.000 ;
        RECT 808.950 364.950 811.050 367.050 ;
        RECT 800.400 344.400 804.600 345.600 ;
        RECT 793.950 341.100 796.050 343.200 ;
        RECT 787.950 337.950 790.050 340.050 ;
        RECT 793.950 337.950 796.050 340.050 ;
        RECT 799.950 339.000 802.050 343.050 ;
        RECT 803.400 340.050 804.600 344.400 ;
        RECT 805.950 343.950 808.050 346.050 ;
        RECT 794.400 337.050 795.600 337.950 ;
        RECT 800.400 337.050 801.600 339.000 ;
        RECT 802.950 337.950 805.050 340.050 ;
        RECT 790.950 334.950 793.050 337.050 ;
        RECT 793.950 334.950 796.050 337.050 ;
        RECT 796.950 334.950 799.050 337.050 ;
        RECT 799.950 334.950 802.050 337.050 ;
        RECT 791.400 333.900 792.600 334.950 ;
        RECT 797.400 333.900 798.600 334.950 ;
        RECT 790.950 331.800 793.050 333.900 ;
        RECT 796.950 331.800 799.050 333.900 ;
        RECT 802.950 331.950 805.050 334.050 ;
        RECT 803.400 325.050 804.600 331.950 ;
        RECT 802.950 322.950 805.050 325.050 ;
        RECT 799.950 319.950 802.050 322.050 ;
        RECT 790.950 301.950 793.050 304.050 ;
        RECT 784.950 295.950 787.050 298.050 ;
        RECT 785.400 292.050 786.600 295.950 ;
        RECT 791.400 292.050 792.600 301.950 ;
        RECT 784.950 289.950 787.050 292.050 ;
        RECT 787.950 289.950 790.050 292.050 ;
        RECT 790.950 289.950 793.050 292.050 ;
        RECT 793.950 289.950 796.050 292.050 ;
        RECT 788.400 288.900 789.600 289.950 ;
        RECT 787.950 286.800 790.050 288.900 ;
        RECT 788.400 265.050 789.600 286.800 ;
        RECT 790.950 283.950 793.050 286.050 ;
        RECT 791.400 268.050 792.600 283.950 ;
        RECT 794.400 283.050 795.600 289.950 ;
        RECT 800.400 286.050 801.600 319.950 ;
        RECT 806.400 304.050 807.600 343.950 ;
        RECT 805.950 301.950 808.050 304.050 ;
        RECT 809.400 301.050 810.600 364.950 ;
        RECT 812.400 316.050 813.600 400.950 ;
        RECT 815.400 376.050 816.600 409.950 ;
        RECT 817.950 406.950 820.050 411.000 ;
        RECT 823.950 406.950 826.050 411.000 ;
        RECT 823.950 394.950 826.050 397.050 ;
        RECT 814.950 373.950 817.050 376.050 ;
        RECT 817.950 372.000 820.050 376.050 ;
        RECT 818.400 370.050 819.600 372.000 ;
        RECT 824.400 370.050 825.600 394.950 ;
        RECT 829.950 385.950 832.050 388.050 ;
        RECT 817.950 367.950 820.050 370.050 ;
        RECT 820.950 367.950 823.050 370.050 ;
        RECT 823.950 367.950 826.050 370.050 ;
        RECT 814.950 364.950 817.050 367.050 ;
        RECT 815.400 340.050 816.600 364.950 ;
        RECT 821.400 349.050 822.600 367.950 ;
        RECT 830.400 354.600 831.600 385.950 ;
        RECT 833.400 382.050 834.600 415.950 ;
        RECT 839.400 415.050 840.600 424.950 ;
        RECT 842.400 424.050 843.600 448.950 ;
        RECT 848.400 448.050 849.600 460.950 ;
        RECT 850.950 457.950 853.050 460.050 ;
        RECT 851.400 454.050 852.600 457.950 ;
        RECT 854.400 457.050 855.600 484.950 ;
        RECT 857.400 460.050 858.600 490.950 ;
        RECT 866.400 484.050 867.600 496.950 ;
        RECT 869.400 496.050 870.600 500.400 ;
        RECT 868.950 493.950 871.050 496.050 ;
        RECT 874.950 495.000 877.050 499.050 ;
        RECT 881.400 496.200 882.600 562.950 ;
        RECT 883.950 547.950 886.050 550.050 ;
        RECT 875.400 493.050 876.600 495.000 ;
        RECT 880.950 494.100 883.050 496.200 ;
        RECT 884.400 496.050 885.600 547.950 ;
        RECT 881.400 493.050 882.600 494.100 ;
        RECT 883.950 493.950 886.050 496.050 ;
        RECT 886.950 493.950 889.050 496.050 ;
        RECT 871.950 490.950 874.050 493.050 ;
        RECT 874.950 490.950 877.050 493.050 ;
        RECT 877.950 490.950 880.050 493.050 ;
        RECT 880.950 490.950 883.050 493.050 ;
        RECT 868.950 487.950 871.050 490.050 ;
        RECT 872.400 489.900 873.600 490.950 ;
        RECT 865.950 481.950 868.050 484.050 ;
        RECT 859.950 466.950 862.050 469.050 ;
        RECT 856.950 457.950 859.050 460.050 ;
        RECT 853.950 454.950 856.050 457.050 ;
        RECT 850.950 451.950 853.050 454.050 ;
        RECT 854.400 451.050 855.600 454.950 ;
        RECT 857.400 454.050 858.600 457.950 ;
        RECT 856.950 451.950 859.050 454.050 ;
        RECT 853.950 448.950 856.050 451.050 ;
        RECT 847.950 445.950 850.050 448.050 ;
        RECT 850.950 445.950 853.050 448.050 ;
        RECT 851.400 444.900 852.600 445.950 ;
        RECT 850.950 442.800 853.050 444.900 ;
        RECT 844.950 427.950 847.050 430.050 ;
        RECT 853.950 427.950 856.050 430.050 ;
        RECT 841.950 421.950 844.050 424.050 ;
        RECT 845.400 415.050 846.600 427.950 ;
        RECT 850.950 421.950 853.050 424.050 ;
        RECT 838.950 412.950 841.050 415.050 ;
        RECT 841.950 412.950 844.050 415.050 ;
        RECT 844.950 412.950 847.050 415.050 ;
        RECT 832.950 379.950 835.050 382.050 ;
        RECT 842.400 379.050 843.600 412.950 ;
        RECT 832.950 376.800 835.050 378.900 ;
        RECT 841.950 376.950 844.050 379.050 ;
        RECT 833.400 364.050 834.600 376.800 ;
        RECT 847.950 373.200 850.050 376.050 ;
        RECT 841.950 371.100 844.050 373.200 ;
        RECT 847.800 372.000 850.050 373.200 ;
        RECT 851.400 373.050 852.600 421.950 ;
        RECT 854.400 403.050 855.600 427.950 ;
        RECT 857.400 421.050 858.600 451.950 ;
        RECT 860.400 451.050 861.600 466.950 ;
        RECT 866.400 451.200 867.600 481.950 ;
        RECT 859.950 448.950 862.050 451.050 ;
        RECT 865.950 449.100 868.050 451.200 ;
        RECT 869.400 450.600 870.600 487.950 ;
        RECT 871.950 487.800 874.050 489.900 ;
        RECT 872.400 463.050 873.600 487.800 ;
        RECT 878.400 486.600 879.600 490.950 ;
        RECT 883.950 487.950 886.050 490.050 ;
        RECT 875.400 485.400 879.600 486.600 ;
        RECT 875.400 478.050 876.600 485.400 ;
        RECT 874.950 475.950 877.050 478.050 ;
        RECT 874.950 463.950 877.050 466.050 ;
        RECT 871.950 460.950 874.050 463.050 ;
        RECT 869.400 449.400 873.600 450.600 ;
        RECT 866.400 448.050 867.600 449.100 ;
        RECT 862.950 445.950 865.050 448.050 ;
        RECT 865.950 445.950 868.050 448.050 ;
        RECT 859.950 442.950 862.050 445.050 ;
        RECT 863.400 444.000 864.600 445.950 ;
        RECT 860.400 424.050 861.600 442.950 ;
        RECT 862.950 439.950 865.050 444.000 ;
        RECT 872.400 438.600 873.600 449.400 ;
        RECT 875.400 441.600 876.600 463.950 ;
        RECT 880.950 460.950 883.050 463.050 ;
        RECT 881.400 448.050 882.600 460.950 ;
        RECT 884.400 454.050 885.600 487.950 ;
        RECT 887.400 469.050 888.600 493.950 ;
        RECT 886.950 466.950 889.050 469.050 ;
        RECT 890.400 466.050 891.600 583.950 ;
        RECT 889.950 463.950 892.050 466.050 ;
        RECT 883.950 451.950 886.050 454.050 ;
        RECT 886.950 450.000 889.050 454.050 ;
        RECT 893.400 451.050 894.600 589.950 ;
        RECT 896.400 529.050 897.600 595.950 ;
        RECT 895.950 526.950 898.050 529.050 ;
        RECT 895.950 469.950 898.050 472.050 ;
        RECT 887.400 448.050 888.600 450.000 ;
        RECT 892.950 448.950 895.050 451.050 ;
        RECT 880.950 445.950 883.050 448.050 ;
        RECT 883.950 445.950 886.050 448.050 ;
        RECT 886.950 445.950 889.050 448.050 ;
        RECT 889.950 445.950 892.050 448.050 ;
        RECT 884.400 444.900 885.600 445.950 ;
        RECT 883.950 442.800 886.050 444.900 ;
        RECT 875.400 440.400 879.600 441.600 ;
        RECT 869.400 437.400 873.600 438.600 ;
        RECT 859.950 421.950 862.050 424.050 ;
        RECT 869.400 421.050 870.600 437.400 ;
        RECT 874.950 436.950 877.050 439.050 ;
        RECT 871.950 433.950 874.050 436.050 ;
        RECT 856.950 418.950 859.050 421.050 ;
        RECT 868.950 418.950 871.050 421.050 ;
        RECT 857.400 417.600 858.600 418.950 ;
        RECT 857.400 416.400 861.600 417.600 ;
        RECT 860.400 415.050 861.600 416.400 ;
        RECT 865.950 416.100 868.050 418.200 ;
        RECT 872.400 418.050 873.600 433.950 ;
        RECT 866.400 415.050 867.600 416.100 ;
        RECT 871.950 415.950 874.050 418.050 ;
        RECT 859.950 412.950 862.050 415.050 ;
        RECT 862.950 412.950 865.050 415.050 ;
        RECT 865.950 412.950 868.050 415.050 ;
        RECT 868.950 412.950 871.050 415.050 ;
        RECT 863.400 411.000 864.600 412.950 ;
        RECT 862.950 406.950 865.050 411.000 ;
        RECT 853.950 400.950 856.050 403.050 ;
        RECT 869.400 394.050 870.600 412.950 ;
        RECT 875.400 406.050 876.600 436.950 ;
        RECT 874.950 403.950 877.050 406.050 ;
        RECT 868.950 391.950 871.050 394.050 ;
        RECT 862.950 379.950 865.050 382.050 ;
        RECT 847.800 371.100 849.900 372.000 ;
        RECT 842.400 370.050 843.600 371.100 ;
        RECT 848.400 370.050 849.600 371.100 ;
        RECT 850.950 370.950 853.050 373.050 ;
        RECT 856.950 370.950 859.050 373.050 ;
        RECT 838.950 367.950 841.050 370.050 ;
        RECT 841.950 367.950 844.050 370.050 ;
        RECT 844.950 367.950 847.050 370.050 ;
        RECT 847.950 367.950 850.050 370.050 ;
        RECT 835.950 364.950 838.050 367.050 ;
        RECT 839.400 366.000 840.600 367.950 ;
        RECT 832.950 361.950 835.050 364.050 ;
        RECT 836.400 358.050 837.600 364.950 ;
        RECT 838.950 361.950 841.050 366.000 ;
        RECT 835.950 355.950 838.050 358.050 ;
        RECT 830.400 353.400 834.600 354.600 ;
        RECT 820.950 346.950 823.050 349.050 ;
        RECT 820.950 343.800 823.050 345.900 ;
        RECT 814.950 337.950 817.050 340.050 ;
        RECT 821.400 337.050 822.600 343.800 ;
        RECT 826.950 339.000 829.050 343.050 ;
        RECT 827.400 337.050 828.600 339.000 ;
        RECT 817.950 334.950 820.050 337.050 ;
        RECT 820.950 334.950 823.050 337.050 ;
        RECT 823.950 334.950 826.050 337.050 ;
        RECT 826.950 334.950 829.050 337.050 ;
        RECT 818.400 319.050 819.600 334.950 ;
        RECT 824.400 333.900 825.600 334.950 ;
        RECT 823.950 331.800 826.050 333.900 ;
        RECT 820.950 328.950 823.050 331.050 ;
        RECT 817.950 316.950 820.050 319.050 ;
        RECT 811.950 313.950 814.050 316.050 ;
        RECT 808.950 298.950 811.050 301.050 ;
        RECT 817.950 298.950 820.050 301.050 ;
        RECT 802.950 295.950 805.050 298.050 ;
        RECT 799.950 283.950 802.050 286.050 ;
        RECT 793.950 280.950 796.050 283.050 ;
        RECT 790.950 265.950 793.050 268.050 ;
        RECT 781.950 262.950 784.050 265.050 ;
        RECT 787.950 262.950 790.050 265.050 ;
        RECT 794.400 264.600 795.600 280.950 ;
        RECT 799.950 277.950 802.050 280.050 ;
        RECT 796.950 268.950 799.050 271.050 ;
        RECT 791.400 263.400 795.600 264.600 ;
        RECT 773.400 259.050 774.600 261.000 ;
        RECT 778.950 259.950 781.050 262.050 ;
        RECT 769.950 256.950 772.050 259.050 ;
        RECT 772.950 256.950 775.050 259.050 ;
        RECT 775.950 256.950 778.050 259.050 ;
        RECT 770.400 255.900 771.600 256.950 ;
        RECT 763.950 253.800 766.050 255.900 ;
        RECT 769.950 253.800 772.050 255.900 ;
        RECT 776.400 255.000 777.600 256.950 ;
        RECT 769.950 250.650 772.050 252.750 ;
        RECT 775.950 250.950 778.050 255.000 ;
        RECT 778.950 253.950 781.050 256.050 ;
        RECT 766.950 235.950 769.050 238.050 ;
        RECT 767.400 226.050 768.600 235.950 ;
        RECT 766.950 223.950 769.050 226.050 ;
        RECT 770.400 223.050 771.600 250.650 ;
        RECT 779.400 249.600 780.600 253.950 ;
        RECT 782.400 253.050 783.600 262.950 ;
        RECT 791.400 259.050 792.600 263.400 ;
        RECT 797.400 259.050 798.600 268.950 ;
        RECT 800.400 268.050 801.600 277.950 ;
        RECT 799.950 265.950 802.050 268.050 ;
        RECT 787.950 256.950 790.050 259.050 ;
        RECT 790.950 256.950 793.050 259.050 ;
        RECT 793.950 256.950 796.050 259.050 ;
        RECT 796.950 256.950 799.050 259.050 ;
        RECT 788.400 255.900 789.600 256.950 ;
        RECT 787.950 253.800 790.050 255.900 ;
        RECT 794.400 255.000 795.600 256.950 ;
        RECT 781.950 250.950 784.050 253.050 ;
        RECT 793.950 250.950 796.050 255.000 ;
        RECT 799.950 253.950 802.050 256.050 ;
        RECT 796.950 250.950 799.050 253.050 ;
        RECT 776.400 248.400 780.600 249.600 ;
        RECT 769.950 220.950 772.050 223.050 ;
        RECT 760.950 218.100 763.050 220.200 ;
        RECT 760.950 214.950 763.050 217.050 ;
        RECT 766.950 216.000 769.050 220.050 ;
        RECT 770.400 217.050 771.600 220.950 ;
        RECT 772.950 217.950 775.050 220.050 ;
        RECT 761.400 214.050 762.600 214.950 ;
        RECT 767.400 214.050 768.600 216.000 ;
        RECT 769.950 214.950 772.050 217.050 ;
        RECT 757.950 211.950 760.050 214.050 ;
        RECT 760.950 211.950 763.050 214.050 ;
        RECT 763.950 211.950 766.050 214.050 ;
        RECT 766.950 211.950 769.050 214.050 ;
        RECT 758.400 211.050 759.600 211.950 ;
        RECT 754.950 209.400 759.600 211.050 ;
        RECT 764.400 210.900 765.600 211.950 ;
        RECT 754.950 208.950 759.000 209.400 ;
        RECT 763.950 208.800 766.050 210.900 ;
        RECT 757.950 205.950 763.050 208.050 ;
        RECT 769.950 205.950 772.050 211.050 ;
        RECT 769.950 199.950 772.050 202.050 ;
        RECT 752.400 182.400 756.600 183.600 ;
        RECT 739.950 178.950 742.050 181.050 ;
        RECT 742.950 178.950 745.050 181.050 ;
        RECT 745.950 178.950 748.050 181.050 ;
        RECT 748.950 178.950 751.050 181.050 ;
        RECT 736.950 175.950 739.050 178.050 ;
        RECT 743.400 177.900 744.600 178.950 ;
        RECT 733.950 154.950 736.050 157.050 ;
        RECT 725.400 103.050 726.600 104.100 ;
        RECT 730.950 103.950 733.050 106.050 ;
        RECT 721.950 100.950 724.050 103.050 ;
        RECT 724.950 100.950 727.050 103.050 ;
        RECT 727.950 100.950 730.050 103.050 ;
        RECT 709.950 91.950 712.050 94.050 ;
        RECT 715.950 91.950 718.050 94.050 ;
        RECT 722.400 91.050 723.600 100.950 ;
        RECT 728.400 99.900 729.600 100.950 ;
        RECT 727.950 97.800 730.050 99.900 ;
        RECT 730.950 97.950 733.050 100.050 ;
        RECT 721.950 88.950 724.050 91.050 ;
        RECT 691.950 85.950 694.050 88.050 ;
        RECT 703.950 85.950 706.050 88.050 ;
        RECT 688.950 76.950 691.050 79.050 ;
        RECT 683.400 59.400 687.600 60.600 ;
        RECT 664.950 55.950 667.050 58.050 ;
        RECT 667.950 55.950 670.050 58.050 ;
        RECT 670.950 55.950 673.050 58.050 ;
        RECT 673.950 55.950 676.050 58.050 ;
        RECT 616.950 26.100 619.050 28.200 ;
        RECT 607.950 22.950 610.050 25.050 ;
        RECT 610.950 22.950 613.050 25.050 ;
        RECT 613.950 22.950 616.050 25.050 ;
        RECT 608.400 16.050 609.600 22.950 ;
        RECT 614.400 21.900 615.600 22.950 ;
        RECT 620.400 21.900 621.600 52.950 ;
        RECT 628.950 52.800 631.050 54.900 ;
        RECT 640.950 52.800 643.050 54.900 ;
        RECT 646.950 52.800 649.050 54.900 ;
        RECT 652.950 52.800 655.050 54.900 ;
        RECT 625.950 26.100 628.050 28.200 ;
        RECT 631.950 26.100 634.050 28.200 ;
        RECT 641.400 27.600 642.600 52.800 ;
        RECT 665.400 40.050 666.600 55.950 ;
        RECT 671.400 46.050 672.600 55.950 ;
        RECT 680.400 55.050 681.600 59.100 ;
        RECT 679.950 52.950 682.050 55.050 ;
        RECT 670.950 43.950 673.050 46.050 ;
        RECT 664.950 37.950 667.050 40.050 ;
        RECT 646.950 32.400 649.050 34.500 ;
        RECT 667.950 32.400 670.050 34.500 ;
        RECT 683.400 34.050 684.600 59.400 ;
        RECT 692.400 58.050 693.600 85.950 ;
        RECT 718.950 79.950 721.050 82.050 ;
        RECT 712.950 64.950 715.050 67.050 ;
        RECT 697.950 60.000 700.050 64.050 ;
        RECT 698.400 58.050 699.600 60.000 ;
        RECT 703.950 58.950 706.050 64.050 ;
        RECT 688.950 55.950 691.050 58.050 ;
        RECT 691.950 55.950 694.050 58.050 ;
        RECT 694.950 55.950 697.050 58.050 ;
        RECT 697.950 55.950 700.050 58.050 ;
        RECT 689.400 54.900 690.600 55.950 ;
        RECT 695.400 54.900 696.600 55.950 ;
        RECT 688.950 52.800 691.050 54.900 ;
        RECT 694.950 52.800 697.050 54.900 ;
        RECT 700.950 52.950 703.050 55.050 ;
        RECT 691.950 43.950 694.050 46.050 ;
        RECT 641.400 26.400 645.600 27.600 ;
        RECT 626.400 25.050 627.600 26.100 ;
        RECT 632.400 25.050 633.600 26.100 ;
        RECT 644.400 25.050 645.600 26.400 ;
        RECT 625.950 22.950 628.050 25.050 ;
        RECT 628.950 22.950 631.050 25.050 ;
        RECT 631.950 22.950 634.050 25.050 ;
        RECT 634.950 22.950 637.050 25.050 ;
        RECT 643.950 22.950 646.050 25.050 ;
        RECT 613.950 19.800 616.050 21.900 ;
        RECT 619.950 19.800 622.050 21.900 ;
        RECT 622.950 19.950 625.050 22.050 ;
        RECT 629.400 21.900 630.600 22.950 ;
        RECT 623.400 16.050 624.600 19.950 ;
        RECT 628.950 19.800 631.050 21.900 ;
        RECT 635.400 16.050 636.600 22.950 ;
        RECT 647.850 17.400 649.050 32.400 ;
        RECT 652.950 26.100 655.050 28.200 ;
        RECT 653.400 22.050 654.600 26.100 ;
        RECT 661.950 22.950 664.050 25.050 ;
        RECT 652.950 19.950 655.050 22.050 ;
        RECT 662.400 21.600 663.600 22.950 ;
        RECT 661.950 19.500 664.050 21.600 ;
        RECT 607.950 13.950 610.050 16.050 ;
        RECT 622.950 13.950 625.050 16.050 ;
        RECT 634.950 13.950 637.050 16.050 ;
        RECT 646.950 15.300 649.050 17.400 ;
        RECT 647.850 11.700 649.050 15.300 ;
        RECT 668.100 12.600 669.300 32.400 ;
        RECT 682.950 31.950 685.050 34.050 ;
        RECT 683.400 25.050 684.600 31.950 ;
        RECT 692.400 25.050 693.600 43.950 ;
        RECT 670.950 22.950 673.050 25.050 ;
        RECT 682.950 22.950 685.050 25.050 ;
        RECT 688.950 22.950 691.050 25.050 ;
        RECT 691.950 22.950 694.050 25.050 ;
        RECT 694.950 22.950 697.050 25.050 ;
        RECT 671.400 21.600 672.600 22.950 ;
        RECT 689.400 21.900 690.600 22.950 ;
        RECT 695.400 21.900 696.600 22.950 ;
        RECT 701.400 21.900 702.600 52.950 ;
        RECT 670.950 19.500 673.050 21.600 ;
        RECT 688.950 19.800 691.050 21.900 ;
        RECT 694.950 19.800 697.050 21.900 ;
        RECT 700.950 19.800 703.050 21.900 ;
        RECT 704.400 19.050 705.600 58.950 ;
        RECT 713.400 58.050 714.600 64.950 ;
        RECT 709.950 55.950 712.050 58.050 ;
        RECT 712.950 55.950 715.050 58.050 ;
        RECT 710.400 54.900 711.600 55.950 ;
        RECT 719.400 54.900 720.600 79.950 ;
        RECT 731.400 70.050 732.600 97.950 ;
        RECT 734.400 76.050 735.600 154.950 ;
        RECT 737.400 139.050 738.600 175.950 ;
        RECT 742.950 175.800 745.050 177.900 ;
        RECT 749.400 166.050 750.600 178.950 ;
        RECT 748.950 163.950 751.050 166.050 ;
        RECT 751.950 160.950 754.050 163.050 ;
        RECT 736.950 136.950 739.050 139.050 ;
        RECT 742.950 137.100 745.050 139.200 ;
        RECT 748.950 138.000 751.050 142.050 ;
        RECT 752.400 139.050 753.600 160.950 ;
        RECT 743.400 136.050 744.600 137.100 ;
        RECT 749.400 136.050 750.600 138.000 ;
        RECT 751.950 136.950 754.050 139.050 ;
        RECT 739.950 133.950 742.050 136.050 ;
        RECT 742.950 133.950 745.050 136.050 ;
        RECT 745.950 133.950 748.050 136.050 ;
        RECT 748.950 133.950 751.050 136.050 ;
        RECT 740.400 133.050 741.600 133.950 ;
        RECT 736.950 131.400 741.600 133.050 ;
        RECT 736.950 130.950 741.000 131.400 ;
        RECT 736.800 127.800 738.900 129.900 ;
        RECT 739.950 127.950 742.050 130.050 ;
        RECT 737.400 99.900 738.600 127.800 ;
        RECT 736.950 97.800 739.050 99.900 ;
        RECT 733.950 73.950 736.050 76.050 ;
        RECT 730.950 67.950 733.050 70.050 ;
        RECT 737.400 64.050 738.600 97.800 ;
        RECT 740.400 91.050 741.600 127.950 ;
        RECT 746.400 124.050 747.600 133.950 ;
        RECT 745.950 121.950 748.050 124.050 ;
        RECT 755.400 121.050 756.600 182.400 ;
        RECT 757.950 182.100 760.050 184.200 ;
        RECT 763.950 182.100 766.050 184.200 ;
        RECT 770.400 184.050 771.600 199.950 ;
        RECT 758.400 169.050 759.600 182.100 ;
        RECT 764.400 181.050 765.600 182.100 ;
        RECT 769.950 181.950 772.050 184.050 ;
        RECT 763.950 178.950 766.050 181.050 ;
        RECT 766.950 178.950 769.050 181.050 ;
        RECT 757.950 166.950 760.050 169.050 ;
        RECT 758.400 127.050 759.600 166.950 ;
        RECT 760.950 148.950 763.050 151.050 ;
        RECT 757.950 124.950 760.050 127.050 ;
        RECT 754.950 118.950 757.050 121.050 ;
        RECT 752.400 108.900 753.600 111.450 ;
        RECT 748.200 105.900 750.300 107.700 ;
        RECT 752.100 106.800 754.200 108.900 ;
        RECT 755.400 108.300 757.500 110.400 ;
        RECT 761.400 108.600 762.600 148.950 ;
        RECT 767.400 142.050 768.600 178.950 ;
        RECT 769.950 175.950 772.050 178.050 ;
        RECT 770.400 169.050 771.600 175.950 ;
        RECT 769.950 166.950 772.050 169.050 ;
        RECT 769.950 157.950 772.050 160.050 ;
        RECT 766.950 139.950 769.050 142.050 ;
        RECT 770.400 136.050 771.600 157.950 ;
        RECT 773.400 151.050 774.600 217.950 ;
        RECT 776.400 175.050 777.600 248.400 ;
        RECT 793.950 247.800 796.050 249.900 ;
        RECT 794.400 238.050 795.600 247.800 ;
        RECT 797.400 241.050 798.600 250.950 ;
        RECT 796.950 238.950 799.050 241.050 ;
        RECT 793.950 235.950 796.050 238.050 ;
        RECT 796.950 229.950 799.050 232.050 ;
        RECT 787.800 223.950 789.900 226.050 ;
        RECT 790.950 223.950 793.050 226.050 ;
        RECT 781.950 215.100 784.050 217.200 ;
        RECT 788.400 217.050 789.600 223.950 ;
        RECT 782.400 214.050 783.600 215.100 ;
        RECT 787.950 214.950 790.050 217.050 ;
        RECT 781.950 211.950 784.050 214.050 ;
        RECT 784.950 211.950 787.050 214.050 ;
        RECT 785.400 210.900 786.600 211.950 ;
        RECT 784.950 208.800 787.050 210.900 ;
        RECT 785.400 205.050 786.600 208.800 ;
        RECT 784.950 202.950 787.050 205.050 ;
        RECT 791.400 187.200 792.600 223.950 ;
        RECT 797.400 217.200 798.600 229.950 ;
        RECT 800.400 223.050 801.600 253.950 ;
        RECT 803.400 226.050 804.600 295.950 ;
        RECT 805.950 292.950 808.050 295.050 ;
        RECT 814.950 293.100 817.050 295.200 ;
        RECT 818.400 295.050 819.600 298.950 ;
        RECT 806.400 256.050 807.600 292.950 ;
        RECT 815.400 292.050 816.600 293.100 ;
        RECT 817.950 292.950 820.050 295.050 ;
        RECT 811.950 289.950 814.050 292.050 ;
        RECT 814.950 289.950 817.050 292.050 ;
        RECT 812.400 277.050 813.600 289.950 ;
        RECT 817.950 286.800 820.050 288.900 ;
        RECT 811.950 274.950 814.050 277.050 ;
        RECT 818.400 274.050 819.600 286.800 ;
        RECT 808.950 271.950 811.050 274.050 ;
        RECT 817.950 271.950 820.050 274.050 ;
        RECT 805.950 253.950 808.050 256.050 ;
        RECT 805.950 235.950 808.050 238.050 ;
        RECT 806.400 229.050 807.600 235.950 ;
        RECT 805.950 226.950 808.050 229.050 ;
        RECT 802.950 223.950 805.050 226.050 ;
        RECT 799.950 220.950 802.050 223.050 ;
        RECT 800.400 219.600 801.600 220.950 ;
        RECT 800.400 218.400 804.600 219.600 ;
        RECT 796.950 215.100 799.050 217.200 ;
        RECT 797.400 214.050 798.600 215.100 ;
        RECT 803.400 214.050 804.600 218.400 ;
        RECT 796.950 211.950 799.050 214.050 ;
        RECT 799.950 211.950 802.050 214.050 ;
        RECT 802.950 211.950 805.050 214.050 ;
        RECT 793.950 208.950 796.050 211.050 ;
        RECT 784.950 183.000 787.050 187.050 ;
        RECT 790.950 185.100 793.050 187.200 ;
        RECT 794.400 184.050 795.600 208.950 ;
        RECT 800.400 196.050 801.600 211.950 ;
        RECT 809.400 198.600 810.600 271.950 ;
        RECT 821.400 265.050 822.600 328.950 ;
        RECT 829.950 304.950 832.050 307.050 ;
        RECT 823.950 295.950 829.050 298.050 ;
        RECT 830.400 292.050 831.600 304.950 ;
        RECT 833.400 304.050 834.600 353.400 ;
        RECT 835.950 346.950 838.050 349.050 ;
        RECT 836.400 340.050 837.600 346.950 ;
        RECT 845.400 346.050 846.600 367.950 ;
        RECT 844.950 343.950 847.050 346.050 ;
        RECT 835.950 337.950 838.050 340.050 ;
        RECT 838.950 339.000 841.050 343.050 ;
        RECT 839.400 337.050 840.600 339.000 ;
        RECT 844.950 338.100 847.050 340.200 ;
        RECT 845.400 337.050 846.600 338.100 ;
        RECT 853.950 337.950 856.050 340.050 ;
        RECT 838.950 334.950 841.050 337.050 ;
        RECT 841.950 334.950 844.050 337.050 ;
        RECT 844.950 334.950 847.050 337.050 ;
        RECT 847.950 334.950 850.050 337.050 ;
        RECT 842.400 333.900 843.600 334.950 ;
        RECT 841.950 331.800 844.050 333.900 ;
        RECT 848.400 333.000 849.600 334.950 ;
        RECT 847.950 328.950 850.050 333.000 ;
        RECT 854.400 307.050 855.600 337.950 ;
        RECT 853.950 304.950 856.050 307.050 ;
        RECT 832.950 301.950 835.050 304.050 ;
        RECT 847.950 301.950 850.050 304.050 ;
        RECT 835.950 294.000 838.050 298.050 ;
        RECT 836.400 292.050 837.600 294.000 ;
        RECT 844.950 292.950 847.050 295.050 ;
        RECT 829.950 289.950 832.050 292.050 ;
        RECT 832.950 289.950 835.050 292.050 ;
        RECT 835.950 289.950 838.050 292.050 ;
        RECT 838.950 289.950 841.050 292.050 ;
        RECT 823.950 286.950 826.050 289.050 ;
        RECT 826.950 286.950 829.050 289.050 ;
        RECT 811.950 259.950 814.050 265.050 ;
        RECT 820.950 262.950 823.050 265.050 ;
        RECT 817.950 260.100 820.050 262.200 ;
        RECT 818.400 259.050 819.600 260.100 ;
        RECT 824.400 259.050 825.600 286.950 ;
        RECT 827.400 273.600 828.600 286.950 ;
        RECT 833.400 274.050 834.600 289.950 ;
        RECT 839.400 288.900 840.600 289.950 ;
        RECT 838.950 286.800 841.050 288.900 ;
        RECT 838.950 280.950 841.050 283.050 ;
        RECT 827.400 272.400 831.600 273.600 ;
        RECT 826.950 268.950 829.050 271.050 ;
        RECT 830.400 270.600 831.600 272.400 ;
        RECT 832.950 271.950 835.050 274.050 ;
        RECT 830.400 269.400 834.600 270.600 ;
        RECT 827.400 262.050 828.600 268.950 ;
        RECT 829.950 265.950 832.050 268.050 ;
        RECT 826.950 259.950 829.050 262.050 ;
        RECT 814.950 256.950 817.050 259.050 ;
        RECT 817.950 256.950 820.050 259.050 ;
        RECT 820.950 256.950 823.050 259.050 ;
        RECT 823.950 256.950 826.050 259.050 ;
        RECT 815.400 256.050 816.600 256.950 ;
        RECT 811.950 254.400 816.600 256.050 ;
        RECT 811.950 253.950 816.000 254.400 ;
        RECT 814.950 250.950 817.050 253.050 ;
        RECT 811.950 238.950 814.050 241.050 ;
        RECT 806.400 197.400 810.600 198.600 ;
        RECT 799.950 193.950 802.050 196.050 ;
        RECT 796.950 190.950 799.050 193.050 ;
        RECT 785.400 181.050 786.600 183.000 ;
        RECT 790.950 181.950 793.050 184.050 ;
        RECT 793.950 181.950 796.050 184.050 ;
        RECT 791.400 181.050 792.600 181.950 ;
        RECT 781.950 178.950 784.050 181.050 ;
        RECT 784.950 178.950 787.050 181.050 ;
        RECT 787.950 178.950 790.050 181.050 ;
        RECT 790.950 178.950 793.050 181.050 ;
        RECT 775.950 172.950 778.050 175.050 ;
        RECT 778.950 172.950 781.050 178.050 ;
        RECT 782.400 177.900 783.600 178.950 ;
        RECT 781.950 175.800 784.050 177.900 ;
        RECT 781.950 172.650 784.050 174.750 ;
        RECT 775.950 166.950 778.050 169.050 ;
        RECT 772.950 148.950 775.050 151.050 ;
        RECT 776.400 148.050 777.600 166.950 ;
        RECT 778.950 151.950 781.050 154.050 ;
        RECT 775.950 145.950 778.050 148.050 ;
        RECT 775.950 138.000 778.050 142.050 ;
        RECT 779.400 139.050 780.600 151.950 ;
        RECT 776.400 136.050 777.600 138.000 ;
        RECT 778.950 136.950 781.050 139.050 ;
        RECT 766.950 133.950 769.050 136.050 ;
        RECT 769.950 133.950 772.050 136.050 ;
        RECT 772.950 133.950 775.050 136.050 ;
        RECT 775.950 133.950 778.050 136.050 ;
        RECT 763.950 130.950 766.050 133.050 ;
        RECT 767.400 132.900 768.600 133.950 ;
        RECT 773.400 132.900 774.600 133.950 ;
        RECT 764.400 115.050 765.600 130.950 ;
        RECT 766.950 130.800 769.050 132.900 ;
        RECT 772.950 130.800 775.050 132.900 ;
        RECT 778.950 130.950 781.050 133.050 ;
        RECT 766.950 118.950 769.050 121.050 ;
        RECT 763.950 112.950 766.050 115.050 ;
        RECT 746.700 104.700 755.250 105.900 ;
        RECT 743.400 102.900 745.500 103.050 ;
        RECT 742.950 100.950 745.500 102.900 ;
        RECT 742.950 100.800 745.050 100.950 ;
        RECT 743.400 98.400 744.600 100.800 ;
        RECT 746.700 95.700 747.600 104.700 ;
        RECT 753.150 103.800 755.250 104.700 ;
        RECT 756.150 102.900 757.050 108.300 ;
        RECT 761.400 107.400 765.600 108.600 ;
        RECT 758.400 103.050 759.600 105.600 ;
        RECT 750.300 101.700 757.050 102.900 ;
        RECT 750.300 99.300 751.200 101.700 ;
        RECT 749.100 97.200 751.200 99.300 ;
        RECT 752.100 98.100 754.200 100.200 ;
        RECT 745.800 93.600 747.900 95.700 ;
        RECT 752.400 95.550 753.600 98.100 ;
        RECT 756.000 94.500 757.050 101.700 ;
        RECT 757.950 100.950 760.050 103.050 ;
        RECT 764.400 97.050 765.600 107.400 ;
        RECT 767.400 99.900 768.600 118.950 ;
        RECT 769.950 103.950 772.050 109.050 ;
        RECT 779.400 108.600 780.600 130.950 ;
        RECT 782.400 121.050 783.600 172.650 ;
        RECT 788.400 154.050 789.600 178.950 ;
        RECT 793.950 175.950 796.050 178.050 ;
        RECT 787.950 151.950 790.050 154.050 ;
        RECT 794.400 151.050 795.600 175.950 ;
        RECT 793.950 148.950 796.050 151.050 ;
        RECT 784.950 145.950 787.050 148.050 ;
        RECT 785.400 139.050 786.600 145.950 ;
        RECT 797.400 145.050 798.600 190.950 ;
        RECT 806.400 187.050 807.600 197.400 ;
        RECT 808.950 193.950 811.050 196.050 ;
        RECT 799.950 184.950 802.050 187.050 ;
        RECT 802.950 184.950 805.050 187.050 ;
        RECT 805.950 184.950 808.050 187.050 ;
        RECT 790.950 142.950 793.050 145.050 ;
        RECT 796.950 142.950 799.050 145.050 ;
        RECT 784.950 136.950 787.050 139.050 ;
        RECT 791.400 136.050 792.600 142.950 ;
        RECT 796.950 138.000 799.050 141.900 ;
        RECT 800.400 139.050 801.600 184.950 ;
        RECT 797.400 136.050 798.600 138.000 ;
        RECT 799.950 136.950 802.050 139.050 ;
        RECT 787.950 133.950 790.050 136.050 ;
        RECT 790.950 133.950 793.050 136.050 ;
        RECT 793.950 133.950 796.050 136.050 ;
        RECT 796.950 133.950 799.050 136.050 ;
        RECT 784.950 130.950 787.050 133.050 ;
        RECT 788.400 132.900 789.600 133.950 ;
        RECT 781.950 118.950 784.050 121.050 ;
        RECT 785.400 112.050 786.600 130.950 ;
        RECT 787.950 130.800 790.050 132.900 ;
        RECT 787.950 124.950 790.050 127.050 ;
        RECT 784.950 109.950 787.050 112.050 ;
        RECT 776.400 107.400 780.600 108.600 ;
        RECT 776.400 103.050 777.600 107.400 ;
        RECT 781.950 104.100 784.050 109.050 ;
        RECT 782.400 103.050 783.600 104.100 ;
        RECT 772.950 100.950 775.050 103.050 ;
        RECT 775.950 100.950 778.050 103.050 ;
        RECT 778.950 100.950 781.050 103.050 ;
        RECT 781.950 100.950 784.050 103.050 ;
        RECT 773.400 99.900 774.600 100.950 ;
        RECT 766.950 97.800 769.050 99.900 ;
        RECT 772.950 97.800 775.050 99.900 ;
        RECT 779.400 99.000 780.600 100.950 ;
        RECT 763.950 94.950 766.050 97.050 ;
        RECT 755.400 92.400 757.500 94.500 ;
        RECT 739.950 88.950 742.050 91.050 ;
        RECT 745.950 88.950 748.050 91.050 ;
        RECT 736.950 61.950 739.050 64.050 ;
        RECT 742.950 61.950 745.050 64.050 ;
        RECT 721.950 59.100 724.050 61.200 ;
        RECT 727.950 59.100 730.050 61.200 ;
        RECT 733.950 59.100 736.050 61.200 ;
        RECT 709.950 52.800 712.050 54.900 ;
        RECT 718.950 52.800 721.050 54.900 ;
        RECT 722.400 52.050 723.600 59.100 ;
        RECT 728.400 58.050 729.600 59.100 ;
        RECT 734.400 58.050 735.600 59.100 ;
        RECT 727.950 55.950 730.050 58.050 ;
        RECT 730.950 55.950 733.050 58.050 ;
        RECT 733.950 55.950 736.050 58.050 ;
        RECT 736.950 55.950 739.050 58.050 ;
        RECT 731.400 54.900 732.600 55.950 ;
        RECT 730.950 52.800 733.050 54.900 ;
        RECT 721.950 49.950 724.050 52.050 ;
        RECT 737.400 46.050 738.600 55.950 ;
        RECT 739.950 52.950 742.050 55.050 ;
        RECT 736.950 43.950 739.050 46.050 ;
        RECT 733.950 37.950 736.050 40.050 ;
        RECT 734.400 28.200 735.600 37.950 ;
        RECT 740.400 37.050 741.600 52.950 ;
        RECT 739.950 34.950 742.050 37.050 ;
        RECT 712.950 26.100 715.050 28.200 ;
        RECT 718.950 26.100 721.050 28.200 ;
        RECT 733.950 26.100 736.050 28.200 ;
        RECT 713.400 25.050 714.600 26.100 ;
        RECT 719.400 25.050 720.600 26.100 ;
        RECT 734.400 25.050 735.600 26.100 ;
        RECT 709.950 22.950 712.050 25.050 ;
        RECT 712.950 22.950 715.050 25.050 ;
        RECT 715.950 22.950 718.050 25.050 ;
        RECT 718.950 22.950 721.050 25.050 ;
        RECT 730.950 22.950 733.050 25.050 ;
        RECT 733.950 22.950 736.050 25.050 ;
        RECT 736.950 22.950 739.050 25.050 ;
        RECT 710.400 21.000 711.600 22.950 ;
        RECT 703.950 16.950 706.050 19.050 ;
        RECT 709.950 16.950 712.050 21.000 ;
        RECT 716.400 16.050 717.600 22.950 ;
        RECT 731.400 21.600 732.600 22.950 ;
        RECT 737.400 21.900 738.600 22.950 ;
        RECT 728.400 21.000 732.600 21.600 ;
        RECT 727.950 20.400 732.600 21.000 ;
        RECT 727.950 16.950 730.050 20.400 ;
        RECT 736.950 19.800 739.050 21.900 ;
        RECT 743.400 16.050 744.600 61.950 ;
        RECT 746.400 40.050 747.600 88.950 ;
        RECT 751.950 79.950 754.050 85.050 ;
        RECT 748.950 67.950 751.050 70.050 ;
        RECT 760.950 67.950 763.050 70.050 ;
        RECT 745.950 37.950 748.050 40.050 ;
        RECT 745.950 34.800 748.050 36.900 ;
        RECT 746.400 22.050 747.600 34.800 ;
        RECT 749.400 28.200 750.600 67.950 ;
        RECT 754.950 59.100 757.050 61.200 ;
        RECT 755.400 58.050 756.600 59.100 ;
        RECT 761.400 58.050 762.600 67.950 ;
        RECT 764.400 61.050 765.600 94.950 ;
        RECT 763.950 58.950 766.050 61.050 ;
        RECT 754.950 55.950 757.050 58.050 ;
        RECT 757.950 55.950 760.050 58.050 ;
        RECT 760.950 55.950 763.050 58.050 ;
        RECT 758.400 54.000 759.600 55.950 ;
        RECT 757.950 49.950 760.050 54.000 ;
        RECT 767.400 31.050 768.600 97.800 ;
        RECT 773.400 58.050 774.600 97.800 ;
        RECT 778.950 94.950 781.050 99.000 ;
        RECT 784.950 94.950 787.050 97.050 ;
        RECT 785.400 88.050 786.600 94.950 ;
        RECT 784.950 85.950 787.050 88.050 ;
        RECT 778.950 60.000 781.050 64.050 ;
        RECT 779.400 58.050 780.600 60.000 ;
        RECT 772.950 55.950 775.050 58.050 ;
        RECT 775.950 55.950 778.050 58.050 ;
        RECT 778.950 55.950 781.050 58.050 ;
        RECT 781.950 55.950 784.050 58.050 ;
        RECT 769.950 52.950 772.050 55.050 ;
        RECT 776.400 54.900 777.600 55.950 ;
        RECT 766.950 28.950 769.050 31.050 ;
        RECT 748.950 26.100 751.050 28.200 ;
        RECT 760.950 26.100 763.050 28.200 ;
        RECT 761.400 25.050 762.600 26.100 ;
        RECT 754.950 22.950 757.050 25.050 ;
        RECT 760.950 22.950 763.050 25.050 ;
        RECT 763.950 22.950 766.050 25.050 ;
        RECT 745.950 19.950 748.050 22.050 ;
        RECT 755.400 21.900 756.600 22.950 ;
        RECT 764.400 21.900 765.600 22.950 ;
        RECT 770.400 22.050 771.600 52.950 ;
        RECT 775.950 52.800 778.050 54.900 ;
        RECT 782.400 25.050 783.600 55.950 ;
        RECT 784.950 49.950 787.050 54.900 ;
        RECT 788.400 46.050 789.600 124.950 ;
        RECT 794.400 105.600 795.600 133.950 ;
        RECT 803.400 115.050 804.600 184.950 ;
        RECT 809.400 181.050 810.600 193.950 ;
        RECT 812.400 187.050 813.600 238.950 ;
        RECT 815.400 187.200 816.600 250.950 ;
        RECT 821.400 241.050 822.600 256.950 ;
        RECT 826.950 253.950 829.050 256.050 ;
        RECT 820.950 238.950 823.050 241.050 ;
        RECT 820.950 232.950 823.050 235.050 ;
        RECT 821.400 214.050 822.600 232.950 ;
        RECT 827.400 217.050 828.600 253.950 ;
        RECT 830.400 220.050 831.600 265.950 ;
        RECT 833.400 262.050 834.600 269.400 ;
        RECT 832.950 259.950 835.050 262.050 ;
        RECT 839.400 259.050 840.600 280.950 ;
        RECT 845.400 277.050 846.600 292.950 ;
        RECT 844.950 274.950 847.050 277.050 ;
        RECT 848.400 271.050 849.600 301.950 ;
        RECT 853.950 301.800 856.050 303.900 ;
        RECT 850.950 295.950 853.050 298.050 ;
        RECT 847.950 268.950 850.050 271.050 ;
        RECT 844.950 260.100 847.050 262.200 ;
        RECT 845.400 259.050 846.600 260.100 ;
        RECT 835.950 256.950 838.050 259.050 ;
        RECT 838.950 256.950 841.050 259.050 ;
        RECT 841.950 256.950 844.050 259.050 ;
        RECT 844.950 256.950 847.050 259.050 ;
        RECT 832.950 253.950 835.050 256.050 ;
        RECT 833.400 232.050 834.600 253.950 ;
        RECT 836.400 250.050 837.600 256.950 ;
        RECT 838.950 250.950 841.050 253.050 ;
        RECT 835.950 247.950 838.050 250.050 ;
        RECT 839.400 238.050 840.600 250.950 ;
        RECT 842.400 244.050 843.600 256.950 ;
        RECT 847.950 253.950 850.050 256.050 ;
        RECT 848.400 250.050 849.600 253.950 ;
        RECT 847.950 247.950 850.050 250.050 ;
        RECT 841.950 241.950 844.050 244.050 ;
        RECT 838.950 235.950 841.050 238.050 ;
        RECT 832.950 229.950 835.050 232.050 ;
        RECT 838.950 226.950 841.050 229.050 ;
        RECT 829.950 217.950 832.050 220.050 ;
        RECT 835.950 217.950 838.050 220.050 ;
        RECT 826.950 216.600 829.050 217.050 ;
        RECT 826.950 215.400 831.600 216.600 ;
        RECT 826.950 214.950 829.050 215.400 ;
        RECT 830.400 214.050 831.600 215.400 ;
        RECT 820.950 211.950 823.050 214.050 ;
        RECT 823.950 211.950 826.050 214.050 ;
        RECT 829.950 211.950 832.050 214.050 ;
        RECT 824.400 196.050 825.600 211.950 ;
        RECT 826.950 208.950 829.050 211.050 ;
        RECT 836.400 210.900 837.600 217.950 ;
        RECT 839.400 216.600 840.600 226.950 ;
        RECT 851.400 223.050 852.600 295.950 ;
        RECT 854.400 295.050 855.600 301.800 ;
        RECT 857.400 298.050 858.600 370.950 ;
        RECT 863.400 370.050 864.600 379.950 ;
        RECT 868.950 372.000 871.050 376.050 ;
        RECT 869.400 370.050 870.600 372.000 ;
        RECT 862.950 367.950 865.050 370.050 ;
        RECT 865.950 367.950 868.050 370.050 ;
        RECT 868.950 367.950 871.050 370.050 ;
        RECT 871.950 367.950 874.050 370.050 ;
        RECT 866.400 366.900 867.600 367.950 ;
        RECT 865.950 364.800 868.050 366.900 ;
        RECT 865.950 352.950 868.050 355.050 ;
        RECT 859.950 343.950 862.050 346.050 ;
        RECT 860.400 340.050 861.600 343.950 ;
        RECT 866.400 340.200 867.600 352.950 ;
        RECT 872.400 349.050 873.600 367.950 ;
        RECT 871.950 346.950 874.050 349.050 ;
        RECT 859.950 337.950 862.050 340.050 ;
        RECT 865.800 338.100 867.900 340.200 ;
        RECT 871.950 338.100 874.050 340.200 ;
        RECT 866.400 337.050 867.600 338.100 ;
        RECT 872.400 337.050 873.600 338.100 ;
        RECT 862.950 334.950 865.050 337.050 ;
        RECT 865.950 334.950 868.050 337.050 ;
        RECT 868.950 334.950 871.050 337.050 ;
        RECT 871.950 334.950 874.050 337.050 ;
        RECT 863.400 333.900 864.600 334.950 ;
        RECT 862.950 331.800 865.050 333.900 ;
        RECT 869.400 333.000 870.600 334.950 ;
        RECT 859.950 328.950 862.050 331.050 ;
        RECT 860.400 313.050 861.600 328.950 ;
        RECT 859.950 310.950 862.050 313.050 ;
        RECT 856.950 295.950 859.050 298.050 ;
        RECT 853.950 292.950 856.050 295.050 ;
        RECT 860.400 292.050 861.600 310.950 ;
        RECT 863.400 298.050 864.600 331.800 ;
        RECT 865.800 328.950 867.900 331.050 ;
        RECT 868.950 328.950 871.050 333.000 ;
        RECT 878.400 331.050 879.600 440.400 ;
        RECT 886.950 439.950 889.050 442.050 ;
        RECT 880.950 430.950 883.050 433.050 ;
        RECT 881.400 418.050 882.600 430.950 ;
        RECT 887.400 424.050 888.600 439.950 ;
        RECT 886.950 421.950 889.050 424.050 ;
        RECT 890.400 421.050 891.600 445.950 ;
        RECT 892.950 442.950 895.050 445.050 ;
        RECT 893.400 439.050 894.600 442.950 ;
        RECT 892.950 436.950 895.050 439.050 ;
        RECT 896.400 430.050 897.600 469.950 ;
        RECT 895.950 427.950 898.050 430.050 ;
        RECT 889.950 418.950 892.050 421.050 ;
        RECT 880.950 415.950 883.050 418.050 ;
        RECT 886.950 416.100 889.050 418.200 ;
        RECT 887.400 415.050 888.600 416.100 ;
        RECT 895.950 415.950 898.050 418.050 ;
        RECT 883.950 412.950 886.050 415.050 ;
        RECT 886.950 412.950 889.050 415.050 ;
        RECT 889.950 412.950 892.050 415.050 ;
        RECT 884.400 411.900 885.600 412.950 ;
        RECT 890.400 411.900 891.600 412.950 ;
        RECT 883.950 409.800 886.050 411.900 ;
        RECT 889.950 409.800 892.050 411.900 ;
        RECT 880.950 406.950 883.050 409.050 ;
        RECT 877.950 328.950 880.050 331.050 ;
        RECT 866.400 298.050 867.600 328.950 ;
        RECT 869.400 319.050 870.600 328.950 ;
        RECT 868.950 316.950 871.050 319.050 ;
        RECT 881.400 313.050 882.600 406.950 ;
        RECT 883.950 406.650 886.050 408.750 ;
        RECT 880.950 310.950 883.050 313.050 ;
        RECT 868.950 304.950 871.050 307.050 ;
        RECT 862.950 295.950 865.050 298.050 ;
        RECT 865.950 295.950 868.050 298.050 ;
        RECT 866.400 292.050 867.600 295.950 ;
        RECT 869.400 295.050 870.600 304.950 ;
        RECT 871.950 295.950 874.050 298.050 ;
        RECT 868.950 292.950 871.050 295.050 ;
        RECT 856.950 289.950 859.050 292.050 ;
        RECT 859.950 289.950 862.050 292.050 ;
        RECT 862.950 289.950 865.050 292.050 ;
        RECT 865.950 289.950 868.050 292.050 ;
        RECT 857.400 271.050 858.600 289.950 ;
        RECT 863.400 288.900 864.600 289.950 ;
        RECT 862.950 286.800 865.050 288.900 ;
        RECT 872.400 286.050 873.600 295.950 ;
        RECT 877.950 293.100 880.050 298.050 ;
        RECT 881.400 297.600 882.600 310.950 ;
        RECT 884.400 301.050 885.600 406.650 ;
        RECT 886.950 400.950 889.050 403.050 ;
        RECT 887.400 304.050 888.600 400.950 ;
        RECT 890.400 397.050 891.600 409.800 ;
        RECT 892.950 403.950 895.050 406.050 ;
        RECT 889.950 394.950 892.050 397.050 ;
        RECT 890.400 346.050 891.600 394.950 ;
        RECT 889.950 343.950 892.050 346.050 ;
        RECT 889.950 337.950 892.050 340.050 ;
        RECT 886.950 301.950 889.050 304.050 ;
        RECT 883.950 298.950 886.050 301.050 ;
        RECT 881.400 296.400 885.600 297.600 ;
        RECT 878.400 292.050 879.600 293.100 ;
        RECT 884.400 292.050 885.600 296.400 ;
        RECT 890.400 295.050 891.600 337.950 ;
        RECT 889.950 292.950 892.050 295.050 ;
        RECT 877.950 289.950 880.050 292.050 ;
        RECT 880.950 289.950 883.050 292.050 ;
        RECT 883.950 289.950 886.050 292.050 ;
        RECT 886.950 289.950 889.050 292.050 ;
        RECT 881.400 288.000 882.600 289.950 ;
        RECT 871.950 283.950 874.050 286.050 ;
        RECT 880.950 283.950 883.050 288.000 ;
        RECT 868.950 280.950 871.050 283.050 ;
        RECT 877.950 280.950 880.050 283.050 ;
        RECT 859.950 277.950 862.050 280.050 ;
        RECT 853.950 268.950 856.050 271.050 ;
        RECT 856.950 268.950 859.050 271.050 ;
        RECT 854.400 240.600 855.600 268.950 ;
        RECT 857.400 259.050 858.600 268.950 ;
        RECT 860.400 262.050 861.600 277.950 ;
        RECT 862.950 265.950 865.050 268.050 ;
        RECT 859.950 259.950 862.050 262.050 ;
        RECT 863.400 259.050 864.600 265.950 ;
        RECT 869.400 262.200 870.600 280.950 ;
        RECT 868.950 260.100 871.050 262.200 ;
        RECT 869.400 259.050 870.600 260.100 ;
        RECT 856.950 256.950 859.050 259.050 ;
        RECT 862.950 256.950 865.050 259.050 ;
        RECT 865.950 256.950 868.050 259.050 ;
        RECT 868.950 256.950 871.050 259.050 ;
        RECT 871.950 256.950 874.050 259.050 ;
        RECT 862.950 247.950 865.050 250.050 ;
        RECT 854.400 239.400 858.600 240.600 ;
        RECT 853.950 235.950 856.050 238.050 ;
        RECT 850.950 220.950 853.050 223.050 ;
        RECT 839.400 215.400 843.600 216.600 ;
        RECT 847.950 216.000 850.050 220.050 ;
        RECT 854.400 217.050 855.600 235.950 ;
        RECT 842.400 214.050 843.600 215.400 ;
        RECT 848.400 214.050 849.600 216.000 ;
        RECT 853.950 214.950 856.050 217.050 ;
        RECT 841.950 211.950 844.050 214.050 ;
        RECT 844.950 211.950 847.050 214.050 ;
        RECT 847.950 211.950 850.050 214.050 ;
        RECT 850.950 211.950 853.050 214.050 ;
        RECT 845.400 210.900 846.600 211.950 ;
        RECT 823.950 193.950 826.050 196.050 ;
        RECT 811.950 184.950 814.050 187.050 ;
        RECT 814.950 185.100 817.050 187.200 ;
        RECT 820.950 184.950 823.050 187.050 ;
        RECT 814.950 181.950 817.050 184.050 ;
        RECT 815.400 181.050 816.600 181.950 ;
        RECT 808.950 178.950 811.050 181.050 ;
        RECT 811.950 178.950 814.050 181.050 ;
        RECT 814.950 178.950 817.050 181.050 ;
        RECT 805.950 175.950 808.050 178.050 ;
        RECT 812.400 177.000 813.600 178.950 ;
        RECT 806.400 127.050 807.600 175.950 ;
        RECT 811.950 172.950 814.050 177.000 ;
        RECT 817.950 175.950 820.050 178.050 ;
        RECT 818.400 172.050 819.600 175.950 ;
        RECT 817.950 169.950 820.050 172.050 ;
        RECT 817.950 166.800 820.050 168.900 ;
        RECT 818.400 145.050 819.600 166.800 ;
        RECT 817.950 142.950 820.050 145.050 ;
        RECT 811.950 141.600 816.000 142.050 ;
        RECT 811.950 139.950 816.600 141.600 ;
        RECT 808.950 136.950 811.050 139.050 ;
        RECT 805.950 124.950 808.050 127.050 ;
        RECT 805.950 115.950 808.050 118.050 ;
        RECT 796.950 112.950 799.050 115.050 ;
        RECT 802.950 112.950 805.050 115.050 ;
        RECT 797.400 108.600 798.600 112.950 ;
        RECT 806.400 111.600 807.600 115.950 ;
        RECT 800.400 110.400 807.600 111.600 ;
        RECT 809.400 111.600 810.600 136.950 ;
        RECT 815.400 136.050 816.600 139.950 ;
        RECT 821.400 139.050 822.600 184.950 ;
        RECT 824.400 184.050 825.600 193.950 ;
        RECT 827.400 187.050 828.600 208.950 ;
        RECT 835.950 208.800 838.050 210.900 ;
        RECT 844.950 208.800 847.050 210.900 ;
        RECT 835.950 202.950 838.050 205.050 ;
        RECT 829.950 187.950 832.050 190.050 ;
        RECT 826.950 184.950 829.050 187.050 ;
        RECT 823.950 181.950 826.050 184.050 ;
        RECT 830.400 181.050 831.600 187.950 ;
        RECT 836.400 184.050 837.600 202.950 ;
        RECT 838.950 199.950 841.050 202.050 ;
        RECT 835.950 181.950 838.050 184.050 ;
        RECT 826.950 178.950 829.050 181.050 ;
        RECT 829.950 178.950 832.050 181.050 ;
        RECT 832.950 178.950 835.050 181.050 ;
        RECT 827.400 177.900 828.600 178.950 ;
        RECT 833.400 177.900 834.600 178.950 ;
        RECT 826.950 175.800 829.050 177.900 ;
        RECT 832.950 175.800 835.050 177.900 ;
        RECT 835.950 175.950 838.050 178.050 ;
        RECT 836.400 172.050 837.600 175.950 ;
        RECT 835.950 169.950 838.050 172.050 ;
        RECT 823.950 163.950 826.050 166.050 ;
        RECT 824.400 142.050 825.600 163.950 ;
        RECT 826.950 157.950 829.050 160.050 ;
        RECT 823.950 139.950 826.050 142.050 ;
        RECT 820.950 136.950 823.050 139.050 ;
        RECT 814.950 133.950 817.050 136.050 ;
        RECT 817.950 133.950 820.050 136.050 ;
        RECT 818.400 132.000 819.600 133.950 ;
        RECT 817.950 127.950 820.050 132.000 ;
        RECT 820.950 130.950 823.050 133.050 ;
        RECT 821.400 112.050 822.600 130.950 ;
        RECT 824.400 112.050 825.600 139.950 ;
        RECT 827.400 133.050 828.600 157.950 ;
        RECT 829.950 148.950 832.050 151.050 ;
        RECT 830.400 139.050 831.600 148.950 ;
        RECT 839.400 148.050 840.600 199.950 ;
        RECT 851.400 196.050 852.600 211.950 ;
        RECT 853.950 208.950 856.050 211.050 ;
        RECT 850.950 193.950 853.050 196.050 ;
        RECT 841.950 184.950 844.050 190.050 ;
        RECT 854.400 187.050 855.600 208.950 ;
        RECT 857.400 202.050 858.600 239.400 ;
        RECT 863.400 225.600 864.600 247.950 ;
        RECT 866.400 232.050 867.600 256.950 ;
        RECT 872.400 255.900 873.600 256.950 ;
        RECT 871.950 253.800 874.050 255.900 ;
        RECT 868.950 250.950 871.050 253.050 ;
        RECT 865.950 229.950 868.050 232.050 ;
        RECT 863.400 224.400 867.600 225.600 ;
        RECT 862.950 220.950 865.050 223.050 ;
        RECT 859.950 217.950 862.050 220.050 ;
        RECT 856.950 199.950 859.050 202.050 ;
        RECT 856.950 193.950 859.050 196.050 ;
        RECT 853.950 184.950 856.050 187.050 ;
        RECT 841.950 181.800 844.050 183.900 ;
        RECT 850.950 182.100 853.050 184.200 ;
        RECT 857.400 184.050 858.600 193.950 ;
        RECT 842.400 172.050 843.600 181.800 ;
        RECT 851.400 181.050 852.600 182.100 ;
        RECT 856.950 181.950 859.050 184.050 ;
        RECT 847.950 178.950 850.050 181.050 ;
        RECT 850.950 178.950 853.050 181.050 ;
        RECT 853.950 178.950 856.050 181.050 ;
        RECT 848.400 177.900 849.600 178.950 ;
        RECT 847.950 175.800 850.050 177.900 ;
        RECT 850.950 172.950 853.050 175.050 ;
        RECT 842.400 170.400 847.050 172.050 ;
        RECT 843.000 169.950 847.050 170.400 ;
        RECT 838.950 145.950 841.050 148.050 ;
        RECT 847.950 145.950 850.050 148.050 ;
        RECT 829.950 136.950 832.050 139.050 ;
        RECT 832.950 138.000 835.050 142.050 ;
        RECT 835.950 141.600 838.050 145.050 ;
        RECT 835.950 141.000 840.600 141.600 ;
        RECT 836.400 140.400 840.600 141.000 ;
        RECT 833.400 136.050 834.600 138.000 ;
        RECT 839.400 136.050 840.600 140.400 ;
        RECT 832.950 133.950 835.050 136.050 ;
        RECT 835.950 133.950 838.050 136.050 ;
        RECT 838.950 133.950 841.050 136.050 ;
        RECT 841.950 133.950 844.050 136.050 ;
        RECT 826.950 130.950 829.050 133.050 ;
        RECT 829.950 130.950 832.050 133.050 ;
        RECT 836.400 132.900 837.600 133.950 ;
        RECT 842.400 133.050 843.600 133.950 ;
        RECT 809.400 110.400 813.600 111.600 ;
        RECT 800.400 108.600 801.600 110.400 ;
        RECT 797.400 107.400 801.600 108.600 ;
        RECT 791.400 104.400 795.600 105.600 ;
        RECT 791.400 97.050 792.600 104.400 ;
        RECT 800.400 103.050 801.600 107.400 ;
        RECT 805.950 104.100 808.050 106.200 ;
        RECT 806.400 103.050 807.600 104.100 ;
        RECT 796.950 100.950 799.050 103.050 ;
        RECT 799.950 100.950 802.050 103.050 ;
        RECT 802.950 100.950 805.050 103.050 ;
        RECT 805.950 100.950 808.050 103.050 ;
        RECT 797.400 99.900 798.600 100.950 ;
        RECT 796.950 97.800 799.050 99.900 ;
        RECT 790.950 94.950 793.050 97.050 ;
        RECT 790.950 91.800 793.050 93.900 ;
        RECT 787.950 43.950 790.050 46.050 ;
        RECT 791.400 43.050 792.600 91.800 ;
        RECT 797.400 91.050 798.600 97.800 ;
        RECT 799.950 91.950 802.050 97.050 ;
        RECT 803.400 96.600 804.600 100.950 ;
        RECT 803.400 95.400 807.600 96.600 ;
        RECT 796.950 88.950 799.050 91.050 ;
        RECT 799.950 60.000 802.050 64.050 ;
        RECT 800.400 58.050 801.600 60.000 ;
        RECT 796.950 55.950 799.050 58.050 ;
        RECT 799.950 55.950 802.050 58.050 ;
        RECT 793.950 52.950 796.050 55.050 ;
        RECT 797.400 54.900 798.600 55.950 ;
        RECT 794.400 49.050 795.600 52.950 ;
        RECT 796.950 52.800 799.050 54.900 ;
        RECT 793.950 46.950 796.050 49.050 ;
        RECT 790.950 40.950 793.050 43.050 ;
        RECT 793.950 25.950 796.050 28.050 ;
        RECT 797.400 27.600 798.600 52.800 ;
        RECT 806.400 52.050 807.600 95.400 ;
        RECT 808.950 61.950 811.050 64.050 ;
        RECT 805.950 49.950 808.050 52.050 ;
        RECT 809.400 34.050 810.600 61.950 ;
        RECT 812.400 61.050 813.600 110.400 ;
        RECT 817.950 109.950 820.050 112.050 ;
        RECT 820.950 109.950 823.050 112.050 ;
        RECT 823.950 109.950 826.050 112.050 ;
        RECT 818.400 100.050 819.600 109.950 ;
        RECT 830.400 109.200 831.600 130.950 ;
        RECT 835.950 130.800 838.050 132.900 ;
        RECT 842.400 131.400 847.050 133.050 ;
        RECT 843.000 130.950 847.050 131.400 ;
        RECT 844.950 127.800 847.050 129.900 ;
        RECT 838.950 124.950 841.050 127.050 ;
        RECT 835.950 118.950 838.050 121.050 ;
        RECT 829.950 107.100 832.050 109.200 ;
        RECT 823.950 104.100 826.050 106.200 ;
        RECT 824.400 103.050 825.600 104.100 ;
        RECT 829.950 103.950 832.050 106.050 ;
        RECT 830.400 103.050 831.600 103.950 ;
        RECT 823.950 100.950 826.050 103.050 ;
        RECT 826.950 100.950 829.050 103.050 ;
        RECT 829.950 100.950 832.050 103.050 ;
        RECT 817.950 97.950 820.050 100.050 ;
        RECT 827.400 99.900 828.600 100.950 ;
        RECT 826.950 97.800 829.050 99.900 ;
        RECT 832.950 97.950 835.050 100.050 ;
        RECT 823.950 91.950 826.050 94.050 ;
        RECT 811.950 58.950 814.050 61.050 ;
        RECT 817.950 60.000 820.050 64.050 ;
        RECT 818.400 58.050 819.600 60.000 ;
        RECT 814.950 55.950 817.050 58.050 ;
        RECT 817.950 55.950 820.050 58.050 ;
        RECT 815.400 49.050 816.600 55.950 ;
        RECT 824.400 49.050 825.600 91.950 ;
        RECT 833.400 88.050 834.600 97.950 ;
        RECT 836.400 97.050 837.600 118.950 ;
        RECT 839.400 106.050 840.600 124.950 ;
        RECT 841.950 121.950 844.050 124.050 ;
        RECT 842.400 118.050 843.600 121.950 ;
        RECT 841.950 115.950 844.050 118.050 ;
        RECT 841.950 109.950 844.050 112.050 ;
        RECT 838.950 103.950 841.050 106.050 ;
        RECT 842.400 103.050 843.600 109.950 ;
        RECT 845.400 108.600 846.600 127.800 ;
        RECT 848.400 118.050 849.600 145.950 ;
        RECT 851.400 133.050 852.600 172.950 ;
        RECT 854.400 163.050 855.600 178.950 ;
        RECT 853.950 160.950 856.050 163.050 ;
        RECT 856.950 151.950 859.050 154.050 ;
        RECT 857.400 136.050 858.600 151.950 ;
        RECT 860.400 142.050 861.600 217.950 ;
        RECT 859.950 139.950 862.050 142.050 ;
        RECT 863.400 138.600 864.600 220.950 ;
        RECT 866.400 217.050 867.600 224.400 ;
        RECT 865.950 214.950 868.050 217.050 ;
        RECT 869.400 214.050 870.600 250.950 ;
        RECT 872.400 220.050 873.600 253.800 ;
        RECT 874.950 223.950 877.050 226.050 ;
        RECT 871.950 217.950 874.050 220.050 ;
        RECT 875.400 214.050 876.600 223.950 ;
        RECT 878.400 220.050 879.600 280.950 ;
        RECT 880.950 268.950 883.050 271.050 ;
        RECT 881.400 250.050 882.600 268.950 ;
        RECT 883.950 265.950 886.050 268.050 ;
        RECT 880.950 247.950 883.050 250.050 ;
        RECT 884.400 241.050 885.600 265.950 ;
        RECT 883.950 238.950 886.050 241.050 ;
        RECT 880.950 229.950 883.050 232.050 ;
        RECT 877.950 217.950 880.050 220.050 ;
        RECT 881.400 216.600 882.600 229.950 ;
        RECT 887.400 226.050 888.600 289.950 ;
        RECT 889.950 286.950 892.050 289.050 ;
        RECT 890.400 255.900 891.600 286.950 ;
        RECT 889.950 253.800 892.050 255.900 ;
        RECT 889.950 241.950 892.050 244.050 ;
        RECT 886.950 223.950 889.050 226.050 ;
        RECT 881.400 215.400 885.600 216.600 ;
        RECT 868.950 211.950 871.050 214.050 ;
        RECT 871.950 211.950 874.050 214.050 ;
        RECT 874.950 211.950 877.050 214.050 ;
        RECT 877.950 211.950 880.050 214.050 ;
        RECT 865.950 208.950 868.050 211.050 ;
        RECT 872.400 210.900 873.600 211.950 ;
        RECT 866.400 184.050 867.600 208.950 ;
        RECT 871.950 208.800 874.050 210.900 ;
        RECT 878.400 195.600 879.600 211.950 ;
        RECT 884.400 210.600 885.600 215.400 ;
        RECT 881.400 209.400 885.600 210.600 ;
        RECT 881.400 195.600 882.600 209.400 ;
        RECT 883.950 205.950 886.050 208.050 ;
        RECT 878.400 194.400 882.600 195.600 ;
        RECT 871.950 187.950 874.050 190.050 ;
        RECT 865.950 181.950 868.050 184.050 ;
        RECT 872.400 181.050 873.600 187.950 ;
        RECT 868.950 178.950 871.050 181.050 ;
        RECT 871.950 178.950 874.050 181.050 ;
        RECT 874.950 178.950 877.050 181.050 ;
        RECT 865.950 175.950 868.050 178.050 ;
        RECT 869.400 177.000 870.600 178.950 ;
        RECT 866.400 142.050 867.600 175.950 ;
        RECT 868.950 172.950 871.050 177.000 ;
        RECT 875.400 172.050 876.600 178.950 ;
        RECT 877.950 175.950 880.050 178.050 ;
        RECT 874.950 169.950 877.050 172.050 ;
        RECT 871.950 166.950 874.050 169.050 ;
        RECT 865.950 139.950 868.050 142.050 ;
        RECT 872.400 139.200 873.600 166.950 ;
        RECT 878.400 148.050 879.600 175.950 ;
        RECT 881.400 169.050 882.600 194.400 ;
        RECT 880.950 166.950 883.050 169.050 ;
        RECT 877.950 145.950 880.050 148.050 ;
        RECT 863.400 137.400 867.600 138.600 ;
        RECT 856.950 133.950 859.050 136.050 ;
        RECT 859.950 133.950 862.050 136.050 ;
        RECT 850.950 130.800 853.050 133.050 ;
        RECT 860.400 132.900 861.600 133.950 ;
        RECT 859.950 130.800 862.050 132.900 ;
        RECT 847.950 115.950 850.050 118.050 ;
        RECT 866.400 109.050 867.600 137.400 ;
        RECT 871.950 137.100 874.050 139.200 ;
        RECT 877.950 138.000 880.050 142.050 ;
        RECT 884.400 139.050 885.600 205.950 ;
        RECT 886.950 187.950 889.050 190.050 ;
        RECT 887.400 163.050 888.600 187.950 ;
        RECT 886.950 160.950 889.050 163.050 ;
        RECT 886.950 145.950 889.050 148.050 ;
        RECT 872.400 136.050 873.600 137.100 ;
        RECT 878.400 136.050 879.600 138.000 ;
        RECT 883.950 136.950 886.050 139.050 ;
        RECT 871.950 133.950 874.050 136.050 ;
        RECT 874.950 133.950 877.050 136.050 ;
        RECT 877.950 133.950 880.050 136.050 ;
        RECT 880.950 133.950 883.050 136.050 ;
        RECT 875.400 124.050 876.600 133.950 ;
        RECT 881.400 133.050 882.600 133.950 ;
        RECT 881.400 131.400 886.050 133.050 ;
        RECT 882.000 130.950 886.050 131.400 ;
        RECT 877.800 127.950 879.900 130.050 ;
        RECT 880.950 127.950 883.050 130.050 ;
        RECT 868.950 121.950 871.050 124.050 ;
        RECT 874.950 121.950 877.050 124.050 ;
        RECT 845.400 107.400 849.600 108.600 ;
        RECT 848.400 103.050 849.600 107.400 ;
        RECT 853.950 106.950 856.050 109.050 ;
        RECT 856.950 106.950 859.050 109.050 ;
        RECT 841.950 100.950 844.050 103.050 ;
        RECT 844.950 100.950 847.050 103.050 ;
        RECT 847.950 100.950 850.050 103.050 ;
        RECT 838.950 97.950 841.050 100.050 ;
        RECT 835.950 94.950 838.050 97.050 ;
        RECT 832.950 85.950 835.050 88.050 ;
        RECT 839.400 67.050 840.600 97.950 ;
        RECT 841.950 94.950 844.050 97.050 ;
        RECT 826.950 64.950 829.050 67.050 ;
        RECT 838.950 64.950 841.050 67.050 ;
        RECT 814.950 46.950 817.050 49.050 ;
        RECT 823.950 46.950 826.050 49.050 ;
        RECT 827.400 34.050 828.600 64.950 ;
        RECT 842.400 64.050 843.600 94.950 ;
        RECT 845.400 76.050 846.600 100.950 ;
        RECT 850.950 97.950 853.050 100.050 ;
        RECT 851.400 88.050 852.600 97.950 ;
        RECT 854.400 91.050 855.600 106.950 ;
        RECT 853.950 88.950 856.050 91.050 ;
        RECT 850.950 85.950 853.050 88.050 ;
        RECT 844.950 73.950 847.050 76.050 ;
        RECT 857.400 64.050 858.600 106.950 ;
        RECT 862.950 105.000 865.050 109.050 ;
        RECT 865.950 106.950 868.050 109.050 ;
        RECT 863.400 103.050 864.600 105.000 ;
        RECT 869.400 103.050 870.600 121.950 ;
        RECT 874.950 115.950 877.050 118.050 ;
        RECT 862.950 100.950 865.050 103.050 ;
        RECT 865.950 100.950 868.050 103.050 ;
        RECT 868.950 100.950 871.050 103.050 ;
        RECT 866.400 99.900 867.600 100.950 ;
        RECT 865.950 97.800 868.050 99.900 ;
        RECT 871.950 97.950 874.050 100.050 ;
        RECT 865.950 91.950 868.050 94.050 ;
        RECT 859.950 64.950 862.050 67.050 ;
        RECT 841.950 61.950 844.050 64.050 ;
        RECT 847.950 61.950 850.050 64.050 ;
        RECT 856.950 61.950 859.050 64.050 ;
        RECT 844.950 58.950 847.050 61.050 ;
        RECT 832.950 55.950 835.050 58.050 ;
        RECT 833.400 43.050 834.600 55.950 ;
        RECT 832.950 40.950 835.050 43.050 ;
        RECT 845.400 37.050 846.600 58.950 ;
        RECT 848.400 54.900 849.600 61.950 ;
        RECT 853.950 59.100 856.050 61.200 ;
        RECT 854.400 58.050 855.600 59.100 ;
        RECT 860.400 58.050 861.600 64.950 ;
        RECT 866.400 61.050 867.600 91.950 ;
        RECT 865.950 58.950 868.050 61.050 ;
        RECT 868.950 58.950 871.050 61.050 ;
        RECT 853.950 55.950 856.050 58.050 ;
        RECT 856.950 55.950 859.050 58.050 ;
        RECT 859.950 55.950 862.050 58.050 ;
        RECT 862.950 55.950 865.050 58.050 ;
        RECT 857.400 54.900 858.600 55.950 ;
        RECT 863.400 55.050 864.600 55.950 ;
        RECT 847.950 52.800 850.050 54.900 ;
        RECT 856.950 52.800 859.050 54.900 ;
        RECT 863.400 53.400 868.050 55.050 ;
        RECT 864.000 52.950 868.050 53.400 ;
        RECT 844.950 34.950 847.050 37.050 ;
        RECT 808.950 31.950 811.050 34.050 ;
        RECT 814.950 31.950 817.050 34.050 ;
        RECT 826.950 31.950 829.050 34.050 ;
        RECT 835.950 31.950 838.050 34.050 ;
        RECT 797.400 26.400 801.600 27.600 ;
        RECT 778.950 22.950 781.050 25.050 ;
        RECT 781.950 22.950 784.050 25.050 ;
        RECT 787.950 22.950 790.050 25.050 ;
        RECT 754.950 19.800 757.050 21.900 ;
        RECT 763.950 19.800 766.050 21.900 ;
        RECT 769.950 19.950 772.050 22.050 ;
        RECT 779.400 21.900 780.600 22.950 ;
        RECT 788.400 21.900 789.600 22.950 ;
        RECT 794.400 21.900 795.600 25.950 ;
        RECT 800.400 25.050 801.600 26.400 ;
        RECT 805.950 26.100 808.050 28.200 ;
        RECT 806.400 25.050 807.600 26.100 ;
        RECT 815.400 25.050 816.600 31.950 ;
        RECT 823.950 27.000 826.050 31.050 ;
        RECT 824.400 25.050 825.600 27.000 ;
        RECT 799.950 22.950 802.050 25.050 ;
        RECT 802.950 22.950 805.050 25.050 ;
        RECT 805.950 22.950 808.050 25.050 ;
        RECT 808.950 22.950 811.050 25.050 ;
        RECT 814.950 22.950 817.050 25.050 ;
        RECT 823.950 22.950 826.050 25.050 ;
        RECT 826.950 22.950 829.050 25.050 ;
        RECT 803.400 21.900 804.600 22.950 ;
        RECT 809.400 21.900 810.600 22.950 ;
        RECT 827.400 21.900 828.600 22.950 ;
        RECT 836.400 21.900 837.600 31.950 ;
        RECT 848.400 30.600 849.600 52.800 ;
        RECT 850.950 43.950 853.050 46.050 ;
        RECT 845.400 29.400 849.600 30.600 ;
        RECT 845.400 25.050 846.600 29.400 ;
        RECT 851.400 25.050 852.600 43.950 ;
        RECT 869.400 31.050 870.600 58.950 ;
        RECT 872.400 54.900 873.600 97.950 ;
        RECT 875.400 64.050 876.600 115.950 ;
        RECT 878.400 100.050 879.600 127.950 ;
        RECT 881.400 106.050 882.600 127.950 ;
        RECT 883.950 112.950 886.050 115.050 ;
        RECT 880.950 103.950 883.050 106.050 ;
        RECT 884.400 103.050 885.600 112.950 ;
        RECT 887.400 109.050 888.600 145.950 ;
        RECT 890.400 133.050 891.600 241.950 ;
        RECT 889.950 130.950 892.050 133.050 ;
        RECT 886.950 106.950 889.050 109.050 ;
        RECT 883.950 100.950 886.050 103.050 ;
        RECT 886.950 100.950 889.050 103.050 ;
        RECT 877.950 97.950 880.050 100.050 ;
        RECT 887.400 99.900 888.600 100.950 ;
        RECT 886.950 97.800 889.050 99.900 ;
        RECT 883.950 94.950 886.050 97.050 ;
        RECT 880.950 73.950 883.050 76.050 ;
        RECT 874.950 61.950 877.050 64.050 ;
        RECT 881.400 58.050 882.600 73.950 ;
        RECT 884.400 61.050 885.600 94.950 ;
        RECT 886.950 61.950 889.050 64.050 ;
        RECT 883.950 58.950 886.050 61.050 ;
        RECT 877.950 55.950 880.050 58.050 ;
        RECT 880.950 55.950 883.050 58.050 ;
        RECT 878.400 54.900 879.600 55.950 ;
        RECT 871.950 52.800 874.050 54.900 ;
        RECT 877.950 52.800 880.050 54.900 ;
        RECT 883.950 52.950 886.050 55.050 ;
        RECT 871.950 46.950 874.050 49.050 ;
        RECT 856.950 28.950 859.050 31.050 ;
        RECT 868.950 28.950 871.050 31.050 ;
        RECT 841.950 22.950 844.050 25.050 ;
        RECT 844.950 22.950 847.050 25.050 ;
        RECT 847.950 22.950 850.050 25.050 ;
        RECT 850.950 22.950 853.050 25.050 ;
        RECT 842.400 21.900 843.600 22.950 ;
        RECT 848.400 21.900 849.600 22.950 ;
        RECT 857.400 21.900 858.600 28.950 ;
        RECT 872.400 25.050 873.600 46.950 ;
        RECT 884.400 46.050 885.600 52.950 ;
        RECT 883.950 43.950 886.050 46.050 ;
        RECT 877.950 34.950 880.050 37.050 ;
        RECT 878.400 25.050 879.600 34.950 ;
        RECT 868.950 22.950 871.050 25.050 ;
        RECT 871.950 22.950 874.050 25.050 ;
        RECT 874.950 22.950 877.050 25.050 ;
        RECT 877.950 22.950 880.050 25.050 ;
        RECT 869.400 21.900 870.600 22.950 ;
        RECT 778.950 19.800 781.050 21.900 ;
        RECT 787.950 19.800 790.050 21.900 ;
        RECT 793.950 19.800 796.050 21.900 ;
        RECT 802.950 19.800 805.050 21.900 ;
        RECT 808.950 19.800 811.050 21.900 ;
        RECT 826.950 19.800 829.050 21.900 ;
        RECT 835.950 19.800 838.050 21.900 ;
        RECT 841.950 19.800 844.050 21.900 ;
        RECT 847.950 19.800 850.050 21.900 ;
        RECT 856.950 19.800 859.050 21.900 ;
        RECT 868.950 19.800 871.050 21.900 ;
        RECT 715.950 13.950 718.050 16.050 ;
        RECT 742.950 13.950 745.050 16.050 ;
        RECT 646.950 9.600 649.050 11.700 ;
        RECT 667.950 10.500 670.050 12.600 ;
        RECT 875.400 7.050 876.600 22.950 ;
        RECT 887.400 21.900 888.600 61.950 ;
        RECT 893.400 49.050 894.600 403.950 ;
        RECT 896.400 366.900 897.600 415.950 ;
        RECT 895.950 364.800 898.050 366.900 ;
        RECT 895.950 343.950 898.050 346.050 ;
        RECT 896.400 271.050 897.600 343.950 ;
        RECT 895.950 268.950 898.050 271.050 ;
        RECT 895.950 259.950 898.050 262.050 ;
        RECT 896.400 124.050 897.600 259.950 ;
        RECT 895.950 121.950 898.050 124.050 ;
        RECT 892.950 46.950 895.050 49.050 ;
        RECT 886.950 19.800 889.050 21.900 ;
        RECT 226.950 4.950 229.050 7.050 ;
        RECT 232.950 4.950 235.050 7.050 ;
        RECT 454.950 4.950 457.050 7.050 ;
        RECT 598.950 4.950 601.050 7.050 ;
        RECT 874.950 4.950 877.050 7.050 ;
      LAYER metal3 ;
        RECT 256.950 894.600 259.050 895.050 ;
        RECT 268.950 894.600 271.050 895.050 ;
        RECT 256.950 893.400 271.050 894.600 ;
        RECT 256.950 892.950 259.050 893.400 ;
        RECT 268.950 892.950 271.050 893.400 ;
        RECT 310.950 894.600 313.050 895.050 ;
        RECT 322.950 894.600 325.050 895.050 ;
        RECT 310.950 893.400 325.050 894.600 ;
        RECT 310.950 892.950 313.050 893.400 ;
        RECT 322.950 892.950 325.050 893.400 ;
        RECT 334.950 894.600 337.050 895.050 ;
        RECT 364.950 894.600 367.050 895.050 ;
        RECT 334.950 893.400 367.050 894.600 ;
        RECT 334.950 892.950 337.050 893.400 ;
        RECT 364.950 892.950 367.050 893.400 ;
        RECT 370.950 894.600 373.050 895.050 ;
        RECT 394.950 894.600 397.050 895.050 ;
        RECT 370.950 893.400 397.050 894.600 ;
        RECT 370.950 892.950 373.050 893.400 ;
        RECT 394.950 892.950 397.050 893.400 ;
        RECT 562.950 894.600 565.050 895.050 ;
        RECT 679.950 894.600 682.050 895.050 ;
        RECT 562.950 893.400 682.050 894.600 ;
        RECT 562.950 892.950 565.050 893.400 ;
        RECT 679.950 892.950 682.050 893.400 ;
        RECT 688.950 894.600 691.050 895.050 ;
        RECT 778.950 894.600 781.050 895.050 ;
        RECT 688.950 893.400 781.050 894.600 ;
        RECT 688.950 892.950 691.050 893.400 ;
        RECT 778.950 892.950 781.050 893.400 ;
        RECT 166.950 891.600 169.050 892.050 ;
        RECT 196.950 891.600 199.050 892.050 ;
        RECT 166.950 890.400 199.050 891.600 ;
        RECT 166.950 889.950 169.050 890.400 ;
        RECT 196.950 889.950 199.050 890.400 ;
        RECT 226.950 891.600 229.050 892.050 ;
        RECT 244.950 891.600 247.050 892.050 ;
        RECT 316.950 891.600 319.050 892.050 ;
        RECT 367.950 891.600 370.050 892.050 ;
        RECT 226.950 890.400 319.050 891.600 ;
        RECT 226.950 889.950 229.050 890.400 ;
        RECT 244.950 889.950 247.050 890.400 ;
        RECT 316.950 889.950 319.050 890.400 ;
        RECT 338.400 890.400 370.050 891.600 ;
        RECT 338.400 889.050 339.600 890.400 ;
        RECT 367.950 889.950 370.050 890.400 ;
        RECT 490.950 891.600 493.050 892.050 ;
        RECT 541.950 891.600 544.050 892.050 ;
        RECT 490.950 890.400 544.050 891.600 ;
        RECT 490.950 889.950 493.050 890.400 ;
        RECT 541.950 889.950 544.050 890.400 ;
        RECT 601.950 891.600 604.050 892.050 ;
        RECT 613.950 891.600 616.050 892.050 ;
        RECT 601.950 890.400 616.050 891.600 ;
        RECT 601.950 889.950 604.050 890.400 ;
        RECT 613.950 889.950 616.050 890.400 ;
        RECT 640.950 891.600 643.050 892.050 ;
        RECT 667.950 891.600 670.050 892.050 ;
        RECT 640.950 890.400 670.050 891.600 ;
        RECT 640.950 889.950 643.050 890.400 ;
        RECT 667.950 889.950 670.050 890.400 ;
        RECT 820.950 891.600 823.050 892.050 ;
        RECT 886.950 891.600 889.050 892.050 ;
        RECT 820.950 890.400 889.050 891.600 ;
        RECT 820.950 889.950 823.050 890.400 ;
        RECT 886.950 889.950 889.050 890.400 ;
        RECT 22.950 888.600 25.050 889.050 ;
        RECT 31.950 888.600 34.050 889.050 ;
        RECT 22.950 887.400 34.050 888.600 ;
        RECT 22.950 886.950 25.050 887.400 ;
        RECT 31.950 886.950 34.050 887.400 ;
        RECT 331.950 888.600 334.050 889.050 ;
        RECT 337.950 888.600 340.050 889.050 ;
        RECT 331.950 887.400 340.050 888.600 ;
        RECT 331.950 886.950 334.050 887.400 ;
        RECT 337.950 886.950 340.050 887.400 ;
        RECT 16.950 885.600 19.050 886.200 ;
        RECT 43.950 885.600 46.050 886.500 ;
        RECT 16.950 884.400 46.050 885.600 ;
        RECT 55.950 886.050 58.050 886.500 ;
        RECT 79.950 886.050 82.050 886.500 ;
        RECT 55.950 884.850 82.050 886.050 ;
        RECT 55.950 884.400 58.050 884.850 ;
        RECT 79.950 884.400 82.050 884.850 ;
        RECT 181.950 885.600 184.050 886.050 ;
        RECT 217.950 885.600 220.050 886.200 ;
        RECT 181.950 884.400 220.050 885.600 ;
        RECT 16.950 884.100 19.050 884.400 ;
        RECT 17.400 882.600 18.600 884.100 ;
        RECT 181.950 883.950 184.050 884.400 ;
        RECT 217.950 884.100 220.050 884.400 ;
        RECT 229.950 885.600 232.050 886.050 ;
        RECT 238.950 885.600 241.050 886.200 ;
        RECT 262.950 885.600 265.050 886.200 ;
        RECT 289.950 885.600 292.050 886.200 ;
        RECT 304.950 885.600 307.050 886.200 ;
        RECT 229.950 884.400 265.050 885.600 ;
        RECT 229.950 883.950 232.050 884.400 ;
        RECT 238.950 884.100 241.050 884.400 ;
        RECT 262.950 884.100 265.050 884.400 ;
        RECT 272.400 884.400 307.050 885.600 ;
        RECT 17.400 881.400 30.600 882.600 ;
        RECT 29.400 879.900 30.600 881.400 ;
        RECT 13.950 879.450 16.050 879.900 ;
        RECT 25.800 879.450 27.900 879.900 ;
        RECT 13.950 878.250 27.900 879.450 ;
        RECT 13.950 877.800 16.050 878.250 ;
        RECT 25.800 877.800 27.900 878.250 ;
        RECT 28.950 877.800 31.050 879.900 ;
        RECT 34.950 879.600 37.050 879.900 ;
        RECT 55.950 879.600 58.050 880.050 ;
        RECT 34.950 878.400 58.050 879.600 ;
        RECT 34.950 877.800 37.050 878.400 ;
        RECT 55.950 877.950 58.050 878.400 ;
        RECT 109.950 879.600 112.050 880.050 ;
        RECT 272.400 879.900 273.600 884.400 ;
        RECT 289.950 884.100 292.050 884.400 ;
        RECT 304.950 884.100 307.050 884.400 ;
        RECT 316.950 885.600 319.050 886.050 ;
        RECT 334.950 885.600 337.050 886.050 ;
        RECT 316.950 884.400 337.050 885.600 ;
        RECT 316.950 883.950 319.050 884.400 ;
        RECT 334.950 883.950 337.050 884.400 ;
        RECT 340.950 885.600 343.050 886.050 ;
        RECT 346.950 885.600 349.050 886.200 ;
        RECT 340.950 884.400 349.050 885.600 ;
        RECT 340.950 883.950 343.050 884.400 ;
        RECT 346.950 884.100 349.050 884.400 ;
        RECT 352.950 885.750 355.050 886.200 ;
        RECT 358.950 885.750 361.050 886.200 ;
        RECT 352.950 884.550 361.050 885.750 ;
        RECT 352.950 884.100 355.050 884.550 ;
        RECT 358.950 884.100 361.050 884.550 ;
        RECT 373.950 885.600 376.050 886.200 ;
        RECT 388.950 885.600 391.050 886.050 ;
        RECT 373.950 884.400 391.050 885.600 ;
        RECT 373.950 884.100 376.050 884.400 ;
        RECT 388.950 883.950 391.050 884.400 ;
        RECT 400.950 884.100 403.050 886.200 ;
        RECT 409.950 885.750 412.050 886.200 ;
        RECT 415.950 885.750 418.050 886.200 ;
        RECT 409.950 884.550 418.050 885.750 ;
        RECT 409.950 884.100 412.050 884.550 ;
        RECT 415.950 884.100 418.050 884.550 ;
        RECT 439.950 884.100 442.050 886.200 ;
        RECT 445.950 885.600 448.050 886.200 ;
        RECT 454.950 885.750 457.050 886.200 ;
        RECT 463.950 885.750 466.050 886.200 ;
        RECT 454.950 885.600 466.050 885.750 ;
        RECT 445.950 884.550 466.050 885.600 ;
        RECT 445.950 884.400 457.050 884.550 ;
        RECT 445.950 884.100 448.050 884.400 ;
        RECT 454.950 884.100 457.050 884.400 ;
        RECT 463.950 884.100 466.050 884.550 ;
        RECT 469.950 885.600 472.050 886.200 ;
        RECT 475.800 885.600 477.900 886.050 ;
        RECT 469.950 884.400 477.900 885.600 ;
        RECT 469.950 884.100 472.050 884.400 ;
        RECT 401.400 882.600 402.600 884.100 ;
        RECT 440.400 882.600 441.600 884.100 ;
        RECT 475.800 883.950 477.900 884.400 ;
        RECT 478.950 885.750 481.050 886.200 ;
        RECT 484.950 885.750 487.050 886.200 ;
        RECT 478.950 884.550 487.050 885.750 ;
        RECT 478.950 884.100 481.050 884.550 ;
        RECT 484.950 884.100 487.050 884.550 ;
        RECT 499.950 885.600 502.050 886.050 ;
        RECT 508.950 885.600 511.050 886.200 ;
        RECT 499.950 884.400 511.050 885.600 ;
        RECT 499.950 883.950 502.050 884.400 ;
        RECT 508.950 884.100 511.050 884.400 ;
        RECT 520.950 885.600 523.050 886.050 ;
        RECT 529.950 885.600 532.050 886.200 ;
        RECT 520.950 884.400 532.050 885.600 ;
        RECT 520.950 883.950 523.050 884.400 ;
        RECT 529.950 884.100 532.050 884.400 ;
        RECT 535.950 885.600 538.050 886.200 ;
        RECT 544.950 885.600 547.050 886.050 ;
        RECT 535.950 884.400 547.050 885.600 ;
        RECT 535.950 884.100 538.050 884.400 ;
        RECT 544.950 883.950 547.050 884.400 ;
        RECT 574.950 885.750 577.050 886.200 ;
        RECT 580.950 885.750 583.050 886.200 ;
        RECT 574.950 884.550 583.050 885.750 ;
        RECT 574.950 884.100 577.050 884.550 ;
        RECT 580.950 884.100 583.050 884.550 ;
        RECT 586.950 885.600 589.050 886.200 ;
        RECT 592.950 885.600 595.050 889.050 ;
        RECT 670.950 888.600 673.050 889.050 ;
        RECT 703.950 888.600 706.050 889.050 ;
        RECT 670.950 887.400 706.050 888.600 ;
        RECT 670.950 886.950 673.050 887.400 ;
        RECT 703.950 886.950 706.050 887.400 ;
        RECT 847.950 888.600 850.050 889.050 ;
        RECT 853.950 888.600 856.050 889.050 ;
        RECT 847.950 887.400 856.050 888.600 ;
        RECT 847.950 886.950 850.050 887.400 ;
        RECT 853.950 886.950 856.050 887.400 ;
        RECT 586.950 885.000 595.050 885.600 ;
        RECT 595.950 885.600 598.050 886.050 ;
        RECT 607.950 885.600 610.050 886.200 ;
        RECT 586.950 884.400 594.600 885.000 ;
        RECT 595.950 884.400 610.050 885.600 ;
        RECT 586.950 884.100 589.050 884.400 ;
        RECT 595.950 883.950 598.050 884.400 ;
        RECT 607.950 884.100 610.050 884.400 ;
        RECT 622.950 885.600 625.050 886.050 ;
        RECT 634.950 885.600 637.050 886.200 ;
        RECT 622.950 884.400 637.050 885.600 ;
        RECT 622.950 883.950 625.050 884.400 ;
        RECT 634.950 884.100 637.050 884.400 ;
        RECT 649.950 885.600 652.050 886.050 ;
        RECT 655.950 885.600 658.050 886.200 ;
        RECT 649.950 884.400 658.050 885.600 ;
        RECT 649.950 883.950 652.050 884.400 ;
        RECT 655.950 884.100 658.050 884.400 ;
        RECT 661.950 884.100 664.050 886.200 ;
        RECT 667.950 885.600 670.050 886.050 ;
        RECT 700.950 885.600 703.050 886.200 ;
        RECT 667.950 884.400 703.050 885.600 ;
        RECT 500.400 882.600 501.600 883.950 ;
        RECT 401.400 881.400 501.600 882.600 ;
        RECT 662.400 882.600 663.600 884.100 ;
        RECT 667.950 883.950 670.050 884.400 ;
        RECT 700.950 884.100 703.050 884.400 ;
        RECT 706.950 883.950 709.050 886.050 ;
        RECT 730.950 884.100 733.050 886.200 ;
        RECT 739.950 885.600 742.050 886.050 ;
        RECT 748.950 885.600 751.050 886.200 ;
        RECT 739.950 884.400 751.050 885.600 ;
        RECT 707.400 882.600 708.600 883.950 ;
        RECT 731.400 882.600 732.600 884.100 ;
        RECT 739.950 883.950 742.050 884.400 ;
        RECT 748.950 884.100 751.050 884.400 ;
        RECT 754.950 885.600 757.050 886.200 ;
        RECT 763.950 885.750 766.050 886.200 ;
        RECT 772.950 885.750 775.050 886.200 ;
        RECT 763.950 885.600 775.050 885.750 ;
        RECT 754.950 884.550 775.050 885.600 ;
        RECT 754.950 884.400 766.050 884.550 ;
        RECT 754.950 884.100 757.050 884.400 ;
        RECT 763.950 884.100 766.050 884.400 ;
        RECT 772.950 884.100 775.050 884.550 ;
        RECT 790.950 885.750 793.050 886.200 ;
        RECT 799.950 885.750 802.050 886.200 ;
        RECT 790.950 884.550 802.050 885.750 ;
        RECT 790.950 884.100 793.050 884.550 ;
        RECT 799.950 884.100 802.050 884.550 ;
        RECT 805.950 885.750 808.050 886.200 ;
        RECT 811.950 885.750 814.050 886.200 ;
        RECT 805.950 884.550 814.050 885.750 ;
        RECT 805.950 884.100 808.050 884.550 ;
        RECT 811.950 884.100 814.050 884.550 ;
        RECT 823.950 885.750 826.050 886.200 ;
        RECT 832.950 885.750 835.050 886.200 ;
        RECT 823.950 884.550 835.050 885.750 ;
        RECT 823.950 884.100 826.050 884.550 ;
        RECT 832.950 884.100 835.050 884.550 ;
        RECT 838.950 885.600 841.050 886.200 ;
        RECT 844.950 885.600 847.050 886.050 ;
        RECT 838.950 884.400 847.050 885.600 ;
        RECT 838.950 884.100 841.050 884.400 ;
        RECT 844.950 883.950 847.050 884.400 ;
        RECT 859.950 885.600 862.050 886.200 ;
        RECT 871.950 885.600 874.050 886.050 ;
        RECT 880.950 885.600 883.050 886.200 ;
        RECT 859.950 884.400 883.050 885.600 ;
        RECT 859.950 884.100 862.050 884.400 ;
        RECT 871.950 883.950 874.050 884.400 ;
        RECT 880.950 884.100 883.050 884.400 ;
        RECT 662.400 881.400 681.600 882.600 ;
        RECT 707.400 881.400 732.600 882.600 ;
        RECT 145.950 879.600 148.050 879.900 ;
        RECT 109.950 878.400 148.050 879.600 ;
        RECT 109.950 877.950 112.050 878.400 ;
        RECT 145.950 877.800 148.050 878.400 ;
        RECT 214.950 879.450 217.050 879.900 ;
        RECT 226.950 879.450 229.050 879.900 ;
        RECT 214.950 878.250 229.050 879.450 ;
        RECT 214.950 877.800 217.050 878.250 ;
        RECT 226.950 877.800 229.050 878.250 ;
        RECT 271.950 877.800 274.050 879.900 ;
        RECT 295.950 879.450 298.050 879.900 ;
        RECT 307.950 879.450 310.050 879.900 ;
        RECT 295.950 878.250 310.050 879.450 ;
        RECT 295.950 877.800 298.050 878.250 ;
        RECT 307.950 877.800 310.050 878.250 ;
        RECT 313.950 879.600 316.050 879.900 ;
        RECT 328.950 879.600 331.050 879.900 ;
        RECT 313.950 878.400 331.050 879.600 ;
        RECT 313.950 877.800 316.050 878.400 ;
        RECT 328.950 877.800 331.050 878.400 ;
        RECT 388.950 879.450 391.050 879.900 ;
        RECT 442.950 879.450 445.050 879.900 ;
        RECT 388.950 878.250 445.050 879.450 ;
        RECT 388.950 877.800 391.050 878.250 ;
        RECT 442.950 877.800 445.050 878.250 ;
        RECT 448.950 879.600 451.050 879.900 ;
        RECT 460.950 879.600 463.050 879.900 ;
        RECT 448.950 878.400 463.050 879.600 ;
        RECT 448.950 877.800 451.050 878.400 ;
        RECT 460.950 877.800 463.050 878.400 ;
        RECT 475.950 879.450 478.050 879.900 ;
        RECT 487.950 879.450 490.050 879.900 ;
        RECT 475.950 878.250 490.050 879.450 ;
        RECT 475.950 877.800 478.050 878.250 ;
        RECT 487.950 877.800 490.050 878.250 ;
        RECT 511.950 879.600 514.050 879.900 ;
        RECT 532.950 879.600 535.050 879.900 ;
        RECT 511.950 878.400 535.050 879.600 ;
        RECT 511.950 877.800 514.050 878.400 ;
        RECT 532.950 877.800 535.050 878.400 ;
        RECT 568.950 879.450 571.050 879.900 ;
        RECT 583.950 879.450 586.050 879.900 ;
        RECT 568.950 878.250 586.050 879.450 ;
        RECT 568.950 877.800 571.050 878.250 ;
        RECT 583.950 877.800 586.050 878.250 ;
        RECT 589.950 879.450 592.050 879.900 ;
        RECT 595.950 879.450 598.050 879.900 ;
        RECT 589.950 878.250 598.050 879.450 ;
        RECT 589.950 877.800 592.050 878.250 ;
        RECT 595.950 877.800 598.050 878.250 ;
        RECT 616.950 879.450 619.050 879.900 ;
        RECT 649.950 879.450 652.050 879.900 ;
        RECT 616.950 878.250 652.050 879.450 ;
        RECT 616.950 877.800 619.050 878.250 ;
        RECT 649.950 877.800 652.050 878.250 ;
        RECT 664.950 879.600 667.050 879.900 ;
        RECT 670.950 879.600 673.050 879.900 ;
        RECT 664.950 879.450 673.050 879.600 ;
        RECT 676.950 879.450 679.050 879.900 ;
        RECT 664.950 878.400 679.050 879.450 ;
        RECT 680.400 879.600 681.600 881.400 ;
        RECT 682.950 879.600 685.050 879.900 ;
        RECT 680.400 878.400 685.050 879.600 ;
        RECT 664.950 877.800 667.050 878.400 ;
        RECT 670.950 878.250 679.050 878.400 ;
        RECT 670.950 877.800 673.050 878.250 ;
        RECT 676.950 877.800 679.050 878.250 ;
        RECT 682.950 877.800 685.050 878.400 ;
        RECT 709.950 879.600 712.050 879.900 ;
        RECT 727.950 879.600 730.050 879.900 ;
        RECT 709.950 878.400 730.050 879.600 ;
        RECT 731.400 879.600 732.600 881.400 ;
        RECT 736.950 879.600 739.050 880.050 ;
        RECT 731.400 878.400 739.050 879.600 ;
        RECT 709.950 877.800 712.050 878.400 ;
        RECT 727.950 877.800 730.050 878.400 ;
        RECT 736.950 877.950 739.050 878.400 ;
        RECT 751.950 879.600 754.050 879.900 ;
        RECT 769.950 879.600 772.050 879.900 ;
        RECT 751.950 878.400 772.050 879.600 ;
        RECT 751.950 877.800 754.050 878.400 ;
        RECT 769.950 877.800 772.050 878.400 ;
        RECT 775.950 879.600 778.050 879.900 ;
        RECT 796.950 879.600 799.050 879.900 ;
        RECT 775.950 878.400 799.050 879.600 ;
        RECT 775.950 877.800 778.050 878.400 ;
        RECT 796.950 877.800 799.050 878.400 ;
        RECT 814.950 879.600 817.050 879.900 ;
        RECT 835.950 879.600 838.050 879.900 ;
        RECT 814.950 878.400 838.050 879.600 ;
        RECT 814.950 877.800 817.050 878.400 ;
        RECT 835.950 877.800 838.050 878.400 ;
        RECT 70.950 876.600 73.050 877.050 ;
        RECT 76.950 876.600 79.050 877.050 ;
        RECT 106.950 876.600 109.050 877.050 ;
        RECT 70.950 875.400 109.050 876.600 ;
        RECT 70.950 874.950 73.050 875.400 ;
        RECT 76.950 874.950 79.050 875.400 ;
        RECT 106.950 874.950 109.050 875.400 ;
        RECT 397.950 876.600 400.050 877.050 ;
        RECT 406.950 876.600 409.050 877.050 ;
        RECT 397.950 875.400 409.050 876.600 ;
        RECT 397.950 874.950 400.050 875.400 ;
        RECT 406.950 874.950 409.050 875.400 ;
        RECT 493.950 876.600 496.050 877.050 ;
        RECT 499.950 876.600 502.050 877.050 ;
        RECT 493.950 875.400 502.050 876.600 ;
        RECT 493.950 874.950 496.050 875.400 ;
        RECT 499.950 874.950 502.050 875.400 ;
        RECT 544.950 876.600 547.050 877.050 ;
        RECT 574.950 876.600 577.050 877.050 ;
        RECT 544.950 875.400 577.050 876.600 ;
        RECT 544.950 874.950 547.050 875.400 ;
        RECT 574.950 874.950 577.050 875.400 ;
        RECT 634.950 876.600 637.050 877.050 ;
        RECT 658.950 876.600 661.050 877.050 ;
        RECT 634.950 875.400 661.050 876.600 ;
        RECT 634.950 874.950 637.050 875.400 ;
        RECT 658.950 874.950 661.050 875.400 ;
        RECT 703.950 876.600 706.050 877.050 ;
        RECT 733.950 876.600 736.050 877.050 ;
        RECT 703.950 875.400 736.050 876.600 ;
        RECT 703.950 874.950 706.050 875.400 ;
        RECT 733.950 874.950 736.050 875.400 ;
        RECT 199.950 873.600 202.050 874.050 ;
        RECT 229.950 873.600 232.050 874.050 ;
        RECT 199.950 872.400 232.050 873.600 ;
        RECT 199.950 871.950 202.050 872.400 ;
        RECT 229.950 871.950 232.050 872.400 ;
        RECT 241.950 873.600 244.050 874.050 ;
        RECT 340.950 873.600 343.050 874.050 ;
        RECT 601.950 873.600 604.050 874.050 ;
        RECT 241.950 872.400 604.050 873.600 ;
        RECT 241.950 871.950 244.050 872.400 ;
        RECT 340.950 871.950 343.050 872.400 ;
        RECT 601.950 871.950 604.050 872.400 ;
        RECT 682.950 873.600 685.050 874.050 ;
        RECT 730.800 873.600 732.900 874.050 ;
        RECT 682.950 872.400 732.900 873.600 ;
        RECT 734.400 873.600 735.600 874.950 ;
        RECT 790.950 873.600 793.050 874.050 ;
        RECT 829.950 873.600 832.050 874.050 ;
        RECT 734.400 872.400 832.050 873.600 ;
        RECT 682.950 871.950 685.050 872.400 ;
        RECT 730.800 871.950 732.900 872.400 ;
        RECT 790.950 871.950 793.050 872.400 ;
        RECT 829.950 871.950 832.050 872.400 ;
        RECT 856.950 873.600 859.050 874.050 ;
        RECT 862.950 873.600 865.050 874.050 ;
        RECT 856.950 872.400 865.050 873.600 ;
        RECT 856.950 871.950 859.050 872.400 ;
        RECT 862.950 871.950 865.050 872.400 ;
        RECT 352.950 870.600 355.050 871.050 ;
        RECT 370.950 870.600 373.050 871.050 ;
        RECT 352.950 869.400 373.050 870.600 ;
        RECT 352.950 868.950 355.050 869.400 ;
        RECT 370.950 868.950 373.050 869.400 ;
        RECT 403.950 870.600 406.050 871.050 ;
        RECT 409.950 870.600 412.050 871.050 ;
        RECT 421.950 870.600 424.050 871.050 ;
        RECT 478.950 870.600 481.050 871.050 ;
        RECT 403.950 869.400 481.050 870.600 ;
        RECT 403.950 868.950 406.050 869.400 ;
        RECT 409.950 868.950 412.050 869.400 ;
        RECT 421.950 868.950 424.050 869.400 ;
        RECT 478.950 868.950 481.050 869.400 ;
        RECT 637.950 870.600 640.050 871.050 ;
        RECT 688.950 870.600 691.050 871.050 ;
        RECT 637.950 869.400 691.050 870.600 ;
        RECT 637.950 868.950 640.050 869.400 ;
        RECT 688.950 868.950 691.050 869.400 ;
        RECT 763.950 870.600 766.050 871.050 ;
        RECT 772.950 870.600 775.050 871.050 ;
        RECT 763.950 869.400 775.050 870.600 ;
        RECT 763.950 868.950 766.050 869.400 ;
        RECT 772.950 868.950 775.050 869.400 ;
        RECT 172.950 867.600 175.050 868.050 ;
        RECT 193.950 867.600 196.050 868.050 ;
        RECT 226.950 867.600 229.050 868.050 ;
        RECT 235.950 867.600 238.050 868.050 ;
        RECT 172.950 866.400 238.050 867.600 ;
        RECT 172.950 865.950 175.050 866.400 ;
        RECT 193.950 865.950 196.050 866.400 ;
        RECT 226.950 865.950 229.050 866.400 ;
        RECT 235.950 865.950 238.050 866.400 ;
        RECT 301.950 867.600 304.050 868.050 ;
        RECT 322.950 867.600 325.050 868.050 ;
        RECT 376.950 867.600 379.050 868.050 ;
        RECT 301.950 866.400 379.050 867.600 ;
        RECT 301.950 865.950 304.050 866.400 ;
        RECT 322.950 865.950 325.050 866.400 ;
        RECT 376.950 865.950 379.050 866.400 ;
        RECT 406.950 867.600 409.050 868.050 ;
        RECT 520.950 867.600 523.050 868.050 ;
        RECT 406.950 866.400 523.050 867.600 ;
        RECT 406.950 865.950 409.050 866.400 ;
        RECT 520.950 865.950 523.050 866.400 ;
        RECT 550.950 867.600 553.050 868.050 ;
        RECT 634.950 867.600 637.050 868.050 ;
        RECT 550.950 866.400 637.050 867.600 ;
        RECT 550.950 865.950 553.050 866.400 ;
        RECT 634.950 865.950 637.050 866.400 ;
        RECT 727.950 867.600 730.050 868.050 ;
        RECT 823.950 867.600 826.050 868.050 ;
        RECT 727.950 866.400 826.050 867.600 ;
        RECT 727.950 865.950 730.050 866.400 ;
        RECT 823.950 865.950 826.050 866.400 ;
        RECT 97.950 861.600 100.050 862.050 ;
        RECT 106.950 861.600 109.050 862.050 ;
        RECT 97.950 860.400 109.050 861.600 ;
        RECT 97.950 859.950 100.050 860.400 ;
        RECT 106.950 859.950 109.050 860.400 ;
        RECT 265.950 861.600 268.050 862.050 ;
        RECT 325.950 861.600 328.050 862.050 ;
        RECT 265.950 860.400 328.050 861.600 ;
        RECT 265.950 859.950 268.050 860.400 ;
        RECT 325.950 859.950 328.050 860.400 ;
        RECT 358.950 861.600 361.050 862.050 ;
        RECT 559.950 861.600 562.050 862.050 ;
        RECT 358.950 860.400 562.050 861.600 ;
        RECT 358.950 859.950 361.050 860.400 ;
        RECT 559.950 859.950 562.050 860.400 ;
        RECT 574.950 861.600 577.050 862.050 ;
        RECT 631.950 861.600 634.050 862.050 ;
        RECT 574.950 860.400 634.050 861.600 ;
        RECT 574.950 859.950 577.050 860.400 ;
        RECT 631.950 859.950 634.050 860.400 ;
        RECT 658.950 861.600 661.050 862.050 ;
        RECT 685.950 861.600 688.050 862.050 ;
        RECT 658.950 860.400 688.050 861.600 ;
        RECT 658.950 859.950 661.050 860.400 ;
        RECT 685.950 859.950 688.050 860.400 ;
        RECT 97.950 855.600 100.050 856.050 ;
        RECT 151.950 855.600 154.050 856.050 ;
        RECT 97.950 854.400 154.050 855.600 ;
        RECT 97.950 853.950 100.050 854.400 ;
        RECT 151.950 853.950 154.050 854.400 ;
        RECT 220.950 855.600 223.050 856.050 ;
        RECT 247.950 855.600 250.050 856.050 ;
        RECT 427.800 855.600 429.900 856.050 ;
        RECT 220.950 854.400 429.900 855.600 ;
        RECT 220.950 853.950 223.050 854.400 ;
        RECT 247.950 853.950 250.050 854.400 ;
        RECT 427.800 853.950 429.900 854.400 ;
        RECT 430.950 855.600 433.050 856.050 ;
        RECT 439.950 855.600 442.050 856.050 ;
        RECT 526.950 855.600 529.050 856.050 ;
        RECT 430.950 854.400 529.050 855.600 ;
        RECT 430.950 853.950 433.050 854.400 ;
        RECT 439.950 853.950 442.050 854.400 ;
        RECT 526.950 853.950 529.050 854.400 ;
        RECT 616.950 855.600 619.050 856.050 ;
        RECT 715.950 855.600 718.050 856.050 ;
        RECT 616.950 854.400 718.050 855.600 ;
        RECT 616.950 853.950 619.050 854.400 ;
        RECT 715.950 853.950 718.050 854.400 ;
        RECT 733.950 855.600 736.050 856.050 ;
        RECT 793.950 855.600 796.050 856.050 ;
        RECT 805.950 855.600 808.050 856.050 ;
        RECT 733.950 854.400 808.050 855.600 ;
        RECT 733.950 853.950 736.050 854.400 ;
        RECT 793.950 853.950 796.050 854.400 ;
        RECT 805.950 853.950 808.050 854.400 ;
        RECT 160.950 852.600 163.050 853.050 ;
        RECT 169.950 852.600 172.050 853.050 ;
        RECT 160.950 851.400 172.050 852.600 ;
        RECT 160.950 850.950 163.050 851.400 ;
        RECT 169.950 850.950 172.050 851.400 ;
        RECT 223.950 852.600 226.050 853.050 ;
        RECT 349.950 852.600 352.050 853.050 ;
        RECT 223.950 851.400 352.050 852.600 ;
        RECT 223.950 850.950 226.050 851.400 ;
        RECT 349.950 850.950 352.050 851.400 ;
        RECT 463.950 852.600 466.050 853.050 ;
        RECT 544.950 852.600 547.050 853.050 ;
        RECT 463.950 851.400 547.050 852.600 ;
        RECT 463.950 850.950 466.050 851.400 ;
        RECT 544.950 850.950 547.050 851.400 ;
        RECT 559.950 852.600 562.050 853.050 ;
        RECT 607.950 852.600 610.050 853.050 ;
        RECT 559.950 851.400 610.050 852.600 ;
        RECT 559.950 850.950 562.050 851.400 ;
        RECT 607.950 850.950 610.050 851.400 ;
        RECT 148.950 849.600 151.050 850.050 ;
        RECT 595.950 849.600 598.050 850.050 ;
        RECT 148.950 848.400 598.050 849.600 ;
        RECT 148.950 847.950 151.050 848.400 ;
        RECT 595.950 847.950 598.050 848.400 ;
        RECT 835.950 849.600 838.050 850.050 ;
        RECT 844.950 849.600 847.050 850.050 ;
        RECT 835.950 848.400 847.050 849.600 ;
        RECT 835.950 847.950 838.050 848.400 ;
        RECT 844.950 847.950 847.050 848.400 ;
        RECT 151.950 846.600 154.050 847.050 ;
        RECT 223.950 846.600 226.050 847.050 ;
        RECT 151.950 845.400 226.050 846.600 ;
        RECT 151.950 844.950 154.050 845.400 ;
        RECT 223.950 844.950 226.050 845.400 ;
        RECT 268.950 846.600 271.050 847.050 ;
        RECT 286.800 846.600 288.900 847.050 ;
        RECT 268.950 845.400 288.900 846.600 ;
        RECT 268.950 844.950 271.050 845.400 ;
        RECT 286.800 844.950 288.900 845.400 ;
        RECT 289.950 846.600 292.050 847.050 ;
        RECT 313.950 846.600 316.050 847.050 ;
        RECT 319.950 846.600 322.050 847.050 ;
        RECT 289.950 845.400 322.050 846.600 ;
        RECT 289.950 844.950 292.050 845.400 ;
        RECT 313.950 844.950 316.050 845.400 ;
        RECT 319.950 844.950 322.050 845.400 ;
        RECT 367.950 846.600 370.050 847.050 ;
        RECT 385.950 846.600 388.050 847.050 ;
        RECT 394.950 846.600 397.050 847.050 ;
        RECT 367.950 845.400 397.050 846.600 ;
        RECT 367.950 844.950 370.050 845.400 ;
        RECT 385.950 844.950 388.050 845.400 ;
        RECT 394.950 844.950 397.050 845.400 ;
        RECT 433.950 846.600 436.050 847.050 ;
        RECT 469.950 846.600 472.050 847.050 ;
        RECT 433.950 845.400 472.050 846.600 ;
        RECT 433.950 844.950 436.050 845.400 ;
        RECT 469.950 844.950 472.050 845.400 ;
        RECT 484.950 846.600 487.050 847.050 ;
        RECT 502.950 846.600 505.050 847.050 ;
        RECT 514.950 846.600 517.050 847.050 ;
        RECT 484.950 845.400 517.050 846.600 ;
        RECT 484.950 844.950 487.050 845.400 ;
        RECT 502.950 844.950 505.050 845.400 ;
        RECT 514.950 844.950 517.050 845.400 ;
        RECT 541.950 846.600 544.050 847.050 ;
        RECT 553.950 846.600 556.050 847.050 ;
        RECT 541.950 845.400 556.050 846.600 ;
        RECT 541.950 844.950 544.050 845.400 ;
        RECT 553.950 844.950 556.050 845.400 ;
        RECT 724.950 846.600 727.050 847.050 ;
        RECT 799.950 846.600 802.050 847.050 ;
        RECT 724.950 845.400 802.050 846.600 ;
        RECT 724.950 844.950 727.050 845.400 ;
        RECT 799.950 844.950 802.050 845.400 ;
        RECT 871.950 844.050 874.050 844.200 ;
        RECT 76.950 843.600 79.050 844.050 ;
        RECT 82.950 843.600 85.050 844.050 ;
        RECT 76.950 842.400 85.050 843.600 ;
        RECT 76.950 841.950 79.050 842.400 ;
        RECT 82.950 841.950 85.050 842.400 ;
        RECT 124.950 843.600 127.050 844.050 ;
        RECT 133.950 843.600 136.050 844.050 ;
        RECT 124.950 842.400 136.050 843.600 ;
        RECT 124.950 841.950 127.050 842.400 ;
        RECT 133.950 841.950 136.050 842.400 ;
        RECT 313.950 843.600 316.050 843.900 ;
        RECT 322.950 843.600 325.050 844.050 ;
        RECT 334.950 843.600 337.050 844.050 ;
        RECT 349.950 843.600 352.050 844.050 ;
        RECT 313.950 842.400 333.600 843.600 ;
        RECT 313.950 841.800 316.050 842.400 ;
        RECT 322.950 841.950 325.050 842.400 ;
        RECT 10.950 839.100 13.050 841.200 ;
        RECT 19.800 840.600 21.900 841.200 ;
        RECT 14.250 839.400 21.900 840.600 ;
        RECT 11.400 837.600 12.600 839.100 ;
        RECT 8.400 837.000 12.600 837.600 ;
        RECT 7.950 836.400 12.600 837.000 ;
        RECT 7.950 832.950 10.050 836.400 ;
        RECT 14.250 835.050 15.450 839.400 ;
        RECT 19.800 839.100 21.900 839.400 ;
        RECT 22.950 840.600 25.050 841.050 ;
        RECT 28.950 840.600 31.050 841.050 ;
        RECT 22.950 839.400 31.050 840.600 ;
        RECT 22.950 838.950 25.050 839.400 ;
        RECT 28.950 838.950 31.050 839.400 ;
        RECT 37.950 839.100 40.050 841.200 ;
        RECT 64.950 839.400 67.050 841.500 ;
        RECT 91.950 840.600 94.050 841.200 ;
        RECT 109.950 840.750 112.050 841.200 ;
        RECT 118.950 840.750 121.050 841.200 ;
        RECT 109.950 840.600 121.050 840.750 ;
        RECT 142.950 840.600 145.050 841.200 ;
        RECT 166.950 840.600 169.050 841.200 ;
        RECT 91.950 839.550 169.050 840.600 ;
        RECT 91.950 839.400 112.050 839.550 ;
        RECT 13.800 832.950 15.900 835.050 ;
        RECT 16.950 834.450 19.050 834.900 ;
        RECT 22.950 834.450 25.050 835.050 ;
        RECT 28.950 834.450 31.050 834.900 ;
        RECT 16.950 833.250 31.050 834.450 ;
        RECT 38.400 834.600 39.600 839.100 ;
        RECT 43.950 834.600 46.050 835.050 ;
        RECT 38.400 833.400 46.050 834.600 ;
        RECT 65.400 834.600 66.600 839.400 ;
        RECT 91.950 839.100 94.050 839.400 ;
        RECT 109.950 839.100 112.050 839.400 ;
        RECT 118.950 839.400 169.050 839.550 ;
        RECT 118.950 839.100 121.050 839.400 ;
        RECT 142.950 839.100 145.050 839.400 ;
        RECT 166.950 839.100 169.050 839.400 ;
        RECT 193.950 839.100 196.050 841.200 ;
        RECT 199.950 840.600 202.050 841.200 ;
        RECT 211.950 840.600 214.050 841.200 ;
        RECT 199.950 839.400 214.050 840.600 ;
        RECT 199.950 839.100 202.050 839.400 ;
        RECT 211.950 839.100 214.050 839.400 ;
        RECT 217.950 839.100 220.050 841.200 ;
        RECT 229.950 840.750 232.050 841.200 ;
        RECT 235.950 840.750 238.050 841.200 ;
        RECT 229.950 839.550 238.050 840.750 ;
        RECT 229.950 839.100 232.050 839.550 ;
        RECT 235.950 839.100 238.050 839.550 ;
        RECT 241.950 840.750 244.050 841.200 ;
        RECT 250.950 840.750 253.050 841.200 ;
        RECT 241.950 839.550 253.050 840.750 ;
        RECT 241.950 839.100 244.050 839.550 ;
        RECT 250.950 839.100 253.050 839.550 ;
        RECT 280.950 840.750 283.050 841.200 ;
        RECT 295.950 840.750 298.050 841.200 ;
        RECT 280.950 840.600 298.050 840.750 ;
        RECT 307.950 840.600 310.050 841.200 ;
        RECT 319.950 840.600 322.050 841.050 ;
        RECT 280.950 839.550 310.050 840.600 ;
        RECT 280.950 839.100 283.050 839.550 ;
        RECT 295.950 839.400 310.050 839.550 ;
        RECT 295.950 839.100 298.050 839.400 ;
        RECT 307.950 839.100 310.050 839.400 ;
        RECT 311.400 839.400 322.050 840.600 ;
        RECT 332.400 840.600 333.600 842.400 ;
        RECT 334.950 842.400 352.050 843.600 ;
        RECT 334.950 841.950 337.050 842.400 ;
        RECT 349.950 841.950 352.050 842.400 ;
        RECT 397.950 843.600 400.050 844.050 ;
        RECT 412.950 843.600 415.050 844.050 ;
        RECT 397.950 842.400 415.050 843.600 ;
        RECT 397.950 841.950 400.050 842.400 ;
        RECT 412.950 841.950 415.050 842.400 ;
        RECT 634.950 843.600 637.050 844.050 ;
        RECT 640.950 843.600 643.050 844.050 ;
        RECT 667.950 843.600 670.050 844.050 ;
        RECT 634.950 842.400 670.050 843.600 ;
        RECT 634.950 841.950 637.050 842.400 ;
        RECT 640.950 841.950 643.050 842.400 ;
        RECT 667.950 841.950 670.050 842.400 ;
        RECT 685.950 843.600 688.050 844.050 ;
        RECT 691.950 843.600 694.050 844.050 ;
        RECT 870.000 843.600 874.050 844.050 ;
        RECT 685.950 842.400 694.050 843.600 ;
        RECT 685.950 841.950 688.050 842.400 ;
        RECT 691.950 841.950 694.050 842.400 ;
        RECT 869.400 842.100 874.050 843.600 ;
        RECT 869.400 841.950 873.000 842.100 ;
        RECT 340.950 840.600 343.050 841.200 ;
        RECT 332.400 839.400 343.050 840.600 ;
        RECT 184.950 837.600 187.050 838.050 ;
        RECT 194.400 837.600 195.600 839.100 ;
        RECT 184.950 836.400 195.600 837.600 ;
        RECT 205.950 837.600 208.050 838.050 ;
        RECT 218.400 837.600 219.600 839.100 ;
        RECT 205.950 836.400 219.600 837.600 ;
        RECT 184.950 835.950 187.050 836.400 ;
        RECT 205.950 835.950 208.050 836.400 ;
        RECT 94.950 834.600 97.050 834.900 ;
        RECT 65.400 833.400 97.050 834.600 ;
        RECT 16.950 832.800 19.050 833.250 ;
        RECT 22.950 832.950 25.050 833.250 ;
        RECT 28.950 832.800 31.050 833.250 ;
        RECT 43.950 832.950 46.050 833.400 ;
        RECT 94.950 832.800 97.050 833.400 ;
        RECT 106.950 834.450 109.050 834.900 ;
        RECT 121.950 834.450 124.050 834.900 ;
        RECT 106.950 833.250 124.050 834.450 ;
        RECT 106.950 832.800 109.050 833.250 ;
        RECT 121.950 832.800 124.050 833.250 ;
        RECT 196.950 834.600 199.050 834.900 ;
        RECT 214.950 834.600 217.050 834.900 ;
        RECT 196.950 833.400 217.050 834.600 ;
        RECT 196.950 832.800 199.050 833.400 ;
        RECT 214.950 832.800 217.050 833.400 ;
        RECT 220.950 834.600 223.050 834.900 ;
        RECT 226.950 834.600 229.050 835.050 ;
        RECT 220.950 833.400 229.050 834.600 ;
        RECT 220.950 832.800 223.050 833.400 ;
        RECT 226.950 832.950 229.050 833.400 ;
        RECT 244.950 834.600 247.050 834.900 ;
        RECT 253.950 834.600 256.050 835.050 ;
        RECT 311.400 834.900 312.600 839.400 ;
        RECT 319.950 838.950 322.050 839.400 ;
        RECT 340.950 839.100 343.050 839.400 ;
        RECT 376.950 837.600 379.050 841.050 ;
        RECT 406.950 839.100 409.050 841.200 ;
        RECT 376.950 837.000 387.600 837.600 ;
        RECT 377.400 836.400 387.600 837.000 ;
        RECT 244.950 833.400 256.050 834.600 ;
        RECT 244.950 832.800 247.050 833.400 ;
        RECT 253.950 832.950 256.050 833.400 ;
        RECT 271.950 834.600 274.050 834.900 ;
        RECT 286.950 834.600 289.050 834.900 ;
        RECT 271.950 833.400 289.050 834.600 ;
        RECT 271.950 832.800 274.050 833.400 ;
        RECT 286.950 832.800 289.050 833.400 ;
        RECT 292.950 834.450 295.050 834.900 ;
        RECT 301.950 834.450 304.050 834.900 ;
        RECT 292.950 833.250 304.050 834.450 ;
        RECT 292.950 832.800 295.050 833.250 ;
        RECT 301.950 832.800 304.050 833.250 ;
        RECT 310.950 832.800 313.050 834.900 ;
        RECT 325.950 834.600 328.050 835.050 ;
        RECT 337.950 834.600 340.050 834.900 ;
        RECT 325.950 833.400 340.050 834.600 ;
        RECT 325.950 832.950 328.050 833.400 ;
        RECT 337.950 832.800 340.050 833.400 ;
        RECT 343.950 834.600 346.050 834.900 ;
        RECT 352.950 834.600 355.050 835.050 ;
        RECT 358.950 834.600 361.050 834.900 ;
        RECT 343.950 833.400 361.050 834.600 ;
        RECT 343.950 832.800 346.050 833.400 ;
        RECT 352.950 832.950 355.050 833.400 ;
        RECT 358.950 832.800 361.050 833.400 ;
        RECT 370.950 834.450 373.050 834.900 ;
        RECT 382.950 834.450 385.050 834.900 ;
        RECT 370.950 833.250 385.050 834.450 ;
        RECT 386.400 834.600 387.600 836.400 ;
        RECT 388.950 834.600 391.050 834.900 ;
        RECT 386.400 833.400 391.050 834.600 ;
        RECT 370.950 832.800 373.050 833.250 ;
        RECT 382.950 832.800 385.050 833.250 ;
        RECT 388.950 832.800 391.050 833.400 ;
        RECT 400.950 834.600 403.050 835.050 ;
        RECT 407.400 834.600 408.600 839.100 ;
        RECT 427.950 838.950 430.050 841.050 ;
        RECT 445.950 840.750 448.050 841.200 ;
        RECT 457.950 840.750 460.050 841.200 ;
        RECT 445.950 839.550 460.050 840.750 ;
        RECT 445.950 839.100 448.050 839.550 ;
        RECT 457.950 839.100 460.050 839.550 ;
        RECT 466.950 840.750 469.050 841.200 ;
        RECT 478.950 840.750 481.050 841.200 ;
        RECT 466.950 839.550 481.050 840.750 ;
        RECT 466.950 839.100 469.050 839.550 ;
        RECT 478.950 839.100 481.050 839.550 ;
        RECT 493.950 840.750 496.050 841.200 ;
        RECT 508.950 840.750 511.050 841.200 ;
        RECT 493.950 839.550 511.050 840.750 ;
        RECT 493.950 839.100 496.050 839.550 ;
        RECT 508.950 839.100 511.050 839.550 ;
        RECT 529.950 839.100 532.050 841.200 ;
        RECT 535.950 840.750 538.050 841.200 ;
        RECT 541.950 840.750 544.050 841.200 ;
        RECT 535.950 839.550 544.050 840.750 ;
        RECT 535.950 839.100 538.050 839.550 ;
        RECT 541.950 839.100 544.050 839.550 ;
        RECT 559.950 839.100 562.050 841.200 ;
        RECT 595.950 840.750 598.050 841.200 ;
        RECT 628.950 840.750 631.050 841.200 ;
        RECT 595.950 839.550 631.050 840.750 ;
        RECT 595.950 839.100 598.050 839.550 ;
        RECT 628.950 839.100 631.050 839.550 ;
        RECT 679.950 840.600 682.050 841.200 ;
        RECT 697.950 840.600 700.050 841.200 ;
        RECT 724.950 840.600 727.050 841.200 ;
        RECT 679.950 839.400 727.050 840.600 ;
        RECT 679.950 839.100 682.050 839.400 ;
        RECT 697.950 839.100 700.050 839.400 ;
        RECT 724.950 839.100 727.050 839.400 ;
        RECT 748.950 839.100 751.050 841.200 ;
        RECT 754.950 840.750 757.050 841.200 ;
        RECT 760.950 840.750 763.050 841.200 ;
        RECT 754.950 839.550 763.050 840.750 ;
        RECT 754.950 839.100 757.050 839.550 ;
        RECT 760.950 839.100 763.050 839.550 ;
        RECT 766.950 839.100 769.050 841.200 ;
        RECT 787.950 840.600 790.050 841.200 ;
        RECT 773.400 839.400 790.050 840.600 ;
        RECT 400.950 833.400 408.600 834.600 ;
        RECT 428.400 834.600 429.600 838.950 ;
        RECT 430.950 834.600 433.050 834.900 ;
        RECT 428.400 833.400 433.050 834.600 ;
        RECT 400.950 832.950 403.050 833.400 ;
        RECT 430.950 832.800 433.050 833.400 ;
        RECT 436.950 834.450 439.050 834.900 ;
        RECT 442.950 834.450 445.050 834.900 ;
        RECT 436.950 833.250 445.050 834.450 ;
        RECT 436.950 832.800 439.050 833.250 ;
        RECT 442.950 832.800 445.050 833.250 ;
        RECT 469.950 834.600 472.050 835.050 ;
        RECT 481.950 834.600 484.050 834.900 ;
        RECT 469.950 833.400 484.050 834.600 ;
        RECT 469.950 832.950 472.050 833.400 ;
        RECT 481.950 832.800 484.050 833.400 ;
        RECT 514.950 834.600 517.050 835.050 ;
        RECT 526.950 834.600 529.050 834.900 ;
        RECT 514.950 833.400 529.050 834.600 ;
        RECT 530.400 834.600 531.600 839.100 ;
        RECT 560.400 835.050 561.600 839.100 ;
        RECT 664.950 837.600 667.050 838.050 ;
        RECT 656.400 836.400 667.050 837.600 ;
        RECT 749.400 837.600 750.600 839.100 ;
        RECT 749.400 836.400 753.600 837.600 ;
        RECT 538.950 834.600 541.050 835.050 ;
        RECT 530.400 833.400 541.050 834.600 ;
        RECT 514.950 832.950 517.050 833.400 ;
        RECT 526.950 832.800 529.050 833.400 ;
        RECT 538.950 832.950 541.050 833.400 ;
        RECT 544.950 834.600 547.050 835.050 ;
        RECT 550.950 834.600 553.050 834.900 ;
        RECT 544.950 833.400 553.050 834.600 ;
        RECT 560.400 833.400 564.900 835.050 ;
        RECT 544.950 832.950 547.050 833.400 ;
        RECT 550.950 832.800 553.050 833.400 ;
        RECT 561.000 832.950 564.900 833.400 ;
        RECT 565.950 834.600 568.050 835.050 ;
        RECT 622.950 834.600 625.050 835.050 ;
        RECT 656.400 834.900 657.600 836.400 ;
        RECT 664.950 835.950 667.050 836.400 ;
        RECT 565.950 833.400 625.050 834.600 ;
        RECT 565.950 832.950 568.050 833.400 ;
        RECT 622.950 832.950 625.050 833.400 ;
        RECT 655.950 832.800 658.050 834.900 ;
        RECT 667.950 834.600 670.050 835.050 ;
        RECT 676.950 834.600 679.050 834.900 ;
        RECT 667.950 833.400 679.050 834.600 ;
        RECT 667.950 832.950 670.050 833.400 ;
        RECT 676.950 832.800 679.050 833.400 ;
        RECT 685.950 834.600 688.050 835.050 ;
        RECT 733.950 834.600 736.050 835.050 ;
        RECT 739.950 834.600 742.050 834.900 ;
        RECT 685.950 833.400 693.600 834.600 ;
        RECT 685.950 832.950 688.050 833.400 ;
        RECT 37.950 831.600 40.050 832.050 ;
        RECT 46.950 831.600 49.050 832.050 ;
        RECT 37.950 830.400 49.050 831.600 ;
        RECT 37.950 829.950 40.050 830.400 ;
        RECT 46.950 829.950 49.050 830.400 ;
        RECT 100.950 831.600 103.050 832.050 ;
        RECT 145.950 831.600 148.050 832.050 ;
        RECT 100.950 830.400 148.050 831.600 ;
        RECT 100.950 829.950 103.050 830.400 ;
        RECT 145.950 829.950 148.050 830.400 ;
        RECT 229.950 831.600 232.050 832.050 ;
        RECT 238.950 831.600 241.050 832.050 ;
        RECT 229.950 830.400 241.050 831.600 ;
        RECT 229.950 829.950 232.050 830.400 ;
        RECT 238.950 829.950 241.050 830.400 ;
        RECT 397.950 831.600 400.050 832.050 ;
        RECT 406.950 831.600 409.050 832.050 ;
        RECT 397.950 830.400 409.050 831.600 ;
        RECT 397.950 829.950 400.050 830.400 ;
        RECT 406.950 829.950 409.050 830.400 ;
        RECT 448.950 831.600 453.000 832.050 ;
        RECT 460.950 831.600 463.050 832.050 ;
        RECT 448.950 830.400 463.050 831.600 ;
        RECT 448.950 829.950 453.600 830.400 ;
        RECT 460.950 829.950 463.050 830.400 ;
        RECT 505.950 831.600 508.050 832.050 ;
        RECT 511.950 831.600 514.050 832.050 ;
        RECT 505.950 830.400 514.050 831.600 ;
        RECT 505.950 829.950 508.050 830.400 ;
        RECT 511.950 829.950 514.050 830.400 ;
        RECT 565.950 831.600 568.050 831.900 ;
        RECT 580.950 831.600 583.050 832.050 ;
        RECT 565.950 830.400 583.050 831.600 ;
        RECT 13.950 828.600 16.050 829.050 ;
        RECT 19.950 828.600 22.050 829.050 ;
        RECT 13.950 827.400 22.050 828.600 ;
        RECT 13.950 826.950 16.050 827.400 ;
        RECT 19.950 826.950 22.050 827.400 ;
        RECT 148.950 828.600 151.050 829.050 ;
        RECT 184.950 828.600 187.050 829.050 ;
        RECT 205.950 828.600 208.050 829.050 ;
        RECT 148.950 827.400 208.050 828.600 ;
        RECT 148.950 826.950 151.050 827.400 ;
        RECT 184.950 826.950 187.050 827.400 ;
        RECT 205.950 826.950 208.050 827.400 ;
        RECT 214.950 828.600 217.050 829.050 ;
        RECT 265.950 828.600 268.050 829.050 ;
        RECT 214.950 827.400 268.050 828.600 ;
        RECT 214.950 826.950 217.050 827.400 ;
        RECT 265.950 826.950 268.050 827.400 ;
        RECT 394.950 828.600 397.050 829.050 ;
        RECT 409.950 828.600 412.050 829.050 ;
        RECT 394.950 827.400 412.050 828.600 ;
        RECT 394.950 826.950 397.050 827.400 ;
        RECT 409.950 826.950 412.050 827.400 ;
        RECT 439.950 828.600 442.050 829.050 ;
        RECT 452.400 828.600 453.600 829.950 ;
        RECT 565.950 829.800 568.050 830.400 ;
        RECT 580.950 829.950 583.050 830.400 ;
        RECT 604.950 831.600 607.050 832.050 ;
        RECT 616.950 831.600 619.050 832.050 ;
        RECT 604.950 830.400 619.050 831.600 ;
        RECT 692.400 831.600 693.600 833.400 ;
        RECT 733.950 833.400 742.050 834.600 ;
        RECT 752.400 834.600 753.600 836.400 ;
        RECT 763.950 834.600 766.050 834.900 ;
        RECT 752.400 833.400 766.050 834.600 ;
        RECT 733.950 832.950 736.050 833.400 ;
        RECT 739.950 832.800 742.050 833.400 ;
        RECT 763.950 832.800 766.050 833.400 ;
        RECT 767.400 832.050 768.600 839.100 ;
        RECT 773.400 837.600 774.600 839.400 ;
        RECT 787.950 839.100 790.050 839.400 ;
        RECT 808.950 839.100 811.050 841.200 ;
        RECT 814.950 840.750 817.050 841.200 ;
        RECT 820.950 840.750 823.050 841.200 ;
        RECT 814.950 839.550 823.050 840.750 ;
        RECT 814.950 839.100 817.050 839.550 ;
        RECT 820.950 839.100 823.050 839.550 ;
        RECT 841.950 839.100 844.050 841.200 ;
        RECT 809.400 837.600 810.600 839.100 ;
        RECT 770.400 836.400 774.600 837.600 ;
        RECT 797.400 836.400 810.600 837.600 ;
        RECT 770.400 834.900 771.600 836.400 ;
        RECT 769.950 832.800 772.050 834.900 ;
        RECT 775.950 834.450 778.050 835.050 ;
        RECT 784.950 834.450 787.050 834.900 ;
        RECT 775.950 833.250 787.050 834.450 ;
        RECT 775.950 832.950 778.050 833.250 ;
        RECT 784.950 832.800 787.050 833.250 ;
        RECT 790.950 834.600 793.050 834.900 ;
        RECT 797.400 834.600 798.600 836.400 ;
        RECT 790.950 833.400 798.600 834.600 ;
        RECT 799.950 834.600 802.050 835.050 ;
        RECT 838.950 834.600 841.050 834.900 ;
        RECT 799.950 833.400 841.050 834.600 ;
        RECT 842.400 834.600 843.600 839.100 ;
        RECT 869.400 834.900 870.600 841.950 ;
        RECT 871.950 840.600 874.050 841.050 ;
        RECT 883.950 840.600 886.050 841.050 ;
        RECT 892.950 840.600 895.050 841.050 ;
        RECT 871.950 839.400 895.050 840.600 ;
        RECT 871.950 838.950 874.050 839.400 ;
        RECT 883.950 838.950 886.050 839.400 ;
        RECT 892.950 838.950 895.050 839.400 ;
        RECT 862.950 834.600 865.050 834.900 ;
        RECT 842.400 833.400 865.050 834.600 ;
        RECT 790.950 832.800 793.050 833.400 ;
        RECT 799.950 832.950 802.050 833.400 ;
        RECT 838.950 832.800 841.050 833.400 ;
        RECT 862.950 832.800 865.050 833.400 ;
        RECT 868.950 832.800 871.050 834.900 ;
        RECT 706.950 831.600 709.050 831.900 ;
        RECT 692.400 830.400 709.050 831.600 ;
        RECT 604.950 829.950 607.050 830.400 ;
        RECT 616.950 829.950 619.050 830.400 ;
        RECT 706.950 829.800 709.050 830.400 ;
        RECT 766.950 829.950 769.050 832.050 ;
        RECT 439.950 827.400 453.600 828.600 ;
        RECT 463.950 828.600 466.050 829.050 ;
        RECT 487.950 828.600 490.050 829.050 ;
        RECT 499.950 828.600 502.050 829.050 ;
        RECT 463.950 827.400 502.050 828.600 ;
        RECT 439.950 826.950 442.050 827.400 ;
        RECT 463.950 826.950 466.050 827.400 ;
        RECT 487.950 826.950 490.050 827.400 ;
        RECT 499.950 826.950 502.050 827.400 ;
        RECT 532.950 828.600 535.050 829.050 ;
        RECT 556.950 828.600 559.050 829.050 ;
        RECT 628.950 828.600 631.050 829.050 ;
        RECT 532.950 827.400 631.050 828.600 ;
        RECT 532.950 826.950 535.050 827.400 ;
        RECT 556.950 826.950 559.050 827.400 ;
        RECT 628.950 826.950 631.050 827.400 ;
        RECT 748.950 828.600 751.050 829.050 ;
        RECT 754.950 828.600 757.050 829.050 ;
        RECT 748.950 827.400 757.050 828.600 ;
        RECT 748.950 826.950 751.050 827.400 ;
        RECT 754.950 826.950 757.050 827.400 ;
        RECT 7.950 825.600 10.050 826.050 ;
        RECT 13.950 825.600 16.050 825.900 ;
        RECT 7.950 824.400 16.050 825.600 ;
        RECT 7.950 823.950 10.050 824.400 ;
        RECT 13.950 823.800 16.050 824.400 ;
        RECT 40.950 825.600 43.050 826.050 ;
        RECT 88.950 825.600 91.050 826.050 ;
        RECT 40.950 824.400 91.050 825.600 ;
        RECT 40.950 823.950 43.050 824.400 ;
        RECT 88.950 823.950 91.050 824.400 ;
        RECT 133.950 825.600 136.050 826.050 ;
        RECT 169.950 825.600 172.050 826.050 ;
        RECT 133.950 824.400 172.050 825.600 ;
        RECT 133.950 823.950 136.050 824.400 ;
        RECT 169.950 823.950 172.050 824.400 ;
        RECT 316.950 825.600 319.050 826.050 ;
        RECT 445.950 825.600 448.050 826.050 ;
        RECT 316.950 824.400 448.050 825.600 ;
        RECT 316.950 823.950 319.050 824.400 ;
        RECT 445.950 823.950 448.050 824.400 ;
        RECT 535.950 825.600 538.050 826.050 ;
        RECT 565.950 825.600 568.050 826.050 ;
        RECT 535.950 824.400 568.050 825.600 ;
        RECT 535.950 823.950 538.050 824.400 ;
        RECT 565.950 823.950 568.050 824.400 ;
        RECT 571.950 825.600 574.050 826.050 ;
        RECT 610.950 825.600 613.050 826.050 ;
        RECT 571.950 824.400 613.050 825.600 ;
        RECT 571.950 823.950 574.050 824.400 ;
        RECT 610.950 823.950 613.050 824.400 ;
        RECT 625.950 825.600 628.050 826.050 ;
        RECT 694.950 825.600 697.050 826.050 ;
        RECT 625.950 824.400 697.050 825.600 ;
        RECT 625.950 823.950 628.050 824.400 ;
        RECT 694.950 823.950 697.050 824.400 ;
        RECT 853.950 825.600 856.050 826.050 ;
        RECT 895.950 825.600 898.050 826.050 ;
        RECT 853.950 824.400 898.050 825.600 ;
        RECT 853.950 823.950 856.050 824.400 ;
        RECT 895.950 823.950 898.050 824.400 ;
        RECT 127.950 822.600 130.050 823.050 ;
        RECT 190.950 822.600 193.050 823.050 ;
        RECT 127.950 821.400 193.050 822.600 ;
        RECT 127.950 820.950 130.050 821.400 ;
        RECT 190.950 820.950 193.050 821.400 ;
        RECT 286.950 822.600 289.050 823.050 ;
        RECT 295.950 822.600 298.050 823.050 ;
        RECT 397.950 822.600 400.050 823.050 ;
        RECT 286.950 821.400 400.050 822.600 ;
        RECT 446.400 822.600 447.600 823.950 ;
        RECT 493.950 822.600 496.050 823.050 ;
        RECT 446.400 821.400 496.050 822.600 ;
        RECT 286.950 820.950 289.050 821.400 ;
        RECT 295.950 820.950 298.050 821.400 ;
        RECT 397.950 820.950 400.050 821.400 ;
        RECT 493.950 820.950 496.050 821.400 ;
        RECT 514.950 822.600 517.050 823.050 ;
        RECT 538.950 822.600 541.050 823.050 ;
        RECT 562.950 822.600 565.050 823.050 ;
        RECT 697.950 822.600 700.050 823.050 ;
        RECT 514.950 821.400 700.050 822.600 ;
        RECT 514.950 820.950 517.050 821.400 ;
        RECT 538.950 820.950 541.050 821.400 ;
        RECT 562.950 820.950 565.050 821.400 ;
        RECT 697.950 820.950 700.050 821.400 ;
        RECT 811.950 822.600 814.050 823.050 ;
        RECT 868.950 822.600 871.050 823.050 ;
        RECT 811.950 821.400 871.050 822.600 ;
        RECT 811.950 820.950 814.050 821.400 ;
        RECT 868.950 820.950 871.050 821.400 ;
        RECT 34.950 819.600 37.050 820.050 ;
        RECT 55.950 819.600 58.050 820.050 ;
        RECT 34.950 818.400 58.050 819.600 ;
        RECT 34.950 817.950 37.050 818.400 ;
        RECT 55.950 817.950 58.050 818.400 ;
        RECT 364.950 819.600 367.050 820.050 ;
        RECT 373.950 819.600 376.050 820.050 ;
        RECT 364.950 818.400 376.050 819.600 ;
        RECT 364.950 817.950 367.050 818.400 ;
        RECT 373.950 817.950 376.050 818.400 ;
        RECT 388.950 819.600 391.050 820.050 ;
        RECT 400.950 819.600 403.050 820.050 ;
        RECT 388.950 818.400 403.050 819.600 ;
        RECT 388.950 817.950 391.050 818.400 ;
        RECT 400.950 817.950 403.050 818.400 ;
        RECT 430.950 819.600 433.050 820.050 ;
        RECT 535.950 819.600 538.050 820.050 ;
        RECT 430.950 818.400 538.050 819.600 ;
        RECT 430.950 817.950 433.050 818.400 ;
        RECT 535.950 817.950 538.050 818.400 ;
        RECT 544.950 819.600 547.050 820.050 ;
        RECT 580.950 819.600 583.050 820.050 ;
        RECT 544.950 818.400 583.050 819.600 ;
        RECT 544.950 817.950 547.050 818.400 ;
        RECT 580.950 817.950 583.050 818.400 ;
        RECT 703.950 819.600 706.050 820.050 ;
        RECT 712.950 819.600 715.050 820.050 ;
        RECT 703.950 818.400 715.050 819.600 ;
        RECT 703.950 817.950 706.050 818.400 ;
        RECT 712.950 817.950 715.050 818.400 ;
        RECT 748.950 819.600 751.050 820.050 ;
        RECT 796.950 819.600 799.050 820.050 ;
        RECT 748.950 818.400 799.050 819.600 ;
        RECT 748.950 817.950 751.050 818.400 ;
        RECT 796.950 817.950 799.050 818.400 ;
        RECT 343.950 816.600 346.050 817.050 ;
        RECT 376.950 816.600 379.050 817.050 ;
        RECT 343.950 815.400 379.050 816.600 ;
        RECT 343.950 814.950 346.050 815.400 ;
        RECT 376.950 814.950 379.050 815.400 ;
        RECT 553.950 816.600 556.050 817.050 ;
        RECT 604.950 816.600 607.050 817.050 ;
        RECT 553.950 815.400 607.050 816.600 ;
        RECT 553.950 814.950 556.050 815.400 ;
        RECT 604.950 814.950 607.050 815.400 ;
        RECT 706.950 816.600 709.050 817.050 ;
        RECT 718.950 816.600 721.050 817.050 ;
        RECT 817.950 816.600 820.050 817.050 ;
        RECT 706.950 815.400 820.050 816.600 ;
        RECT 706.950 814.950 709.050 815.400 ;
        RECT 718.950 814.950 721.050 815.400 ;
        RECT 817.950 814.950 820.050 815.400 ;
        RECT 85.950 813.600 88.050 814.050 ;
        RECT 109.950 813.600 112.050 814.050 ;
        RECT 127.950 813.600 130.050 814.050 ;
        RECT 85.950 812.400 130.050 813.600 ;
        RECT 85.950 811.950 88.050 812.400 ;
        RECT 109.950 811.950 112.050 812.400 ;
        RECT 127.950 811.950 130.050 812.400 ;
        RECT 232.950 813.600 235.050 814.050 ;
        RECT 415.950 813.600 418.050 814.050 ;
        RECT 232.950 812.400 418.050 813.600 ;
        RECT 232.950 811.950 235.050 812.400 ;
        RECT 415.950 811.950 418.050 812.400 ;
        RECT 478.950 813.600 481.050 814.050 ;
        RECT 526.950 813.600 529.050 814.050 ;
        RECT 478.950 812.400 529.050 813.600 ;
        RECT 478.950 811.950 481.050 812.400 ;
        RECT 526.950 811.950 529.050 812.400 ;
        RECT 538.950 813.600 541.050 814.050 ;
        RECT 652.950 813.600 655.050 814.050 ;
        RECT 538.950 812.400 655.050 813.600 ;
        RECT 538.950 811.950 541.050 812.400 ;
        RECT 652.950 811.950 655.050 812.400 ;
        RECT 703.950 813.600 706.050 814.050 ;
        RECT 745.950 813.600 748.050 814.050 ;
        RECT 766.950 813.600 769.050 814.050 ;
        RECT 703.950 812.400 769.050 813.600 ;
        RECT 703.950 811.950 706.050 812.400 ;
        RECT 745.950 811.950 748.050 812.400 ;
        RECT 766.950 811.950 769.050 812.400 ;
        RECT 850.950 813.600 853.050 814.050 ;
        RECT 889.950 813.600 892.050 814.050 ;
        RECT 850.950 812.400 892.050 813.600 ;
        RECT 850.950 811.950 853.050 812.400 ;
        RECT 889.950 811.950 892.050 812.400 ;
        RECT 157.950 810.600 160.050 811.050 ;
        RECT 184.950 810.600 187.050 811.050 ;
        RECT 157.950 809.400 187.050 810.600 ;
        RECT 157.950 808.950 160.050 809.400 ;
        RECT 184.950 808.950 187.050 809.400 ;
        RECT 304.950 810.600 307.050 811.050 ;
        RECT 328.950 810.600 331.050 811.050 ;
        RECT 304.950 809.400 331.050 810.600 ;
        RECT 304.950 808.950 307.050 809.400 ;
        RECT 328.950 808.950 331.050 809.400 ;
        RECT 454.950 810.600 457.050 811.050 ;
        RECT 469.950 810.600 472.050 811.050 ;
        RECT 539.400 810.600 540.600 811.950 ;
        RECT 454.950 809.400 540.600 810.600 ;
        RECT 622.950 810.600 625.050 811.050 ;
        RECT 631.950 810.600 634.050 811.050 ;
        RECT 622.950 809.400 634.050 810.600 ;
        RECT 454.950 808.950 457.050 809.400 ;
        RECT 469.950 808.950 472.050 809.400 ;
        RECT 622.950 808.950 625.050 809.400 ;
        RECT 631.950 808.950 634.050 809.400 ;
        RECT 811.950 810.600 814.050 811.050 ;
        RECT 820.950 810.600 823.050 811.050 ;
        RECT 811.950 809.400 823.050 810.600 ;
        RECT 811.950 808.950 814.050 809.400 ;
        RECT 820.950 808.950 823.050 809.400 ;
        RECT 4.950 807.750 7.050 808.200 ;
        RECT 31.950 807.750 34.050 808.200 ;
        RECT 4.950 807.600 34.050 807.750 ;
        RECT 37.950 807.600 40.050 808.050 ;
        RECT 4.950 806.550 40.050 807.600 ;
        RECT 4.950 806.100 7.050 806.550 ;
        RECT 31.950 806.400 40.050 806.550 ;
        RECT 31.950 806.100 34.050 806.400 ;
        RECT 37.950 805.950 40.050 806.400 ;
        RECT 61.950 807.750 64.050 808.200 ;
        RECT 85.950 807.750 88.050 808.200 ;
        RECT 61.950 806.550 88.050 807.750 ;
        RECT 61.950 806.100 64.050 806.550 ;
        RECT 85.950 806.100 88.050 806.550 ;
        RECT 94.950 807.600 97.050 808.500 ;
        RECT 103.950 807.750 106.050 808.200 ;
        RECT 109.950 807.750 112.050 808.200 ;
        RECT 103.950 807.600 112.050 807.750 ;
        RECT 94.950 806.550 112.050 807.600 ;
        RECT 94.950 806.400 106.050 806.550 ;
        RECT 103.950 806.100 106.050 806.400 ;
        RECT 109.950 806.100 112.050 806.550 ;
        RECT 127.950 806.100 130.050 808.200 ;
        RECT 133.950 807.750 136.050 808.200 ;
        RECT 142.950 807.750 145.050 808.200 ;
        RECT 133.950 806.550 145.050 807.750 ;
        RECT 133.950 806.100 136.050 806.550 ;
        RECT 142.950 806.100 145.050 806.550 ;
        RECT 166.950 807.600 169.050 808.050 ;
        RECT 175.950 807.600 178.050 808.200 ;
        RECT 166.950 806.400 178.050 807.600 ;
        RECT 128.400 804.600 129.600 806.100 ;
        RECT 166.950 805.950 169.050 806.400 ;
        RECT 175.950 806.100 178.050 806.400 ;
        RECT 196.950 806.100 199.050 808.200 ;
        RECT 208.950 807.600 211.050 808.050 ;
        RECT 214.950 807.600 217.050 808.200 ;
        RECT 208.950 806.400 217.050 807.600 ;
        RECT 128.400 803.400 162.600 804.600 ;
        RECT 34.950 801.450 37.050 801.900 ;
        RECT 40.950 801.450 43.050 802.050 ;
        RECT 34.950 800.250 43.050 801.450 ;
        RECT 34.950 799.800 37.050 800.250 ;
        RECT 40.950 799.950 43.050 800.250 ;
        RECT 112.950 801.600 115.050 801.900 ;
        RECT 130.950 801.600 133.050 801.900 ;
        RECT 112.950 800.400 133.050 801.600 ;
        RECT 112.950 799.800 115.050 800.400 ;
        RECT 130.950 799.800 133.050 800.400 ;
        RECT 148.950 801.600 151.050 802.050 ;
        RECT 154.950 801.600 157.050 801.900 ;
        RECT 148.950 800.400 157.050 801.600 ;
        RECT 161.400 801.600 162.600 803.400 ;
        RECT 178.950 801.600 181.050 801.900 ;
        RECT 161.400 800.400 181.050 801.600 ;
        RECT 197.400 801.600 198.600 806.100 ;
        RECT 208.950 805.950 211.050 806.400 ;
        RECT 214.950 806.100 217.050 806.400 ;
        RECT 220.950 806.100 223.050 808.200 ;
        RECT 241.950 807.600 244.050 808.200 ;
        RECT 253.950 807.750 256.050 808.200 ;
        RECT 268.950 807.750 271.050 808.200 ;
        RECT 253.950 807.600 271.050 807.750 ;
        RECT 304.950 807.600 307.050 808.200 ;
        RECT 241.950 806.550 271.050 807.600 ;
        RECT 241.950 806.400 256.050 806.550 ;
        RECT 241.950 806.100 244.050 806.400 ;
        RECT 253.950 806.100 256.050 806.400 ;
        RECT 268.950 806.100 271.050 806.550 ;
        RECT 290.400 806.400 307.050 807.600 ;
        RECT 221.400 801.600 222.600 806.100 ;
        RECT 290.400 801.900 291.600 806.400 ;
        RECT 304.950 806.100 307.050 806.400 ;
        RECT 310.950 807.600 313.050 808.200 ;
        RECT 322.950 807.600 325.050 808.050 ;
        RECT 310.950 806.400 325.050 807.600 ;
        RECT 310.950 806.100 313.050 806.400 ;
        RECT 322.950 805.950 325.050 806.400 ;
        RECT 334.950 807.750 337.050 808.200 ;
        RECT 343.950 807.750 346.050 808.200 ;
        RECT 334.950 806.550 346.050 807.750 ;
        RECT 334.950 806.100 337.050 806.550 ;
        RECT 343.950 806.100 346.050 806.550 ;
        RECT 355.950 807.600 358.050 808.200 ;
        RECT 385.950 807.750 388.050 808.200 ;
        RECT 403.950 807.750 406.050 808.200 ;
        RECT 385.950 807.600 406.050 807.750 ;
        RECT 355.950 806.550 406.050 807.600 ;
        RECT 355.950 806.400 388.050 806.550 ;
        RECT 355.950 806.100 358.050 806.400 ;
        RECT 385.950 806.100 388.050 806.400 ;
        RECT 403.950 806.100 406.050 806.550 ;
        RECT 415.950 807.600 420.000 808.050 ;
        RECT 433.950 807.750 436.050 808.200 ;
        RECT 445.950 807.750 448.050 808.200 ;
        RECT 415.950 805.950 420.600 807.600 ;
        RECT 433.950 806.550 448.050 807.750 ;
        RECT 433.950 806.100 436.050 806.550 ;
        RECT 445.950 806.100 448.050 806.550 ;
        RECT 490.950 806.100 493.050 808.200 ;
        RECT 526.950 807.600 529.050 808.050 ;
        RECT 553.950 807.600 556.050 808.200 ;
        RECT 526.950 806.400 556.050 807.600 ;
        RECT 262.950 801.600 265.050 801.900 ;
        RECT 197.400 800.400 265.050 801.600 ;
        RECT 148.950 799.950 151.050 800.400 ;
        RECT 154.950 799.800 157.050 800.400 ;
        RECT 178.950 799.800 181.050 800.400 ;
        RECT 262.950 799.800 265.050 800.400 ;
        RECT 289.950 799.800 292.050 801.900 ;
        RECT 295.950 801.450 298.050 801.900 ;
        RECT 301.950 801.450 304.050 801.900 ;
        RECT 295.950 800.250 304.050 801.450 ;
        RECT 295.950 799.800 298.050 800.250 ;
        RECT 301.950 799.800 304.050 800.250 ;
        RECT 343.950 801.600 346.050 802.050 ;
        RECT 352.950 801.600 355.050 801.900 ;
        RECT 343.950 800.400 355.050 801.600 ;
        RECT 343.950 799.950 346.050 800.400 ;
        RECT 352.950 799.800 355.050 800.400 ;
        RECT 388.950 801.600 391.050 802.050 ;
        RECT 419.400 801.900 420.600 805.950 ;
        RECT 400.950 801.600 403.050 801.900 ;
        RECT 388.950 800.400 403.050 801.600 ;
        RECT 388.950 799.950 391.050 800.400 ;
        RECT 400.950 799.800 403.050 800.400 ;
        RECT 418.950 799.800 421.050 801.900 ;
        RECT 448.950 801.450 451.050 801.900 ;
        RECT 454.950 801.450 457.050 801.900 ;
        RECT 448.950 800.250 457.050 801.450 ;
        RECT 448.950 799.800 451.050 800.250 ;
        RECT 454.950 799.800 457.050 800.250 ;
        RECT 472.950 801.450 475.050 801.900 ;
        RECT 478.950 801.450 481.050 801.900 ;
        RECT 472.950 800.250 481.050 801.450 ;
        RECT 491.400 801.600 492.600 806.100 ;
        RECT 526.950 805.950 529.050 806.400 ;
        RECT 553.950 806.100 556.050 806.400 ;
        RECT 586.950 807.600 589.050 808.200 ;
        RECT 598.950 807.750 601.050 808.200 ;
        RECT 613.950 807.750 616.050 808.200 ;
        RECT 598.950 807.600 616.050 807.750 ;
        RECT 586.950 806.550 616.050 807.600 ;
        RECT 586.950 806.400 601.050 806.550 ;
        RECT 586.950 806.100 589.050 806.400 ;
        RECT 598.950 806.100 601.050 806.400 ;
        RECT 613.950 806.100 616.050 806.550 ;
        RECT 634.950 807.750 637.050 808.200 ;
        RECT 643.950 807.750 646.050 808.200 ;
        RECT 634.950 806.550 646.050 807.750 ;
        RECT 634.950 806.100 637.050 806.550 ;
        RECT 643.950 806.100 646.050 806.550 ;
        RECT 652.950 806.100 655.050 808.200 ;
        RECT 658.950 807.600 661.050 808.200 ;
        RECT 667.950 807.600 670.050 808.050 ;
        RECT 676.950 807.600 679.050 808.200 ;
        RECT 658.950 806.400 679.050 807.600 ;
        RECT 658.950 806.100 661.050 806.400 ;
        RECT 653.400 804.600 654.600 806.100 ;
        RECT 667.950 805.950 670.050 806.400 ;
        RECT 676.950 806.100 679.050 806.400 ;
        RECT 682.950 807.600 685.050 808.200 ;
        RECT 688.950 807.600 691.050 808.050 ;
        RECT 682.950 806.400 691.050 807.600 ;
        RECT 682.950 806.100 685.050 806.400 ;
        RECT 688.950 805.950 691.050 806.400 ;
        RECT 733.950 807.600 736.050 808.200 ;
        RECT 781.950 807.600 784.050 808.200 ;
        RECT 733.950 806.400 784.050 807.600 ;
        RECT 733.950 806.100 736.050 806.400 ;
        RECT 781.950 806.100 784.050 806.400 ;
        RECT 790.950 807.750 793.050 808.200 ;
        RECT 802.950 807.750 805.050 808.200 ;
        RECT 790.950 806.550 805.050 807.750 ;
        RECT 826.950 807.600 829.050 808.200 ;
        RECT 790.950 806.100 793.050 806.550 ;
        RECT 802.950 806.100 805.050 806.550 ;
        RECT 806.400 806.400 829.050 807.600 ;
        RECT 782.400 804.600 783.600 806.100 ;
        RECT 806.400 804.600 807.600 806.400 ;
        RECT 826.950 806.100 829.050 806.400 ;
        RECT 850.950 807.600 853.050 808.200 ;
        RECT 874.950 807.750 877.050 808.200 ;
        RECT 883.950 807.750 886.050 808.200 ;
        RECT 874.950 807.600 886.050 807.750 ;
        RECT 850.950 806.550 886.050 807.600 ;
        RECT 850.950 806.400 877.050 806.550 ;
        RECT 850.950 806.100 853.050 806.400 ;
        RECT 874.950 806.100 877.050 806.400 ;
        RECT 883.950 806.100 886.050 806.550 ;
        RECT 653.400 803.400 705.600 804.600 ;
        RECT 782.400 803.400 807.600 804.600 ;
        RECT 517.950 801.600 520.050 801.900 ;
        RECT 491.400 800.400 520.050 801.600 ;
        RECT 472.950 799.800 475.050 800.250 ;
        RECT 478.950 799.800 481.050 800.250 ;
        RECT 517.950 799.800 520.050 800.400 ;
        RECT 535.950 801.600 538.050 801.900 ;
        RECT 556.950 801.600 559.050 801.900 ;
        RECT 535.950 800.400 559.050 801.600 ;
        RECT 535.950 799.800 538.050 800.400 ;
        RECT 556.950 799.800 559.050 800.400 ;
        RECT 583.950 801.600 586.050 801.900 ;
        RECT 601.950 801.600 604.050 801.900 ;
        RECT 583.950 800.400 604.050 801.600 ;
        RECT 583.950 799.800 586.050 800.400 ;
        RECT 601.950 799.800 604.050 800.400 ;
        RECT 607.950 801.600 610.050 801.900 ;
        RECT 631.950 801.600 634.050 801.900 ;
        RECT 607.950 800.400 634.050 801.600 ;
        RECT 607.950 799.800 610.050 800.400 ;
        RECT 631.950 799.800 634.050 800.400 ;
        RECT 643.950 801.600 646.050 802.050 ;
        RECT 655.950 801.600 658.050 801.900 ;
        RECT 643.950 800.400 658.050 801.600 ;
        RECT 643.950 799.950 646.050 800.400 ;
        RECT 655.950 799.800 658.050 800.400 ;
        RECT 688.950 801.450 691.050 801.900 ;
        RECT 700.950 801.450 703.050 801.900 ;
        RECT 688.950 800.250 703.050 801.450 ;
        RECT 704.400 801.600 705.600 803.400 ;
        RECT 706.950 801.600 709.050 801.900 ;
        RECT 704.400 800.400 709.050 801.600 ;
        RECT 688.950 799.800 691.050 800.250 ;
        RECT 700.950 799.800 703.050 800.250 ;
        RECT 706.950 799.800 709.050 800.400 ;
        RECT 745.950 801.450 748.050 801.900 ;
        RECT 760.950 801.450 763.050 801.900 ;
        RECT 745.950 800.250 763.050 801.450 ;
        RECT 745.950 799.800 748.050 800.250 ;
        RECT 760.950 799.800 763.050 800.250 ;
        RECT 799.950 801.600 802.050 801.900 ;
        RECT 823.950 801.600 826.050 801.900 ;
        RECT 799.950 800.400 826.050 801.600 ;
        RECT 799.950 799.800 802.050 800.400 ;
        RECT 823.950 799.800 826.050 800.400 ;
        RECT 853.950 801.600 856.050 801.900 ;
        RECT 871.950 801.600 874.050 801.900 ;
        RECT 853.950 800.400 874.050 801.600 ;
        RECT 853.950 799.800 856.050 800.400 ;
        RECT 871.950 799.800 874.050 800.400 ;
        RECT 10.950 798.600 13.050 799.050 ;
        RECT 25.950 798.600 28.050 799.050 ;
        RECT 46.950 798.600 49.050 799.050 ;
        RECT 58.950 798.600 61.050 799.050 ;
        RECT 10.950 797.400 61.050 798.600 ;
        RECT 10.950 796.950 13.050 797.400 ;
        RECT 25.950 796.950 28.050 797.400 ;
        RECT 46.950 796.950 49.050 797.400 ;
        RECT 58.950 796.950 61.050 797.400 ;
        RECT 67.950 798.600 70.050 799.050 ;
        RECT 82.950 798.600 85.050 799.050 ;
        RECT 67.950 797.400 85.050 798.600 ;
        RECT 67.950 796.950 70.050 797.400 ;
        RECT 82.950 796.950 85.050 797.400 ;
        RECT 661.950 798.600 664.050 799.050 ;
        RECT 679.950 798.600 682.050 799.050 ;
        RECT 661.950 797.400 682.050 798.600 ;
        RECT 661.950 796.950 664.050 797.400 ;
        RECT 679.950 796.950 682.050 797.400 ;
        RECT 790.950 798.600 793.050 799.050 ;
        RECT 808.950 798.600 811.050 799.050 ;
        RECT 790.950 797.400 811.050 798.600 ;
        RECT 790.950 796.950 793.050 797.400 ;
        RECT 808.950 796.950 811.050 797.400 ;
        RECT 847.950 798.600 850.050 799.050 ;
        RECT 877.950 798.600 880.050 799.050 ;
        RECT 847.950 797.400 880.050 798.600 ;
        RECT 847.950 796.950 850.050 797.400 ;
        RECT 877.950 796.950 880.050 797.400 ;
        RECT 127.950 795.600 130.050 796.050 ;
        RECT 136.950 795.600 139.050 796.050 ;
        RECT 127.950 794.400 139.050 795.600 ;
        RECT 127.950 793.950 130.050 794.400 ;
        RECT 136.950 793.950 139.050 794.400 ;
        RECT 193.950 795.600 196.050 796.050 ;
        RECT 247.950 795.600 250.050 796.050 ;
        RECT 193.950 794.400 250.050 795.600 ;
        RECT 193.950 793.950 196.050 794.400 ;
        RECT 247.950 793.950 250.050 794.400 ;
        RECT 262.950 795.600 265.050 796.050 ;
        RECT 313.950 795.600 316.050 796.050 ;
        RECT 262.950 794.400 316.050 795.600 ;
        RECT 262.950 793.950 265.050 794.400 ;
        RECT 313.950 793.950 316.050 794.400 ;
        RECT 331.950 795.600 334.050 796.050 ;
        RECT 373.950 795.600 376.050 796.050 ;
        RECT 331.950 794.400 376.050 795.600 ;
        RECT 331.950 793.950 334.050 794.400 ;
        RECT 373.950 793.950 376.050 794.400 ;
        RECT 442.950 795.600 445.050 796.050 ;
        RECT 478.950 795.600 481.050 796.050 ;
        RECT 442.950 794.400 481.050 795.600 ;
        RECT 442.950 793.950 445.050 794.400 ;
        RECT 478.950 793.950 481.050 794.400 ;
        RECT 637.950 795.600 640.050 796.050 ;
        RECT 667.950 795.600 670.050 796.050 ;
        RECT 694.950 795.600 697.050 796.050 ;
        RECT 637.950 794.400 697.050 795.600 ;
        RECT 637.950 793.950 640.050 794.400 ;
        RECT 667.950 793.950 670.050 794.400 ;
        RECT 694.950 793.950 697.050 794.400 ;
        RECT 724.950 795.600 727.050 796.050 ;
        RECT 751.950 795.600 754.050 796.050 ;
        RECT 724.950 794.400 754.050 795.600 ;
        RECT 724.950 793.950 727.050 794.400 ;
        RECT 751.950 793.950 754.050 794.400 ;
        RECT 76.950 792.600 79.050 793.050 ;
        RECT 142.950 792.600 145.050 793.050 ;
        RECT 76.950 791.400 145.050 792.600 ;
        RECT 76.950 790.950 79.050 791.400 ;
        RECT 142.950 790.950 145.050 791.400 ;
        RECT 346.950 792.600 349.050 793.050 ;
        RECT 388.950 792.600 391.050 793.050 ;
        RECT 346.950 791.400 391.050 792.600 ;
        RECT 346.950 790.950 349.050 791.400 ;
        RECT 388.950 790.950 391.050 791.400 ;
        RECT 622.950 792.600 625.050 793.050 ;
        RECT 637.950 792.600 640.050 792.900 ;
        RECT 622.950 791.400 640.050 792.600 ;
        RECT 622.950 790.950 625.050 791.400 ;
        RECT 637.950 790.800 640.050 791.400 ;
        RECT 778.950 792.600 781.050 793.050 ;
        RECT 835.950 792.600 838.050 793.050 ;
        RECT 778.950 791.400 838.050 792.600 ;
        RECT 778.950 790.950 781.050 791.400 ;
        RECT 835.950 790.950 838.050 791.400 ;
        RECT 172.950 789.600 175.050 790.050 ;
        RECT 184.950 789.600 187.050 790.050 ;
        RECT 196.950 789.600 199.050 790.050 ;
        RECT 172.950 788.400 199.050 789.600 ;
        RECT 172.950 787.950 175.050 788.400 ;
        RECT 184.950 787.950 187.050 788.400 ;
        RECT 196.950 787.950 199.050 788.400 ;
        RECT 256.950 789.600 259.050 790.050 ;
        RECT 274.950 789.600 277.050 790.050 ;
        RECT 256.950 788.400 277.050 789.600 ;
        RECT 256.950 787.950 259.050 788.400 ;
        RECT 274.950 787.950 277.050 788.400 ;
        RECT 433.950 789.600 436.050 790.050 ;
        RECT 466.950 789.600 469.050 790.050 ;
        RECT 487.950 789.600 490.050 790.050 ;
        RECT 550.950 789.600 553.050 790.050 ;
        RECT 433.950 788.400 553.050 789.600 ;
        RECT 433.950 787.950 436.050 788.400 ;
        RECT 466.950 787.950 469.050 788.400 ;
        RECT 487.950 787.950 490.050 788.400 ;
        RECT 550.950 787.950 553.050 788.400 ;
        RECT 556.950 789.600 559.050 790.050 ;
        RECT 571.950 789.600 574.050 790.050 ;
        RECT 556.950 788.400 574.050 789.600 ;
        RECT 556.950 787.950 559.050 788.400 ;
        RECT 571.950 787.950 574.050 788.400 ;
        RECT 577.950 789.600 580.050 790.050 ;
        RECT 649.950 789.600 652.050 790.050 ;
        RECT 661.950 789.600 664.050 790.050 ;
        RECT 577.950 788.400 664.050 789.600 ;
        RECT 577.950 787.950 580.050 788.400 ;
        RECT 649.950 787.950 652.050 788.400 ;
        RECT 661.950 787.950 664.050 788.400 ;
        RECT 325.950 786.600 328.050 787.050 ;
        RECT 361.950 786.600 364.050 787.050 ;
        RECT 325.950 785.400 364.050 786.600 ;
        RECT 325.950 784.950 328.050 785.400 ;
        RECT 361.950 784.950 364.050 785.400 ;
        RECT 496.950 786.600 499.050 787.050 ;
        RECT 511.950 786.600 514.050 787.050 ;
        RECT 559.950 786.600 562.050 787.050 ;
        RECT 496.950 785.400 562.050 786.600 ;
        RECT 496.950 784.950 499.050 785.400 ;
        RECT 511.950 784.950 514.050 785.400 ;
        RECT 559.950 784.950 562.050 785.400 ;
        RECT 565.950 786.600 568.050 787.050 ;
        RECT 724.950 786.600 727.050 787.050 ;
        RECT 565.950 785.400 727.050 786.600 ;
        RECT 565.950 784.950 568.050 785.400 ;
        RECT 724.950 784.950 727.050 785.400 ;
        RECT 730.950 786.600 733.050 787.050 ;
        RECT 778.950 786.600 781.050 787.050 ;
        RECT 730.950 785.400 781.050 786.600 ;
        RECT 730.950 784.950 733.050 785.400 ;
        RECT 778.950 784.950 781.050 785.400 ;
        RECT 805.950 786.600 808.050 787.050 ;
        RECT 811.950 786.600 814.050 787.050 ;
        RECT 874.950 786.600 877.050 787.050 ;
        RECT 805.950 785.400 877.050 786.600 ;
        RECT 805.950 784.950 808.050 785.400 ;
        RECT 811.950 784.950 814.050 785.400 ;
        RECT 874.950 784.950 877.050 785.400 ;
        RECT 526.950 783.600 529.050 784.050 ;
        RECT 556.950 783.600 559.050 784.050 ;
        RECT 526.950 782.400 559.050 783.600 ;
        RECT 526.950 781.950 529.050 782.400 ;
        RECT 556.950 781.950 559.050 782.400 ;
        RECT 601.950 783.600 604.050 784.050 ;
        RECT 667.950 783.600 670.050 784.050 ;
        RECT 601.950 782.400 670.050 783.600 ;
        RECT 601.950 781.950 604.050 782.400 ;
        RECT 667.950 781.950 670.050 782.400 ;
        RECT 877.950 783.600 880.050 784.050 ;
        RECT 883.950 783.600 886.050 784.050 ;
        RECT 877.950 782.400 886.050 783.600 ;
        RECT 877.950 781.950 880.050 782.400 ;
        RECT 883.950 781.950 886.050 782.400 ;
        RECT 16.950 780.600 19.050 781.050 ;
        RECT 43.950 780.600 46.050 781.050 ;
        RECT 52.950 780.600 55.050 781.050 ;
        RECT 118.950 780.600 121.050 781.050 ;
        RECT 16.950 779.400 121.050 780.600 ;
        RECT 16.950 778.950 19.050 779.400 ;
        RECT 43.950 778.950 46.050 779.400 ;
        RECT 52.950 778.950 55.050 779.400 ;
        RECT 118.950 778.950 121.050 779.400 ;
        RECT 337.950 780.600 340.050 781.050 ;
        RECT 403.950 780.600 406.050 781.050 ;
        RECT 409.950 780.600 412.050 781.050 ;
        RECT 337.950 779.400 412.050 780.600 ;
        RECT 337.950 778.950 340.050 779.400 ;
        RECT 403.950 778.950 406.050 779.400 ;
        RECT 409.950 778.950 412.050 779.400 ;
        RECT 424.950 780.600 427.050 781.050 ;
        RECT 571.950 780.600 574.050 781.050 ;
        RECT 424.950 779.400 574.050 780.600 ;
        RECT 424.950 778.950 427.050 779.400 ;
        RECT 571.950 778.950 574.050 779.400 ;
        RECT 613.950 780.600 616.050 781.050 ;
        RECT 613.950 779.400 651.600 780.600 ;
        RECT 613.950 778.950 616.050 779.400 ;
        RECT 373.950 777.600 376.050 778.050 ;
        RECT 382.950 777.600 385.050 778.050 ;
        RECT 373.950 776.400 385.050 777.600 ;
        RECT 373.950 775.950 376.050 776.400 ;
        RECT 382.950 775.950 385.050 776.400 ;
        RECT 400.950 777.600 403.050 778.050 ;
        RECT 460.950 777.600 463.050 778.050 ;
        RECT 400.950 776.400 463.050 777.600 ;
        RECT 400.950 775.950 403.050 776.400 ;
        RECT 460.950 775.950 463.050 776.400 ;
        RECT 472.950 777.600 475.050 778.050 ;
        RECT 550.950 777.600 553.050 778.050 ;
        RECT 472.950 776.400 553.050 777.600 ;
        RECT 650.400 777.600 651.600 779.400 ;
        RECT 718.950 777.600 721.050 778.050 ;
        RECT 650.400 776.400 721.050 777.600 ;
        RECT 472.950 775.950 475.050 776.400 ;
        RECT 550.950 775.950 553.050 776.400 ;
        RECT 718.950 775.950 721.050 776.400 ;
        RECT 307.950 774.600 310.050 775.050 ;
        RECT 316.950 774.600 319.050 775.050 ;
        RECT 307.950 773.400 319.050 774.600 ;
        RECT 307.950 772.950 310.050 773.400 ;
        RECT 316.950 772.950 319.050 773.400 ;
        RECT 589.950 774.600 592.050 775.050 ;
        RECT 712.950 774.600 715.050 775.050 ;
        RECT 589.950 773.400 715.050 774.600 ;
        RECT 589.950 772.950 592.050 773.400 ;
        RECT 712.950 772.950 715.050 773.400 ;
        RECT 763.950 774.600 766.050 775.050 ;
        RECT 805.950 774.600 808.050 775.050 ;
        RECT 847.950 774.600 850.050 775.050 ;
        RECT 763.950 773.400 850.050 774.600 ;
        RECT 763.950 772.950 766.050 773.400 ;
        RECT 805.950 772.950 808.050 773.400 ;
        RECT 847.950 772.950 850.050 773.400 ;
        RECT 166.950 771.600 169.050 772.050 ;
        RECT 184.950 771.600 187.050 772.050 ;
        RECT 166.950 770.400 187.050 771.600 ;
        RECT 166.950 769.950 169.050 770.400 ;
        RECT 184.950 769.950 187.050 770.400 ;
        RECT 358.950 771.600 361.050 772.050 ;
        RECT 373.950 771.600 376.050 772.050 ;
        RECT 358.950 770.400 376.050 771.600 ;
        RECT 358.950 769.950 361.050 770.400 ;
        RECT 373.950 769.950 376.050 770.400 ;
        RECT 385.950 771.600 388.050 772.050 ;
        RECT 424.950 771.600 427.050 772.050 ;
        RECT 385.950 770.400 427.050 771.600 ;
        RECT 385.950 769.950 388.050 770.400 ;
        RECT 424.950 769.950 427.050 770.400 ;
        RECT 556.950 771.600 559.050 772.050 ;
        RECT 577.950 771.600 580.050 772.050 ;
        RECT 556.950 770.400 580.050 771.600 ;
        RECT 556.950 769.950 559.050 770.400 ;
        RECT 577.950 769.950 580.050 770.400 ;
        RECT 607.950 771.600 610.050 772.050 ;
        RECT 676.950 771.600 679.050 772.050 ;
        RECT 607.950 770.400 679.050 771.600 ;
        RECT 607.950 769.950 610.050 770.400 ;
        RECT 676.950 769.950 679.050 770.400 ;
        RECT 715.950 771.600 718.050 772.050 ;
        RECT 748.950 771.600 751.050 772.050 ;
        RECT 715.950 770.400 751.050 771.600 ;
        RECT 715.950 769.950 718.050 770.400 ;
        RECT 748.950 769.950 751.050 770.400 ;
        RECT 1.950 768.600 4.050 769.050 ;
        RECT 34.950 768.600 37.050 769.050 ;
        RECT 1.950 767.400 37.050 768.600 ;
        RECT 1.950 766.950 4.050 767.400 ;
        RECT 34.950 766.950 37.050 767.400 ;
        RECT 82.950 768.600 85.050 769.050 ;
        RECT 109.950 768.600 112.050 769.050 ;
        RECT 82.950 767.400 112.050 768.600 ;
        RECT 82.950 766.950 85.050 767.400 ;
        RECT 109.950 766.950 112.050 767.400 ;
        RECT 151.950 768.600 154.050 769.050 ;
        RECT 163.950 768.600 166.050 769.050 ;
        RECT 151.950 767.400 166.050 768.600 ;
        RECT 151.950 766.950 154.050 767.400 ;
        RECT 163.950 766.950 166.050 767.400 ;
        RECT 193.950 768.600 196.050 769.050 ;
        RECT 214.950 768.600 217.050 769.050 ;
        RECT 193.950 767.400 217.050 768.600 ;
        RECT 193.950 766.950 196.050 767.400 ;
        RECT 214.950 766.950 217.050 767.400 ;
        RECT 238.950 768.600 241.050 769.050 ;
        RECT 268.950 768.600 271.050 769.050 ;
        RECT 469.950 768.600 472.050 769.050 ;
        RECT 238.950 767.400 472.050 768.600 ;
        RECT 238.950 766.950 241.050 767.400 ;
        RECT 268.950 766.950 271.050 767.400 ;
        RECT 469.950 766.950 472.050 767.400 ;
        RECT 553.950 768.600 556.050 769.050 ;
        RECT 562.950 768.600 565.050 769.050 ;
        RECT 553.950 767.400 565.050 768.600 ;
        RECT 553.950 766.950 556.050 767.400 ;
        RECT 562.950 766.950 565.050 767.400 ;
        RECT 682.950 768.600 685.050 769.050 ;
        RECT 706.950 768.600 709.050 769.050 ;
        RECT 682.950 767.400 709.050 768.600 ;
        RECT 682.950 766.950 685.050 767.400 ;
        RECT 706.950 766.950 709.050 767.400 ;
        RECT 79.950 765.600 82.050 766.050 ;
        RECT 85.950 765.600 88.050 766.050 ;
        RECT 79.950 764.400 88.050 765.600 ;
        RECT 79.950 763.950 82.050 764.400 ;
        RECT 85.950 763.950 88.050 764.400 ;
        RECT 319.950 765.600 322.050 766.050 ;
        RECT 367.950 765.600 370.050 766.050 ;
        RECT 319.950 764.400 370.050 765.600 ;
        RECT 319.950 763.950 322.050 764.400 ;
        RECT 367.950 763.950 370.050 764.400 ;
        RECT 481.950 765.600 484.050 766.050 ;
        RECT 595.950 765.600 598.050 766.050 ;
        RECT 610.950 765.600 613.050 766.050 ;
        RECT 481.950 764.400 567.600 765.600 ;
        RECT 481.950 763.950 484.050 764.400 ;
        RECT 566.400 763.200 567.600 764.400 ;
        RECT 595.950 764.400 613.050 765.600 ;
        RECT 595.950 763.950 598.050 764.400 ;
        RECT 610.950 763.950 613.050 764.400 ;
        RECT 712.950 765.600 715.050 766.050 ;
        RECT 730.950 765.600 733.050 766.050 ;
        RECT 712.950 764.400 733.050 765.600 ;
        RECT 712.950 763.950 715.050 764.400 ;
        RECT 730.950 763.950 733.050 764.400 ;
        RECT 7.950 762.600 10.050 763.050 ;
        RECT 13.950 762.600 16.050 763.200 ;
        RECT 28.950 762.600 31.050 763.200 ;
        RECT 7.950 761.400 16.050 762.600 ;
        RECT 7.950 760.950 10.050 761.400 ;
        RECT 13.950 761.100 16.050 761.400 ;
        RECT 17.400 761.400 31.050 762.600 ;
        RECT 17.400 756.900 18.600 761.400 ;
        RECT 28.950 761.100 31.050 761.400 ;
        RECT 34.950 761.100 37.050 763.200 ;
        RECT 43.950 762.750 46.050 763.200 ;
        RECT 58.950 762.750 61.050 763.200 ;
        RECT 43.950 762.600 61.050 762.750 ;
        RECT 73.950 762.600 76.050 763.200 ;
        RECT 43.950 761.550 76.050 762.600 ;
        RECT 43.950 761.100 46.050 761.550 ;
        RECT 58.950 761.400 76.050 761.550 ;
        RECT 58.950 761.100 61.050 761.400 ;
        RECT 73.950 761.100 76.050 761.400 ;
        RECT 88.950 762.600 91.050 763.050 ;
        RECT 97.950 762.600 100.050 763.200 ;
        RECT 118.950 762.600 121.050 763.200 ;
        RECT 88.950 761.400 100.050 762.600 ;
        RECT 35.400 759.600 36.600 761.100 ;
        RECT 88.950 760.950 91.050 761.400 ;
        RECT 97.950 761.100 100.050 761.400 ;
        RECT 101.400 761.400 121.050 762.600 ;
        RECT 64.950 759.600 67.050 760.050 ;
        RECT 101.400 759.600 102.600 761.400 ;
        RECT 118.950 761.100 121.050 761.400 ;
        RECT 139.950 762.600 142.050 763.200 ;
        RECT 148.950 762.600 151.050 763.050 ;
        RECT 139.950 761.400 151.050 762.600 ;
        RECT 139.950 761.100 142.050 761.400 ;
        RECT 148.950 760.950 151.050 761.400 ;
        RECT 160.950 762.750 163.050 763.200 ;
        RECT 166.950 762.750 169.050 763.200 ;
        RECT 160.950 761.550 169.050 762.750 ;
        RECT 160.950 761.100 163.050 761.550 ;
        RECT 166.950 761.100 169.050 761.550 ;
        RECT 178.950 761.100 181.050 763.200 ;
        RECT 199.950 762.600 202.050 763.050 ;
        RECT 208.950 762.600 211.050 763.200 ;
        RECT 199.950 761.400 211.050 762.600 ;
        RECT 35.400 758.400 67.050 759.600 ;
        RECT 64.950 757.950 67.050 758.400 ;
        RECT 95.400 758.400 102.600 759.600 ;
        RECT 16.950 754.800 19.050 756.900 ;
        RECT 31.950 756.600 34.050 756.900 ;
        RECT 43.950 756.600 46.050 757.050 ;
        RECT 95.400 756.900 96.600 758.400 ;
        RECT 31.950 755.400 46.050 756.600 ;
        RECT 31.950 754.800 34.050 755.400 ;
        RECT 43.950 754.950 46.050 755.400 ;
        RECT 94.950 754.800 97.050 756.900 ;
        RECT 106.950 756.600 109.050 757.050 ;
        RECT 115.950 756.600 118.050 756.900 ;
        RECT 106.950 755.400 118.050 756.600 ;
        RECT 106.950 754.950 109.050 755.400 ;
        RECT 115.950 754.800 118.050 755.400 ;
        RECT 130.950 756.600 133.050 757.050 ;
        RECT 136.950 756.600 139.050 756.900 ;
        RECT 130.950 755.400 139.050 756.600 ;
        RECT 130.950 754.950 133.050 755.400 ;
        RECT 136.950 754.800 139.050 755.400 ;
        RECT 142.950 756.600 145.050 756.900 ;
        RECT 166.950 756.600 169.050 757.050 ;
        RECT 175.950 756.600 178.050 756.900 ;
        RECT 142.950 755.400 178.050 756.600 ;
        RECT 142.950 754.800 145.050 755.400 ;
        RECT 166.950 754.950 169.050 755.400 ;
        RECT 175.950 754.800 178.050 755.400 ;
        RECT 179.400 751.050 180.600 761.100 ;
        RECT 199.950 760.950 202.050 761.400 ;
        RECT 208.950 761.100 211.050 761.400 ;
        RECT 232.950 762.750 235.050 763.200 ;
        RECT 244.950 762.750 247.050 763.200 ;
        RECT 232.950 761.550 247.050 762.750 ;
        RECT 259.950 762.600 262.050 763.200 ;
        RECT 232.950 761.100 235.050 761.550 ;
        RECT 244.950 761.100 247.050 761.550 ;
        RECT 257.400 761.400 262.050 762.600 ;
        RECT 247.950 759.600 250.050 760.050 ;
        RECT 257.400 759.600 258.600 761.400 ;
        RECT 259.950 761.100 262.050 761.400 ;
        RECT 265.950 761.100 268.050 763.200 ;
        RECT 271.950 762.750 274.050 763.200 ;
        RECT 283.950 762.750 286.050 763.200 ;
        RECT 271.950 761.550 286.050 762.750 ;
        RECT 271.950 761.100 274.050 761.550 ;
        RECT 283.950 761.100 286.050 761.550 ;
        RECT 295.950 762.750 298.050 763.200 ;
        RECT 307.950 762.750 310.050 763.200 ;
        RECT 295.950 761.550 310.050 762.750 ;
        RECT 295.950 761.100 298.050 761.550 ;
        RECT 307.950 761.100 310.050 761.550 ;
        RECT 247.950 758.400 258.600 759.600 ;
        RECT 247.950 757.950 250.050 758.400 ;
        RECT 266.400 757.050 267.600 761.100 ;
        RECT 313.950 760.950 316.050 763.050 ;
        RECT 343.950 762.600 346.050 763.050 ;
        RECT 349.950 762.600 352.050 763.200 ;
        RECT 343.950 761.400 352.050 762.600 ;
        RECT 343.950 760.950 346.050 761.400 ;
        RECT 349.950 761.100 352.050 761.400 ;
        RECT 364.950 760.950 367.050 763.050 ;
        RECT 424.950 762.750 427.050 763.200 ;
        RECT 436.950 762.750 439.050 763.200 ;
        RECT 424.950 761.550 439.050 762.750 ;
        RECT 424.950 761.100 427.050 761.550 ;
        RECT 436.950 761.100 439.050 761.550 ;
        RECT 442.950 761.100 445.050 763.200 ;
        RECT 487.950 762.750 490.050 763.200 ;
        RECT 496.950 762.750 499.050 763.200 ;
        RECT 487.950 761.550 499.050 762.750 ;
        RECT 487.950 761.100 490.050 761.550 ;
        RECT 496.950 761.100 499.050 761.550 ;
        RECT 523.950 762.600 526.050 763.050 ;
        RECT 532.950 762.600 535.050 763.200 ;
        RECT 523.950 761.400 535.050 762.600 ;
        RECT 196.950 756.600 199.050 757.050 ;
        RECT 205.950 756.600 208.050 756.900 ;
        RECT 196.950 755.400 208.050 756.600 ;
        RECT 196.950 754.950 199.050 755.400 ;
        RECT 205.950 754.800 208.050 755.400 ;
        RECT 235.950 756.600 238.050 756.900 ;
        RECT 256.950 756.600 259.050 756.900 ;
        RECT 235.950 755.400 259.050 756.600 ;
        RECT 266.400 755.400 271.050 757.050 ;
        RECT 235.950 754.800 238.050 755.400 ;
        RECT 256.950 754.800 259.050 755.400 ;
        RECT 267.000 754.950 271.050 755.400 ;
        RECT 274.950 756.600 277.050 757.050 ;
        RECT 280.950 756.600 283.050 756.900 ;
        RECT 274.950 755.400 283.050 756.600 ;
        RECT 274.950 754.950 277.050 755.400 ;
        RECT 280.950 754.800 283.050 755.400 ;
        RECT 286.950 756.600 289.050 756.900 ;
        RECT 304.950 756.600 307.050 756.900 ;
        RECT 286.950 755.400 307.050 756.600 ;
        RECT 286.950 754.800 289.050 755.400 ;
        RECT 304.950 754.800 307.050 755.400 ;
        RECT 310.950 756.600 313.050 756.900 ;
        RECT 314.400 756.600 315.600 760.950 ;
        RECT 310.950 755.400 315.600 756.600 ;
        RECT 352.950 756.450 355.050 756.900 ;
        RECT 358.950 756.450 361.050 756.900 ;
        RECT 310.950 754.800 313.050 755.400 ;
        RECT 352.950 755.250 361.050 756.450 ;
        RECT 365.400 756.600 366.600 760.950 ;
        RECT 443.400 759.600 444.600 761.100 ;
        RECT 523.950 760.950 526.050 761.400 ;
        RECT 532.950 761.100 535.050 761.400 ;
        RECT 541.950 762.750 544.050 763.200 ;
        RECT 547.950 762.750 550.050 763.200 ;
        RECT 541.950 761.550 550.050 762.750 ;
        RECT 541.950 761.100 544.050 761.550 ;
        RECT 547.950 761.100 550.050 761.550 ;
        RECT 559.950 760.950 562.050 763.050 ;
        RECT 565.950 762.750 568.050 763.200 ;
        RECT 580.950 762.750 583.050 763.200 ;
        RECT 565.950 761.550 583.050 762.750 ;
        RECT 565.950 761.100 568.050 761.550 ;
        RECT 580.950 761.100 583.050 761.550 ;
        RECT 616.950 761.100 619.050 763.200 ;
        RECT 622.950 762.750 625.050 763.200 ;
        RECT 631.950 762.750 634.050 763.200 ;
        RECT 622.950 761.550 634.050 762.750 ;
        RECT 648.000 762.600 652.050 763.050 ;
        RECT 622.950 761.100 625.050 761.550 ;
        RECT 631.950 761.100 634.050 761.550 ;
        RECT 443.400 758.400 453.600 759.600 ;
        RECT 370.950 756.600 373.050 756.900 ;
        RECT 365.400 755.400 373.050 756.600 ;
        RECT 352.950 754.800 355.050 755.250 ;
        RECT 358.950 754.800 361.050 755.250 ;
        RECT 370.950 754.800 373.050 755.400 ;
        RECT 397.950 756.600 400.050 756.900 ;
        RECT 403.950 756.600 406.050 757.050 ;
        RECT 452.400 756.900 453.600 758.400 ;
        RECT 412.950 756.600 415.050 756.900 ;
        RECT 433.950 756.600 436.050 756.900 ;
        RECT 397.950 755.400 436.050 756.600 ;
        RECT 397.950 754.800 400.050 755.400 ;
        RECT 403.950 754.950 406.050 755.400 ;
        RECT 412.950 754.800 415.050 755.400 ;
        RECT 433.950 754.800 436.050 755.400 ;
        RECT 451.950 756.450 454.050 756.900 ;
        RECT 463.950 756.450 466.050 756.900 ;
        RECT 451.950 755.250 466.050 756.450 ;
        RECT 451.950 754.800 454.050 755.250 ;
        RECT 463.950 754.800 466.050 755.250 ;
        RECT 484.950 756.600 487.050 756.900 ;
        RECT 490.950 756.600 493.050 757.050 ;
        RECT 484.950 755.400 493.050 756.600 ;
        RECT 484.950 754.800 487.050 755.400 ;
        RECT 490.950 754.950 493.050 755.400 ;
        RECT 514.950 756.600 517.050 756.900 ;
        RECT 520.950 756.600 523.050 757.050 ;
        RECT 529.950 756.600 532.050 757.050 ;
        RECT 514.950 755.400 532.050 756.600 ;
        RECT 514.950 754.800 517.050 755.400 ;
        RECT 520.950 754.950 523.050 755.400 ;
        RECT 529.950 754.950 532.050 755.400 ;
        RECT 556.950 756.600 559.050 756.900 ;
        RECT 560.400 756.600 561.600 760.950 ;
        RECT 556.950 755.400 561.600 756.600 ;
        RECT 562.950 756.600 565.050 757.050 ;
        RECT 577.950 756.600 580.050 756.900 ;
        RECT 562.950 755.400 580.050 756.600 ;
        RECT 556.950 754.800 559.050 755.400 ;
        RECT 562.950 754.950 565.050 755.400 ;
        RECT 577.950 754.800 580.050 755.400 ;
        RECT 598.950 756.600 601.050 756.900 ;
        RECT 617.400 756.600 618.600 761.100 ;
        RECT 647.400 760.950 652.050 762.600 ;
        RECT 655.950 762.600 658.050 763.050 ;
        RECT 661.950 762.600 664.050 763.200 ;
        RECT 682.950 762.600 685.050 763.200 ;
        RECT 655.950 761.400 664.050 762.600 ;
        RECT 655.950 760.950 658.050 761.400 ;
        RECT 661.950 761.100 664.050 761.400 ;
        RECT 665.400 761.400 685.050 762.600 ;
        RECT 640.950 756.600 643.050 757.050 ;
        RECT 647.400 756.900 648.600 760.950 ;
        RECT 665.400 759.600 666.600 761.400 ;
        RECT 682.950 761.100 685.050 761.400 ;
        RECT 697.950 762.750 700.050 763.200 ;
        RECT 706.950 762.750 709.050 763.200 ;
        RECT 697.950 761.550 709.050 762.750 ;
        RECT 697.950 761.100 700.050 761.550 ;
        RECT 706.950 761.100 709.050 761.550 ;
        RECT 724.950 761.100 727.050 763.200 ;
        RECT 730.950 762.750 733.050 763.200 ;
        RECT 742.950 762.750 745.050 763.200 ;
        RECT 730.950 761.550 745.050 762.750 ;
        RECT 730.950 761.100 733.050 761.550 ;
        RECT 742.950 761.100 745.050 761.550 ;
        RECT 754.950 761.100 757.050 763.200 ;
        RECT 766.950 762.750 769.050 763.200 ;
        RECT 772.950 762.750 775.050 763.200 ;
        RECT 766.950 761.550 775.050 762.750 ;
        RECT 766.950 761.100 769.050 761.550 ;
        RECT 772.950 761.100 775.050 761.550 ;
        RECT 778.950 761.100 781.050 763.200 ;
        RECT 784.950 762.600 787.050 763.050 ;
        RECT 790.950 762.600 793.050 763.200 ;
        RECT 784.950 761.400 793.050 762.600 ;
        RECT 659.400 759.000 666.600 759.600 ;
        RECT 658.950 758.400 666.600 759.000 ;
        RECT 598.950 755.400 643.050 756.600 ;
        RECT 598.950 754.800 601.050 755.400 ;
        RECT 640.950 754.950 643.050 755.400 ;
        RECT 646.950 754.800 649.050 756.900 ;
        RECT 658.950 754.950 661.050 758.400 ;
        RECT 694.950 756.450 697.050 756.900 ;
        RECT 703.950 756.450 706.050 756.900 ;
        RECT 694.950 755.250 706.050 756.450 ;
        RECT 694.950 754.800 697.050 755.250 ;
        RECT 703.950 754.800 706.050 755.250 ;
        RECT 709.950 756.600 712.050 756.900 ;
        RECT 725.400 756.600 726.600 761.100 ;
        RECT 739.950 759.600 742.050 760.050 ;
        RECT 755.400 759.600 756.600 761.100 ;
        RECT 779.400 759.600 780.600 761.100 ;
        RECT 784.950 760.950 787.050 761.400 ;
        RECT 790.950 761.100 793.050 761.400 ;
        RECT 799.950 762.600 802.050 763.200 ;
        RECT 814.950 762.600 817.050 763.200 ;
        RECT 799.950 761.400 817.050 762.600 ;
        RECT 799.950 761.100 802.050 761.400 ;
        RECT 814.950 761.100 817.050 761.400 ;
        RECT 820.950 762.750 823.050 763.200 ;
        RECT 826.950 762.750 829.050 763.200 ;
        RECT 820.950 761.550 829.050 762.750 ;
        RECT 820.950 761.100 823.050 761.550 ;
        RECT 826.950 761.100 829.050 761.550 ;
        RECT 832.950 762.600 835.050 763.050 ;
        RECT 850.950 762.600 853.050 763.050 ;
        RECT 832.950 761.400 853.050 762.600 ;
        RECT 832.950 760.950 835.050 761.400 ;
        RECT 850.950 760.950 853.050 761.400 ;
        RECT 859.950 761.100 862.050 763.200 ;
        RECT 739.950 758.400 780.600 759.600 ;
        RECT 739.950 757.950 742.050 758.400 ;
        RECT 709.950 755.400 726.600 756.600 ;
        RECT 751.950 756.600 754.050 756.900 ;
        RECT 763.950 756.600 766.050 757.050 ;
        RECT 751.950 755.400 766.050 756.600 ;
        RECT 779.400 756.600 780.600 758.400 ;
        RECT 853.950 759.600 856.050 760.050 ;
        RECT 860.400 759.600 861.600 761.100 ;
        RECT 853.950 758.400 861.600 759.600 ;
        RECT 853.950 757.950 856.050 758.400 ;
        RECT 796.950 756.600 799.050 756.900 ;
        RECT 779.400 755.400 799.050 756.600 ;
        RECT 709.950 754.800 712.050 755.400 ;
        RECT 751.950 754.800 754.050 755.400 ;
        RECT 763.950 754.950 766.050 755.400 ;
        RECT 796.950 754.800 799.050 755.400 ;
        RECT 811.950 756.450 814.050 756.900 ;
        RECT 817.950 756.450 820.050 756.900 ;
        RECT 811.950 755.250 820.050 756.450 ;
        RECT 811.950 754.800 814.050 755.250 ;
        RECT 817.950 754.800 820.050 755.250 ;
        RECT 823.950 756.600 826.050 756.900 ;
        RECT 832.950 756.600 835.050 757.050 ;
        RECT 823.950 755.400 835.050 756.600 ;
        RECT 823.950 754.800 826.050 755.400 ;
        RECT 832.950 754.950 835.050 755.400 ;
        RECT 868.950 756.600 871.050 756.900 ;
        RECT 892.950 756.600 895.050 757.050 ;
        RECT 868.950 755.400 895.050 756.600 ;
        RECT 868.950 754.800 871.050 755.400 ;
        RECT 892.950 754.950 895.050 755.400 ;
        RECT 688.950 753.600 691.050 754.050 ;
        RECT 494.400 752.400 576.600 753.600 ;
        RECT 494.400 751.050 495.600 752.400 ;
        RECT 13.950 750.600 16.050 751.050 ;
        RECT 85.950 750.600 88.050 751.050 ;
        RECT 13.950 749.400 88.050 750.600 ;
        RECT 13.950 748.950 16.050 749.400 ;
        RECT 85.950 748.950 88.050 749.400 ;
        RECT 121.950 750.600 124.050 751.050 ;
        RECT 157.950 750.600 160.050 751.050 ;
        RECT 121.950 749.400 160.050 750.600 ;
        RECT 121.950 748.950 124.050 749.400 ;
        RECT 157.950 748.950 160.050 749.400 ;
        RECT 175.950 749.400 180.600 751.050 ;
        RECT 262.950 750.600 265.050 751.050 ;
        RECT 295.950 750.600 298.050 751.050 ;
        RECT 373.950 750.600 376.050 751.050 ;
        RECT 262.950 749.400 376.050 750.600 ;
        RECT 175.950 748.950 180.000 749.400 ;
        RECT 262.950 748.950 265.050 749.400 ;
        RECT 295.950 748.950 298.050 749.400 ;
        RECT 373.950 748.950 376.050 749.400 ;
        RECT 478.950 750.600 481.050 751.050 ;
        RECT 493.950 750.600 496.050 751.050 ;
        RECT 478.950 749.400 496.050 750.600 ;
        RECT 478.950 748.950 481.050 749.400 ;
        RECT 493.950 748.950 496.050 749.400 ;
        RECT 508.950 750.600 511.050 751.050 ;
        RECT 523.950 750.600 526.050 751.050 ;
        RECT 508.950 749.400 526.050 750.600 ;
        RECT 508.950 748.950 511.050 749.400 ;
        RECT 523.950 748.950 526.050 749.400 ;
        RECT 535.950 750.600 538.050 751.050 ;
        RECT 541.950 750.600 544.050 751.050 ;
        RECT 562.950 750.600 565.050 751.050 ;
        RECT 535.950 749.400 565.050 750.600 ;
        RECT 575.400 750.600 576.600 752.400 ;
        RECT 650.400 752.400 691.050 753.600 ;
        RECT 583.950 750.600 586.050 751.050 ;
        RECT 575.400 749.400 586.050 750.600 ;
        RECT 535.950 748.950 538.050 749.400 ;
        RECT 541.950 748.950 544.050 749.400 ;
        RECT 562.950 748.950 565.050 749.400 ;
        RECT 583.950 748.950 586.050 749.400 ;
        RECT 598.950 750.600 601.050 751.050 ;
        RECT 610.950 750.600 613.050 751.050 ;
        RECT 598.950 749.400 613.050 750.600 ;
        RECT 598.950 748.950 601.050 749.400 ;
        RECT 610.950 748.950 613.050 749.400 ;
        RECT 625.950 750.600 628.050 751.050 ;
        RECT 650.400 750.600 651.600 752.400 ;
        RECT 688.950 751.950 691.050 752.400 ;
        RECT 712.950 753.600 715.050 754.050 ;
        RECT 727.950 753.600 730.050 754.050 ;
        RECT 712.950 752.400 730.050 753.600 ;
        RECT 712.950 751.950 715.050 752.400 ;
        RECT 727.950 751.950 730.050 752.400 ;
        RECT 736.950 753.600 739.050 754.050 ;
        RECT 766.950 753.600 769.050 754.050 ;
        RECT 784.950 753.600 787.050 754.050 ;
        RECT 736.950 752.400 787.050 753.600 ;
        RECT 736.950 751.950 739.050 752.400 ;
        RECT 766.950 751.950 769.050 752.400 ;
        RECT 784.950 751.950 787.050 752.400 ;
        RECT 856.950 753.600 859.050 754.050 ;
        RECT 862.950 753.600 865.050 754.050 ;
        RECT 856.950 752.400 865.050 753.600 ;
        RECT 856.950 751.950 859.050 752.400 ;
        RECT 862.950 751.950 865.050 752.400 ;
        RECT 625.950 749.400 651.600 750.600 ;
        RECT 655.950 750.600 658.050 751.050 ;
        RECT 679.950 750.600 682.050 751.050 ;
        RECT 655.950 749.400 682.050 750.600 ;
        RECT 625.950 748.950 628.050 749.400 ;
        RECT 655.950 748.950 658.050 749.400 ;
        RECT 679.950 748.950 682.050 749.400 ;
        RECT 697.950 750.600 700.050 751.050 ;
        RECT 713.400 750.600 714.600 751.950 ;
        RECT 697.950 749.400 714.600 750.600 ;
        RECT 757.950 750.600 760.050 751.050 ;
        RECT 811.950 750.600 814.050 751.050 ;
        RECT 757.950 749.400 814.050 750.600 ;
        RECT 697.950 748.950 700.050 749.400 ;
        RECT 757.950 748.950 760.050 749.400 ;
        RECT 811.950 748.950 814.050 749.400 ;
        RECT 817.950 750.600 820.050 751.050 ;
        RECT 835.950 750.600 838.050 751.050 ;
        RECT 817.950 749.400 838.050 750.600 ;
        RECT 817.950 748.950 820.050 749.400 ;
        RECT 835.950 748.950 838.050 749.400 ;
        RECT 127.950 747.600 130.050 748.050 ;
        RECT 142.950 747.600 145.050 748.050 ;
        RECT 127.950 746.400 145.050 747.600 ;
        RECT 127.950 745.950 130.050 746.400 ;
        RECT 142.950 745.950 145.050 746.400 ;
        RECT 211.950 747.600 214.050 748.050 ;
        RECT 223.950 747.600 226.050 748.050 ;
        RECT 229.950 747.600 232.050 748.050 ;
        RECT 211.950 746.400 232.050 747.600 ;
        RECT 211.950 745.950 214.050 746.400 ;
        RECT 223.950 745.950 226.050 746.400 ;
        RECT 229.950 745.950 232.050 746.400 ;
        RECT 244.950 747.600 247.050 748.050 ;
        RECT 259.950 747.600 262.050 748.050 ;
        RECT 244.950 746.400 262.050 747.600 ;
        RECT 244.950 745.950 247.050 746.400 ;
        RECT 259.950 745.950 262.050 746.400 ;
        RECT 268.950 747.600 271.050 748.050 ;
        RECT 286.950 747.600 289.050 748.050 ;
        RECT 268.950 746.400 289.050 747.600 ;
        RECT 268.950 745.950 271.050 746.400 ;
        RECT 286.950 745.950 289.050 746.400 ;
        RECT 316.950 747.600 319.050 748.050 ;
        RECT 352.950 747.600 355.050 748.050 ;
        RECT 316.950 746.400 355.050 747.600 ;
        RECT 316.950 745.950 319.050 746.400 ;
        RECT 352.950 745.950 355.050 746.400 ;
        RECT 415.950 747.600 418.050 748.050 ;
        RECT 445.950 747.600 448.050 748.050 ;
        RECT 457.950 747.600 460.050 748.050 ;
        RECT 415.950 746.400 460.050 747.600 ;
        RECT 415.950 745.950 418.050 746.400 ;
        RECT 445.950 745.950 448.050 746.400 ;
        RECT 457.950 745.950 460.050 746.400 ;
        RECT 565.950 747.600 568.050 748.050 ;
        RECT 571.800 747.600 573.900 748.050 ;
        RECT 565.950 746.400 573.900 747.600 ;
        RECT 565.950 745.950 568.050 746.400 ;
        RECT 571.800 745.950 573.900 746.400 ;
        RECT 574.950 747.600 577.050 748.050 ;
        RECT 607.950 747.600 610.050 748.050 ;
        RECT 574.950 746.400 610.050 747.600 ;
        RECT 574.950 745.950 577.050 746.400 ;
        RECT 607.950 745.950 610.050 746.400 ;
        RECT 685.950 747.600 688.050 748.050 ;
        RECT 739.950 747.600 742.050 748.050 ;
        RECT 685.950 746.400 742.050 747.600 ;
        RECT 685.950 745.950 688.050 746.400 ;
        RECT 739.950 745.950 742.050 746.400 ;
        RECT 187.950 744.600 190.050 745.050 ;
        RECT 208.950 744.600 211.050 745.050 ;
        RECT 187.950 743.400 211.050 744.600 ;
        RECT 187.950 742.950 190.050 743.400 ;
        RECT 208.950 742.950 211.050 743.400 ;
        RECT 475.950 744.600 478.050 745.050 ;
        RECT 550.950 744.600 553.050 745.050 ;
        RECT 475.950 743.400 553.050 744.600 ;
        RECT 475.950 742.950 478.050 743.400 ;
        RECT 550.950 742.950 553.050 743.400 ;
        RECT 640.950 744.600 643.050 745.050 ;
        RECT 664.950 744.600 667.050 745.050 ;
        RECT 640.950 743.400 667.050 744.600 ;
        RECT 640.950 742.950 643.050 743.400 ;
        RECT 664.950 742.950 667.050 743.400 ;
        RECT 688.950 744.600 691.050 745.050 ;
        RECT 736.950 744.600 739.050 745.050 ;
        RECT 688.950 743.400 739.050 744.600 ;
        RECT 688.950 742.950 691.050 743.400 ;
        RECT 736.950 742.950 739.050 743.400 ;
        RECT 805.950 744.600 808.050 745.050 ;
        RECT 829.950 744.600 832.050 745.050 ;
        RECT 805.950 743.400 832.050 744.600 ;
        RECT 805.950 742.950 808.050 743.400 ;
        RECT 829.950 742.950 832.050 743.400 ;
        RECT 79.950 741.600 82.050 742.050 ;
        RECT 94.950 741.600 97.050 742.050 ;
        RECT 79.950 740.400 97.050 741.600 ;
        RECT 79.950 739.950 82.050 740.400 ;
        RECT 94.950 739.950 97.050 740.400 ;
        RECT 145.950 741.600 148.050 742.050 ;
        RECT 151.950 741.600 154.050 742.050 ;
        RECT 145.950 740.400 154.050 741.600 ;
        RECT 145.950 739.950 148.050 740.400 ;
        RECT 151.950 739.950 154.050 740.400 ;
        RECT 274.950 741.600 277.050 742.050 ;
        RECT 427.950 741.600 430.050 742.050 ;
        RECT 274.950 740.400 430.050 741.600 ;
        RECT 274.950 739.950 277.050 740.400 ;
        RECT 427.950 739.950 430.050 740.400 ;
        RECT 439.950 741.600 442.050 742.050 ;
        RECT 472.950 741.600 475.050 742.050 ;
        RECT 439.950 740.400 475.050 741.600 ;
        RECT 439.950 739.950 442.050 740.400 ;
        RECT 472.950 739.950 475.050 740.400 ;
        RECT 478.950 741.600 481.050 742.050 ;
        RECT 520.950 741.600 523.050 742.050 ;
        RECT 478.950 740.400 523.050 741.600 ;
        RECT 478.950 739.950 481.050 740.400 ;
        RECT 520.950 739.950 523.050 740.400 ;
        RECT 553.950 741.600 556.050 742.050 ;
        RECT 589.950 741.600 592.050 742.050 ;
        RECT 553.950 740.400 592.050 741.600 ;
        RECT 553.950 739.950 556.050 740.400 ;
        RECT 589.950 739.950 592.050 740.400 ;
        RECT 622.950 741.600 625.050 742.050 ;
        RECT 637.950 741.600 640.050 742.050 ;
        RECT 622.950 740.400 640.050 741.600 ;
        RECT 622.950 739.950 625.050 740.400 ;
        RECT 637.950 739.950 640.050 740.400 ;
        RECT 709.950 741.600 712.050 742.050 ;
        RECT 715.950 741.600 718.050 742.050 ;
        RECT 709.950 740.400 718.050 741.600 ;
        RECT 709.950 739.950 712.050 740.400 ;
        RECT 715.950 739.950 718.050 740.400 ;
        RECT 772.950 741.600 775.050 742.050 ;
        RECT 832.950 741.600 835.050 742.050 ;
        RECT 772.950 740.400 835.050 741.600 ;
        RECT 772.950 739.950 775.050 740.400 ;
        RECT 832.950 739.950 835.050 740.400 ;
        RECT 847.950 741.600 850.050 742.050 ;
        RECT 865.950 741.600 868.050 742.050 ;
        RECT 847.950 740.400 868.050 741.600 ;
        RECT 847.950 739.950 850.050 740.400 ;
        RECT 865.950 739.950 868.050 740.400 ;
        RECT 97.950 738.600 100.050 739.050 ;
        RECT 100.950 738.600 103.050 739.050 ;
        RECT 148.950 738.600 151.050 739.050 ;
        RECT 97.950 737.400 151.050 738.600 ;
        RECT 97.950 736.950 100.050 737.400 ;
        RECT 100.950 736.950 103.050 737.400 ;
        RECT 148.950 736.950 151.050 737.400 ;
        RECT 220.950 738.600 223.050 739.050 ;
        RECT 235.950 738.600 238.050 739.050 ;
        RECT 220.950 737.400 238.050 738.600 ;
        RECT 220.950 736.950 223.050 737.400 ;
        RECT 235.950 736.950 238.050 737.400 ;
        RECT 532.950 738.600 535.050 739.050 ;
        RECT 604.950 738.600 607.050 739.050 ;
        RECT 532.950 737.400 607.050 738.600 ;
        RECT 532.950 736.950 535.050 737.400 ;
        RECT 604.950 736.950 607.050 737.400 ;
        RECT 610.950 738.600 613.050 739.050 ;
        RECT 631.950 738.600 634.050 739.050 ;
        RECT 610.950 737.400 634.050 738.600 ;
        RECT 610.950 736.950 613.050 737.400 ;
        RECT 631.950 736.950 634.050 737.400 ;
        RECT 775.950 738.600 778.050 739.050 ;
        RECT 775.950 737.400 825.600 738.600 ;
        RECT 775.950 736.950 778.050 737.400 ;
        RECT 824.400 736.050 825.600 737.400 ;
        RECT 76.950 735.600 79.050 736.050 ;
        RECT 85.950 735.600 88.050 736.050 ;
        RECT 76.950 734.400 88.050 735.600 ;
        RECT 76.950 733.950 79.050 734.400 ;
        RECT 85.950 733.950 88.050 734.400 ;
        RECT 115.950 735.600 118.050 736.050 ;
        RECT 148.950 735.600 151.050 735.900 ;
        RECT 115.950 734.400 151.050 735.600 ;
        RECT 115.950 733.950 118.050 734.400 ;
        RECT 148.950 733.800 151.050 734.400 ;
        RECT 268.950 735.600 271.050 736.050 ;
        RECT 328.950 735.600 331.050 736.050 ;
        RECT 334.950 735.600 337.050 736.050 ;
        RECT 376.950 735.600 379.050 736.050 ;
        RECT 268.950 734.400 379.050 735.600 ;
        RECT 268.950 733.950 271.050 734.400 ;
        RECT 328.950 733.950 331.050 734.400 ;
        RECT 334.950 733.950 337.050 734.400 ;
        RECT 376.950 733.950 379.050 734.400 ;
        RECT 388.950 735.600 391.050 736.050 ;
        RECT 460.950 735.600 463.050 736.050 ;
        RECT 388.950 734.400 463.050 735.600 ;
        RECT 388.950 733.950 391.050 734.400 ;
        RECT 460.950 733.950 463.050 734.400 ;
        RECT 472.950 735.600 475.050 736.050 ;
        RECT 550.950 735.600 553.050 736.050 ;
        RECT 559.950 735.600 562.050 736.050 ;
        RECT 472.950 734.400 495.600 735.600 ;
        RECT 472.950 733.950 475.050 734.400 ;
        RECT 31.950 732.600 34.050 733.050 ;
        RECT 64.950 732.600 67.050 733.050 ;
        RECT 73.950 732.600 76.050 733.050 ;
        RECT 31.950 731.400 76.050 732.600 ;
        RECT 31.950 730.950 34.050 731.400 ;
        RECT 64.950 730.950 67.050 731.400 ;
        RECT 73.950 730.950 76.050 731.400 ;
        RECT 181.950 730.950 184.050 733.050 ;
        RECT 494.400 732.600 495.600 734.400 ;
        RECT 550.950 734.400 562.050 735.600 ;
        RECT 550.950 733.950 553.050 734.400 ;
        RECT 559.950 733.950 562.050 734.400 ;
        RECT 781.950 735.600 784.050 736.050 ;
        RECT 793.950 735.600 796.050 736.050 ;
        RECT 811.950 735.600 814.050 736.050 ;
        RECT 781.950 734.400 814.050 735.600 ;
        RECT 781.950 733.950 784.050 734.400 ;
        RECT 793.950 733.950 796.050 734.400 ;
        RECT 811.950 733.950 814.050 734.400 ;
        RECT 823.950 735.600 826.050 736.050 ;
        RECT 859.950 735.600 862.050 736.050 ;
        RECT 823.950 734.400 862.050 735.600 ;
        RECT 823.950 733.950 826.050 734.400 ;
        RECT 859.950 733.950 862.050 734.400 ;
        RECT 496.950 732.600 499.050 733.050 ;
        RECT 541.950 732.600 544.050 733.050 ;
        RECT 494.400 731.400 544.050 732.600 ;
        RECT 496.950 730.950 499.050 731.400 ;
        RECT 541.950 730.950 544.050 731.400 ;
        RECT 646.950 732.600 649.050 733.050 ;
        RECT 652.950 732.600 655.050 733.050 ;
        RECT 646.950 731.400 655.050 732.600 ;
        RECT 646.950 730.950 649.050 731.400 ;
        RECT 652.950 730.950 655.050 731.400 ;
        RECT 670.950 732.600 673.050 733.050 ;
        RECT 706.950 732.600 709.050 733.050 ;
        RECT 670.950 731.400 709.050 732.600 ;
        RECT 670.950 730.950 673.050 731.400 ;
        RECT 706.950 730.950 709.050 731.400 ;
        RECT 850.950 732.600 853.050 733.050 ;
        RECT 895.950 732.600 898.050 733.050 ;
        RECT 850.950 731.400 898.050 732.600 ;
        RECT 850.950 730.950 853.050 731.400 ;
        RECT 895.950 730.950 898.050 731.400 ;
        RECT 7.950 729.600 12.000 730.050 ;
        RECT 55.950 729.600 58.050 730.200 ;
        RECT 103.950 730.050 106.050 730.500 ;
        RECT 136.950 730.050 139.050 730.500 ;
        RECT 61.950 729.600 64.050 730.050 ;
        RECT 7.950 727.950 12.600 729.600 ;
        RECT 55.950 728.400 64.050 729.600 ;
        RECT 103.950 728.850 139.050 730.050 ;
        RECT 103.950 728.400 106.050 728.850 ;
        RECT 136.950 728.400 139.050 728.850 ;
        RECT 145.950 729.600 148.050 730.050 ;
        RECT 145.950 728.400 156.600 729.600 ;
        RECT 55.950 728.100 58.050 728.400 ;
        RECT 61.950 727.950 64.050 728.400 ;
        RECT 145.950 727.950 148.050 728.400 ;
        RECT 11.400 723.900 12.600 727.950 ;
        RECT 10.950 721.800 13.050 723.900 ;
        RECT 16.950 723.600 19.050 723.900 ;
        RECT 34.950 723.600 37.050 723.900 ;
        RECT 16.950 722.400 37.050 723.600 ;
        RECT 16.950 721.800 19.050 722.400 ;
        RECT 34.950 721.800 37.050 722.400 ;
        RECT 115.950 723.600 118.050 724.050 ;
        RECT 155.400 723.900 156.600 728.400 ;
        RECT 157.950 728.100 160.050 730.200 ;
        RECT 115.950 722.400 124.050 723.600 ;
        RECT 115.950 721.950 118.050 722.400 ;
        RECT 121.950 721.500 124.050 722.400 ;
        RECT 154.950 721.800 157.050 723.900 ;
        RECT 158.400 721.050 159.600 728.100 ;
        RECT 182.400 723.600 183.600 730.950 ;
        RECT 199.950 729.750 202.050 730.200 ;
        RECT 214.950 729.750 217.050 730.200 ;
        RECT 199.950 728.550 217.050 729.750 ;
        RECT 199.950 728.100 202.050 728.550 ;
        RECT 214.950 728.100 217.050 728.550 ;
        RECT 241.950 729.600 244.050 730.200 ;
        RECT 253.950 729.600 256.050 730.200 ;
        RECT 280.950 729.600 283.050 730.200 ;
        RECT 241.950 728.400 283.050 729.600 ;
        RECT 241.950 728.100 244.050 728.400 ;
        RECT 253.950 728.100 256.050 728.400 ;
        RECT 280.950 728.100 283.050 728.400 ;
        RECT 286.950 729.600 289.050 730.200 ;
        RECT 310.950 729.600 313.050 730.200 ;
        RECT 346.950 729.600 349.050 730.200 ;
        RECT 286.950 728.400 349.050 729.600 ;
        RECT 286.950 728.100 289.050 728.400 ;
        RECT 310.950 728.100 313.050 728.400 ;
        RECT 346.950 728.100 349.050 728.400 ;
        RECT 358.950 729.750 361.050 730.200 ;
        RECT 367.950 729.750 370.050 730.200 ;
        RECT 358.950 728.550 370.050 729.750 ;
        RECT 358.950 728.100 361.050 728.550 ;
        RECT 367.950 728.100 370.050 728.550 ;
        RECT 385.950 729.750 388.050 730.200 ;
        RECT 391.950 729.750 394.050 730.200 ;
        RECT 385.950 728.550 394.050 729.750 ;
        RECT 385.950 728.100 388.050 728.550 ;
        RECT 391.950 728.100 394.050 728.550 ;
        RECT 397.950 729.600 400.050 730.200 ;
        RECT 415.950 729.600 418.050 730.200 ;
        RECT 397.950 728.400 418.050 729.600 ;
        RECT 397.950 728.100 400.050 728.400 ;
        RECT 415.950 728.100 418.050 728.400 ;
        RECT 466.950 729.750 469.050 730.200 ;
        RECT 478.950 729.750 481.050 730.200 ;
        RECT 466.950 728.550 481.050 729.750 ;
        RECT 466.950 728.100 469.050 728.550 ;
        RECT 478.950 728.100 481.050 728.550 ;
        RECT 484.950 729.750 487.050 730.200 ;
        RECT 490.950 729.750 493.050 730.200 ;
        RECT 484.950 728.550 493.050 729.750 ;
        RECT 484.950 728.100 487.050 728.550 ;
        RECT 490.950 728.100 493.050 728.550 ;
        RECT 511.950 729.600 514.050 730.050 ;
        RECT 526.950 729.600 529.050 730.050 ;
        RECT 511.950 728.400 529.050 729.600 ;
        RECT 511.950 727.950 514.050 728.400 ;
        RECT 526.950 727.950 529.050 728.400 ;
        RECT 682.950 729.600 685.050 730.200 ;
        RECT 691.950 729.750 694.050 730.200 ;
        RECT 700.950 729.750 703.050 730.200 ;
        RECT 691.950 729.600 703.050 729.750 ;
        RECT 682.950 728.550 703.050 729.600 ;
        RECT 682.950 728.400 694.050 728.550 ;
        RECT 682.950 728.100 685.050 728.400 ;
        RECT 691.950 728.100 694.050 728.400 ;
        RECT 700.950 728.100 703.050 728.550 ;
        RECT 727.950 729.600 730.050 730.200 ;
        RECT 733.950 729.600 736.050 730.200 ;
        RECT 742.950 729.600 745.050 730.050 ;
        RECT 748.950 729.600 751.050 730.200 ;
        RECT 766.950 729.600 769.050 730.200 ;
        RECT 787.950 729.600 790.050 730.200 ;
        RECT 727.950 728.400 732.600 729.600 ;
        RECT 727.950 728.100 730.050 728.400 ;
        RECT 238.950 723.600 241.050 723.900 ;
        RECT 256.950 723.600 259.050 723.900 ;
        RECT 181.950 721.500 184.050 723.600 ;
        RECT 238.950 722.400 259.050 723.600 ;
        RECT 238.950 721.800 241.050 722.400 ;
        RECT 256.950 721.800 259.050 722.400 ;
        RECT 262.950 723.600 265.050 723.900 ;
        RECT 271.950 723.600 274.050 724.050 ;
        RECT 262.950 722.400 274.050 723.600 ;
        RECT 262.950 721.800 265.050 722.400 ;
        RECT 271.950 721.950 274.050 722.400 ;
        RECT 289.950 723.600 292.050 723.900 ;
        RECT 307.950 723.600 310.050 723.900 ;
        RECT 289.950 722.400 310.050 723.600 ;
        RECT 289.950 721.800 292.050 722.400 ;
        RECT 307.950 721.800 310.050 722.400 ;
        RECT 313.950 723.600 316.050 723.900 ;
        RECT 328.950 723.600 331.050 723.900 ;
        RECT 343.950 723.600 346.050 723.900 ;
        RECT 313.950 722.400 346.050 723.600 ;
        RECT 313.950 721.800 316.050 722.400 ;
        RECT 328.950 721.800 331.050 722.400 ;
        RECT 343.950 721.800 346.050 722.400 ;
        RECT 349.950 723.600 352.050 723.900 ;
        RECT 370.950 723.600 373.050 723.900 ;
        RECT 349.950 722.400 373.050 723.600 ;
        RECT 349.950 721.800 352.050 722.400 ;
        RECT 370.950 721.800 373.050 722.400 ;
        RECT 469.950 723.450 472.050 723.900 ;
        RECT 481.950 723.450 484.050 723.900 ;
        RECT 469.950 722.250 484.050 723.450 ;
        RECT 469.950 721.800 472.050 722.250 ;
        RECT 481.950 721.800 484.050 722.250 ;
        RECT 607.950 721.800 610.050 723.900 ;
        RECT 613.950 723.600 616.050 723.900 ;
        RECT 631.950 723.600 634.050 723.900 ;
        RECT 652.950 723.600 655.050 723.900 ;
        RECT 613.950 722.400 655.050 723.600 ;
        RECT 613.950 721.800 616.050 722.400 ;
        RECT 631.950 721.800 634.050 722.400 ;
        RECT 652.950 721.800 655.050 722.400 ;
        RECT 703.950 723.600 706.050 723.900 ;
        RECT 724.950 723.600 727.050 723.900 ;
        RECT 703.950 722.400 727.050 723.600 ;
        RECT 731.400 723.600 732.600 728.400 ;
        RECT 733.950 728.400 769.050 729.600 ;
        RECT 733.950 728.100 736.050 728.400 ;
        RECT 742.950 727.950 745.050 728.400 ;
        RECT 748.950 728.100 751.050 728.400 ;
        RECT 766.950 728.100 769.050 728.400 ;
        RECT 770.400 728.400 790.050 729.600 ;
        RECT 760.950 726.600 763.050 727.050 ;
        RECT 770.400 726.600 771.600 728.400 ;
        RECT 787.950 728.100 790.050 728.400 ;
        RECT 826.950 729.750 829.050 730.200 ;
        RECT 838.950 729.750 841.050 730.200 ;
        RECT 826.950 728.550 841.050 729.750 ;
        RECT 826.950 728.100 829.050 728.550 ;
        RECT 838.950 728.100 841.050 728.550 ;
        RECT 844.950 729.600 847.050 730.200 ;
        RECT 874.950 729.600 877.050 730.050 ;
        RECT 844.950 728.400 877.050 729.600 ;
        RECT 844.950 728.100 847.050 728.400 ;
        RECT 760.950 725.400 771.600 726.600 ;
        RECT 760.950 724.950 763.050 725.400 ;
        RECT 736.950 723.600 739.050 724.050 ;
        RECT 731.400 722.400 739.050 723.600 ;
        RECT 703.950 721.800 706.050 722.400 ;
        RECT 724.950 721.800 727.050 722.400 ;
        RECT 736.950 721.950 739.050 722.400 ;
        RECT 814.950 723.600 817.050 723.900 ;
        RECT 823.950 723.600 826.050 724.050 ;
        RECT 869.400 723.900 870.600 728.400 ;
        RECT 874.950 727.950 877.050 728.400 ;
        RECT 814.950 722.400 826.050 723.600 ;
        RECT 814.950 721.800 817.050 722.400 ;
        RECT 823.950 721.950 826.050 722.400 ;
        RECT 868.950 721.800 871.050 723.900 ;
        RECT 70.950 720.600 73.050 721.050 ;
        RECT 94.950 720.600 97.050 721.050 ;
        RECT 70.950 719.400 97.050 720.600 ;
        RECT 70.950 718.950 73.050 719.400 ;
        RECT 94.950 718.950 97.050 719.400 ;
        RECT 157.950 718.950 160.050 721.050 ;
        RECT 283.950 720.600 286.050 721.050 ;
        RECT 313.950 720.600 316.050 721.050 ;
        RECT 283.950 719.400 316.050 720.600 ;
        RECT 283.950 718.950 286.050 719.400 ;
        RECT 313.950 718.950 316.050 719.400 ;
        RECT 424.950 720.600 427.050 721.050 ;
        RECT 433.950 720.600 436.050 721.050 ;
        RECT 424.950 719.400 436.050 720.600 ;
        RECT 424.950 718.950 427.050 719.400 ;
        RECT 433.950 718.950 436.050 719.400 ;
        RECT 562.950 720.600 565.050 721.050 ;
        RECT 571.950 720.600 574.050 721.050 ;
        RECT 608.400 720.600 609.600 721.800 ;
        RECT 562.950 719.400 609.600 720.600 ;
        RECT 685.950 720.600 688.050 721.050 ;
        RECT 703.950 720.600 706.050 721.050 ;
        RECT 685.950 719.400 706.050 720.600 ;
        RECT 562.950 718.950 565.050 719.400 ;
        RECT 571.950 718.950 574.050 719.400 ;
        RECT 685.950 718.950 688.050 719.400 ;
        RECT 703.950 718.950 706.050 719.400 ;
        RECT 802.950 720.600 805.050 721.050 ;
        RECT 841.950 720.600 844.050 721.050 ;
        RECT 802.950 719.400 844.050 720.600 ;
        RECT 802.950 718.950 805.050 719.400 ;
        RECT 841.950 718.950 844.050 719.400 ;
        RECT 112.950 717.600 115.050 718.050 ;
        RECT 121.950 717.600 124.050 718.050 ;
        RECT 130.950 717.600 133.050 718.050 ;
        RECT 190.950 717.600 193.050 718.050 ;
        RECT 112.950 716.400 193.050 717.600 ;
        RECT 112.950 715.950 115.050 716.400 ;
        RECT 121.950 715.950 124.050 716.400 ;
        RECT 130.950 715.950 133.050 716.400 ;
        RECT 190.950 715.950 193.050 716.400 ;
        RECT 196.950 717.600 199.050 718.050 ;
        RECT 211.950 717.600 214.050 718.050 ;
        RECT 196.950 716.400 214.050 717.600 ;
        RECT 196.950 715.950 199.050 716.400 ;
        RECT 211.950 715.950 214.050 716.400 ;
        RECT 235.950 717.600 238.050 718.050 ;
        RECT 247.950 717.600 250.050 718.050 ;
        RECT 235.950 716.400 250.050 717.600 ;
        RECT 235.950 715.950 238.050 716.400 ;
        RECT 247.950 715.950 250.050 716.400 ;
        RECT 334.950 717.600 337.050 718.050 ;
        RECT 376.950 717.600 379.050 718.050 ;
        RECT 334.950 716.400 379.050 717.600 ;
        RECT 334.950 715.950 337.050 716.400 ;
        RECT 376.950 715.950 379.050 716.400 ;
        RECT 385.950 717.600 388.050 718.050 ;
        RECT 394.950 717.600 397.050 718.050 ;
        RECT 385.950 716.400 397.050 717.600 ;
        RECT 385.950 715.950 388.050 716.400 ;
        RECT 394.950 715.950 397.050 716.400 ;
        RECT 475.950 717.600 478.050 718.050 ;
        RECT 493.950 717.600 496.050 718.050 ;
        RECT 475.950 716.400 496.050 717.600 ;
        RECT 475.950 715.950 478.050 716.400 ;
        RECT 493.950 715.950 496.050 716.400 ;
        RECT 679.950 717.600 682.050 718.050 ;
        RECT 697.950 717.600 700.050 718.050 ;
        RECT 769.950 717.600 772.050 718.050 ;
        RECT 679.950 716.400 772.050 717.600 ;
        RECT 679.950 715.950 682.050 716.400 ;
        RECT 697.950 715.950 700.050 716.400 ;
        RECT 769.950 715.950 772.050 716.400 ;
        RECT 805.950 717.600 808.050 718.050 ;
        RECT 862.950 717.600 865.050 718.050 ;
        RECT 805.950 716.400 865.050 717.600 ;
        RECT 805.950 715.950 808.050 716.400 ;
        RECT 862.950 715.950 865.050 716.400 ;
        RECT 154.950 714.600 157.050 715.050 ;
        RECT 175.950 714.600 178.050 715.050 ;
        RECT 154.950 713.400 178.050 714.600 ;
        RECT 154.950 712.950 157.050 713.400 ;
        RECT 175.950 712.950 178.050 713.400 ;
        RECT 382.950 714.600 385.050 715.050 ;
        RECT 418.950 714.600 421.050 715.050 ;
        RECT 382.950 713.400 421.050 714.600 ;
        RECT 382.950 712.950 385.050 713.400 ;
        RECT 418.950 712.950 421.050 713.400 ;
        RECT 463.950 714.600 466.050 715.050 ;
        RECT 472.950 714.600 475.050 715.050 ;
        RECT 463.950 713.400 475.050 714.600 ;
        RECT 463.950 712.950 466.050 713.400 ;
        RECT 472.950 712.950 475.050 713.400 ;
        RECT 517.950 714.600 520.050 715.050 ;
        RECT 559.950 714.600 562.050 715.050 ;
        RECT 565.950 714.600 568.050 715.050 ;
        RECT 517.950 713.400 568.050 714.600 ;
        RECT 517.950 712.950 520.050 713.400 ;
        RECT 559.950 712.950 562.050 713.400 ;
        RECT 565.950 712.950 568.050 713.400 ;
        RECT 571.950 714.600 574.050 715.050 ;
        RECT 607.950 714.600 610.050 715.050 ;
        RECT 571.950 713.400 610.050 714.600 ;
        RECT 571.950 712.950 574.050 713.400 ;
        RECT 607.950 712.950 610.050 713.400 ;
        RECT 721.950 714.600 724.050 715.050 ;
        RECT 790.950 714.600 793.050 715.050 ;
        RECT 721.950 713.400 793.050 714.600 ;
        RECT 721.950 712.950 724.050 713.400 ;
        RECT 790.950 712.950 793.050 713.400 ;
        RECT 370.950 711.600 373.050 712.050 ;
        RECT 391.950 711.600 394.050 712.050 ;
        RECT 370.950 710.400 394.050 711.600 ;
        RECT 370.950 709.950 373.050 710.400 ;
        RECT 391.950 709.950 394.050 710.400 ;
        RECT 421.950 711.600 424.050 712.050 ;
        RECT 436.950 711.600 439.050 712.050 ;
        RECT 421.950 710.400 439.050 711.600 ;
        RECT 421.950 709.950 424.050 710.400 ;
        RECT 436.950 709.950 439.050 710.400 ;
        RECT 520.950 711.600 523.050 712.050 ;
        RECT 532.950 711.600 535.050 712.050 ;
        RECT 520.950 710.400 535.050 711.600 ;
        RECT 791.400 711.600 792.600 712.950 ;
        RECT 808.950 711.600 811.050 712.050 ;
        RECT 791.400 710.400 811.050 711.600 ;
        RECT 520.950 709.950 523.050 710.400 ;
        RECT 532.950 709.950 535.050 710.400 ;
        RECT 808.950 709.950 811.050 710.400 ;
        RECT 130.950 708.600 133.050 709.050 ;
        RECT 136.950 708.600 139.050 709.050 ;
        RECT 130.950 707.400 139.050 708.600 ;
        RECT 130.950 706.950 133.050 707.400 ;
        RECT 136.950 706.950 139.050 707.400 ;
        RECT 451.950 708.600 454.050 709.050 ;
        RECT 472.950 708.600 475.050 709.050 ;
        RECT 451.950 707.400 475.050 708.600 ;
        RECT 451.950 706.950 454.050 707.400 ;
        RECT 472.950 706.950 475.050 707.400 ;
        RECT 538.950 708.600 541.050 709.050 ;
        RECT 589.950 708.600 592.050 709.050 ;
        RECT 598.950 708.600 601.050 709.050 ;
        RECT 538.950 707.400 601.050 708.600 ;
        RECT 538.950 706.950 541.050 707.400 ;
        RECT 589.950 706.950 592.050 707.400 ;
        RECT 598.950 706.950 601.050 707.400 ;
        RECT 610.950 708.600 613.050 709.050 ;
        RECT 622.950 708.600 625.050 709.050 ;
        RECT 610.950 707.400 625.050 708.600 ;
        RECT 610.950 706.950 613.050 707.400 ;
        RECT 622.950 706.950 625.050 707.400 ;
        RECT 631.950 708.600 634.050 709.050 ;
        RECT 655.950 708.600 658.050 709.050 ;
        RECT 631.950 707.400 658.050 708.600 ;
        RECT 631.950 706.950 634.050 707.400 ;
        RECT 655.950 706.950 658.050 707.400 ;
        RECT 832.950 708.600 835.050 709.050 ;
        RECT 886.950 708.600 889.050 709.050 ;
        RECT 832.950 707.400 889.050 708.600 ;
        RECT 832.950 706.950 835.050 707.400 ;
        RECT 886.950 706.950 889.050 707.400 ;
        RECT 490.950 705.600 493.050 706.050 ;
        RECT 539.400 705.600 540.600 706.950 ;
        RECT 490.950 704.400 540.600 705.600 ;
        RECT 544.950 705.600 547.050 706.050 ;
        RECT 550.950 705.600 553.050 706.050 ;
        RECT 583.950 705.600 586.050 706.050 ;
        RECT 544.950 704.400 586.050 705.600 ;
        RECT 490.950 703.950 493.050 704.400 ;
        RECT 544.950 703.950 547.050 704.400 ;
        RECT 550.950 703.950 553.050 704.400 ;
        RECT 583.950 703.950 586.050 704.400 ;
        RECT 622.950 705.600 625.050 705.900 ;
        RECT 658.800 705.600 660.900 706.050 ;
        RECT 622.950 704.400 660.900 705.600 ;
        RECT 622.950 703.800 625.050 704.400 ;
        RECT 658.800 703.950 660.900 704.400 ;
        RECT 661.950 705.600 664.050 706.050 ;
        RECT 661.950 704.400 714.600 705.600 ;
        RECT 661.950 703.950 664.050 704.400 ;
        RECT 355.950 702.600 358.050 703.050 ;
        RECT 505.950 702.600 508.050 703.050 ;
        RECT 538.800 702.600 540.900 702.900 ;
        RECT 355.950 701.400 414.600 702.600 ;
        RECT 355.950 700.950 358.050 701.400 ;
        RECT 413.400 700.050 414.600 701.400 ;
        RECT 505.950 701.400 540.900 702.600 ;
        RECT 505.950 700.950 508.050 701.400 ;
        RECT 538.800 700.800 540.900 701.400 ;
        RECT 541.950 702.600 544.050 703.050 ;
        RECT 553.950 702.600 556.050 703.050 ;
        RECT 541.950 701.400 556.050 702.600 ;
        RECT 541.950 700.950 544.050 701.400 ;
        RECT 553.950 700.950 556.050 701.400 ;
        RECT 586.950 702.600 589.050 703.050 ;
        RECT 685.950 702.600 688.050 703.050 ;
        RECT 691.950 702.600 694.050 703.050 ;
        RECT 586.950 701.400 694.050 702.600 ;
        RECT 713.400 702.600 714.600 704.400 ;
        RECT 724.950 702.600 727.050 703.050 ;
        RECT 713.400 701.400 727.050 702.600 ;
        RECT 586.950 700.950 589.050 701.400 ;
        RECT 685.950 700.950 688.050 701.400 ;
        RECT 691.950 700.950 694.050 701.400 ;
        RECT 724.950 700.950 727.050 701.400 ;
        RECT 736.950 702.600 739.050 703.050 ;
        RECT 793.950 702.600 796.050 703.050 ;
        RECT 826.950 702.600 829.050 703.050 ;
        RECT 736.950 701.400 829.050 702.600 ;
        RECT 736.950 700.950 739.050 701.400 ;
        RECT 793.950 700.950 796.050 701.400 ;
        RECT 826.950 700.950 829.050 701.400 ;
        RECT 19.950 699.600 22.050 700.050 ;
        RECT 43.950 699.600 46.050 700.050 ;
        RECT 52.950 699.600 55.050 700.050 ;
        RECT 19.950 698.400 55.050 699.600 ;
        RECT 19.950 697.950 22.050 698.400 ;
        RECT 43.950 697.950 46.050 698.400 ;
        RECT 52.950 697.950 55.050 698.400 ;
        RECT 328.950 699.600 331.050 700.050 ;
        RECT 397.950 699.600 400.050 700.050 ;
        RECT 328.950 698.400 400.050 699.600 ;
        RECT 328.950 697.950 331.050 698.400 ;
        RECT 397.950 697.950 400.050 698.400 ;
        RECT 412.950 699.600 415.050 700.050 ;
        RECT 427.950 699.600 430.050 700.050 ;
        RECT 571.950 699.600 574.050 700.050 ;
        RECT 412.950 698.400 574.050 699.600 ;
        RECT 412.950 697.950 415.050 698.400 ;
        RECT 427.950 697.950 430.050 698.400 ;
        RECT 571.950 697.950 574.050 698.400 ;
        RECT 709.950 699.600 712.050 700.050 ;
        RECT 730.950 699.600 733.050 700.050 ;
        RECT 709.950 698.400 733.050 699.600 ;
        RECT 709.950 697.950 712.050 698.400 ;
        RECT 730.950 697.950 733.050 698.400 ;
        RECT 760.950 699.600 763.050 700.050 ;
        RECT 775.950 699.600 778.050 700.050 ;
        RECT 760.950 698.400 778.050 699.600 ;
        RECT 760.950 697.950 763.050 698.400 ;
        RECT 775.950 697.950 778.050 698.400 ;
        RECT 247.950 696.600 250.050 697.050 ;
        RECT 322.950 696.600 325.050 697.050 ;
        RECT 247.950 695.400 325.050 696.600 ;
        RECT 247.950 694.950 250.050 695.400 ;
        RECT 322.950 694.950 325.050 695.400 ;
        RECT 373.950 696.600 376.050 697.050 ;
        RECT 388.950 696.600 391.050 697.050 ;
        RECT 406.950 696.600 409.050 697.050 ;
        RECT 373.950 695.400 409.050 696.600 ;
        RECT 373.950 694.950 376.050 695.400 ;
        RECT 388.950 694.950 391.050 695.400 ;
        RECT 406.950 694.950 409.050 695.400 ;
        RECT 448.950 696.600 451.050 697.050 ;
        RECT 457.950 696.600 460.050 697.050 ;
        RECT 448.950 695.400 460.050 696.600 ;
        RECT 448.950 694.950 451.050 695.400 ;
        RECT 457.950 694.950 460.050 695.400 ;
        RECT 472.950 696.600 475.050 697.050 ;
        RECT 640.950 696.600 643.050 697.050 ;
        RECT 472.950 695.400 643.050 696.600 ;
        RECT 472.950 694.950 475.050 695.400 ;
        RECT 640.950 694.950 643.050 695.400 ;
        RECT 691.950 696.600 694.050 697.050 ;
        RECT 715.800 696.600 717.900 697.050 ;
        RECT 691.950 695.400 717.900 696.600 ;
        RECT 691.950 694.950 694.050 695.400 ;
        RECT 715.800 694.950 717.900 695.400 ;
        RECT 718.950 696.600 721.050 697.050 ;
        RECT 736.950 696.600 739.050 697.050 ;
        RECT 718.950 695.400 739.050 696.600 ;
        RECT 718.950 694.950 721.050 695.400 ;
        RECT 736.950 694.950 739.050 695.400 ;
        RECT 13.950 693.600 16.050 694.050 ;
        RECT 46.950 693.600 49.050 694.050 ;
        RECT 13.950 692.400 49.050 693.600 ;
        RECT 13.950 691.950 16.050 692.400 ;
        RECT 46.950 691.950 49.050 692.400 ;
        RECT 64.950 693.600 67.050 694.050 ;
        RECT 76.950 693.600 79.050 694.050 ;
        RECT 64.950 692.400 79.050 693.600 ;
        RECT 64.950 691.950 67.050 692.400 ;
        RECT 76.950 691.950 79.050 692.400 ;
        RECT 232.950 693.600 235.050 694.050 ;
        RECT 274.950 693.600 277.050 694.050 ;
        RECT 232.950 692.400 277.050 693.600 ;
        RECT 232.950 691.950 235.050 692.400 ;
        RECT 274.950 691.950 277.050 692.400 ;
        RECT 310.950 693.600 313.050 694.050 ;
        RECT 325.950 693.600 328.050 694.050 ;
        RECT 331.950 693.600 334.050 694.050 ;
        RECT 310.950 692.400 334.050 693.600 ;
        RECT 310.950 691.950 313.050 692.400 ;
        RECT 325.950 691.950 328.050 692.400 ;
        RECT 331.950 691.950 334.050 692.400 ;
        RECT 361.950 693.600 364.050 694.050 ;
        RECT 421.950 693.600 424.050 693.900 ;
        RECT 361.950 692.400 424.050 693.600 ;
        RECT 361.950 691.950 364.050 692.400 ;
        RECT 421.950 691.800 424.050 692.400 ;
        RECT 514.950 693.600 517.050 694.050 ;
        RECT 544.950 693.600 547.050 694.050 ;
        RECT 514.950 692.400 547.050 693.600 ;
        RECT 514.950 691.950 517.050 692.400 ;
        RECT 544.950 691.950 547.050 692.400 ;
        RECT 574.950 693.600 577.050 694.050 ;
        RECT 583.950 693.600 586.050 694.050 ;
        RECT 574.950 692.400 586.050 693.600 ;
        RECT 574.950 691.950 577.050 692.400 ;
        RECT 583.950 691.950 586.050 692.400 ;
        RECT 607.950 693.600 610.050 694.050 ;
        RECT 631.950 693.600 634.050 694.050 ;
        RECT 607.950 692.400 634.050 693.600 ;
        RECT 607.950 691.950 610.050 692.400 ;
        RECT 631.950 691.950 634.050 692.400 ;
        RECT 724.950 693.600 727.050 694.050 ;
        RECT 745.950 693.600 748.050 694.050 ;
        RECT 724.950 692.400 748.050 693.600 ;
        RECT 724.950 691.950 727.050 692.400 ;
        RECT 745.950 691.950 748.050 692.400 ;
        RECT 775.950 693.600 778.050 694.050 ;
        RECT 835.950 693.600 838.050 694.050 ;
        RECT 775.950 692.400 838.050 693.600 ;
        RECT 775.950 691.950 778.050 692.400 ;
        RECT 835.950 691.950 838.050 692.400 ;
        RECT 88.950 690.600 91.050 691.050 ;
        RECT 103.950 690.600 106.050 691.050 ;
        RECT 88.950 689.400 106.050 690.600 ;
        RECT 88.950 688.950 91.050 689.400 ;
        RECT 103.950 688.950 106.050 689.400 ;
        RECT 202.950 690.600 205.050 691.050 ;
        RECT 229.950 690.600 232.050 691.050 ;
        RECT 376.950 690.600 379.050 691.050 ;
        RECT 382.950 690.600 385.050 691.050 ;
        RECT 415.950 690.600 418.050 691.050 ;
        RECT 595.950 690.600 598.050 691.050 ;
        RECT 202.950 689.400 321.600 690.600 ;
        RECT 202.950 688.950 205.050 689.400 ;
        RECT 229.950 688.950 232.050 689.400 ;
        RECT 43.950 685.950 46.050 688.050 ;
        RECT 52.950 687.600 55.050 688.050 ;
        RECT 61.950 687.600 64.050 688.050 ;
        RECT 52.950 686.400 64.050 687.600 ;
        RECT 320.400 687.600 321.600 689.400 ;
        RECT 376.950 689.400 418.050 690.600 ;
        RECT 376.950 688.950 379.050 689.400 ;
        RECT 382.950 688.950 385.050 689.400 ;
        RECT 415.950 688.950 418.050 689.400 ;
        RECT 491.400 689.400 598.050 690.600 ;
        RECT 491.400 688.050 492.600 689.400 ;
        RECT 595.950 688.950 598.050 689.400 ;
        RECT 646.950 690.600 649.050 691.050 ;
        RECT 652.950 690.600 655.050 691.050 ;
        RECT 646.950 689.400 655.050 690.600 ;
        RECT 646.950 688.950 649.050 689.400 ;
        RECT 652.950 688.950 655.050 689.400 ;
        RECT 664.950 690.600 667.050 691.050 ;
        RECT 748.950 690.600 751.050 691.050 ;
        RECT 664.950 689.400 751.050 690.600 ;
        RECT 664.950 688.950 667.050 689.400 ;
        RECT 748.950 688.950 751.050 689.400 ;
        RECT 328.950 687.600 331.050 688.050 ;
        RECT 320.400 686.400 331.050 687.600 ;
        RECT 52.950 685.950 55.050 686.400 ;
        RECT 61.950 685.950 64.050 686.400 ;
        RECT 328.950 685.950 331.050 686.400 ;
        RECT 367.950 687.600 370.050 688.050 ;
        RECT 373.950 687.600 376.050 688.050 ;
        RECT 367.950 686.400 376.050 687.600 ;
        RECT 367.950 685.950 370.050 686.400 ;
        RECT 373.950 685.950 376.050 686.400 ;
        RECT 457.950 687.600 460.050 688.050 ;
        RECT 481.950 687.600 484.050 688.050 ;
        RECT 490.950 687.600 493.050 688.050 ;
        RECT 457.950 686.400 493.050 687.600 ;
        RECT 457.950 685.950 460.050 686.400 ;
        RECT 481.950 685.950 484.050 686.400 ;
        RECT 490.950 685.950 493.050 686.400 ;
        RECT 721.950 685.950 724.050 688.050 ;
        RECT 787.950 687.600 790.050 688.050 ;
        RECT 802.950 687.600 805.050 688.050 ;
        RECT 787.950 686.400 805.050 687.600 ;
        RECT 787.950 685.950 790.050 686.400 ;
        RECT 802.950 685.950 805.050 686.400 ;
        RECT 841.950 687.600 844.050 688.050 ;
        RECT 859.950 687.600 862.050 688.050 ;
        RECT 841.950 686.400 862.050 687.600 ;
        RECT 841.950 685.950 844.050 686.400 ;
        RECT 859.950 685.950 862.050 686.400 ;
        RECT 28.950 684.750 31.050 685.200 ;
        RECT 37.950 684.750 40.050 685.200 ;
        RECT 28.950 683.550 40.050 684.750 ;
        RECT 28.950 683.100 31.050 683.550 ;
        RECT 37.950 683.100 40.050 683.550 ;
        RECT 22.950 678.600 25.050 678.900 ;
        RECT 28.950 678.600 31.050 679.050 ;
        RECT 22.950 677.400 31.050 678.600 ;
        RECT 22.950 676.800 25.050 677.400 ;
        RECT 28.950 676.950 31.050 677.400 ;
        RECT 44.400 676.050 45.600 685.950 ;
        RECT 58.950 682.950 61.050 685.050 ;
        RECT 73.950 684.600 76.050 685.050 ;
        RECT 88.950 684.600 91.050 685.200 ;
        RECT 73.950 683.400 91.050 684.600 ;
        RECT 73.950 682.950 76.050 683.400 ;
        RECT 88.950 683.100 91.050 683.400 ;
        RECT 97.950 684.600 100.050 685.200 ;
        RECT 109.950 684.600 112.050 685.200 ;
        RECT 115.950 684.600 118.050 685.200 ;
        RECT 124.950 684.750 127.050 685.200 ;
        RECT 130.950 684.750 133.050 685.200 ;
        RECT 124.950 684.600 133.050 684.750 ;
        RECT 97.950 683.400 114.600 684.600 ;
        RECT 97.950 683.100 100.050 683.400 ;
        RECT 109.950 683.100 112.050 683.400 ;
        RECT 59.400 679.050 60.600 682.950 ;
        RECT 113.400 681.600 114.600 683.400 ;
        RECT 115.950 683.550 133.050 684.600 ;
        RECT 115.950 683.400 127.050 683.550 ;
        RECT 115.950 683.100 118.050 683.400 ;
        RECT 124.950 683.100 127.050 683.400 ;
        RECT 130.950 683.100 133.050 683.550 ;
        RECT 136.950 684.750 139.050 685.200 ;
        RECT 157.950 684.750 160.050 685.050 ;
        RECT 166.950 684.750 169.050 685.200 ;
        RECT 136.950 683.550 169.050 684.750 ;
        RECT 136.950 683.100 139.050 683.550 ;
        RECT 157.950 682.950 160.050 683.550 ;
        RECT 166.950 683.100 169.050 683.550 ;
        RECT 175.950 684.600 178.050 685.200 ;
        RECT 187.950 684.600 190.050 685.050 ;
        RECT 214.950 684.600 217.050 685.200 ;
        RECT 175.950 683.400 217.050 684.600 ;
        RECT 175.950 683.100 178.050 683.400 ;
        RECT 187.950 682.950 190.050 683.400 ;
        RECT 214.950 683.100 217.050 683.400 ;
        RECT 220.950 683.100 223.050 685.200 ;
        RECT 241.950 684.750 244.050 685.200 ;
        RECT 256.950 684.750 259.050 685.200 ;
        RECT 241.950 683.550 259.050 684.750 ;
        RECT 241.950 683.100 244.050 683.550 ;
        RECT 256.950 683.100 259.050 683.550 ;
        RECT 113.400 681.000 120.600 681.600 ;
        RECT 113.400 680.400 121.050 681.000 ;
        RECT 58.950 676.950 61.050 679.050 ;
        RECT 67.950 678.600 70.050 679.050 ;
        RECT 79.950 678.600 82.050 679.050 ;
        RECT 67.950 677.400 82.050 678.600 ;
        RECT 67.950 676.950 70.050 677.400 ;
        RECT 79.950 676.950 82.050 677.400 ;
        RECT 118.950 676.950 121.050 680.400 ;
        RECT 133.950 678.600 136.050 678.900 ;
        RECT 148.950 678.600 151.050 679.050 ;
        RECT 133.950 677.400 151.050 678.600 ;
        RECT 133.950 676.800 136.050 677.400 ;
        RECT 148.950 676.950 151.050 677.400 ;
        RECT 166.950 678.600 169.050 679.050 ;
        RECT 211.950 678.600 214.050 679.050 ;
        RECT 166.950 677.400 214.050 678.600 ;
        RECT 166.950 676.950 169.050 677.400 ;
        RECT 211.950 676.950 214.050 677.400 ;
        RECT 221.400 676.050 222.600 683.100 ;
        RECT 262.950 682.950 265.050 685.050 ;
        RECT 274.950 684.750 277.050 685.200 ;
        RECT 283.950 684.750 286.050 685.200 ;
        RECT 274.950 683.550 286.050 684.750 ;
        RECT 274.950 683.100 277.050 683.550 ;
        RECT 283.950 683.100 286.050 683.550 ;
        RECT 295.950 684.750 298.050 685.200 ;
        RECT 301.950 684.750 304.050 685.200 ;
        RECT 295.950 683.550 304.050 684.750 ;
        RECT 295.950 683.100 298.050 683.550 ;
        RECT 301.950 683.100 304.050 683.550 ;
        RECT 316.950 683.100 319.050 685.200 ;
        RECT 340.950 684.600 343.050 685.200 ;
        RECT 349.950 684.600 352.050 685.050 ;
        RECT 355.950 684.600 358.050 685.200 ;
        RECT 340.950 683.400 358.050 684.600 ;
        RECT 340.950 683.100 343.050 683.400 ;
        RECT 223.950 678.600 226.050 678.900 ;
        RECT 235.950 678.600 238.050 679.050 ;
        RECT 223.950 677.400 238.050 678.600 ;
        RECT 223.950 676.800 226.050 677.400 ;
        RECT 235.950 676.950 238.050 677.400 ;
        RECT 244.950 678.600 247.050 678.900 ;
        RECT 263.400 678.600 264.600 682.950 ;
        RECT 317.400 681.600 318.600 683.100 ;
        RECT 349.950 682.950 352.050 683.400 ;
        RECT 355.950 683.100 358.050 683.400 ;
        RECT 403.950 683.100 406.050 685.200 ;
        RECT 409.950 683.100 412.050 685.200 ;
        RECT 415.950 684.600 418.050 685.050 ;
        RECT 439.950 684.750 442.050 685.200 ;
        RECT 445.950 684.750 448.050 685.200 ;
        RECT 415.950 683.400 432.600 684.600 ;
        RECT 346.950 681.600 349.050 682.050 ;
        RECT 404.400 681.600 405.600 683.100 ;
        RECT 317.400 680.400 349.050 681.600 ;
        RECT 346.950 679.950 349.050 680.400 ;
        RECT 395.400 680.400 405.600 681.600 ;
        RECT 244.950 677.400 264.600 678.600 ;
        RECT 271.950 678.450 274.050 678.900 ;
        RECT 280.950 678.450 283.050 678.900 ;
        RECT 244.950 676.800 247.050 677.400 ;
        RECT 271.950 677.250 283.050 678.450 ;
        RECT 271.950 676.800 274.050 677.250 ;
        RECT 280.950 676.800 283.050 677.250 ;
        RECT 304.950 678.600 307.050 679.050 ;
        RECT 313.950 678.600 316.050 678.900 ;
        RECT 304.950 677.400 316.050 678.600 ;
        RECT 304.950 676.950 307.050 677.400 ;
        RECT 313.950 676.800 316.050 677.400 ;
        RECT 334.950 678.600 337.050 678.900 ;
        RECT 358.950 678.600 361.050 678.900 ;
        RECT 334.950 678.450 361.050 678.600 ;
        RECT 376.950 678.450 379.050 678.900 ;
        RECT 334.950 677.400 379.050 678.450 ;
        RECT 334.950 676.800 337.050 677.400 ;
        RECT 358.950 677.250 379.050 677.400 ;
        RECT 358.950 676.800 361.050 677.250 ;
        RECT 376.950 676.800 379.050 677.250 ;
        RECT 385.950 678.600 388.050 678.900 ;
        RECT 395.400 678.600 396.600 680.400 ;
        RECT 385.950 677.400 396.600 678.600 ;
        RECT 397.950 678.600 400.050 679.050 ;
        RECT 406.950 678.600 409.050 678.900 ;
        RECT 397.950 677.400 409.050 678.600 ;
        RECT 410.400 678.600 411.600 683.100 ;
        RECT 415.950 682.950 418.050 683.400 ;
        RECT 415.950 678.600 418.050 679.050 ;
        RECT 410.400 677.400 418.050 678.600 ;
        RECT 431.400 678.600 432.600 683.400 ;
        RECT 439.950 683.550 448.050 684.750 ;
        RECT 439.950 683.100 442.050 683.550 ;
        RECT 445.950 683.100 448.050 683.550 ;
        RECT 463.950 683.100 466.050 685.200 ;
        RECT 487.950 684.600 490.050 685.200 ;
        RECT 499.950 684.600 502.050 685.050 ;
        RECT 505.950 684.600 508.050 685.200 ;
        RECT 510.000 684.600 514.050 685.050 ;
        RECT 487.950 683.400 508.050 684.600 ;
        RECT 487.950 683.100 490.050 683.400 ;
        RECT 436.950 678.600 439.050 678.900 ;
        RECT 431.400 677.400 439.050 678.600 ;
        RECT 385.950 676.800 388.050 677.400 ;
        RECT 397.950 676.950 400.050 677.400 ;
        RECT 406.950 676.800 409.050 677.400 ;
        RECT 415.950 676.950 418.050 677.400 ;
        RECT 436.950 676.800 439.050 677.400 ;
        RECT 448.950 678.600 451.050 679.050 ;
        RECT 460.950 678.600 463.050 678.900 ;
        RECT 448.950 677.400 463.050 678.600 ;
        RECT 448.950 676.950 451.050 677.400 ;
        RECT 460.950 676.800 463.050 677.400 ;
        RECT 43.950 673.950 46.050 676.050 ;
        RECT 94.950 675.600 97.050 676.050 ;
        RECT 124.950 675.600 127.050 676.050 ;
        RECT 94.950 674.400 127.050 675.600 ;
        RECT 94.950 673.950 97.050 674.400 ;
        RECT 124.950 673.950 127.050 674.400 ;
        RECT 187.950 675.600 190.050 676.050 ;
        RECT 199.950 675.600 202.050 676.050 ;
        RECT 187.950 674.400 202.050 675.600 ;
        RECT 187.950 673.950 190.050 674.400 ;
        RECT 199.950 673.950 202.050 674.400 ;
        RECT 220.950 673.950 223.050 676.050 ;
        RECT 259.950 675.600 262.050 676.050 ;
        RECT 265.950 675.600 268.050 676.050 ;
        RECT 259.950 674.400 268.050 675.600 ;
        RECT 259.950 673.950 262.050 674.400 ;
        RECT 265.950 673.950 268.050 674.400 ;
        RECT 289.950 675.600 292.050 676.050 ;
        RECT 301.950 675.600 304.050 676.050 ;
        RECT 289.950 674.400 304.050 675.600 ;
        RECT 289.950 673.950 292.050 674.400 ;
        RECT 301.950 673.950 304.050 674.400 ;
        RECT 418.950 675.600 421.050 676.050 ;
        RECT 427.950 675.600 430.050 676.050 ;
        RECT 418.950 674.400 430.050 675.600 ;
        RECT 418.950 673.950 421.050 674.400 ;
        RECT 427.950 673.950 430.050 674.400 ;
        RECT 439.950 675.600 442.050 676.050 ;
        RECT 454.950 675.600 457.050 676.050 ;
        RECT 439.950 674.400 457.050 675.600 ;
        RECT 464.400 675.600 465.600 683.100 ;
        RECT 499.950 682.950 502.050 683.400 ;
        RECT 505.950 683.100 508.050 683.400 ;
        RECT 509.400 682.950 514.050 684.600 ;
        RECT 529.950 683.100 532.050 685.200 ;
        RECT 544.950 684.750 547.050 685.200 ;
        RECT 550.950 684.750 553.050 685.200 ;
        RECT 544.950 683.550 553.050 684.750 ;
        RECT 544.950 683.100 547.050 683.550 ;
        RECT 550.950 683.100 553.050 683.550 ;
        RECT 562.950 684.750 565.050 685.200 ;
        RECT 574.950 684.750 577.050 685.200 ;
        RECT 562.950 683.550 577.050 684.750 ;
        RECT 562.950 683.100 565.050 683.550 ;
        RECT 574.950 683.100 577.050 683.550 ;
        RECT 580.950 683.100 583.050 685.200 ;
        RECT 604.950 684.600 607.050 685.200 ;
        RECT 622.950 684.600 625.050 685.200 ;
        RECT 604.950 683.400 625.050 684.600 ;
        RECT 604.950 683.100 607.050 683.400 ;
        RECT 622.950 683.100 625.050 683.400 ;
        RECT 640.950 684.600 645.000 685.050 ;
        RECT 484.950 678.600 487.050 678.900 ;
        RECT 493.950 678.600 496.050 679.050 ;
        RECT 484.950 677.400 496.050 678.600 ;
        RECT 484.950 676.800 487.050 677.400 ;
        RECT 493.950 676.950 496.050 677.400 ;
        RECT 509.400 676.050 510.600 682.950 ;
        RECT 530.400 676.050 531.600 683.100 ;
        RECT 532.950 678.450 535.050 678.900 ;
        RECT 541.950 678.450 544.050 678.900 ;
        RECT 532.950 677.250 544.050 678.450 ;
        RECT 532.950 676.800 535.050 677.250 ;
        RECT 541.950 676.800 544.050 677.250 ;
        RECT 553.950 678.600 556.050 678.900 ;
        RECT 581.400 678.600 582.600 683.100 ;
        RECT 640.950 682.950 645.600 684.600 ;
        RECT 652.950 682.950 655.050 685.050 ;
        RECT 667.950 684.750 670.050 685.200 ;
        RECT 673.950 684.750 676.050 685.200 ;
        RECT 667.950 683.550 676.050 684.750 ;
        RECT 667.950 683.100 670.050 683.550 ;
        RECT 673.950 683.100 676.050 683.550 ;
        RECT 697.950 683.100 700.050 685.200 ;
        RECT 703.950 683.100 706.050 685.200 ;
        RECT 644.400 681.600 645.600 682.950 ;
        RECT 635.400 681.000 645.600 681.600 ;
        RECT 634.950 680.400 645.600 681.000 ;
        RECT 553.950 677.400 582.600 678.600 ;
        RECT 601.950 678.600 604.050 678.900 ;
        RECT 616.950 678.600 619.050 679.050 ;
        RECT 601.950 677.400 619.050 678.600 ;
        RECT 553.950 676.800 556.050 677.400 ;
        RECT 601.950 676.800 604.050 677.400 ;
        RECT 616.950 676.950 619.050 677.400 ;
        RECT 634.950 676.950 637.050 680.400 ;
        RECT 644.400 678.900 645.600 680.400 ;
        RECT 653.400 679.050 654.600 682.950 ;
        RECT 643.950 676.800 646.050 678.900 ;
        RECT 652.950 676.950 655.050 679.050 ;
        RECT 664.950 678.450 667.050 678.900 ;
        RECT 670.950 678.450 673.050 678.900 ;
        RECT 664.950 677.250 673.050 678.450 ;
        RECT 664.950 676.800 667.050 677.250 ;
        RECT 670.950 676.800 673.050 677.250 ;
        RECT 676.950 678.450 679.050 678.900 ;
        RECT 685.950 678.450 688.050 678.900 ;
        RECT 676.950 677.250 688.050 678.450 ;
        RECT 676.950 676.800 679.050 677.250 ;
        RECT 685.950 676.800 688.050 677.250 ;
        RECT 691.950 678.600 694.050 679.050 ;
        RECT 698.400 678.600 699.600 683.100 ;
        RECT 691.950 677.400 699.600 678.600 ;
        RECT 704.400 679.050 705.600 683.100 ;
        RECT 704.400 677.400 709.050 679.050 ;
        RECT 722.400 678.900 723.600 685.950 ;
        RECT 724.950 684.600 727.050 685.200 ;
        RECT 733.950 684.750 736.050 685.200 ;
        RECT 742.950 684.750 745.050 685.200 ;
        RECT 733.950 684.600 745.050 684.750 ;
        RECT 724.950 683.550 745.050 684.600 ;
        RECT 724.950 683.400 736.050 683.550 ;
        RECT 724.950 683.100 727.050 683.400 ;
        RECT 733.950 683.100 736.050 683.400 ;
        RECT 742.950 683.100 745.050 683.550 ;
        RECT 748.950 684.600 751.050 685.200 ;
        RECT 769.950 684.600 772.050 685.200 ;
        RECT 748.950 683.400 772.050 684.600 ;
        RECT 748.950 683.100 751.050 683.400 ;
        RECT 769.950 683.100 772.050 683.400 ;
        RECT 775.950 683.100 778.050 685.200 ;
        RECT 814.950 683.100 817.050 685.200 ;
        RECT 820.950 684.750 823.050 685.200 ;
        RECT 826.950 684.750 829.050 685.200 ;
        RECT 820.950 683.550 829.050 684.750 ;
        RECT 820.950 683.100 823.050 683.550 ;
        RECT 826.950 683.100 829.050 683.550 ;
        RECT 691.950 676.950 694.050 677.400 ;
        RECT 705.000 676.950 709.050 677.400 ;
        RECT 721.950 676.800 724.050 678.900 ;
        RECT 727.950 678.600 730.050 678.900 ;
        RECT 739.950 678.600 742.050 678.900 ;
        RECT 727.950 677.400 742.050 678.600 ;
        RECT 727.950 676.800 730.050 677.400 ;
        RECT 739.950 676.800 742.050 677.400 ;
        RECT 745.950 678.600 748.050 678.900 ;
        RECT 757.950 678.600 760.050 679.050 ;
        RECT 745.950 677.400 760.050 678.600 ;
        RECT 776.400 678.600 777.600 683.100 ;
        RECT 790.950 678.600 793.050 678.900 ;
        RECT 776.400 677.400 793.050 678.600 ;
        RECT 815.400 678.600 816.600 683.100 ;
        RECT 850.950 682.950 853.050 685.050 ;
        RECT 865.950 684.750 868.050 685.200 ;
        RECT 874.950 684.750 877.050 685.200 ;
        RECT 865.950 683.550 877.050 684.750 ;
        RECT 865.950 683.100 868.050 683.550 ;
        RECT 874.950 683.100 877.050 683.550 ;
        RECT 851.400 679.050 852.600 682.950 ;
        RECT 880.950 681.600 883.050 685.050 ;
        RECT 880.950 681.000 885.600 681.600 ;
        RECT 881.400 680.400 885.600 681.000 ;
        RECT 838.950 678.600 841.050 678.900 ;
        RECT 815.400 677.400 841.050 678.600 ;
        RECT 745.950 676.800 748.050 677.400 ;
        RECT 757.950 676.950 760.050 677.400 ;
        RECT 790.950 676.800 793.050 677.400 ;
        RECT 838.950 676.800 841.050 677.400 ;
        RECT 850.950 676.950 853.050 679.050 ;
        RECT 884.400 678.600 885.600 680.400 ;
        RECT 892.950 678.600 895.050 679.050 ;
        RECT 884.400 677.400 895.050 678.600 ;
        RECT 892.950 676.950 895.050 677.400 ;
        RECT 469.800 675.600 471.900 675.900 ;
        RECT 464.400 674.400 471.900 675.600 ;
        RECT 439.950 673.950 442.050 674.400 ;
        RECT 454.950 673.950 457.050 674.400 ;
        RECT 469.800 673.800 471.900 674.400 ;
        RECT 472.950 675.600 475.050 676.050 ;
        RECT 478.950 675.600 481.050 676.050 ;
        RECT 472.950 674.400 481.050 675.600 ;
        RECT 472.950 673.950 475.050 674.400 ;
        RECT 478.950 673.950 481.050 674.400 ;
        RECT 508.950 673.950 511.050 676.050 ;
        RECT 520.950 675.600 523.050 676.050 ;
        RECT 526.800 675.600 528.900 676.050 ;
        RECT 520.950 674.400 528.900 675.600 ;
        RECT 520.950 673.950 523.050 674.400 ;
        RECT 526.800 673.950 528.900 674.400 ;
        RECT 529.950 673.950 532.050 676.050 ;
        RECT 544.950 675.600 547.050 676.050 ;
        RECT 550.950 675.600 553.050 676.050 ;
        RECT 544.950 674.400 553.050 675.600 ;
        RECT 544.950 673.950 547.050 674.400 ;
        RECT 550.950 673.950 553.050 674.400 ;
        RECT 556.950 675.600 559.050 676.050 ;
        RECT 562.950 675.600 565.050 676.050 ;
        RECT 556.950 674.400 565.050 675.600 ;
        RECT 556.950 673.950 559.050 674.400 ;
        RECT 562.950 673.950 565.050 674.400 ;
        RECT 580.950 675.600 583.050 676.050 ;
        RECT 586.950 675.600 589.050 676.050 ;
        RECT 580.950 674.400 589.050 675.600 ;
        RECT 580.950 673.950 583.050 674.400 ;
        RECT 586.950 673.950 589.050 674.400 ;
        RECT 772.950 675.600 775.050 676.050 ;
        RECT 796.950 675.600 799.050 676.050 ;
        RECT 802.950 675.600 805.050 676.050 ;
        RECT 772.950 674.400 805.050 675.600 ;
        RECT 772.950 673.950 775.050 674.400 ;
        RECT 796.950 673.950 799.050 674.400 ;
        RECT 802.950 673.950 805.050 674.400 ;
        RECT 811.950 675.600 814.050 676.050 ;
        RECT 823.950 675.600 826.050 676.050 ;
        RECT 832.950 675.600 835.050 676.050 ;
        RECT 811.950 674.400 835.050 675.600 ;
        RECT 811.950 673.950 814.050 674.400 ;
        RECT 823.950 673.950 826.050 674.400 ;
        RECT 832.950 673.950 835.050 674.400 ;
        RECT 859.950 675.600 862.050 676.050 ;
        RECT 874.950 675.600 877.050 676.050 ;
        RECT 859.950 674.400 877.050 675.600 ;
        RECT 859.950 673.950 862.050 674.400 ;
        RECT 874.950 673.950 877.050 674.400 ;
        RECT 880.950 675.600 883.050 676.050 ;
        RECT 889.950 675.600 892.050 676.050 ;
        RECT 880.950 674.400 892.050 675.600 ;
        RECT 880.950 673.950 883.050 674.400 ;
        RECT 889.950 673.950 892.050 674.400 ;
        RECT 55.950 672.600 58.050 673.050 ;
        RECT 64.950 672.600 67.050 673.050 ;
        RECT 112.950 672.600 115.050 673.050 ;
        RECT 55.950 671.400 115.050 672.600 ;
        RECT 55.950 670.950 58.050 671.400 ;
        RECT 64.950 670.950 67.050 671.400 ;
        RECT 112.950 670.950 115.050 671.400 ;
        RECT 358.950 672.600 361.050 673.050 ;
        RECT 394.950 672.600 397.050 673.050 ;
        RECT 409.800 672.600 411.900 673.050 ;
        RECT 358.950 671.400 411.900 672.600 ;
        RECT 358.950 670.950 361.050 671.400 ;
        RECT 394.950 670.950 397.050 671.400 ;
        RECT 409.800 670.950 411.900 671.400 ;
        RECT 412.950 672.600 415.050 673.050 ;
        RECT 466.950 672.600 469.050 673.050 ;
        RECT 412.950 671.400 469.050 672.600 ;
        RECT 412.950 670.950 415.050 671.400 ;
        RECT 466.950 670.950 469.050 671.400 ;
        RECT 487.950 672.600 490.050 673.050 ;
        RECT 499.950 672.600 502.050 673.050 ;
        RECT 487.950 671.400 502.050 672.600 ;
        RECT 487.950 670.950 490.050 671.400 ;
        RECT 499.950 670.950 502.050 671.400 ;
        RECT 577.950 672.600 580.050 673.050 ;
        RECT 583.950 672.600 586.050 673.050 ;
        RECT 577.950 671.400 586.050 672.600 ;
        RECT 577.950 670.950 580.050 671.400 ;
        RECT 583.950 670.950 586.050 671.400 ;
        RECT 649.950 672.600 652.050 673.050 ;
        RECT 691.950 672.600 694.050 673.050 ;
        RECT 649.950 671.400 694.050 672.600 ;
        RECT 649.950 670.950 652.050 671.400 ;
        RECT 691.950 670.950 694.050 671.400 ;
        RECT 700.950 670.950 703.050 673.050 ;
        RECT 826.950 672.600 829.050 673.050 ;
        RECT 841.950 672.600 844.050 673.050 ;
        RECT 826.950 671.400 844.050 672.600 ;
        RECT 826.950 670.950 829.050 671.400 ;
        RECT 841.950 670.950 844.050 671.400 ;
        RECT 4.950 669.600 7.050 670.050 ;
        RECT 28.950 669.600 31.050 670.050 ;
        RECT 4.950 668.400 31.050 669.600 ;
        RECT 4.950 667.950 7.050 668.400 ;
        RECT 28.950 667.950 31.050 668.400 ;
        RECT 49.950 669.600 52.050 670.050 ;
        RECT 70.950 669.600 73.050 670.050 ;
        RECT 49.950 668.400 73.050 669.600 ;
        RECT 49.950 667.950 52.050 668.400 ;
        RECT 70.950 667.950 73.050 668.400 ;
        RECT 178.950 669.600 181.050 670.050 ;
        RECT 250.950 669.600 253.050 670.050 ;
        RECT 292.950 669.600 295.050 670.050 ;
        RECT 313.950 669.600 316.050 670.050 ;
        RECT 178.950 668.400 295.050 669.600 ;
        RECT 178.950 667.950 181.050 668.400 ;
        RECT 250.950 667.950 253.050 668.400 ;
        RECT 292.950 667.950 295.050 668.400 ;
        RECT 296.400 668.400 316.050 669.600 ;
        RECT 217.950 666.600 220.050 667.050 ;
        RECT 229.950 666.600 232.050 667.050 ;
        RECT 217.950 665.400 232.050 666.600 ;
        RECT 217.950 664.950 220.050 665.400 ;
        RECT 229.950 664.950 232.050 665.400 ;
        RECT 256.950 666.600 259.050 667.050 ;
        RECT 296.400 666.600 297.600 668.400 ;
        RECT 313.950 667.950 316.050 668.400 ;
        RECT 355.950 669.600 358.050 670.050 ;
        RECT 364.950 669.600 367.050 670.050 ;
        RECT 355.950 668.400 367.050 669.600 ;
        RECT 355.950 667.950 358.050 668.400 ;
        RECT 364.950 667.950 367.050 668.400 ;
        RECT 385.950 669.600 388.050 670.050 ;
        RECT 424.950 669.600 427.050 669.900 ;
        RECT 385.950 668.400 427.050 669.600 ;
        RECT 385.950 667.950 388.050 668.400 ;
        RECT 424.950 667.800 427.050 668.400 ;
        RECT 457.950 669.600 460.050 670.050 ;
        RECT 484.950 669.600 487.050 670.050 ;
        RECT 457.950 668.400 487.050 669.600 ;
        RECT 457.950 667.950 460.050 668.400 ;
        RECT 484.950 667.950 487.050 668.400 ;
        RECT 529.950 669.600 532.050 670.050 ;
        RECT 553.950 669.600 556.050 670.050 ;
        RECT 529.950 668.400 556.050 669.600 ;
        RECT 529.950 667.950 532.050 668.400 ;
        RECT 553.950 667.950 556.050 668.400 ;
        RECT 701.400 667.050 702.600 670.950 ;
        RECT 703.950 669.600 706.050 670.050 ;
        RECT 712.950 669.600 715.050 670.050 ;
        RECT 703.950 668.400 715.050 669.600 ;
        RECT 703.950 667.950 706.050 668.400 ;
        RECT 712.950 667.950 715.050 668.400 ;
        RECT 730.950 669.600 733.050 670.050 ;
        RECT 760.950 669.600 763.050 670.050 ;
        RECT 730.950 668.400 763.050 669.600 ;
        RECT 730.950 667.950 733.050 668.400 ;
        RECT 760.950 667.950 763.050 668.400 ;
        RECT 766.950 669.600 769.050 670.050 ;
        RECT 781.950 669.600 784.050 670.050 ;
        RECT 766.950 668.400 784.050 669.600 ;
        RECT 766.950 667.950 769.050 668.400 ;
        RECT 781.950 667.950 784.050 668.400 ;
        RECT 844.950 669.600 847.050 670.050 ;
        RECT 853.950 669.600 856.050 670.050 ;
        RECT 862.950 669.600 865.050 670.050 ;
        RECT 844.950 668.400 865.050 669.600 ;
        RECT 844.950 667.950 847.050 668.400 ;
        RECT 853.950 667.950 856.050 668.400 ;
        RECT 862.950 667.950 865.050 668.400 ;
        RECT 256.950 665.400 297.600 666.600 ;
        RECT 304.950 666.600 307.050 667.050 ;
        RECT 322.950 666.600 325.050 667.050 ;
        RECT 328.950 666.600 331.050 667.050 ;
        RECT 304.950 665.400 331.050 666.600 ;
        RECT 256.950 664.950 259.050 665.400 ;
        RECT 304.950 664.950 307.050 665.400 ;
        RECT 322.950 664.950 325.050 665.400 ;
        RECT 328.950 664.950 331.050 665.400 ;
        RECT 379.950 666.600 382.050 667.050 ;
        RECT 421.950 666.600 424.050 667.050 ;
        RECT 511.950 666.600 514.050 667.050 ;
        RECT 589.950 666.600 592.050 667.050 ;
        RECT 379.950 665.400 592.050 666.600 ;
        RECT 701.400 666.900 705.000 667.050 ;
        RECT 701.400 665.400 706.050 666.900 ;
        RECT 379.950 664.950 382.050 665.400 ;
        RECT 421.950 664.950 424.050 665.400 ;
        RECT 511.950 664.950 514.050 665.400 ;
        RECT 589.950 664.950 592.050 665.400 ;
        RECT 702.000 664.950 706.050 665.400 ;
        RECT 772.950 666.600 775.050 667.050 ;
        RECT 790.950 666.600 793.050 667.050 ;
        RECT 772.950 665.400 793.050 666.600 ;
        RECT 772.950 664.950 775.050 665.400 ;
        RECT 790.950 664.950 793.050 665.400 ;
        RECT 805.950 666.600 808.050 667.050 ;
        RECT 829.950 666.600 832.050 667.050 ;
        RECT 805.950 665.400 832.050 666.600 ;
        RECT 805.950 664.950 808.050 665.400 ;
        RECT 829.950 664.950 832.050 665.400 ;
        RECT 841.950 666.600 844.050 667.050 ;
        RECT 868.950 666.600 871.050 667.050 ;
        RECT 877.950 666.600 880.050 667.050 ;
        RECT 841.950 665.400 880.050 666.600 ;
        RECT 841.950 664.950 844.050 665.400 ;
        RECT 868.950 664.950 871.050 665.400 ;
        RECT 877.950 664.950 880.050 665.400 ;
        RECT 4.950 663.600 7.050 664.050 ;
        RECT 55.950 663.600 58.050 664.050 ;
        RECT 4.950 662.400 58.050 663.600 ;
        RECT 4.950 661.950 7.050 662.400 ;
        RECT 55.950 661.950 58.050 662.400 ;
        RECT 160.950 663.600 163.050 664.050 ;
        RECT 190.950 663.600 193.050 664.050 ;
        RECT 160.950 662.400 193.050 663.600 ;
        RECT 160.950 661.950 163.050 662.400 ;
        RECT 190.950 661.950 193.050 662.400 ;
        RECT 205.950 663.600 208.050 664.050 ;
        RECT 257.400 663.600 258.600 664.950 ;
        RECT 703.950 664.800 706.050 664.950 ;
        RECT 205.950 662.400 258.600 663.600 ;
        RECT 325.950 663.600 328.050 664.050 ;
        RECT 454.950 663.600 457.050 664.050 ;
        RECT 463.950 663.600 466.050 664.050 ;
        RECT 325.950 662.400 378.600 663.600 ;
        RECT 205.950 661.950 208.050 662.400 ;
        RECT 325.950 661.950 328.050 662.400 ;
        RECT 106.950 660.600 109.050 661.050 ;
        RECT 115.950 660.600 118.050 661.050 ;
        RECT 106.950 659.400 118.050 660.600 ;
        RECT 106.950 658.950 109.050 659.400 ;
        RECT 115.950 658.950 118.050 659.400 ;
        RECT 214.950 660.600 217.050 661.050 ;
        RECT 274.950 660.600 277.050 661.050 ;
        RECT 214.950 659.400 277.050 660.600 ;
        RECT 214.950 658.950 217.050 659.400 ;
        RECT 274.950 658.950 277.050 659.400 ;
        RECT 280.950 660.600 283.050 661.050 ;
        RECT 307.950 660.600 310.050 661.050 ;
        RECT 280.950 659.400 310.050 660.600 ;
        RECT 280.950 658.950 283.050 659.400 ;
        RECT 307.950 658.950 310.050 659.400 ;
        RECT 313.950 660.600 316.050 661.050 ;
        RECT 340.950 660.600 343.050 661.050 ;
        RECT 313.950 659.400 343.050 660.600 ;
        RECT 377.400 660.600 378.600 662.400 ;
        RECT 454.950 662.400 466.050 663.600 ;
        RECT 454.950 661.950 457.050 662.400 ;
        RECT 463.950 661.950 466.050 662.400 ;
        RECT 469.950 663.600 472.050 664.050 ;
        RECT 520.950 663.600 523.050 664.050 ;
        RECT 571.950 663.600 574.050 664.050 ;
        RECT 469.950 662.400 523.050 663.600 ;
        RECT 469.950 661.950 472.050 662.400 ;
        RECT 520.950 661.950 523.050 662.400 ;
        RECT 548.400 662.400 574.050 663.600 ;
        RECT 385.950 660.600 388.050 661.050 ;
        RECT 377.400 659.400 388.050 660.600 ;
        RECT 313.950 658.950 316.050 659.400 ;
        RECT 340.950 658.950 343.050 659.400 ;
        RECT 385.950 658.950 388.050 659.400 ;
        RECT 400.950 660.600 403.050 661.050 ;
        RECT 523.950 660.600 526.050 661.050 ;
        RECT 548.400 660.600 549.600 662.400 ;
        RECT 571.950 661.950 574.050 662.400 ;
        RECT 622.950 663.600 625.050 664.050 ;
        RECT 682.800 663.600 684.900 664.050 ;
        RECT 622.950 662.400 684.900 663.600 ;
        RECT 622.950 661.950 625.050 662.400 ;
        RECT 682.800 661.950 684.900 662.400 ;
        RECT 685.950 663.600 688.050 664.050 ;
        RECT 832.950 663.600 835.050 664.050 ;
        RECT 685.950 662.400 835.050 663.600 ;
        RECT 685.950 661.950 688.050 662.400 ;
        RECT 832.950 661.950 835.050 662.400 ;
        RECT 856.950 663.600 859.050 664.050 ;
        RECT 883.950 663.600 886.050 664.050 ;
        RECT 856.950 662.400 886.050 663.600 ;
        RECT 856.950 661.950 859.050 662.400 ;
        RECT 883.950 661.950 886.050 662.400 ;
        RECT 400.950 659.400 549.600 660.600 ;
        RECT 553.950 660.600 556.050 661.050 ;
        RECT 565.950 660.600 568.050 661.050 ;
        RECT 553.950 659.400 568.050 660.600 ;
        RECT 400.950 658.950 403.050 659.400 ;
        RECT 523.950 658.950 526.050 659.400 ;
        RECT 553.950 658.950 556.050 659.400 ;
        RECT 565.950 658.950 568.050 659.400 ;
        RECT 652.950 660.600 655.050 661.050 ;
        RECT 676.950 660.600 679.050 661.050 ;
        RECT 652.950 659.400 679.050 660.600 ;
        RECT 652.950 658.950 655.050 659.400 ;
        RECT 676.950 658.950 679.050 659.400 ;
        RECT 691.950 660.600 694.050 661.050 ;
        RECT 709.950 660.600 712.050 661.050 ;
        RECT 691.950 659.400 712.050 660.600 ;
        RECT 691.950 658.950 694.050 659.400 ;
        RECT 709.950 658.950 712.050 659.400 ;
        RECT 760.950 660.600 763.050 661.050 ;
        RECT 811.950 660.600 814.050 661.050 ;
        RECT 760.950 659.400 814.050 660.600 ;
        RECT 760.950 658.950 763.050 659.400 ;
        RECT 811.950 658.950 814.050 659.400 ;
        RECT 16.950 657.600 19.050 658.050 ;
        RECT 25.950 657.600 28.050 658.050 ;
        RECT 16.950 656.400 28.050 657.600 ;
        RECT 16.950 655.950 19.050 656.400 ;
        RECT 25.950 655.950 28.050 656.400 ;
        RECT 31.950 657.600 34.050 658.050 ;
        RECT 52.950 657.600 55.050 658.050 ;
        RECT 31.950 656.400 55.050 657.600 ;
        RECT 31.950 655.950 34.050 656.400 ;
        RECT 52.950 655.950 55.050 656.400 ;
        RECT 58.950 657.600 61.050 658.050 ;
        RECT 145.950 657.600 148.050 658.050 ;
        RECT 181.950 657.600 184.050 658.050 ;
        RECT 58.950 657.000 78.600 657.600 ;
        RECT 58.950 656.400 79.050 657.000 ;
        RECT 58.950 655.950 61.050 656.400 ;
        RECT 53.400 654.600 54.600 655.950 ;
        RECT 53.400 653.400 75.600 654.600 ;
        RECT 19.950 651.600 22.050 652.200 ;
        RECT 22.950 651.600 25.050 652.050 ;
        RECT 49.950 651.600 52.050 652.200 ;
        RECT 19.950 650.400 52.050 651.600 ;
        RECT 74.400 651.600 75.600 653.400 ;
        RECT 76.950 652.800 79.050 656.400 ;
        RECT 145.950 656.400 184.050 657.600 ;
        RECT 145.950 655.950 148.050 656.400 ;
        RECT 181.950 655.950 184.050 656.400 ;
        RECT 220.950 657.600 223.050 658.050 ;
        RECT 310.950 657.600 313.050 658.050 ;
        RECT 220.950 656.400 313.050 657.600 ;
        RECT 220.950 655.950 223.050 656.400 ;
        RECT 310.950 655.950 313.050 656.400 ;
        RECT 319.950 657.600 322.050 658.050 ;
        RECT 388.950 657.600 391.050 658.050 ;
        RECT 319.950 656.400 391.050 657.600 ;
        RECT 319.950 655.950 322.050 656.400 ;
        RECT 388.950 655.950 391.050 656.400 ;
        RECT 445.950 657.600 448.050 658.050 ;
        RECT 505.950 657.600 508.050 658.050 ;
        RECT 445.950 656.400 508.050 657.600 ;
        RECT 445.950 655.950 448.050 656.400 ;
        RECT 505.950 655.950 508.050 656.400 ;
        RECT 763.950 657.600 766.050 658.050 ;
        RECT 781.950 657.600 784.050 658.050 ;
        RECT 763.950 656.400 784.050 657.600 ;
        RECT 763.950 655.950 766.050 656.400 ;
        RECT 781.950 655.950 784.050 656.400 ;
        RECT 832.950 657.600 835.050 658.050 ;
        RECT 856.950 657.600 859.050 658.050 ;
        RECT 832.950 656.400 859.050 657.600 ;
        RECT 832.950 655.950 835.050 656.400 ;
        RECT 856.950 655.950 859.050 656.400 ;
        RECT 103.950 654.600 106.050 655.050 ;
        RECT 112.950 654.600 115.050 655.050 ;
        RECT 103.950 653.400 115.050 654.600 ;
        RECT 103.950 652.950 106.050 653.400 ;
        RECT 112.950 652.950 115.050 653.400 ;
        RECT 127.950 654.600 130.050 655.050 ;
        RECT 133.950 654.600 136.050 655.050 ;
        RECT 127.950 653.400 136.050 654.600 ;
        RECT 127.950 652.950 130.050 653.400 ;
        RECT 133.950 652.950 136.050 653.400 ;
        RECT 238.950 654.600 241.050 655.050 ;
        RECT 250.950 654.600 253.050 655.050 ;
        RECT 268.950 654.600 271.050 655.050 ;
        RECT 238.950 653.400 271.050 654.600 ;
        RECT 238.950 652.950 241.050 653.400 ;
        RECT 250.950 652.950 253.050 653.400 ;
        RECT 268.950 652.950 271.050 653.400 ;
        RECT 286.950 654.600 289.050 655.050 ;
        RECT 298.950 654.600 301.050 655.050 ;
        RECT 286.950 653.400 301.050 654.600 ;
        RECT 286.950 652.950 289.050 653.400 ;
        RECT 298.950 652.950 301.050 653.400 ;
        RECT 367.950 654.600 370.050 655.050 ;
        RECT 421.950 654.600 424.050 655.050 ;
        RECT 367.950 653.400 424.050 654.600 ;
        RECT 367.950 652.950 370.050 653.400 ;
        RECT 421.950 652.950 424.050 653.400 ;
        RECT 433.950 654.600 436.050 655.050 ;
        RECT 457.800 654.600 459.900 655.050 ;
        RECT 433.950 653.400 459.900 654.600 ;
        RECT 433.950 652.950 436.050 653.400 ;
        RECT 457.800 652.950 459.900 653.400 ;
        RECT 460.950 654.600 463.050 655.050 ;
        RECT 496.950 654.600 499.050 655.050 ;
        RECT 547.950 654.600 550.050 655.050 ;
        RECT 559.950 654.600 562.050 655.050 ;
        RECT 460.950 653.400 562.050 654.600 ;
        RECT 460.950 652.950 463.050 653.400 ;
        RECT 496.950 652.950 499.050 653.400 ;
        RECT 547.950 652.950 550.050 653.400 ;
        RECT 559.950 652.950 562.050 653.400 ;
        RECT 571.950 654.600 574.050 655.050 ;
        RECT 616.950 654.600 619.050 655.050 ;
        RECT 571.950 653.400 619.050 654.600 ;
        RECT 571.950 652.950 574.050 653.400 ;
        RECT 616.950 652.950 619.050 653.400 ;
        RECT 628.950 654.600 631.050 655.050 ;
        RECT 637.950 654.600 640.050 655.050 ;
        RECT 628.950 653.400 640.050 654.600 ;
        RECT 628.950 652.950 631.050 653.400 ;
        RECT 637.950 652.950 640.050 653.400 ;
        RECT 667.950 654.600 670.050 655.050 ;
        RECT 688.950 654.600 691.050 655.050 ;
        RECT 667.950 653.400 691.050 654.600 ;
        RECT 667.950 652.950 670.050 653.400 ;
        RECT 688.950 652.950 691.050 653.400 ;
        RECT 721.950 654.600 724.050 655.050 ;
        RECT 727.950 654.600 730.050 655.050 ;
        RECT 745.950 654.600 748.050 655.050 ;
        RECT 721.950 653.400 748.050 654.600 ;
        RECT 721.950 652.950 724.050 653.400 ;
        RECT 727.950 652.950 730.050 653.400 ;
        RECT 745.950 652.950 748.050 653.400 ;
        RECT 817.950 654.600 820.050 655.050 ;
        RECT 829.950 654.600 832.050 655.050 ;
        RECT 817.950 653.400 832.050 654.600 ;
        RECT 817.950 652.950 820.050 653.400 ;
        RECT 829.950 652.950 832.050 653.400 ;
        RECT 82.950 651.600 85.050 652.050 ;
        RECT 74.400 650.400 85.050 651.600 ;
        RECT 19.950 650.100 22.050 650.400 ;
        RECT 22.950 649.950 25.050 650.400 ;
        RECT 49.950 650.100 52.050 650.400 ;
        RECT 50.400 648.600 51.600 650.100 ;
        RECT 82.950 649.950 85.050 650.400 ;
        RECT 91.950 651.750 94.050 652.200 ;
        RECT 100.950 651.750 103.050 652.200 ;
        RECT 91.950 650.550 103.050 651.750 ;
        RECT 91.950 650.100 94.050 650.550 ;
        RECT 100.950 650.100 103.050 650.550 ;
        RECT 121.950 651.600 124.050 652.050 ;
        RECT 166.950 651.750 169.050 652.200 ;
        RECT 175.950 651.750 178.050 652.200 ;
        RECT 121.950 650.400 159.600 651.600 ;
        RECT 121.950 649.950 124.050 650.400 ;
        RECT 41.400 647.400 51.600 648.600 ;
        RECT 34.950 645.600 37.050 645.900 ;
        RECT 41.400 645.600 42.600 647.400 ;
        RECT 34.950 644.400 42.600 645.600 ;
        RECT 43.950 645.450 46.050 645.900 ;
        RECT 52.950 645.450 55.050 645.900 ;
        RECT 34.950 643.800 37.050 644.400 ;
        RECT 43.950 644.250 55.050 645.450 ;
        RECT 43.950 643.800 46.050 644.250 ;
        RECT 52.950 643.800 55.050 644.250 ;
        RECT 64.950 645.450 67.050 645.900 ;
        RECT 103.950 645.450 106.050 645.900 ;
        RECT 64.950 644.250 106.050 645.450 ;
        RECT 64.950 643.800 67.050 644.250 ;
        RECT 103.950 643.800 106.050 644.250 ;
        RECT 145.950 645.600 148.050 646.050 ;
        RECT 158.400 645.600 159.600 650.400 ;
        RECT 166.950 650.550 178.050 651.750 ;
        RECT 166.950 650.100 169.050 650.550 ;
        RECT 175.950 650.100 178.050 650.550 ;
        RECT 208.950 649.950 211.050 652.050 ;
        RECT 214.950 651.600 217.050 651.900 ;
        RECT 223.950 651.600 226.050 652.200 ;
        RECT 214.950 650.400 226.050 651.600 ;
        RECT 202.950 645.600 205.050 645.900 ;
        RECT 209.400 645.600 210.600 649.950 ;
        RECT 214.950 649.800 217.050 650.400 ;
        RECT 223.950 650.100 226.050 650.400 ;
        RECT 229.950 651.600 232.050 652.200 ;
        RECT 244.950 651.600 247.050 652.200 ;
        RECT 229.950 650.400 247.050 651.600 ;
        RECT 229.950 650.100 232.050 650.400 ;
        RECT 244.950 650.100 247.050 650.400 ;
        RECT 292.950 651.600 297.000 652.050 ;
        RECT 292.950 649.950 297.600 651.600 ;
        RECT 316.950 650.100 319.050 652.200 ;
        RECT 322.950 651.750 325.050 652.200 ;
        RECT 358.950 651.750 361.050 652.200 ;
        RECT 322.950 650.550 361.050 651.750 ;
        RECT 322.950 650.100 325.050 650.550 ;
        RECT 358.950 650.100 361.050 650.550 ;
        RECT 394.950 651.750 397.050 652.200 ;
        RECT 400.950 651.750 403.050 652.200 ;
        RECT 394.950 650.550 403.050 651.750 ;
        RECT 394.950 650.100 397.050 650.550 ;
        RECT 400.950 650.100 403.050 650.550 ;
        RECT 424.950 651.600 429.000 652.050 ;
        RECT 463.950 651.600 466.050 652.050 ;
        RECT 469.950 651.600 472.050 652.050 ;
        RECT 296.400 645.900 297.600 649.950 ;
        RECT 226.950 645.600 229.050 645.900 ;
        RECT 145.950 644.400 154.050 645.600 ;
        RECT 158.400 644.400 163.050 645.600 ;
        RECT 145.950 643.950 148.050 644.400 ;
        RECT 151.950 643.500 154.050 644.400 ;
        RECT 160.950 643.500 163.050 644.400 ;
        RECT 202.950 644.400 229.050 645.600 ;
        RECT 202.950 643.800 205.050 644.400 ;
        RECT 226.950 643.800 229.050 644.400 ;
        RECT 253.950 645.600 256.050 645.900 ;
        RECT 271.950 645.600 274.050 645.900 ;
        RECT 253.950 645.450 274.050 645.600 ;
        RECT 286.950 645.450 289.050 645.900 ;
        RECT 253.950 644.400 289.050 645.450 ;
        RECT 253.950 643.800 256.050 644.400 ;
        RECT 271.950 644.250 289.050 644.400 ;
        RECT 271.950 643.800 274.050 644.250 ;
        RECT 286.950 643.800 289.050 644.250 ;
        RECT 295.950 643.800 298.050 645.900 ;
        RECT 307.950 645.600 310.050 646.050 ;
        RECT 317.400 645.600 318.600 650.100 ;
        RECT 424.950 649.950 429.600 651.600 ;
        RECT 463.950 650.400 472.050 651.600 ;
        RECT 463.950 649.950 466.050 650.400 ;
        RECT 469.950 649.950 472.050 650.400 ;
        RECT 484.950 651.600 487.050 652.050 ;
        RECT 499.950 651.600 502.050 652.200 ;
        RECT 484.950 650.400 502.050 651.600 ;
        RECT 484.950 649.950 487.050 650.400 ;
        RECT 499.950 650.100 502.050 650.400 ;
        RECT 428.400 648.600 429.600 649.950 ;
        RECT 500.400 648.600 501.600 650.100 ;
        RECT 505.950 649.950 508.050 652.050 ;
        RECT 529.950 651.750 532.050 652.200 ;
        RECT 541.950 651.750 544.050 652.200 ;
        RECT 529.950 650.550 544.050 651.750 ;
        RECT 529.950 650.100 532.050 650.550 ;
        RECT 541.950 650.100 544.050 650.550 ;
        RECT 586.950 651.600 589.050 652.200 ;
        RECT 586.950 650.400 591.600 651.600 ;
        RECT 586.950 650.100 589.050 650.400 ;
        RECT 428.400 647.400 453.600 648.600 ;
        RECT 352.950 645.600 355.050 646.050 ;
        RECT 428.400 645.900 429.600 647.400 ;
        RECT 452.400 645.900 453.600 647.400 ;
        RECT 479.400 647.400 501.600 648.600 ;
        RECT 361.950 645.600 364.050 645.900 ;
        RECT 385.950 645.600 388.050 645.900 ;
        RECT 307.950 644.400 318.600 645.600 ;
        RECT 350.400 644.400 388.050 645.600 ;
        RECT 307.950 643.950 310.050 644.400 ;
        RECT 58.950 642.600 61.050 643.050 ;
        RECT 70.950 642.600 73.050 643.050 ;
        RECT 58.950 641.400 73.050 642.600 ;
        RECT 58.950 640.950 61.050 641.400 ;
        RECT 70.950 640.950 73.050 641.400 ;
        RECT 343.950 642.600 346.050 643.050 ;
        RECT 350.400 642.600 351.600 644.400 ;
        RECT 352.950 643.950 355.050 644.400 ;
        RECT 361.950 643.800 364.050 644.400 ;
        RECT 385.950 643.800 388.050 644.400 ;
        RECT 391.950 645.450 394.050 645.900 ;
        RECT 403.950 645.450 406.050 645.900 ;
        RECT 391.950 644.250 406.050 645.450 ;
        RECT 391.950 643.800 394.050 644.250 ;
        RECT 403.950 643.800 406.050 644.250 ;
        RECT 412.950 645.450 415.050 645.900 ;
        RECT 421.950 645.450 424.050 645.900 ;
        RECT 412.950 644.250 424.050 645.450 ;
        RECT 412.950 643.800 415.050 644.250 ;
        RECT 421.950 643.800 424.050 644.250 ;
        RECT 427.950 643.800 430.050 645.900 ;
        RECT 451.950 643.800 454.050 645.900 ;
        RECT 457.950 645.450 460.050 645.900 ;
        RECT 463.950 645.450 466.050 645.900 ;
        RECT 457.950 644.250 466.050 645.450 ;
        RECT 457.950 643.800 460.050 644.250 ;
        RECT 463.950 643.800 466.050 644.250 ;
        RECT 475.950 645.600 478.050 645.900 ;
        RECT 479.400 645.600 480.600 647.400 ;
        RECT 475.950 644.400 480.600 645.600 ;
        RECT 502.950 645.600 505.050 645.900 ;
        RECT 506.400 645.600 507.600 649.950 ;
        RECT 502.950 644.400 507.600 645.600 ;
        RECT 511.950 645.600 514.050 646.050 ;
        RECT 517.950 645.600 520.050 645.900 ;
        RECT 511.950 644.400 520.050 645.600 ;
        RECT 475.950 643.800 478.050 644.400 ;
        RECT 502.950 643.800 505.050 644.400 ;
        RECT 511.950 643.950 514.050 644.400 ;
        RECT 517.950 643.800 520.050 644.400 ;
        RECT 550.950 645.600 553.050 646.050 ;
        RECT 562.950 645.600 565.050 645.900 ;
        RECT 550.950 644.400 565.050 645.600 ;
        RECT 550.950 643.950 553.050 644.400 ;
        RECT 562.950 643.800 565.050 644.400 ;
        RECT 571.950 645.450 574.050 645.900 ;
        RECT 577.950 645.450 580.050 645.900 ;
        RECT 571.950 644.250 580.050 645.450 ;
        RECT 590.400 645.600 591.600 650.400 ;
        RECT 610.950 649.950 613.050 652.050 ;
        RECT 633.000 651.600 637.050 652.050 ;
        RECT 632.400 649.950 637.050 651.600 ;
        RECT 691.950 649.950 694.050 652.050 ;
        RECT 697.950 651.750 700.050 652.200 ;
        RECT 703.950 651.750 706.050 652.200 ;
        RECT 697.950 650.550 706.050 651.750 ;
        RECT 697.950 650.100 700.050 650.550 ;
        RECT 703.950 650.100 706.050 650.550 ;
        RECT 748.950 649.950 751.050 652.050 ;
        RECT 766.950 650.100 769.050 652.200 ;
        RECT 790.950 651.600 793.050 652.200 ;
        RECT 802.950 651.600 805.050 652.050 ;
        RECT 790.950 650.400 805.050 651.600 ;
        RECT 790.950 650.100 793.050 650.400 ;
        RECT 611.400 646.050 612.600 649.950 ;
        RECT 616.950 648.600 619.050 649.050 ;
        RECT 632.400 648.600 633.600 649.950 ;
        RECT 616.950 647.400 633.600 648.600 ;
        RECT 637.950 648.600 640.050 649.050 ;
        RECT 692.400 648.600 693.600 649.950 ;
        RECT 637.950 647.400 693.600 648.600 ;
        RECT 616.950 646.950 619.050 647.400 ;
        RECT 598.950 645.600 601.050 646.050 ;
        RECT 590.400 644.400 601.050 645.600 ;
        RECT 571.950 643.800 574.050 644.250 ;
        RECT 577.950 643.800 580.050 644.250 ;
        RECT 598.950 643.950 601.050 644.400 ;
        RECT 610.950 643.950 613.050 646.050 ;
        RECT 626.400 645.900 627.600 647.400 ;
        RECT 637.950 646.950 640.050 647.400 ;
        RECT 625.950 643.800 628.050 645.900 ;
        RECT 643.950 645.600 646.050 646.050 ;
        RECT 652.950 645.600 655.050 645.900 ;
        RECT 688.950 645.600 691.050 645.900 ;
        RECT 643.950 644.400 691.050 645.600 ;
        RECT 643.950 643.950 646.050 644.400 ;
        RECT 652.950 643.800 655.050 644.400 ;
        RECT 688.950 643.800 691.050 644.400 ;
        RECT 700.950 645.600 703.050 645.900 ;
        RECT 706.950 645.600 709.050 646.050 ;
        RECT 712.950 645.600 715.050 645.900 ;
        RECT 700.950 644.400 715.050 645.600 ;
        RECT 700.950 643.800 703.050 644.400 ;
        RECT 706.950 643.950 709.050 644.400 ;
        RECT 712.950 643.800 715.050 644.400 ;
        RECT 718.950 645.600 721.050 645.900 ;
        RECT 733.950 645.600 736.050 646.050 ;
        RECT 718.950 644.400 736.050 645.600 ;
        RECT 718.950 643.800 721.050 644.400 ;
        RECT 733.950 643.950 736.050 644.400 ;
        RECT 749.400 643.050 750.600 649.950 ;
        RECT 751.950 645.600 754.050 645.900 ;
        RECT 760.950 645.600 763.050 646.050 ;
        RECT 767.400 645.600 768.600 650.100 ;
        RECT 802.950 649.950 805.050 650.400 ;
        RECT 835.950 650.100 838.050 652.200 ;
        RECT 865.950 650.100 868.050 652.200 ;
        RECT 874.950 651.750 877.050 652.200 ;
        RECT 883.950 651.750 886.050 652.200 ;
        RECT 874.950 650.550 886.050 651.750 ;
        RECT 874.950 650.100 877.050 650.550 ;
        RECT 883.950 650.100 886.050 650.550 ;
        RECT 751.950 644.400 768.600 645.600 ;
        RECT 781.950 645.600 784.050 646.050 ;
        RECT 787.950 645.600 790.050 645.900 ;
        RECT 781.950 644.400 790.050 645.600 ;
        RECT 751.950 643.800 754.050 644.400 ;
        RECT 760.950 643.950 763.050 644.400 ;
        RECT 781.950 643.950 784.050 644.400 ;
        RECT 787.950 643.800 790.050 644.400 ;
        RECT 836.400 643.050 837.600 650.100 ;
        RECT 866.400 645.600 867.600 650.100 ;
        RECT 892.950 649.950 895.050 652.050 ;
        RECT 893.400 646.050 894.600 649.950 ;
        RECT 886.950 645.600 889.050 645.900 ;
        RECT 866.400 644.400 889.050 645.600 ;
        RECT 886.950 643.800 889.050 644.400 ;
        RECT 892.950 643.950 895.050 646.050 ;
        RECT 343.950 641.400 351.600 642.600 ;
        RECT 442.950 642.600 445.050 643.050 ;
        RECT 481.950 642.600 484.050 643.050 ;
        RECT 442.950 641.400 484.050 642.600 ;
        RECT 343.950 640.950 346.050 641.400 ;
        RECT 442.950 640.950 445.050 641.400 ;
        RECT 481.950 640.950 484.050 641.400 ;
        RECT 541.950 642.600 544.050 643.050 ;
        RECT 547.950 642.600 550.050 643.050 ;
        RECT 541.950 641.400 550.050 642.600 ;
        RECT 541.950 640.950 544.050 641.400 ;
        RECT 547.950 640.950 550.050 641.400 ;
        RECT 661.950 642.600 664.050 643.050 ;
        RECT 673.950 642.600 676.050 643.050 ;
        RECT 661.950 641.400 676.050 642.600 ;
        RECT 661.950 640.950 664.050 641.400 ;
        RECT 673.950 640.950 676.050 641.400 ;
        RECT 748.950 640.950 751.050 643.050 ;
        RECT 835.950 640.950 838.050 643.050 ;
        RECT 16.950 639.600 19.050 640.050 ;
        RECT 97.950 639.600 100.050 640.050 ;
        RECT 16.950 638.400 100.050 639.600 ;
        RECT 16.950 637.950 19.050 638.400 ;
        RECT 97.950 637.950 100.050 638.400 ;
        RECT 160.950 639.600 163.050 640.050 ;
        RECT 184.950 639.600 187.050 640.050 ;
        RECT 160.950 638.400 187.050 639.600 ;
        RECT 160.950 637.950 163.050 638.400 ;
        RECT 184.950 637.950 187.050 638.400 ;
        RECT 193.950 639.600 196.050 640.050 ;
        RECT 238.950 639.600 241.050 640.050 ;
        RECT 193.950 638.400 241.050 639.600 ;
        RECT 193.950 637.950 196.050 638.400 ;
        RECT 238.950 637.950 241.050 638.400 ;
        RECT 370.950 639.600 373.050 640.050 ;
        RECT 376.950 639.600 379.050 640.050 ;
        RECT 406.950 639.600 409.050 640.050 ;
        RECT 370.950 638.400 409.050 639.600 ;
        RECT 370.950 637.950 373.050 638.400 ;
        RECT 376.950 637.950 379.050 638.400 ;
        RECT 406.950 637.950 409.050 638.400 ;
        RECT 466.950 639.600 469.050 640.050 ;
        RECT 478.950 639.600 481.050 640.050 ;
        RECT 466.950 638.400 481.050 639.600 ;
        RECT 466.950 637.950 469.050 638.400 ;
        RECT 478.950 637.950 481.050 638.400 ;
        RECT 508.950 639.600 511.050 640.050 ;
        RECT 520.950 639.600 523.050 640.050 ;
        RECT 529.950 639.600 532.050 640.050 ;
        RECT 508.950 638.400 519.600 639.600 ;
        RECT 508.950 637.950 511.050 638.400 ;
        RECT 31.950 636.600 34.050 637.050 ;
        RECT 67.950 636.600 70.050 637.050 ;
        RECT 31.950 635.400 70.050 636.600 ;
        RECT 31.950 634.950 34.050 635.400 ;
        RECT 67.950 634.950 70.050 635.400 ;
        RECT 124.950 636.600 127.050 637.050 ;
        RECT 175.950 636.600 178.050 637.050 ;
        RECT 124.950 635.400 178.050 636.600 ;
        RECT 124.950 634.950 127.050 635.400 ;
        RECT 175.950 634.950 178.050 635.400 ;
        RECT 301.950 636.600 304.050 637.050 ;
        RECT 310.950 636.600 313.050 637.050 ;
        RECT 319.950 636.600 322.050 637.050 ;
        RECT 301.950 635.400 322.050 636.600 ;
        RECT 301.950 634.950 304.050 635.400 ;
        RECT 310.950 634.950 313.050 635.400 ;
        RECT 319.950 634.950 322.050 635.400 ;
        RECT 409.950 636.600 412.050 637.050 ;
        RECT 415.950 636.600 418.050 637.050 ;
        RECT 463.950 636.600 466.050 637.050 ;
        RECT 409.950 635.400 466.050 636.600 ;
        RECT 409.950 634.950 412.050 635.400 ;
        RECT 415.950 634.950 418.050 635.400 ;
        RECT 463.950 634.950 466.050 635.400 ;
        RECT 502.950 636.600 505.050 637.050 ;
        RECT 518.400 636.600 519.600 638.400 ;
        RECT 520.950 638.400 532.050 639.600 ;
        RECT 548.400 639.600 549.600 640.950 ;
        RECT 595.950 639.600 598.050 640.050 ;
        RECT 548.400 638.400 598.050 639.600 ;
        RECT 520.950 637.950 523.050 638.400 ;
        RECT 529.950 637.950 532.050 638.400 ;
        RECT 595.950 637.950 598.050 638.400 ;
        RECT 601.950 639.600 604.050 640.050 ;
        RECT 637.950 639.600 640.050 640.050 ;
        RECT 646.950 639.600 649.050 640.050 ;
        RECT 601.950 638.400 649.050 639.600 ;
        RECT 601.950 637.950 604.050 638.400 ;
        RECT 637.950 637.950 640.050 638.400 ;
        RECT 646.950 637.950 649.050 638.400 ;
        RECT 658.950 639.600 661.050 640.050 ;
        RECT 673.950 639.600 676.050 639.900 ;
        RECT 658.950 638.400 676.050 639.600 ;
        RECT 658.950 637.950 661.050 638.400 ;
        RECT 673.950 637.800 676.050 638.400 ;
        RECT 688.950 639.600 691.050 640.050 ;
        RECT 703.950 639.600 706.050 640.050 ;
        RECT 688.950 638.400 706.050 639.600 ;
        RECT 688.950 637.950 691.050 638.400 ;
        RECT 703.950 637.950 706.050 638.400 ;
        RECT 721.950 639.600 724.050 640.050 ;
        RECT 727.950 639.600 730.050 640.050 ;
        RECT 745.950 639.600 748.050 639.900 ;
        RECT 721.950 638.400 730.050 639.600 ;
        RECT 721.950 637.950 724.050 638.400 ;
        RECT 727.950 637.950 730.050 638.400 ;
        RECT 734.400 638.400 748.050 639.600 ;
        RECT 529.950 636.600 532.050 636.900 ;
        RECT 502.950 635.400 513.600 636.600 ;
        RECT 518.400 635.400 532.050 636.600 ;
        RECT 502.950 634.950 505.050 635.400 ;
        RECT 247.950 633.600 250.050 634.050 ;
        RECT 265.950 633.600 268.050 634.050 ;
        RECT 295.950 633.600 298.050 634.050 ;
        RECT 247.950 632.400 298.050 633.600 ;
        RECT 247.950 631.950 250.050 632.400 ;
        RECT 265.950 631.950 268.050 632.400 ;
        RECT 295.950 631.950 298.050 632.400 ;
        RECT 328.950 633.600 331.050 634.050 ;
        RECT 385.950 633.600 388.050 634.050 ;
        RECT 328.950 632.400 388.050 633.600 ;
        RECT 328.950 631.950 331.050 632.400 ;
        RECT 385.950 631.950 388.050 632.400 ;
        RECT 481.950 633.600 484.050 634.050 ;
        RECT 493.950 633.600 496.050 634.050 ;
        RECT 505.950 633.600 508.050 634.050 ;
        RECT 481.950 632.400 508.050 633.600 ;
        RECT 512.400 633.600 513.600 635.400 ;
        RECT 529.950 634.800 532.050 635.400 ;
        RECT 583.950 636.600 586.050 637.050 ;
        RECT 589.950 636.600 592.050 637.050 ;
        RECT 583.950 635.400 592.050 636.600 ;
        RECT 583.950 634.950 586.050 635.400 ;
        RECT 589.950 634.950 592.050 635.400 ;
        RECT 679.950 636.600 682.050 637.050 ;
        RECT 694.950 636.600 697.050 637.050 ;
        RECT 679.950 635.400 697.050 636.600 ;
        RECT 679.950 634.950 682.050 635.400 ;
        RECT 694.950 634.950 697.050 635.400 ;
        RECT 706.950 636.600 709.050 637.050 ;
        RECT 734.400 636.600 735.600 638.400 ;
        RECT 745.950 637.800 748.050 638.400 ;
        RECT 814.950 639.600 817.050 640.050 ;
        RECT 823.950 639.600 826.050 640.050 ;
        RECT 814.950 638.400 826.050 639.600 ;
        RECT 814.950 637.950 817.050 638.400 ;
        RECT 823.950 637.950 826.050 638.400 ;
        RECT 832.950 639.600 835.050 640.050 ;
        RECT 844.950 639.600 847.050 640.050 ;
        RECT 832.950 638.400 847.050 639.600 ;
        RECT 832.950 637.950 835.050 638.400 ;
        RECT 844.950 637.950 847.050 638.400 ;
        RECT 883.950 639.600 886.050 640.050 ;
        RECT 892.950 639.600 895.050 640.050 ;
        RECT 883.950 638.400 895.050 639.600 ;
        RECT 883.950 637.950 886.050 638.400 ;
        RECT 892.950 637.950 895.050 638.400 ;
        RECT 706.950 635.400 735.600 636.600 ;
        RECT 748.950 636.600 751.050 637.050 ;
        RECT 769.950 636.600 772.050 637.050 ;
        RECT 748.950 635.400 772.050 636.600 ;
        RECT 706.950 634.950 709.050 635.400 ;
        RECT 748.950 634.950 751.050 635.400 ;
        RECT 769.950 634.950 772.050 635.400 ;
        RECT 664.950 633.600 667.050 634.050 ;
        RECT 512.400 632.400 667.050 633.600 ;
        RECT 481.950 631.950 484.050 632.400 ;
        RECT 493.950 631.950 496.050 632.400 ;
        RECT 505.950 631.950 508.050 632.400 ;
        RECT 664.950 631.950 667.050 632.400 ;
        RECT 742.950 633.600 745.050 634.050 ;
        RECT 754.950 633.600 757.050 634.050 ;
        RECT 742.950 632.400 757.050 633.600 ;
        RECT 742.950 631.950 745.050 632.400 ;
        RECT 754.950 631.950 757.050 632.400 ;
        RECT 805.950 633.600 808.050 634.050 ;
        RECT 877.950 633.600 880.050 634.050 ;
        RECT 805.950 632.400 880.050 633.600 ;
        RECT 805.950 631.950 808.050 632.400 ;
        RECT 877.950 631.950 880.050 632.400 ;
        RECT 22.950 630.600 25.050 631.050 ;
        RECT 94.950 630.600 97.050 631.050 ;
        RECT 22.950 629.400 97.050 630.600 ;
        RECT 22.950 628.950 25.050 629.400 ;
        RECT 94.950 628.950 97.050 629.400 ;
        RECT 136.950 630.600 139.050 631.050 ;
        RECT 142.950 630.600 145.050 631.050 ;
        RECT 136.950 629.400 145.050 630.600 ;
        RECT 136.950 628.950 139.050 629.400 ;
        RECT 142.950 628.950 145.050 629.400 ;
        RECT 175.950 630.600 178.050 631.050 ;
        RECT 190.950 630.600 193.050 631.050 ;
        RECT 175.950 629.400 193.050 630.600 ;
        RECT 175.950 628.950 178.050 629.400 ;
        RECT 190.950 628.950 193.050 629.400 ;
        RECT 424.950 630.600 427.050 631.050 ;
        RECT 436.950 630.600 439.050 631.050 ;
        RECT 424.950 629.400 439.050 630.600 ;
        RECT 424.950 628.950 427.050 629.400 ;
        RECT 436.950 628.950 439.050 629.400 ;
        RECT 487.950 630.600 490.050 631.050 ;
        RECT 526.950 630.600 529.050 631.050 ;
        RECT 487.950 629.400 529.050 630.600 ;
        RECT 487.950 628.950 490.050 629.400 ;
        RECT 526.950 628.950 529.050 629.400 ;
        RECT 679.950 630.600 682.050 631.050 ;
        RECT 727.950 630.600 730.050 631.050 ;
        RECT 679.950 629.400 730.050 630.600 ;
        RECT 679.950 628.950 682.050 629.400 ;
        RECT 727.950 628.950 730.050 629.400 ;
        RECT 739.950 630.600 742.050 631.050 ;
        RECT 757.950 630.600 760.050 631.050 ;
        RECT 739.950 629.400 760.050 630.600 ;
        RECT 739.950 628.950 742.050 629.400 ;
        RECT 757.950 628.950 760.050 629.400 ;
        RECT 766.950 630.600 769.050 631.050 ;
        RECT 793.950 630.600 796.050 631.050 ;
        RECT 766.950 629.400 796.050 630.600 ;
        RECT 766.950 628.950 769.050 629.400 ;
        RECT 793.950 628.950 796.050 629.400 ;
        RECT 868.950 630.600 871.050 631.050 ;
        RECT 874.950 630.600 877.050 631.050 ;
        RECT 880.950 630.600 883.050 631.050 ;
        RECT 868.950 629.400 883.050 630.600 ;
        RECT 868.950 628.950 871.050 629.400 ;
        RECT 874.950 628.950 877.050 629.400 ;
        RECT 880.950 628.950 883.050 629.400 ;
        RECT 355.950 627.600 358.050 628.050 ;
        RECT 397.950 627.600 400.050 628.050 ;
        RECT 355.950 626.400 400.050 627.600 ;
        RECT 355.950 625.950 358.050 626.400 ;
        RECT 397.950 625.950 400.050 626.400 ;
        RECT 427.950 627.600 430.050 628.050 ;
        RECT 469.950 627.600 472.050 628.050 ;
        RECT 427.950 626.400 472.050 627.600 ;
        RECT 427.950 625.950 430.050 626.400 ;
        RECT 469.950 625.950 472.050 626.400 ;
        RECT 607.950 627.600 610.050 628.050 ;
        RECT 631.950 627.600 634.050 628.050 ;
        RECT 607.950 626.400 634.050 627.600 ;
        RECT 607.950 625.950 610.050 626.400 ;
        RECT 631.950 625.950 634.050 626.400 ;
        RECT 745.950 627.600 748.050 628.050 ;
        RECT 757.950 627.600 760.050 627.900 ;
        RECT 745.950 626.400 760.050 627.600 ;
        RECT 745.950 625.950 748.050 626.400 ;
        RECT 757.950 625.800 760.050 626.400 ;
        RECT 40.950 624.600 43.050 625.050 ;
        RECT 85.950 624.600 88.050 625.050 ;
        RECT 40.950 623.400 88.050 624.600 ;
        RECT 40.950 622.950 43.050 623.400 ;
        RECT 85.950 622.950 88.050 623.400 ;
        RECT 349.950 624.600 352.050 625.050 ;
        RECT 370.950 624.600 373.050 625.050 ;
        RECT 412.950 624.600 415.050 625.050 ;
        RECT 349.950 623.400 373.050 624.600 ;
        RECT 349.950 622.950 352.050 623.400 ;
        RECT 370.950 622.950 373.050 623.400 ;
        RECT 374.400 623.400 415.050 624.600 ;
        RECT 13.950 621.600 16.050 622.050 ;
        RECT 91.950 621.600 94.050 622.050 ;
        RECT 13.950 620.400 94.050 621.600 ;
        RECT 13.950 619.950 16.050 620.400 ;
        RECT 91.950 619.950 94.050 620.400 ;
        RECT 115.950 621.600 118.050 622.050 ;
        RECT 124.950 621.600 127.050 622.050 ;
        RECT 115.950 620.400 127.050 621.600 ;
        RECT 115.950 619.950 118.050 620.400 ;
        RECT 124.950 619.950 127.050 620.400 ;
        RECT 163.950 621.600 166.050 622.050 ;
        RECT 220.950 621.600 223.050 622.050 ;
        RECT 232.950 621.600 235.050 622.050 ;
        RECT 163.950 620.400 235.050 621.600 ;
        RECT 163.950 619.950 166.050 620.400 ;
        RECT 220.950 619.950 223.050 620.400 ;
        RECT 232.950 619.950 235.050 620.400 ;
        RECT 283.950 621.600 286.050 622.050 ;
        RECT 374.400 621.600 375.600 623.400 ;
        RECT 412.950 622.950 415.050 623.400 ;
        RECT 436.950 624.600 439.050 625.050 ;
        RECT 550.950 624.600 553.050 625.050 ;
        RECT 436.950 623.400 553.050 624.600 ;
        RECT 436.950 622.950 439.050 623.400 ;
        RECT 550.950 622.950 553.050 623.400 ;
        RECT 646.950 624.600 649.050 625.050 ;
        RECT 706.950 624.600 709.050 625.050 ;
        RECT 646.950 623.400 709.050 624.600 ;
        RECT 646.950 622.950 649.050 623.400 ;
        RECT 706.950 622.950 709.050 623.400 ;
        RECT 283.950 620.400 375.600 621.600 ;
        RECT 391.950 621.600 394.050 622.050 ;
        RECT 406.950 621.600 409.050 622.050 ;
        RECT 424.950 621.600 427.050 622.050 ;
        RECT 391.950 620.400 427.050 621.600 ;
        RECT 283.950 619.950 286.050 620.400 ;
        RECT 391.950 619.950 394.050 620.400 ;
        RECT 406.950 619.950 409.050 620.400 ;
        RECT 424.950 619.950 427.050 620.400 ;
        RECT 433.950 621.600 436.050 622.050 ;
        RECT 553.950 621.600 556.050 622.050 ;
        RECT 433.950 620.400 556.050 621.600 ;
        RECT 433.950 619.950 436.050 620.400 ;
        RECT 553.950 619.950 556.050 620.400 ;
        RECT 634.950 621.600 637.050 622.050 ;
        RECT 667.950 621.600 670.050 622.050 ;
        RECT 634.950 620.400 670.050 621.600 ;
        RECT 634.950 619.950 637.050 620.400 ;
        RECT 667.950 619.950 670.050 620.400 ;
        RECT 712.950 621.600 715.050 622.050 ;
        RECT 718.950 621.600 721.050 622.050 ;
        RECT 712.950 620.400 721.050 621.600 ;
        RECT 712.950 619.950 715.050 620.400 ;
        RECT 718.950 619.950 721.050 620.400 ;
        RECT 724.950 621.600 727.050 622.050 ;
        RECT 742.950 621.600 745.050 622.050 ;
        RECT 769.950 621.600 772.050 622.050 ;
        RECT 724.950 620.400 745.050 621.600 ;
        RECT 724.950 619.950 727.050 620.400 ;
        RECT 742.950 619.950 745.050 620.400 ;
        RECT 752.400 620.400 772.050 621.600 ;
        RECT 94.950 618.600 97.050 619.050 ;
        RECT 145.950 618.600 148.050 619.050 ;
        RECT 94.950 617.400 148.050 618.600 ;
        RECT 94.950 616.950 97.050 617.400 ;
        RECT 145.950 616.950 148.050 617.400 ;
        RECT 157.950 618.600 160.050 619.050 ;
        RECT 184.950 618.600 187.050 619.050 ;
        RECT 157.950 617.400 187.050 618.600 ;
        RECT 157.950 616.950 160.050 617.400 ;
        RECT 184.950 616.950 187.050 617.400 ;
        RECT 451.950 618.600 454.050 619.050 ;
        RECT 475.950 618.600 478.050 619.050 ;
        RECT 451.950 617.400 478.050 618.600 ;
        RECT 451.950 616.950 454.050 617.400 ;
        RECT 475.950 616.950 478.050 617.400 ;
        RECT 484.950 618.600 487.050 619.050 ;
        RECT 547.950 618.600 550.050 619.050 ;
        RECT 484.950 617.400 550.050 618.600 ;
        RECT 484.950 616.950 487.050 617.400 ;
        RECT 547.950 616.950 550.050 617.400 ;
        RECT 586.950 618.600 589.050 619.050 ;
        RECT 598.950 618.600 601.050 619.050 ;
        RECT 622.950 618.600 625.050 619.050 ;
        RECT 586.950 617.400 625.050 618.600 ;
        RECT 586.950 616.950 589.050 617.400 ;
        RECT 598.950 616.950 601.050 617.400 ;
        RECT 622.950 616.950 625.050 617.400 ;
        RECT 631.950 618.600 634.050 619.050 ;
        RECT 694.950 618.600 697.050 619.050 ;
        RECT 631.950 617.400 697.050 618.600 ;
        RECT 631.950 616.950 634.050 617.400 ;
        RECT 694.950 616.950 697.050 617.400 ;
        RECT 703.950 618.600 706.050 619.050 ;
        RECT 752.400 618.600 753.600 620.400 ;
        RECT 769.950 619.950 772.050 620.400 ;
        RECT 787.950 621.600 790.050 622.050 ;
        RECT 871.950 621.600 874.050 622.050 ;
        RECT 787.950 620.400 874.050 621.600 ;
        RECT 787.950 619.950 790.050 620.400 ;
        RECT 871.950 619.950 874.050 620.400 ;
        RECT 703.950 617.400 753.600 618.600 ;
        RECT 793.950 618.600 796.050 619.050 ;
        RECT 805.950 618.600 808.050 619.050 ;
        RECT 817.950 618.600 820.050 619.050 ;
        RECT 793.950 617.400 820.050 618.600 ;
        RECT 703.950 616.950 706.050 617.400 ;
        RECT 793.950 616.950 796.050 617.400 ;
        RECT 805.950 616.950 808.050 617.400 ;
        RECT 817.950 616.950 820.050 617.400 ;
        RECT 79.950 615.600 82.050 616.050 ;
        RECT 85.950 615.600 88.050 615.900 ;
        RECT 79.950 614.400 88.050 615.600 ;
        RECT 79.950 613.950 82.050 614.400 ;
        RECT 85.950 613.800 88.050 614.400 ;
        RECT 289.950 615.600 292.050 616.050 ;
        RECT 358.950 615.600 361.050 616.050 ;
        RECT 424.950 615.600 427.050 616.050 ;
        RECT 433.950 615.600 436.050 616.050 ;
        RECT 289.950 614.400 436.050 615.600 ;
        RECT 289.950 613.950 292.050 614.400 ;
        RECT 358.950 613.950 361.050 614.400 ;
        RECT 424.950 613.950 427.050 614.400 ;
        RECT 433.950 613.950 436.050 614.400 ;
        RECT 733.950 615.600 736.050 616.050 ;
        RECT 763.950 615.600 766.050 616.050 ;
        RECT 793.950 615.600 796.050 615.900 ;
        RECT 811.950 615.600 814.050 616.050 ;
        RECT 733.950 614.400 814.050 615.600 ;
        RECT 733.950 613.950 736.050 614.400 ;
        RECT 763.950 613.950 766.050 614.400 ;
        RECT 793.950 613.800 796.050 614.400 ;
        RECT 811.950 613.950 814.050 614.400 ;
        RECT 859.950 615.600 862.050 616.050 ;
        RECT 874.950 615.600 877.050 616.050 ;
        RECT 886.950 615.600 889.050 616.050 ;
        RECT 859.950 614.400 889.050 615.600 ;
        RECT 859.950 613.950 862.050 614.400 ;
        RECT 874.950 613.950 877.050 614.400 ;
        RECT 886.950 613.950 889.050 614.400 ;
        RECT 154.950 612.600 157.050 613.050 ;
        RECT 187.950 612.600 190.050 613.050 ;
        RECT 154.950 611.400 190.050 612.600 ;
        RECT 154.950 610.950 157.050 611.400 ;
        RECT 187.950 610.950 190.050 611.400 ;
        RECT 214.950 612.600 217.050 613.050 ;
        RECT 229.950 612.600 232.050 613.050 ;
        RECT 214.950 611.400 232.050 612.600 ;
        RECT 214.950 610.950 217.050 611.400 ;
        RECT 229.950 610.950 232.050 611.400 ;
        RECT 382.950 612.600 385.050 613.050 ;
        RECT 421.950 612.600 424.050 613.050 ;
        RECT 430.950 612.600 433.050 613.050 ;
        RECT 559.950 612.600 562.050 613.050 ;
        RECT 382.950 611.400 433.050 612.600 ;
        RECT 382.950 610.950 385.050 611.400 ;
        RECT 421.950 610.950 424.050 611.400 ;
        RECT 430.950 610.950 433.050 611.400 ;
        RECT 548.400 611.400 562.050 612.600 ;
        RECT 61.950 609.600 64.050 610.050 ;
        RECT 163.950 609.600 166.050 610.050 ;
        RECT 61.950 608.400 166.050 609.600 ;
        RECT 61.950 607.950 64.050 608.400 ;
        RECT 163.950 607.950 166.050 608.400 ;
        RECT 184.950 609.600 187.050 610.050 ;
        RECT 196.950 609.600 199.050 610.050 ;
        RECT 184.950 608.400 199.050 609.600 ;
        RECT 184.950 607.950 187.050 608.400 ;
        RECT 196.950 607.950 199.050 608.400 ;
        RECT 235.950 609.600 238.050 610.050 ;
        RECT 247.950 609.600 250.050 610.050 ;
        RECT 235.950 608.400 250.050 609.600 ;
        RECT 235.950 607.950 238.050 608.400 ;
        RECT 247.950 607.950 250.050 608.400 ;
        RECT 322.950 609.600 325.050 610.050 ;
        RECT 346.950 609.600 349.050 610.050 ;
        RECT 379.950 609.600 382.050 610.050 ;
        RECT 322.950 608.400 382.050 609.600 ;
        RECT 322.950 607.950 325.050 608.400 ;
        RECT 346.950 607.950 349.050 608.400 ;
        RECT 379.950 607.950 382.050 608.400 ;
        RECT 502.950 609.600 505.050 610.050 ;
        RECT 535.950 609.600 538.050 610.050 ;
        RECT 548.400 609.600 549.600 611.400 ;
        RECT 559.950 610.950 562.050 611.400 ;
        RECT 640.950 612.600 643.050 613.050 ;
        RECT 655.950 612.600 658.050 613.050 ;
        RECT 640.950 611.400 658.050 612.600 ;
        RECT 640.950 610.950 643.050 611.400 ;
        RECT 655.950 610.950 658.050 611.400 ;
        RECT 775.950 612.600 778.050 613.050 ;
        RECT 790.950 612.600 793.050 613.050 ;
        RECT 775.950 611.400 793.050 612.600 ;
        RECT 775.950 610.950 778.050 611.400 ;
        RECT 790.950 610.950 793.050 611.400 ;
        RECT 502.950 608.400 538.050 609.600 ;
        RECT 502.950 607.950 505.050 608.400 ;
        RECT 535.950 607.950 538.050 608.400 ;
        RECT 545.400 608.400 549.600 609.600 ;
        RECT 682.950 609.600 685.050 610.050 ;
        RECT 748.950 609.600 751.050 610.050 ;
        RECT 757.950 609.600 760.050 610.050 ;
        RECT 682.950 608.400 693.600 609.600 ;
        RECT 25.950 606.600 28.050 607.050 ;
        RECT 14.400 605.400 28.050 606.600 ;
        RECT 14.400 598.050 15.600 605.400 ;
        RECT 25.950 604.950 28.050 605.400 ;
        RECT 91.950 606.600 94.050 607.050 ;
        RECT 100.950 606.750 103.050 607.200 ;
        RECT 109.950 606.750 112.050 607.200 ;
        RECT 91.950 605.400 99.600 606.600 ;
        RECT 91.950 604.950 94.050 605.400 ;
        RECT 25.950 600.600 28.050 601.050 ;
        RECT 31.950 600.600 34.050 601.050 ;
        RECT 98.400 600.900 99.600 605.400 ;
        RECT 100.950 605.550 112.050 606.750 ;
        RECT 100.950 605.100 103.050 605.550 ;
        RECT 109.950 605.100 112.050 605.550 ;
        RECT 118.950 605.100 121.050 607.200 ;
        RECT 205.950 607.050 208.050 607.500 ;
        RECT 214.950 607.050 217.050 607.500 ;
        RECT 205.950 605.850 217.050 607.050 ;
        RECT 205.950 605.400 208.050 605.850 ;
        RECT 214.950 605.400 217.050 605.850 ;
        RECT 316.950 605.100 319.050 607.200 ;
        RECT 358.950 605.100 361.050 607.200 ;
        RECT 451.950 606.600 454.050 607.200 ;
        RECT 440.400 605.400 454.050 606.600 ;
        RECT 25.950 599.400 34.050 600.600 ;
        RECT 25.950 598.950 28.050 599.400 ;
        RECT 31.950 598.950 34.050 599.400 ;
        RECT 97.950 598.800 100.050 600.900 ;
        RECT 103.950 600.600 106.050 600.900 ;
        RECT 119.400 600.600 120.600 605.100 ;
        RECT 103.950 599.400 120.600 600.600 ;
        RECT 121.950 600.600 124.050 600.900 ;
        RECT 133.950 600.600 136.050 601.050 ;
        RECT 121.950 599.400 136.050 600.600 ;
        RECT 103.950 598.800 106.050 599.400 ;
        RECT 121.950 598.800 124.050 599.400 ;
        RECT 133.950 598.950 136.050 599.400 ;
        RECT 148.950 600.450 151.050 600.900 ;
        RECT 154.950 600.600 157.050 600.900 ;
        RECT 160.950 600.600 163.050 601.050 ;
        RECT 154.950 600.450 163.050 600.600 ;
        RECT 148.950 599.400 163.050 600.450 ;
        RECT 148.950 599.250 157.050 599.400 ;
        RECT 148.950 598.800 151.050 599.250 ;
        RECT 154.950 598.800 157.050 599.250 ;
        RECT 160.950 598.950 163.050 599.400 ;
        RECT 169.950 600.450 172.050 600.900 ;
        RECT 175.950 600.450 178.050 601.050 ;
        RECT 208.950 600.450 211.050 600.900 ;
        RECT 169.950 599.250 211.050 600.450 ;
        RECT 169.950 598.800 172.050 599.250 ;
        RECT 175.950 598.950 178.050 599.250 ;
        RECT 208.950 598.800 211.050 599.250 ;
        RECT 214.950 600.600 217.050 601.050 ;
        RECT 244.950 600.600 247.050 600.900 ;
        RECT 214.950 599.400 247.050 600.600 ;
        RECT 317.400 600.600 318.600 605.100 ;
        RECT 325.950 600.600 328.050 601.050 ;
        RECT 317.400 599.400 328.050 600.600 ;
        RECT 214.950 598.950 217.050 599.400 ;
        RECT 244.950 598.800 247.050 599.400 ;
        RECT 325.950 598.950 328.050 599.400 ;
        RECT 359.400 598.050 360.600 605.100 ;
        RECT 440.400 603.600 441.600 605.400 ;
        RECT 451.950 605.100 454.050 605.400 ;
        RECT 472.950 605.100 475.050 607.200 ;
        RECT 496.950 605.400 499.050 607.500 ;
        RECT 422.400 602.400 441.600 603.600 ;
        RECT 373.950 600.450 376.050 600.900 ;
        RECT 382.950 600.450 385.050 600.900 ;
        RECT 373.950 599.250 385.050 600.450 ;
        RECT 373.950 598.800 376.050 599.250 ;
        RECT 382.950 598.800 385.050 599.250 ;
        RECT 397.950 600.600 400.050 601.050 ;
        RECT 412.950 600.600 415.050 600.900 ;
        RECT 422.400 600.600 423.600 602.400 ;
        RECT 397.950 599.400 423.600 600.600 ;
        RECT 397.950 598.950 400.050 599.400 ;
        RECT 412.950 598.800 415.050 599.400 ;
        RECT 473.400 598.050 474.600 605.100 ;
        RECT 475.950 600.600 478.050 600.900 ;
        RECT 497.400 600.600 498.600 605.400 ;
        RECT 517.950 604.950 520.050 607.050 ;
        RECT 518.400 600.600 519.600 604.950 ;
        RECT 475.950 599.400 498.600 600.600 ;
        RECT 514.950 599.400 519.600 600.600 ;
        RECT 538.950 600.600 541.050 600.900 ;
        RECT 545.400 600.600 546.600 608.400 ;
        RECT 682.950 607.950 685.050 608.400 ;
        RECT 550.950 605.400 553.050 607.500 ;
        RECT 568.950 606.600 571.050 607.050 ;
        RECT 601.950 606.750 604.050 607.200 ;
        RECT 628.950 606.750 631.050 607.200 ;
        RECT 601.950 606.600 631.050 606.750 ;
        RECT 568.950 605.550 631.050 606.600 ;
        RECT 568.950 605.400 604.050 605.550 ;
        RECT 538.950 599.400 546.600 600.600 ;
        RECT 475.950 598.800 478.050 599.400 ;
        RECT 514.950 598.500 517.050 599.400 ;
        RECT 538.950 598.800 541.050 599.400 ;
        RECT 13.950 595.950 16.050 598.050 ;
        RECT 211.950 597.600 214.050 598.050 ;
        RECT 250.950 597.600 253.050 598.050 ;
        RECT 256.950 597.600 259.050 598.050 ;
        RECT 211.950 596.400 259.050 597.600 ;
        RECT 211.950 595.950 214.050 596.400 ;
        RECT 250.950 595.950 253.050 596.400 ;
        RECT 256.950 595.950 259.050 596.400 ;
        RECT 331.950 597.600 334.050 598.050 ;
        RECT 331.950 596.400 345.600 597.600 ;
        RECT 331.950 595.950 334.050 596.400 ;
        RECT 28.950 594.600 31.050 595.050 ;
        RECT 55.950 594.600 58.050 595.050 ;
        RECT 103.950 594.600 106.050 595.050 ;
        RECT 28.950 593.400 106.050 594.600 ;
        RECT 28.950 592.950 31.050 593.400 ;
        RECT 55.950 592.950 58.050 593.400 ;
        RECT 103.950 592.950 106.050 593.400 ;
        RECT 226.950 594.600 229.050 595.050 ;
        RECT 238.950 594.600 241.050 595.050 ;
        RECT 226.950 593.400 241.050 594.600 ;
        RECT 226.950 592.950 229.050 593.400 ;
        RECT 238.950 592.950 241.050 593.400 ;
        RECT 268.950 594.600 271.050 595.050 ;
        RECT 292.950 594.600 295.050 595.050 ;
        RECT 322.950 594.600 325.050 595.050 ;
        RECT 268.950 593.400 312.600 594.600 ;
        RECT 268.950 592.950 271.050 593.400 ;
        RECT 292.950 592.950 295.050 593.400 ;
        RECT 16.950 591.600 19.050 592.050 ;
        RECT 19.950 591.600 22.050 592.050 ;
        RECT 49.950 591.600 52.050 592.050 ;
        RECT 73.950 591.600 76.050 592.050 ;
        RECT 16.950 590.400 76.050 591.600 ;
        RECT 16.950 589.950 19.050 590.400 ;
        RECT 19.950 589.950 22.050 590.400 ;
        RECT 49.950 589.950 52.050 590.400 ;
        RECT 73.950 589.950 76.050 590.400 ;
        RECT 109.950 591.600 112.050 592.050 ;
        RECT 151.950 591.600 154.050 592.050 ;
        RECT 109.950 590.400 154.050 591.600 ;
        RECT 311.400 591.600 312.600 593.400 ;
        RECT 317.400 593.400 325.050 594.600 ;
        RECT 344.400 594.600 345.600 596.400 ;
        RECT 358.950 595.950 361.050 598.050 ;
        RECT 472.950 595.950 475.050 598.050 ;
        RECT 520.950 597.600 523.050 597.900 ;
        RECT 526.950 597.600 529.050 598.050 ;
        RECT 520.950 596.400 529.050 597.600 ;
        RECT 551.400 597.600 552.600 605.400 ;
        RECT 568.950 604.950 571.050 605.400 ;
        RECT 601.950 605.100 604.050 605.400 ;
        RECT 628.950 605.100 631.050 605.550 ;
        RECT 640.950 605.100 643.050 607.200 ;
        RECT 646.950 605.100 649.050 607.200 ;
        RECT 661.950 605.100 664.050 607.200 ;
        RECT 679.950 606.600 682.050 607.050 ;
        RECT 674.400 605.400 682.050 606.600 ;
        RECT 565.950 603.600 568.050 604.050 ;
        RECT 641.400 603.600 642.600 605.100 ;
        RECT 565.950 602.400 642.600 603.600 ;
        RECT 565.950 601.950 568.050 602.400 ;
        RECT 578.400 600.600 579.600 602.400 ;
        RECT 598.950 600.600 601.050 600.900 ;
        RECT 610.950 600.600 613.050 601.050 ;
        RECT 577.950 598.500 580.050 600.600 ;
        RECT 598.950 599.400 613.050 600.600 ;
        RECT 598.950 598.800 601.050 599.400 ;
        RECT 610.950 598.950 613.050 599.400 ;
        RECT 625.950 600.600 628.050 600.900 ;
        RECT 647.400 600.600 648.600 605.100 ;
        RECT 655.950 600.600 658.050 601.050 ;
        RECT 625.950 599.400 658.050 600.600 ;
        RECT 662.400 600.600 663.600 605.100 ;
        RECT 670.950 600.600 673.050 601.050 ;
        RECT 662.400 599.400 673.050 600.600 ;
        RECT 625.950 598.800 628.050 599.400 ;
        RECT 559.950 597.600 562.050 598.050 ;
        RECT 551.400 596.400 562.050 597.600 ;
        RECT 520.950 595.800 523.050 596.400 ;
        RECT 526.950 595.950 529.050 596.400 ;
        RECT 559.950 595.950 562.050 596.400 ;
        RECT 628.950 595.950 631.050 599.400 ;
        RECT 655.950 598.950 658.050 599.400 ;
        RECT 670.950 598.950 673.050 599.400 ;
        RECT 664.950 597.600 667.050 598.050 ;
        RECT 674.400 597.600 675.600 605.400 ;
        RECT 679.950 604.950 682.050 605.400 ;
        RECT 692.400 601.050 693.600 608.400 ;
        RECT 748.950 608.400 760.050 609.600 ;
        RECT 748.950 607.950 751.050 608.400 ;
        RECT 757.950 607.950 760.050 608.400 ;
        RECT 796.950 609.600 799.050 610.050 ;
        RECT 823.950 609.600 826.050 610.050 ;
        RECT 796.950 608.400 826.050 609.600 ;
        RECT 796.950 607.950 799.050 608.400 ;
        RECT 823.950 607.950 826.050 608.400 ;
        RECT 709.950 606.600 712.050 607.200 ;
        RECT 707.400 605.400 712.050 606.600 ;
        RECT 707.400 601.050 708.600 605.400 ;
        RECT 709.950 605.100 712.050 605.400 ;
        RECT 766.950 603.600 769.050 607.050 ;
        RECT 781.950 605.100 784.050 607.200 ;
        RECT 755.400 603.000 769.050 603.600 ;
        RECT 782.400 603.600 783.600 605.100 ;
        RECT 793.950 603.600 796.050 607.050 ;
        RECT 802.950 606.600 805.050 607.050 ;
        RECT 808.950 606.600 811.050 607.050 ;
        RECT 802.950 605.400 811.050 606.600 ;
        RECT 802.950 604.950 805.050 605.400 ;
        RECT 808.950 604.950 811.050 605.400 ;
        RECT 814.950 604.950 817.050 607.050 ;
        RECT 838.950 605.100 841.050 607.200 ;
        RECT 844.950 605.100 847.050 607.200 ;
        RECT 850.950 606.600 853.050 607.050 ;
        RECT 856.950 606.600 859.050 607.050 ;
        RECT 850.950 605.400 859.050 606.600 ;
        RECT 782.400 603.000 786.600 603.600 ;
        RECT 793.950 603.000 798.600 603.600 ;
        RECT 755.400 602.400 768.600 603.000 ;
        RECT 782.400 602.400 787.050 603.000 ;
        RECT 794.400 602.400 798.600 603.000 ;
        RECT 691.950 598.950 694.050 601.050 ;
        RECT 706.950 598.950 709.050 601.050 ;
        RECT 755.400 600.900 756.600 602.400 ;
        RECT 727.950 600.450 730.050 600.900 ;
        RECT 733.950 600.450 736.050 600.900 ;
        RECT 727.950 599.250 736.050 600.450 ;
        RECT 727.950 598.800 730.050 599.250 ;
        RECT 733.950 598.800 736.050 599.250 ;
        RECT 754.950 598.800 757.050 600.900 ;
        RECT 784.950 598.950 787.050 602.400 ;
        RECT 797.400 600.900 798.600 602.400 ;
        RECT 664.950 596.400 675.600 597.600 ;
        RECT 682.950 597.600 685.050 598.050 ;
        RECT 694.950 597.600 697.050 598.050 ;
        RECT 682.950 596.400 697.050 597.600 ;
        RECT 664.950 595.950 667.050 596.400 ;
        RECT 682.950 595.950 685.050 596.400 ;
        RECT 694.950 595.950 697.050 596.400 ;
        RECT 742.950 597.600 745.050 598.050 ;
        RECT 785.400 597.600 786.600 598.950 ;
        RECT 796.950 598.800 799.050 600.900 ;
        RECT 802.950 600.600 805.050 601.050 ;
        RECT 815.400 600.600 816.600 604.950 ;
        RECT 839.400 601.050 840.600 605.100 ;
        RECT 826.950 600.600 829.050 600.900 ;
        RECT 802.950 599.400 816.600 600.600 ;
        RECT 818.400 599.400 829.050 600.600 ;
        RECT 802.950 598.950 805.050 599.400 ;
        RECT 742.950 596.400 753.600 597.600 ;
        RECT 742.950 595.950 745.050 596.400 ;
        RECT 361.950 594.600 364.050 595.050 ;
        RECT 344.400 593.400 364.050 594.600 ;
        RECT 317.400 591.600 318.600 593.400 ;
        RECT 322.950 592.950 325.050 593.400 ;
        RECT 361.950 592.950 364.050 593.400 ;
        RECT 484.950 594.600 487.050 595.050 ;
        RECT 529.950 594.600 532.050 595.050 ;
        RECT 484.950 593.400 532.050 594.600 ;
        RECT 484.950 592.950 487.050 593.400 ;
        RECT 529.950 592.950 532.050 593.400 ;
        RECT 616.950 594.600 619.050 595.050 ;
        RECT 625.950 594.600 628.050 595.050 ;
        RECT 616.950 593.400 628.050 594.600 ;
        RECT 616.950 592.950 619.050 593.400 ;
        RECT 625.950 592.950 628.050 593.400 ;
        RECT 634.950 594.600 637.050 595.050 ;
        RECT 643.950 594.600 646.050 595.050 ;
        RECT 634.950 593.400 646.050 594.600 ;
        RECT 634.950 592.950 637.050 593.400 ;
        RECT 643.950 592.950 646.050 593.400 ;
        RECT 670.950 594.600 673.050 595.050 ;
        RECT 679.950 594.600 682.050 595.050 ;
        RECT 670.950 593.400 682.050 594.600 ;
        RECT 670.950 592.950 673.050 593.400 ;
        RECT 679.950 592.950 682.050 593.400 ;
        RECT 706.950 594.600 709.050 595.050 ;
        RECT 724.950 594.600 727.050 595.050 ;
        RECT 706.950 593.400 727.050 594.600 ;
        RECT 706.950 592.950 709.050 593.400 ;
        RECT 724.950 592.950 727.050 593.400 ;
        RECT 733.950 594.600 736.050 594.900 ;
        RECT 739.950 594.600 742.050 595.050 ;
        RECT 733.950 593.400 742.050 594.600 ;
        RECT 752.400 594.600 753.600 596.400 ;
        RECT 764.400 596.400 786.600 597.600 ;
        RECT 811.950 597.600 814.050 598.050 ;
        RECT 818.400 597.600 819.600 599.400 ;
        RECT 826.950 598.800 829.050 599.400 ;
        RECT 835.950 599.400 840.600 601.050 ;
        RECT 835.950 598.950 840.000 599.400 ;
        RECT 811.950 596.400 819.600 597.600 ;
        RECT 764.400 594.600 765.600 596.400 ;
        RECT 811.950 595.950 814.050 596.400 ;
        RECT 845.400 595.050 846.600 605.100 ;
        RECT 850.950 604.950 853.050 605.400 ;
        RECT 856.950 604.950 859.050 605.400 ;
        RECT 862.950 604.950 865.050 607.050 ;
        RECT 877.950 604.950 880.050 607.050 ;
        RECT 847.950 600.600 850.050 600.900 ;
        RECT 853.950 600.600 856.050 601.050 ;
        RECT 847.950 599.400 856.050 600.600 ;
        RECT 863.400 600.600 864.600 604.950 ;
        RECT 878.400 601.050 879.600 604.950 ;
        RECT 871.950 600.600 874.050 600.900 ;
        RECT 863.400 599.400 874.050 600.600 ;
        RECT 847.950 598.800 850.050 599.400 ;
        RECT 853.950 598.950 856.050 599.400 ;
        RECT 871.950 598.800 874.050 599.400 ;
        RECT 877.950 598.950 880.050 601.050 ;
        RECT 880.950 597.600 883.050 598.050 ;
        RECT 895.950 597.600 898.050 598.050 ;
        RECT 880.950 596.400 898.050 597.600 ;
        RECT 880.950 595.950 883.050 596.400 ;
        RECT 895.950 595.950 898.050 596.400 ;
        RECT 752.400 593.400 765.600 594.600 ;
        RECT 772.950 594.600 775.050 595.050 ;
        RECT 787.950 594.600 790.050 595.050 ;
        RECT 772.950 593.400 790.050 594.600 ;
        RECT 733.950 592.800 736.050 593.400 ;
        RECT 739.950 592.950 742.050 593.400 ;
        RECT 772.950 592.950 775.050 593.400 ;
        RECT 787.950 592.950 790.050 593.400 ;
        RECT 841.950 593.400 846.600 595.050 ;
        RECT 865.950 594.600 868.050 595.050 ;
        RECT 871.950 594.600 874.050 595.050 ;
        RECT 865.950 593.400 874.050 594.600 ;
        RECT 841.950 592.950 846.000 593.400 ;
        RECT 865.950 592.950 868.050 593.400 ;
        RECT 871.950 592.950 874.050 593.400 ;
        RECT 311.400 590.400 318.600 591.600 ;
        RECT 328.950 591.600 331.050 592.050 ;
        RECT 340.950 591.600 343.050 592.050 ;
        RECT 388.950 591.600 391.050 592.050 ;
        RECT 589.950 591.600 592.050 592.050 ;
        RECT 328.950 590.400 391.050 591.600 ;
        RECT 109.950 589.950 112.050 590.400 ;
        RECT 151.950 589.950 154.050 590.400 ;
        RECT 328.950 589.950 331.050 590.400 ;
        RECT 340.950 589.950 343.050 590.400 ;
        RECT 388.950 589.950 391.050 590.400 ;
        RECT 488.400 590.400 592.050 591.600 ;
        RECT 79.950 588.600 82.050 589.050 ;
        RECT 85.950 588.600 88.050 589.050 ;
        RECT 79.950 587.400 88.050 588.600 ;
        RECT 79.950 586.950 82.050 587.400 ;
        RECT 85.950 586.950 88.050 587.400 ;
        RECT 214.950 588.600 217.050 589.050 ;
        RECT 229.950 588.600 232.050 589.050 ;
        RECT 214.950 587.400 232.050 588.600 ;
        RECT 214.950 586.950 217.050 587.400 ;
        RECT 229.950 586.950 232.050 587.400 ;
        RECT 235.950 588.600 238.050 589.050 ;
        RECT 247.950 588.600 250.050 589.050 ;
        RECT 235.950 587.400 250.050 588.600 ;
        RECT 235.950 586.950 238.050 587.400 ;
        RECT 247.950 586.950 250.050 587.400 ;
        RECT 286.950 588.600 289.050 589.050 ;
        RECT 298.950 588.600 301.050 589.050 ;
        RECT 307.950 588.600 310.050 589.050 ;
        RECT 319.950 588.600 322.050 589.050 ;
        RECT 488.400 588.600 489.600 590.400 ;
        RECT 589.950 589.950 592.050 590.400 ;
        RECT 619.950 591.600 622.050 592.050 ;
        RECT 631.950 591.600 634.050 592.050 ;
        RECT 619.950 590.400 634.050 591.600 ;
        RECT 619.950 589.950 622.050 590.400 ;
        RECT 631.950 589.950 634.050 590.400 ;
        RECT 667.950 591.600 670.050 592.050 ;
        RECT 676.950 591.600 679.050 592.050 ;
        RECT 721.950 591.600 724.050 592.050 ;
        RECT 667.950 590.400 724.050 591.600 ;
        RECT 667.950 589.950 670.050 590.400 ;
        RECT 676.950 589.950 679.050 590.400 ;
        RECT 721.950 589.950 724.050 590.400 ;
        RECT 748.950 591.600 751.050 592.050 ;
        RECT 760.950 591.600 763.050 592.050 ;
        RECT 778.950 591.600 781.050 592.050 ;
        RECT 748.950 590.400 781.050 591.600 ;
        RECT 748.950 589.950 751.050 590.400 ;
        RECT 760.950 589.950 763.050 590.400 ;
        RECT 778.950 589.950 781.050 590.400 ;
        RECT 820.950 591.600 823.050 592.050 ;
        RECT 826.800 591.600 828.900 592.050 ;
        RECT 820.950 590.400 828.900 591.600 ;
        RECT 820.950 589.950 823.050 590.400 ;
        RECT 826.800 589.950 828.900 590.400 ;
        RECT 829.950 591.600 832.050 592.050 ;
        RECT 844.950 591.600 847.050 592.050 ;
        RECT 829.950 590.400 847.050 591.600 ;
        RECT 829.950 589.950 832.050 590.400 ;
        RECT 844.950 589.950 847.050 590.400 ;
        RECT 883.950 591.600 886.050 592.050 ;
        RECT 892.950 591.600 895.050 592.050 ;
        RECT 883.950 590.400 895.050 591.600 ;
        RECT 883.950 589.950 886.050 590.400 ;
        RECT 892.950 589.950 895.050 590.400 ;
        RECT 286.950 587.400 322.050 588.600 ;
        RECT 286.950 586.950 289.050 587.400 ;
        RECT 298.950 586.950 301.050 587.400 ;
        RECT 307.950 586.950 310.050 587.400 ;
        RECT 319.950 586.950 322.050 587.400 ;
        RECT 407.400 587.400 489.600 588.600 ;
        RECT 544.950 588.600 547.050 589.050 ;
        RECT 568.950 588.600 571.050 589.050 ;
        RECT 544.950 587.400 571.050 588.600 ;
        RECT 58.950 585.600 61.050 586.050 ;
        RECT 268.950 585.600 271.050 586.050 ;
        RECT 58.950 584.400 271.050 585.600 ;
        RECT 58.950 583.950 61.050 584.400 ;
        RECT 268.950 583.950 271.050 584.400 ;
        RECT 385.950 585.600 388.050 586.050 ;
        RECT 403.950 585.600 406.050 586.050 ;
        RECT 407.400 585.600 408.600 587.400 ;
        RECT 544.950 586.950 547.050 587.400 ;
        RECT 568.950 586.950 571.050 587.400 ;
        RECT 592.950 588.600 595.050 589.050 ;
        RECT 727.950 588.600 730.050 589.050 ;
        RECT 592.950 587.400 730.050 588.600 ;
        RECT 592.950 586.950 595.050 587.400 ;
        RECT 727.950 586.950 730.050 587.400 ;
        RECT 832.950 588.600 835.050 589.050 ;
        RECT 838.950 588.600 841.050 589.050 ;
        RECT 832.950 587.400 841.050 588.600 ;
        RECT 832.950 586.950 835.050 587.400 ;
        RECT 838.950 586.950 841.050 587.400 ;
        RECT 385.950 584.400 408.600 585.600 ;
        RECT 532.950 585.600 535.050 586.050 ;
        RECT 562.950 585.600 565.050 586.050 ;
        RECT 532.950 584.400 565.050 585.600 ;
        RECT 385.950 583.950 388.050 584.400 ;
        RECT 403.950 583.950 406.050 584.400 ;
        RECT 532.950 583.950 535.050 584.400 ;
        RECT 562.950 583.950 565.050 584.400 ;
        RECT 664.950 585.600 667.050 586.050 ;
        RECT 670.950 585.600 673.050 586.050 ;
        RECT 664.950 584.400 673.050 585.600 ;
        RECT 664.950 583.950 667.050 584.400 ;
        RECT 670.950 583.950 673.050 584.400 ;
        RECT 679.950 585.600 682.050 586.050 ;
        RECT 712.950 585.600 715.050 586.050 ;
        RECT 679.950 584.400 715.050 585.600 ;
        RECT 679.950 583.950 682.050 584.400 ;
        RECT 712.950 583.950 715.050 584.400 ;
        RECT 736.950 585.600 739.050 586.050 ;
        RECT 751.950 585.600 754.050 586.050 ;
        RECT 736.950 584.400 754.050 585.600 ;
        RECT 736.950 583.950 739.050 584.400 ;
        RECT 751.950 583.950 754.050 584.400 ;
        RECT 784.950 585.600 787.050 586.050 ;
        RECT 805.950 585.600 808.050 586.050 ;
        RECT 784.950 584.400 808.050 585.600 ;
        RECT 784.950 583.950 787.050 584.400 ;
        RECT 805.950 583.950 808.050 584.400 ;
        RECT 826.950 585.600 829.050 586.050 ;
        RECT 862.950 585.600 865.050 586.050 ;
        RECT 826.950 584.400 865.050 585.600 ;
        RECT 826.950 583.950 829.050 584.400 ;
        RECT 862.950 583.950 865.050 584.400 ;
        RECT 868.950 585.600 871.050 586.050 ;
        RECT 889.950 585.600 892.050 586.050 ;
        RECT 868.950 584.400 892.050 585.600 ;
        RECT 868.950 583.950 871.050 584.400 ;
        RECT 889.950 583.950 892.050 584.400 ;
        RECT 82.950 582.600 85.050 583.050 ;
        RECT 100.950 582.600 103.050 583.050 ;
        RECT 106.950 582.600 109.050 583.050 ;
        RECT 82.950 581.400 109.050 582.600 ;
        RECT 82.950 580.950 85.050 581.400 ;
        RECT 100.950 580.950 103.050 581.400 ;
        RECT 106.950 580.950 109.050 581.400 ;
        RECT 181.950 582.600 184.050 583.050 ;
        RECT 190.950 582.600 193.050 583.050 ;
        RECT 199.950 582.600 202.050 583.050 ;
        RECT 181.950 581.400 202.050 582.600 ;
        RECT 181.950 580.950 184.050 581.400 ;
        RECT 190.950 580.950 193.050 581.400 ;
        RECT 199.950 580.950 202.050 581.400 ;
        RECT 658.950 582.600 661.050 583.050 ;
        RECT 673.950 582.600 676.050 583.050 ;
        RECT 658.950 581.400 676.050 582.600 ;
        RECT 658.950 580.950 661.050 581.400 ;
        RECT 673.950 580.950 676.050 581.400 ;
        RECT 721.950 582.600 724.050 583.050 ;
        RECT 754.950 582.600 757.050 583.050 ;
        RECT 781.950 582.600 784.050 583.050 ;
        RECT 721.950 581.400 784.050 582.600 ;
        RECT 721.950 580.950 724.050 581.400 ;
        RECT 754.950 580.950 757.050 581.400 ;
        RECT 781.950 580.950 784.050 581.400 ;
        RECT 817.950 582.600 820.050 583.050 ;
        RECT 865.950 582.600 868.050 583.050 ;
        RECT 817.950 581.400 868.050 582.600 ;
        RECT 817.950 580.950 820.050 581.400 ;
        RECT 865.950 580.950 868.050 581.400 ;
        RECT 28.950 579.600 31.050 580.050 ;
        RECT 43.950 579.600 46.050 580.050 ;
        RECT 28.950 578.400 46.050 579.600 ;
        RECT 28.950 577.950 31.050 578.400 ;
        RECT 43.950 577.950 46.050 578.400 ;
        RECT 85.950 579.600 88.050 580.050 ;
        RECT 97.950 579.600 100.050 580.050 ;
        RECT 85.950 578.400 100.050 579.600 ;
        RECT 85.950 577.950 88.050 578.400 ;
        RECT 97.950 577.950 100.050 578.400 ;
        RECT 127.950 579.600 130.050 580.050 ;
        RECT 145.950 579.600 148.050 580.050 ;
        RECT 127.950 578.400 148.050 579.600 ;
        RECT 127.950 577.950 130.050 578.400 ;
        RECT 145.950 577.950 148.050 578.400 ;
        RECT 541.950 579.600 544.050 580.050 ;
        RECT 619.950 579.600 622.050 580.050 ;
        RECT 700.950 579.600 703.050 580.050 ;
        RECT 541.950 578.400 579.600 579.600 ;
        RECT 541.950 577.950 544.050 578.400 ;
        RECT 52.950 576.600 55.050 577.050 ;
        RECT 61.950 576.600 64.050 577.200 ;
        RECT 52.950 575.400 64.050 576.600 ;
        RECT 52.950 574.950 55.050 575.400 ;
        RECT 61.950 575.100 64.050 575.400 ;
        RECT 88.950 576.600 91.050 577.050 ;
        RECT 94.950 576.600 97.050 577.050 ;
        RECT 88.950 575.400 97.050 576.600 ;
        RECT 88.950 574.950 91.050 575.400 ;
        RECT 94.950 574.950 97.050 575.400 ;
        RECT 166.950 576.600 169.050 577.050 ;
        RECT 175.950 576.600 178.050 577.050 ;
        RECT 190.950 576.600 193.050 577.050 ;
        RECT 166.950 575.400 193.050 576.600 ;
        RECT 166.950 574.950 169.050 575.400 ;
        RECT 175.950 574.950 178.050 575.400 ;
        RECT 190.950 574.950 193.050 575.400 ;
        RECT 271.950 576.600 274.050 577.050 ;
        RECT 277.950 576.600 280.050 577.050 ;
        RECT 271.950 575.400 280.050 576.600 ;
        RECT 271.950 574.950 274.050 575.400 ;
        RECT 277.950 574.950 280.050 575.400 ;
        RECT 493.950 576.600 496.050 577.050 ;
        RECT 499.950 576.600 502.050 577.050 ;
        RECT 493.950 575.400 502.050 576.600 ;
        RECT 578.400 576.600 579.600 578.400 ;
        RECT 608.400 578.400 622.050 579.600 ;
        RECT 608.400 577.050 609.600 578.400 ;
        RECT 619.950 577.950 622.050 578.400 ;
        RECT 689.400 578.400 703.050 579.600 ;
        RECT 583.950 576.600 586.050 577.050 ;
        RECT 607.950 576.600 610.050 577.050 ;
        RECT 578.400 575.400 586.050 576.600 ;
        RECT 493.950 574.950 496.050 575.400 ;
        RECT 499.950 574.950 502.050 575.400 ;
        RECT 583.950 574.950 586.050 575.400 ;
        RECT 593.400 575.400 610.050 576.600 ;
        RECT 13.950 573.600 16.050 574.200 ;
        RECT 37.950 573.600 40.050 574.200 ;
        RECT 46.950 573.600 49.050 574.050 ;
        RECT 61.950 573.600 64.050 574.050 ;
        RECT 13.950 572.400 36.600 573.600 ;
        RECT 13.950 572.100 16.050 572.400 ;
        RECT 35.400 567.900 36.600 572.400 ;
        RECT 37.950 572.400 45.600 573.600 ;
        RECT 37.950 572.100 40.050 572.400 ;
        RECT 44.400 571.050 45.600 572.400 ;
        RECT 46.950 572.400 64.050 573.600 ;
        RECT 46.950 571.950 49.050 572.400 ;
        RECT 61.950 571.950 64.050 572.400 ;
        RECT 67.950 573.600 70.050 574.200 ;
        RECT 103.950 573.600 106.050 574.050 ;
        RECT 67.950 572.400 93.600 573.600 ;
        RECT 67.950 572.100 70.050 572.400 ;
        RECT 44.400 570.900 48.000 571.050 ;
        RECT 44.400 569.400 49.050 570.900 ;
        RECT 92.400 570.600 93.600 572.400 ;
        RECT 103.950 572.400 123.600 573.600 ;
        RECT 103.950 571.950 106.050 572.400 ;
        RECT 122.400 570.600 123.600 572.400 ;
        RECT 142.950 571.950 145.050 574.050 ;
        RECT 157.950 573.600 160.050 574.050 ;
        RECT 163.950 573.600 166.050 574.050 ;
        RECT 157.950 572.400 166.050 573.600 ;
        RECT 157.950 571.950 160.050 572.400 ;
        RECT 163.950 571.950 166.050 572.400 ;
        RECT 178.950 571.950 181.050 574.050 ;
        RECT 184.950 571.950 187.050 574.050 ;
        RECT 334.950 573.600 337.050 574.200 ;
        RECT 340.950 573.600 343.050 574.050 ;
        RECT 334.950 572.400 343.050 573.600 ;
        RECT 334.950 572.100 337.050 572.400 ;
        RECT 340.950 571.950 343.050 572.400 ;
        RECT 388.950 573.600 391.050 574.050 ;
        RECT 394.950 573.600 397.050 574.200 ;
        RECT 388.950 572.400 397.050 573.600 ;
        RECT 388.950 571.950 391.050 572.400 ;
        RECT 394.950 572.100 397.050 572.400 ;
        RECT 424.950 573.750 427.050 574.200 ;
        RECT 433.950 573.750 436.050 574.200 ;
        RECT 424.950 572.550 436.050 573.750 ;
        RECT 424.950 572.100 427.050 572.550 ;
        RECT 433.950 572.100 436.050 572.550 ;
        RECT 448.950 573.600 451.050 574.200 ;
        RECT 463.950 573.600 466.050 574.050 ;
        RECT 448.950 572.400 466.050 573.600 ;
        RECT 448.950 572.100 451.050 572.400 ;
        RECT 92.400 569.400 111.600 570.600 ;
        RECT 122.400 569.400 132.600 570.600 ;
        RECT 45.000 568.950 49.050 569.400 ;
        RECT 46.950 568.800 49.050 568.950 ;
        RECT 110.400 567.900 111.600 569.400 ;
        RECT 131.400 567.900 132.600 569.400 ;
        RECT 34.950 565.800 37.050 567.900 ;
        RECT 40.950 567.450 43.050 567.900 ;
        RECT 49.950 567.450 52.050 567.900 ;
        RECT 40.950 566.250 52.050 567.450 ;
        RECT 40.950 565.800 43.050 566.250 ;
        RECT 49.950 565.800 52.050 566.250 ;
        RECT 55.950 567.450 58.050 567.900 ;
        RECT 64.950 567.450 67.050 567.900 ;
        RECT 55.950 566.250 67.050 567.450 ;
        RECT 55.950 565.800 58.050 566.250 ;
        RECT 64.950 565.800 67.050 566.250 ;
        RECT 109.950 565.800 112.050 567.900 ;
        RECT 130.950 565.800 133.050 567.900 ;
        RECT 143.400 567.600 144.600 571.950 ;
        RECT 172.950 567.600 175.050 567.900 ;
        RECT 143.400 566.400 175.050 567.600 ;
        RECT 172.950 565.800 175.050 566.400 ;
        RECT 179.400 565.050 180.600 571.950 ;
        RECT 185.400 567.600 186.600 571.950 ;
        RECT 193.950 567.600 196.050 567.900 ;
        RECT 238.950 567.600 241.050 568.050 ;
        RECT 244.950 567.600 247.050 567.900 ;
        RECT 185.400 566.400 247.050 567.600 ;
        RECT 193.950 565.800 196.050 566.400 ;
        RECT 238.950 565.950 241.050 566.400 ;
        RECT 244.950 565.800 247.050 566.400 ;
        RECT 271.950 567.450 274.050 567.900 ;
        RECT 298.950 567.450 301.050 567.900 ;
        RECT 271.950 566.250 301.050 567.450 ;
        RECT 395.400 567.600 396.600 572.100 ;
        RECT 463.950 571.950 466.050 572.400 ;
        RECT 511.950 573.600 514.050 574.200 ;
        RECT 526.950 573.600 529.050 574.050 ;
        RECT 511.950 572.400 529.050 573.600 ;
        RECT 511.950 572.100 514.050 572.400 ;
        RECT 526.950 571.950 529.050 572.400 ;
        RECT 535.950 572.100 538.050 574.200 ;
        RECT 536.400 570.600 537.600 572.100 ;
        RECT 559.950 571.950 562.050 574.050 ;
        RECT 574.950 573.600 577.050 574.500 ;
        RECT 589.950 573.600 592.050 574.200 ;
        RECT 593.400 573.600 594.600 575.400 ;
        RECT 607.950 574.950 610.050 575.400 ;
        RECT 652.950 576.600 657.000 577.050 ;
        RECT 652.950 574.950 657.600 576.600 ;
        RECT 574.950 572.400 594.600 573.600 ;
        RECT 610.950 573.750 613.050 574.200 ;
        RECT 622.950 573.750 625.050 574.200 ;
        RECT 610.950 572.550 625.050 573.750 ;
        RECT 589.950 572.100 592.050 572.400 ;
        RECT 610.950 572.100 613.050 572.550 ;
        RECT 622.950 572.100 625.050 572.550 ;
        RECT 631.950 573.600 634.050 574.200 ;
        RECT 640.950 573.600 643.050 574.050 ;
        RECT 631.950 572.400 643.050 573.600 ;
        RECT 631.950 572.100 634.050 572.400 ;
        RECT 640.950 571.950 643.050 572.400 ;
        RECT 536.400 569.400 552.600 570.600 ;
        RECT 551.400 568.050 552.600 569.400 ;
        RECT 560.400 568.050 561.600 571.950 ;
        RECT 656.400 568.050 657.600 574.950 ;
        RECT 673.950 573.750 676.050 574.200 ;
        RECT 685.950 573.750 688.050 574.200 ;
        RECT 673.950 572.550 688.050 573.750 ;
        RECT 673.950 572.100 676.050 572.550 ;
        RECT 685.950 572.100 688.050 572.550 ;
        RECT 689.400 570.600 690.600 578.400 ;
        RECT 700.950 577.950 703.050 578.400 ;
        RECT 790.950 579.600 793.050 580.050 ;
        RECT 799.950 579.600 802.050 580.050 ;
        RECT 790.950 578.400 802.050 579.600 ;
        RECT 790.950 577.950 793.050 578.400 ;
        RECT 799.950 577.950 802.050 578.400 ;
        RECT 823.950 579.600 826.050 580.050 ;
        RECT 829.950 579.600 832.050 579.900 ;
        RECT 823.950 578.400 832.050 579.600 ;
        RECT 823.950 577.950 826.050 578.400 ;
        RECT 829.950 577.800 832.050 578.400 ;
        RECT 838.950 579.600 841.050 580.050 ;
        RECT 850.950 579.600 853.050 580.050 ;
        RECT 838.950 578.400 853.050 579.600 ;
        RECT 838.950 577.950 841.050 578.400 ;
        RECT 850.950 577.950 853.050 578.400 ;
        RECT 736.950 576.600 739.050 577.050 ;
        RECT 775.950 576.600 778.050 577.050 ;
        RECT 784.950 576.600 787.050 577.050 ;
        RECT 736.950 575.400 759.600 576.600 ;
        RECT 736.950 574.950 739.050 575.400 ;
        RECT 697.950 573.600 700.050 574.200 ;
        RECT 733.950 573.600 736.050 574.050 ;
        RECT 697.950 572.400 736.050 573.600 ;
        RECT 697.950 572.100 700.050 572.400 ;
        RECT 671.400 569.400 690.600 570.600 ;
        RECT 409.950 567.600 412.050 567.900 ;
        RECT 395.400 566.400 412.050 567.600 ;
        RECT 271.950 565.800 274.050 566.250 ;
        RECT 298.950 565.800 301.050 566.250 ;
        RECT 409.950 565.800 412.050 566.400 ;
        RECT 430.950 567.450 433.050 567.900 ;
        RECT 436.950 567.450 439.050 567.900 ;
        RECT 430.950 566.250 439.050 567.450 ;
        RECT 430.950 565.800 433.050 566.250 ;
        RECT 436.950 565.800 439.050 566.250 ;
        RECT 451.950 565.800 454.050 567.900 ;
        RECT 475.950 567.600 478.050 567.900 ;
        RECT 481.950 567.600 484.050 568.050 ;
        RECT 496.950 567.600 499.050 567.900 ;
        RECT 475.950 566.400 499.050 567.600 ;
        RECT 475.950 565.800 478.050 566.400 ;
        RECT 481.950 565.950 484.050 566.400 ;
        RECT 496.950 565.800 499.050 566.400 ;
        RECT 526.950 567.450 529.050 567.900 ;
        RECT 532.950 567.450 535.050 567.900 ;
        RECT 526.950 566.250 535.050 567.450 ;
        RECT 551.400 566.400 556.050 568.050 ;
        RECT 526.950 565.800 529.050 566.250 ;
        RECT 532.950 565.800 535.050 566.250 ;
        RECT 552.000 565.950 556.050 566.400 ;
        RECT 559.950 565.950 562.050 568.050 ;
        RECT 583.950 567.450 586.050 567.900 ;
        RECT 592.950 567.450 595.050 567.900 ;
        RECT 583.950 566.250 595.050 567.450 ;
        RECT 583.950 565.800 586.050 566.250 ;
        RECT 592.950 565.800 595.050 566.250 ;
        RECT 655.950 565.950 658.050 568.050 ;
        RECT 671.400 567.600 672.600 569.400 ;
        RECT 722.400 567.900 723.600 572.400 ;
        RECT 733.950 571.950 736.050 572.400 ;
        RECT 742.950 572.100 745.050 574.200 ;
        RECT 758.400 573.600 759.600 575.400 ;
        RECT 775.950 575.400 787.050 576.600 ;
        RECT 775.950 574.950 778.050 575.400 ;
        RECT 784.950 574.950 787.050 575.400 ;
        RECT 796.950 576.600 799.050 577.050 ;
        RECT 805.950 576.600 808.050 577.050 ;
        RECT 796.950 575.400 808.050 576.600 ;
        RECT 796.950 574.950 799.050 575.400 ;
        RECT 805.950 574.950 808.050 575.400 ;
        RECT 835.950 574.950 838.050 577.050 ;
        RECT 844.950 576.600 847.050 577.050 ;
        RECT 868.950 576.600 871.050 577.050 ;
        RECT 844.950 575.400 871.050 576.600 ;
        RECT 844.950 574.950 847.050 575.400 ;
        RECT 868.950 574.950 871.050 575.400 ;
        RECT 760.950 573.600 763.050 574.200 ;
        RECT 769.950 573.600 772.050 574.050 ;
        RECT 787.950 573.600 790.050 574.200 ;
        RECT 758.400 572.400 772.050 573.600 ;
        RECT 760.950 572.100 763.050 572.400 ;
        RECT 743.400 570.600 744.600 572.100 ;
        RECT 769.950 571.950 772.050 572.400 ;
        RECT 779.400 572.400 790.050 573.600 ;
        RECT 775.950 570.600 778.050 571.050 ;
        RECT 743.400 569.400 778.050 570.600 ;
        RECT 775.950 568.950 778.050 569.400 ;
        RECT 668.400 566.400 672.600 567.600 ;
        RECT 694.950 567.450 697.050 567.900 ;
        RECT 703.950 567.450 706.050 567.900 ;
        RECT 94.950 564.600 97.050 565.050 ;
        RECT 100.950 564.600 103.050 565.050 ;
        RECT 124.950 564.600 127.050 565.050 ;
        RECT 94.950 563.400 127.050 564.600 ;
        RECT 94.950 562.950 97.050 563.400 ;
        RECT 100.950 562.950 103.050 563.400 ;
        RECT 124.950 562.950 127.050 563.400 ;
        RECT 148.950 564.600 151.050 565.050 ;
        RECT 160.950 564.600 163.050 565.050 ;
        RECT 148.950 563.400 163.050 564.600 ;
        RECT 148.950 562.950 151.050 563.400 ;
        RECT 160.950 562.950 163.050 563.400 ;
        RECT 175.950 563.400 180.600 565.050 ;
        RECT 235.950 564.600 238.050 565.050 ;
        RECT 265.950 564.600 268.050 565.050 ;
        RECT 328.950 564.600 331.050 565.050 ;
        RECT 235.950 563.400 331.050 564.600 ;
        RECT 175.950 562.950 180.000 563.400 ;
        RECT 235.950 562.950 238.050 563.400 ;
        RECT 265.950 562.950 268.050 563.400 ;
        RECT 328.950 562.950 331.050 563.400 ;
        RECT 442.950 564.600 445.050 565.050 ;
        RECT 452.400 564.600 453.600 565.800 ;
        RECT 472.950 564.600 475.050 565.050 ;
        RECT 514.950 564.600 517.050 565.050 ;
        RECT 442.950 563.400 517.050 564.600 ;
        RECT 442.950 562.950 445.050 563.400 ;
        RECT 472.950 562.950 475.050 563.400 ;
        RECT 514.950 562.950 517.050 563.400 ;
        RECT 577.950 564.600 580.050 565.050 ;
        RECT 668.400 564.600 669.600 566.400 ;
        RECT 694.950 566.250 706.050 567.450 ;
        RECT 694.950 565.800 697.050 566.250 ;
        RECT 703.950 565.800 706.050 566.250 ;
        RECT 721.950 565.800 724.050 567.900 ;
        RECT 769.950 567.600 772.050 568.050 ;
        RECT 761.400 566.400 772.050 567.600 ;
        RECT 577.950 563.400 669.600 564.600 ;
        RECT 745.950 564.600 748.050 565.050 ;
        RECT 761.400 564.600 762.600 566.400 ;
        RECT 769.950 565.950 772.050 566.400 ;
        RECT 779.400 565.050 780.600 572.400 ;
        RECT 787.950 572.100 790.050 572.400 ;
        RECT 793.950 573.750 796.050 574.200 ;
        RECT 808.950 573.750 811.050 574.050 ;
        RECT 793.950 572.550 811.050 573.750 ;
        RECT 793.950 572.100 796.050 572.550 ;
        RECT 808.950 571.950 811.050 572.550 ;
        RECT 826.950 571.950 829.050 574.050 ;
        RECT 790.950 567.600 793.050 567.900 ;
        RECT 814.950 567.600 817.050 567.900 ;
        RECT 827.400 567.600 828.600 571.950 ;
        RECT 836.400 570.600 837.600 574.950 ;
        RECT 856.950 573.600 859.050 574.050 ;
        RECT 833.400 570.000 837.600 570.600 ;
        RECT 790.950 566.400 828.600 567.600 ;
        RECT 832.950 569.400 837.600 570.000 ;
        RECT 848.400 572.400 859.050 573.600 ;
        RECT 790.950 565.800 793.050 566.400 ;
        RECT 814.950 565.800 817.050 566.400 ;
        RECT 832.950 565.950 835.050 569.400 ;
        RECT 848.400 568.050 849.600 572.400 ;
        RECT 856.950 571.950 859.050 572.400 ;
        RECT 847.950 565.950 850.050 568.050 ;
        RECT 745.950 563.400 762.600 564.600 ;
        RECT 766.950 564.600 769.050 565.050 ;
        RECT 779.400 564.900 783.000 565.050 ;
        RECT 779.400 564.600 784.050 564.900 ;
        RECT 766.950 563.400 784.050 564.600 ;
        RECT 577.950 562.950 580.050 563.400 ;
        RECT 745.950 562.950 748.050 563.400 ;
        RECT 766.950 562.950 769.050 563.400 ;
        RECT 780.000 562.950 784.050 563.400 ;
        RECT 805.950 564.600 808.050 565.050 ;
        RECT 820.950 564.600 823.050 565.050 ;
        RECT 838.950 564.600 841.050 565.050 ;
        RECT 805.950 563.400 841.050 564.600 ;
        RECT 805.950 562.950 808.050 563.400 ;
        RECT 820.950 562.950 823.050 563.400 ;
        RECT 838.950 562.950 841.050 563.400 ;
        RECT 859.950 564.600 862.050 565.050 ;
        RECT 880.950 564.600 883.050 565.050 ;
        RECT 859.950 563.400 883.050 564.600 ;
        RECT 859.950 562.950 862.050 563.400 ;
        RECT 880.950 562.950 883.050 563.400 ;
        RECT 7.950 561.600 10.050 562.050 ;
        RECT 55.950 561.600 58.050 562.050 ;
        RECT 7.950 560.400 58.050 561.600 ;
        RECT 7.950 559.950 10.050 560.400 ;
        RECT 55.950 559.950 58.050 560.400 ;
        RECT 229.950 561.600 232.050 562.050 ;
        RECT 310.950 561.600 313.050 562.050 ;
        RECT 229.950 560.400 313.050 561.600 ;
        RECT 229.950 559.950 232.050 560.400 ;
        RECT 310.950 559.950 313.050 560.400 ;
        RECT 325.950 561.600 328.050 562.050 ;
        RECT 355.950 561.600 358.050 562.050 ;
        RECT 325.950 560.400 358.050 561.600 ;
        RECT 325.950 559.950 328.050 560.400 ;
        RECT 355.950 559.950 358.050 560.400 ;
        RECT 385.950 561.600 388.050 562.050 ;
        RECT 391.950 561.600 394.050 562.050 ;
        RECT 385.950 560.400 394.050 561.600 ;
        RECT 515.400 561.600 516.600 562.950 ;
        RECT 781.950 562.800 784.050 562.950 ;
        RECT 538.950 561.600 541.050 562.050 ;
        RECT 515.400 560.400 541.050 561.600 ;
        RECT 385.950 559.950 388.050 560.400 ;
        RECT 391.950 559.950 394.050 560.400 ;
        RECT 538.950 559.950 541.050 560.400 ;
        RECT 547.950 561.600 550.050 562.050 ;
        RECT 559.950 561.600 562.050 562.050 ;
        RECT 547.950 560.400 562.050 561.600 ;
        RECT 502.950 558.600 505.050 559.050 ;
        RECT 532.950 558.600 535.050 559.050 ;
        RECT 502.950 557.400 535.050 558.600 ;
        RECT 502.950 556.950 505.050 557.400 ;
        RECT 532.950 556.950 535.050 557.400 ;
        RECT 538.950 558.600 541.050 558.900 ;
        RECT 547.950 558.600 550.050 560.400 ;
        RECT 559.950 559.950 562.050 560.400 ;
        RECT 565.950 561.600 568.050 562.050 ;
        RECT 634.950 561.600 637.050 562.050 ;
        RECT 565.950 560.400 637.050 561.600 ;
        RECT 565.950 559.950 568.050 560.400 ;
        RECT 634.950 559.950 637.050 560.400 ;
        RECT 652.950 561.600 655.050 562.050 ;
        RECT 685.950 561.600 688.050 562.050 ;
        RECT 652.950 560.400 688.050 561.600 ;
        RECT 652.950 559.950 655.050 560.400 ;
        RECT 685.950 559.950 688.050 560.400 ;
        RECT 715.950 561.600 718.050 562.050 ;
        RECT 724.950 561.600 727.050 562.050 ;
        RECT 715.950 560.400 727.050 561.600 ;
        RECT 715.950 559.950 718.050 560.400 ;
        RECT 724.950 559.950 727.050 560.400 ;
        RECT 739.950 561.600 742.050 562.050 ;
        RECT 754.950 561.600 757.050 562.050 ;
        RECT 739.950 560.400 757.050 561.600 ;
        RECT 739.950 559.950 742.050 560.400 ;
        RECT 754.950 559.950 757.050 560.400 ;
        RECT 763.950 561.600 766.050 562.050 ;
        RECT 784.950 561.600 787.050 562.050 ;
        RECT 763.950 560.400 787.050 561.600 ;
        RECT 763.950 559.950 766.050 560.400 ;
        RECT 784.950 559.950 787.050 560.400 ;
        RECT 538.950 558.000 550.050 558.600 ;
        RECT 607.950 558.600 610.050 559.050 ;
        RECT 616.800 558.600 618.900 559.050 ;
        RECT 538.950 557.400 549.600 558.000 ;
        RECT 607.950 557.400 618.900 558.600 ;
        RECT 538.950 556.800 541.050 557.400 ;
        RECT 607.950 556.950 610.050 557.400 ;
        RECT 616.800 556.950 618.900 557.400 ;
        RECT 619.950 558.600 622.050 559.050 ;
        RECT 673.950 558.600 676.050 559.050 ;
        RECT 679.950 558.600 682.050 559.050 ;
        RECT 700.950 558.600 703.050 559.050 ;
        RECT 619.950 557.400 703.050 558.600 ;
        RECT 619.950 556.950 622.050 557.400 ;
        RECT 673.950 556.950 676.050 557.400 ;
        RECT 679.950 556.950 682.050 557.400 ;
        RECT 700.950 556.950 703.050 557.400 ;
        RECT 748.950 558.600 751.050 559.050 ;
        RECT 775.950 558.600 778.050 559.050 ;
        RECT 802.950 558.600 805.050 559.050 ;
        RECT 748.950 557.400 805.050 558.600 ;
        RECT 748.950 556.950 751.050 557.400 ;
        RECT 775.950 556.950 778.050 557.400 ;
        RECT 802.950 556.950 805.050 557.400 ;
        RECT 811.950 558.600 814.050 559.050 ;
        RECT 847.950 558.600 850.050 559.050 ;
        RECT 811.950 557.400 850.050 558.600 ;
        RECT 811.950 556.950 814.050 557.400 ;
        RECT 847.950 556.950 850.050 557.400 ;
        RECT 865.950 558.600 868.050 559.050 ;
        RECT 874.950 558.600 877.050 559.050 ;
        RECT 865.950 557.400 877.050 558.600 ;
        RECT 865.950 556.950 868.050 557.400 ;
        RECT 874.950 556.950 877.050 557.400 ;
        RECT 37.950 555.600 40.050 556.050 ;
        RECT 46.950 555.600 49.050 556.050 ;
        RECT 37.950 554.400 49.050 555.600 ;
        RECT 37.950 553.950 40.050 554.400 ;
        RECT 46.950 553.950 49.050 554.400 ;
        RECT 211.950 555.600 214.050 556.050 ;
        RECT 241.950 555.600 244.050 556.050 ;
        RECT 211.950 554.400 244.050 555.600 ;
        RECT 211.950 553.950 214.050 554.400 ;
        RECT 241.950 553.950 244.050 554.400 ;
        RECT 367.950 555.600 370.050 556.050 ;
        RECT 391.950 555.600 394.050 556.050 ;
        RECT 367.950 554.400 394.050 555.600 ;
        RECT 367.950 553.950 370.050 554.400 ;
        RECT 391.950 553.950 394.050 554.400 ;
        RECT 424.950 555.600 427.050 556.050 ;
        RECT 466.950 555.600 469.050 556.050 ;
        RECT 424.950 554.400 469.050 555.600 ;
        RECT 424.950 553.950 427.050 554.400 ;
        RECT 466.950 553.950 469.050 554.400 ;
        RECT 478.950 555.600 481.050 556.050 ;
        RECT 652.950 555.600 655.050 556.050 ;
        RECT 745.950 555.600 748.050 556.050 ;
        RECT 478.950 554.400 612.600 555.600 ;
        RECT 478.950 553.950 481.050 554.400 ;
        RECT 611.400 553.050 612.600 554.400 ;
        RECT 652.950 554.400 748.050 555.600 ;
        RECT 652.950 553.950 655.050 554.400 ;
        RECT 745.950 553.950 748.050 554.400 ;
        RECT 835.950 555.600 838.050 556.050 ;
        RECT 844.950 555.600 847.050 556.050 ;
        RECT 835.950 554.400 847.050 555.600 ;
        RECT 835.950 553.950 838.050 554.400 ;
        RECT 844.950 553.950 847.050 554.400 ;
        RECT 502.950 552.600 505.050 553.050 ;
        RECT 520.800 552.600 522.900 553.050 ;
        RECT 502.950 551.400 522.900 552.600 ;
        RECT 502.950 550.950 505.050 551.400 ;
        RECT 520.800 550.950 522.900 551.400 ;
        RECT 610.950 552.600 613.050 553.050 ;
        RECT 631.950 552.600 634.050 553.050 ;
        RECT 748.950 552.600 751.050 553.050 ;
        RECT 610.950 551.400 751.050 552.600 ;
        RECT 610.950 550.950 613.050 551.400 ;
        RECT 631.950 550.950 634.050 551.400 ;
        RECT 748.950 550.950 751.050 551.400 ;
        RECT 754.950 552.600 757.050 553.050 ;
        RECT 766.950 552.600 769.050 553.050 ;
        RECT 754.950 551.400 769.050 552.600 ;
        RECT 754.950 550.950 757.050 551.400 ;
        RECT 766.950 550.950 769.050 551.400 ;
        RECT 787.950 552.600 790.050 553.050 ;
        RECT 808.950 552.600 811.050 553.050 ;
        RECT 787.950 551.400 811.050 552.600 ;
        RECT 787.950 550.950 790.050 551.400 ;
        RECT 808.950 550.950 811.050 551.400 ;
        RECT 52.950 549.600 55.050 549.900 ;
        RECT 115.950 549.600 118.050 550.050 ;
        RECT 52.950 548.400 118.050 549.600 ;
        RECT 52.950 547.800 55.050 548.400 ;
        RECT 115.950 547.950 118.050 548.400 ;
        RECT 163.950 549.600 166.050 550.050 ;
        RECT 178.950 549.600 181.050 550.050 ;
        RECT 163.950 548.400 181.050 549.600 ;
        RECT 163.950 547.950 166.050 548.400 ;
        RECT 178.950 547.950 181.050 548.400 ;
        RECT 187.950 549.600 190.050 550.050 ;
        RECT 196.950 549.600 199.050 550.050 ;
        RECT 187.950 548.400 199.050 549.600 ;
        RECT 187.950 547.950 190.050 548.400 ;
        RECT 196.950 547.950 199.050 548.400 ;
        RECT 250.950 549.600 253.050 550.050 ;
        RECT 259.950 549.600 262.050 550.050 ;
        RECT 250.950 548.400 262.050 549.600 ;
        RECT 250.950 547.950 253.050 548.400 ;
        RECT 259.950 547.950 262.050 548.400 ;
        RECT 388.950 549.600 391.050 550.050 ;
        RECT 442.950 549.600 445.050 550.050 ;
        RECT 388.950 548.400 445.050 549.600 ;
        RECT 388.950 547.950 391.050 548.400 ;
        RECT 442.950 547.950 445.050 548.400 ;
        RECT 622.950 549.600 625.050 550.050 ;
        RECT 664.950 549.600 667.050 550.050 ;
        RECT 670.950 549.600 673.050 550.050 ;
        RECT 622.950 548.400 673.050 549.600 ;
        RECT 622.950 547.950 625.050 548.400 ;
        RECT 664.950 547.950 667.050 548.400 ;
        RECT 670.950 547.950 673.050 548.400 ;
        RECT 679.950 549.600 682.050 550.050 ;
        RECT 715.950 549.600 718.050 550.050 ;
        RECT 679.950 548.400 718.050 549.600 ;
        RECT 679.950 547.950 682.050 548.400 ;
        RECT 715.950 547.950 718.050 548.400 ;
        RECT 742.950 549.600 745.050 550.050 ;
        RECT 766.950 549.600 769.050 549.900 ;
        RECT 742.950 548.400 769.050 549.600 ;
        RECT 742.950 547.950 745.050 548.400 ;
        RECT 766.950 547.800 769.050 548.400 ;
        RECT 850.950 549.600 853.050 550.050 ;
        RECT 883.950 549.600 886.050 550.050 ;
        RECT 850.950 548.400 886.050 549.600 ;
        RECT 850.950 547.950 853.050 548.400 ;
        RECT 883.950 547.950 886.050 548.400 ;
        RECT 460.950 546.600 463.050 547.050 ;
        RECT 712.950 546.600 715.050 547.050 ;
        RECT 460.950 545.400 715.050 546.600 ;
        RECT 460.950 544.950 463.050 545.400 ;
        RECT 712.950 544.950 715.050 545.400 ;
        RECT 763.950 546.600 766.050 547.050 ;
        RECT 772.950 546.600 775.050 547.050 ;
        RECT 763.950 545.400 775.050 546.600 ;
        RECT 763.950 544.950 766.050 545.400 ;
        RECT 772.950 544.950 775.050 545.400 ;
        RECT 781.950 546.600 784.050 547.050 ;
        RECT 808.950 546.600 811.050 547.050 ;
        RECT 781.950 545.400 811.050 546.600 ;
        RECT 781.950 544.950 784.050 545.400 ;
        RECT 808.950 544.950 811.050 545.400 ;
        RECT 820.950 546.600 823.050 547.050 ;
        RECT 853.950 546.600 856.050 547.050 ;
        RECT 820.950 545.400 856.050 546.600 ;
        RECT 820.950 544.950 823.050 545.400 ;
        RECT 853.950 544.950 856.050 545.400 ;
        RECT 4.950 543.600 7.050 544.050 ;
        RECT 82.950 543.600 85.050 544.050 ;
        RECT 4.950 542.400 85.050 543.600 ;
        RECT 4.950 541.950 7.050 542.400 ;
        RECT 82.950 541.950 85.050 542.400 ;
        RECT 97.950 543.600 100.050 544.050 ;
        RECT 112.950 543.600 115.050 544.050 ;
        RECT 97.950 542.400 115.050 543.600 ;
        RECT 97.950 541.950 100.050 542.400 ;
        RECT 112.950 541.950 115.050 542.400 ;
        RECT 175.950 543.600 178.050 544.050 ;
        RECT 211.950 543.600 214.050 544.050 ;
        RECT 175.950 542.400 214.050 543.600 ;
        RECT 175.950 541.950 178.050 542.400 ;
        RECT 211.950 541.950 214.050 542.400 ;
        RECT 391.950 543.600 394.050 544.050 ;
        RECT 439.950 543.600 442.050 544.050 ;
        RECT 391.950 542.400 442.050 543.600 ;
        RECT 391.950 541.950 394.050 542.400 ;
        RECT 439.950 541.950 442.050 542.400 ;
        RECT 463.950 543.600 466.050 544.050 ;
        RECT 469.950 543.600 472.050 544.050 ;
        RECT 463.950 542.400 472.050 543.600 ;
        RECT 463.950 541.950 466.050 542.400 ;
        RECT 469.950 541.950 472.050 542.400 ;
        RECT 484.950 543.600 487.050 544.050 ;
        RECT 496.950 543.600 499.050 544.050 ;
        RECT 484.950 542.400 499.050 543.600 ;
        RECT 484.950 541.950 487.050 542.400 ;
        RECT 496.950 541.950 499.050 542.400 ;
        RECT 730.950 543.600 733.050 544.050 ;
        RECT 736.950 543.600 739.050 544.050 ;
        RECT 754.950 543.600 757.050 544.050 ;
        RECT 730.950 542.400 757.050 543.600 ;
        RECT 730.950 541.950 733.050 542.400 ;
        RECT 736.950 541.950 739.050 542.400 ;
        RECT 754.950 541.950 757.050 542.400 ;
        RECT 790.950 543.600 793.050 544.050 ;
        RECT 811.950 543.600 814.050 544.050 ;
        RECT 790.950 542.400 814.050 543.600 ;
        RECT 790.950 541.950 793.050 542.400 ;
        RECT 811.950 541.950 814.050 542.400 ;
        RECT 25.950 540.600 28.050 541.050 ;
        RECT 76.950 540.600 79.050 541.050 ;
        RECT 25.950 539.400 79.050 540.600 ;
        RECT 25.950 538.950 28.050 539.400 ;
        RECT 76.950 538.950 79.050 539.400 ;
        RECT 145.950 540.600 148.050 541.050 ;
        RECT 235.950 540.600 238.050 541.050 ;
        RECT 145.950 539.400 238.050 540.600 ;
        RECT 145.950 538.950 148.050 539.400 ;
        RECT 235.950 538.950 238.050 539.400 ;
        RECT 280.950 540.600 283.050 541.050 ;
        RECT 313.950 540.600 316.050 541.050 ;
        RECT 388.950 540.600 391.050 541.050 ;
        RECT 280.950 539.400 391.050 540.600 ;
        RECT 280.950 538.950 283.050 539.400 ;
        RECT 313.950 538.950 316.050 539.400 ;
        RECT 388.950 538.950 391.050 539.400 ;
        RECT 466.950 540.600 469.050 541.050 ;
        RECT 481.950 540.600 484.050 541.050 ;
        RECT 466.950 539.400 484.050 540.600 ;
        RECT 466.950 538.950 469.050 539.400 ;
        RECT 481.950 538.950 484.050 539.400 ;
        RECT 532.950 540.600 535.050 541.050 ;
        RECT 577.950 540.600 580.050 541.050 ;
        RECT 532.950 539.400 580.050 540.600 ;
        RECT 532.950 538.950 535.050 539.400 ;
        RECT 577.950 538.950 580.050 539.400 ;
        RECT 685.950 540.600 688.050 541.050 ;
        RECT 760.950 540.600 763.050 541.050 ;
        RECT 772.950 540.600 775.050 541.050 ;
        RECT 787.950 540.600 790.050 541.050 ;
        RECT 685.950 539.400 790.050 540.600 ;
        RECT 685.950 538.950 688.050 539.400 ;
        RECT 760.950 538.950 763.050 539.400 ;
        RECT 772.950 538.950 775.050 539.400 ;
        RECT 787.950 538.950 790.050 539.400 ;
        RECT 823.950 540.600 826.050 541.050 ;
        RECT 877.950 540.600 880.050 541.050 ;
        RECT 823.950 539.400 880.050 540.600 ;
        RECT 823.950 538.950 826.050 539.400 ;
        RECT 877.950 538.950 880.050 539.400 ;
        RECT 88.950 537.600 91.050 538.050 ;
        RECT 68.400 536.400 91.050 537.600 ;
        RECT 16.950 531.600 19.050 532.050 ;
        RECT 11.400 530.400 19.050 531.600 ;
        RECT 11.400 522.900 12.600 530.400 ;
        RECT 16.950 529.950 19.050 530.400 ;
        RECT 13.950 527.100 16.050 529.200 ;
        RECT 19.950 528.750 22.050 529.200 ;
        RECT 25.950 528.750 28.050 529.200 ;
        RECT 19.950 527.550 28.050 528.750 ;
        RECT 19.950 527.100 22.050 527.550 ;
        RECT 25.950 527.100 28.050 527.550 ;
        RECT 10.950 520.800 13.050 522.900 ;
        RECT 14.400 522.600 15.600 527.100 ;
        RECT 40.950 522.600 43.050 522.900 ;
        RECT 14.400 521.400 43.050 522.600 ;
        RECT 40.950 520.800 43.050 521.400 ;
        RECT 68.400 517.050 69.600 536.400 ;
        RECT 88.950 535.950 91.050 536.400 ;
        RECT 109.950 537.600 112.050 538.050 ;
        RECT 124.950 537.600 127.050 538.050 ;
        RECT 109.950 536.400 127.050 537.600 ;
        RECT 109.950 535.950 112.050 536.400 ;
        RECT 124.950 535.950 127.050 536.400 ;
        RECT 136.950 537.600 139.050 538.050 ;
        RECT 193.950 537.600 196.050 538.050 ;
        RECT 136.950 536.400 196.050 537.600 ;
        RECT 136.950 535.950 139.050 536.400 ;
        RECT 193.950 535.950 196.050 536.400 ;
        RECT 262.950 537.600 265.050 538.050 ;
        RECT 277.950 537.600 280.050 538.050 ;
        RECT 262.950 536.400 280.050 537.600 ;
        RECT 262.950 535.950 265.050 536.400 ;
        RECT 277.950 535.950 280.050 536.400 ;
        RECT 334.950 537.600 337.050 538.050 ;
        RECT 340.950 537.600 343.050 538.050 ;
        RECT 334.950 536.400 343.050 537.600 ;
        RECT 334.950 535.950 337.050 536.400 ;
        RECT 340.950 535.950 343.050 536.400 ;
        RECT 358.950 537.600 361.050 538.050 ;
        RECT 373.950 537.600 376.050 538.050 ;
        RECT 400.950 537.600 403.050 538.050 ;
        RECT 430.950 537.600 433.050 538.050 ;
        RECT 358.950 536.400 387.600 537.600 ;
        RECT 358.950 535.950 361.050 536.400 ;
        RECT 373.950 535.950 376.050 536.400 ;
        RECT 91.950 534.600 94.050 535.050 ;
        RECT 71.400 533.400 94.050 534.600 ;
        RECT 71.400 520.050 72.600 533.400 ;
        RECT 91.950 532.950 94.050 533.400 ;
        RECT 109.950 534.600 112.050 534.900 ;
        RECT 178.950 534.600 181.050 535.050 ;
        RECT 187.950 534.600 190.050 535.050 ;
        RECT 109.950 533.400 190.050 534.600 ;
        RECT 109.950 532.800 112.050 533.400 ;
        RECT 178.950 532.950 181.050 533.400 ;
        RECT 187.950 532.950 190.050 533.400 ;
        RECT 205.950 534.600 208.050 535.050 ;
        RECT 223.950 534.600 226.050 535.050 ;
        RECT 205.950 533.400 226.050 534.600 ;
        RECT 205.950 532.950 208.050 533.400 ;
        RECT 223.950 532.950 226.050 533.400 ;
        RECT 274.950 534.600 277.050 535.050 ;
        RECT 304.950 534.600 307.050 535.050 ;
        RECT 274.950 533.400 307.050 534.600 ;
        RECT 274.950 532.950 277.050 533.400 ;
        RECT 304.950 532.950 307.050 533.400 ;
        RECT 310.950 534.600 313.050 535.050 ;
        RECT 349.950 534.600 352.050 535.050 ;
        RECT 310.950 533.400 352.050 534.600 ;
        RECT 386.400 534.600 387.600 536.400 ;
        RECT 400.950 536.400 433.050 537.600 ;
        RECT 400.950 535.950 403.050 536.400 ;
        RECT 430.950 535.950 433.050 536.400 ;
        RECT 457.950 537.600 460.050 538.050 ;
        RECT 493.950 537.600 496.050 538.050 ;
        RECT 457.950 536.400 496.050 537.600 ;
        RECT 457.950 535.950 460.050 536.400 ;
        RECT 493.950 535.950 496.050 536.400 ;
        RECT 505.950 537.600 508.050 538.050 ;
        RECT 520.950 537.600 523.050 538.050 ;
        RECT 505.950 536.400 523.050 537.600 ;
        RECT 505.950 535.950 508.050 536.400 ;
        RECT 520.950 535.950 523.050 536.400 ;
        RECT 700.950 537.600 703.050 538.050 ;
        RECT 757.950 537.600 760.050 538.050 ;
        RECT 700.950 536.400 760.050 537.600 ;
        RECT 700.950 535.950 703.050 536.400 ;
        RECT 757.950 535.950 760.050 536.400 ;
        RECT 766.950 537.600 769.050 538.050 ;
        RECT 790.950 537.600 793.050 538.050 ;
        RECT 766.950 536.400 793.050 537.600 ;
        RECT 766.950 535.950 769.050 536.400 ;
        RECT 790.950 535.950 793.050 536.400 ;
        RECT 421.950 534.600 424.050 535.050 ;
        RECT 386.400 533.400 424.050 534.600 ;
        RECT 310.950 532.950 313.050 533.400 ;
        RECT 349.950 532.950 352.050 533.400 ;
        RECT 421.950 532.950 424.050 533.400 ;
        RECT 475.950 534.600 478.050 535.050 ;
        RECT 517.950 534.600 520.050 535.050 ;
        RECT 475.950 533.400 520.050 534.600 ;
        RECT 475.950 532.950 478.050 533.400 ;
        RECT 517.950 532.950 520.050 533.400 ;
        RECT 523.950 534.600 526.050 535.050 ;
        RECT 532.950 534.600 535.050 535.050 ;
        RECT 523.950 533.400 535.050 534.600 ;
        RECT 523.950 532.950 526.050 533.400 ;
        RECT 532.950 532.950 535.050 533.400 ;
        RECT 625.950 534.600 628.050 535.050 ;
        RECT 640.950 534.600 643.050 535.050 ;
        RECT 625.950 533.400 643.050 534.600 ;
        RECT 625.950 532.950 628.050 533.400 ;
        RECT 640.950 532.950 643.050 533.400 ;
        RECT 793.950 534.600 796.050 535.050 ;
        RECT 811.950 534.600 814.050 535.050 ;
        RECT 793.950 533.400 814.050 534.600 ;
        RECT 793.950 532.950 796.050 533.400 ;
        RECT 811.950 532.950 814.050 533.400 ;
        RECT 829.950 534.600 832.050 535.050 ;
        RECT 847.950 534.600 850.050 535.050 ;
        RECT 829.950 533.400 850.050 534.600 ;
        RECT 829.950 532.950 832.050 533.400 ;
        RECT 847.950 532.950 850.050 533.400 ;
        RECT 862.950 534.600 865.050 535.050 ;
        RECT 877.950 534.600 880.050 535.050 ;
        RECT 862.950 533.400 880.050 534.600 ;
        RECT 862.950 532.950 865.050 533.400 ;
        RECT 877.950 532.950 880.050 533.400 ;
        RECT 76.950 528.600 79.050 529.050 ;
        RECT 88.950 528.600 91.050 529.050 ;
        RECT 93.000 528.600 97.050 529.050 ;
        RECT 74.400 528.000 91.050 528.600 ;
        RECT 73.950 527.400 91.050 528.000 ;
        RECT 73.950 523.800 76.050 527.400 ;
        RECT 76.950 526.950 79.050 527.400 ;
        RECT 88.950 526.950 91.050 527.400 ;
        RECT 92.400 526.950 97.050 528.600 ;
        RECT 100.950 528.600 103.050 529.050 ;
        RECT 115.950 528.600 118.050 529.050 ;
        RECT 145.950 528.600 148.050 529.200 ;
        RECT 100.950 527.400 118.050 528.600 ;
        RECT 100.950 526.950 103.050 527.400 ;
        RECT 115.950 526.950 118.050 527.400 ;
        RECT 122.400 527.400 148.050 528.600 ;
        RECT 92.400 525.600 93.600 526.950 ;
        RECT 80.400 524.400 93.600 525.600 ;
        RECT 80.400 522.600 81.600 524.400 ;
        RECT 122.400 522.900 123.600 527.400 ;
        RECT 145.950 527.100 148.050 527.400 ;
        RECT 151.950 528.750 154.050 529.200 ;
        RECT 169.800 528.750 171.900 529.200 ;
        RECT 151.950 527.550 171.900 528.750 ;
        RECT 151.950 527.100 154.050 527.550 ;
        RECT 169.800 527.100 171.900 527.550 ;
        RECT 172.950 528.600 175.050 529.050 ;
        RECT 178.950 528.600 181.050 529.500 ;
        RECT 172.950 527.400 181.050 528.600 ;
        RECT 220.950 528.600 223.050 532.050 ;
        RECT 229.950 531.600 232.050 532.050 ;
        RECT 235.950 531.600 238.050 532.050 ;
        RECT 229.950 530.400 238.050 531.600 ;
        RECT 229.950 529.950 232.050 530.400 ;
        RECT 235.950 529.950 238.050 530.400 ;
        RECT 382.950 531.600 385.050 532.050 ;
        RECT 406.950 531.600 409.050 532.050 ;
        RECT 382.950 530.400 409.050 531.600 ;
        RECT 382.950 529.950 385.050 530.400 ;
        RECT 406.950 529.950 409.050 530.400 ;
        RECT 454.950 531.600 457.050 531.900 ;
        RECT 469.950 531.600 472.050 532.050 ;
        RECT 454.950 530.400 472.050 531.600 ;
        RECT 454.950 529.800 457.050 530.400 ;
        RECT 469.950 529.950 472.050 530.400 ;
        RECT 601.950 531.600 604.050 531.900 ;
        RECT 658.950 531.600 661.050 532.050 ;
        RECT 601.950 530.400 661.050 531.600 ;
        RECT 601.950 529.800 604.050 530.400 ;
        RECT 658.950 529.950 661.050 530.400 ;
        RECT 682.950 529.950 685.050 532.050 ;
        RECT 739.950 531.600 742.050 532.050 ;
        RECT 751.950 531.600 754.050 532.050 ;
        RECT 739.950 530.400 754.050 531.600 ;
        RECT 739.950 529.950 742.050 530.400 ;
        RECT 751.950 529.950 754.050 530.400 ;
        RECT 238.950 528.600 241.050 529.050 ;
        RECT 253.950 528.600 256.050 529.200 ;
        RECT 268.950 528.600 271.050 529.200 ;
        RECT 220.950 528.000 228.600 528.600 ;
        RECT 221.400 527.400 228.600 528.000 ;
        RECT 172.950 526.950 175.050 527.400 ;
        RECT 79.950 520.500 82.050 522.600 ;
        RECT 121.950 520.800 124.050 522.900 ;
        RECT 136.950 522.600 139.050 523.050 ;
        RECT 227.400 522.900 228.600 527.400 ;
        RECT 238.950 527.400 271.050 528.600 ;
        RECT 238.950 526.950 241.050 527.400 ;
        RECT 253.950 527.100 256.050 527.400 ;
        RECT 268.950 527.100 271.050 527.400 ;
        RECT 292.950 528.600 295.050 529.200 ;
        RECT 292.950 527.400 330.600 528.600 ;
        RECT 340.950 527.400 343.050 529.500 ;
        RECT 373.950 528.750 376.050 529.200 ;
        RECT 379.950 528.750 382.050 529.200 ;
        RECT 373.950 527.550 382.050 528.750 ;
        RECT 292.950 527.100 295.050 527.400 ;
        RECT 329.400 526.050 330.600 527.400 ;
        RECT 329.400 524.400 334.050 526.050 ;
        RECT 330.000 523.950 334.050 524.400 ;
        RECT 341.400 523.050 342.600 527.400 ;
        RECT 373.950 527.100 376.050 527.550 ;
        RECT 379.950 527.100 382.050 527.550 ;
        RECT 412.950 527.100 415.050 529.200 ;
        RECT 397.950 525.600 400.050 526.050 ;
        RECT 413.400 525.600 414.600 527.100 ;
        RECT 472.950 526.950 475.050 529.050 ;
        RECT 481.950 528.750 484.050 529.200 ;
        RECT 487.950 528.750 490.050 529.200 ;
        RECT 481.950 527.550 490.050 528.750 ;
        RECT 481.950 527.100 484.050 527.550 ;
        RECT 487.950 527.100 490.050 527.550 ;
        RECT 493.950 528.600 496.050 529.050 ;
        RECT 499.950 528.600 502.050 529.050 ;
        RECT 493.950 527.400 502.050 528.600 ;
        RECT 493.950 526.950 496.050 527.400 ;
        RECT 499.950 526.950 502.050 527.400 ;
        RECT 505.950 528.600 508.050 529.050 ;
        RECT 505.950 527.400 513.600 528.600 ;
        RECT 523.950 527.400 526.050 529.500 ;
        RECT 559.950 528.600 562.050 529.050 ;
        RECT 568.950 528.600 571.050 529.200 ;
        RECT 559.950 527.400 571.050 528.600 ;
        RECT 505.950 526.950 508.050 527.400 ;
        RECT 397.950 524.400 414.600 525.600 ;
        RECT 397.950 523.950 400.050 524.400 ;
        RECT 148.950 522.600 151.050 522.900 ;
        RECT 136.950 521.400 151.050 522.600 ;
        RECT 136.950 520.950 139.050 521.400 ;
        RECT 148.950 520.800 151.050 521.400 ;
        RECT 196.950 522.450 199.050 522.900 ;
        RECT 202.950 522.450 205.050 522.900 ;
        RECT 196.950 521.250 205.050 522.450 ;
        RECT 196.950 520.800 199.050 521.250 ;
        RECT 202.950 520.800 205.050 521.250 ;
        RECT 226.950 520.800 229.050 522.900 ;
        RECT 250.950 522.600 253.050 523.050 ;
        RECT 283.950 522.600 286.050 523.050 ;
        RECT 250.950 521.400 286.050 522.600 ;
        RECT 250.950 520.950 253.050 521.400 ;
        RECT 283.950 520.950 286.050 521.400 ;
        RECT 337.950 521.400 342.600 523.050 ;
        RECT 400.950 522.600 403.050 523.050 ;
        RECT 409.950 522.600 412.050 522.900 ;
        RECT 400.950 521.400 412.050 522.600 ;
        RECT 413.400 522.600 414.600 524.400 ;
        RECT 473.400 523.050 474.600 526.950 ;
        RECT 418.950 522.600 421.050 523.050 ;
        RECT 457.950 522.600 460.050 523.050 ;
        RECT 466.950 522.600 469.050 522.900 ;
        RECT 413.400 521.400 421.050 522.600 ;
        RECT 337.950 520.950 342.000 521.400 ;
        RECT 400.950 520.950 403.050 521.400 ;
        RECT 409.950 520.800 412.050 521.400 ;
        RECT 418.950 520.950 421.050 521.400 ;
        RECT 439.950 522.150 442.050 522.600 ;
        RECT 448.950 522.150 451.050 522.600 ;
        RECT 439.950 520.950 451.050 522.150 ;
        RECT 457.950 521.400 469.050 522.600 ;
        RECT 457.950 520.950 460.050 521.400 ;
        RECT 439.950 520.500 442.050 520.950 ;
        RECT 448.950 520.500 451.050 520.950 ;
        RECT 466.950 520.800 469.050 521.400 ;
        RECT 472.950 520.950 475.050 523.050 ;
        RECT 512.400 522.900 513.600 527.400 ;
        RECT 524.400 525.600 525.600 527.400 ;
        RECT 559.950 526.950 562.050 527.400 ;
        RECT 568.950 527.100 571.050 527.400 ;
        RECT 619.950 527.100 622.050 529.200 ;
        RECT 625.950 528.600 628.050 529.200 ;
        RECT 640.950 528.600 643.050 529.200 ;
        RECT 646.950 528.600 649.050 529.050 ;
        RECT 655.950 528.600 658.050 529.050 ;
        RECT 625.950 527.400 639.600 528.600 ;
        RECT 625.950 527.100 628.050 527.400 ;
        RECT 538.950 525.600 541.050 526.050 ;
        RECT 620.400 525.600 621.600 527.100 ;
        RECT 524.400 524.400 541.050 525.600 ;
        RECT 538.950 523.950 541.050 524.400 ;
        RECT 593.400 524.400 621.600 525.600 ;
        RECT 511.950 520.800 514.050 522.900 ;
        RECT 517.950 522.450 520.050 522.900 ;
        RECT 538.950 522.450 541.050 522.900 ;
        RECT 571.950 522.600 574.050 522.900 ;
        RECT 593.400 522.600 594.600 524.400 ;
        RECT 638.400 522.900 639.600 527.400 ;
        RECT 640.950 527.400 649.050 528.600 ;
        RECT 640.950 527.100 643.050 527.400 ;
        RECT 646.950 526.950 649.050 527.400 ;
        RECT 650.400 527.400 658.050 528.600 ;
        RECT 517.950 521.250 541.050 522.450 ;
        RECT 517.950 520.800 520.050 521.250 ;
        RECT 538.950 520.800 541.050 521.250 ;
        RECT 550.950 522.150 553.050 522.600 ;
        RECT 556.950 522.150 559.050 522.600 ;
        RECT 550.950 520.950 559.050 522.150 ;
        RECT 550.950 520.500 553.050 520.950 ;
        RECT 556.950 520.500 559.050 520.950 ;
        RECT 571.950 521.400 594.600 522.600 ;
        RECT 571.950 520.800 574.050 521.400 ;
        RECT 637.950 520.800 640.050 522.900 ;
        RECT 643.950 522.600 646.050 523.050 ;
        RECT 650.400 522.600 651.600 527.400 ;
        RECT 655.950 526.950 658.050 527.400 ;
        RECT 664.950 527.100 667.050 529.200 ;
        RECT 643.950 521.400 651.600 522.600 ;
        RECT 643.950 520.950 646.050 521.400 ;
        RECT 665.400 520.050 666.600 527.100 ;
        RECT 673.950 526.950 676.050 529.050 ;
        RECT 674.400 523.050 675.600 526.950 ;
        RECT 673.950 520.950 676.050 523.050 ;
        RECT 683.400 522.900 684.600 529.950 ;
        RECT 706.950 528.600 709.050 529.200 ;
        RECT 706.950 527.400 717.600 528.600 ;
        RECT 706.950 527.100 709.050 527.400 ;
        RECT 716.400 523.050 717.600 527.400 ;
        RECT 742.950 526.950 745.050 529.050 ;
        RECT 766.950 528.750 769.050 529.200 ;
        RECT 793.950 528.750 796.050 529.200 ;
        RECT 766.950 527.550 796.050 528.750 ;
        RECT 766.950 527.100 769.050 527.550 ;
        RECT 793.950 527.100 796.050 527.550 ;
        RECT 799.950 527.100 802.050 529.200 ;
        RECT 808.950 528.600 811.050 529.050 ;
        RECT 808.950 527.400 816.600 528.600 ;
        RECT 743.400 523.050 744.600 526.950 ;
        RECT 800.400 523.050 801.600 527.100 ;
        RECT 808.950 526.950 811.050 527.400 ;
        RECT 815.400 523.050 816.600 527.400 ;
        RECT 823.950 526.950 826.050 529.050 ;
        RECT 835.950 526.950 838.050 529.050 ;
        RECT 841.950 527.100 844.050 529.200 ;
        RECT 853.950 528.750 856.050 529.200 ;
        RECT 868.950 528.750 871.050 529.200 ;
        RECT 853.950 528.600 871.050 528.750 ;
        RECT 895.950 528.600 898.050 529.050 ;
        RECT 853.950 527.550 898.050 528.600 ;
        RECT 853.950 527.100 856.050 527.550 ;
        RECT 868.950 527.400 898.050 527.550 ;
        RECT 868.950 527.100 871.050 527.400 ;
        RECT 824.400 523.050 825.600 526.950 ;
        RECT 836.400 523.050 837.600 526.950 ;
        RECT 842.400 525.600 843.600 527.100 ;
        RECT 895.950 526.950 898.050 527.400 ;
        RECT 842.400 524.400 867.600 525.600 ;
        RECT 682.950 520.800 685.050 522.900 ;
        RECT 716.400 521.400 721.050 523.050 ;
        RECT 717.000 520.950 721.050 521.400 ;
        RECT 742.950 520.950 745.050 523.050 ;
        RECT 775.950 522.450 778.050 522.900 ;
        RECT 784.950 522.450 787.050 523.050 ;
        RECT 790.950 522.450 793.050 522.900 ;
        RECT 775.950 521.250 793.050 522.450 ;
        RECT 800.400 521.400 805.050 523.050 ;
        RECT 775.950 520.800 778.050 521.250 ;
        RECT 784.950 520.950 787.050 521.250 ;
        RECT 790.950 520.800 793.050 521.250 ;
        RECT 801.000 520.950 805.050 521.400 ;
        RECT 814.950 520.950 817.050 523.050 ;
        RECT 823.950 520.950 826.050 523.050 ;
        RECT 835.950 520.950 838.050 523.050 ;
        RECT 866.400 520.050 867.600 524.400 ;
        RECT 71.400 519.900 75.000 520.050 ;
        RECT 71.400 518.400 76.050 519.900 ;
        RECT 72.000 517.950 76.050 518.400 ;
        RECT 241.950 519.600 244.050 520.050 ;
        RECT 247.950 519.600 250.050 520.050 ;
        RECT 241.950 518.400 250.050 519.600 ;
        RECT 241.950 517.950 244.050 518.400 ;
        RECT 247.950 517.950 250.050 518.400 ;
        RECT 379.950 519.600 382.050 520.050 ;
        RECT 397.950 519.600 400.050 520.050 ;
        RECT 379.950 518.400 400.050 519.600 ;
        RECT 379.950 517.950 382.050 518.400 ;
        RECT 397.950 517.950 400.050 518.400 ;
        RECT 664.950 517.950 667.050 520.050 ;
        RECT 808.950 519.600 811.050 520.050 ;
        RECT 832.950 519.600 835.050 520.050 ;
        RECT 859.800 519.600 861.900 520.050 ;
        RECT 808.950 518.400 861.900 519.600 ;
        RECT 808.950 517.950 811.050 518.400 ;
        RECT 832.950 517.950 835.050 518.400 ;
        RECT 859.800 517.950 861.900 518.400 ;
        RECT 862.950 518.400 867.600 520.050 ;
        RECT 862.950 517.950 867.000 518.400 ;
        RECT 73.950 517.800 76.050 517.950 ;
        RECT 25.950 516.600 28.050 517.050 ;
        RECT 49.950 516.600 52.050 517.050 ;
        RECT 25.950 515.400 52.050 516.600 ;
        RECT 68.400 515.400 73.050 517.050 ;
        RECT 25.950 514.950 28.050 515.400 ;
        RECT 49.950 514.950 52.050 515.400 ;
        RECT 69.000 514.950 73.050 515.400 ;
        RECT 115.950 516.600 118.050 517.050 ;
        RECT 127.950 516.600 130.050 517.050 ;
        RECT 115.950 515.400 130.050 516.600 ;
        RECT 115.950 514.950 118.050 515.400 ;
        RECT 127.950 514.950 130.050 515.400 ;
        RECT 139.950 516.600 142.050 517.050 ;
        RECT 178.950 516.600 181.050 517.050 ;
        RECT 139.950 515.400 181.050 516.600 ;
        RECT 139.950 514.950 142.050 515.400 ;
        RECT 178.950 514.950 181.050 515.400 ;
        RECT 202.950 516.600 205.050 517.050 ;
        RECT 211.950 516.600 214.050 517.050 ;
        RECT 202.950 515.400 214.050 516.600 ;
        RECT 202.950 514.950 205.050 515.400 ;
        RECT 211.950 514.950 214.050 515.400 ;
        RECT 220.950 516.600 223.050 517.050 ;
        RECT 238.950 516.600 241.050 517.050 ;
        RECT 220.950 515.400 241.050 516.600 ;
        RECT 220.950 514.950 223.050 515.400 ;
        RECT 238.950 514.950 241.050 515.400 ;
        RECT 250.950 516.600 253.050 517.050 ;
        RECT 280.950 516.600 283.050 517.050 ;
        RECT 250.950 515.400 283.050 516.600 ;
        RECT 250.950 514.950 253.050 515.400 ;
        RECT 280.950 514.950 283.050 515.400 ;
        RECT 286.950 516.600 289.050 517.050 ;
        RECT 298.950 516.600 301.050 517.050 ;
        RECT 286.950 515.400 301.050 516.600 ;
        RECT 286.950 514.950 289.050 515.400 ;
        RECT 298.950 514.950 301.050 515.400 ;
        RECT 316.950 516.600 319.050 517.050 ;
        RECT 352.950 516.600 355.050 517.050 ;
        RECT 316.950 515.400 355.050 516.600 ;
        RECT 316.950 514.950 319.050 515.400 ;
        RECT 352.950 514.950 355.050 515.400 ;
        RECT 616.950 516.600 619.050 517.050 ;
        RECT 718.950 516.600 721.050 517.050 ;
        RECT 751.950 516.600 754.050 517.050 ;
        RECT 778.950 516.600 781.050 517.050 ;
        RECT 616.950 515.400 672.600 516.600 ;
        RECT 616.950 514.950 619.050 515.400 ;
        RECT 61.950 513.600 64.050 514.050 ;
        RECT 73.950 513.600 76.050 514.050 ;
        RECT 61.950 512.400 76.050 513.600 ;
        RECT 61.950 511.950 64.050 512.400 ;
        RECT 73.950 511.950 76.050 512.400 ;
        RECT 193.950 513.600 196.050 514.050 ;
        RECT 229.950 513.600 232.050 514.050 ;
        RECT 193.950 512.400 232.050 513.600 ;
        RECT 193.950 511.950 196.050 512.400 ;
        RECT 229.950 511.950 232.050 512.400 ;
        RECT 253.950 513.600 256.050 514.050 ;
        RECT 262.950 513.600 265.050 514.050 ;
        RECT 499.950 513.600 502.050 514.050 ;
        RECT 505.950 513.600 508.050 514.050 ;
        RECT 253.950 512.400 265.050 513.600 ;
        RECT 253.950 511.950 256.050 512.400 ;
        RECT 262.950 511.950 265.050 512.400 ;
        RECT 497.400 512.400 508.050 513.600 ;
        RECT 235.950 510.600 238.050 511.050 ;
        RECT 271.950 510.600 274.050 511.050 ;
        RECT 235.950 509.400 274.050 510.600 ;
        RECT 235.950 508.950 238.050 509.400 ;
        RECT 271.950 508.950 274.050 509.400 ;
        RECT 337.950 510.600 340.050 511.050 ;
        RECT 346.950 510.600 349.050 511.050 ;
        RECT 337.950 509.400 349.050 510.600 ;
        RECT 337.950 508.950 340.050 509.400 ;
        RECT 346.950 508.950 349.050 509.400 ;
        RECT 388.950 510.600 391.050 511.050 ;
        RECT 418.950 510.600 421.050 511.050 ;
        RECT 388.950 509.400 421.050 510.600 ;
        RECT 388.950 508.950 391.050 509.400 ;
        RECT 418.950 508.950 421.050 509.400 ;
        RECT 433.950 510.600 436.050 511.050 ;
        RECT 497.400 510.600 498.600 512.400 ;
        RECT 499.950 511.950 502.050 512.400 ;
        RECT 505.950 511.950 508.050 512.400 ;
        RECT 562.950 513.600 565.050 514.050 ;
        RECT 580.950 513.600 583.050 514.050 ;
        RECT 562.950 512.400 583.050 513.600 ;
        RECT 562.950 511.950 565.050 512.400 ;
        RECT 580.950 511.950 583.050 512.400 ;
        RECT 661.950 513.600 666.000 514.050 ;
        RECT 671.400 513.600 672.600 515.400 ;
        RECT 718.950 515.400 781.050 516.600 ;
        RECT 718.950 514.950 721.050 515.400 ;
        RECT 751.950 514.950 754.050 515.400 ;
        RECT 778.950 514.950 781.050 515.400 ;
        RECT 826.950 516.600 829.050 517.050 ;
        RECT 838.950 516.600 841.050 517.050 ;
        RECT 826.950 515.400 841.050 516.600 ;
        RECT 826.950 514.950 829.050 515.400 ;
        RECT 838.950 514.950 841.050 515.400 ;
        RECT 694.950 513.600 697.050 514.050 ;
        RECT 661.950 511.950 666.600 513.600 ;
        RECT 671.400 512.400 697.050 513.600 ;
        RECT 694.950 511.950 697.050 512.400 ;
        RECT 700.950 513.600 703.050 514.050 ;
        RECT 712.950 513.600 715.050 514.050 ;
        RECT 700.950 512.400 715.050 513.600 ;
        RECT 700.950 511.950 703.050 512.400 ;
        RECT 712.950 511.950 715.050 512.400 ;
        RECT 739.950 513.600 742.050 514.050 ;
        RECT 748.950 513.600 751.050 514.050 ;
        RECT 739.950 512.400 751.050 513.600 ;
        RECT 739.950 511.950 742.050 512.400 ;
        RECT 748.950 511.950 751.050 512.400 ;
        RECT 775.950 513.600 778.050 514.050 ;
        RECT 781.950 513.600 784.050 514.050 ;
        RECT 775.950 512.400 784.050 513.600 ;
        RECT 775.950 511.950 778.050 512.400 ;
        RECT 781.950 511.950 784.050 512.400 ;
        RECT 433.950 509.400 498.600 510.600 ;
        RECT 665.400 510.600 666.600 511.950 ;
        RECT 691.950 510.600 694.050 511.050 ;
        RECT 665.400 509.400 694.050 510.600 ;
        RECT 433.950 508.950 436.050 509.400 ;
        RECT 691.950 508.950 694.050 509.400 ;
        RECT 769.950 510.600 772.050 511.050 ;
        RECT 802.950 510.600 805.050 511.050 ;
        RECT 817.950 510.600 820.050 511.050 ;
        RECT 769.950 509.400 820.050 510.600 ;
        RECT 769.950 508.950 772.050 509.400 ;
        RECT 802.950 508.950 805.050 509.400 ;
        RECT 817.950 508.950 820.050 509.400 ;
        RECT 28.950 507.600 31.050 508.050 ;
        RECT 37.950 507.600 40.050 508.050 ;
        RECT 28.950 506.400 40.050 507.600 ;
        RECT 28.950 505.950 31.050 506.400 ;
        RECT 37.950 505.950 40.050 506.400 ;
        RECT 169.950 507.600 172.050 508.050 ;
        RECT 319.950 507.600 322.050 508.050 ;
        RECT 328.950 507.600 331.050 508.050 ;
        RECT 169.950 506.400 331.050 507.600 ;
        RECT 169.950 505.950 172.050 506.400 ;
        RECT 319.950 505.950 322.050 506.400 ;
        RECT 328.950 505.950 331.050 506.400 ;
        RECT 358.950 507.600 361.050 508.050 ;
        RECT 370.950 507.600 373.050 508.050 ;
        RECT 358.950 506.400 373.050 507.600 ;
        RECT 358.950 505.950 361.050 506.400 ;
        RECT 370.950 505.950 373.050 506.400 ;
        RECT 490.950 507.600 493.050 508.050 ;
        RECT 499.950 507.600 502.050 508.050 ;
        RECT 490.950 506.400 502.050 507.600 ;
        RECT 490.950 505.950 493.050 506.400 ;
        RECT 499.950 505.950 502.050 506.400 ;
        RECT 511.950 507.600 514.050 508.050 ;
        RECT 523.950 507.600 526.050 508.050 ;
        RECT 511.950 506.400 526.050 507.600 ;
        RECT 511.950 505.950 514.050 506.400 ;
        RECT 523.950 505.950 526.050 506.400 ;
        RECT 532.950 507.600 535.050 508.050 ;
        RECT 565.950 507.600 568.050 508.050 ;
        RECT 532.950 506.400 568.050 507.600 ;
        RECT 532.950 505.950 535.050 506.400 ;
        RECT 565.950 505.950 568.050 506.400 ;
        RECT 589.950 507.600 592.050 508.050 ;
        RECT 634.950 507.600 637.050 508.050 ;
        RECT 589.950 506.400 637.050 507.600 ;
        RECT 589.950 505.950 592.050 506.400 ;
        RECT 634.950 505.950 637.050 506.400 ;
        RECT 682.950 507.600 685.050 508.050 ;
        RECT 715.950 507.600 718.050 508.050 ;
        RECT 682.950 506.400 718.050 507.600 ;
        RECT 682.950 505.950 685.050 506.400 ;
        RECT 715.950 505.950 718.050 506.400 ;
        RECT 739.950 507.600 742.050 508.050 ;
        RECT 799.950 507.600 802.050 508.050 ;
        RECT 805.950 507.600 808.050 508.050 ;
        RECT 739.950 506.400 808.050 507.600 ;
        RECT 739.950 505.950 742.050 506.400 ;
        RECT 799.950 505.950 802.050 506.400 ;
        RECT 805.950 505.950 808.050 506.400 ;
        RECT 820.950 507.600 823.050 508.050 ;
        RECT 835.950 507.600 838.050 508.050 ;
        RECT 820.950 506.400 838.050 507.600 ;
        RECT 820.950 505.950 823.050 506.400 ;
        RECT 835.950 505.950 838.050 506.400 ;
        RECT 847.950 507.600 850.050 508.050 ;
        RECT 877.950 507.600 880.050 508.050 ;
        RECT 847.950 506.400 880.050 507.600 ;
        RECT 847.950 505.950 850.050 506.400 ;
        RECT 877.950 505.950 880.050 506.400 ;
        RECT 172.950 504.600 175.050 505.050 ;
        RECT 184.950 504.600 187.050 505.050 ;
        RECT 172.950 503.400 187.050 504.600 ;
        RECT 172.950 502.950 175.050 503.400 ;
        RECT 184.950 502.950 187.050 503.400 ;
        RECT 193.950 504.600 196.050 505.050 ;
        RECT 217.950 504.600 220.050 505.050 ;
        RECT 193.950 503.400 220.050 504.600 ;
        RECT 193.950 502.950 196.050 503.400 ;
        RECT 217.950 502.950 220.050 503.400 ;
        RECT 226.950 504.600 229.050 505.050 ;
        RECT 250.950 504.600 253.050 505.050 ;
        RECT 226.950 503.400 253.050 504.600 ;
        RECT 226.950 502.950 229.050 503.400 ;
        RECT 250.950 502.950 253.050 503.400 ;
        RECT 391.950 504.600 394.050 505.050 ;
        RECT 409.950 504.600 412.050 505.050 ;
        RECT 391.950 503.400 412.050 504.600 ;
        RECT 391.950 502.950 394.050 503.400 ;
        RECT 409.950 502.950 412.050 503.400 ;
        RECT 457.950 504.600 460.050 505.050 ;
        RECT 520.950 504.600 523.050 505.050 ;
        RECT 589.950 504.600 592.050 504.900 ;
        RECT 457.950 503.400 592.050 504.600 ;
        RECT 457.950 502.950 460.050 503.400 ;
        RECT 520.950 502.950 523.050 503.400 ;
        RECT 589.950 502.800 592.050 503.400 ;
        RECT 595.950 504.600 598.050 505.050 ;
        RECT 604.950 504.600 607.050 505.050 ;
        RECT 595.950 503.400 607.050 504.600 ;
        RECT 595.950 502.950 598.050 503.400 ;
        RECT 604.950 502.950 607.050 503.400 ;
        RECT 610.950 504.600 613.050 505.050 ;
        RECT 628.950 504.600 631.050 505.050 ;
        RECT 610.950 503.400 631.050 504.600 ;
        RECT 610.950 502.950 613.050 503.400 ;
        RECT 628.950 502.950 631.050 503.400 ;
        RECT 640.950 504.600 643.050 505.050 ;
        RECT 649.950 504.600 652.050 505.050 ;
        RECT 640.950 503.400 652.050 504.600 ;
        RECT 640.950 502.950 643.050 503.400 ;
        RECT 649.950 502.950 652.050 503.400 ;
        RECT 664.950 504.600 667.050 505.050 ;
        RECT 676.950 504.600 679.050 505.050 ;
        RECT 664.950 503.400 679.050 504.600 ;
        RECT 664.950 502.950 667.050 503.400 ;
        RECT 676.950 502.950 679.050 503.400 ;
        RECT 685.950 504.600 688.050 505.050 ;
        RECT 697.950 504.600 700.050 505.050 ;
        RECT 685.950 503.400 700.050 504.600 ;
        RECT 685.950 502.950 688.050 503.400 ;
        RECT 697.950 502.950 700.050 503.400 ;
        RECT 703.950 504.600 706.050 505.050 ;
        RECT 766.950 504.600 769.050 505.050 ;
        RECT 703.950 503.400 769.050 504.600 ;
        RECT 703.950 502.950 706.050 503.400 ;
        RECT 766.950 502.950 769.050 503.400 ;
        RECT 811.950 504.600 814.050 505.050 ;
        RECT 832.950 504.600 835.050 505.050 ;
        RECT 811.950 503.400 835.050 504.600 ;
        RECT 811.950 502.950 814.050 503.400 ;
        RECT 832.950 502.950 835.050 503.400 ;
        RECT 853.950 504.600 856.050 505.050 ;
        RECT 871.950 504.600 874.050 505.050 ;
        RECT 853.950 503.400 874.050 504.600 ;
        RECT 853.950 502.950 856.050 503.400 ;
        RECT 871.950 502.950 874.050 503.400 ;
        RECT 118.950 501.600 121.050 502.050 ;
        RECT 157.950 501.600 160.050 502.050 ;
        RECT 169.950 501.600 172.050 502.050 ;
        RECT 118.950 500.400 172.050 501.600 ;
        RECT 118.950 499.950 121.050 500.400 ;
        RECT 157.950 499.950 160.050 500.400 ;
        RECT 169.950 499.950 172.050 500.400 ;
        RECT 208.950 501.600 211.050 502.050 ;
        RECT 214.950 501.600 217.050 502.050 ;
        RECT 208.950 500.400 217.050 501.600 ;
        RECT 208.950 499.950 211.050 500.400 ;
        RECT 214.950 499.950 217.050 500.400 ;
        RECT 238.950 501.600 241.050 502.050 ;
        RECT 247.800 501.600 249.900 502.050 ;
        RECT 238.950 500.400 249.900 501.600 ;
        RECT 238.950 499.950 241.050 500.400 ;
        RECT 247.800 499.950 249.900 500.400 ;
        RECT 250.950 501.600 253.050 501.900 ;
        RECT 262.950 501.600 265.050 502.050 ;
        RECT 250.950 500.400 265.050 501.600 ;
        RECT 250.950 499.800 253.050 500.400 ;
        RECT 262.950 499.950 265.050 500.400 ;
        RECT 352.950 501.600 355.050 502.050 ;
        RECT 397.950 501.600 400.050 502.050 ;
        RECT 352.950 500.400 400.050 501.600 ;
        RECT 352.950 499.950 355.050 500.400 ;
        RECT 397.950 499.950 400.050 500.400 ;
        RECT 415.950 501.600 418.050 502.050 ;
        RECT 433.950 501.600 436.050 502.050 ;
        RECT 415.950 500.400 436.050 501.600 ;
        RECT 415.950 499.950 418.050 500.400 ;
        RECT 433.950 499.950 436.050 500.400 ;
        RECT 442.950 501.600 445.050 502.050 ;
        RECT 451.950 501.600 454.050 502.050 ;
        RECT 442.950 500.400 454.050 501.600 ;
        RECT 442.950 499.950 445.050 500.400 ;
        RECT 451.950 499.950 454.050 500.400 ;
        RECT 523.950 501.600 526.050 502.050 ;
        RECT 547.950 501.600 550.050 502.050 ;
        RECT 523.950 500.400 550.050 501.600 ;
        RECT 523.950 499.950 526.050 500.400 ;
        RECT 547.950 499.950 550.050 500.400 ;
        RECT 592.950 501.600 595.050 502.050 ;
        RECT 670.950 501.600 673.050 502.050 ;
        RECT 706.950 501.600 709.050 502.050 ;
        RECT 592.950 500.400 709.050 501.600 ;
        RECT 592.950 499.950 595.050 500.400 ;
        RECT 670.950 499.950 673.050 500.400 ;
        RECT 706.950 499.950 709.050 500.400 ;
        RECT 721.950 501.600 724.050 502.050 ;
        RECT 763.950 501.600 766.050 502.050 ;
        RECT 721.950 500.400 766.050 501.600 ;
        RECT 721.950 499.950 724.050 500.400 ;
        RECT 763.950 499.950 766.050 500.400 ;
        RECT 796.950 501.600 799.050 502.050 ;
        RECT 808.950 501.600 811.050 502.050 ;
        RECT 796.950 500.400 811.050 501.600 ;
        RECT 796.950 499.950 799.050 500.400 ;
        RECT 808.950 499.950 811.050 500.400 ;
        RECT 115.950 498.600 118.050 499.050 ;
        RECT 133.950 498.600 136.050 499.050 ;
        RECT 115.950 497.400 136.050 498.600 ;
        RECT 115.950 496.950 118.050 497.400 ;
        RECT 133.950 496.950 136.050 497.400 ;
        RECT 205.950 498.600 208.050 499.050 ;
        RECT 259.950 498.600 262.050 499.050 ;
        RECT 268.950 498.600 271.050 499.050 ;
        RECT 205.950 497.400 271.050 498.600 ;
        RECT 205.950 496.950 208.050 497.400 ;
        RECT 259.950 496.950 262.050 497.400 ;
        RECT 268.950 496.950 271.050 497.400 ;
        RECT 322.950 498.600 325.050 499.050 ;
        RECT 331.950 498.600 334.050 498.900 ;
        RECT 322.950 497.400 334.050 498.600 ;
        RECT 322.950 496.950 325.050 497.400 ;
        RECT 331.950 496.800 334.050 497.400 ;
        RECT 409.950 498.600 412.050 499.050 ;
        RECT 427.950 498.600 430.050 499.050 ;
        RECT 454.950 498.600 457.050 499.050 ;
        RECT 472.950 498.600 475.050 499.050 ;
        RECT 409.950 497.400 430.050 498.600 ;
        RECT 409.950 496.950 412.050 497.400 ;
        RECT 427.950 496.950 430.050 497.400 ;
        RECT 449.400 497.400 457.050 498.600 ;
        RECT 31.950 496.050 34.050 496.500 ;
        RECT 40.950 496.050 43.050 496.500 ;
        RECT 31.950 494.850 43.050 496.050 ;
        RECT 31.950 494.400 34.050 494.850 ;
        RECT 40.950 494.400 43.050 494.850 ;
        RECT 82.950 494.400 85.050 496.500 ;
        RECT 94.950 495.600 97.050 496.050 ;
        RECT 112.950 495.600 115.050 496.050 ;
        RECT 127.950 495.600 130.050 496.200 ;
        RECT 94.950 494.400 115.050 495.600 ;
        RECT 40.950 489.600 43.050 490.050 ;
        RECT 46.950 489.600 49.050 489.900 ;
        RECT 13.950 489.150 16.050 489.600 ;
        RECT 19.950 489.150 22.050 489.600 ;
        RECT 13.950 487.950 22.050 489.150 ;
        RECT 40.950 488.400 49.050 489.600 ;
        RECT 40.950 487.950 43.050 488.400 ;
        RECT 13.950 487.500 16.050 487.950 ;
        RECT 19.950 487.500 22.050 487.950 ;
        RECT 46.950 487.800 49.050 488.400 ;
        RECT 52.950 489.600 55.050 489.900 ;
        RECT 70.950 489.600 73.050 489.900 ;
        RECT 52.950 488.400 73.050 489.600 ;
        RECT 52.950 487.800 55.050 488.400 ;
        RECT 70.950 487.800 73.050 488.400 ;
        RECT 76.950 489.600 79.050 489.900 ;
        RECT 83.400 489.600 84.600 494.400 ;
        RECT 94.950 493.950 97.050 494.400 ;
        RECT 112.950 493.950 115.050 494.400 ;
        RECT 116.400 494.400 130.050 495.600 ;
        RECT 91.950 492.600 94.050 493.050 ;
        RECT 116.400 492.600 117.600 494.400 ;
        RECT 127.950 494.100 130.050 494.400 ;
        RECT 142.950 495.600 145.050 496.050 ;
        RECT 148.950 495.600 151.050 496.200 ;
        RECT 142.950 494.400 151.050 495.600 ;
        RECT 142.950 493.950 145.050 494.400 ;
        RECT 148.950 494.100 151.050 494.400 ;
        RECT 154.950 495.600 157.050 496.200 ;
        RECT 160.950 495.600 163.050 496.050 ;
        RECT 154.950 494.400 163.050 495.600 ;
        RECT 154.950 494.100 157.050 494.400 ;
        RECT 160.950 493.950 163.050 494.400 ;
        RECT 181.950 495.600 184.050 496.050 ;
        RECT 199.950 495.600 202.050 496.050 ;
        RECT 181.950 494.400 202.050 495.600 ;
        RECT 181.950 493.950 184.050 494.400 ;
        RECT 199.950 493.950 202.050 494.400 ;
        RECT 211.950 495.600 214.050 496.050 ;
        RECT 226.950 495.600 229.050 496.050 ;
        RECT 211.950 494.400 229.050 495.600 ;
        RECT 211.950 493.950 214.050 494.400 ;
        RECT 226.950 493.950 229.050 494.400 ;
        RECT 238.950 495.600 241.050 496.200 ;
        RECT 274.950 496.050 277.050 496.500 ;
        RECT 286.950 496.050 289.050 496.500 ;
        RECT 238.950 494.400 261.600 495.600 ;
        RECT 274.950 494.850 289.050 496.050 ;
        RECT 303.000 495.600 307.050 496.050 ;
        RECT 274.950 494.400 277.050 494.850 ;
        RECT 286.950 494.400 289.050 494.850 ;
        RECT 238.950 494.100 241.050 494.400 ;
        RECT 91.950 491.400 117.600 492.600 ;
        RECT 91.950 490.950 94.050 491.400 ;
        RECT 130.950 489.600 133.050 489.900 ;
        RECT 151.950 489.600 154.050 489.900 ;
        RECT 76.950 488.400 84.600 489.600 ;
        RECT 94.950 489.150 97.050 489.600 ;
        RECT 100.950 489.150 103.050 489.600 ;
        RECT 76.950 487.800 79.050 488.400 ;
        RECT 94.950 487.950 103.050 489.150 ;
        RECT 94.950 487.500 97.050 487.950 ;
        RECT 100.950 487.500 103.050 487.950 ;
        RECT 130.950 488.400 154.050 489.600 ;
        RECT 130.950 487.800 133.050 488.400 ;
        RECT 151.950 487.800 154.050 488.400 ;
        RECT 160.950 489.450 163.050 489.900 ;
        RECT 172.950 489.600 175.050 489.900 ;
        RECT 190.950 489.600 193.050 489.900 ;
        RECT 172.950 489.450 193.050 489.600 ;
        RECT 160.950 488.400 193.050 489.450 ;
        RECT 160.950 488.250 175.050 488.400 ;
        RECT 160.950 487.800 163.050 488.250 ;
        RECT 172.950 487.800 175.050 488.250 ;
        RECT 190.950 487.800 193.050 488.400 ;
        RECT 208.950 489.450 211.050 489.900 ;
        RECT 223.800 489.450 225.900 489.900 ;
        RECT 208.950 488.250 225.900 489.450 ;
        RECT 208.950 487.800 211.050 488.250 ;
        RECT 223.800 487.800 225.900 488.250 ;
        RECT 226.950 489.450 229.050 489.900 ;
        RECT 235.950 489.450 238.050 489.900 ;
        RECT 226.950 488.250 238.050 489.450 ;
        RECT 226.950 487.800 229.050 488.250 ;
        RECT 235.950 487.800 238.050 488.250 ;
        RECT 244.950 489.600 247.050 490.050 ;
        RECT 250.950 489.600 253.050 490.050 ;
        RECT 260.400 489.900 261.600 494.400 ;
        RECT 302.400 493.950 307.050 495.600 ;
        RECT 328.950 493.950 331.050 496.050 ;
        RECT 352.950 494.100 355.050 496.200 ;
        RECT 406.950 495.600 409.050 496.200 ;
        RECT 406.950 494.400 426.600 495.600 ;
        RECT 406.950 494.100 409.050 494.400 ;
        RECT 244.950 488.400 253.050 489.600 ;
        RECT 244.950 487.950 247.050 488.400 ;
        RECT 250.950 487.950 253.050 488.400 ;
        RECT 259.950 487.800 262.050 489.900 ;
        RECT 302.400 489.600 303.600 493.950 ;
        RECT 329.400 490.050 330.600 493.950 ;
        RECT 337.950 492.600 340.050 493.050 ;
        RECT 337.950 491.400 351.600 492.600 ;
        RECT 337.950 490.950 340.050 491.400 ;
        RECT 301.950 489.000 318.600 489.600 ;
        RECT 301.950 488.400 319.050 489.000 ;
        RECT 301.950 487.500 304.050 488.400 ;
        RECT 4.950 486.600 7.050 487.050 ;
        RECT 109.950 486.600 112.050 487.050 ;
        RECT 4.950 485.400 112.050 486.600 ;
        RECT 4.950 484.950 7.050 485.400 ;
        RECT 109.950 484.950 112.050 485.400 ;
        RECT 202.950 486.600 205.050 487.050 ;
        RECT 202.950 485.400 219.600 486.600 ;
        RECT 202.950 484.950 205.050 485.400 ;
        RECT 184.950 483.600 187.050 484.050 ;
        RECT 214.950 483.600 217.050 484.050 ;
        RECT 184.950 482.400 217.050 483.600 ;
        RECT 218.400 483.600 219.600 485.400 ;
        RECT 316.950 484.950 319.050 488.400 ;
        RECT 328.950 487.950 331.050 490.050 ;
        RECT 350.400 489.900 351.600 491.400 ;
        RECT 353.400 490.050 354.600 494.100 ;
        RECT 349.950 487.800 352.050 489.900 ;
        RECT 353.400 488.400 358.050 490.050 ;
        RECT 425.400 489.900 426.600 494.400 ;
        RECT 354.000 487.950 358.050 488.400 ;
        RECT 370.950 489.150 373.050 489.600 ;
        RECT 385.950 489.150 388.050 489.600 ;
        RECT 370.950 487.950 388.050 489.150 ;
        RECT 370.950 487.500 373.050 487.950 ;
        RECT 385.950 487.500 388.050 487.950 ;
        RECT 424.950 487.800 427.050 489.900 ;
        RECT 430.950 489.600 433.050 489.900 ;
        RECT 439.950 489.600 442.050 490.050 ;
        RECT 449.400 489.900 450.600 497.400 ;
        RECT 454.950 496.950 457.050 497.400 ;
        RECT 461.400 497.400 475.050 498.600 ;
        RECT 461.400 495.600 462.600 497.400 ;
        RECT 472.950 496.950 475.050 497.400 ;
        RECT 523.950 498.600 526.050 498.900 ;
        RECT 643.950 498.600 646.050 499.050 ;
        RECT 523.950 497.400 588.600 498.600 ;
        RECT 523.950 496.800 526.050 497.400 ;
        RECT 455.400 494.400 462.600 495.600 ;
        RECT 478.950 496.050 481.050 496.500 ;
        RECT 490.950 496.050 493.050 496.500 ;
        RECT 478.950 494.850 493.050 496.050 ;
        RECT 478.950 494.400 481.050 494.850 ;
        RECT 490.950 494.400 493.050 494.850 ;
        RECT 455.400 489.900 456.600 494.400 ;
        RECT 502.950 493.950 505.050 496.050 ;
        RECT 532.950 495.600 535.050 496.200 ;
        RECT 509.400 494.400 535.050 495.600 ;
        RECT 503.400 490.050 504.600 493.950 ;
        RECT 430.950 488.400 442.050 489.600 ;
        RECT 430.950 487.800 433.050 488.400 ;
        RECT 439.950 487.950 442.050 488.400 ;
        RECT 448.950 487.800 451.050 489.900 ;
        RECT 454.950 487.800 457.050 489.900 ;
        RECT 502.950 487.950 505.050 490.050 ;
        RECT 509.400 489.900 510.600 494.400 ;
        RECT 532.950 494.100 535.050 494.400 ;
        RECT 556.950 492.600 559.050 496.050 ;
        RECT 574.950 495.600 577.050 496.200 ;
        RECT 580.950 495.600 583.050 496.050 ;
        RECT 574.950 494.400 583.050 495.600 ;
        RECT 587.400 495.600 588.600 497.400 ;
        RECT 617.400 497.400 646.050 498.600 ;
        RECT 601.950 495.600 604.050 496.200 ;
        RECT 613.950 495.600 616.050 496.200 ;
        RECT 587.400 494.400 616.050 495.600 ;
        RECT 574.950 494.100 577.050 494.400 ;
        RECT 580.950 493.950 583.050 494.400 ;
        RECT 601.950 494.100 604.050 494.400 ;
        RECT 613.950 494.100 616.050 494.400 ;
        RECT 583.950 492.600 586.050 493.050 ;
        RECT 617.400 492.600 618.600 497.400 ;
        RECT 643.950 496.950 646.050 497.400 ;
        RECT 772.950 498.600 775.050 499.050 ;
        RECT 832.950 498.600 835.050 499.050 ;
        RECT 853.950 498.600 856.050 499.050 ;
        RECT 772.950 497.400 810.600 498.600 ;
        RECT 772.950 496.950 775.050 497.400 ;
        RECT 634.950 495.600 639.000 496.050 ;
        RECT 646.950 495.750 649.050 496.200 ;
        RECT 661.950 495.750 664.050 496.200 ;
        RECT 634.950 493.950 639.600 495.600 ;
        RECT 646.950 494.550 664.050 495.750 ;
        RECT 646.950 494.100 649.050 494.550 ;
        RECT 661.950 494.100 664.050 494.550 ;
        RECT 667.950 495.600 670.050 496.200 ;
        RECT 694.950 495.600 697.050 496.050 ;
        RECT 667.950 494.400 697.050 495.600 ;
        RECT 667.950 494.100 670.050 494.400 ;
        RECT 694.950 493.950 697.050 494.400 ;
        RECT 712.950 495.600 715.050 496.200 ;
        RECT 727.950 495.750 730.050 496.200 ;
        RECT 733.950 495.750 736.050 496.200 ;
        RECT 712.950 494.400 726.600 495.600 ;
        RECT 712.950 494.100 715.050 494.400 ;
        RECT 556.950 492.000 586.050 492.600 ;
        RECT 605.400 492.000 618.600 492.600 ;
        RECT 557.400 491.400 586.050 492.000 ;
        RECT 583.950 490.950 586.050 491.400 ;
        RECT 604.950 491.400 618.600 492.000 ;
        RECT 508.950 489.600 511.050 489.900 ;
        RECT 526.950 489.600 529.050 490.050 ;
        RECT 508.950 488.400 529.050 489.600 ;
        RECT 508.950 487.800 511.050 488.400 ;
        RECT 526.950 487.950 529.050 488.400 ;
        RECT 604.950 487.950 607.050 491.400 ;
        RECT 638.400 489.900 639.600 493.950 ;
        RECT 725.400 492.600 726.600 494.400 ;
        RECT 727.950 494.550 736.050 495.750 ;
        RECT 727.950 494.100 730.050 494.550 ;
        RECT 733.950 494.100 736.050 494.550 ;
        RECT 754.950 493.950 757.050 496.050 ;
        RECT 769.950 493.950 772.050 496.050 ;
        RECT 775.950 493.950 778.050 496.050 ;
        RECT 809.400 495.600 810.600 497.400 ;
        RECT 832.950 497.400 856.050 498.600 ;
        RECT 832.950 496.950 835.050 497.400 ;
        RECT 853.950 496.950 856.050 497.400 ;
        RECT 865.950 498.600 868.050 499.050 ;
        RECT 874.950 498.600 877.050 499.050 ;
        RECT 865.950 497.400 877.050 498.600 ;
        RECT 865.950 496.950 868.050 497.400 ;
        RECT 874.950 496.950 877.050 497.400 ;
        RECT 811.950 495.600 814.050 496.200 ;
        RECT 809.400 494.400 814.050 495.600 ;
        RECT 811.950 494.100 814.050 494.400 ;
        RECT 823.950 493.950 826.050 496.050 ;
        RECT 829.950 495.600 832.050 496.200 ;
        RECT 838.950 495.600 841.050 496.050 ;
        RECT 829.950 494.400 841.050 495.600 ;
        RECT 829.950 494.100 832.050 494.400 ;
        RECT 838.950 493.950 841.050 494.400 ;
        RECT 847.950 493.950 850.050 496.050 ;
        RECT 859.800 495.600 861.900 496.200 ;
        RECT 854.400 494.400 861.900 495.600 ;
        RECT 725.400 491.400 732.600 492.600 ;
        RECT 637.950 487.800 640.050 489.900 ;
        RECT 649.950 489.450 652.050 489.900 ;
        RECT 664.950 489.600 667.050 489.900 ;
        RECT 682.950 489.600 685.050 489.900 ;
        RECT 664.950 489.450 685.050 489.600 ;
        RECT 649.950 488.400 685.050 489.450 ;
        RECT 649.950 488.250 667.050 488.400 ;
        RECT 649.950 487.800 652.050 488.250 ;
        RECT 664.950 487.800 667.050 488.250 ;
        RECT 682.950 487.800 685.050 488.400 ;
        RECT 688.950 489.450 691.050 489.900 ;
        RECT 694.950 489.450 697.050 489.900 ;
        RECT 688.950 488.250 697.050 489.450 ;
        RECT 688.950 487.800 691.050 488.250 ;
        RECT 694.950 487.800 697.050 488.250 ;
        RECT 700.950 489.600 703.050 490.050 ;
        RECT 731.400 489.900 732.600 491.400 ;
        RECT 755.400 490.050 756.600 493.950 ;
        RECT 709.950 489.600 712.050 489.900 ;
        RECT 700.950 488.400 712.050 489.600 ;
        RECT 700.950 487.950 703.050 488.400 ;
        RECT 709.950 487.800 712.050 488.400 ;
        RECT 730.950 487.800 733.050 489.900 ;
        RECT 754.950 487.950 757.050 490.050 ;
        RECT 770.400 489.600 771.600 493.950 ;
        RECT 776.400 490.050 777.600 493.950 ;
        RECT 824.400 490.050 825.600 493.950 ;
        RECT 770.400 488.400 774.600 489.600 ;
        RECT 773.400 487.050 774.600 488.400 ;
        RECT 775.950 487.950 778.050 490.050 ;
        RECT 784.950 489.600 787.050 489.900 ;
        RECT 814.950 489.600 817.050 490.050 ;
        RECT 784.950 488.400 817.050 489.600 ;
        RECT 784.950 487.800 787.050 488.400 ;
        RECT 814.950 487.950 817.050 488.400 ;
        RECT 823.950 487.950 826.050 490.050 ;
        RECT 835.950 489.600 838.050 490.050 ;
        RECT 848.400 489.600 849.600 493.950 ;
        RECT 835.950 488.400 849.600 489.600 ;
        RECT 835.950 487.950 838.050 488.400 ;
        RECT 854.400 487.050 855.600 494.400 ;
        RECT 859.800 494.100 861.900 494.400 ;
        RECT 862.950 493.950 865.050 496.050 ;
        RECT 880.950 495.600 883.050 496.200 ;
        RECT 886.950 495.600 889.050 496.050 ;
        RECT 880.950 494.400 889.050 495.600 ;
        RECT 880.950 494.100 883.050 494.400 ;
        RECT 886.950 493.950 889.050 494.400 ;
        RECT 863.400 489.600 864.600 493.950 ;
        RECT 871.950 489.600 874.050 489.900 ;
        RECT 863.400 488.400 874.050 489.600 ;
        RECT 871.950 487.800 874.050 488.400 ;
        RECT 331.950 486.600 334.050 487.050 ;
        RECT 343.950 486.600 346.050 487.050 ;
        RECT 331.950 485.400 346.050 486.600 ;
        RECT 331.950 484.950 334.050 485.400 ;
        RECT 343.950 484.950 346.050 485.400 ;
        RECT 529.950 486.600 532.050 487.050 ;
        RECT 562.950 486.600 565.050 487.050 ;
        RECT 577.950 486.600 580.050 487.050 ;
        RECT 634.950 486.600 637.050 487.050 ;
        RECT 529.950 485.400 637.050 486.600 ;
        RECT 529.950 484.950 532.050 485.400 ;
        RECT 562.950 484.950 565.050 485.400 ;
        RECT 577.950 484.950 580.050 485.400 ;
        RECT 634.950 484.950 637.050 485.400 ;
        RECT 736.950 486.600 739.050 487.050 ;
        RECT 769.950 486.600 772.050 487.050 ;
        RECT 736.950 485.400 772.050 486.600 ;
        RECT 773.400 486.900 777.000 487.050 ;
        RECT 773.400 485.400 778.050 486.900 ;
        RECT 736.950 484.950 739.050 485.400 ;
        RECT 769.950 484.950 772.050 485.400 ;
        RECT 774.000 484.950 778.050 485.400 ;
        RECT 787.950 486.600 790.050 487.050 ;
        RECT 796.950 486.600 799.050 487.050 ;
        RECT 787.950 485.400 799.050 486.600 ;
        RECT 787.950 484.950 790.050 485.400 ;
        RECT 796.950 484.950 799.050 485.400 ;
        RECT 853.950 484.950 856.050 487.050 ;
        RECT 775.950 484.800 778.050 484.950 ;
        RECT 262.950 483.600 265.050 484.050 ;
        RECT 218.400 482.400 265.050 483.600 ;
        RECT 184.950 481.950 187.050 482.400 ;
        RECT 214.950 481.950 217.050 482.400 ;
        RECT 262.950 481.950 265.050 482.400 ;
        RECT 376.950 483.600 379.050 484.050 ;
        RECT 391.950 483.600 394.050 484.050 ;
        RECT 376.950 482.400 394.050 483.600 ;
        RECT 376.950 481.950 379.050 482.400 ;
        RECT 391.950 481.950 394.050 482.400 ;
        RECT 442.950 483.600 445.050 484.050 ;
        RECT 472.950 483.600 475.050 484.050 ;
        RECT 442.950 482.400 475.050 483.600 ;
        RECT 442.950 481.950 445.050 482.400 ;
        RECT 472.950 481.950 475.050 482.400 ;
        RECT 499.950 483.600 502.050 484.050 ;
        RECT 514.950 483.600 517.050 484.050 ;
        RECT 499.950 482.400 517.050 483.600 ;
        RECT 499.950 481.950 502.050 482.400 ;
        RECT 514.950 481.950 517.050 482.400 ;
        RECT 586.950 483.600 589.050 483.900 ;
        RECT 598.950 483.600 601.050 484.050 ;
        RECT 616.950 483.600 619.050 484.050 ;
        RECT 586.950 482.400 619.050 483.600 ;
        RECT 586.950 481.800 589.050 482.400 ;
        RECT 598.950 481.950 601.050 482.400 ;
        RECT 616.950 481.950 619.050 482.400 ;
        RECT 715.950 483.600 718.050 484.050 ;
        RECT 757.950 483.600 760.050 484.050 ;
        RECT 715.950 482.400 760.050 483.600 ;
        RECT 715.950 481.950 718.050 482.400 ;
        RECT 757.950 481.950 760.050 482.400 ;
        RECT 763.950 483.600 766.050 484.050 ;
        RECT 778.950 483.600 781.050 484.050 ;
        RECT 763.950 482.400 781.050 483.600 ;
        RECT 763.950 481.950 766.050 482.400 ;
        RECT 778.950 481.950 781.050 482.400 ;
        RECT 805.950 483.600 808.050 484.050 ;
        RECT 832.950 483.600 835.050 484.050 ;
        RECT 805.950 482.400 835.050 483.600 ;
        RECT 805.950 481.950 808.050 482.400 ;
        RECT 832.950 481.950 835.050 482.400 ;
        RECT 844.950 483.600 847.050 484.050 ;
        RECT 865.950 483.600 868.050 484.050 ;
        RECT 844.950 482.400 868.050 483.600 ;
        RECT 844.950 481.950 847.050 482.400 ;
        RECT 865.950 481.950 868.050 482.400 ;
        RECT 292.950 480.600 295.050 481.050 ;
        RECT 304.950 480.600 307.050 481.050 ;
        RECT 292.950 479.400 307.050 480.600 ;
        RECT 292.950 478.950 295.050 479.400 ;
        RECT 304.950 478.950 307.050 479.400 ;
        RECT 397.950 480.600 400.050 481.050 ;
        RECT 409.950 480.600 412.050 481.050 ;
        RECT 397.950 479.400 412.050 480.600 ;
        RECT 397.950 478.950 400.050 479.400 ;
        RECT 409.950 478.950 412.050 479.400 ;
        RECT 634.950 480.600 637.050 481.050 ;
        RECT 670.950 480.600 673.050 481.050 ;
        RECT 634.950 479.400 673.050 480.600 ;
        RECT 634.950 478.950 637.050 479.400 ;
        RECT 670.950 478.950 673.050 479.400 ;
        RECT 697.950 480.600 700.050 481.050 ;
        RECT 784.950 480.600 787.050 481.050 ;
        RECT 697.950 479.400 787.050 480.600 ;
        RECT 697.950 478.950 700.050 479.400 ;
        RECT 784.950 478.950 787.050 479.400 ;
        RECT 196.950 477.600 199.050 478.050 ;
        RECT 205.950 477.600 208.050 478.050 ;
        RECT 241.950 477.600 244.050 478.050 ;
        RECT 196.950 476.400 244.050 477.600 ;
        RECT 196.950 475.950 199.050 476.400 ;
        RECT 205.950 475.950 208.050 476.400 ;
        RECT 241.950 475.950 244.050 476.400 ;
        RECT 253.950 477.600 256.050 478.050 ;
        RECT 265.950 477.600 268.050 478.050 ;
        RECT 253.950 476.400 268.050 477.600 ;
        RECT 253.950 475.950 256.050 476.400 ;
        RECT 265.950 475.950 268.050 476.400 ;
        RECT 310.950 477.600 313.050 478.050 ;
        RECT 319.950 477.600 322.050 478.050 ;
        RECT 325.950 477.600 328.050 478.050 ;
        RECT 337.950 477.600 340.050 478.050 ;
        RECT 310.950 476.400 340.050 477.600 ;
        RECT 310.950 475.950 313.050 476.400 ;
        RECT 319.950 475.950 322.050 476.400 ;
        RECT 325.950 475.950 328.050 476.400 ;
        RECT 337.950 475.950 340.050 476.400 ;
        RECT 418.950 477.600 421.050 478.050 ;
        RECT 493.950 477.600 496.050 478.050 ;
        RECT 418.950 476.400 496.050 477.600 ;
        RECT 418.950 475.950 421.050 476.400 ;
        RECT 493.950 475.950 496.050 476.400 ;
        RECT 631.950 477.600 634.050 478.050 ;
        RECT 649.950 477.600 652.050 478.050 ;
        RECT 691.950 477.600 694.050 478.050 ;
        RECT 631.950 476.400 694.050 477.600 ;
        RECT 631.950 475.950 634.050 476.400 ;
        RECT 649.950 475.950 652.050 476.400 ;
        RECT 691.950 475.950 694.050 476.400 ;
        RECT 706.950 477.600 709.050 478.050 ;
        RECT 775.950 477.600 778.050 478.050 ;
        RECT 706.950 476.400 778.050 477.600 ;
        RECT 706.950 475.950 709.050 476.400 ;
        RECT 775.950 475.950 778.050 476.400 ;
        RECT 781.950 477.600 784.050 478.050 ;
        RECT 829.950 477.600 832.050 478.050 ;
        RECT 781.950 476.400 832.050 477.600 ;
        RECT 781.950 475.950 784.050 476.400 ;
        RECT 829.950 475.950 832.050 476.400 ;
        RECT 838.950 477.600 841.050 478.050 ;
        RECT 874.950 477.600 877.050 478.050 ;
        RECT 838.950 476.400 877.050 477.600 ;
        RECT 838.950 475.950 841.050 476.400 ;
        RECT 874.950 475.950 877.050 476.400 ;
        RECT 298.950 474.600 301.050 475.050 ;
        RECT 307.950 474.600 310.050 475.050 ;
        RECT 298.950 473.400 310.050 474.600 ;
        RECT 298.950 472.950 301.050 473.400 ;
        RECT 307.950 472.950 310.050 473.400 ;
        RECT 370.950 474.600 373.050 475.050 ;
        RECT 421.950 474.600 424.050 475.050 ;
        RECT 370.950 473.400 424.050 474.600 ;
        RECT 370.950 472.950 373.050 473.400 ;
        RECT 421.950 472.950 424.050 473.400 ;
        RECT 502.950 474.600 505.050 475.050 ;
        RECT 544.950 474.600 547.050 475.050 ;
        RECT 502.950 473.400 547.050 474.600 ;
        RECT 502.950 472.950 505.050 473.400 ;
        RECT 544.950 472.950 547.050 473.400 ;
        RECT 754.950 474.600 757.050 475.050 ;
        RECT 763.950 474.600 766.050 475.050 ;
        RECT 772.950 474.600 775.050 475.050 ;
        RECT 754.950 473.400 775.050 474.600 ;
        RECT 754.950 472.950 757.050 473.400 ;
        RECT 763.950 472.950 766.050 473.400 ;
        RECT 772.950 472.950 775.050 473.400 ;
        RECT 778.950 474.600 781.050 475.050 ;
        RECT 790.950 474.600 793.050 475.050 ;
        RECT 778.950 473.400 793.050 474.600 ;
        RECT 778.950 472.950 781.050 473.400 ;
        RECT 790.950 472.950 793.050 473.400 ;
        RECT 175.950 471.600 178.050 472.050 ;
        RECT 196.950 471.600 199.050 472.050 ;
        RECT 175.950 470.400 199.050 471.600 ;
        RECT 175.950 469.950 178.050 470.400 ;
        RECT 196.950 469.950 199.050 470.400 ;
        RECT 304.950 471.600 307.050 472.050 ;
        RECT 346.950 471.600 349.050 472.050 ;
        RECT 304.950 470.400 349.050 471.600 ;
        RECT 304.950 469.950 307.050 470.400 ;
        RECT 346.950 469.950 349.050 470.400 ;
        RECT 361.950 471.600 364.050 472.050 ;
        RECT 427.950 471.600 430.050 472.050 ;
        RECT 361.950 470.400 430.050 471.600 ;
        RECT 361.950 469.950 364.050 470.400 ;
        RECT 427.950 469.950 430.050 470.400 ;
        RECT 556.950 471.600 559.050 472.050 ;
        RECT 673.950 471.600 676.050 472.050 ;
        RECT 556.950 470.400 676.050 471.600 ;
        RECT 556.950 469.950 559.050 470.400 ;
        RECT 673.950 469.950 676.050 470.400 ;
        RECT 724.950 471.600 727.050 472.050 ;
        RECT 745.950 471.600 748.050 472.050 ;
        RECT 724.950 470.400 748.050 471.600 ;
        RECT 724.950 469.950 727.050 470.400 ;
        RECT 745.950 469.950 748.050 470.400 ;
        RECT 841.950 471.600 844.050 472.050 ;
        RECT 895.950 471.600 898.050 472.050 ;
        RECT 841.950 470.400 898.050 471.600 ;
        RECT 841.950 469.950 844.050 470.400 ;
        RECT 895.950 469.950 898.050 470.400 ;
        RECT 286.950 468.600 289.050 469.050 ;
        RECT 301.950 468.600 304.050 469.050 ;
        RECT 286.950 467.400 304.050 468.600 ;
        RECT 286.950 466.950 289.050 467.400 ;
        RECT 301.950 466.950 304.050 467.400 ;
        RECT 493.950 468.600 496.050 469.050 ;
        RECT 523.950 468.600 526.050 469.050 ;
        RECT 493.950 467.400 526.050 468.600 ;
        RECT 493.950 466.950 496.050 467.400 ;
        RECT 523.950 466.950 526.050 467.400 ;
        RECT 589.950 468.600 592.050 469.050 ;
        RECT 700.950 468.600 703.050 469.050 ;
        RECT 589.950 467.400 703.050 468.600 ;
        RECT 589.950 466.950 592.050 467.400 ;
        RECT 700.950 466.950 703.050 467.400 ;
        RECT 799.950 468.600 802.050 469.050 ;
        RECT 811.950 468.600 814.050 469.050 ;
        RECT 799.950 467.400 814.050 468.600 ;
        RECT 799.950 466.950 802.050 467.400 ;
        RECT 811.950 466.950 814.050 467.400 ;
        RECT 859.950 468.600 862.050 469.050 ;
        RECT 886.950 468.600 889.050 469.050 ;
        RECT 859.950 467.400 889.050 468.600 ;
        RECT 859.950 466.950 862.050 467.400 ;
        RECT 886.950 466.950 889.050 467.400 ;
        RECT 229.950 465.600 232.050 466.050 ;
        RECT 238.950 465.600 241.050 466.050 ;
        RECT 229.950 464.400 241.050 465.600 ;
        RECT 229.950 463.950 232.050 464.400 ;
        RECT 238.950 463.950 241.050 464.400 ;
        RECT 259.950 465.600 262.050 466.050 ;
        RECT 316.950 465.600 319.050 466.050 ;
        RECT 259.950 464.400 319.050 465.600 ;
        RECT 259.950 463.950 262.050 464.400 ;
        RECT 316.950 463.950 319.050 464.400 ;
        RECT 355.950 465.600 358.050 466.050 ;
        RECT 370.950 465.600 373.050 466.050 ;
        RECT 355.950 464.400 373.050 465.600 ;
        RECT 355.950 463.950 358.050 464.400 ;
        RECT 370.950 463.950 373.050 464.400 ;
        RECT 415.950 465.600 418.050 466.050 ;
        RECT 436.950 465.600 439.050 466.050 ;
        RECT 415.950 464.400 439.050 465.600 ;
        RECT 415.950 463.950 418.050 464.400 ;
        RECT 436.950 463.950 439.050 464.400 ;
        RECT 550.950 465.600 553.050 466.050 ;
        RECT 559.950 465.600 562.050 466.050 ;
        RECT 550.950 464.400 562.050 465.600 ;
        RECT 550.950 463.950 553.050 464.400 ;
        RECT 559.950 463.950 562.050 464.400 ;
        RECT 748.950 465.600 751.050 466.050 ;
        RECT 781.950 465.600 784.050 466.050 ;
        RECT 748.950 464.400 784.050 465.600 ;
        RECT 748.950 463.950 751.050 464.400 ;
        RECT 781.950 463.950 784.050 464.400 ;
        RECT 829.950 465.600 832.050 466.050 ;
        RECT 844.950 465.600 847.050 466.050 ;
        RECT 850.950 465.600 853.050 466.050 ;
        RECT 829.950 464.400 853.050 465.600 ;
        RECT 829.950 463.950 832.050 464.400 ;
        RECT 844.950 463.950 847.050 464.400 ;
        RECT 850.950 463.950 853.050 464.400 ;
        RECT 874.950 465.600 877.050 466.050 ;
        RECT 889.950 465.600 892.050 466.050 ;
        RECT 874.950 464.400 892.050 465.600 ;
        RECT 874.950 463.950 877.050 464.400 ;
        RECT 889.950 463.950 892.050 464.400 ;
        RECT 283.950 462.600 286.050 463.050 ;
        RECT 319.950 462.600 322.050 463.050 ;
        RECT 283.950 461.400 322.050 462.600 ;
        RECT 283.950 460.950 286.050 461.400 ;
        RECT 319.950 460.950 322.050 461.400 ;
        RECT 496.950 462.600 499.050 463.050 ;
        RECT 505.950 462.600 508.050 463.050 ;
        RECT 496.950 461.400 508.050 462.600 ;
        RECT 496.950 460.950 499.050 461.400 ;
        RECT 505.950 460.950 508.050 461.400 ;
        RECT 538.950 462.600 541.050 463.050 ;
        RECT 568.950 462.600 571.050 463.050 ;
        RECT 676.950 462.600 679.050 463.050 ;
        RECT 697.800 462.600 699.900 463.050 ;
        RECT 538.950 461.400 699.900 462.600 ;
        RECT 538.950 460.950 541.050 461.400 ;
        RECT 568.950 460.950 571.050 461.400 ;
        RECT 676.950 460.950 679.050 461.400 ;
        RECT 697.800 460.950 699.900 461.400 ;
        RECT 700.950 462.600 703.050 463.050 ;
        RECT 727.950 462.600 730.050 463.050 ;
        RECT 778.950 462.600 781.050 463.050 ;
        RECT 700.950 461.400 781.050 462.600 ;
        RECT 700.950 460.950 703.050 461.400 ;
        RECT 727.950 460.950 730.050 461.400 ;
        RECT 778.950 460.950 781.050 461.400 ;
        RECT 808.950 462.600 811.050 463.050 ;
        RECT 817.950 462.600 820.050 463.050 ;
        RECT 808.950 461.400 820.050 462.600 ;
        RECT 808.950 460.950 811.050 461.400 ;
        RECT 817.950 460.950 820.050 461.400 ;
        RECT 847.950 462.600 850.050 463.050 ;
        RECT 871.950 462.600 874.050 463.050 ;
        RECT 880.950 462.600 883.050 463.050 ;
        RECT 847.950 461.400 883.050 462.600 ;
        RECT 847.950 460.950 850.050 461.400 ;
        RECT 871.950 460.950 874.050 461.400 ;
        RECT 880.950 460.950 883.050 461.400 ;
        RECT 136.950 459.600 139.050 460.050 ;
        RECT 145.950 459.600 148.050 460.050 ;
        RECT 136.950 458.400 148.050 459.600 ;
        RECT 136.950 457.950 139.050 458.400 ;
        RECT 145.950 457.950 148.050 458.400 ;
        RECT 208.950 459.600 211.050 460.050 ;
        RECT 220.950 459.600 223.050 460.050 ;
        RECT 331.950 459.600 334.050 460.050 ;
        RECT 208.950 458.400 223.050 459.600 ;
        RECT 208.950 457.950 211.050 458.400 ;
        RECT 220.950 457.950 223.050 458.400 ;
        RECT 323.400 458.400 334.050 459.600 ;
        RECT 4.950 456.600 7.050 457.050 ;
        RECT 22.950 456.600 25.050 457.050 ;
        RECT 4.950 455.400 25.050 456.600 ;
        RECT 4.950 454.950 7.050 455.400 ;
        RECT 22.950 454.950 25.050 455.400 ;
        RECT 154.950 456.600 157.050 457.050 ;
        RECT 199.950 456.600 202.050 457.050 ;
        RECT 154.950 455.400 202.050 456.600 ;
        RECT 154.950 454.950 157.050 455.400 ;
        RECT 199.950 454.950 202.050 455.400 ;
        RECT 301.950 456.600 304.050 457.050 ;
        RECT 323.400 456.600 324.600 458.400 ;
        RECT 331.950 457.950 334.050 458.400 ;
        RECT 502.950 459.600 505.050 460.050 ;
        RECT 529.950 459.600 532.050 460.050 ;
        RECT 502.950 458.400 532.050 459.600 ;
        RECT 502.950 457.950 505.050 458.400 ;
        RECT 529.950 457.950 532.050 458.400 ;
        RECT 541.950 459.600 544.050 460.050 ;
        RECT 556.950 459.600 559.050 460.050 ;
        RECT 541.950 458.400 559.050 459.600 ;
        RECT 541.950 457.950 544.050 458.400 ;
        RECT 556.950 457.950 559.050 458.400 ;
        RECT 610.950 459.600 613.050 460.050 ;
        RECT 658.950 459.600 661.050 460.050 ;
        RECT 610.950 458.400 661.050 459.600 ;
        RECT 610.950 457.950 613.050 458.400 ;
        RECT 658.950 457.950 661.050 458.400 ;
        RECT 736.950 459.600 739.050 460.050 ;
        RECT 742.950 459.600 745.050 460.050 ;
        RECT 736.950 458.400 745.050 459.600 ;
        RECT 736.950 457.950 739.050 458.400 ;
        RECT 742.950 457.950 745.050 458.400 ;
        RECT 757.950 459.600 760.050 460.050 ;
        RECT 805.950 459.600 808.050 460.050 ;
        RECT 757.950 458.400 808.050 459.600 ;
        RECT 757.950 457.950 760.050 458.400 ;
        RECT 805.950 457.950 808.050 458.400 ;
        RECT 823.950 459.600 826.050 460.050 ;
        RECT 832.950 459.600 835.050 460.050 ;
        RECT 823.950 458.400 835.050 459.600 ;
        RECT 823.950 457.950 826.050 458.400 ;
        RECT 832.950 457.950 835.050 458.400 ;
        RECT 301.950 455.400 324.600 456.600 ;
        RECT 349.950 456.600 352.050 457.050 ;
        RECT 361.950 456.600 364.050 457.050 ;
        RECT 349.950 455.400 364.050 456.600 ;
        RECT 301.950 454.950 304.050 455.400 ;
        RECT 349.950 454.950 352.050 455.400 ;
        RECT 361.950 454.950 364.050 455.400 ;
        RECT 421.950 456.600 424.050 457.050 ;
        RECT 460.950 456.600 463.050 457.050 ;
        RECT 475.950 456.600 478.050 457.050 ;
        RECT 481.950 456.600 484.050 457.050 ;
        RECT 421.950 455.400 484.050 456.600 ;
        RECT 421.950 454.950 424.050 455.400 ;
        RECT 460.950 454.950 463.050 455.400 ;
        RECT 475.950 454.950 478.050 455.400 ;
        RECT 481.950 454.950 484.050 455.400 ;
        RECT 496.950 456.600 499.050 457.050 ;
        RECT 607.950 456.600 610.050 457.050 ;
        RECT 496.950 455.400 610.050 456.600 ;
        RECT 496.950 454.950 499.050 455.400 ;
        RECT 607.950 454.950 610.050 455.400 ;
        RECT 664.950 456.600 667.050 457.050 ;
        RECT 676.950 456.600 679.050 457.050 ;
        RECT 820.800 456.600 822.900 457.050 ;
        RECT 664.950 455.400 679.050 456.600 ;
        RECT 664.950 454.950 667.050 455.400 ;
        RECT 676.950 454.950 679.050 455.400 ;
        RECT 770.400 455.400 822.900 456.600 ;
        RECT 55.950 453.600 58.050 454.050 ;
        RECT 64.950 453.600 67.050 454.050 ;
        RECT 55.950 452.400 67.050 453.600 ;
        RECT 55.950 451.950 58.050 452.400 ;
        RECT 64.950 451.950 67.050 452.400 ;
        RECT 76.950 453.600 79.050 454.050 ;
        RECT 85.950 453.600 88.050 454.050 ;
        RECT 76.950 452.400 88.050 453.600 ;
        RECT 76.950 451.950 79.050 452.400 ;
        RECT 85.950 451.950 88.050 452.400 ;
        RECT 214.950 453.600 217.050 454.050 ;
        RECT 241.950 453.600 244.050 454.050 ;
        RECT 247.950 453.600 250.050 454.050 ;
        RECT 271.950 453.600 274.050 454.050 ;
        RECT 334.950 453.600 337.050 454.050 ;
        RECT 214.950 452.400 274.050 453.600 ;
        RECT 214.950 451.950 217.050 452.400 ;
        RECT 241.950 451.950 244.050 452.400 ;
        RECT 247.950 451.950 250.050 452.400 ;
        RECT 271.950 451.950 274.050 452.400 ;
        RECT 329.400 452.400 337.050 453.600 ;
        RECT 13.950 451.050 16.050 451.500 ;
        RECT 19.950 451.050 22.050 451.500 ;
        RECT 13.950 449.850 22.050 451.050 ;
        RECT 13.950 449.400 16.050 449.850 ;
        RECT 19.950 449.400 22.050 449.850 ;
        RECT 49.950 449.100 52.050 451.200 ;
        RECT 67.950 450.600 70.050 451.050 ;
        RECT 73.950 450.600 76.050 451.200 ;
        RECT 67.950 449.400 76.050 450.600 ;
        RECT 31.950 444.150 34.050 444.600 ;
        RECT 40.950 444.150 43.050 444.600 ;
        RECT 31.950 442.950 43.050 444.150 ;
        RECT 31.950 442.500 34.050 442.950 ;
        RECT 40.950 442.500 43.050 442.950 ;
        RECT 50.400 442.050 51.600 449.100 ;
        RECT 67.950 448.950 70.050 449.400 ;
        RECT 73.950 449.100 76.050 449.400 ;
        RECT 142.950 450.750 145.050 451.200 ;
        RECT 154.950 450.750 157.050 451.200 ;
        RECT 142.950 449.550 157.050 450.750 ;
        RECT 142.950 449.100 145.050 449.550 ;
        RECT 154.950 449.100 157.050 449.550 ;
        RECT 184.950 450.750 187.050 451.200 ;
        RECT 193.950 450.750 196.050 451.200 ;
        RECT 184.950 449.550 196.050 450.750 ;
        RECT 214.950 450.600 217.050 451.200 ;
        RECT 184.950 449.100 187.050 449.550 ;
        RECT 193.950 449.100 196.050 449.550 ;
        RECT 203.400 449.400 217.050 450.600 ;
        RECT 58.950 444.450 61.050 444.900 ;
        RECT 67.950 444.450 70.050 444.900 ;
        RECT 58.950 443.250 70.050 444.450 ;
        RECT 58.950 442.800 61.050 443.250 ;
        RECT 67.950 442.800 70.050 443.250 ;
        RECT 139.950 444.450 142.050 444.900 ;
        RECT 151.950 444.450 154.050 445.050 ;
        RECT 203.400 444.900 204.600 449.400 ;
        RECT 214.950 449.100 217.050 449.400 ;
        RECT 226.950 448.950 229.050 451.050 ;
        RECT 277.950 450.750 280.050 451.200 ;
        RECT 295.950 450.750 298.050 451.200 ;
        RECT 277.950 449.550 298.050 450.750 ;
        RECT 277.950 449.100 280.050 449.550 ;
        RECT 295.950 449.100 298.050 449.550 ;
        RECT 304.950 449.400 307.050 451.500 ;
        RECT 227.400 445.050 228.600 448.950 ;
        RECT 157.950 444.450 160.050 444.900 ;
        RECT 139.950 443.250 160.050 444.450 ;
        RECT 139.950 442.800 142.050 443.250 ;
        RECT 151.950 442.950 154.050 443.250 ;
        RECT 157.950 442.800 160.050 443.250 ;
        RECT 202.950 442.800 205.050 444.900 ;
        RECT 226.950 442.950 229.050 445.050 ;
        RECT 238.950 444.600 241.050 445.050 ;
        RECT 283.950 444.600 286.050 445.050 ;
        RECT 238.950 443.400 286.050 444.600 ;
        RECT 305.400 444.600 306.600 449.400 ;
        RECT 329.400 445.050 330.600 452.400 ;
        RECT 334.950 451.950 337.050 452.400 ;
        RECT 400.950 453.600 403.050 454.050 ;
        RECT 409.950 453.600 412.050 454.050 ;
        RECT 400.950 452.400 412.050 453.600 ;
        RECT 400.950 451.950 403.050 452.400 ;
        RECT 409.950 451.950 412.050 452.400 ;
        RECT 544.950 453.600 547.050 454.050 ;
        RECT 586.950 453.600 589.050 454.050 ;
        RECT 544.950 452.400 589.050 453.600 ;
        RECT 544.950 451.950 547.050 452.400 ;
        RECT 586.950 451.950 589.050 452.400 ;
        RECT 355.950 449.100 358.050 451.200 ;
        RECT 382.950 450.600 385.050 451.200 ;
        RECT 466.950 450.600 469.050 451.500 ;
        RECT 481.950 450.600 484.050 451.050 ;
        RECT 382.950 449.400 408.600 450.600 ;
        RECT 466.950 449.400 484.050 450.600 ;
        RECT 382.950 449.100 385.050 449.400 ;
        RECT 356.400 447.600 357.600 449.100 ;
        RECT 344.400 446.400 357.600 447.600 ;
        RECT 316.950 444.600 319.050 445.050 ;
        RECT 305.400 443.400 319.050 444.600 ;
        RECT 238.950 442.950 241.050 443.400 ;
        RECT 283.950 442.950 286.050 443.400 ;
        RECT 316.950 442.950 319.050 443.400 ;
        RECT 328.950 442.950 331.050 445.050 ;
        RECT 334.950 444.600 337.050 444.900 ;
        RECT 344.400 444.600 345.600 446.400 ;
        RECT 407.400 445.050 408.600 449.400 ;
        RECT 481.950 448.950 484.050 449.400 ;
        RECT 559.950 450.600 562.050 451.200 ;
        RECT 589.950 450.600 592.050 451.200 ;
        RECT 559.950 449.400 592.050 450.600 ;
        RECT 559.950 449.100 562.050 449.400 ;
        RECT 589.950 449.100 592.050 449.400 ;
        RECT 601.950 450.600 604.050 451.050 ;
        RECT 616.950 450.600 619.050 451.200 ;
        RECT 601.950 449.400 619.050 450.600 ;
        RECT 601.950 448.950 604.050 449.400 ;
        RECT 616.950 449.100 619.050 449.400 ;
        RECT 640.950 450.600 643.050 451.200 ;
        RECT 652.800 450.600 654.900 451.050 ;
        RECT 640.950 449.400 654.900 450.600 ;
        RECT 640.950 449.100 643.050 449.400 ;
        RECT 652.800 448.950 654.900 449.400 ;
        RECT 655.800 450.000 657.900 451.050 ;
        RECT 658.950 450.750 661.050 451.200 ;
        RECT 673.950 450.750 676.050 451.200 ;
        RECT 658.950 450.600 676.050 450.750 ;
        RECT 679.950 450.600 682.050 451.050 ;
        RECT 712.950 450.600 715.050 451.200 ;
        RECT 757.950 450.600 760.050 451.200 ;
        RECT 655.800 448.950 658.050 450.000 ;
        RECT 658.950 449.550 682.050 450.600 ;
        RECT 658.950 449.100 661.050 449.550 ;
        RECT 673.950 449.400 682.050 449.550 ;
        RECT 673.950 449.100 676.050 449.400 ;
        RECT 679.950 448.950 682.050 449.400 ;
        RECT 695.400 449.400 715.050 450.600 ;
        RECT 655.950 447.600 658.050 448.950 ;
        RECT 695.400 447.600 696.600 449.400 ;
        RECT 712.950 449.100 715.050 449.400 ;
        RECT 728.400 449.400 747.600 450.600 ;
        RECT 635.400 447.000 658.050 447.600 ;
        RECT 634.950 446.400 657.450 447.000 ;
        RECT 692.400 446.400 696.600 447.600 ;
        RECT 634.950 445.050 637.050 446.400 ;
        RECT 334.950 443.400 345.600 444.600 ;
        RECT 346.950 444.600 349.050 445.050 ;
        RECT 358.950 444.600 361.050 444.900 ;
        RECT 346.950 443.400 361.050 444.600 ;
        RECT 334.950 442.800 337.050 443.400 ;
        RECT 346.950 442.950 349.050 443.400 ;
        RECT 358.950 442.800 361.050 443.400 ;
        RECT 373.950 444.600 376.050 445.050 ;
        RECT 379.950 444.600 382.050 444.900 ;
        RECT 373.950 443.400 394.050 444.600 ;
        RECT 373.950 442.950 376.050 443.400 ;
        RECT 379.950 442.800 382.050 443.400 ;
        RECT 391.950 442.500 394.050 443.400 ;
        RECT 406.950 442.950 409.050 445.050 ;
        RECT 439.950 444.150 442.050 444.600 ;
        RECT 448.950 444.150 451.050 444.600 ;
        RECT 439.950 442.950 451.050 444.150 ;
        RECT 634.800 444.000 637.050 445.050 ;
        RECT 688.950 444.600 691.050 444.900 ;
        RECT 692.400 444.600 693.600 446.400 ;
        RECT 728.400 445.050 729.600 449.400 ;
        RECT 746.400 447.600 747.600 449.400 ;
        RECT 752.400 449.400 760.050 450.600 ;
        RECT 752.400 447.600 753.600 449.400 ;
        RECT 757.950 449.100 760.050 449.400 ;
        RECT 746.400 446.400 753.600 447.600 ;
        RECT 770.400 445.050 771.600 455.400 ;
        RECT 820.800 454.950 822.900 455.400 ;
        RECT 823.950 456.600 826.050 456.900 ;
        RECT 853.950 456.600 856.050 457.050 ;
        RECT 823.950 455.400 856.050 456.600 ;
        RECT 823.950 454.800 826.050 455.400 ;
        RECT 853.950 454.950 856.050 455.400 ;
        RECT 817.950 453.600 820.050 454.050 ;
        RECT 850.950 453.600 853.050 454.050 ;
        RECT 817.950 452.400 853.050 453.600 ;
        RECT 817.950 451.950 820.050 452.400 ;
        RECT 850.950 451.950 853.050 452.400 ;
        RECT 856.950 453.600 859.050 454.050 ;
        RECT 886.950 453.600 889.050 454.050 ;
        RECT 856.950 452.400 889.050 453.600 ;
        RECT 856.950 451.950 859.050 452.400 ;
        RECT 886.950 451.950 889.050 452.400 ;
        RECT 781.950 448.950 784.050 451.050 ;
        RECT 814.950 450.750 817.050 451.200 ;
        RECT 823.950 450.750 826.050 451.200 ;
        RECT 814.950 449.550 826.050 450.750 ;
        RECT 814.950 449.100 817.050 449.550 ;
        RECT 823.950 449.100 826.050 449.550 ;
        RECT 829.950 450.750 832.050 451.200 ;
        RECT 838.950 450.750 841.050 451.200 ;
        RECT 829.950 449.550 841.050 450.750 ;
        RECT 829.950 449.100 832.050 449.550 ;
        RECT 838.950 449.100 841.050 449.550 ;
        RECT 844.950 450.600 847.050 451.050 ;
        RECT 844.950 449.400 852.600 450.600 ;
        RECT 844.950 448.950 847.050 449.400 ;
        RECT 782.400 445.050 783.600 448.950 ;
        RECT 634.800 442.950 636.900 444.000 ;
        RECT 688.950 443.400 693.600 444.600 ;
        RECT 697.950 444.450 700.050 444.900 ;
        RECT 703.950 444.450 706.050 444.900 ;
        RECT 439.950 442.500 442.050 442.950 ;
        RECT 448.950 442.500 451.050 442.950 ;
        RECT 688.950 442.800 691.050 443.400 ;
        RECT 697.950 443.250 706.050 444.450 ;
        RECT 697.950 442.800 700.050 443.250 ;
        RECT 703.950 442.800 706.050 443.250 ;
        RECT 724.950 443.400 729.600 445.050 ;
        RECT 742.950 444.600 745.050 445.050 ;
        RECT 754.950 444.600 757.050 444.900 ;
        RECT 742.950 443.400 757.050 444.600 ;
        RECT 724.950 442.950 729.000 443.400 ;
        RECT 742.950 442.950 745.050 443.400 ;
        RECT 754.950 442.800 757.050 443.400 ;
        RECT 769.950 442.950 772.050 445.050 ;
        RECT 781.950 442.950 784.050 445.050 ;
        RECT 832.950 444.600 835.050 445.050 ;
        RECT 851.400 444.900 852.600 449.400 ;
        RECT 859.950 448.950 862.050 451.050 ;
        RECT 865.950 450.600 868.050 451.200 ;
        RECT 865.950 449.400 870.600 450.600 ;
        RECT 865.950 449.100 868.050 449.400 ;
        RECT 860.400 445.050 861.600 448.950 ;
        RECT 850.950 444.600 853.050 444.900 ;
        RECT 832.950 443.400 853.050 444.600 ;
        RECT 832.950 442.950 835.050 443.400 ;
        RECT 850.950 442.800 853.050 443.400 ;
        RECT 859.950 442.950 862.050 445.050 ;
        RECT 869.400 444.600 870.600 449.400 ;
        RECT 892.950 448.950 895.050 451.050 ;
        RECT 893.400 445.050 894.600 448.950 ;
        RECT 883.950 444.600 886.050 444.900 ;
        RECT 869.400 443.400 886.050 444.600 ;
        RECT 883.950 442.800 886.050 443.400 ;
        RECT 892.950 442.950 895.050 445.050 ;
        RECT 49.950 439.950 52.050 442.050 ;
        RECT 79.950 441.600 82.050 442.050 ;
        RECT 169.950 441.600 172.050 442.050 ;
        RECT 79.950 440.400 172.050 441.600 ;
        RECT 79.950 439.950 82.050 440.400 ;
        RECT 169.950 439.950 172.050 440.400 ;
        RECT 112.950 438.600 115.050 439.050 ;
        RECT 130.950 438.600 133.050 438.900 ;
        RECT 112.950 437.400 133.050 438.600 ;
        RECT 112.950 436.950 115.050 437.400 ;
        RECT 130.950 436.800 133.050 437.400 ;
        RECT 172.950 438.600 175.050 439.050 ;
        RECT 181.950 438.600 184.050 439.050 ;
        RECT 172.950 437.400 184.050 438.600 ;
        RECT 172.950 436.950 175.050 437.400 ;
        RECT 181.950 436.950 184.050 437.400 ;
        RECT 187.950 438.600 190.050 439.050 ;
        RECT 217.950 438.600 220.050 439.050 ;
        RECT 187.950 437.400 220.050 438.600 ;
        RECT 286.950 438.600 289.050 442.050 ;
        RECT 340.950 441.600 343.050 442.050 ;
        RECT 364.950 441.600 367.050 442.050 ;
        RECT 340.950 440.400 367.050 441.600 ;
        RECT 340.950 439.950 343.050 440.400 ;
        RECT 364.950 439.950 367.050 440.400 ;
        RECT 370.950 441.600 373.050 442.050 ;
        RECT 379.950 441.600 382.050 441.750 ;
        RECT 370.950 440.400 382.050 441.600 ;
        RECT 370.950 439.950 373.050 440.400 ;
        RECT 379.950 439.650 382.050 440.400 ;
        RECT 514.950 441.600 517.050 442.050 ;
        RECT 544.950 441.600 547.050 442.050 ;
        RECT 514.950 440.400 547.050 441.600 ;
        RECT 514.950 439.950 517.050 440.400 ;
        RECT 544.950 439.950 547.050 440.400 ;
        RECT 556.950 441.600 559.050 442.050 ;
        RECT 562.950 441.600 565.050 442.050 ;
        RECT 568.950 441.600 571.050 442.050 ;
        RECT 595.950 441.600 598.050 442.050 ;
        RECT 556.950 440.400 598.050 441.600 ;
        RECT 556.950 439.950 559.050 440.400 ;
        RECT 562.950 439.950 565.050 440.400 ;
        RECT 568.950 439.950 571.050 440.400 ;
        RECT 595.950 439.950 598.050 440.400 ;
        RECT 607.950 441.600 610.050 442.050 ;
        RECT 619.950 441.600 622.050 442.050 ;
        RECT 607.950 440.400 622.050 441.600 ;
        RECT 607.950 439.950 610.050 440.400 ;
        RECT 619.950 439.950 622.050 440.400 ;
        RECT 766.950 441.600 769.050 442.050 ;
        RECT 775.950 441.600 778.050 442.050 ;
        RECT 814.950 441.600 817.050 442.050 ;
        RECT 766.950 440.400 817.050 441.600 ;
        RECT 766.950 439.950 769.050 440.400 ;
        RECT 775.950 439.950 778.050 440.400 ;
        RECT 814.950 439.950 817.050 440.400 ;
        RECT 298.950 438.600 301.050 439.050 ;
        RECT 337.950 438.600 340.050 439.050 ;
        RECT 286.950 438.000 340.050 438.600 ;
        RECT 287.400 437.400 340.050 438.000 ;
        RECT 187.950 436.950 190.050 437.400 ;
        RECT 217.950 436.950 220.050 437.400 ;
        RECT 298.950 436.950 301.050 437.400 ;
        RECT 337.950 436.950 340.050 437.400 ;
        RECT 367.950 438.600 370.050 439.050 ;
        RECT 487.950 438.600 490.050 439.050 ;
        RECT 367.950 437.400 490.050 438.600 ;
        RECT 367.950 436.950 370.050 437.400 ;
        RECT 487.950 436.950 490.050 437.400 ;
        RECT 709.950 438.600 712.050 439.050 ;
        RECT 736.950 438.600 739.050 439.050 ;
        RECT 709.950 437.400 739.050 438.600 ;
        RECT 709.950 436.950 712.050 437.400 ;
        RECT 736.950 436.950 739.050 437.400 ;
        RECT 874.950 438.600 877.050 439.050 ;
        RECT 892.950 438.600 895.050 439.050 ;
        RECT 874.950 437.400 895.050 438.600 ;
        RECT 874.950 436.950 877.050 437.400 ;
        RECT 892.950 436.950 895.050 437.400 ;
        RECT 19.950 435.600 22.050 436.050 ;
        RECT 52.950 435.600 55.050 436.050 ;
        RECT 19.950 434.400 55.050 435.600 ;
        RECT 19.950 433.950 22.050 434.400 ;
        RECT 52.950 433.950 55.050 434.400 ;
        RECT 184.950 435.600 187.050 436.050 ;
        RECT 274.950 435.600 277.050 436.050 ;
        RECT 184.950 434.400 277.050 435.600 ;
        RECT 184.950 433.950 187.050 434.400 ;
        RECT 274.950 433.950 277.050 434.400 ;
        RECT 319.950 435.600 322.050 436.050 ;
        RECT 358.950 435.600 361.050 436.050 ;
        RECT 319.950 434.400 361.050 435.600 ;
        RECT 319.950 433.950 322.050 434.400 ;
        RECT 358.950 433.950 361.050 434.400 ;
        RECT 520.950 435.600 523.050 436.050 ;
        RECT 538.950 435.600 541.050 436.050 ;
        RECT 520.950 434.400 541.050 435.600 ;
        RECT 520.950 433.950 523.050 434.400 ;
        RECT 538.950 433.950 541.050 434.400 ;
        RECT 688.950 435.600 691.050 436.050 ;
        RECT 790.950 435.600 793.050 436.050 ;
        RECT 688.950 434.400 793.050 435.600 ;
        RECT 688.950 433.950 691.050 434.400 ;
        RECT 790.950 433.950 793.050 434.400 ;
        RECT 820.950 435.600 823.050 436.050 ;
        RECT 832.800 435.600 834.900 436.050 ;
        RECT 820.950 434.400 834.900 435.600 ;
        RECT 820.950 433.950 823.050 434.400 ;
        RECT 832.800 433.950 834.900 434.400 ;
        RECT 835.950 435.600 838.050 436.050 ;
        RECT 871.950 435.600 874.050 436.050 ;
        RECT 835.950 434.400 874.050 435.600 ;
        RECT 835.950 433.950 838.050 434.400 ;
        RECT 871.950 433.950 874.050 434.400 ;
        RECT 97.950 432.600 100.050 433.050 ;
        RECT 145.950 432.600 148.050 433.050 ;
        RECT 181.950 432.600 184.050 433.050 ;
        RECT 97.950 431.400 184.050 432.600 ;
        RECT 97.950 430.950 100.050 431.400 ;
        RECT 145.950 430.950 148.050 431.400 ;
        RECT 181.950 430.950 184.050 431.400 ;
        RECT 295.950 432.600 298.050 433.050 ;
        RECT 373.950 432.600 376.050 433.050 ;
        RECT 295.950 431.400 376.050 432.600 ;
        RECT 295.950 430.950 298.050 431.400 ;
        RECT 373.950 430.950 376.050 431.400 ;
        RECT 760.950 432.600 763.050 433.050 ;
        RECT 778.950 432.600 781.050 433.050 ;
        RECT 880.950 432.600 883.050 433.050 ;
        RECT 760.950 431.400 781.050 432.600 ;
        RECT 760.950 430.950 763.050 431.400 ;
        RECT 778.950 430.950 781.050 431.400 ;
        RECT 845.400 431.400 883.050 432.600 ;
        RECT 845.400 430.050 846.600 431.400 ;
        RECT 880.950 430.950 883.050 431.400 ;
        RECT 208.950 429.600 211.050 430.050 ;
        RECT 235.950 429.600 238.050 430.050 ;
        RECT 208.950 428.400 238.050 429.600 ;
        RECT 208.950 427.950 211.050 428.400 ;
        RECT 235.950 427.950 238.050 428.400 ;
        RECT 265.950 429.600 268.050 430.050 ;
        RECT 295.950 429.600 298.050 429.900 ;
        RECT 265.950 428.400 298.050 429.600 ;
        RECT 265.950 427.950 268.050 428.400 ;
        RECT 295.950 427.800 298.050 428.400 ;
        RECT 385.950 429.600 388.050 430.050 ;
        RECT 424.950 429.600 427.050 430.050 ;
        RECT 457.950 429.600 460.050 430.050 ;
        RECT 508.950 429.600 511.050 430.050 ;
        RECT 385.950 428.400 447.600 429.600 ;
        RECT 385.950 427.950 388.050 428.400 ;
        RECT 424.950 427.950 427.050 428.400 ;
        RECT 100.950 426.600 103.050 427.050 ;
        RECT 109.950 426.600 112.050 427.050 ;
        RECT 100.950 425.400 112.050 426.600 ;
        RECT 100.950 424.950 103.050 425.400 ;
        RECT 109.950 424.950 112.050 425.400 ;
        RECT 241.950 426.600 244.050 427.050 ;
        RECT 259.950 426.600 262.050 427.050 ;
        RECT 241.950 425.400 262.050 426.600 ;
        RECT 241.950 424.950 244.050 425.400 ;
        RECT 259.950 424.950 262.050 425.400 ;
        RECT 424.950 426.600 427.050 426.900 ;
        RECT 442.950 426.600 445.050 427.050 ;
        RECT 424.950 425.400 445.050 426.600 ;
        RECT 446.400 426.600 447.600 428.400 ;
        RECT 457.950 428.400 511.050 429.600 ;
        RECT 457.950 427.950 460.050 428.400 ;
        RECT 508.950 427.950 511.050 428.400 ;
        RECT 574.950 429.600 577.050 430.050 ;
        RECT 613.950 429.600 616.050 430.050 ;
        RECT 619.800 429.600 621.900 430.050 ;
        RECT 574.950 428.400 621.900 429.600 ;
        RECT 574.950 427.950 577.050 428.400 ;
        RECT 613.950 427.950 616.050 428.400 ;
        RECT 619.800 427.950 621.900 428.400 ;
        RECT 622.950 429.600 625.050 430.050 ;
        RECT 655.950 429.600 658.050 430.050 ;
        RECT 622.950 428.400 658.050 429.600 ;
        RECT 622.950 427.950 625.050 428.400 ;
        RECT 655.950 427.950 658.050 428.400 ;
        RECT 715.950 429.600 718.050 430.050 ;
        RECT 739.950 429.600 742.050 430.050 ;
        RECT 715.950 428.400 742.050 429.600 ;
        RECT 715.950 427.950 718.050 428.400 ;
        RECT 739.950 427.950 742.050 428.400 ;
        RECT 745.950 429.600 748.050 430.050 ;
        RECT 763.950 429.600 766.050 430.050 ;
        RECT 745.950 428.400 766.050 429.600 ;
        RECT 745.950 427.950 748.050 428.400 ;
        RECT 763.950 427.950 766.050 428.400 ;
        RECT 799.950 429.600 802.050 430.050 ;
        RECT 805.950 429.600 808.050 430.050 ;
        RECT 844.950 429.600 847.050 430.050 ;
        RECT 799.950 428.400 847.050 429.600 ;
        RECT 799.950 427.950 802.050 428.400 ;
        RECT 805.950 427.950 808.050 428.400 ;
        RECT 844.950 427.950 847.050 428.400 ;
        RECT 853.950 429.600 856.050 430.050 ;
        RECT 895.950 429.600 898.050 430.050 ;
        RECT 853.950 428.400 898.050 429.600 ;
        RECT 853.950 427.950 856.050 428.400 ;
        RECT 895.950 427.950 898.050 428.400 ;
        RECT 469.950 426.600 472.050 427.050 ;
        RECT 446.400 425.400 472.050 426.600 ;
        RECT 424.950 424.800 427.050 425.400 ;
        RECT 442.950 424.950 445.050 425.400 ;
        RECT 469.950 424.950 472.050 425.400 ;
        RECT 481.950 426.600 484.050 427.050 ;
        RECT 520.950 426.600 523.050 427.050 ;
        RECT 481.950 425.400 523.050 426.600 ;
        RECT 481.950 424.950 484.050 425.400 ;
        RECT 520.950 424.950 523.050 425.400 ;
        RECT 544.950 426.600 547.050 427.050 ;
        RECT 571.950 426.600 574.050 427.050 ;
        RECT 544.950 425.400 574.050 426.600 ;
        RECT 544.950 424.950 547.050 425.400 ;
        RECT 571.950 424.950 574.050 425.400 ;
        RECT 679.950 426.600 682.050 427.050 ;
        RECT 718.950 426.600 721.050 427.050 ;
        RECT 724.950 426.600 727.050 427.050 ;
        RECT 679.950 425.400 727.050 426.600 ;
        RECT 679.950 424.950 682.050 425.400 ;
        RECT 718.950 424.950 721.050 425.400 ;
        RECT 724.950 424.950 727.050 425.400 ;
        RECT 826.950 426.600 829.050 427.050 ;
        RECT 838.950 426.600 841.050 427.050 ;
        RECT 826.950 425.400 841.050 426.600 ;
        RECT 826.950 424.950 829.050 425.400 ;
        RECT 838.950 424.950 841.050 425.400 ;
        RECT 19.950 423.600 22.050 424.050 ;
        RECT 73.950 423.600 76.050 424.050 ;
        RECT 19.950 422.400 76.050 423.600 ;
        RECT 19.950 421.950 22.050 422.400 ;
        RECT 73.950 421.950 76.050 422.400 ;
        RECT 82.950 423.600 85.050 424.050 ;
        RECT 106.950 423.600 109.050 424.050 ;
        RECT 82.950 422.400 109.050 423.600 ;
        RECT 82.950 421.950 85.050 422.400 ;
        RECT 106.950 421.950 109.050 422.400 ;
        RECT 148.950 423.600 151.050 424.050 ;
        RECT 196.950 423.600 199.050 424.050 ;
        RECT 148.950 422.400 199.050 423.600 ;
        RECT 148.950 421.950 151.050 422.400 ;
        RECT 196.950 421.950 199.050 422.400 ;
        RECT 304.950 423.600 307.050 424.050 ;
        RECT 349.950 423.600 352.050 424.050 ;
        RECT 304.950 422.400 352.050 423.600 ;
        RECT 304.950 421.950 307.050 422.400 ;
        RECT 349.950 421.950 352.050 422.400 ;
        RECT 364.950 423.600 367.050 424.050 ;
        RECT 385.950 423.600 388.050 424.050 ;
        RECT 364.950 422.400 388.050 423.600 ;
        RECT 364.950 421.950 367.050 422.400 ;
        RECT 385.950 421.950 388.050 422.400 ;
        RECT 439.950 423.600 442.050 424.050 ;
        RECT 502.950 423.600 505.050 424.050 ;
        RECT 439.950 422.400 505.050 423.600 ;
        RECT 439.950 421.950 442.050 422.400 ;
        RECT 502.950 421.950 505.050 422.400 ;
        RECT 523.950 423.600 526.050 424.050 ;
        RECT 628.950 423.600 631.050 424.050 ;
        RECT 523.950 422.400 631.050 423.600 ;
        RECT 523.950 421.950 526.050 422.400 ;
        RECT 628.950 421.950 631.050 422.400 ;
        RECT 652.950 423.600 655.050 424.050 ;
        RECT 661.950 423.600 664.050 424.050 ;
        RECT 652.950 422.400 664.050 423.600 ;
        RECT 652.950 421.950 655.050 422.400 ;
        RECT 661.950 421.950 664.050 422.400 ;
        RECT 673.950 423.600 676.050 424.050 ;
        RECT 688.950 423.600 691.050 424.050 ;
        RECT 673.950 422.400 691.050 423.600 ;
        RECT 673.950 421.950 676.050 422.400 ;
        RECT 688.950 421.950 691.050 422.400 ;
        RECT 751.950 423.600 754.050 424.050 ;
        RECT 808.950 423.600 811.050 424.050 ;
        RECT 751.950 422.400 811.050 423.600 ;
        RECT 751.950 421.950 754.050 422.400 ;
        RECT 808.950 421.950 811.050 422.400 ;
        RECT 814.950 423.600 817.050 424.050 ;
        RECT 841.950 423.600 844.050 424.050 ;
        RECT 814.950 422.400 844.050 423.600 ;
        RECT 814.950 421.950 817.050 422.400 ;
        RECT 841.950 421.950 844.050 422.400 ;
        RECT 850.950 423.600 853.050 424.050 ;
        RECT 859.950 423.600 862.050 424.050 ;
        RECT 850.950 422.400 862.050 423.600 ;
        RECT 850.950 421.950 853.050 422.400 ;
        RECT 859.950 421.950 862.050 422.400 ;
        RECT 886.950 423.600 889.050 424.050 ;
        RECT 886.950 422.400 900.600 423.600 ;
        RECT 886.950 421.950 889.050 422.400 ;
        RECT 88.950 420.600 91.050 421.050 ;
        RECT 103.950 420.600 106.050 421.050 ;
        RECT 88.950 419.400 106.050 420.600 ;
        RECT 88.950 418.950 91.050 419.400 ;
        RECT 103.950 418.950 106.050 419.400 ;
        RECT 328.950 420.600 331.050 421.050 ;
        RECT 334.950 420.600 337.050 421.050 ;
        RECT 328.950 419.400 337.050 420.600 ;
        RECT 328.950 418.950 331.050 419.400 ;
        RECT 334.950 418.950 337.050 419.400 ;
        RECT 379.950 420.600 382.050 421.050 ;
        RECT 391.950 420.600 394.050 421.050 ;
        RECT 379.950 419.400 394.050 420.600 ;
        RECT 379.950 418.950 382.050 419.400 ;
        RECT 391.950 418.950 394.050 419.400 ;
        RECT 445.950 420.600 448.050 421.050 ;
        RECT 481.950 420.600 484.050 421.050 ;
        RECT 490.950 420.600 493.050 421.050 ;
        RECT 445.950 419.400 493.050 420.600 ;
        RECT 445.950 418.950 448.050 419.400 ;
        RECT 481.950 418.950 484.050 419.400 ;
        RECT 490.950 418.950 493.050 419.400 ;
        RECT 592.950 420.600 597.000 421.050 ;
        RECT 610.950 420.600 613.050 421.050 ;
        RECT 616.950 420.600 619.050 421.050 ;
        RECT 592.950 418.950 597.600 420.600 ;
        RECT 610.950 419.400 619.050 420.600 ;
        RECT 610.950 418.950 613.050 419.400 ;
        RECT 616.950 418.950 619.050 419.400 ;
        RECT 730.950 420.600 733.050 421.050 ;
        RECT 739.950 420.600 742.050 421.050 ;
        RECT 730.950 419.400 742.050 420.600 ;
        RECT 730.950 418.950 733.050 419.400 ;
        RECT 739.950 418.950 742.050 419.400 ;
        RECT 757.950 420.600 760.050 421.050 ;
        RECT 772.800 420.600 774.900 421.050 ;
        RECT 757.950 419.400 774.900 420.600 ;
        RECT 757.950 418.950 760.050 419.400 ;
        RECT 772.800 418.950 774.900 419.400 ;
        RECT 775.950 420.600 778.050 421.050 ;
        RECT 826.950 420.600 829.050 421.050 ;
        RECT 856.950 420.600 859.050 421.050 ;
        RECT 775.950 419.400 789.600 420.600 ;
        RECT 775.950 418.950 778.050 419.400 ;
        RECT 31.950 416.400 34.050 418.500 ;
        RECT 91.950 417.600 94.050 418.050 ;
        RECT 97.950 417.600 100.050 418.200 ;
        RECT 91.950 416.400 100.050 417.600 ;
        RECT 151.950 418.050 154.050 418.500 ;
        RECT 160.950 418.050 163.050 418.500 ;
        RECT 151.950 416.850 163.050 418.050 ;
        RECT 151.950 416.400 154.050 416.850 ;
        RECT 160.950 416.400 163.050 416.850 ;
        RECT 196.950 417.750 199.050 418.200 ;
        RECT 202.950 417.750 205.050 418.200 ;
        RECT 196.950 416.550 205.050 417.750 ;
        RECT 32.400 414.600 33.600 416.400 ;
        RECT 91.950 415.950 94.050 416.400 ;
        RECT 97.950 416.100 100.050 416.400 ;
        RECT 196.950 416.100 199.050 416.550 ;
        RECT 202.950 416.100 205.050 416.550 ;
        RECT 208.950 417.600 211.050 418.200 ;
        RECT 214.800 417.600 216.900 418.050 ;
        RECT 208.950 416.400 216.900 417.600 ;
        RECT 208.950 416.100 211.050 416.400 ;
        RECT 214.800 415.950 216.900 416.400 ;
        RECT 217.950 417.600 220.050 418.050 ;
        RECT 226.950 417.600 229.050 418.200 ;
        RECT 217.950 416.400 229.050 417.600 ;
        RECT 217.950 415.950 220.050 416.400 ;
        RECT 226.950 416.100 229.050 416.400 ;
        RECT 232.950 417.750 235.050 418.200 ;
        RECT 244.950 417.750 247.050 418.200 ;
        RECT 232.950 416.550 247.050 417.750 ;
        RECT 232.950 416.100 235.050 416.550 ;
        RECT 244.950 416.100 247.050 416.550 ;
        RECT 250.950 416.400 253.050 418.500 ;
        RECT 307.950 417.750 310.050 418.200 ;
        RECT 313.950 417.750 316.050 418.200 ;
        RECT 307.950 416.550 316.050 417.750 ;
        RECT 346.950 417.600 349.050 418.200 ;
        RECT 112.950 414.600 115.050 415.050 ;
        RECT 32.400 413.400 115.050 414.600 ;
        RECT 112.950 412.950 115.050 413.400 ;
        RECT 40.950 411.600 43.050 412.050 ;
        RECT 46.950 411.600 49.050 411.900 ;
        RECT 13.950 411.150 16.050 411.600 ;
        RECT 19.950 411.150 22.050 411.600 ;
        RECT 13.950 409.950 22.050 411.150 ;
        RECT 40.950 410.400 49.050 411.600 ;
        RECT 40.950 409.950 43.050 410.400 ;
        RECT 13.950 409.500 16.050 409.950 ;
        RECT 19.950 409.500 22.050 409.950 ;
        RECT 46.950 409.800 49.050 410.400 ;
        RECT 52.950 411.450 55.050 411.900 ;
        RECT 58.800 411.450 60.900 411.900 ;
        RECT 52.950 410.250 60.900 411.450 ;
        RECT 52.950 409.800 55.050 410.250 ;
        RECT 58.800 409.800 60.900 410.250 ;
        RECT 61.950 411.450 64.050 411.900 ;
        RECT 70.950 411.450 73.050 411.900 ;
        RECT 61.950 410.250 73.050 411.450 ;
        RECT 61.950 409.800 64.050 410.250 ;
        RECT 70.950 409.800 73.050 410.250 ;
        RECT 76.950 411.450 79.050 411.900 ;
        RECT 82.950 411.450 85.050 411.900 ;
        RECT 76.950 410.250 85.050 411.450 ;
        RECT 76.950 409.800 79.050 410.250 ;
        RECT 82.950 409.800 85.050 410.250 ;
        RECT 100.950 411.450 103.050 411.900 ;
        RECT 109.950 411.450 112.050 411.900 ;
        RECT 148.950 411.600 151.050 412.050 ;
        RECT 100.950 410.250 112.050 411.450 ;
        RECT 100.950 409.800 103.050 410.250 ;
        RECT 109.950 409.800 112.050 410.250 ;
        RECT 142.950 410.400 151.050 411.600 ;
        RECT 142.950 409.500 145.050 410.400 ;
        RECT 148.950 409.950 151.050 410.400 ;
        RECT 163.950 411.450 166.050 411.900 ;
        RECT 178.950 411.450 181.050 411.900 ;
        RECT 163.950 410.250 181.050 411.450 ;
        RECT 163.950 409.800 166.050 410.250 ;
        RECT 178.950 409.800 181.050 410.250 ;
        RECT 184.950 411.600 187.050 411.900 ;
        RECT 196.950 411.600 199.050 412.050 ;
        RECT 223.950 411.600 226.050 411.900 ;
        RECT 184.950 410.400 226.050 411.600 ;
        RECT 184.950 409.800 187.050 410.400 ;
        RECT 196.950 409.950 199.050 410.400 ;
        RECT 223.950 409.800 226.050 410.400 ;
        RECT 238.950 411.600 241.050 412.050 ;
        RECT 251.400 411.600 252.600 416.400 ;
        RECT 307.950 416.100 310.050 416.550 ;
        RECT 313.950 416.100 316.050 416.550 ;
        RECT 323.400 416.400 349.050 417.600 ;
        RECT 323.400 411.900 324.600 416.400 ;
        RECT 346.950 416.100 349.050 416.400 ;
        RECT 352.950 416.100 355.050 418.200 ;
        RECT 370.950 417.600 373.050 418.200 ;
        RECT 382.950 417.600 385.050 418.050 ;
        RECT 370.950 416.400 385.050 417.600 ;
        RECT 370.950 416.100 373.050 416.400 ;
        RECT 238.950 410.400 252.600 411.600 ;
        RECT 262.950 411.150 265.050 411.600 ;
        RECT 277.950 411.150 280.050 411.600 ;
        RECT 238.950 409.950 241.050 410.400 ;
        RECT 262.950 409.950 280.050 411.150 ;
        RECT 262.950 409.500 265.050 409.950 ;
        RECT 277.950 409.500 280.050 409.950 ;
        RECT 304.950 411.450 307.050 411.900 ;
        RECT 316.950 411.450 319.050 411.900 ;
        RECT 304.950 410.250 319.050 411.450 ;
        RECT 304.950 409.800 307.050 410.250 ;
        RECT 316.950 409.800 319.050 410.250 ;
        RECT 322.950 409.800 325.050 411.900 ;
        RECT 337.950 411.600 340.050 412.050 ;
        RECT 343.950 411.600 346.050 411.900 ;
        RECT 337.950 410.400 346.050 411.600 ;
        RECT 353.400 411.600 354.600 416.100 ;
        RECT 382.950 415.950 385.050 416.400 ;
        RECT 409.950 417.600 412.050 418.050 ;
        RECT 418.950 417.600 421.050 418.200 ;
        RECT 457.950 418.050 460.050 418.500 ;
        RECT 463.950 418.050 466.050 418.500 ;
        RECT 427.950 417.600 430.050 418.050 ;
        RECT 409.950 416.400 421.050 417.600 ;
        RECT 409.950 415.950 412.050 416.400 ;
        RECT 418.950 416.100 421.050 416.400 ;
        RECT 422.400 416.400 430.050 417.600 ;
        RECT 422.400 411.900 423.600 416.400 ;
        RECT 427.950 415.950 430.050 416.400 ;
        RECT 442.950 417.600 445.050 418.050 ;
        RECT 448.950 417.600 451.050 418.050 ;
        RECT 442.950 416.400 451.050 417.600 ;
        RECT 457.950 416.850 466.050 418.050 ;
        RECT 457.950 416.400 460.050 416.850 ;
        RECT 463.950 416.400 466.050 416.850 ;
        RECT 496.950 417.600 499.050 418.200 ;
        RECT 502.950 417.600 505.050 418.050 ;
        RECT 496.950 416.400 505.050 417.600 ;
        RECT 442.950 415.950 445.050 416.400 ;
        RECT 448.950 415.950 451.050 416.400 ;
        RECT 496.950 416.100 499.050 416.400 ;
        RECT 502.950 415.950 505.050 416.400 ;
        RECT 526.950 417.600 529.050 418.200 ;
        RECT 532.950 417.600 535.050 418.050 ;
        RECT 526.950 416.400 535.050 417.600 ;
        RECT 526.950 416.100 529.050 416.400 ;
        RECT 532.950 415.950 535.050 416.400 ;
        RECT 538.950 417.600 541.050 418.200 ;
        RECT 553.950 417.600 556.050 418.050 ;
        RECT 538.950 416.400 556.050 417.600 ;
        RECT 538.950 416.100 541.050 416.400 ;
        RECT 553.950 415.950 556.050 416.400 ;
        RECT 568.950 417.750 571.050 418.200 ;
        RECT 574.950 417.750 577.050 418.200 ;
        RECT 568.950 416.550 577.050 417.750 ;
        RECT 568.950 416.100 571.050 416.550 ;
        RECT 574.950 416.100 577.050 416.550 ;
        RECT 580.950 417.600 583.050 418.050 ;
        RECT 589.950 417.600 592.050 418.200 ;
        RECT 580.950 416.400 592.050 417.600 ;
        RECT 580.950 415.950 583.050 416.400 ;
        RECT 589.950 416.100 592.050 416.400 ;
        RECT 596.400 414.600 597.600 418.950 ;
        RECT 604.950 415.950 607.050 418.050 ;
        RECT 619.950 417.750 622.050 418.050 ;
        RECT 634.950 417.750 637.050 418.200 ;
        RECT 619.950 416.550 637.050 417.750 ;
        RECT 619.950 415.950 622.050 416.550 ;
        RECT 634.950 416.100 637.050 416.550 ;
        RECT 679.950 417.600 682.050 418.200 ;
        RECT 685.800 417.600 687.900 418.050 ;
        RECT 679.950 416.400 687.900 417.600 ;
        RECT 679.950 416.100 682.050 416.400 ;
        RECT 685.800 415.950 687.900 416.400 ;
        RECT 688.950 417.750 691.050 418.200 ;
        RECT 697.950 417.750 700.050 418.200 ;
        RECT 688.950 416.550 700.050 417.750 ;
        RECT 688.950 416.100 691.050 416.550 ;
        RECT 697.950 416.100 700.050 416.550 ;
        RECT 703.950 417.750 706.050 418.200 ;
        RECT 712.950 417.750 715.050 418.200 ;
        RECT 703.950 416.550 715.050 417.750 ;
        RECT 703.950 416.100 706.050 416.550 ;
        RECT 712.950 416.100 715.050 416.550 ;
        RECT 721.950 417.600 724.050 418.050 ;
        RECT 742.950 417.600 745.050 418.050 ;
        RECT 721.950 416.400 745.050 417.600 ;
        RECT 721.950 415.950 724.050 416.400 ;
        RECT 742.950 415.950 745.050 416.400 ;
        RECT 760.950 415.950 763.050 418.050 ;
        RECT 596.400 414.000 600.600 414.600 ;
        RECT 596.400 413.400 601.050 414.000 ;
        RECT 388.950 411.600 391.050 411.900 ;
        RECT 353.400 410.400 391.050 411.600 ;
        RECT 337.950 409.950 340.050 410.400 ;
        RECT 343.950 409.800 346.050 410.400 ;
        RECT 388.950 409.800 391.050 410.400 ;
        RECT 394.950 411.450 397.050 411.900 ;
        RECT 406.950 411.450 409.050 411.900 ;
        RECT 394.950 410.250 409.050 411.450 ;
        RECT 394.950 409.800 397.050 410.250 ;
        RECT 406.950 409.800 409.050 410.250 ;
        RECT 421.950 409.800 424.050 411.900 ;
        RECT 469.950 411.600 472.050 412.050 ;
        RECT 475.950 411.600 478.050 411.900 ;
        RECT 469.950 410.400 478.050 411.600 ;
        RECT 469.950 409.950 472.050 410.400 ;
        RECT 475.950 409.800 478.050 410.400 ;
        RECT 508.950 411.450 511.050 411.900 ;
        RECT 523.950 411.450 526.050 411.900 ;
        RECT 508.950 410.250 526.050 411.450 ;
        RECT 508.950 409.800 511.050 410.250 ;
        RECT 523.950 409.800 526.050 410.250 ;
        RECT 541.950 411.450 544.050 411.900 ;
        RECT 556.950 411.450 559.050 411.900 ;
        RECT 541.950 410.250 559.050 411.450 ;
        RECT 541.950 409.800 544.050 410.250 ;
        RECT 556.950 409.800 559.050 410.250 ;
        RECT 598.950 409.950 601.050 413.400 ;
        RECT 605.400 412.050 606.600 415.950 ;
        RECT 680.400 413.400 696.600 414.600 ;
        RECT 604.950 409.950 607.050 412.050 ;
        RECT 670.950 411.600 673.050 411.900 ;
        RECT 680.400 411.600 681.600 413.400 ;
        RECT 695.400 411.900 696.600 413.400 ;
        RECT 761.400 412.050 762.600 415.950 ;
        RECT 766.950 414.600 769.050 418.050 ;
        RECT 788.400 417.600 789.600 419.400 ;
        RECT 826.950 419.400 859.050 420.600 ;
        RECT 826.950 418.950 829.050 419.400 ;
        RECT 856.950 418.950 859.050 419.400 ;
        RECT 820.950 417.600 823.050 418.200 ;
        RECT 788.400 416.400 792.600 417.600 ;
        RECT 766.950 414.000 777.600 414.600 ;
        RECT 767.400 413.400 777.600 414.000 ;
        RECT 670.950 410.400 681.600 411.600 ;
        RECT 670.950 409.800 673.050 410.400 ;
        RECT 694.950 409.800 697.050 411.900 ;
        RECT 718.950 411.450 721.050 411.900 ;
        RECT 733.950 411.450 736.050 411.900 ;
        RECT 718.950 410.250 736.050 411.450 ;
        RECT 718.950 409.800 721.050 410.250 ;
        RECT 733.950 409.800 736.050 410.250 ;
        RECT 760.950 409.950 763.050 412.050 ;
        RECT 776.400 411.900 777.600 413.400 ;
        RECT 791.400 411.900 792.600 416.400 ;
        RECT 797.400 416.400 823.050 417.600 ;
        RECT 797.400 412.050 798.600 416.400 ;
        RECT 820.950 416.100 823.050 416.400 ;
        RECT 832.950 417.600 835.050 418.050 ;
        RECT 865.950 417.600 868.050 418.200 ;
        RECT 832.950 416.400 868.050 417.600 ;
        RECT 868.950 417.600 871.050 421.050 ;
        RECT 889.950 420.600 892.050 421.050 ;
        RECT 884.400 419.400 892.050 420.600 ;
        RECT 868.950 417.000 879.600 417.600 ;
        RECT 869.400 416.400 879.600 417.000 ;
        RECT 832.950 415.950 835.050 416.400 ;
        RECT 865.950 416.100 868.050 416.400 ;
        RECT 775.950 409.800 778.050 411.900 ;
        RECT 790.950 409.800 793.050 411.900 ;
        RECT 796.950 409.950 799.050 412.050 ;
        RECT 88.950 408.600 91.050 409.050 ;
        RECT 94.950 408.600 97.050 409.050 ;
        RECT 88.950 407.400 97.050 408.600 ;
        RECT 88.950 406.950 91.050 407.400 ;
        RECT 94.950 406.950 97.050 407.400 ;
        RECT 112.950 408.600 115.050 409.050 ;
        RECT 118.950 408.600 121.050 409.050 ;
        RECT 112.950 407.400 121.050 408.600 ;
        RECT 112.950 406.950 115.050 407.400 ;
        RECT 118.950 406.950 121.050 407.400 ;
        RECT 127.950 408.600 130.050 409.050 ;
        RECT 133.950 408.600 136.050 409.050 ;
        RECT 127.950 407.400 136.050 408.600 ;
        RECT 127.950 406.950 130.050 407.400 ;
        RECT 133.950 406.950 136.050 407.400 ;
        RECT 328.950 408.600 331.050 409.050 ;
        RECT 349.950 408.600 352.050 409.050 ;
        RECT 367.950 408.600 370.050 409.050 ;
        RECT 328.950 407.400 370.050 408.600 ;
        RECT 328.950 406.950 331.050 407.400 ;
        RECT 349.950 406.950 352.050 407.400 ;
        RECT 367.950 406.950 370.050 407.400 ;
        RECT 424.950 408.600 427.050 409.050 ;
        RECT 430.950 408.600 433.050 409.050 ;
        RECT 424.950 407.400 433.050 408.600 ;
        RECT 424.950 406.950 427.050 407.400 ;
        RECT 430.950 406.950 433.050 407.400 ;
        RECT 499.950 408.600 502.050 409.050 ;
        RECT 509.400 408.600 510.600 409.800 ;
        RECT 499.950 407.400 510.600 408.600 ;
        RECT 557.400 408.600 558.600 409.800 ;
        RECT 878.400 409.050 879.600 416.400 ;
        RECT 880.950 415.950 883.050 418.050 ;
        RECT 881.400 411.600 882.600 415.950 ;
        RECT 884.400 414.600 885.600 419.400 ;
        RECT 889.950 418.950 892.050 419.400 ;
        RECT 886.950 417.600 889.050 418.200 ;
        RECT 895.950 417.600 898.050 418.050 ;
        RECT 886.950 416.400 898.050 417.600 ;
        RECT 886.950 416.100 889.050 416.400 ;
        RECT 895.950 415.950 898.050 416.400 ;
        RECT 899.400 414.600 900.600 422.400 ;
        RECT 884.400 413.400 891.600 414.600 ;
        RECT 890.400 411.900 891.600 413.400 ;
        RECT 896.400 413.400 900.600 414.600 ;
        RECT 883.950 411.600 886.050 411.900 ;
        RECT 881.400 410.400 886.050 411.600 ;
        RECT 883.950 409.800 886.050 410.400 ;
        RECT 889.950 409.800 892.050 411.900 ;
        RECT 592.950 408.600 595.050 409.050 ;
        RECT 557.400 407.400 595.050 408.600 ;
        RECT 499.950 406.950 502.050 407.400 ;
        RECT 592.950 406.950 595.050 407.400 ;
        RECT 682.950 408.600 685.050 409.050 ;
        RECT 715.950 408.600 718.050 409.050 ;
        RECT 682.950 407.400 718.050 408.600 ;
        RECT 682.950 406.950 685.050 407.400 ;
        RECT 715.950 406.950 718.050 407.400 ;
        RECT 739.950 408.600 742.050 409.050 ;
        RECT 754.950 408.600 757.050 409.050 ;
        RECT 739.950 407.400 757.050 408.600 ;
        RECT 739.950 406.950 742.050 407.400 ;
        RECT 754.950 406.950 757.050 407.400 ;
        RECT 811.950 408.600 814.050 409.050 ;
        RECT 823.950 408.600 826.050 409.050 ;
        RECT 862.950 408.600 865.050 409.050 ;
        RECT 811.950 407.400 865.050 408.600 ;
        RECT 878.400 407.400 883.050 409.050 ;
        RECT 811.950 406.950 814.050 407.400 ;
        RECT 823.950 406.950 826.050 407.400 ;
        RECT 862.950 406.950 865.050 407.400 ;
        RECT 879.000 406.950 883.050 407.400 ;
        RECT 4.950 405.600 7.050 406.050 ;
        RECT 22.950 405.600 25.050 406.050 ;
        RECT 4.950 404.400 25.050 405.600 ;
        RECT 4.950 403.950 7.050 404.400 ;
        RECT 22.950 403.950 25.050 404.400 ;
        RECT 37.950 405.600 40.050 406.050 ;
        RECT 55.950 405.600 58.050 406.050 ;
        RECT 37.950 404.400 58.050 405.600 ;
        RECT 37.950 403.950 40.050 404.400 ;
        RECT 55.950 403.950 58.050 404.400 ;
        RECT 64.950 405.600 67.050 406.050 ;
        RECT 91.950 405.600 94.050 406.050 ;
        RECT 64.950 404.400 94.050 405.600 ;
        RECT 64.950 403.950 67.050 404.400 ;
        RECT 91.950 403.950 94.050 404.400 ;
        RECT 193.950 405.600 196.050 406.050 ;
        RECT 214.950 405.600 217.050 406.050 ;
        RECT 241.950 405.600 244.050 406.050 ;
        RECT 247.950 405.600 250.050 406.050 ;
        RECT 193.950 404.400 250.050 405.600 ;
        RECT 193.950 403.950 196.050 404.400 ;
        RECT 214.950 403.950 217.050 404.400 ;
        RECT 241.950 403.950 244.050 404.400 ;
        RECT 247.950 403.950 250.050 404.400 ;
        RECT 382.950 405.600 385.050 406.050 ;
        RECT 415.950 405.600 418.050 406.050 ;
        RECT 382.950 404.400 418.050 405.600 ;
        RECT 382.950 403.950 385.050 404.400 ;
        RECT 415.950 403.950 418.050 404.400 ;
        RECT 535.950 405.600 538.050 406.050 ;
        RECT 547.950 405.600 550.050 406.050 ;
        RECT 535.950 404.400 550.050 405.600 ;
        RECT 535.950 403.950 538.050 404.400 ;
        RECT 547.950 403.950 550.050 404.400 ;
        RECT 607.950 405.600 610.050 406.050 ;
        RECT 640.950 405.600 643.050 406.050 ;
        RECT 607.950 404.400 643.050 405.600 ;
        RECT 607.950 403.950 610.050 404.400 ;
        RECT 640.950 403.950 643.050 404.400 ;
        RECT 667.950 405.600 670.050 406.050 ;
        RECT 676.950 405.600 679.050 406.050 ;
        RECT 667.950 404.400 679.050 405.600 ;
        RECT 667.950 403.950 670.050 404.400 ;
        RECT 676.950 403.950 679.050 404.400 ;
        RECT 688.950 405.600 691.050 406.050 ;
        RECT 724.950 405.600 727.050 406.050 ;
        RECT 688.950 404.400 727.050 405.600 ;
        RECT 688.950 403.950 691.050 404.400 ;
        RECT 724.950 403.950 727.050 404.400 ;
        RECT 874.950 405.600 877.050 406.050 ;
        RECT 892.950 405.600 895.050 406.050 ;
        RECT 874.950 404.400 895.050 405.600 ;
        RECT 874.950 403.950 877.050 404.400 ;
        RECT 892.950 403.950 895.050 404.400 ;
        RECT 58.950 402.600 61.050 403.050 ;
        RECT 124.950 402.600 127.050 403.050 ;
        RECT 58.950 401.400 127.050 402.600 ;
        RECT 58.950 400.950 61.050 401.400 ;
        RECT 124.950 400.950 127.050 401.400 ;
        RECT 298.950 402.600 301.050 403.050 ;
        RECT 361.950 402.600 364.050 403.050 ;
        RECT 298.950 401.400 364.050 402.600 ;
        RECT 298.950 400.950 301.050 401.400 ;
        RECT 361.950 400.950 364.050 401.400 ;
        RECT 367.950 402.600 370.050 403.050 ;
        RECT 373.950 402.600 376.050 403.050 ;
        RECT 463.950 402.600 466.050 403.050 ;
        RECT 367.950 401.400 466.050 402.600 ;
        RECT 367.950 400.950 370.050 401.400 ;
        RECT 373.950 400.950 376.050 401.400 ;
        RECT 463.950 400.950 466.050 401.400 ;
        RECT 616.950 402.600 619.050 403.050 ;
        RECT 634.950 402.600 637.050 403.050 ;
        RECT 616.950 401.400 637.050 402.600 ;
        RECT 616.950 400.950 619.050 401.400 ;
        RECT 634.950 400.950 637.050 401.400 ;
        RECT 736.950 402.600 739.050 403.050 ;
        RECT 769.950 402.600 772.050 403.050 ;
        RECT 736.950 401.400 772.050 402.600 ;
        RECT 736.950 400.950 739.050 401.400 ;
        RECT 769.950 400.950 772.050 401.400 ;
        RECT 811.950 402.600 814.050 403.050 ;
        RECT 853.950 402.600 856.050 403.050 ;
        RECT 811.950 401.400 856.050 402.600 ;
        RECT 811.950 400.950 814.050 401.400 ;
        RECT 853.950 400.950 856.050 401.400 ;
        RECT 886.950 402.600 889.050 403.050 ;
        RECT 896.400 402.600 897.600 413.400 ;
        RECT 886.950 401.400 897.600 402.600 ;
        RECT 886.950 400.950 889.050 401.400 ;
        RECT 124.950 399.600 127.050 399.900 ;
        RECT 169.950 399.600 172.050 400.050 ;
        RECT 124.950 398.400 172.050 399.600 ;
        RECT 124.950 397.800 127.050 398.400 ;
        RECT 169.950 397.950 172.050 398.400 ;
        RECT 220.950 399.600 223.050 400.050 ;
        RECT 232.950 399.600 235.050 400.050 ;
        RECT 220.950 398.400 235.050 399.600 ;
        RECT 220.950 397.950 223.050 398.400 ;
        RECT 232.950 397.950 235.050 398.400 ;
        RECT 358.950 399.600 361.050 400.050 ;
        RECT 364.950 399.600 367.050 400.050 ;
        RECT 358.950 398.400 367.050 399.600 ;
        RECT 358.950 397.950 361.050 398.400 ;
        RECT 364.950 397.950 367.050 398.400 ;
        RECT 409.950 399.600 412.050 400.050 ;
        RECT 439.950 399.600 442.050 400.050 ;
        RECT 409.950 398.400 442.050 399.600 ;
        RECT 409.950 397.950 412.050 398.400 ;
        RECT 439.950 397.950 442.050 398.400 ;
        RECT 508.950 399.600 511.050 400.050 ;
        RECT 577.950 399.600 580.050 400.050 ;
        RECT 643.950 399.600 646.050 400.050 ;
        RECT 508.950 398.400 646.050 399.600 ;
        RECT 508.950 397.950 511.050 398.400 ;
        RECT 577.950 397.950 580.050 398.400 ;
        RECT 643.950 397.950 646.050 398.400 ;
        RECT 37.950 396.600 40.050 397.050 ;
        RECT 190.950 396.600 193.050 397.050 ;
        RECT 445.950 396.600 448.050 397.050 ;
        RECT 37.950 395.400 448.050 396.600 ;
        RECT 37.950 394.950 40.050 395.400 ;
        RECT 190.950 394.950 193.050 395.400 ;
        RECT 445.950 394.950 448.050 395.400 ;
        RECT 604.950 396.600 607.050 397.050 ;
        RECT 616.950 396.600 619.050 397.050 ;
        RECT 604.950 395.400 619.050 396.600 ;
        RECT 604.950 394.950 607.050 395.400 ;
        RECT 616.950 394.950 619.050 395.400 ;
        RECT 700.950 396.600 703.050 397.050 ;
        RECT 712.950 396.600 715.050 397.050 ;
        RECT 700.950 395.400 715.050 396.600 ;
        RECT 700.950 394.950 703.050 395.400 ;
        RECT 712.950 394.950 715.050 395.400 ;
        RECT 733.950 396.600 736.050 397.050 ;
        RECT 799.950 396.600 802.050 397.050 ;
        RECT 733.950 395.400 802.050 396.600 ;
        RECT 733.950 394.950 736.050 395.400 ;
        RECT 799.950 394.950 802.050 395.400 ;
        RECT 823.950 396.600 826.050 397.050 ;
        RECT 889.950 396.600 892.050 397.050 ;
        RECT 823.950 395.400 892.050 396.600 ;
        RECT 823.950 394.950 826.050 395.400 ;
        RECT 889.950 394.950 892.050 395.400 ;
        RECT 187.950 393.600 190.050 394.050 ;
        RECT 205.950 393.600 208.050 394.050 ;
        RECT 187.950 392.400 208.050 393.600 ;
        RECT 187.950 391.950 190.050 392.400 ;
        RECT 205.950 391.950 208.050 392.400 ;
        RECT 277.950 393.600 280.050 394.050 ;
        RECT 292.950 393.600 295.050 394.050 ;
        RECT 277.950 392.400 295.050 393.600 ;
        RECT 277.950 391.950 280.050 392.400 ;
        RECT 292.950 391.950 295.050 392.400 ;
        RECT 367.950 393.600 370.050 394.050 ;
        RECT 388.950 393.600 391.050 394.050 ;
        RECT 367.950 392.400 391.050 393.600 ;
        RECT 367.950 391.950 370.050 392.400 ;
        RECT 388.950 391.950 391.050 392.400 ;
        RECT 679.950 393.600 682.050 394.050 ;
        RECT 685.950 393.600 688.050 394.050 ;
        RECT 706.950 393.600 709.050 394.050 ;
        RECT 748.800 393.600 750.900 394.050 ;
        RECT 679.950 392.400 750.900 393.600 ;
        RECT 679.950 391.950 682.050 392.400 ;
        RECT 685.950 391.950 688.050 392.400 ;
        RECT 706.950 391.950 709.050 392.400 ;
        RECT 748.800 391.950 750.900 392.400 ;
        RECT 751.950 393.600 754.050 394.050 ;
        RECT 763.950 393.600 766.050 394.050 ;
        RECT 868.950 393.600 871.050 394.050 ;
        RECT 751.950 392.400 766.050 393.600 ;
        RECT 751.950 391.950 754.050 392.400 ;
        RECT 763.950 391.950 766.050 392.400 ;
        RECT 827.400 392.400 871.050 393.600 ;
        RECT 88.950 390.600 91.050 391.050 ;
        RECT 103.950 390.600 106.050 391.050 ;
        RECT 88.950 389.400 106.050 390.600 ;
        RECT 88.950 388.950 91.050 389.400 ;
        RECT 103.950 388.950 106.050 389.400 ;
        RECT 511.950 390.600 514.050 391.050 ;
        RECT 550.950 390.600 553.050 391.050 ;
        RECT 511.950 389.400 553.050 390.600 ;
        RECT 511.950 388.950 514.050 389.400 ;
        RECT 550.950 388.950 553.050 389.400 ;
        RECT 625.950 390.600 628.050 391.050 ;
        RECT 658.950 390.600 661.050 391.050 ;
        RECT 625.950 389.400 661.050 390.600 ;
        RECT 625.950 388.950 628.050 389.400 ;
        RECT 658.950 388.950 661.050 389.400 ;
        RECT 808.950 390.600 811.050 391.050 ;
        RECT 827.400 390.600 828.600 392.400 ;
        RECT 868.950 391.950 871.050 392.400 ;
        RECT 808.950 389.400 828.600 390.600 ;
        RECT 808.950 388.950 811.050 389.400 ;
        RECT 70.950 387.600 73.050 388.050 ;
        RECT 85.950 387.600 88.050 388.050 ;
        RECT 70.950 386.400 88.050 387.600 ;
        RECT 70.950 385.950 73.050 386.400 ;
        RECT 85.950 385.950 88.050 386.400 ;
        RECT 586.950 387.600 589.050 388.050 ;
        RECT 622.950 387.600 625.050 388.050 ;
        RECT 586.950 386.400 625.050 387.600 ;
        RECT 586.950 385.950 589.050 386.400 ;
        RECT 622.950 385.950 625.050 386.400 ;
        RECT 715.950 387.600 718.050 388.050 ;
        RECT 766.950 387.600 769.050 388.050 ;
        RECT 715.950 386.400 769.050 387.600 ;
        RECT 715.950 385.950 718.050 386.400 ;
        RECT 766.950 385.950 769.050 386.400 ;
        RECT 781.950 387.600 784.050 388.050 ;
        RECT 829.950 387.600 832.050 388.050 ;
        RECT 781.950 386.400 832.050 387.600 ;
        RECT 781.950 385.950 784.050 386.400 ;
        RECT 829.950 385.950 832.050 386.400 ;
        RECT 244.950 384.600 247.050 385.050 ;
        RECT 259.950 384.600 262.050 385.050 ;
        RECT 244.950 383.400 262.050 384.600 ;
        RECT 244.950 382.950 247.050 383.400 ;
        RECT 259.950 382.950 262.050 383.400 ;
        RECT 283.950 384.600 286.050 385.050 ;
        RECT 316.950 384.600 319.050 385.050 ;
        RECT 283.950 383.400 319.050 384.600 ;
        RECT 283.950 382.950 286.050 383.400 ;
        RECT 316.950 382.950 319.050 383.400 ;
        RECT 340.950 384.600 343.050 385.050 ;
        RECT 400.950 384.600 403.050 385.050 ;
        RECT 340.950 383.400 403.050 384.600 ;
        RECT 340.950 382.950 343.050 383.400 ;
        RECT 400.950 382.950 403.050 383.400 ;
        RECT 538.950 384.600 541.050 385.050 ;
        RECT 574.950 384.600 577.050 385.050 ;
        RECT 538.950 383.400 577.050 384.600 ;
        RECT 538.950 382.950 541.050 383.400 ;
        RECT 574.950 382.950 577.050 383.400 ;
        RECT 631.950 384.600 634.050 385.050 ;
        RECT 706.950 384.600 709.050 385.050 ;
        RECT 787.950 384.600 790.050 385.050 ;
        RECT 631.950 383.400 790.050 384.600 ;
        RECT 631.950 382.950 634.050 383.400 ;
        RECT 706.950 382.950 709.050 383.400 ;
        RECT 787.950 382.950 790.050 383.400 ;
        RECT 97.950 381.600 100.050 382.050 ;
        RECT 172.950 381.600 175.050 382.050 ;
        RECT 97.950 380.400 175.050 381.600 ;
        RECT 97.950 379.950 100.050 380.400 ;
        RECT 172.950 379.950 175.050 380.400 ;
        RECT 238.950 381.600 241.050 382.050 ;
        RECT 262.950 381.600 265.050 382.050 ;
        RECT 424.950 381.600 427.050 382.050 ;
        RECT 238.950 380.400 427.050 381.600 ;
        RECT 238.950 379.950 241.050 380.400 ;
        RECT 262.950 379.950 265.050 380.400 ;
        RECT 67.950 378.600 70.050 379.050 ;
        RECT 79.950 378.600 82.050 379.050 ;
        RECT 142.950 378.600 145.050 379.050 ;
        RECT 67.950 377.400 82.050 378.600 ;
        RECT 67.950 376.950 70.050 377.400 ;
        RECT 79.950 376.950 82.050 377.400 ;
        RECT 128.400 377.400 145.050 378.600 ;
        RECT 128.400 376.050 129.600 377.400 ;
        RECT 142.950 376.950 145.050 377.400 ;
        RECT 382.950 376.950 385.050 380.400 ;
        RECT 424.950 379.950 427.050 380.400 ;
        RECT 487.950 381.600 490.050 382.050 ;
        RECT 493.950 381.600 496.050 382.050 ;
        RECT 511.950 381.600 514.050 382.050 ;
        RECT 487.950 380.400 514.050 381.600 ;
        RECT 487.950 379.950 490.050 380.400 ;
        RECT 493.950 379.950 496.050 380.400 ;
        RECT 511.950 379.950 514.050 380.400 ;
        RECT 589.950 381.600 592.050 382.050 ;
        RECT 604.950 381.600 607.050 382.050 ;
        RECT 589.950 380.400 607.050 381.600 ;
        RECT 589.950 379.950 592.050 380.400 ;
        RECT 604.950 379.950 607.050 380.400 ;
        RECT 649.950 381.600 652.050 382.050 ;
        RECT 736.950 381.600 739.050 382.050 ;
        RECT 649.950 380.400 739.050 381.600 ;
        RECT 649.950 379.950 652.050 380.400 ;
        RECT 736.950 379.950 739.050 380.400 ;
        RECT 832.950 381.600 835.050 382.050 ;
        RECT 862.950 381.600 865.050 382.050 ;
        RECT 832.950 380.400 865.050 381.600 ;
        RECT 832.950 379.950 835.050 380.400 ;
        RECT 862.950 379.950 865.050 380.400 ;
        RECT 616.950 378.600 619.050 379.050 ;
        RECT 622.950 378.600 625.050 379.050 ;
        RECT 649.950 378.600 652.050 378.900 ;
        RECT 616.950 377.400 652.050 378.600 ;
        RECT 616.950 376.950 619.050 377.400 ;
        RECT 622.950 376.950 625.050 377.400 ;
        RECT 649.950 376.800 652.050 377.400 ;
        RECT 664.950 378.600 667.050 379.050 ;
        RECT 718.950 378.600 721.050 379.050 ;
        RECT 664.950 377.400 721.050 378.600 ;
        RECT 664.950 376.950 667.050 377.400 ;
        RECT 718.950 376.950 721.050 377.400 ;
        RECT 832.950 378.600 835.050 378.900 ;
        RECT 841.950 378.600 844.050 379.050 ;
        RECT 832.950 377.400 844.050 378.600 ;
        RECT 832.950 376.800 835.050 377.400 ;
        RECT 841.950 376.950 844.050 377.400 ;
        RECT 4.950 375.600 7.050 376.050 ;
        RECT 22.950 375.600 25.050 376.050 ;
        RECT 112.950 375.600 115.050 376.050 ;
        RECT 127.950 375.600 130.050 376.050 ;
        RECT 4.950 374.400 130.050 375.600 ;
        RECT 4.950 373.950 7.050 374.400 ;
        RECT 22.950 373.950 25.050 374.400 ;
        RECT 112.950 373.950 115.050 374.400 ;
        RECT 127.950 373.950 130.050 374.400 ;
        RECT 265.950 375.600 268.050 376.050 ;
        RECT 298.950 375.600 301.050 376.050 ;
        RECT 265.950 374.400 301.050 375.600 ;
        RECT 265.950 373.950 268.050 374.400 ;
        RECT 298.950 373.950 301.050 374.400 ;
        RECT 334.950 375.600 337.050 376.050 ;
        RECT 346.950 375.600 349.050 376.050 ;
        RECT 334.950 374.400 349.050 375.600 ;
        RECT 334.950 373.950 337.050 374.400 ;
        RECT 346.950 373.950 349.050 374.400 ;
        RECT 517.950 375.600 520.050 376.050 ;
        RECT 529.950 375.600 532.050 376.050 ;
        RECT 517.950 374.400 532.050 375.600 ;
        RECT 517.950 373.950 520.050 374.400 ;
        RECT 529.950 373.950 532.050 374.400 ;
        RECT 541.950 375.600 544.050 376.050 ;
        RECT 553.950 375.600 556.050 376.050 ;
        RECT 541.950 374.400 556.050 375.600 ;
        RECT 541.950 373.950 544.050 374.400 ;
        RECT 553.950 373.950 556.050 374.400 ;
        RECT 601.950 375.600 604.050 376.050 ;
        RECT 631.950 375.600 634.050 376.050 ;
        RECT 601.950 374.400 634.050 375.600 ;
        RECT 601.950 373.950 604.050 374.400 ;
        RECT 631.950 373.950 634.050 374.400 ;
        RECT 742.950 375.600 745.050 376.050 ;
        RECT 757.950 375.600 760.050 376.050 ;
        RECT 814.950 375.600 817.050 376.050 ;
        RECT 742.950 374.400 760.050 375.600 ;
        RECT 742.950 373.950 745.050 374.400 ;
        RECT 757.950 373.950 760.050 374.400 ;
        RECT 809.400 374.400 817.050 375.600 ;
        RECT 13.950 373.050 16.050 373.500 ;
        RECT 19.950 373.050 22.050 373.500 ;
        RECT 13.950 371.850 22.050 373.050 ;
        RECT 13.950 371.400 16.050 371.850 ;
        RECT 19.950 371.400 22.050 371.850 ;
        RECT 49.950 371.100 52.050 373.200 ;
        RECT 73.950 372.600 76.050 373.200 ;
        RECT 94.950 372.600 97.050 373.050 ;
        RECT 121.950 372.600 124.050 373.050 ;
        RECT 130.950 372.600 133.050 373.200 ;
        RECT 73.950 371.400 133.050 372.600 ;
        RECT 73.950 371.100 76.050 371.400 ;
        RECT 50.400 364.050 51.600 371.100 ;
        RECT 74.400 369.600 75.600 371.100 ;
        RECT 94.950 370.950 97.050 371.400 ;
        RECT 121.950 370.950 124.050 371.400 ;
        RECT 130.950 371.100 133.050 371.400 ;
        RECT 145.950 372.600 148.050 373.050 ;
        RECT 154.950 372.600 157.050 373.200 ;
        RECT 145.950 371.400 157.050 372.600 ;
        RECT 145.950 370.950 148.050 371.400 ;
        RECT 154.950 371.100 157.050 371.400 ;
        RECT 172.950 371.100 175.050 373.200 ;
        RECT 178.950 371.100 181.050 373.200 ;
        RECT 184.950 372.600 187.050 373.050 ;
        RECT 199.950 372.600 202.050 373.200 ;
        RECT 184.950 371.400 202.050 372.600 ;
        RECT 226.950 372.600 229.050 373.500 ;
        RECT 247.950 372.750 250.050 373.200 ;
        RECT 253.950 372.750 256.050 373.200 ;
        RECT 226.950 371.400 240.600 372.600 ;
        RECT 59.400 368.400 75.600 369.600 ;
        RECT 59.400 366.900 60.600 368.400 ;
        RECT 58.950 364.800 61.050 366.900 ;
        RECT 67.950 366.150 70.050 367.050 ;
        RECT 82.950 366.150 85.050 367.050 ;
        RECT 85.950 366.150 88.050 366.600 ;
        RECT 67.950 364.950 88.050 366.150 ;
        RECT 85.950 364.500 88.050 364.950 ;
        RECT 31.950 360.600 34.050 364.050 ;
        RECT 49.950 361.950 52.050 364.050 ;
        RECT 157.950 363.600 160.050 364.050 ;
        RECT 173.400 363.600 174.600 371.100 ;
        RECT 179.400 367.050 180.600 371.100 ;
        RECT 184.950 370.950 187.050 371.400 ;
        RECT 199.950 371.100 202.050 371.400 ;
        RECT 239.400 367.050 240.600 371.400 ;
        RECT 247.950 371.550 256.050 372.750 ;
        RECT 247.950 371.100 250.050 371.550 ;
        RECT 253.950 371.100 256.050 371.550 ;
        RECT 259.950 372.750 262.050 373.200 ;
        RECT 271.950 372.750 274.050 373.200 ;
        RECT 259.950 371.550 274.050 372.750 ;
        RECT 259.950 371.100 262.050 371.550 ;
        RECT 271.950 371.100 274.050 371.550 ;
        RECT 322.950 372.600 325.050 373.200 ;
        RECT 373.950 372.600 376.050 373.500 ;
        RECT 322.950 371.400 327.600 372.600 ;
        RECT 322.950 371.100 325.050 371.400 ;
        RECT 179.400 365.400 184.050 367.050 ;
        RECT 180.000 364.950 184.050 365.400 ;
        RECT 190.950 366.600 193.050 367.050 ;
        RECT 205.950 366.600 208.050 367.050 ;
        RECT 190.950 365.400 208.050 366.600 ;
        RECT 190.950 364.950 193.050 365.400 ;
        RECT 205.950 364.950 208.050 365.400 ;
        RECT 238.950 364.950 241.050 367.050 ;
        RECT 244.950 366.450 247.050 366.900 ;
        RECT 250.950 366.450 253.050 366.900 ;
        RECT 244.950 365.250 253.050 366.450 ;
        RECT 244.950 364.800 247.050 365.250 ;
        RECT 250.950 364.800 253.050 365.250 ;
        RECT 271.950 366.600 274.050 367.050 ;
        RECT 280.950 366.600 283.050 366.900 ;
        RECT 271.950 365.400 283.050 366.600 ;
        RECT 326.400 366.600 327.600 371.400 ;
        RECT 344.400 371.400 376.050 372.600 ;
        RECT 344.400 366.900 345.600 371.400 ;
        RECT 385.950 370.950 388.050 373.050 ;
        RECT 409.950 371.400 412.050 373.500 ;
        RECT 418.950 372.600 421.050 373.500 ;
        RECT 427.950 372.600 430.050 373.500 ;
        RECT 418.950 371.400 430.050 372.600 ;
        RECT 436.950 373.050 439.050 373.500 ;
        RECT 460.950 373.050 463.050 373.500 ;
        RECT 436.950 371.850 463.050 373.050 ;
        RECT 436.950 371.400 439.050 371.850 ;
        RECT 460.950 371.400 463.050 371.850 ;
        RECT 472.950 372.600 475.050 373.200 ;
        RECT 499.950 372.600 502.050 373.200 ;
        RECT 472.950 371.400 502.050 372.600 ;
        RECT 337.950 366.600 340.050 366.900 ;
        RECT 326.400 365.400 340.050 366.600 ;
        RECT 271.950 364.950 274.050 365.400 ;
        RECT 280.950 364.800 283.050 365.400 ;
        RECT 337.950 364.800 340.050 365.400 ;
        RECT 343.950 364.800 346.050 366.900 ;
        RECT 370.950 366.600 373.050 367.050 ;
        RECT 386.400 366.600 387.600 370.950 ;
        RECT 370.950 365.400 387.600 366.600 ;
        RECT 370.950 364.950 373.050 365.400 ;
        RECT 410.400 364.050 411.600 371.400 ;
        RECT 419.400 367.050 420.600 371.400 ;
        RECT 472.950 371.100 475.050 371.400 ;
        RECT 499.950 371.100 502.050 371.400 ;
        RECT 505.950 372.600 508.050 373.050 ;
        RECT 514.950 372.600 517.050 373.050 ;
        RECT 523.950 372.600 526.050 373.200 ;
        RECT 505.950 371.400 517.050 372.600 ;
        RECT 505.950 370.950 508.050 371.400 ;
        RECT 514.950 370.950 517.050 371.400 ;
        RECT 518.400 371.400 526.050 372.600 ;
        RECT 419.400 365.400 424.050 367.050 ;
        RECT 475.950 366.600 478.050 366.900 ;
        RECT 496.950 366.600 499.050 366.900 ;
        RECT 420.000 364.950 424.050 365.400 ;
        RECT 454.950 366.150 457.050 366.600 ;
        RECT 466.950 366.150 469.050 366.600 ;
        RECT 454.950 364.950 469.050 366.150 ;
        RECT 454.950 364.500 457.050 364.950 ;
        RECT 466.950 364.500 469.050 364.950 ;
        RECT 475.950 365.400 499.050 366.600 ;
        RECT 475.950 364.800 478.050 365.400 ;
        RECT 496.950 364.800 499.050 365.400 ;
        RECT 505.950 366.600 508.050 367.050 ;
        RECT 518.400 366.600 519.600 371.400 ;
        RECT 523.950 371.100 526.050 371.400 ;
        RECT 565.950 372.600 568.050 372.900 ;
        RECT 574.950 372.600 577.050 373.200 ;
        RECT 598.950 372.600 601.050 373.200 ;
        RECT 565.950 371.400 601.050 372.600 ;
        RECT 565.950 370.800 568.050 371.400 ;
        RECT 574.950 371.100 577.050 371.400 ;
        RECT 598.950 371.100 601.050 371.400 ;
        RECT 619.950 372.600 622.050 373.050 ;
        RECT 625.950 372.600 628.050 373.200 ;
        RECT 619.950 371.400 628.050 372.600 ;
        RECT 619.950 370.950 622.050 371.400 ;
        RECT 625.950 371.100 628.050 371.400 ;
        RECT 709.950 372.750 712.050 373.200 ;
        RECT 721.950 372.750 724.050 373.200 ;
        RECT 709.950 371.550 724.050 372.750 ;
        RECT 709.950 371.100 712.050 371.550 ;
        RECT 721.950 371.100 724.050 371.550 ;
        RECT 727.950 372.750 730.050 373.200 ;
        RECT 739.950 372.750 742.050 373.200 ;
        RECT 727.950 371.550 742.050 372.750 ;
        RECT 727.950 371.100 730.050 371.550 ;
        RECT 739.950 371.100 742.050 371.550 ;
        RECT 745.950 372.600 748.050 373.200 ;
        RECT 754.950 372.600 757.050 373.050 ;
        RECT 796.950 372.600 799.050 373.200 ;
        RECT 745.950 371.400 757.050 372.600 ;
        RECT 745.950 371.100 748.050 371.400 ;
        RECT 754.950 370.950 757.050 371.400 ;
        RECT 794.400 371.400 799.050 372.600 ;
        RECT 613.950 369.600 616.050 370.050 ;
        RECT 530.400 368.400 616.050 369.600 ;
        RECT 530.400 366.900 531.600 368.400 ;
        RECT 572.400 366.900 573.600 368.400 ;
        RECT 596.400 366.900 597.600 368.400 ;
        RECT 613.950 367.950 616.050 368.400 ;
        RECT 794.400 367.050 795.600 371.400 ;
        RECT 796.950 371.100 799.050 371.400 ;
        RECT 802.950 371.100 805.050 373.200 ;
        RECT 505.950 365.400 519.600 366.600 ;
        RECT 505.950 364.950 508.050 365.400 ;
        RECT 529.950 364.800 532.050 366.900 ;
        RECT 571.950 364.800 574.050 366.900 ;
        RECT 595.950 364.800 598.050 366.900 ;
        RECT 622.950 366.450 625.050 366.900 ;
        RECT 631.950 366.450 634.050 366.900 ;
        RECT 622.950 365.250 634.050 366.450 ;
        RECT 622.950 364.800 625.050 365.250 ;
        RECT 631.950 364.800 634.050 365.250 ;
        RECT 736.950 366.450 739.050 366.900 ;
        RECT 742.950 366.450 745.050 366.900 ;
        RECT 736.950 365.250 745.050 366.450 ;
        RECT 736.950 364.800 739.050 365.250 ;
        RECT 742.950 364.800 745.050 365.250 ;
        RECT 793.950 364.950 796.050 367.050 ;
        RECT 184.950 363.600 187.050 364.050 ;
        RECT 157.950 362.400 187.050 363.600 ;
        RECT 157.950 361.950 160.050 362.400 ;
        RECT 184.950 361.950 187.050 362.400 ;
        RECT 202.950 363.600 205.050 364.050 ;
        RECT 208.950 363.600 211.050 364.050 ;
        RECT 220.950 363.600 223.050 364.050 ;
        RECT 202.950 362.400 223.050 363.600 ;
        RECT 202.950 361.950 205.050 362.400 ;
        RECT 208.950 361.950 211.050 362.400 ;
        RECT 220.950 361.950 223.050 362.400 ;
        RECT 301.950 363.600 304.050 364.050 ;
        RECT 331.950 363.600 334.050 364.050 ;
        RECT 355.950 363.600 358.050 364.050 ;
        RECT 301.950 362.400 334.050 363.600 ;
        RECT 301.950 361.950 304.050 362.400 ;
        RECT 331.950 361.950 334.050 362.400 ;
        RECT 347.400 362.400 358.050 363.600 ;
        RECT 37.950 360.600 40.050 361.050 ;
        RECT 31.950 360.000 40.050 360.600 ;
        RECT 32.400 359.400 40.050 360.000 ;
        RECT 37.950 358.950 40.050 359.400 ;
        RECT 124.950 360.600 127.050 361.050 ;
        RECT 139.950 360.600 142.050 361.050 ;
        RECT 124.950 359.400 142.050 360.600 ;
        RECT 124.950 358.950 127.050 359.400 ;
        RECT 139.950 358.950 142.050 359.400 ;
        RECT 196.950 360.600 199.050 361.050 ;
        RECT 217.950 360.600 220.050 361.050 ;
        RECT 196.950 359.400 220.050 360.600 ;
        RECT 196.950 358.950 199.050 359.400 ;
        RECT 217.950 358.950 220.050 359.400 ;
        RECT 238.950 360.600 241.050 361.050 ;
        RECT 256.950 360.600 259.050 361.050 ;
        RECT 238.950 359.400 259.050 360.600 ;
        RECT 238.950 358.950 241.050 359.400 ;
        RECT 256.950 358.950 259.050 359.400 ;
        RECT 325.950 360.600 328.050 361.050 ;
        RECT 347.400 360.600 348.600 362.400 ;
        RECT 355.950 361.950 358.050 362.400 ;
        RECT 409.950 361.950 412.050 364.050 ;
        RECT 532.950 363.600 535.050 364.050 ;
        RECT 541.950 363.600 544.050 364.050 ;
        RECT 547.950 363.600 550.050 364.050 ;
        RECT 532.950 362.400 550.050 363.600 ;
        RECT 532.950 361.950 535.050 362.400 ;
        RECT 541.950 361.950 544.050 362.400 ;
        RECT 547.950 361.950 550.050 362.400 ;
        RECT 643.950 363.600 646.050 364.050 ;
        RECT 709.950 363.600 712.050 364.050 ;
        RECT 643.950 362.400 712.050 363.600 ;
        RECT 643.950 361.950 646.050 362.400 ;
        RECT 709.950 361.950 712.050 362.400 ;
        RECT 730.950 363.600 733.050 364.050 ;
        RECT 748.950 363.600 751.050 364.050 ;
        RECT 730.950 362.400 751.050 363.600 ;
        RECT 730.950 361.950 733.050 362.400 ;
        RECT 748.950 361.950 751.050 362.400 ;
        RECT 763.950 363.600 766.050 363.900 ;
        RECT 803.400 363.600 804.600 371.100 ;
        RECT 809.400 367.050 810.600 374.400 ;
        RECT 814.950 373.950 817.050 374.400 ;
        RECT 841.950 371.100 844.050 373.200 ;
        RECT 847.800 371.100 849.900 373.200 ;
        RECT 850.950 372.600 853.050 373.050 ;
        RECT 856.950 372.600 859.050 373.050 ;
        RECT 850.950 371.400 859.050 372.600 ;
        RECT 842.400 369.600 843.600 371.100 ;
        RECT 836.400 369.000 843.600 369.600 ;
        RECT 835.950 368.400 843.600 369.000 ;
        RECT 808.950 364.950 811.050 367.050 ;
        RECT 835.950 364.950 838.050 368.400 ;
        RECT 763.950 362.400 804.600 363.600 ;
        RECT 763.950 361.800 766.050 362.400 ;
        RECT 325.950 359.400 348.600 360.600 ;
        RECT 460.950 360.600 463.050 361.050 ;
        RECT 502.950 360.600 505.050 361.050 ;
        RECT 583.950 360.600 586.050 361.050 ;
        RECT 460.950 359.400 505.050 360.600 ;
        RECT 325.950 358.950 328.050 359.400 ;
        RECT 460.950 358.950 463.050 359.400 ;
        RECT 502.950 358.950 505.050 359.400 ;
        RECT 554.400 359.400 586.050 360.600 ;
        RECT 19.950 357.600 22.050 358.050 ;
        RECT 52.950 357.600 55.050 358.050 ;
        RECT 19.950 356.400 55.050 357.600 ;
        RECT 19.950 355.950 22.050 356.400 ;
        RECT 52.950 355.950 55.050 356.400 ;
        RECT 64.950 357.600 67.050 358.050 ;
        RECT 76.950 357.600 79.050 358.050 ;
        RECT 64.950 356.400 79.050 357.600 ;
        RECT 64.950 355.950 67.050 356.400 ;
        RECT 76.950 355.950 79.050 356.400 ;
        RECT 151.950 357.600 154.050 358.050 ;
        RECT 169.950 357.600 172.050 358.050 ;
        RECT 187.950 357.600 190.050 358.050 ;
        RECT 151.950 356.400 190.050 357.600 ;
        RECT 151.950 355.950 154.050 356.400 ;
        RECT 169.950 355.950 172.050 356.400 ;
        RECT 187.950 355.950 190.050 356.400 ;
        RECT 256.950 357.600 259.050 357.900 ;
        RECT 268.950 357.600 271.050 358.050 ;
        RECT 256.950 356.400 271.050 357.600 ;
        RECT 256.950 355.800 259.050 356.400 ;
        RECT 268.950 355.950 271.050 356.400 ;
        RECT 289.950 357.600 292.050 358.050 ;
        RECT 388.950 357.600 391.050 358.050 ;
        RECT 289.950 356.400 391.050 357.600 ;
        RECT 289.950 355.950 292.050 356.400 ;
        RECT 388.950 355.950 391.050 356.400 ;
        RECT 514.950 357.600 517.050 358.050 ;
        RECT 554.400 357.600 555.600 359.400 ;
        RECT 583.950 358.950 586.050 359.400 ;
        RECT 631.950 360.600 634.050 361.050 ;
        RECT 652.950 360.600 655.050 361.050 ;
        RECT 667.950 360.600 670.050 361.050 ;
        RECT 631.950 359.400 670.050 360.600 ;
        RECT 803.400 360.600 804.600 362.400 ;
        RECT 805.950 363.600 808.050 364.050 ;
        RECT 832.950 363.600 835.050 364.050 ;
        RECT 838.950 363.600 841.050 364.050 ;
        RECT 805.950 362.400 841.050 363.600 ;
        RECT 805.950 361.950 808.050 362.400 ;
        RECT 832.950 361.950 835.050 362.400 ;
        RECT 838.950 361.950 841.050 362.400 ;
        RECT 848.400 360.600 849.600 371.100 ;
        RECT 850.950 370.950 853.050 371.400 ;
        RECT 856.950 370.950 859.050 371.400 ;
        RECT 865.950 366.450 868.050 366.900 ;
        RECT 895.950 366.450 898.050 366.900 ;
        RECT 865.950 365.250 898.050 366.450 ;
        RECT 865.950 364.800 868.050 365.250 ;
        RECT 895.950 364.800 898.050 365.250 ;
        RECT 803.400 359.400 849.600 360.600 ;
        RECT 631.950 358.950 634.050 359.400 ;
        RECT 652.950 358.950 655.050 359.400 ;
        RECT 667.950 358.950 670.050 359.400 ;
        RECT 514.950 356.400 555.600 357.600 ;
        RECT 613.950 357.600 616.050 358.050 ;
        RECT 634.950 357.600 637.050 358.050 ;
        RECT 613.950 356.400 637.050 357.600 ;
        RECT 514.950 355.950 517.050 356.400 ;
        RECT 613.950 355.950 616.050 356.400 ;
        RECT 634.950 355.950 637.050 356.400 ;
        RECT 697.950 357.600 700.050 358.050 ;
        RECT 763.950 357.600 766.050 358.050 ;
        RECT 697.950 356.400 766.050 357.600 ;
        RECT 697.950 355.950 700.050 356.400 ;
        RECT 763.950 355.950 766.050 356.400 ;
        RECT 778.950 357.600 781.050 358.050 ;
        RECT 835.950 357.600 838.050 358.050 ;
        RECT 778.950 356.400 838.050 357.600 ;
        RECT 778.950 355.950 781.050 356.400 ;
        RECT 835.950 355.950 838.050 356.400 ;
        RECT 229.950 354.600 232.050 355.050 ;
        RECT 241.950 354.600 244.050 355.050 ;
        RECT 229.950 353.400 244.050 354.600 ;
        RECT 229.950 352.950 232.050 353.400 ;
        RECT 241.950 352.950 244.050 353.400 ;
        RECT 361.950 354.600 364.050 355.050 ;
        RECT 370.950 354.600 373.050 355.050 ;
        RECT 361.950 353.400 373.050 354.600 ;
        RECT 361.950 352.950 364.050 353.400 ;
        RECT 370.950 352.950 373.050 353.400 ;
        RECT 478.950 354.600 481.050 355.050 ;
        RECT 538.950 354.600 541.050 355.050 ;
        RECT 478.950 353.400 541.050 354.600 ;
        RECT 478.950 352.950 481.050 353.400 ;
        RECT 538.950 352.950 541.050 353.400 ;
        RECT 556.950 354.600 559.050 355.050 ;
        RECT 646.950 354.600 649.050 355.050 ;
        RECT 556.950 353.400 649.050 354.600 ;
        RECT 556.950 352.950 559.050 353.400 ;
        RECT 646.950 352.950 649.050 353.400 ;
        RECT 652.950 354.600 655.050 355.050 ;
        RECT 688.950 354.600 691.050 355.050 ;
        RECT 754.950 354.600 757.050 355.050 ;
        RECT 652.950 353.400 757.050 354.600 ;
        RECT 652.950 352.950 655.050 353.400 ;
        RECT 688.950 352.950 691.050 353.400 ;
        RECT 754.950 352.950 757.050 353.400 ;
        RECT 775.950 354.600 778.050 355.050 ;
        RECT 865.950 354.600 868.050 355.050 ;
        RECT 775.950 353.400 868.050 354.600 ;
        RECT 775.950 352.950 778.050 353.400 ;
        RECT 865.950 352.950 868.050 353.400 ;
        RECT 181.950 351.600 184.050 352.050 ;
        RECT 196.950 351.600 199.050 352.050 ;
        RECT 181.950 350.400 199.050 351.600 ;
        RECT 181.950 349.950 184.050 350.400 ;
        RECT 196.950 349.950 199.050 350.400 ;
        RECT 262.950 351.600 265.050 352.050 ;
        RECT 307.950 351.600 310.050 352.050 ;
        RECT 262.950 350.400 310.050 351.600 ;
        RECT 262.950 349.950 265.050 350.400 ;
        RECT 307.950 349.950 310.050 350.400 ;
        RECT 463.950 351.600 466.050 352.050 ;
        RECT 475.950 351.600 478.050 352.050 ;
        RECT 463.950 350.400 478.050 351.600 ;
        RECT 463.950 349.950 466.050 350.400 ;
        RECT 475.950 349.950 478.050 350.400 ;
        RECT 571.950 351.600 574.050 352.050 ;
        RECT 643.950 351.600 646.050 352.050 ;
        RECT 571.950 350.400 646.050 351.600 ;
        RECT 571.950 349.950 574.050 350.400 ;
        RECT 643.950 349.950 646.050 350.400 ;
        RECT 121.950 348.600 124.050 349.050 ;
        RECT 133.950 348.600 136.050 349.050 ;
        RECT 121.950 347.400 136.050 348.600 ;
        RECT 121.950 346.950 124.050 347.400 ;
        RECT 133.950 346.950 136.050 347.400 ;
        RECT 241.950 348.600 244.050 349.050 ;
        RECT 277.950 348.600 280.050 349.050 ;
        RECT 337.950 348.600 340.050 349.050 ;
        RECT 241.950 347.400 340.050 348.600 ;
        RECT 241.950 346.950 244.050 347.400 ;
        RECT 277.950 346.950 280.050 347.400 ;
        RECT 337.950 346.950 340.050 347.400 ;
        RECT 379.950 348.600 382.050 349.050 ;
        RECT 421.950 348.600 424.050 349.050 ;
        RECT 379.950 347.400 424.050 348.600 ;
        RECT 379.950 346.950 382.050 347.400 ;
        RECT 421.950 346.950 424.050 347.400 ;
        RECT 496.950 348.600 499.050 349.050 ;
        RECT 508.950 348.600 511.050 349.050 ;
        RECT 496.950 347.400 511.050 348.600 ;
        RECT 496.950 346.950 499.050 347.400 ;
        RECT 508.950 346.950 511.050 347.400 ;
        RECT 517.950 348.600 520.050 349.050 ;
        RECT 541.950 348.600 544.050 349.050 ;
        RECT 517.950 347.400 544.050 348.600 ;
        RECT 517.950 346.950 520.050 347.400 ;
        RECT 541.950 346.950 544.050 347.400 ;
        RECT 586.950 348.600 589.050 349.050 ;
        RECT 601.950 348.600 604.050 349.050 ;
        RECT 586.950 347.400 604.050 348.600 ;
        RECT 586.950 346.950 589.050 347.400 ;
        RECT 601.950 346.950 604.050 347.400 ;
        RECT 718.950 348.600 721.050 349.050 ;
        RECT 724.950 348.600 727.050 349.050 ;
        RECT 718.950 347.400 727.050 348.600 ;
        RECT 718.950 346.950 721.050 347.400 ;
        RECT 724.950 346.950 727.050 347.400 ;
        RECT 748.950 348.600 751.050 349.050 ;
        RECT 760.950 348.600 763.050 349.050 ;
        RECT 787.950 348.600 790.050 349.050 ;
        RECT 820.950 348.600 823.050 349.050 ;
        RECT 748.950 347.400 823.050 348.600 ;
        RECT 748.950 346.950 751.050 347.400 ;
        RECT 760.950 346.950 763.050 347.400 ;
        RECT 787.950 346.950 790.050 347.400 ;
        RECT 820.950 346.950 823.050 347.400 ;
        RECT 835.950 348.600 838.050 349.050 ;
        RECT 871.950 348.600 874.050 349.050 ;
        RECT 835.950 347.400 874.050 348.600 ;
        RECT 835.950 346.950 838.050 347.400 ;
        RECT 871.950 346.950 874.050 347.400 ;
        RECT 187.950 345.600 190.050 346.050 ;
        RECT 199.950 345.600 202.050 346.050 ;
        RECT 217.950 345.600 220.050 346.050 ;
        RECT 187.950 344.400 220.050 345.600 ;
        RECT 187.950 343.950 190.050 344.400 ;
        RECT 199.950 343.950 202.050 344.400 ;
        RECT 217.950 343.950 220.050 344.400 ;
        RECT 490.950 345.600 493.050 346.050 ;
        RECT 514.950 345.600 517.050 346.050 ;
        RECT 706.950 345.600 709.050 346.050 ;
        RECT 490.950 344.400 517.050 345.600 ;
        RECT 490.950 343.950 493.050 344.400 ;
        RECT 514.950 343.950 517.050 344.400 ;
        RECT 698.400 344.400 709.050 345.600 ;
        RECT 40.950 342.600 43.050 343.050 ;
        RECT 76.950 342.600 79.050 343.050 ;
        RECT 40.950 341.400 79.050 342.600 ;
        RECT 40.950 340.950 43.050 341.400 ;
        RECT 76.950 340.950 79.050 341.400 ;
        RECT 103.950 339.600 106.050 340.200 ;
        RECT 115.950 339.600 118.050 340.050 ;
        RECT 103.950 338.400 118.050 339.600 ;
        RECT 121.950 339.600 124.050 343.050 ;
        RECT 145.950 342.600 148.050 343.050 ;
        RECT 160.950 342.600 163.050 343.050 ;
        RECT 145.950 341.400 163.050 342.600 ;
        RECT 145.950 340.950 148.050 341.400 ;
        RECT 160.950 340.950 163.050 341.400 ;
        RECT 175.950 342.600 178.050 343.050 ;
        RECT 181.950 342.600 184.050 343.050 ;
        RECT 175.950 341.400 184.050 342.600 ;
        RECT 175.950 340.950 178.050 341.400 ;
        RECT 181.950 340.950 184.050 341.400 ;
        RECT 364.950 342.600 367.050 343.050 ;
        RECT 451.950 342.600 454.050 343.050 ;
        RECT 466.950 342.600 469.050 343.050 ;
        RECT 364.950 341.400 469.050 342.600 ;
        RECT 364.950 340.950 367.050 341.400 ;
        RECT 451.950 340.950 454.050 341.400 ;
        RECT 466.950 340.950 469.050 341.400 ;
        RECT 610.950 342.600 613.050 343.050 ;
        RECT 622.950 342.600 625.050 343.050 ;
        RECT 610.950 341.400 625.050 342.600 ;
        RECT 610.950 340.950 613.050 341.400 ;
        RECT 622.950 340.950 625.050 341.400 ;
        RECT 676.950 342.600 679.050 343.050 ;
        RECT 698.400 342.600 699.600 344.400 ;
        RECT 706.950 343.950 709.050 344.400 ;
        RECT 715.950 345.600 718.050 346.050 ;
        RECT 727.950 345.600 730.050 346.050 ;
        RECT 715.950 344.400 730.050 345.600 ;
        RECT 715.950 343.950 718.050 344.400 ;
        RECT 727.950 343.950 730.050 344.400 ;
        RECT 805.950 345.600 808.050 346.050 ;
        RECT 820.950 345.600 823.050 345.900 ;
        RECT 805.950 344.400 823.050 345.600 ;
        RECT 805.950 343.950 808.050 344.400 ;
        RECT 820.950 343.800 823.050 344.400 ;
        RECT 844.950 345.600 847.050 346.050 ;
        RECT 859.950 345.600 862.050 346.050 ;
        RECT 844.950 344.400 862.050 345.600 ;
        RECT 844.950 343.950 847.050 344.400 ;
        RECT 859.950 343.950 862.050 344.400 ;
        RECT 889.950 345.600 892.050 346.050 ;
        RECT 895.950 345.600 898.050 346.050 ;
        RECT 889.950 344.400 898.050 345.600 ;
        RECT 889.950 343.950 892.050 344.400 ;
        RECT 895.950 343.950 898.050 344.400 ;
        RECT 676.950 341.400 699.600 342.600 ;
        RECT 724.950 342.600 727.050 343.050 ;
        RECT 736.950 342.600 739.050 343.050 ;
        RECT 724.950 341.400 739.050 342.600 ;
        RECT 676.950 340.950 679.050 341.400 ;
        RECT 724.950 340.950 727.050 341.400 ;
        RECT 736.950 340.950 739.050 341.400 ;
        RECT 772.950 342.600 775.050 343.050 ;
        RECT 799.950 342.600 802.050 343.050 ;
        RECT 826.950 342.600 829.050 343.050 ;
        RECT 838.950 342.600 841.050 343.050 ;
        RECT 772.950 341.400 798.600 342.600 ;
        RECT 772.950 340.950 775.050 341.400 ;
        RECT 127.950 339.600 130.050 340.200 ;
        RECT 151.950 339.600 154.050 340.200 ;
        RECT 121.950 339.000 130.050 339.600 ;
        RECT 122.400 338.400 130.050 339.000 ;
        RECT 103.950 338.100 106.050 338.400 ;
        RECT 115.950 337.950 118.050 338.400 ;
        RECT 127.950 338.100 130.050 338.400 ;
        RECT 131.400 338.400 154.050 339.600 ;
        RECT 59.400 335.400 108.600 336.600 ;
        RECT 22.950 333.600 25.050 334.050 ;
        RECT 59.400 333.900 60.600 335.400 ;
        RECT 107.400 333.900 108.600 335.400 ;
        RECT 131.400 333.900 132.600 338.400 ;
        RECT 151.950 338.100 154.050 338.400 ;
        RECT 163.950 339.600 166.050 340.050 ;
        RECT 172.950 339.600 175.050 340.200 ;
        RECT 163.950 338.400 175.050 339.600 ;
        RECT 163.950 337.950 166.050 338.400 ;
        RECT 172.950 338.100 175.050 338.400 ;
        RECT 223.950 339.750 226.050 340.200 ;
        RECT 235.950 339.750 238.050 340.200 ;
        RECT 223.950 338.550 238.050 339.750 ;
        RECT 223.950 338.100 226.050 338.550 ;
        RECT 235.950 338.100 238.050 338.550 ;
        RECT 250.950 339.750 253.050 340.200 ;
        RECT 262.950 339.750 265.050 340.200 ;
        RECT 250.950 338.550 265.050 339.750 ;
        RECT 250.950 338.100 253.050 338.550 ;
        RECT 262.950 338.100 265.050 338.550 ;
        RECT 271.950 339.600 274.050 340.200 ;
        RECT 304.950 339.600 307.050 340.050 ;
        RECT 271.950 338.400 307.050 339.600 ;
        RECT 313.950 339.600 316.050 340.500 ;
        RECT 328.950 339.600 331.050 340.200 ;
        RECT 313.950 338.400 331.050 339.600 ;
        RECT 271.950 338.100 274.050 338.400 ;
        RECT 304.950 337.950 307.050 338.400 ;
        RECT 328.950 338.100 331.050 338.400 ;
        RECT 367.950 339.600 370.050 340.050 ;
        RECT 394.950 339.750 397.050 340.200 ;
        RECT 403.950 339.750 406.050 340.200 ;
        RECT 394.950 339.600 406.050 339.750 ;
        RECT 367.950 338.550 406.050 339.600 ;
        RECT 367.950 338.400 397.050 338.550 ;
        RECT 367.950 337.950 370.050 338.400 ;
        RECT 394.950 338.100 397.050 338.400 ;
        RECT 403.950 338.100 406.050 338.550 ;
        RECT 415.950 339.750 418.050 340.200 ;
        RECT 424.950 339.750 427.050 340.200 ;
        RECT 415.950 338.550 427.050 339.750 ;
        RECT 415.950 338.100 418.050 338.550 ;
        RECT 424.950 338.100 427.050 338.550 ;
        RECT 502.950 339.600 505.050 340.200 ;
        RECT 517.950 339.750 520.050 340.200 ;
        RECT 532.950 339.750 535.050 340.050 ;
        RECT 502.950 338.400 516.600 339.600 ;
        RECT 502.950 338.100 505.050 338.400 ;
        RECT 515.400 336.600 516.600 338.400 ;
        RECT 517.950 338.550 535.050 339.750 ;
        RECT 517.950 338.100 520.050 338.550 ;
        RECT 532.950 337.950 535.050 338.550 ;
        RECT 547.950 339.600 550.050 340.200 ;
        RECT 625.950 339.600 628.050 340.200 ;
        RECT 637.950 339.600 640.050 340.050 ;
        RECT 646.950 339.600 649.050 340.200 ;
        RECT 547.950 338.400 570.600 339.600 ;
        RECT 547.950 338.100 550.050 338.400 ;
        RECT 532.950 336.600 535.050 336.900 ;
        RECT 515.400 335.400 535.050 336.600 ;
        RECT 532.950 334.800 535.050 335.400 ;
        RECT 4.950 332.400 25.050 333.600 ;
        RECT 4.950 331.500 7.050 332.400 ;
        RECT 22.950 331.950 25.050 332.400 ;
        RECT 52.950 333.450 55.050 333.900 ;
        RECT 58.950 333.450 61.050 333.900 ;
        RECT 52.950 332.250 61.050 333.450 ;
        RECT 52.950 331.800 55.050 332.250 ;
        RECT 58.950 331.800 61.050 332.250 ;
        RECT 73.950 333.450 76.050 333.900 ;
        RECT 94.950 333.450 97.050 333.900 ;
        RECT 73.950 332.250 97.050 333.450 ;
        RECT 73.950 331.800 76.050 332.250 ;
        RECT 94.950 331.800 97.050 332.250 ;
        RECT 106.950 331.800 109.050 333.900 ;
        RECT 115.950 333.450 118.050 333.900 ;
        RECT 124.950 333.450 127.050 333.900 ;
        RECT 115.950 332.250 127.050 333.450 ;
        RECT 115.950 331.800 118.050 332.250 ;
        RECT 124.950 331.800 127.050 332.250 ;
        RECT 130.950 331.800 133.050 333.900 ;
        RECT 232.950 333.600 235.050 333.900 ;
        RECT 253.950 333.600 256.050 333.900 ;
        RECT 298.950 333.600 301.050 334.050 ;
        RECT 304.950 333.600 307.050 333.900 ;
        RECT 232.950 332.400 256.050 333.600 ;
        RECT 232.950 331.800 235.050 332.400 ;
        RECT 253.950 331.800 256.050 332.400 ;
        RECT 280.950 333.150 283.050 333.600 ;
        RECT 286.950 333.150 289.050 333.600 ;
        RECT 280.950 331.950 289.050 333.150 ;
        RECT 298.950 333.450 307.050 333.600 ;
        RECT 331.950 333.450 334.050 333.900 ;
        RECT 298.950 332.400 334.050 333.450 ;
        RECT 298.950 331.950 301.050 332.400 ;
        RECT 304.950 332.250 334.050 332.400 ;
        RECT 280.950 331.500 283.050 331.950 ;
        RECT 286.950 331.500 289.050 331.950 ;
        RECT 304.950 331.800 307.050 332.250 ;
        RECT 331.950 331.800 334.050 332.250 ;
        RECT 391.950 333.600 394.050 333.900 ;
        RECT 412.950 333.600 415.050 333.900 ;
        RECT 391.950 332.400 415.050 333.600 ;
        RECT 391.950 331.800 394.050 332.400 ;
        RECT 412.950 331.800 415.050 332.400 ;
        RECT 448.950 333.600 451.050 334.050 ;
        RECT 466.950 333.600 469.050 334.050 ;
        RECT 448.950 332.400 469.050 333.600 ;
        RECT 448.950 331.950 451.050 332.400 ;
        RECT 466.950 331.950 469.050 332.400 ;
        RECT 499.950 333.450 502.050 333.900 ;
        RECT 508.950 333.450 511.050 333.900 ;
        RECT 499.950 332.250 511.050 333.450 ;
        RECT 499.950 331.800 502.050 332.250 ;
        RECT 508.950 331.800 511.050 332.250 ;
        RECT 535.950 333.450 538.050 333.900 ;
        RECT 544.950 333.450 547.050 333.900 ;
        RECT 535.950 332.250 547.050 333.450 ;
        RECT 535.950 331.800 538.050 332.250 ;
        RECT 544.950 331.800 547.050 332.250 ;
        RECT 550.950 333.450 553.050 333.900 ;
        RECT 556.950 333.450 559.050 334.050 ;
        RECT 569.400 333.900 570.600 338.400 ;
        RECT 625.950 338.400 636.600 339.600 ;
        RECT 625.950 338.100 628.050 338.400 ;
        RECT 635.400 336.600 636.600 338.400 ;
        RECT 637.950 338.400 649.050 339.600 ;
        RECT 637.950 337.950 640.050 338.400 ;
        RECT 646.950 338.100 649.050 338.400 ;
        RECT 670.950 338.100 673.050 340.200 ;
        RECT 700.950 339.600 703.050 340.200 ;
        RECT 718.950 339.600 721.050 340.200 ;
        RECT 700.950 338.400 721.050 339.600 ;
        RECT 700.950 338.100 703.050 338.400 ;
        RECT 718.950 338.100 721.050 338.400 ;
        RECT 730.950 339.600 733.050 340.050 ;
        RECT 742.950 339.600 745.050 340.200 ;
        RECT 769.950 339.600 772.050 340.200 ;
        RECT 730.950 338.400 745.050 339.600 ;
        RECT 661.950 336.600 664.050 337.050 ;
        RECT 671.400 336.600 672.600 338.100 ;
        RECT 730.950 337.950 733.050 338.400 ;
        RECT 742.950 338.100 745.050 338.400 ;
        RECT 752.400 338.400 772.050 339.600 ;
        RECT 635.400 335.400 654.600 336.600 ;
        RECT 550.950 332.250 559.050 333.450 ;
        RECT 550.950 331.800 553.050 332.250 ;
        RECT 556.950 331.950 559.050 332.250 ;
        RECT 568.950 331.800 571.050 333.900 ;
        RECT 616.950 333.450 619.050 333.900 ;
        RECT 628.950 333.450 631.050 333.900 ;
        RECT 616.950 332.250 631.050 333.450 ;
        RECT 616.950 331.800 619.050 332.250 ;
        RECT 628.950 331.800 631.050 332.250 ;
        RECT 37.950 330.600 40.050 331.050 ;
        RECT 46.950 330.600 49.050 331.050 ;
        RECT 37.950 329.400 49.050 330.600 ;
        RECT 37.950 328.950 40.050 329.400 ;
        RECT 46.950 328.950 49.050 329.400 ;
        RECT 148.950 330.600 151.050 331.050 ;
        RECT 163.950 330.600 166.050 331.050 ;
        RECT 148.950 329.400 166.050 330.600 ;
        RECT 148.950 328.950 151.050 329.400 ;
        RECT 163.950 328.950 166.050 329.400 ;
        RECT 211.950 330.600 214.050 331.050 ;
        RECT 223.950 330.600 226.050 331.050 ;
        RECT 229.950 330.600 232.050 331.050 ;
        RECT 247.950 330.600 250.050 331.050 ;
        RECT 211.950 329.400 250.050 330.600 ;
        RECT 211.950 328.950 214.050 329.400 ;
        RECT 223.950 328.950 226.050 329.400 ;
        RECT 229.950 328.950 232.050 329.400 ;
        RECT 247.950 328.950 250.050 329.400 ;
        RECT 256.950 330.600 259.050 331.050 ;
        RECT 265.950 330.600 268.050 331.050 ;
        RECT 256.950 329.400 268.050 330.600 ;
        RECT 256.950 328.950 259.050 329.400 ;
        RECT 265.950 328.950 268.050 329.400 ;
        RECT 478.950 330.600 481.050 331.050 ;
        RECT 493.950 330.600 496.050 331.050 ;
        RECT 478.950 329.400 496.050 330.600 ;
        RECT 478.950 328.950 481.050 329.400 ;
        RECT 493.950 328.950 496.050 329.400 ;
        RECT 520.950 330.600 523.050 331.050 ;
        RECT 536.400 330.600 537.600 331.800 ;
        RECT 653.400 331.050 654.600 335.400 ;
        RECT 661.950 335.400 672.600 336.600 ;
        RECT 661.950 334.950 664.050 335.400 ;
        RECT 752.400 333.900 753.600 338.400 ;
        RECT 769.950 338.100 772.050 338.400 ;
        RECT 787.950 339.600 790.050 340.050 ;
        RECT 793.950 339.600 796.050 340.050 ;
        RECT 787.950 338.400 796.050 339.600 ;
        RECT 787.950 337.950 790.050 338.400 ;
        RECT 793.950 337.950 796.050 338.400 ;
        RECT 797.400 333.900 798.600 341.400 ;
        RECT 799.950 341.400 841.050 342.600 ;
        RECT 799.950 340.950 802.050 341.400 ;
        RECT 826.950 340.950 829.050 341.400 ;
        RECT 838.950 340.950 841.050 341.400 ;
        RECT 802.950 337.950 805.050 340.050 ;
        RECT 814.950 339.600 817.050 340.050 ;
        RECT 814.950 338.400 822.600 339.600 ;
        RECT 814.950 337.950 817.050 338.400 ;
        RECT 803.400 334.050 804.600 337.950 ;
        RECT 673.950 333.450 676.050 333.900 ;
        RECT 688.950 333.450 691.050 333.900 ;
        RECT 673.950 332.250 691.050 333.450 ;
        RECT 673.950 331.800 676.050 332.250 ;
        RECT 688.950 331.800 691.050 332.250 ;
        RECT 703.950 333.600 706.050 333.900 ;
        RECT 715.950 333.600 718.050 333.900 ;
        RECT 703.950 332.400 718.050 333.600 ;
        RECT 703.950 331.800 706.050 332.400 ;
        RECT 715.950 331.800 718.050 332.400 ;
        RECT 721.950 333.450 724.050 333.900 ;
        RECT 730.950 333.450 733.050 333.900 ;
        RECT 721.950 332.250 733.050 333.450 ;
        RECT 721.950 331.800 724.050 332.250 ;
        RECT 730.950 331.800 733.050 332.250 ;
        RECT 751.950 331.800 754.050 333.900 ;
        RECT 760.950 333.450 763.050 333.900 ;
        RECT 766.950 333.450 769.050 333.900 ;
        RECT 760.950 332.250 769.050 333.450 ;
        RECT 760.950 331.800 763.050 332.250 ;
        RECT 766.950 331.800 769.050 332.250 ;
        RECT 772.950 333.600 775.050 333.900 ;
        RECT 781.950 333.600 784.050 333.900 ;
        RECT 772.950 333.450 784.050 333.600 ;
        RECT 790.950 333.450 793.050 333.900 ;
        RECT 772.950 332.400 793.050 333.450 ;
        RECT 772.950 331.800 775.050 332.400 ;
        RECT 781.950 332.250 793.050 332.400 ;
        RECT 781.950 331.800 784.050 332.250 ;
        RECT 790.950 331.800 793.050 332.250 ;
        RECT 796.950 331.800 799.050 333.900 ;
        RECT 802.950 331.950 805.050 334.050 ;
        RECT 821.400 331.050 822.600 338.400 ;
        RECT 835.950 336.600 838.050 340.050 ;
        RECT 844.950 339.600 847.050 340.200 ;
        RECT 853.950 339.600 856.050 340.050 ;
        RECT 844.950 338.400 856.050 339.600 ;
        RECT 844.950 338.100 847.050 338.400 ;
        RECT 853.950 337.950 856.050 338.400 ;
        RECT 859.950 336.600 862.050 340.050 ;
        RECT 865.800 338.100 867.900 340.200 ;
        RECT 871.950 339.600 874.050 340.200 ;
        RECT 889.950 339.600 892.050 340.050 ;
        RECT 871.950 338.400 892.050 339.600 ;
        RECT 871.950 338.100 874.050 338.400 ;
        RECT 835.950 336.000 840.600 336.600 ;
        RECT 859.950 336.000 864.600 336.600 ;
        RECT 836.400 335.400 840.600 336.000 ;
        RECT 860.400 335.400 864.600 336.000 ;
        RECT 823.950 333.600 826.050 333.900 ;
        RECT 839.400 333.600 840.600 335.400 ;
        RECT 863.400 333.900 864.600 335.400 ;
        RECT 841.950 333.600 844.050 333.900 ;
        RECT 823.950 332.400 844.050 333.600 ;
        RECT 823.950 331.800 826.050 332.400 ;
        RECT 841.950 331.800 844.050 332.400 ;
        RECT 862.950 331.800 865.050 333.900 ;
        RECT 866.250 331.050 867.450 338.100 ;
        RECT 889.950 337.950 892.050 338.400 ;
        RECT 520.950 329.400 537.600 330.600 ;
        RECT 547.950 330.600 550.050 331.050 ;
        RECT 562.950 330.600 565.050 331.050 ;
        RECT 547.950 329.400 565.050 330.600 ;
        RECT 520.950 328.950 523.050 329.400 ;
        RECT 547.950 328.950 550.050 329.400 ;
        RECT 562.950 328.950 565.050 329.400 ;
        RECT 652.950 328.950 655.050 331.050 ;
        RECT 820.950 328.950 823.050 331.050 ;
        RECT 865.800 328.950 867.900 331.050 ;
        RECT 868.950 330.600 871.050 331.050 ;
        RECT 877.950 330.600 880.050 331.050 ;
        RECT 868.950 329.400 880.050 330.600 ;
        RECT 868.950 328.950 871.050 329.400 ;
        RECT 877.950 328.950 880.050 329.400 ;
        RECT 73.950 327.600 76.050 328.050 ;
        RECT 79.950 327.600 82.050 328.050 ;
        RECT 73.950 326.400 82.050 327.600 ;
        RECT 73.950 325.950 76.050 326.400 ;
        RECT 79.950 325.950 82.050 326.400 ;
        RECT 175.950 327.600 178.050 328.050 ;
        RECT 199.950 327.600 202.050 328.050 ;
        RECT 175.950 326.400 202.050 327.600 ;
        RECT 175.950 325.950 178.050 326.400 ;
        RECT 199.950 325.950 202.050 326.400 ;
        RECT 538.950 327.600 541.050 328.050 ;
        RECT 574.950 327.600 577.050 328.050 ;
        RECT 622.950 327.600 625.050 328.050 ;
        RECT 655.950 327.600 658.050 328.050 ;
        RECT 538.950 326.400 658.050 327.600 ;
        RECT 538.950 325.950 541.050 326.400 ;
        RECT 574.950 325.950 577.050 326.400 ;
        RECT 622.950 325.950 625.050 326.400 ;
        RECT 655.950 325.950 658.050 326.400 ;
        RECT 676.950 327.600 679.050 328.050 ;
        RECT 745.950 327.600 748.050 328.050 ;
        RECT 778.950 327.600 781.050 328.050 ;
        RECT 676.950 326.400 781.050 327.600 ;
        RECT 676.950 325.950 679.050 326.400 ;
        RECT 745.950 325.950 748.050 326.400 ;
        RECT 778.950 325.950 781.050 326.400 ;
        RECT 64.950 324.600 67.050 325.050 ;
        RECT 85.950 324.600 88.050 325.050 ;
        RECT 91.950 324.600 94.050 325.050 ;
        RECT 148.950 324.600 151.050 325.050 ;
        RECT 211.950 324.600 214.050 325.050 ;
        RECT 64.950 323.400 214.050 324.600 ;
        RECT 64.950 322.950 67.050 323.400 ;
        RECT 85.950 322.950 88.050 323.400 ;
        RECT 91.950 322.950 94.050 323.400 ;
        RECT 148.950 322.950 151.050 323.400 ;
        RECT 211.950 322.950 214.050 323.400 ;
        RECT 217.950 324.600 220.050 325.050 ;
        RECT 274.950 324.600 277.050 325.050 ;
        RECT 217.950 323.400 277.050 324.600 ;
        RECT 217.950 322.950 220.050 323.400 ;
        RECT 274.950 322.950 277.050 323.400 ;
        RECT 424.950 324.600 427.050 325.050 ;
        RECT 445.950 324.600 448.050 325.050 ;
        RECT 478.950 324.600 481.050 325.050 ;
        RECT 424.950 323.400 481.050 324.600 ;
        RECT 424.950 322.950 427.050 323.400 ;
        RECT 445.950 322.950 448.050 323.400 ;
        RECT 478.950 322.950 481.050 323.400 ;
        RECT 568.950 324.600 571.050 325.050 ;
        RECT 649.950 324.600 652.050 325.050 ;
        RECT 667.950 324.600 670.050 325.050 ;
        RECT 568.950 323.400 670.050 324.600 ;
        RECT 568.950 322.950 571.050 323.400 ;
        RECT 649.950 322.950 652.050 323.400 ;
        RECT 667.950 322.950 670.050 323.400 ;
        RECT 697.950 324.600 700.050 325.050 ;
        RECT 745.950 324.600 748.050 324.900 ;
        RECT 802.950 324.600 805.050 325.050 ;
        RECT 697.950 323.400 805.050 324.600 ;
        RECT 697.950 322.950 700.050 323.400 ;
        RECT 745.950 322.800 748.050 323.400 ;
        RECT 802.950 322.950 805.050 323.400 ;
        RECT 76.950 321.600 79.050 322.050 ;
        RECT 44.400 320.400 79.050 321.600 ;
        RECT 44.400 319.050 45.600 320.400 ;
        RECT 76.950 319.950 79.050 320.400 ;
        RECT 154.950 321.600 157.050 322.050 ;
        RECT 181.950 321.600 184.050 322.050 ;
        RECT 154.950 320.400 184.050 321.600 ;
        RECT 154.950 319.950 157.050 320.400 ;
        RECT 181.950 319.950 184.050 320.400 ;
        RECT 400.950 321.600 403.050 322.050 ;
        RECT 436.950 321.600 439.050 322.050 ;
        RECT 457.950 321.600 460.050 322.050 ;
        RECT 400.950 320.400 460.050 321.600 ;
        RECT 400.950 319.950 403.050 320.400 ;
        RECT 436.950 319.950 439.050 320.400 ;
        RECT 457.950 319.950 460.050 320.400 ;
        RECT 763.950 321.600 766.050 322.050 ;
        RECT 799.950 321.600 802.050 322.050 ;
        RECT 763.950 320.400 802.050 321.600 ;
        RECT 763.950 319.950 766.050 320.400 ;
        RECT 799.950 319.950 802.050 320.400 ;
        RECT 40.950 317.400 45.600 319.050 ;
        RECT 403.950 318.600 406.050 319.050 ;
        RECT 418.950 318.600 421.050 319.050 ;
        RECT 433.950 318.600 436.050 319.050 ;
        RECT 403.950 317.400 436.050 318.600 ;
        RECT 40.950 316.950 45.000 317.400 ;
        RECT 403.950 316.950 406.050 317.400 ;
        RECT 418.950 316.950 421.050 317.400 ;
        RECT 433.950 316.950 436.050 317.400 ;
        RECT 817.950 318.600 820.050 319.050 ;
        RECT 868.950 318.600 871.050 319.050 ;
        RECT 817.950 317.400 871.050 318.600 ;
        RECT 817.950 316.950 820.050 317.400 ;
        RECT 868.950 316.950 871.050 317.400 ;
        RECT 73.950 315.600 76.050 316.050 ;
        RECT 139.950 315.600 142.050 316.050 ;
        RECT 304.950 315.600 307.050 316.050 ;
        RECT 73.950 314.400 307.050 315.600 ;
        RECT 73.950 313.950 76.050 314.400 ;
        RECT 139.950 313.950 142.050 314.400 ;
        RECT 304.950 313.950 307.050 314.400 ;
        RECT 586.950 315.600 589.050 316.050 ;
        RECT 619.950 315.600 622.050 316.050 ;
        RECT 586.950 314.400 622.050 315.600 ;
        RECT 586.950 313.950 589.050 314.400 ;
        RECT 619.950 313.950 622.050 314.400 ;
        RECT 637.950 315.600 640.050 316.050 ;
        RECT 703.950 315.600 706.050 316.050 ;
        RECT 637.950 314.400 706.050 315.600 ;
        RECT 637.950 313.950 640.050 314.400 ;
        RECT 703.950 313.950 706.050 314.400 ;
        RECT 778.950 315.600 781.050 316.050 ;
        RECT 811.950 315.600 814.050 316.050 ;
        RECT 778.950 314.400 814.050 315.600 ;
        RECT 778.950 313.950 781.050 314.400 ;
        RECT 811.950 313.950 814.050 314.400 ;
        RECT 235.950 312.600 238.050 313.050 ;
        RECT 241.950 312.600 244.050 313.050 ;
        RECT 235.950 311.400 244.050 312.600 ;
        RECT 235.950 310.950 238.050 311.400 ;
        RECT 241.950 310.950 244.050 311.400 ;
        RECT 583.950 312.600 586.050 313.050 ;
        RECT 625.950 312.600 628.050 313.050 ;
        RECT 685.950 312.600 688.050 313.050 ;
        RECT 583.950 311.400 628.050 312.600 ;
        RECT 583.950 310.950 586.050 311.400 ;
        RECT 625.950 310.950 628.050 311.400 ;
        RECT 629.400 311.400 688.050 312.600 ;
        RECT 76.950 309.600 79.050 310.050 ;
        RECT 100.950 309.600 103.050 310.050 ;
        RECT 76.950 308.400 103.050 309.600 ;
        RECT 76.950 307.950 79.050 308.400 ;
        RECT 100.950 307.950 103.050 308.400 ;
        RECT 109.950 309.600 112.050 310.050 ;
        RECT 118.950 309.600 121.050 310.050 ;
        RECT 109.950 308.400 121.050 309.600 ;
        RECT 109.950 307.950 112.050 308.400 ;
        RECT 118.950 307.950 121.050 308.400 ;
        RECT 190.950 309.600 193.050 310.050 ;
        RECT 196.950 309.600 199.050 310.050 ;
        RECT 214.950 309.600 217.050 310.050 ;
        RECT 190.950 308.400 217.050 309.600 ;
        RECT 190.950 307.950 193.050 308.400 ;
        RECT 196.950 307.950 199.050 308.400 ;
        RECT 214.950 307.950 217.050 308.400 ;
        RECT 370.950 309.600 373.050 310.050 ;
        RECT 379.950 309.600 382.050 310.050 ;
        RECT 370.950 308.400 382.050 309.600 ;
        RECT 370.950 307.950 373.050 308.400 ;
        RECT 379.950 307.950 382.050 308.400 ;
        RECT 595.950 309.600 598.050 310.050 ;
        RECT 629.400 309.600 630.600 311.400 ;
        RECT 685.950 310.950 688.050 311.400 ;
        RECT 859.950 312.600 862.050 313.050 ;
        RECT 880.950 312.600 883.050 313.050 ;
        RECT 859.950 311.400 883.050 312.600 ;
        RECT 859.950 310.950 862.050 311.400 ;
        RECT 880.950 310.950 883.050 311.400 ;
        RECT 595.950 308.400 630.600 309.600 ;
        RECT 652.950 309.600 655.050 310.050 ;
        RECT 751.950 309.600 754.050 310.050 ;
        RECT 652.950 308.400 754.050 309.600 ;
        RECT 595.950 307.950 598.050 308.400 ;
        RECT 652.950 307.950 655.050 308.400 ;
        RECT 751.950 307.950 754.050 308.400 ;
        RECT 1.950 306.600 4.050 307.050 ;
        RECT 13.950 306.600 16.050 307.050 ;
        RECT 1.950 305.400 16.050 306.600 ;
        RECT 1.950 304.950 4.050 305.400 ;
        RECT 13.950 304.950 16.050 305.400 ;
        RECT 241.950 306.600 244.050 307.050 ;
        RECT 292.950 306.600 295.050 307.050 ;
        RECT 829.950 306.600 832.050 307.050 ;
        RECT 241.950 305.400 295.050 306.600 ;
        RECT 241.950 304.950 244.050 305.400 ;
        RECT 292.950 304.950 295.050 305.400 ;
        RECT 806.400 305.400 832.050 306.600 ;
        RECT 806.400 304.050 807.600 305.400 ;
        RECT 829.950 304.950 832.050 305.400 ;
        RECT 853.950 306.600 856.050 307.050 ;
        RECT 868.950 306.600 871.050 307.050 ;
        RECT 853.950 305.400 871.050 306.600 ;
        RECT 853.950 304.950 856.050 305.400 ;
        RECT 868.950 304.950 871.050 305.400 ;
        RECT 127.950 303.600 130.050 304.050 ;
        RECT 142.950 303.600 145.050 304.050 ;
        RECT 127.950 302.400 145.050 303.600 ;
        RECT 127.950 301.950 130.050 302.400 ;
        RECT 142.950 301.950 145.050 302.400 ;
        RECT 340.950 303.600 343.050 304.050 ;
        RECT 397.950 303.600 400.050 304.050 ;
        RECT 340.950 302.400 400.050 303.600 ;
        RECT 340.950 301.950 343.050 302.400 ;
        RECT 397.950 301.950 400.050 302.400 ;
        RECT 442.950 303.600 445.050 304.050 ;
        RECT 469.950 303.600 472.050 304.050 ;
        RECT 442.950 302.400 472.050 303.600 ;
        RECT 442.950 301.950 445.050 302.400 ;
        RECT 469.950 301.950 472.050 302.400 ;
        RECT 652.950 303.600 655.050 304.050 ;
        RECT 715.950 303.600 718.050 304.050 ;
        RECT 652.950 302.400 718.050 303.600 ;
        RECT 652.950 301.950 655.050 302.400 ;
        RECT 715.950 301.950 718.050 302.400 ;
        RECT 757.950 303.600 760.050 304.050 ;
        RECT 775.950 303.600 778.050 304.050 ;
        RECT 757.950 302.400 778.050 303.600 ;
        RECT 757.950 301.950 760.050 302.400 ;
        RECT 775.950 301.950 778.050 302.400 ;
        RECT 790.950 303.600 793.050 304.050 ;
        RECT 805.950 303.600 808.050 304.050 ;
        RECT 790.950 302.400 808.050 303.600 ;
        RECT 790.950 301.950 793.050 302.400 ;
        RECT 805.950 301.950 808.050 302.400 ;
        RECT 832.950 303.600 835.050 304.050 ;
        RECT 847.950 303.600 850.050 304.050 ;
        RECT 832.950 302.400 850.050 303.600 ;
        RECT 832.950 301.950 835.050 302.400 ;
        RECT 847.950 301.950 850.050 302.400 ;
        RECT 853.950 303.600 856.050 303.900 ;
        RECT 886.950 303.600 889.050 304.050 ;
        RECT 853.950 302.400 889.050 303.600 ;
        RECT 853.950 301.800 856.050 302.400 ;
        RECT 886.950 301.950 889.050 302.400 ;
        RECT 70.950 300.600 73.050 301.050 ;
        RECT 85.950 300.600 88.050 301.050 ;
        RECT 70.950 299.400 88.050 300.600 ;
        RECT 70.950 298.950 73.050 299.400 ;
        RECT 85.950 298.950 88.050 299.400 ;
        RECT 265.950 300.600 268.050 301.050 ;
        RECT 283.950 300.600 286.050 301.050 ;
        RECT 265.950 299.400 286.050 300.600 ;
        RECT 265.950 298.950 268.050 299.400 ;
        RECT 283.950 298.950 286.050 299.400 ;
        RECT 292.950 300.600 295.050 301.050 ;
        RECT 298.950 300.600 301.050 301.050 ;
        RECT 292.950 299.400 301.050 300.600 ;
        RECT 292.950 298.950 295.050 299.400 ;
        RECT 298.950 298.950 301.050 299.400 ;
        RECT 319.950 300.600 322.050 301.050 ;
        RECT 331.950 300.600 334.050 301.050 ;
        RECT 319.950 299.400 334.050 300.600 ;
        RECT 319.950 298.950 322.050 299.400 ;
        RECT 331.950 298.950 334.050 299.400 ;
        RECT 463.950 300.600 466.050 301.050 ;
        RECT 472.950 300.600 475.050 301.050 ;
        RECT 463.950 299.400 475.050 300.600 ;
        RECT 463.950 298.950 466.050 299.400 ;
        RECT 472.950 298.950 475.050 299.400 ;
        RECT 550.950 300.600 553.050 301.050 ;
        RECT 589.950 300.600 592.050 301.050 ;
        RECT 550.950 299.400 592.050 300.600 ;
        RECT 550.950 298.950 553.050 299.400 ;
        RECT 589.950 298.950 592.050 299.400 ;
        RECT 736.950 300.600 739.050 301.050 ;
        RECT 754.950 300.600 757.050 301.050 ;
        RECT 736.950 299.400 757.050 300.600 ;
        RECT 736.950 298.950 739.050 299.400 ;
        RECT 754.950 298.950 757.050 299.400 ;
        RECT 808.950 300.600 811.050 301.050 ;
        RECT 817.950 300.600 820.050 301.050 ;
        RECT 808.950 299.400 820.050 300.600 ;
        RECT 808.950 298.950 811.050 299.400 ;
        RECT 817.950 298.950 820.050 299.400 ;
        RECT 883.950 298.950 886.050 301.050 ;
        RECT 133.950 297.600 136.050 298.050 ;
        RECT 169.950 297.600 172.050 298.050 ;
        RECT 133.950 296.400 172.050 297.600 ;
        RECT 133.950 295.950 136.050 296.400 ;
        RECT 169.950 295.950 172.050 296.400 ;
        RECT 295.950 295.950 298.050 298.050 ;
        RECT 379.950 297.600 382.050 298.050 ;
        RECT 451.950 297.600 454.050 298.050 ;
        RECT 496.950 297.600 499.050 298.050 ;
        RECT 379.950 296.400 499.050 297.600 ;
        RECT 379.950 295.950 382.050 296.400 ;
        RECT 451.950 295.950 454.050 296.400 ;
        RECT 496.950 295.950 499.050 296.400 ;
        RECT 703.950 297.600 706.050 298.050 ;
        RECT 709.950 297.600 712.050 298.050 ;
        RECT 760.950 297.600 763.050 298.050 ;
        RECT 703.950 296.400 763.050 297.600 ;
        RECT 703.950 295.950 706.050 296.400 ;
        RECT 709.950 295.950 712.050 296.400 ;
        RECT 760.950 295.950 763.050 296.400 ;
        RECT 784.950 297.600 787.050 298.050 ;
        RECT 802.950 297.600 805.050 298.050 ;
        RECT 823.950 297.600 826.050 298.050 ;
        RECT 784.950 296.400 826.050 297.600 ;
        RECT 784.950 295.950 787.050 296.400 ;
        RECT 802.950 295.950 805.050 296.400 ;
        RECT 823.950 295.950 826.050 296.400 ;
        RECT 850.950 297.600 853.050 298.050 ;
        RECT 856.950 297.600 859.050 298.050 ;
        RECT 850.950 296.400 859.050 297.600 ;
        RECT 850.950 295.950 853.050 296.400 ;
        RECT 856.950 295.950 859.050 296.400 ;
        RECT 865.950 297.600 868.050 298.050 ;
        RECT 871.950 297.600 874.050 298.050 ;
        RECT 865.950 296.400 874.050 297.600 ;
        RECT 865.950 295.950 868.050 296.400 ;
        RECT 871.950 295.950 874.050 296.400 ;
        RECT 52.950 294.600 55.050 295.200 ;
        RECT 79.950 294.600 82.050 295.200 ;
        RECT 142.950 295.050 145.050 295.500 ;
        RECT 151.950 295.050 154.050 295.500 ;
        RECT 106.950 294.600 109.050 295.050 ;
        RECT 52.950 293.400 109.050 294.600 ;
        RECT 142.950 293.850 154.050 295.050 ;
        RECT 142.950 293.400 145.050 293.850 ;
        RECT 151.950 293.400 154.050 293.850 ;
        RECT 169.950 293.400 172.050 295.500 ;
        RECT 274.950 295.050 277.050 295.500 ;
        RECT 280.950 295.050 283.050 295.500 ;
        RECT 274.950 293.850 283.050 295.050 ;
        RECT 274.950 293.400 277.050 293.850 ;
        RECT 280.950 293.400 283.050 293.850 ;
        RECT 52.950 293.100 55.050 293.400 ;
        RECT 79.950 293.100 82.050 293.400 ;
        RECT 106.950 292.950 109.050 293.400 ;
        RECT 46.950 291.600 49.050 292.050 ;
        RECT 46.950 290.400 57.600 291.600 ;
        RECT 46.950 289.950 49.050 290.400 ;
        RECT 56.400 288.900 57.600 290.400 ;
        RECT 170.400 289.050 171.600 293.400 ;
        RECT 55.950 286.800 58.050 288.900 ;
        RECT 88.950 288.600 91.050 288.900 ;
        RECT 77.400 288.000 100.050 288.600 ;
        RECT 76.950 287.400 100.050 288.000 ;
        RECT 43.950 285.600 46.050 286.050 ;
        RECT 61.950 285.600 64.050 286.050 ;
        RECT 43.950 284.400 64.050 285.600 ;
        RECT 43.950 283.950 46.050 284.400 ;
        RECT 61.950 283.950 64.050 284.400 ;
        RECT 76.950 283.950 79.050 287.400 ;
        RECT 88.950 286.800 91.050 287.400 ;
        RECT 97.950 286.500 100.050 287.400 ;
        RECT 166.950 287.400 171.600 289.050 ;
        RECT 226.950 288.600 229.050 289.050 ;
        RECT 238.950 288.600 241.050 288.900 ;
        RECT 256.950 288.600 259.050 289.050 ;
        RECT 296.400 288.900 297.600 295.950 ;
        RECT 307.950 294.750 310.050 295.200 ;
        RECT 316.950 294.750 319.050 295.200 ;
        RECT 307.950 293.550 319.050 294.750 ;
        RECT 307.950 293.100 310.050 293.550 ;
        RECT 316.950 293.100 319.050 293.550 ;
        RECT 322.950 293.100 325.050 295.200 ;
        RECT 367.950 293.400 370.050 295.500 ;
        RECT 385.950 294.600 388.050 295.050 ;
        RECT 403.950 294.600 406.050 295.200 ;
        RECT 385.950 293.400 406.050 294.600 ;
        RECT 226.950 287.400 241.050 288.600 ;
        RECT 166.950 286.950 171.000 287.400 ;
        RECT 226.950 286.950 229.050 287.400 ;
        RECT 238.950 286.800 241.050 287.400 ;
        RECT 247.950 287.400 259.050 288.600 ;
        RECT 247.950 286.500 250.050 287.400 ;
        RECT 256.950 286.950 259.050 287.400 ;
        RECT 295.950 286.800 298.050 288.900 ;
        RECT 310.950 288.600 313.050 289.050 ;
        RECT 319.950 288.600 322.050 288.900 ;
        RECT 310.950 287.400 322.050 288.600 ;
        RECT 323.400 288.600 324.600 293.100 ;
        RECT 337.950 288.600 340.050 288.900 ;
        RECT 368.400 288.600 369.600 293.400 ;
        RECT 385.950 292.950 388.050 293.400 ;
        RECT 403.950 293.100 406.050 293.400 ;
        RECT 421.950 294.600 424.050 295.200 ;
        RECT 454.950 294.600 457.050 295.050 ;
        RECT 421.950 293.400 457.050 294.600 ;
        RECT 421.950 293.100 424.050 293.400 ;
        RECT 454.950 292.950 457.050 293.400 ;
        RECT 478.950 293.100 481.050 295.200 ;
        RECT 505.950 293.400 508.050 295.500 ;
        RECT 541.950 294.600 544.050 295.200 ;
        RECT 565.950 294.600 568.050 295.200 ;
        RECT 574.950 294.600 577.050 295.050 ;
        RECT 580.950 294.600 583.050 295.200 ;
        RECT 541.950 293.400 555.600 294.600 ;
        RECT 479.400 289.050 480.600 293.100 ;
        RECT 394.950 288.600 397.050 288.900 ;
        RECT 323.400 287.400 352.050 288.600 ;
        RECT 368.400 287.400 397.050 288.600 ;
        RECT 310.950 286.950 313.050 287.400 ;
        RECT 319.950 286.800 322.050 287.400 ;
        RECT 337.950 286.800 340.050 287.400 ;
        RECT 349.950 286.500 352.050 287.400 ;
        RECT 394.950 286.800 397.050 287.400 ;
        RECT 475.950 287.400 480.600 289.050 ;
        RECT 487.950 288.600 490.050 288.900 ;
        RECT 506.400 288.600 507.600 293.400 ;
        RECT 541.950 293.100 544.050 293.400 ;
        RECT 554.400 289.050 555.600 293.400 ;
        RECT 565.950 293.400 583.050 294.600 ;
        RECT 565.950 293.100 568.050 293.400 ;
        RECT 574.950 292.950 577.050 293.400 ;
        RECT 580.950 293.100 583.050 293.400 ;
        RECT 589.950 294.600 592.050 295.200 ;
        RECT 607.950 294.600 610.050 295.200 ;
        RECT 631.950 294.750 634.050 295.200 ;
        RECT 640.950 294.750 643.050 295.200 ;
        RECT 589.950 293.400 597.600 294.600 ;
        RECT 589.950 293.100 592.050 293.400 ;
        RECT 487.950 287.400 507.600 288.600 ;
        RECT 475.950 286.950 480.000 287.400 ;
        RECT 487.950 286.800 490.050 287.400 ;
        RECT 553.950 286.950 556.050 289.050 ;
        RECT 559.950 288.450 562.050 288.900 ;
        RECT 568.950 288.450 571.050 288.900 ;
        RECT 559.950 287.250 571.050 288.450 ;
        RECT 596.400 288.600 597.600 293.400 ;
        RECT 607.950 293.400 630.600 294.600 ;
        RECT 607.950 293.100 610.050 293.400 ;
        RECT 629.400 291.600 630.600 293.400 ;
        RECT 631.950 293.550 643.050 294.750 ;
        RECT 631.950 293.100 634.050 293.550 ;
        RECT 640.950 293.100 643.050 293.550 ;
        RECT 670.950 294.600 673.050 295.200 ;
        RECT 685.950 294.600 688.050 295.200 ;
        RECT 670.950 293.400 688.050 294.600 ;
        RECT 670.950 293.100 673.050 293.400 ;
        RECT 685.950 293.100 688.050 293.400 ;
        RECT 691.950 294.750 694.050 295.200 ;
        RECT 700.950 294.750 703.050 295.200 ;
        RECT 691.950 293.550 703.050 294.750 ;
        RECT 691.950 293.100 694.050 293.550 ;
        RECT 700.950 293.100 703.050 293.550 ;
        RECT 715.950 294.600 718.050 295.200 ;
        RECT 739.950 294.600 742.050 295.200 ;
        RECT 757.950 294.600 760.050 295.050 ;
        RECT 715.950 293.400 742.050 294.600 ;
        RECT 715.950 293.100 718.050 293.400 ;
        RECT 739.950 293.100 742.050 293.400 ;
        RECT 746.400 293.400 760.050 294.600 ;
        RECT 629.400 291.000 639.600 291.600 ;
        RECT 629.400 290.400 640.050 291.000 ;
        RECT 604.950 288.600 607.050 288.900 ;
        RECT 596.400 287.400 607.050 288.600 ;
        RECT 559.950 286.800 562.050 287.250 ;
        RECT 568.950 286.800 571.050 287.250 ;
        RECT 604.950 286.800 607.050 287.400 ;
        RECT 637.950 286.950 640.050 290.400 ;
        RECT 646.950 288.450 649.050 288.900 ;
        RECT 655.950 288.450 658.050 288.900 ;
        RECT 646.950 287.250 658.050 288.450 ;
        RECT 646.950 286.800 649.050 287.250 ;
        RECT 655.950 286.800 658.050 287.250 ;
        RECT 679.950 288.450 682.050 288.900 ;
        RECT 688.950 288.450 691.050 288.900 ;
        RECT 679.950 287.250 691.050 288.450 ;
        RECT 679.950 286.800 682.050 287.250 ;
        RECT 688.950 286.800 691.050 287.250 ;
        RECT 706.950 288.450 709.050 288.900 ;
        RECT 712.950 288.600 715.050 288.900 ;
        RECT 736.950 288.600 739.050 288.900 ;
        RECT 712.950 288.450 739.050 288.600 ;
        RECT 706.950 287.400 739.050 288.450 ;
        RECT 706.950 287.250 715.050 287.400 ;
        RECT 706.950 286.800 709.050 287.250 ;
        RECT 712.950 286.800 715.050 287.250 ;
        RECT 736.950 286.800 739.050 287.400 ;
        RECT 742.950 288.600 745.050 288.900 ;
        RECT 746.400 288.600 747.600 293.400 ;
        RECT 757.950 292.950 760.050 293.400 ;
        RECT 805.950 294.600 808.050 295.050 ;
        RECT 814.950 294.600 817.050 295.200 ;
        RECT 877.950 294.600 880.050 295.200 ;
        RECT 805.950 293.400 817.050 294.600 ;
        RECT 805.950 292.950 808.050 293.400 ;
        RECT 814.950 293.100 817.050 293.400 ;
        RECT 863.400 293.400 880.050 294.600 ;
        RECT 742.950 287.400 747.600 288.600 ;
        RECT 754.950 288.450 757.050 288.900 ;
        RECT 763.950 288.450 766.050 288.900 ;
        RECT 742.950 286.800 745.050 287.400 ;
        RECT 754.950 287.250 766.050 288.450 ;
        RECT 754.950 286.800 757.050 287.250 ;
        RECT 763.950 286.800 766.050 287.250 ;
        RECT 787.950 288.450 790.050 288.900 ;
        RECT 817.950 288.450 820.050 288.900 ;
        RECT 787.950 287.250 820.050 288.450 ;
        RECT 787.950 286.800 790.050 287.250 ;
        RECT 817.950 286.800 820.050 287.250 ;
        RECT 823.950 288.600 826.050 289.050 ;
        RECT 863.400 288.900 864.600 293.400 ;
        RECT 877.950 293.100 880.050 293.400 ;
        RECT 838.950 288.600 841.050 288.900 ;
        RECT 823.950 287.400 841.050 288.600 ;
        RECT 823.950 286.950 826.050 287.400 ;
        RECT 838.950 286.800 841.050 287.400 ;
        RECT 862.950 286.800 865.050 288.900 ;
        RECT 289.950 285.600 292.050 286.050 ;
        RECT 301.950 285.600 304.050 286.050 ;
        RECT 289.950 284.400 304.050 285.600 ;
        RECT 289.950 283.950 292.050 284.400 ;
        RECT 301.950 283.950 304.050 284.400 ;
        RECT 361.950 285.600 364.050 286.050 ;
        RECT 379.950 285.600 382.050 286.050 ;
        RECT 361.950 284.400 382.050 285.600 ;
        RECT 361.950 283.950 364.050 284.400 ;
        RECT 379.950 283.950 382.050 284.400 ;
        RECT 466.950 285.600 469.050 286.050 ;
        RECT 523.950 285.600 526.050 286.050 ;
        RECT 466.950 284.400 526.050 285.600 ;
        RECT 466.950 283.950 469.050 284.400 ;
        RECT 523.950 283.950 526.050 284.400 ;
        RECT 583.950 285.600 586.050 286.050 ;
        RECT 616.950 285.600 619.050 286.050 ;
        RECT 583.950 284.400 619.050 285.600 ;
        RECT 583.950 283.950 586.050 284.400 ;
        RECT 616.950 283.950 619.050 284.400 ;
        RECT 661.950 285.600 664.050 286.050 ;
        RECT 685.950 285.600 688.050 286.050 ;
        RECT 661.950 284.400 688.050 285.600 ;
        RECT 661.950 283.950 664.050 284.400 ;
        RECT 685.950 283.950 688.050 284.400 ;
        RECT 790.950 285.600 793.050 286.050 ;
        RECT 799.950 285.600 802.050 286.050 ;
        RECT 790.950 284.400 802.050 285.600 ;
        RECT 790.950 283.950 793.050 284.400 ;
        RECT 799.950 283.950 802.050 284.400 ;
        RECT 163.950 282.600 166.050 283.050 ;
        RECT 184.950 282.600 187.050 283.050 ;
        RECT 220.950 282.600 223.050 283.050 ;
        RECT 163.950 281.400 223.050 282.600 ;
        RECT 163.950 280.950 166.050 281.400 ;
        RECT 184.950 280.950 187.050 281.400 ;
        RECT 220.950 280.950 223.050 281.400 ;
        RECT 244.950 282.600 247.050 283.050 ;
        RECT 259.950 282.600 262.050 283.050 ;
        RECT 244.950 281.400 262.050 282.600 ;
        RECT 244.950 280.950 247.050 281.400 ;
        RECT 259.950 280.950 262.050 281.400 ;
        RECT 460.950 282.600 463.050 283.050 ;
        RECT 472.950 282.600 475.050 283.050 ;
        RECT 481.950 282.600 484.050 283.050 ;
        RECT 460.950 281.400 484.050 282.600 ;
        RECT 460.950 280.950 463.050 281.400 ;
        RECT 472.950 280.950 475.050 281.400 ;
        RECT 481.950 280.950 484.050 281.400 ;
        RECT 505.950 282.600 508.050 283.050 ;
        RECT 511.950 282.600 514.050 283.050 ;
        RECT 505.950 281.400 514.050 282.600 ;
        RECT 505.950 280.950 508.050 281.400 ;
        RECT 511.950 280.950 514.050 281.400 ;
        RECT 655.950 282.600 658.050 283.050 ;
        RECT 700.950 282.600 703.050 283.050 ;
        RECT 655.950 281.400 703.050 282.600 ;
        RECT 655.950 280.950 658.050 281.400 ;
        RECT 700.950 280.950 703.050 281.400 ;
        RECT 709.950 282.600 712.050 283.050 ;
        RECT 718.950 282.600 721.050 283.050 ;
        RECT 709.950 281.400 721.050 282.600 ;
        RECT 709.950 280.950 712.050 281.400 ;
        RECT 718.950 280.950 721.050 281.400 ;
        RECT 793.950 282.600 796.050 283.050 ;
        RECT 838.950 282.600 841.050 283.050 ;
        RECT 793.950 281.400 841.050 282.600 ;
        RECT 793.950 280.950 796.050 281.400 ;
        RECT 838.950 280.950 841.050 281.400 ;
        RECT 877.950 282.600 880.050 283.050 ;
        RECT 884.400 282.600 885.600 298.950 ;
        RECT 889.950 292.950 892.050 295.050 ;
        RECT 890.400 289.050 891.600 292.950 ;
        RECT 889.950 286.950 892.050 289.050 ;
        RECT 877.950 281.400 885.600 282.600 ;
        RECT 877.950 280.950 880.050 281.400 ;
        RECT 142.950 279.600 145.050 280.050 ;
        RECT 148.950 279.600 151.050 280.050 ;
        RECT 142.950 278.400 151.050 279.600 ;
        RECT 142.950 277.950 145.050 278.400 ;
        RECT 148.950 277.950 151.050 278.400 ;
        RECT 229.950 279.600 232.050 280.050 ;
        RECT 283.950 279.600 286.050 280.050 ;
        RECT 343.950 279.600 346.050 280.050 ;
        RECT 385.950 279.600 388.050 280.050 ;
        RECT 229.950 279.000 252.600 279.600 ;
        RECT 229.950 278.400 253.050 279.000 ;
        RECT 229.950 277.950 232.050 278.400 ;
        RECT 139.950 276.600 142.050 277.050 ;
        RECT 151.950 276.600 154.050 277.050 ;
        RECT 139.950 275.400 154.050 276.600 ;
        RECT 139.950 274.950 142.050 275.400 ;
        RECT 151.950 274.950 154.050 275.400 ;
        RECT 169.950 276.600 172.050 277.050 ;
        RECT 226.950 276.600 229.050 277.050 ;
        RECT 169.950 275.400 229.050 276.600 ;
        RECT 169.950 274.950 172.050 275.400 ;
        RECT 226.950 274.950 229.050 275.400 ;
        RECT 250.950 274.950 253.050 278.400 ;
        RECT 283.950 278.400 388.050 279.600 ;
        RECT 283.950 277.950 286.050 278.400 ;
        RECT 343.950 277.950 346.050 278.400 ;
        RECT 385.950 277.950 388.050 278.400 ;
        RECT 514.950 279.600 517.050 280.050 ;
        RECT 544.950 279.600 547.050 280.050 ;
        RECT 514.950 278.400 547.050 279.600 ;
        RECT 514.950 277.950 517.050 278.400 ;
        RECT 544.950 277.950 547.050 278.400 ;
        RECT 643.950 279.600 646.050 280.050 ;
        RECT 664.800 279.600 666.900 280.050 ;
        RECT 643.950 278.400 666.900 279.600 ;
        RECT 643.950 277.950 646.050 278.400 ;
        RECT 664.800 277.950 666.900 278.400 ;
        RECT 667.950 279.600 670.050 280.050 ;
        RECT 703.950 279.600 706.050 280.050 ;
        RECT 667.950 278.400 706.050 279.600 ;
        RECT 667.950 277.950 670.050 278.400 ;
        RECT 703.950 277.950 706.050 278.400 ;
        RECT 769.950 279.600 772.050 280.050 ;
        RECT 799.950 279.600 802.050 280.050 ;
        RECT 859.950 279.600 862.050 280.050 ;
        RECT 769.950 278.400 802.050 279.600 ;
        RECT 769.950 277.950 772.050 278.400 ;
        RECT 799.950 277.950 802.050 278.400 ;
        RECT 845.400 278.400 862.050 279.600 ;
        RECT 845.400 277.050 846.600 278.400 ;
        RECT 859.950 277.950 862.050 278.400 ;
        RECT 274.950 276.600 277.050 277.050 ;
        RECT 280.950 276.600 283.050 277.050 ;
        RECT 274.950 275.400 283.050 276.600 ;
        RECT 274.950 274.950 277.050 275.400 ;
        RECT 280.950 274.950 283.050 275.400 ;
        RECT 574.950 276.600 577.050 277.050 ;
        RECT 616.950 276.600 619.050 277.050 ;
        RECT 574.950 275.400 619.050 276.600 ;
        RECT 574.950 274.950 577.050 275.400 ;
        RECT 616.950 274.950 619.050 275.400 ;
        RECT 640.950 276.600 643.050 277.050 ;
        RECT 667.950 276.600 670.050 276.900 ;
        RECT 676.950 276.600 679.050 277.050 ;
        RECT 745.950 276.600 748.050 277.050 ;
        RECT 640.950 275.400 648.600 276.600 ;
        RECT 640.950 274.950 643.050 275.400 ;
        RECT 170.400 273.600 171.600 274.950 ;
        RECT 143.400 272.400 171.600 273.600 ;
        RECT 232.950 273.600 235.050 274.050 ;
        RECT 271.950 273.600 274.050 274.050 ;
        RECT 232.950 272.400 274.050 273.600 ;
        RECT 61.950 270.600 64.050 271.050 ;
        RECT 100.950 270.600 103.050 271.050 ;
        RECT 143.400 270.600 144.600 272.400 ;
        RECT 232.950 271.950 235.050 272.400 ;
        RECT 271.950 271.950 274.050 272.400 ;
        RECT 427.950 273.600 430.050 274.050 ;
        RECT 481.950 273.600 484.050 274.050 ;
        RECT 427.950 272.400 484.050 273.600 ;
        RECT 427.950 271.950 430.050 272.400 ;
        RECT 481.950 271.950 484.050 272.400 ;
        RECT 598.950 273.600 601.050 274.050 ;
        RECT 647.400 273.600 648.600 275.400 ;
        RECT 667.950 275.400 679.050 276.600 ;
        RECT 667.950 274.800 670.050 275.400 ;
        RECT 676.950 274.950 679.050 275.400 ;
        RECT 680.400 275.400 748.050 276.600 ;
        RECT 680.400 273.600 681.600 275.400 ;
        RECT 745.950 274.950 748.050 275.400 ;
        RECT 811.950 276.600 814.050 277.050 ;
        RECT 844.950 276.600 847.050 277.050 ;
        RECT 811.950 275.400 847.050 276.600 ;
        RECT 811.950 274.950 814.050 275.400 ;
        RECT 844.950 274.950 847.050 275.400 ;
        RECT 598.950 272.400 645.600 273.600 ;
        RECT 647.400 272.400 681.600 273.600 ;
        RECT 697.950 273.600 700.050 274.050 ;
        RECT 760.950 273.600 763.050 274.050 ;
        RECT 697.950 272.400 763.050 273.600 ;
        RECT 598.950 271.950 601.050 272.400 ;
        RECT 61.950 269.400 144.600 270.600 ;
        RECT 199.950 270.600 202.050 271.050 ;
        RECT 238.950 270.600 241.050 271.050 ;
        RECT 418.950 270.600 421.050 271.050 ;
        RECT 199.950 269.400 421.050 270.600 ;
        RECT 61.950 268.950 64.050 269.400 ;
        RECT 100.950 268.950 103.050 269.400 ;
        RECT 199.950 268.950 202.050 269.400 ;
        RECT 238.950 268.950 241.050 269.400 ;
        RECT 418.950 268.950 421.050 269.400 ;
        RECT 478.950 270.600 481.050 271.050 ;
        RECT 511.950 270.600 514.050 271.050 ;
        RECT 478.950 269.400 514.050 270.600 ;
        RECT 478.950 268.950 481.050 269.400 ;
        RECT 511.950 268.950 514.050 269.400 ;
        RECT 556.950 270.600 559.050 271.050 ;
        RECT 580.950 270.600 583.050 271.050 ;
        RECT 556.950 269.400 583.050 270.600 ;
        RECT 556.950 268.950 559.050 269.400 ;
        RECT 580.950 268.950 583.050 269.400 ;
        RECT 619.950 270.600 622.050 271.050 ;
        RECT 631.950 270.600 634.050 271.050 ;
        RECT 619.950 269.400 634.050 270.600 ;
        RECT 644.400 270.600 645.600 272.400 ;
        RECT 697.950 271.950 700.050 272.400 ;
        RECT 760.950 271.950 763.050 272.400 ;
        RECT 775.950 273.600 778.050 274.050 ;
        RECT 808.950 273.600 811.050 274.050 ;
        RECT 775.950 272.400 811.050 273.600 ;
        RECT 775.950 271.950 778.050 272.400 ;
        RECT 808.950 271.950 811.050 272.400 ;
        RECT 817.950 273.600 820.050 274.050 ;
        RECT 832.950 273.600 835.050 274.050 ;
        RECT 817.950 272.400 855.600 273.600 ;
        RECT 817.950 271.950 820.050 272.400 ;
        RECT 832.950 271.950 835.050 272.400 ;
        RECT 854.400 271.050 855.600 272.400 ;
        RECT 712.950 270.600 715.050 271.050 ;
        RECT 644.400 269.400 715.050 270.600 ;
        RECT 619.950 268.950 622.050 269.400 ;
        RECT 631.950 268.950 634.050 269.400 ;
        RECT 712.950 268.950 715.050 269.400 ;
        RECT 796.950 270.600 799.050 271.050 ;
        RECT 826.950 270.600 829.050 271.050 ;
        RECT 796.950 269.400 829.050 270.600 ;
        RECT 854.400 269.400 859.050 271.050 ;
        RECT 796.950 268.950 799.050 269.400 ;
        RECT 826.950 268.950 829.050 269.400 ;
        RECT 855.000 268.950 859.050 269.400 ;
        RECT 880.950 270.600 883.050 271.050 ;
        RECT 895.950 270.600 898.050 271.050 ;
        RECT 880.950 269.400 898.050 270.600 ;
        RECT 880.950 268.950 883.050 269.400 ;
        RECT 895.950 268.950 898.050 269.400 ;
        RECT 148.950 267.600 151.050 268.050 ;
        RECT 196.950 267.600 199.050 268.050 ;
        RECT 148.950 266.400 199.050 267.600 ;
        RECT 148.950 265.950 151.050 266.400 ;
        RECT 196.950 265.950 199.050 266.400 ;
        RECT 256.950 267.600 259.050 268.050 ;
        RECT 295.950 267.600 298.050 268.050 ;
        RECT 256.950 266.400 298.050 267.600 ;
        RECT 256.950 265.950 259.050 266.400 ;
        RECT 295.950 265.950 298.050 266.400 ;
        RECT 304.950 267.600 307.050 268.050 ;
        RECT 319.950 267.600 322.050 268.050 ;
        RECT 349.950 267.600 352.050 268.050 ;
        RECT 415.950 267.600 418.050 268.050 ;
        RECT 304.950 266.400 418.050 267.600 ;
        RECT 304.950 265.950 307.050 266.400 ;
        RECT 319.950 265.950 322.050 266.400 ;
        RECT 349.950 265.950 352.050 266.400 ;
        RECT 415.950 265.950 418.050 266.400 ;
        RECT 454.950 267.600 457.050 268.050 ;
        RECT 547.950 267.600 550.050 268.050 ;
        RECT 454.950 266.400 550.050 267.600 ;
        RECT 454.950 265.950 457.050 266.400 ;
        RECT 547.950 265.950 550.050 266.400 ;
        RECT 553.950 267.600 556.050 268.050 ;
        RECT 592.950 267.600 595.050 268.050 ;
        RECT 655.950 267.600 658.050 268.050 ;
        RECT 553.950 266.400 658.050 267.600 ;
        RECT 553.950 265.950 556.050 266.400 ;
        RECT 592.950 265.950 595.050 266.400 ;
        RECT 655.950 265.950 658.050 266.400 ;
        RECT 727.950 267.600 730.050 268.050 ;
        RECT 733.950 267.600 736.050 268.050 ;
        RECT 727.950 266.400 736.050 267.600 ;
        RECT 727.950 265.950 730.050 266.400 ;
        RECT 733.950 265.950 736.050 266.400 ;
        RECT 742.950 267.600 745.050 268.050 ;
        RECT 751.950 267.600 754.050 268.050 ;
        RECT 742.950 266.400 754.050 267.600 ;
        RECT 742.950 265.950 745.050 266.400 ;
        RECT 751.950 265.950 754.050 266.400 ;
        RECT 763.950 267.600 766.050 268.050 ;
        RECT 769.950 267.600 772.050 268.050 ;
        RECT 763.950 266.400 772.050 267.600 ;
        RECT 763.950 265.950 766.050 266.400 ;
        RECT 769.950 265.950 772.050 266.400 ;
        RECT 790.950 267.600 793.050 268.050 ;
        RECT 799.950 267.600 802.050 268.050 ;
        RECT 829.950 267.600 832.050 268.050 ;
        RECT 790.950 266.400 798.600 267.600 ;
        RECT 790.950 265.950 793.050 266.400 ;
        RECT 418.950 264.600 421.050 265.050 ;
        RECT 448.950 264.600 451.050 265.050 ;
        RECT 418.950 263.400 451.050 264.600 ;
        RECT 418.950 262.950 421.050 263.400 ;
        RECT 448.950 262.950 451.050 263.400 ;
        RECT 490.950 264.600 493.050 265.050 ;
        RECT 496.950 264.600 499.050 265.050 ;
        RECT 490.950 263.400 499.050 264.600 ;
        RECT 490.950 262.950 493.050 263.400 ;
        RECT 496.950 262.950 499.050 263.400 ;
        RECT 610.950 264.600 613.050 265.050 ;
        RECT 622.950 264.600 625.050 265.050 ;
        RECT 610.950 263.400 625.050 264.600 ;
        RECT 610.950 262.950 613.050 263.400 ;
        RECT 622.950 262.950 625.050 263.400 ;
        RECT 772.950 264.600 775.050 265.050 ;
        RECT 781.950 264.600 784.050 265.050 ;
        RECT 772.950 263.400 784.050 264.600 ;
        RECT 772.950 262.950 775.050 263.400 ;
        RECT 781.950 262.950 784.050 263.400 ;
        RECT 787.950 262.950 790.050 265.050 ;
        RECT 55.950 261.600 58.050 262.200 ;
        RECT 50.400 260.400 58.050 261.600 ;
        RECT 50.400 256.050 51.600 260.400 ;
        RECT 55.950 260.100 58.050 260.400 ;
        RECT 73.950 261.750 76.050 262.200 ;
        RECT 85.950 261.750 88.050 262.200 ;
        RECT 73.950 260.550 88.050 261.750 ;
        RECT 73.950 260.100 76.050 260.550 ;
        RECT 85.950 260.100 88.050 260.550 ;
        RECT 109.950 261.750 112.050 262.200 ;
        RECT 121.950 261.750 124.050 262.200 ;
        RECT 109.950 260.550 124.050 261.750 ;
        RECT 109.950 260.100 112.050 260.550 ;
        RECT 121.950 260.100 124.050 260.550 ;
        RECT 127.950 261.750 130.050 262.200 ;
        RECT 136.950 261.750 139.050 262.200 ;
        RECT 127.950 260.550 139.050 261.750 ;
        RECT 141.000 261.600 145.050 262.050 ;
        RECT 127.950 260.100 130.050 260.550 ;
        RECT 136.950 260.100 139.050 260.550 ;
        RECT 140.400 259.950 145.050 261.600 ;
        RECT 157.950 260.400 160.050 262.500 ;
        RECT 190.950 261.600 193.050 262.050 ;
        RECT 205.950 261.600 208.050 262.200 ;
        RECT 190.950 260.400 208.050 261.600 ;
        RECT 140.400 258.600 141.600 259.950 ;
        RECT 131.400 257.400 141.600 258.600 ;
        RECT 49.950 253.950 52.050 256.050 ;
        RECT 131.400 255.900 132.600 257.400 ;
        RECT 112.950 255.450 115.050 255.900 ;
        RECT 118.950 255.450 121.050 255.900 ;
        RECT 112.950 254.250 121.050 255.450 ;
        RECT 112.950 253.800 115.050 254.250 ;
        RECT 118.950 253.800 121.050 254.250 ;
        RECT 130.950 253.800 133.050 255.900 ;
        RECT 136.950 255.600 139.050 256.050 ;
        RECT 151.950 255.600 154.050 255.900 ;
        RECT 158.400 255.600 159.600 260.400 ;
        RECT 190.950 259.950 193.050 260.400 ;
        RECT 205.950 260.100 208.050 260.400 ;
        RECT 211.950 260.100 214.050 262.200 ;
        RECT 193.950 258.600 196.050 259.050 ;
        RECT 212.400 258.600 213.600 260.100 ;
        RECT 220.950 259.950 223.050 262.050 ;
        RECT 262.950 261.600 265.050 262.500 ;
        RECT 260.400 260.400 265.050 261.600 ;
        RECT 301.950 261.750 304.050 262.200 ;
        RECT 307.950 261.750 310.050 262.200 ;
        RECT 301.950 260.550 310.050 261.750 ;
        RECT 193.950 257.400 213.600 258.600 ;
        RECT 193.950 256.950 196.050 257.400 ;
        RECT 136.950 254.400 159.600 255.600 ;
        RECT 175.950 255.150 178.050 255.600 ;
        RECT 190.950 255.150 193.050 255.600 ;
        RECT 136.950 253.950 139.050 254.400 ;
        RECT 151.950 253.800 154.050 254.400 ;
        RECT 175.950 253.950 193.050 255.150 ;
        RECT 175.950 253.500 178.050 253.950 ;
        RECT 190.950 253.500 193.050 253.950 ;
        RECT 196.950 255.450 199.050 255.900 ;
        RECT 202.950 255.450 205.050 255.900 ;
        RECT 196.950 254.250 205.050 255.450 ;
        RECT 196.950 253.800 199.050 254.250 ;
        RECT 202.950 253.800 205.050 254.250 ;
        RECT 208.950 255.450 211.050 255.900 ;
        RECT 217.950 255.450 220.050 255.900 ;
        RECT 208.950 254.250 220.050 255.450 ;
        RECT 221.400 255.600 222.600 259.950 ;
        RECT 241.950 258.600 244.050 259.050 ;
        RECT 260.400 258.600 261.600 260.400 ;
        RECT 301.950 260.100 304.050 260.550 ;
        RECT 307.950 260.100 310.050 260.550 ;
        RECT 325.950 261.600 328.050 262.050 ;
        RECT 331.950 261.600 334.050 262.200 ;
        RECT 325.950 260.400 334.050 261.600 ;
        RECT 391.950 261.600 394.050 262.500 ;
        RECT 406.950 261.750 409.050 262.200 ;
        RECT 415.950 261.750 418.050 262.200 ;
        RECT 406.950 261.600 418.050 261.750 ;
        RECT 391.950 260.550 418.050 261.600 ;
        RECT 391.950 260.400 409.050 260.550 ;
        RECT 325.950 259.950 328.050 260.400 ;
        RECT 331.950 260.100 334.050 260.400 ;
        RECT 406.950 260.100 409.050 260.400 ;
        RECT 415.950 260.100 418.050 260.550 ;
        RECT 430.950 261.750 433.050 262.200 ;
        RECT 439.950 261.750 442.050 262.200 ;
        RECT 430.950 260.550 442.050 261.750 ;
        RECT 430.950 260.100 433.050 260.550 ;
        RECT 439.950 260.100 442.050 260.550 ;
        RECT 451.950 261.600 454.050 262.050 ;
        RECT 451.950 260.400 459.600 261.600 ;
        RECT 451.950 259.950 454.050 260.400 ;
        RECT 458.400 258.600 459.600 260.400 ;
        RECT 475.950 259.950 478.050 262.050 ;
        RECT 499.950 261.750 502.050 262.200 ;
        RECT 505.950 261.750 508.050 262.200 ;
        RECT 499.950 260.550 508.050 261.750 ;
        RECT 499.950 260.100 502.050 260.550 ;
        RECT 505.950 260.100 508.050 260.550 ;
        RECT 520.950 261.600 523.050 262.050 ;
        RECT 532.950 261.600 535.050 262.200 ;
        RECT 520.950 260.400 535.050 261.600 ;
        RECT 520.950 259.950 523.050 260.400 ;
        RECT 532.950 260.100 535.050 260.400 ;
        RECT 556.950 261.600 559.050 262.200 ;
        RECT 565.950 261.600 568.050 262.050 ;
        RECT 601.950 261.600 604.050 262.200 ;
        RECT 670.950 261.600 673.050 262.050 ;
        RECT 679.950 261.600 682.050 262.200 ;
        RECT 556.950 260.400 568.050 261.600 ;
        RECT 556.950 260.100 559.050 260.400 ;
        RECT 565.950 259.950 568.050 260.400 ;
        RECT 584.400 260.400 627.600 261.600 ;
        RECT 241.950 257.400 261.600 258.600 ;
        RECT 365.400 257.400 465.600 258.600 ;
        RECT 241.950 256.950 244.050 257.400 ;
        RECT 223.950 255.600 226.050 255.900 ;
        RECT 221.400 254.400 226.050 255.600 ;
        RECT 208.950 253.800 211.050 254.250 ;
        RECT 217.950 253.800 220.050 254.250 ;
        RECT 223.950 253.800 226.050 254.400 ;
        RECT 280.950 255.150 283.050 255.600 ;
        RECT 295.950 255.150 298.050 255.600 ;
        RECT 280.950 253.950 298.050 255.150 ;
        RECT 280.950 253.500 283.050 253.950 ;
        RECT 295.950 253.500 298.050 253.950 ;
        RECT 313.950 255.450 316.050 255.900 ;
        RECT 319.950 255.450 322.050 255.900 ;
        RECT 365.400 255.600 366.600 257.400 ;
        RECT 409.950 255.600 412.050 255.900 ;
        RECT 427.950 255.600 430.050 255.900 ;
        RECT 313.950 254.250 322.050 255.450 ;
        RECT 313.950 253.800 316.050 254.250 ;
        RECT 319.950 253.800 322.050 254.250 ;
        RECT 364.950 253.500 367.050 255.600 ;
        RECT 409.950 254.400 430.050 255.600 ;
        RECT 409.950 253.800 412.050 254.400 ;
        RECT 427.950 253.800 430.050 254.400 ;
        RECT 433.950 255.450 436.050 255.900 ;
        RECT 442.800 255.450 444.900 255.900 ;
        RECT 451.950 255.600 454.050 256.050 ;
        RECT 464.400 255.600 465.600 257.400 ;
        RECT 476.400 256.050 477.600 259.950 ;
        RECT 433.950 254.250 444.900 255.450 ;
        RECT 446.400 255.000 454.050 255.600 ;
        RECT 433.950 253.800 436.050 254.250 ;
        RECT 442.800 253.800 444.900 254.250 ;
        RECT 445.950 254.400 454.050 255.000 ;
        RECT 43.950 252.600 46.050 253.050 ;
        RECT 58.950 252.600 61.050 253.050 ;
        RECT 43.950 251.400 61.050 252.600 ;
        RECT 43.950 250.950 46.050 251.400 ;
        RECT 58.950 250.950 61.050 251.400 ;
        RECT 445.950 250.950 448.050 254.400 ;
        RECT 451.950 253.950 454.050 254.400 ;
        RECT 463.950 253.500 466.050 255.600 ;
        RECT 475.950 253.950 478.050 256.050 ;
        RECT 584.400 255.900 585.600 260.400 ;
        RECT 601.950 260.100 604.050 260.400 ;
        RECT 626.400 255.900 627.600 260.400 ;
        RECT 670.950 260.400 682.050 261.600 ;
        RECT 670.950 259.950 673.050 260.400 ;
        RECT 679.950 260.100 682.050 260.400 ;
        RECT 703.950 261.600 706.050 262.200 ;
        RECT 721.950 261.600 724.050 262.200 ;
        RECT 703.950 260.400 724.050 261.600 ;
        RECT 703.950 260.100 706.050 260.400 ;
        RECT 721.950 260.100 724.050 260.400 ;
        RECT 727.950 261.600 730.050 262.200 ;
        RECT 736.950 261.600 739.050 262.050 ;
        RECT 727.950 260.400 739.050 261.600 ;
        RECT 727.950 260.100 730.050 260.400 ;
        RECT 736.950 259.950 739.050 260.400 ;
        RECT 742.950 258.600 745.050 262.050 ;
        RECT 751.950 260.100 754.050 262.200 ;
        RECT 752.400 258.600 753.600 260.100 ;
        RECT 778.950 259.950 781.050 262.050 ;
        RECT 742.950 258.000 750.600 258.600 ;
        RECT 743.400 257.400 750.600 258.000 ;
        RECT 752.400 258.000 759.600 258.600 ;
        RECT 752.400 257.400 760.050 258.000 ;
        RECT 514.950 255.450 517.050 255.900 ;
        RECT 520.950 255.450 523.050 255.900 ;
        RECT 514.950 254.250 523.050 255.450 ;
        RECT 514.950 253.800 517.050 254.250 ;
        RECT 520.950 253.800 523.050 254.250 ;
        RECT 583.950 253.800 586.050 255.900 ;
        RECT 592.950 255.450 595.050 255.900 ;
        RECT 598.950 255.450 601.050 255.900 ;
        RECT 592.950 254.250 601.050 255.450 ;
        RECT 592.950 253.800 595.050 254.250 ;
        RECT 598.950 253.800 601.050 254.250 ;
        RECT 625.950 253.800 628.050 255.900 ;
        RECT 637.950 255.600 640.050 256.050 ;
        RECT 673.950 255.600 676.050 256.050 ;
        RECT 637.950 254.400 676.050 255.600 ;
        RECT 637.950 253.950 640.050 254.400 ;
        RECT 673.950 253.950 676.050 254.400 ;
        RECT 682.950 255.450 685.050 255.900 ;
        RECT 688.950 255.450 691.050 255.900 ;
        RECT 682.950 254.250 691.050 255.450 ;
        RECT 682.950 253.800 685.050 254.250 ;
        RECT 688.950 253.800 691.050 254.250 ;
        RECT 706.950 255.600 709.050 255.900 ;
        RECT 718.950 255.600 721.050 255.900 ;
        RECT 706.950 255.450 721.050 255.600 ;
        RECT 733.950 255.450 736.050 255.900 ;
        RECT 706.950 254.400 736.050 255.450 ;
        RECT 749.400 255.600 750.600 257.400 ;
        RECT 749.400 255.000 753.600 255.600 ;
        RECT 749.400 254.400 754.050 255.000 ;
        RECT 706.950 253.800 709.050 254.400 ;
        RECT 718.950 254.250 736.050 254.400 ;
        RECT 718.950 253.800 721.050 254.250 ;
        RECT 733.950 253.800 736.050 254.250 ;
        RECT 508.950 252.600 511.050 253.050 ;
        RECT 535.950 252.600 538.050 253.050 ;
        RECT 508.950 251.400 538.050 252.600 ;
        RECT 508.950 250.950 511.050 251.400 ;
        RECT 535.950 250.950 538.050 251.400 ;
        RECT 676.950 252.600 679.050 253.050 ;
        RECT 691.950 252.600 694.050 253.050 ;
        RECT 676.950 251.400 694.050 252.600 ;
        RECT 676.950 250.950 679.050 251.400 ;
        RECT 691.950 250.950 694.050 251.400 ;
        RECT 751.950 250.950 754.050 254.400 ;
        RECT 757.950 253.950 760.050 257.400 ;
        RECT 779.400 256.050 780.600 259.950 ;
        RECT 763.950 255.450 766.050 255.900 ;
        RECT 769.950 255.450 772.050 255.900 ;
        RECT 763.950 254.250 772.050 255.450 ;
        RECT 763.950 253.800 766.050 254.250 ;
        RECT 769.950 253.800 772.050 254.250 ;
        RECT 778.950 253.950 781.050 256.050 ;
        RECT 788.400 255.900 789.600 262.950 ;
        RECT 787.950 253.800 790.050 255.900 ;
        RECT 797.400 253.050 798.600 266.400 ;
        RECT 799.950 266.400 832.050 267.600 ;
        RECT 799.950 265.950 802.050 266.400 ;
        RECT 829.950 265.950 832.050 266.400 ;
        RECT 862.950 267.600 865.050 268.050 ;
        RECT 883.950 267.600 886.050 268.050 ;
        RECT 862.950 266.400 886.050 267.600 ;
        RECT 862.950 265.950 865.050 266.400 ;
        RECT 883.950 265.950 886.050 266.400 ;
        RECT 811.950 261.600 814.050 265.050 ;
        RECT 820.950 262.950 823.050 265.050 ;
        RECT 817.950 261.600 820.050 262.200 ;
        RECT 811.950 261.000 820.050 261.600 ;
        RECT 812.400 260.400 820.050 261.000 ;
        RECT 817.950 260.100 820.050 260.400 ;
        RECT 821.400 258.600 822.600 262.950 ;
        RECT 826.950 259.950 829.050 262.050 ;
        RECT 844.950 261.600 847.050 262.200 ;
        RECT 859.950 261.600 862.050 262.050 ;
        RECT 833.400 260.400 847.050 261.600 ;
        RECT 815.400 257.400 822.600 258.600 ;
        RECT 805.950 255.600 808.050 256.050 ;
        RECT 811.950 255.600 814.050 256.050 ;
        RECT 805.950 254.400 814.050 255.600 ;
        RECT 805.950 253.950 808.050 254.400 ;
        RECT 811.950 253.950 814.050 254.400 ;
        RECT 815.400 253.050 816.600 257.400 ;
        RECT 827.400 256.050 828.600 259.950 ;
        RECT 833.400 256.050 834.600 260.400 ;
        RECT 844.950 260.100 847.050 260.400 ;
        RECT 848.400 260.400 862.050 261.600 ;
        RECT 848.400 256.050 849.600 260.400 ;
        RECT 859.950 259.950 862.050 260.400 ;
        RECT 868.950 261.600 871.050 262.200 ;
        RECT 895.950 261.600 898.050 262.050 ;
        RECT 868.950 260.400 898.050 261.600 ;
        RECT 868.950 260.100 871.050 260.400 ;
        RECT 895.950 259.950 898.050 260.400 ;
        RECT 856.950 256.950 859.050 259.050 ;
        RECT 826.950 253.950 829.050 256.050 ;
        RECT 832.950 253.950 835.050 256.050 ;
        RECT 847.950 253.950 850.050 256.050 ;
        RECT 79.950 249.600 82.050 250.050 ;
        RECT 145.950 249.600 148.050 250.050 ;
        RECT 193.950 249.600 196.050 250.050 ;
        RECT 199.950 249.600 202.050 250.050 ;
        RECT 79.950 248.400 202.050 249.600 ;
        RECT 79.950 247.950 82.050 248.400 ;
        RECT 145.950 247.950 148.050 248.400 ;
        RECT 193.950 247.950 196.050 248.400 ;
        RECT 199.950 247.950 202.050 248.400 ;
        RECT 205.950 249.600 208.050 250.050 ;
        RECT 229.950 249.600 232.050 250.050 ;
        RECT 253.950 249.600 256.050 250.050 ;
        RECT 205.950 248.400 256.050 249.600 ;
        RECT 205.950 247.950 208.050 248.400 ;
        RECT 229.950 247.950 232.050 248.400 ;
        RECT 253.950 247.950 256.050 248.400 ;
        RECT 373.950 249.600 376.050 250.050 ;
        RECT 439.950 249.600 442.050 250.050 ;
        RECT 373.950 248.400 442.050 249.600 ;
        RECT 373.950 247.950 376.050 248.400 ;
        RECT 439.950 247.950 442.050 248.400 ;
        RECT 448.950 249.600 451.050 250.050 ;
        RECT 463.950 249.600 466.050 250.050 ;
        RECT 448.950 248.400 466.050 249.600 ;
        RECT 448.950 247.950 451.050 248.400 ;
        RECT 463.950 247.950 466.050 248.400 ;
        RECT 472.950 249.600 475.050 250.050 ;
        RECT 478.950 249.600 481.050 250.050 ;
        RECT 472.950 248.400 481.050 249.600 ;
        RECT 472.950 247.950 475.050 248.400 ;
        RECT 478.950 247.950 481.050 248.400 ;
        RECT 529.950 249.600 532.050 250.050 ;
        RECT 553.950 249.600 556.050 250.050 ;
        RECT 529.950 248.400 556.050 249.600 ;
        RECT 529.950 247.950 532.050 248.400 ;
        RECT 553.950 247.950 556.050 248.400 ;
        RECT 619.950 249.600 622.050 250.050 ;
        RECT 637.950 249.600 640.050 250.050 ;
        RECT 619.950 248.400 640.050 249.600 ;
        RECT 692.400 249.600 693.600 250.950 ;
        RECT 775.950 249.600 778.050 253.050 ;
        RECT 796.950 250.950 799.050 253.050 ;
        RECT 814.950 250.950 817.050 253.050 ;
        RECT 857.400 252.600 858.600 256.950 ;
        RECT 871.950 255.450 874.050 255.900 ;
        RECT 889.950 255.450 892.050 255.900 ;
        RECT 871.950 254.250 892.050 255.450 ;
        RECT 871.950 253.800 874.050 254.250 ;
        RECT 889.950 253.800 892.050 254.250 ;
        RECT 868.950 252.600 871.050 253.050 ;
        RECT 857.400 251.400 871.050 252.600 ;
        RECT 868.950 250.950 871.050 251.400 ;
        RECT 793.950 249.600 796.050 249.900 ;
        RECT 692.400 248.400 796.050 249.600 ;
        RECT 619.950 247.950 622.050 248.400 ;
        RECT 637.950 247.950 640.050 248.400 ;
        RECT 496.950 246.600 499.050 247.050 ;
        RECT 530.400 246.600 531.600 247.950 ;
        RECT 793.950 247.800 796.050 248.400 ;
        RECT 835.950 249.600 838.050 250.050 ;
        RECT 847.950 249.600 850.050 250.050 ;
        RECT 835.950 248.400 850.050 249.600 ;
        RECT 835.950 247.950 838.050 248.400 ;
        RECT 847.950 247.950 850.050 248.400 ;
        RECT 862.950 249.600 865.050 250.050 ;
        RECT 880.950 249.600 883.050 250.050 ;
        RECT 862.950 248.400 883.050 249.600 ;
        RECT 862.950 247.950 865.050 248.400 ;
        RECT 880.950 247.950 883.050 248.400 ;
        RECT 496.950 245.400 531.600 246.600 ;
        RECT 604.950 246.600 607.050 247.050 ;
        RECT 631.950 246.600 634.050 247.050 ;
        RECT 604.950 245.400 634.050 246.600 ;
        RECT 496.950 244.950 499.050 245.400 ;
        RECT 604.950 244.950 607.050 245.400 ;
        RECT 631.950 244.950 634.050 245.400 ;
        RECT 103.950 243.600 106.050 244.050 ;
        RECT 139.950 243.600 142.050 244.050 ;
        RECT 190.950 243.600 193.050 244.050 ;
        RECT 241.950 243.600 244.050 244.050 ;
        RECT 103.950 242.400 244.050 243.600 ;
        RECT 103.950 241.950 106.050 242.400 ;
        RECT 139.950 241.950 142.050 242.400 ;
        RECT 190.950 241.950 193.050 242.400 ;
        RECT 241.950 241.950 244.050 242.400 ;
        RECT 271.950 243.600 274.050 244.050 ;
        RECT 433.950 243.600 436.050 244.050 ;
        RECT 271.950 242.400 436.050 243.600 ;
        RECT 271.950 241.950 274.050 242.400 ;
        RECT 433.950 241.950 436.050 242.400 ;
        RECT 841.950 243.600 844.050 244.050 ;
        RECT 889.950 243.600 892.050 244.050 ;
        RECT 841.950 242.400 892.050 243.600 ;
        RECT 841.950 241.950 844.050 242.400 ;
        RECT 889.950 241.950 892.050 242.400 ;
        RECT 244.950 240.600 247.050 241.050 ;
        RECT 256.950 240.600 259.050 241.050 ;
        RECT 244.950 239.400 259.050 240.600 ;
        RECT 244.950 238.950 247.050 239.400 ;
        RECT 256.950 238.950 259.050 239.400 ;
        RECT 367.950 240.600 370.050 241.050 ;
        RECT 379.950 240.600 382.050 241.050 ;
        RECT 367.950 239.400 382.050 240.600 ;
        RECT 367.950 238.950 370.050 239.400 ;
        RECT 379.950 238.950 382.050 239.400 ;
        RECT 400.950 240.600 403.050 241.050 ;
        RECT 445.950 240.600 448.050 241.050 ;
        RECT 400.950 239.400 448.050 240.600 ;
        RECT 400.950 238.950 403.050 239.400 ;
        RECT 445.950 238.950 448.050 239.400 ;
        RECT 466.950 240.600 469.050 241.050 ;
        RECT 475.950 240.600 478.050 241.050 ;
        RECT 466.950 239.400 478.050 240.600 ;
        RECT 466.950 238.950 469.050 239.400 ;
        RECT 475.950 238.950 478.050 239.400 ;
        RECT 517.950 240.600 520.050 241.050 ;
        RECT 559.950 240.600 562.050 241.050 ;
        RECT 595.950 240.600 598.050 241.050 ;
        RECT 517.950 239.400 598.050 240.600 ;
        RECT 517.950 238.950 520.050 239.400 ;
        RECT 559.950 238.950 562.050 239.400 ;
        RECT 595.950 238.950 598.050 239.400 ;
        RECT 670.950 240.600 673.050 241.050 ;
        RECT 721.950 240.600 724.050 241.050 ;
        RECT 670.950 239.400 724.050 240.600 ;
        RECT 670.950 238.950 673.050 239.400 ;
        RECT 721.950 238.950 724.050 239.400 ;
        RECT 796.950 240.600 799.050 241.050 ;
        RECT 811.950 240.600 814.050 241.050 ;
        RECT 796.950 239.400 814.050 240.600 ;
        RECT 796.950 238.950 799.050 239.400 ;
        RECT 811.950 238.950 814.050 239.400 ;
        RECT 820.950 240.600 823.050 241.050 ;
        RECT 883.950 240.600 886.050 241.050 ;
        RECT 820.950 239.400 886.050 240.600 ;
        RECT 820.950 238.950 823.050 239.400 ;
        RECT 883.950 238.950 886.050 239.400 ;
        RECT 52.950 237.600 55.050 238.050 ;
        RECT 64.950 237.600 67.050 238.050 ;
        RECT 205.950 237.600 208.050 238.050 ;
        RECT 52.950 236.400 208.050 237.600 ;
        RECT 52.950 235.950 55.050 236.400 ;
        RECT 64.950 235.950 67.050 236.400 ;
        RECT 205.950 235.950 208.050 236.400 ;
        RECT 268.950 237.600 271.050 238.050 ;
        RECT 355.950 237.600 358.050 238.050 ;
        RECT 268.950 236.400 358.050 237.600 ;
        RECT 446.400 237.600 447.600 238.950 ;
        RECT 499.950 237.600 502.050 238.050 ;
        RECT 446.400 236.400 502.050 237.600 ;
        RECT 268.950 235.950 271.050 236.400 ;
        RECT 355.950 235.950 358.050 236.400 ;
        RECT 499.950 235.950 502.050 236.400 ;
        RECT 739.950 237.600 742.050 238.050 ;
        RECT 766.950 237.600 769.050 238.050 ;
        RECT 739.950 236.400 769.050 237.600 ;
        RECT 739.950 235.950 742.050 236.400 ;
        RECT 766.950 235.950 769.050 236.400 ;
        RECT 793.950 237.600 796.050 238.050 ;
        RECT 805.950 237.600 808.050 238.050 ;
        RECT 793.950 236.400 808.050 237.600 ;
        RECT 793.950 235.950 796.050 236.400 ;
        RECT 805.950 235.950 808.050 236.400 ;
        RECT 838.950 237.600 841.050 238.050 ;
        RECT 853.950 237.600 856.050 238.050 ;
        RECT 838.950 236.400 856.050 237.600 ;
        RECT 838.950 235.950 841.050 236.400 ;
        RECT 853.950 235.950 856.050 236.400 ;
        RECT 433.950 234.600 436.050 235.050 ;
        RECT 508.950 234.600 511.050 235.050 ;
        RECT 433.950 233.400 511.050 234.600 ;
        RECT 433.950 232.950 436.050 233.400 ;
        RECT 508.950 232.950 511.050 233.400 ;
        RECT 664.950 234.600 667.050 235.050 ;
        RECT 688.950 234.600 691.050 235.050 ;
        RECT 664.950 233.400 691.050 234.600 ;
        RECT 664.950 232.950 667.050 233.400 ;
        RECT 688.950 232.950 691.050 233.400 ;
        RECT 718.950 234.600 721.050 235.050 ;
        RECT 748.950 234.600 751.050 235.050 ;
        RECT 820.950 234.600 823.050 235.050 ;
        RECT 718.950 233.400 823.050 234.600 ;
        RECT 718.950 232.950 721.050 233.400 ;
        RECT 748.950 232.950 751.050 233.400 ;
        RECT 820.950 232.950 823.050 233.400 ;
        RECT 22.950 231.600 25.050 232.050 ;
        RECT 79.950 231.600 82.050 232.050 ;
        RECT 22.950 230.400 82.050 231.600 ;
        RECT 22.950 229.950 25.050 230.400 ;
        RECT 79.950 229.950 82.050 230.400 ;
        RECT 454.950 231.600 457.050 232.050 ;
        RECT 469.950 231.600 472.050 232.050 ;
        RECT 454.950 230.400 472.050 231.600 ;
        RECT 454.950 229.950 457.050 230.400 ;
        RECT 469.950 229.950 472.050 230.400 ;
        RECT 652.950 231.600 655.050 232.050 ;
        RECT 691.950 231.600 694.050 232.050 ;
        RECT 652.950 230.400 694.050 231.600 ;
        RECT 652.950 229.950 655.050 230.400 ;
        RECT 691.950 229.950 694.050 230.400 ;
        RECT 754.950 231.600 757.050 232.050 ;
        RECT 796.950 231.600 799.050 232.050 ;
        RECT 832.950 231.600 835.050 232.050 ;
        RECT 754.950 230.400 835.050 231.600 ;
        RECT 754.950 229.950 757.050 230.400 ;
        RECT 796.950 229.950 799.050 230.400 ;
        RECT 832.950 229.950 835.050 230.400 ;
        RECT 865.950 231.600 868.050 232.050 ;
        RECT 880.950 231.600 883.050 232.050 ;
        RECT 865.950 230.400 883.050 231.600 ;
        RECT 865.950 229.950 868.050 230.400 ;
        RECT 880.950 229.950 883.050 230.400 ;
        RECT 13.950 228.600 16.050 229.050 ;
        RECT 127.950 228.600 130.050 229.050 ;
        RECT 166.950 228.600 169.050 229.050 ;
        RECT 187.950 228.600 190.050 229.050 ;
        RECT 250.950 228.600 253.050 229.050 ;
        RECT 274.950 228.600 277.050 229.050 ;
        RECT 292.950 228.600 295.050 229.050 ;
        RECT 13.950 227.400 295.050 228.600 ;
        RECT 13.950 226.950 16.050 227.400 ;
        RECT 127.950 226.950 130.050 227.400 ;
        RECT 166.950 226.950 169.050 227.400 ;
        RECT 187.950 226.950 190.050 227.400 ;
        RECT 250.950 226.950 253.050 227.400 ;
        RECT 274.950 226.950 277.050 227.400 ;
        RECT 292.950 226.950 295.050 227.400 ;
        RECT 547.950 228.600 550.050 229.050 ;
        RECT 583.950 228.600 586.050 229.050 ;
        RECT 547.950 227.400 586.050 228.600 ;
        RECT 547.950 226.950 550.050 227.400 ;
        RECT 583.950 226.950 586.050 227.400 ;
        RECT 736.950 228.600 739.050 229.050 ;
        RECT 748.950 228.600 751.050 229.050 ;
        RECT 736.950 227.400 751.050 228.600 ;
        RECT 736.950 226.950 739.050 227.400 ;
        RECT 748.950 226.950 751.050 227.400 ;
        RECT 805.950 228.600 808.050 229.050 ;
        RECT 838.950 228.600 841.050 229.050 ;
        RECT 805.950 227.400 841.050 228.600 ;
        RECT 805.950 226.950 808.050 227.400 ;
        RECT 838.950 226.950 841.050 227.400 ;
        RECT 232.950 225.600 235.050 226.050 ;
        RECT 238.950 225.600 241.050 226.050 ;
        RECT 232.950 224.400 241.050 225.600 ;
        RECT 232.950 223.950 235.050 224.400 ;
        RECT 238.950 223.950 241.050 224.400 ;
        RECT 442.950 225.600 445.050 226.050 ;
        RECT 487.950 225.600 490.050 226.050 ;
        RECT 442.950 224.400 490.050 225.600 ;
        RECT 442.950 223.950 445.050 224.400 ;
        RECT 487.950 223.950 490.050 224.400 ;
        RECT 574.950 225.600 577.050 226.050 ;
        RECT 622.950 225.600 625.050 226.050 ;
        RECT 646.950 225.600 649.050 226.050 ;
        RECT 574.950 224.400 649.050 225.600 ;
        RECT 574.950 223.950 577.050 224.400 ;
        RECT 622.950 223.950 625.050 224.400 ;
        RECT 646.950 223.950 649.050 224.400 ;
        RECT 766.950 225.600 769.050 226.050 ;
        RECT 787.800 225.600 789.900 226.050 ;
        RECT 766.950 224.400 789.900 225.600 ;
        RECT 766.950 223.950 769.050 224.400 ;
        RECT 787.800 223.950 789.900 224.400 ;
        RECT 790.950 225.600 793.050 226.050 ;
        RECT 802.950 225.600 805.050 226.050 ;
        RECT 790.950 224.400 805.050 225.600 ;
        RECT 790.950 223.950 793.050 224.400 ;
        RECT 802.950 223.950 805.050 224.400 ;
        RECT 874.950 225.600 877.050 226.050 ;
        RECT 886.950 225.600 889.050 226.050 ;
        RECT 874.950 224.400 889.050 225.600 ;
        RECT 874.950 223.950 877.050 224.400 ;
        RECT 886.950 223.950 889.050 224.400 ;
        RECT 4.950 222.600 7.050 223.050 ;
        RECT 13.950 222.600 16.050 223.050 ;
        RECT 4.950 221.400 16.050 222.600 ;
        RECT 4.950 220.950 7.050 221.400 ;
        RECT 13.950 220.950 16.050 221.400 ;
        RECT 67.950 222.600 70.050 223.050 ;
        RECT 91.950 222.600 94.050 223.050 ;
        RECT 67.950 221.400 94.050 222.600 ;
        RECT 67.950 220.950 70.050 221.400 ;
        RECT 91.950 220.950 94.050 221.400 ;
        RECT 124.950 222.600 127.050 223.050 ;
        RECT 157.950 222.600 160.050 223.050 ;
        RECT 124.950 221.400 160.050 222.600 ;
        RECT 124.950 220.950 127.050 221.400 ;
        RECT 157.950 220.950 160.050 221.400 ;
        RECT 241.950 222.600 244.050 223.050 ;
        RECT 277.950 222.600 280.050 223.050 ;
        RECT 241.950 221.400 280.050 222.600 ;
        RECT 241.950 220.950 244.050 221.400 ;
        RECT 277.950 220.950 280.050 221.400 ;
        RECT 481.950 222.600 484.050 223.050 ;
        RECT 517.950 222.600 520.050 223.050 ;
        RECT 481.950 221.400 520.050 222.600 ;
        RECT 481.950 220.950 484.050 221.400 ;
        RECT 517.950 220.950 520.050 221.400 ;
        RECT 550.950 222.600 553.050 223.050 ;
        RECT 571.950 222.600 574.050 223.050 ;
        RECT 550.950 221.400 574.050 222.600 ;
        RECT 550.950 220.950 553.050 221.400 ;
        RECT 571.950 220.950 574.050 221.400 ;
        RECT 769.950 222.600 772.050 223.050 ;
        RECT 799.950 222.600 802.050 223.050 ;
        RECT 769.950 221.400 802.050 222.600 ;
        RECT 769.950 220.950 772.050 221.400 ;
        RECT 799.950 220.950 802.050 221.400 ;
        RECT 850.950 222.600 853.050 223.050 ;
        RECT 862.950 222.600 865.050 223.050 ;
        RECT 850.950 221.400 865.050 222.600 ;
        RECT 850.950 220.950 853.050 221.400 ;
        RECT 862.950 220.950 865.050 221.400 ;
        RECT 49.950 219.600 52.050 220.050 ;
        RECT 55.950 219.600 58.050 220.050 ;
        RECT 49.950 218.400 58.050 219.600 ;
        RECT 49.950 217.950 52.050 218.400 ;
        RECT 55.950 217.950 58.050 218.400 ;
        RECT 97.950 219.600 100.050 220.050 ;
        RECT 124.950 219.600 127.050 219.900 ;
        RECT 97.950 218.400 127.050 219.600 ;
        RECT 97.950 217.950 100.050 218.400 ;
        RECT 124.950 217.800 127.050 218.400 ;
        RECT 316.950 219.600 319.050 220.050 ;
        RECT 328.950 219.600 331.050 220.050 ;
        RECT 334.950 219.600 337.050 220.050 ;
        RECT 316.950 218.400 337.050 219.600 ;
        RECT 316.950 217.950 319.050 218.400 ;
        RECT 328.950 217.950 331.050 218.400 ;
        RECT 334.950 217.950 337.050 218.400 ;
        RECT 433.950 219.600 436.050 220.050 ;
        RECT 448.950 219.600 451.050 220.050 ;
        RECT 511.950 219.600 514.050 220.050 ;
        RECT 559.950 219.600 562.050 220.050 ;
        RECT 766.950 219.600 769.050 220.050 ;
        RECT 433.950 218.400 562.050 219.600 ;
        RECT 433.950 217.950 436.050 218.400 ;
        RECT 448.950 217.950 451.050 218.400 ;
        RECT 511.950 217.950 514.050 218.400 ;
        RECT 559.950 217.950 562.050 218.400 ;
        RECT 758.400 218.400 769.050 219.600 ;
        RECT 13.950 215.400 16.050 217.500 ;
        RECT 73.950 216.750 76.050 217.200 ;
        RECT 79.800 216.750 81.900 217.200 ;
        RECT 73.950 215.550 81.900 216.750 ;
        RECT 14.400 211.050 15.600 215.400 ;
        RECT 73.950 215.100 76.050 215.550 ;
        RECT 79.800 215.100 81.900 215.550 ;
        RECT 82.950 216.600 85.050 217.050 ;
        RECT 115.950 216.600 118.050 217.200 ;
        RECT 82.950 215.400 118.050 216.600 ;
        RECT 82.950 214.950 85.050 215.400 ;
        RECT 115.950 215.100 118.050 215.400 ;
        RECT 130.950 216.600 133.050 217.050 ;
        RECT 139.950 216.600 142.050 217.200 ;
        RECT 130.950 215.400 142.050 216.600 ;
        RECT 130.950 214.950 133.050 215.400 ;
        RECT 139.950 215.100 142.050 215.400 ;
        RECT 163.950 216.750 166.050 217.200 ;
        RECT 169.950 216.750 172.050 217.200 ;
        RECT 163.950 215.550 172.050 216.750 ;
        RECT 181.950 216.600 184.050 217.200 ;
        RECT 163.950 215.100 166.050 215.550 ;
        RECT 169.950 215.100 172.050 215.550 ;
        RECT 173.400 215.400 184.050 216.600 ;
        RECT 173.400 213.600 174.600 215.400 ;
        RECT 181.950 215.100 184.050 215.400 ;
        RECT 211.950 216.600 214.050 217.200 ;
        RECT 229.950 216.600 232.050 217.050 ;
        RECT 262.950 216.600 265.050 217.200 ;
        RECT 211.950 215.400 265.050 216.600 ;
        RECT 211.950 215.100 214.050 215.400 ;
        RECT 229.950 214.950 232.050 215.400 ;
        RECT 262.950 215.100 265.050 215.400 ;
        RECT 268.950 216.600 271.050 217.200 ;
        RECT 274.950 216.600 277.050 217.050 ;
        RECT 268.950 215.400 277.050 216.600 ;
        RECT 268.950 215.100 271.050 215.400 ;
        RECT 274.950 214.950 277.050 215.400 ;
        RECT 280.950 216.750 283.050 217.200 ;
        RECT 286.950 216.750 289.050 217.200 ;
        RECT 280.950 215.550 289.050 216.750 ;
        RECT 280.950 215.100 283.050 215.550 ;
        RECT 286.950 215.100 289.050 215.550 ;
        RECT 292.950 216.750 295.050 217.200 ;
        RECT 301.800 216.750 303.900 217.200 ;
        RECT 292.950 215.550 303.900 216.750 ;
        RECT 292.950 215.100 295.050 215.550 ;
        RECT 301.800 215.100 303.900 215.550 ;
        RECT 304.950 216.750 307.050 217.200 ;
        RECT 310.950 216.750 313.050 217.200 ;
        RECT 304.950 215.550 313.050 216.750 ;
        RECT 337.950 216.600 340.050 217.200 ;
        RECT 304.950 215.100 307.050 215.550 ;
        RECT 310.950 215.100 313.050 215.550 ;
        RECT 314.400 215.400 340.050 216.600 ;
        RECT 190.950 213.600 193.050 214.050 ;
        RECT 314.400 213.600 315.600 215.400 ;
        RECT 337.950 215.100 340.050 215.400 ;
        RECT 349.950 216.600 352.050 217.050 ;
        RECT 355.950 216.600 358.050 217.200 ;
        RECT 349.950 215.400 358.050 216.600 ;
        RECT 349.950 214.950 352.050 215.400 ;
        RECT 355.950 215.100 358.050 215.400 ;
        RECT 364.950 216.600 367.050 217.050 ;
        RECT 373.950 216.600 376.050 217.200 ;
        RECT 364.950 215.400 376.050 216.600 ;
        RECT 364.950 214.950 367.050 215.400 ;
        RECT 373.950 215.100 376.050 215.400 ;
        RECT 382.950 216.600 385.050 217.200 ;
        RECT 397.950 216.600 400.050 217.200 ;
        RECT 382.950 215.400 400.050 216.600 ;
        RECT 382.950 215.100 385.050 215.400 ;
        RECT 397.950 215.100 400.050 215.400 ;
        RECT 406.950 216.600 409.050 217.200 ;
        RECT 418.950 216.600 421.050 217.050 ;
        RECT 406.950 215.400 421.050 216.600 ;
        RECT 406.950 215.100 409.050 215.400 ;
        RECT 418.950 214.950 421.050 215.400 ;
        RECT 424.950 215.100 427.050 217.200 ;
        RECT 478.950 216.600 481.050 217.200 ;
        RECT 496.950 216.600 499.050 217.200 ;
        RECT 478.950 215.400 499.050 216.600 ;
        RECT 478.950 215.100 481.050 215.400 ;
        RECT 496.950 215.100 499.050 215.400 ;
        RECT 568.950 216.600 571.050 217.050 ;
        RECT 577.950 216.600 580.050 217.200 ;
        RECT 568.950 215.400 580.050 216.600 ;
        RECT 167.400 212.400 174.600 213.600 ;
        RECT 179.400 212.400 193.050 213.600 ;
        RECT 14.400 209.400 19.050 211.050 ;
        RECT 167.400 210.900 168.600 212.400 ;
        RECT 179.400 210.900 180.600 212.400 ;
        RECT 190.950 211.950 193.050 212.400 ;
        RECT 299.400 212.400 315.600 213.600 ;
        RECT 15.000 208.950 19.050 209.400 ;
        RECT 31.950 210.150 34.050 210.600 ;
        RECT 43.950 210.150 46.050 210.600 ;
        RECT 31.950 208.950 46.050 210.150 ;
        RECT 31.950 208.500 34.050 208.950 ;
        RECT 43.950 208.500 46.050 208.950 ;
        RECT 58.950 210.450 61.050 210.900 ;
        RECT 82.950 210.450 85.050 210.900 ;
        RECT 58.950 209.250 85.050 210.450 ;
        RECT 58.950 208.800 61.050 209.250 ;
        RECT 82.950 208.800 85.050 209.250 ;
        RECT 106.950 210.450 109.050 210.900 ;
        RECT 112.950 210.450 115.050 210.900 ;
        RECT 106.950 209.250 115.050 210.450 ;
        RECT 106.950 208.800 109.050 209.250 ;
        RECT 112.950 208.800 115.050 209.250 ;
        RECT 118.950 210.450 121.050 210.900 ;
        RECT 154.950 210.450 157.050 210.900 ;
        RECT 118.950 209.250 157.050 210.450 ;
        RECT 118.950 208.800 121.050 209.250 ;
        RECT 154.950 208.800 157.050 209.250 ;
        RECT 166.950 208.800 169.050 210.900 ;
        RECT 178.950 208.800 181.050 210.900 ;
        RECT 265.950 210.600 268.050 210.900 ;
        RECT 280.950 210.600 283.050 211.050 ;
        RECT 220.950 210.150 223.050 210.600 ;
        RECT 229.950 210.150 232.050 210.600 ;
        RECT 220.950 208.950 232.050 210.150 ;
        RECT 220.950 208.500 223.050 208.950 ;
        RECT 229.950 208.500 232.050 208.950 ;
        RECT 265.950 209.400 283.050 210.600 ;
        RECT 265.950 208.800 268.050 209.400 ;
        RECT 280.950 208.950 283.050 209.400 ;
        RECT 295.950 210.600 298.050 210.900 ;
        RECT 299.400 210.600 300.600 212.400 ;
        RECT 295.950 209.400 300.600 210.600 ;
        RECT 301.950 210.600 304.050 211.050 ;
        RECT 313.950 210.600 316.050 210.900 ;
        RECT 301.950 209.400 316.050 210.600 ;
        RECT 295.950 208.800 298.050 209.400 ;
        RECT 301.950 208.950 304.050 209.400 ;
        RECT 313.950 208.800 316.050 209.400 ;
        RECT 325.950 210.450 328.050 210.900 ;
        RECT 334.950 210.450 337.050 210.900 ;
        RECT 325.950 209.250 337.050 210.450 ;
        RECT 325.950 208.800 328.050 209.250 ;
        RECT 334.950 208.800 337.050 209.250 ;
        RECT 340.950 210.600 343.050 210.900 ;
        RECT 358.950 210.600 361.050 210.900 ;
        RECT 340.950 210.450 361.050 210.600 ;
        RECT 364.800 210.450 366.900 210.900 ;
        RECT 340.950 209.400 366.900 210.450 ;
        RECT 340.950 208.800 343.050 209.400 ;
        RECT 358.950 209.250 366.900 209.400 ;
        RECT 358.950 208.800 361.050 209.250 ;
        RECT 364.800 208.800 366.900 209.250 ;
        RECT 367.950 210.600 370.050 211.050 ;
        RECT 379.950 210.600 382.050 211.050 ;
        RECT 367.950 209.400 382.050 210.600 ;
        RECT 367.950 208.950 370.050 209.400 ;
        RECT 379.950 208.950 382.050 209.400 ;
        RECT 403.950 210.600 406.050 210.900 ;
        RECT 425.400 210.600 426.600 215.100 ;
        RECT 568.950 214.950 571.050 215.400 ;
        RECT 577.950 215.100 580.050 215.400 ;
        RECT 589.950 216.750 592.050 217.200 ;
        RECT 601.950 216.750 604.050 217.200 ;
        RECT 589.950 215.550 604.050 216.750 ;
        RECT 589.950 215.100 592.050 215.550 ;
        RECT 601.950 215.100 604.050 215.550 ;
        RECT 607.950 215.100 610.050 217.200 ;
        RECT 631.950 216.600 634.050 217.200 ;
        RECT 640.950 216.600 643.050 217.050 ;
        RECT 631.950 215.400 643.050 216.600 ;
        RECT 631.950 215.100 634.050 215.400 ;
        RECT 475.950 210.600 478.050 210.900 ;
        RECT 403.950 209.400 426.600 210.600 ;
        RECT 460.950 209.400 478.050 210.600 ;
        RECT 403.950 208.800 406.050 209.400 ;
        RECT 181.950 207.600 184.050 207.750 ;
        RECT 208.950 207.600 211.050 208.050 ;
        RECT 181.950 206.400 211.050 207.600 ;
        RECT 181.950 205.650 184.050 206.400 ;
        RECT 208.950 205.950 211.050 206.400 ;
        RECT 280.950 207.600 283.050 207.900 ;
        RECT 326.400 207.600 327.600 208.800 ;
        RECT 280.950 206.400 327.600 207.600 ;
        RECT 407.400 207.600 408.600 209.400 ;
        RECT 460.950 208.500 463.050 209.400 ;
        RECT 475.950 208.800 478.050 209.400 ;
        RECT 484.950 210.450 487.050 211.050 ;
        RECT 493.950 210.450 496.050 210.900 ;
        RECT 484.950 209.250 496.050 210.450 ;
        RECT 484.950 208.950 487.050 209.250 ;
        RECT 493.950 208.800 496.050 209.250 ;
        RECT 505.950 210.600 508.050 211.050 ;
        RECT 571.950 210.600 574.050 211.050 ;
        RECT 604.950 210.600 607.050 210.900 ;
        RECT 505.950 210.150 535.050 210.600 ;
        RECT 568.800 210.150 570.900 210.600 ;
        RECT 505.950 209.400 570.900 210.150 ;
        RECT 505.950 208.950 508.050 209.400 ;
        RECT 532.950 208.950 570.900 209.400 ;
        RECT 571.950 209.400 607.050 210.600 ;
        RECT 608.400 210.600 609.600 215.100 ;
        RECT 640.950 214.950 643.050 215.400 ;
        RECT 655.950 216.600 658.050 217.200 ;
        RECT 664.950 216.600 667.050 217.050 ;
        RECT 655.950 215.400 667.050 216.600 ;
        RECT 655.950 215.100 658.050 215.400 ;
        RECT 664.950 214.950 667.050 215.400 ;
        RECT 682.950 215.100 685.050 217.200 ;
        RECT 694.950 216.600 697.050 217.050 ;
        RECT 758.400 216.600 759.600 218.400 ;
        RECT 766.950 217.950 769.050 218.400 ;
        RECT 829.950 219.600 832.050 220.050 ;
        RECT 835.950 219.600 838.050 220.050 ;
        RECT 829.950 218.400 838.050 219.600 ;
        RECT 829.950 217.950 832.050 218.400 ;
        RECT 835.950 217.950 838.050 218.400 ;
        RECT 847.950 219.600 850.050 220.050 ;
        RECT 859.950 219.600 862.050 220.050 ;
        RECT 871.950 219.600 874.050 220.050 ;
        RECT 847.950 218.400 858.600 219.600 ;
        RECT 847.950 217.950 850.050 218.400 ;
        RECT 694.950 215.400 759.600 216.600 ;
        RECT 683.400 213.600 684.600 215.100 ;
        RECT 694.950 214.950 697.050 215.400 ;
        RECT 760.950 214.950 763.050 217.050 ;
        RECT 745.950 213.600 748.050 214.050 ;
        RECT 683.400 212.400 748.050 213.600 ;
        RECT 745.950 211.950 748.050 212.400 ;
        RECT 613.950 210.600 616.050 211.050 ;
        RECT 608.400 209.400 616.050 210.600 ;
        RECT 571.950 208.950 574.050 209.400 ;
        RECT 532.950 208.500 535.050 208.950 ;
        RECT 568.800 208.500 570.900 208.950 ;
        RECT 604.950 208.800 607.050 209.400 ;
        RECT 613.950 208.950 616.050 209.400 ;
        RECT 761.400 208.050 762.600 214.950 ;
        RECT 769.950 213.600 772.050 217.050 ;
        RECT 781.950 216.600 784.050 217.200 ;
        RECT 796.950 216.600 799.050 217.200 ;
        RECT 764.400 213.000 772.050 213.600 ;
        RECT 773.400 215.400 784.050 216.600 ;
        RECT 764.400 212.400 771.600 213.000 ;
        RECT 764.400 210.900 765.600 212.400 ;
        RECT 773.400 211.050 774.600 215.400 ;
        RECT 781.950 215.100 784.050 215.400 ;
        RECT 785.400 215.400 799.050 216.600 ;
        RECT 763.950 208.800 766.050 210.900 ;
        RECT 769.950 209.400 774.600 211.050 ;
        RECT 785.400 210.900 786.600 215.400 ;
        RECT 796.950 215.100 799.050 215.400 ;
        RECT 826.950 214.950 829.050 217.050 ;
        RECT 853.950 214.950 856.050 217.050 ;
        RECT 827.400 211.050 828.600 214.950 ;
        RECT 854.400 211.050 855.600 214.950 ;
        RECT 857.400 213.600 858.600 218.400 ;
        RECT 859.950 218.400 874.050 219.600 ;
        RECT 859.950 217.950 862.050 218.400 ;
        RECT 871.950 217.950 874.050 218.400 ;
        RECT 877.950 217.950 880.050 220.050 ;
        RECT 857.400 212.400 861.600 213.600 ;
        RECT 769.950 208.950 774.000 209.400 ;
        RECT 784.950 208.800 787.050 210.900 ;
        RECT 826.950 208.950 829.050 211.050 ;
        RECT 835.950 210.450 838.050 210.900 ;
        RECT 844.950 210.450 847.050 210.900 ;
        RECT 835.950 209.250 847.050 210.450 ;
        RECT 835.950 208.800 838.050 209.250 ;
        RECT 844.950 208.800 847.050 209.250 ;
        RECT 853.950 208.950 856.050 211.050 ;
        RECT 860.400 210.600 861.600 212.400 ;
        RECT 871.950 210.600 874.050 210.900 ;
        RECT 860.400 209.400 874.050 210.600 ;
        RECT 871.950 208.800 874.050 209.400 ;
        RECT 481.950 207.600 484.050 208.050 ;
        RECT 407.400 206.400 484.050 207.600 ;
        RECT 280.950 205.800 283.050 206.400 ;
        RECT 481.950 205.950 484.050 206.400 ;
        RECT 514.950 207.600 517.050 208.050 ;
        RECT 520.950 207.600 523.050 208.050 ;
        RECT 514.950 206.400 523.050 207.600 ;
        RECT 514.950 205.950 517.050 206.400 ;
        RECT 520.950 205.950 523.050 206.400 ;
        RECT 616.950 207.600 619.050 208.050 ;
        RECT 628.950 207.600 631.050 208.050 ;
        RECT 616.950 206.400 631.050 207.600 ;
        RECT 616.950 205.950 619.050 206.400 ;
        RECT 628.950 205.950 631.050 206.400 ;
        RECT 757.950 206.400 762.600 208.050 ;
        RECT 878.400 207.600 879.600 217.950 ;
        RECT 883.950 207.600 886.050 208.050 ;
        RECT 878.400 206.400 886.050 207.600 ;
        RECT 757.950 205.950 762.000 206.400 ;
        RECT 883.950 205.950 886.050 206.400 ;
        RECT 34.950 204.600 37.050 205.050 ;
        RECT 52.950 204.600 55.050 205.050 ;
        RECT 34.950 203.400 55.050 204.600 ;
        RECT 34.950 202.950 37.050 203.400 ;
        RECT 52.950 202.950 55.050 203.400 ;
        RECT 67.950 204.600 70.050 205.050 ;
        RECT 79.950 204.600 82.050 205.050 ;
        RECT 100.950 204.600 103.050 205.050 ;
        RECT 136.950 204.600 139.050 205.050 ;
        RECT 67.950 203.400 139.050 204.600 ;
        RECT 67.950 202.950 70.050 203.400 ;
        RECT 79.950 202.950 82.050 203.400 ;
        RECT 100.950 202.950 103.050 203.400 ;
        RECT 136.950 202.950 139.050 203.400 ;
        RECT 142.950 204.600 145.050 205.050 ;
        RECT 151.950 204.600 154.050 205.050 ;
        RECT 172.950 204.600 175.050 205.050 ;
        RECT 142.950 203.400 175.050 204.600 ;
        RECT 142.950 202.950 145.050 203.400 ;
        RECT 151.950 202.950 154.050 203.400 ;
        RECT 172.950 202.950 175.050 203.400 ;
        RECT 196.950 204.600 199.050 205.050 ;
        RECT 463.950 204.600 466.050 205.050 ;
        RECT 196.950 203.400 466.050 204.600 ;
        RECT 196.950 202.950 199.050 203.400 ;
        RECT 463.950 202.950 466.050 203.400 ;
        RECT 490.950 204.600 493.050 205.050 ;
        RECT 505.950 204.600 508.050 205.050 ;
        RECT 490.950 203.400 508.050 204.600 ;
        RECT 490.950 202.950 493.050 203.400 ;
        RECT 505.950 202.950 508.050 203.400 ;
        RECT 580.950 204.600 583.050 205.050 ;
        RECT 589.950 204.600 592.050 205.050 ;
        RECT 580.950 203.400 592.050 204.600 ;
        RECT 580.950 202.950 583.050 203.400 ;
        RECT 589.950 202.950 592.050 203.400 ;
        RECT 631.950 204.600 634.050 205.050 ;
        RECT 658.800 204.600 660.900 205.050 ;
        RECT 631.950 203.400 660.900 204.600 ;
        RECT 631.950 202.950 634.050 203.400 ;
        RECT 658.800 202.950 660.900 203.400 ;
        RECT 661.950 204.600 664.050 205.050 ;
        RECT 733.950 204.600 736.050 204.900 ;
        RECT 661.950 203.400 736.050 204.600 ;
        RECT 661.950 202.950 664.050 203.400 ;
        RECT 733.950 202.800 736.050 203.400 ;
        RECT 784.950 204.600 787.050 205.050 ;
        RECT 835.950 204.600 838.050 205.050 ;
        RECT 784.950 203.400 838.050 204.600 ;
        RECT 784.950 202.950 787.050 203.400 ;
        RECT 835.950 202.950 838.050 203.400 ;
        RECT 79.950 201.600 82.050 201.900 ;
        RECT 97.950 201.600 100.050 202.050 ;
        RECT 79.950 200.400 100.050 201.600 ;
        RECT 79.950 199.800 82.050 200.400 ;
        RECT 97.950 199.950 100.050 200.400 ;
        RECT 178.950 201.600 181.050 202.050 ;
        RECT 184.950 201.600 187.050 202.050 ;
        RECT 178.950 200.400 187.050 201.600 ;
        RECT 178.950 199.950 181.050 200.400 ;
        RECT 184.950 199.950 187.050 200.400 ;
        RECT 277.950 201.600 280.050 202.050 ;
        RECT 289.950 201.600 292.050 202.050 ;
        RECT 277.950 200.400 292.050 201.600 ;
        RECT 277.950 199.950 280.050 200.400 ;
        RECT 289.950 199.950 292.050 200.400 ;
        RECT 376.950 201.600 379.050 202.050 ;
        RECT 415.950 201.600 418.050 202.050 ;
        RECT 421.950 201.600 424.050 202.050 ;
        RECT 376.950 200.400 424.050 201.600 ;
        RECT 376.950 199.950 379.050 200.400 ;
        RECT 415.950 199.950 418.050 200.400 ;
        RECT 421.950 199.950 424.050 200.400 ;
        RECT 487.950 201.600 490.050 202.050 ;
        RECT 499.950 201.600 502.050 202.050 ;
        RECT 487.950 200.400 502.050 201.600 ;
        RECT 487.950 199.950 490.050 200.400 ;
        RECT 499.950 199.950 502.050 200.400 ;
        RECT 508.950 201.600 511.050 202.050 ;
        RECT 514.950 201.600 517.050 202.050 ;
        RECT 508.950 200.400 517.050 201.600 ;
        RECT 508.950 199.950 511.050 200.400 ;
        RECT 514.950 199.950 517.050 200.400 ;
        RECT 640.950 201.600 643.050 202.050 ;
        RECT 679.950 201.600 682.050 202.050 ;
        RECT 700.950 201.600 703.050 202.050 ;
        RECT 721.950 201.600 724.050 202.050 ;
        RECT 640.950 200.400 724.050 201.600 ;
        RECT 640.950 199.950 643.050 200.400 ;
        RECT 679.950 199.950 682.050 200.400 ;
        RECT 700.950 199.950 703.050 200.400 ;
        RECT 721.950 199.950 724.050 200.400 ;
        RECT 748.950 201.600 751.050 202.050 ;
        RECT 769.950 201.600 772.050 202.050 ;
        RECT 748.950 200.400 772.050 201.600 ;
        RECT 748.950 199.950 751.050 200.400 ;
        RECT 769.950 199.950 772.050 200.400 ;
        RECT 838.950 201.600 841.050 202.050 ;
        RECT 856.950 201.600 859.050 202.050 ;
        RECT 838.950 200.400 859.050 201.600 ;
        RECT 838.950 199.950 841.050 200.400 ;
        RECT 856.950 199.950 859.050 200.400 ;
        RECT 40.950 198.600 43.050 199.050 ;
        RECT 52.950 198.600 55.050 199.050 ;
        RECT 40.950 197.400 55.050 198.600 ;
        RECT 40.950 196.950 43.050 197.400 ;
        RECT 52.950 196.950 55.050 197.400 ;
        RECT 73.950 198.600 76.050 199.050 ;
        RECT 94.950 198.600 97.050 199.050 ;
        RECT 73.950 197.400 97.050 198.600 ;
        RECT 73.950 196.950 76.050 197.400 ;
        RECT 94.950 196.950 97.050 197.400 ;
        RECT 124.950 198.600 127.050 199.050 ;
        RECT 166.950 198.600 169.050 199.050 ;
        RECT 124.950 197.400 169.050 198.600 ;
        RECT 124.950 196.950 127.050 197.400 ;
        RECT 166.950 196.950 169.050 197.400 ;
        RECT 475.950 198.600 478.050 199.050 ;
        RECT 523.950 198.600 526.050 199.050 ;
        RECT 538.950 198.600 541.050 199.050 ;
        RECT 475.950 197.400 541.050 198.600 ;
        RECT 475.950 196.950 478.050 197.400 ;
        RECT 523.950 196.950 526.050 197.400 ;
        RECT 538.950 196.950 541.050 197.400 ;
        RECT 610.950 198.600 613.050 199.050 ;
        RECT 631.950 198.600 634.050 199.050 ;
        RECT 610.950 197.400 634.050 198.600 ;
        RECT 610.950 196.950 613.050 197.400 ;
        RECT 631.950 196.950 634.050 197.400 ;
        RECT 643.950 198.600 646.050 199.050 ;
        RECT 703.800 198.600 705.900 199.050 ;
        RECT 643.950 197.400 705.900 198.600 ;
        RECT 643.950 196.950 646.050 197.400 ;
        RECT 703.800 196.950 705.900 197.400 ;
        RECT 706.950 198.600 709.050 199.050 ;
        RECT 745.950 198.600 748.050 199.050 ;
        RECT 706.950 197.400 748.050 198.600 ;
        RECT 706.950 196.950 709.050 197.400 ;
        RECT 745.950 196.950 748.050 197.400 ;
        RECT 28.950 195.600 31.050 196.050 ;
        RECT 34.950 195.600 37.050 196.050 ;
        RECT 28.950 194.400 37.050 195.600 ;
        RECT 28.950 193.950 31.050 194.400 ;
        RECT 34.950 193.950 37.050 194.400 ;
        RECT 97.950 195.600 100.050 196.050 ;
        RECT 142.950 195.600 145.050 196.050 ;
        RECT 97.950 194.400 145.050 195.600 ;
        RECT 97.950 193.950 100.050 194.400 ;
        RECT 142.950 193.950 145.050 194.400 ;
        RECT 172.950 195.600 175.050 196.050 ;
        RECT 214.950 195.600 217.050 196.050 ;
        RECT 172.950 194.400 217.050 195.600 ;
        RECT 172.950 193.950 175.050 194.400 ;
        RECT 214.950 193.950 217.050 194.400 ;
        RECT 313.950 195.600 316.050 196.050 ;
        RECT 319.950 195.600 322.050 196.050 ;
        RECT 349.950 195.600 352.050 196.050 ;
        RECT 361.950 195.600 364.050 196.050 ;
        RECT 313.950 194.400 364.050 195.600 ;
        RECT 313.950 193.950 316.050 194.400 ;
        RECT 319.950 193.950 322.050 194.400 ;
        RECT 349.950 193.950 352.050 194.400 ;
        RECT 361.950 193.950 364.050 194.400 ;
        RECT 565.950 195.600 568.050 196.050 ;
        RECT 577.950 195.600 580.050 196.050 ;
        RECT 565.950 194.400 580.050 195.600 ;
        RECT 565.950 193.950 568.050 194.400 ;
        RECT 577.950 193.950 580.050 194.400 ;
        RECT 613.950 195.600 616.050 196.050 ;
        RECT 634.950 195.600 637.050 196.050 ;
        RECT 613.950 194.400 637.050 195.600 ;
        RECT 613.950 193.950 616.050 194.400 ;
        RECT 634.950 193.950 637.050 194.400 ;
        RECT 664.950 195.600 667.050 196.050 ;
        RECT 682.950 195.600 685.050 196.050 ;
        RECT 664.950 194.400 685.050 195.600 ;
        RECT 664.950 193.950 667.050 194.400 ;
        RECT 682.950 193.950 685.050 194.400 ;
        RECT 715.950 195.600 718.050 196.050 ;
        RECT 799.950 195.600 802.050 196.050 ;
        RECT 808.950 195.600 811.050 196.050 ;
        RECT 715.950 194.400 811.050 195.600 ;
        RECT 715.950 193.950 718.050 194.400 ;
        RECT 799.950 193.950 802.050 194.400 ;
        RECT 808.950 193.950 811.050 194.400 ;
        RECT 823.950 195.600 826.050 196.050 ;
        RECT 850.950 195.600 853.050 196.050 ;
        RECT 856.950 195.600 859.050 196.050 ;
        RECT 823.950 194.400 859.050 195.600 ;
        RECT 823.950 193.950 826.050 194.400 ;
        RECT 850.950 193.950 853.050 194.400 ;
        RECT 856.950 193.950 859.050 194.400 ;
        RECT 22.950 192.600 25.050 193.050 ;
        RECT 46.950 192.600 49.050 193.050 ;
        RECT 22.950 191.400 49.050 192.600 ;
        RECT 22.950 190.950 25.050 191.400 ;
        RECT 46.950 190.950 49.050 191.400 ;
        RECT 307.950 192.600 310.050 193.050 ;
        RECT 358.950 192.600 361.050 193.050 ;
        RECT 307.950 191.400 361.050 192.600 ;
        RECT 307.950 190.950 310.050 191.400 ;
        RECT 358.950 190.950 361.050 191.400 ;
        RECT 364.950 192.600 367.050 193.050 ;
        RECT 409.950 192.600 412.050 193.050 ;
        RECT 364.950 191.400 412.050 192.600 ;
        RECT 364.950 190.950 367.050 191.400 ;
        RECT 409.950 190.950 412.050 191.400 ;
        RECT 421.950 192.600 424.050 193.050 ;
        RECT 451.950 192.600 454.050 193.050 ;
        RECT 421.950 191.400 454.050 192.600 ;
        RECT 421.950 190.950 424.050 191.400 ;
        RECT 451.950 190.950 454.050 191.400 ;
        RECT 469.950 192.600 472.050 193.050 ;
        RECT 535.950 192.600 538.050 193.050 ;
        RECT 469.950 191.400 538.050 192.600 ;
        RECT 469.950 190.950 472.050 191.400 ;
        RECT 535.950 190.950 538.050 191.400 ;
        RECT 544.950 192.600 547.050 193.050 ;
        RECT 574.950 192.600 577.050 193.050 ;
        RECT 610.950 192.600 613.050 193.050 ;
        RECT 544.950 191.400 613.050 192.600 ;
        RECT 544.950 190.950 547.050 191.400 ;
        RECT 574.950 190.950 577.050 191.400 ;
        RECT 610.950 190.950 613.050 191.400 ;
        RECT 637.950 192.600 640.050 193.050 ;
        RECT 796.950 192.600 799.050 193.050 ;
        RECT 637.950 191.400 799.050 192.600 ;
        RECT 637.950 190.950 640.050 191.400 ;
        RECT 796.950 190.950 799.050 191.400 ;
        RECT 211.950 189.600 214.050 190.050 ;
        RECT 259.950 189.600 262.050 190.050 ;
        RECT 211.950 188.400 262.050 189.600 ;
        RECT 211.950 187.950 214.050 188.400 ;
        RECT 259.950 187.950 262.050 188.400 ;
        RECT 442.950 189.600 445.050 190.050 ;
        RECT 451.950 189.600 454.050 189.900 ;
        RECT 547.950 189.600 550.050 190.050 ;
        RECT 442.950 188.400 550.050 189.600 ;
        RECT 442.950 187.950 445.050 188.400 ;
        RECT 451.950 187.800 454.050 188.400 ;
        RECT 547.950 187.950 550.050 188.400 ;
        RECT 619.950 189.600 622.050 190.050 ;
        RECT 652.950 189.600 655.050 190.050 ;
        RECT 619.950 188.400 655.050 189.600 ;
        RECT 619.950 187.950 622.050 188.400 ;
        RECT 652.950 187.950 655.050 188.400 ;
        RECT 694.950 189.600 697.050 190.050 ;
        RECT 715.950 189.600 718.050 190.050 ;
        RECT 694.950 188.400 718.050 189.600 ;
        RECT 694.950 187.950 697.050 188.400 ;
        RECT 715.950 187.950 718.050 188.400 ;
        RECT 829.950 189.600 832.050 190.050 ;
        RECT 841.950 189.600 844.050 190.050 ;
        RECT 829.950 188.400 844.050 189.600 ;
        RECT 829.950 187.950 832.050 188.400 ;
        RECT 841.950 187.950 844.050 188.400 ;
        RECT 871.950 189.600 874.050 190.050 ;
        RECT 886.950 189.600 889.050 190.050 ;
        RECT 871.950 188.400 889.050 189.600 ;
        RECT 871.950 187.950 874.050 188.400 ;
        RECT 886.950 187.950 889.050 188.400 ;
        RECT 37.950 183.600 40.050 184.200 ;
        RECT 32.400 182.400 40.050 183.600 ;
        RECT 32.400 180.600 33.600 182.400 ;
        RECT 37.950 182.100 40.050 182.400 ;
        RECT 43.950 180.600 46.050 184.050 ;
        RECT 49.950 183.750 52.050 184.200 ;
        RECT 61.950 183.750 64.050 184.200 ;
        RECT 49.950 182.550 64.050 183.750 ;
        RECT 85.950 183.600 88.050 184.200 ;
        RECT 49.950 182.100 52.050 182.550 ;
        RECT 61.950 182.100 64.050 182.550 ;
        RECT 65.400 182.400 88.050 183.600 ;
        RECT 97.950 182.400 100.050 184.500 ;
        RECT 126.000 183.600 130.050 184.050 ;
        RECT 14.400 179.400 33.600 180.600 ;
        RECT 38.400 180.000 46.050 180.600 ;
        RECT 38.400 179.400 45.600 180.000 ;
        RECT 14.400 177.900 15.600 179.400 ;
        RECT 13.950 175.800 16.050 177.900 ;
        RECT 34.950 177.600 37.050 177.900 ;
        RECT 38.400 177.600 39.600 179.400 ;
        RECT 65.400 177.900 66.600 182.400 ;
        RECT 85.950 182.100 88.050 182.400 ;
        RECT 34.950 176.400 39.600 177.600 ;
        RECT 52.950 177.450 55.050 177.900 ;
        RECT 58.950 177.450 61.050 177.900 ;
        RECT 34.950 175.800 37.050 176.400 ;
        RECT 52.950 176.250 61.050 177.450 ;
        RECT 52.950 175.800 55.050 176.250 ;
        RECT 58.950 175.800 61.050 176.250 ;
        RECT 64.950 175.800 67.050 177.900 ;
        RECT 82.950 177.600 85.050 177.900 ;
        RECT 98.400 177.600 99.600 182.400 ;
        RECT 125.400 181.950 130.050 183.600 ;
        RECT 133.950 183.600 136.050 184.050 ;
        RECT 142.950 183.600 145.050 184.200 ;
        RECT 133.950 182.400 145.050 183.600 ;
        RECT 181.950 183.600 184.050 187.050 ;
        RECT 328.950 186.600 331.050 187.050 ;
        RECT 352.950 186.600 355.050 187.050 ;
        RECT 328.950 185.400 355.050 186.600 ;
        RECT 328.950 184.950 331.050 185.400 ;
        RECT 352.950 184.950 355.050 185.400 ;
        RECT 400.950 186.600 403.050 187.050 ;
        RECT 412.950 186.600 415.050 187.050 ;
        RECT 400.950 185.400 415.050 186.600 ;
        RECT 400.950 184.950 403.050 185.400 ;
        RECT 412.950 184.950 415.050 185.400 ;
        RECT 424.950 186.600 427.050 187.050 ;
        RECT 430.950 186.600 433.050 187.050 ;
        RECT 517.950 186.600 520.050 187.050 ;
        RECT 424.950 185.400 520.050 186.600 ;
        RECT 424.950 184.950 427.050 185.400 ;
        RECT 430.950 184.950 433.050 185.400 ;
        RECT 517.950 184.950 520.050 185.400 ;
        RECT 595.950 186.600 598.050 187.050 ;
        RECT 613.950 186.600 616.050 187.050 ;
        RECT 649.950 186.600 652.050 187.050 ;
        RECT 595.950 185.400 652.050 186.600 ;
        RECT 595.950 184.950 598.050 185.400 ;
        RECT 613.950 184.950 616.050 185.400 ;
        RECT 649.950 184.950 652.050 185.400 ;
        RECT 658.950 186.600 661.050 187.050 ;
        RECT 676.950 186.600 679.050 187.050 ;
        RECT 658.950 185.400 679.050 186.600 ;
        RECT 658.950 184.950 661.050 185.400 ;
        RECT 676.950 184.950 679.050 185.400 ;
        RECT 724.950 186.600 727.050 187.050 ;
        RECT 730.950 186.600 733.050 187.050 ;
        RECT 724.950 185.400 733.050 186.600 ;
        RECT 724.950 184.950 727.050 185.400 ;
        RECT 730.950 184.950 733.050 185.400 ;
        RECT 739.950 186.600 742.050 187.050 ;
        RECT 790.950 186.600 793.050 187.200 ;
        RECT 802.950 186.600 805.050 187.050 ;
        RECT 811.950 186.600 814.050 187.050 ;
        RECT 739.950 185.400 759.600 186.600 ;
        RECT 739.950 184.950 742.050 185.400 ;
        RECT 187.950 183.600 190.050 184.200 ;
        RECT 220.950 183.600 223.050 184.500 ;
        RECT 268.950 183.600 271.050 184.200 ;
        RECT 181.950 183.000 190.050 183.600 ;
        RECT 182.400 182.400 190.050 183.000 ;
        RECT 133.950 181.950 136.050 182.400 ;
        RECT 142.950 182.100 145.050 182.400 ;
        RECT 187.950 182.100 190.050 182.400 ;
        RECT 218.400 182.400 223.050 183.600 ;
        RECT 239.400 182.400 271.050 183.600 ;
        RECT 125.400 177.600 126.600 181.950 ;
        RECT 152.400 179.400 183.600 180.600 ;
        RECT 152.400 177.900 153.600 179.400 ;
        RECT 82.950 176.400 99.600 177.600 ;
        RECT 82.950 175.800 85.050 176.400 ;
        RECT 124.950 175.500 127.050 177.600 ;
        RECT 139.950 177.450 142.050 177.900 ;
        RECT 151.950 177.450 154.050 177.900 ;
        RECT 139.950 176.250 154.050 177.450 ;
        RECT 139.950 175.800 142.050 176.250 ;
        RECT 151.950 175.800 154.050 176.250 ;
        RECT 163.950 177.450 166.050 177.900 ;
        RECT 175.950 177.450 178.050 177.900 ;
        RECT 163.950 176.250 178.050 177.450 ;
        RECT 182.400 177.600 183.600 179.400 ;
        RECT 184.950 177.600 187.050 177.900 ;
        RECT 182.400 176.400 187.050 177.600 ;
        RECT 163.950 175.800 166.050 176.250 ;
        RECT 175.950 175.800 178.050 176.250 ;
        RECT 184.950 175.800 187.050 176.400 ;
        RECT 214.950 177.600 217.050 177.900 ;
        RECT 218.400 177.600 219.600 182.400 ;
        RECT 239.400 177.600 240.600 182.400 ;
        RECT 268.950 182.100 271.050 182.400 ;
        RECT 274.950 182.100 277.050 184.200 ;
        RECT 283.950 183.600 286.050 184.050 ;
        RECT 289.950 183.600 292.050 184.200 ;
        RECT 283.950 182.400 292.050 183.600 ;
        RECT 275.400 180.600 276.600 182.100 ;
        RECT 283.950 181.950 286.050 182.400 ;
        RECT 289.950 182.100 292.050 182.400 ;
        RECT 295.950 182.100 298.050 184.200 ;
        RECT 319.950 183.750 322.050 184.200 ;
        RECT 325.950 183.750 328.050 184.200 ;
        RECT 319.950 182.550 328.050 183.750 ;
        RECT 319.950 182.100 322.050 182.550 ;
        RECT 325.950 182.100 328.050 182.550 ;
        RECT 358.950 183.600 361.050 184.050 ;
        RECT 367.950 183.600 370.050 184.200 ;
        RECT 358.950 182.400 370.050 183.600 ;
        RECT 272.400 179.400 276.600 180.600 ;
        RECT 214.950 176.400 219.600 177.600 ;
        RECT 214.950 175.800 217.050 176.400 ;
        RECT 238.950 175.500 241.050 177.600 ;
        RECT 247.950 177.150 250.050 177.600 ;
        RECT 253.950 177.150 256.050 177.600 ;
        RECT 247.950 175.950 256.050 177.150 ;
        RECT 247.950 175.500 250.050 175.950 ;
        RECT 253.950 175.500 256.050 175.950 ;
        RECT 259.950 177.450 262.050 177.900 ;
        RECT 265.950 177.450 268.050 177.900 ;
        RECT 259.950 176.250 268.050 177.450 ;
        RECT 259.950 175.800 262.050 176.250 ;
        RECT 265.950 175.800 268.050 176.250 ;
        RECT 272.400 175.050 273.600 179.400 ;
        RECT 296.400 177.600 297.600 182.100 ;
        RECT 358.950 181.950 361.050 182.400 ;
        RECT 367.950 182.100 370.050 182.400 ;
        RECT 391.950 183.750 394.050 184.200 ;
        RECT 397.950 183.750 400.050 184.200 ;
        RECT 391.950 182.550 400.050 183.750 ;
        RECT 391.950 182.100 394.050 182.550 ;
        RECT 397.950 182.100 400.050 182.550 ;
        RECT 436.950 182.100 439.050 184.200 ;
        RECT 510.000 183.600 514.050 184.050 ;
        RECT 316.950 177.600 319.050 177.900 ;
        RECT 296.400 176.400 319.050 177.600 ;
        RECT 316.950 175.800 319.050 176.400 ;
        RECT 352.950 177.450 355.050 177.900 ;
        RECT 364.950 177.450 367.050 177.900 ;
        RECT 352.950 176.250 367.050 177.450 ;
        RECT 352.950 175.800 355.050 176.250 ;
        RECT 364.950 175.800 367.050 176.250 ;
        RECT 370.950 177.450 373.050 177.900 ;
        RECT 376.950 177.450 379.050 177.900 ;
        RECT 370.950 176.250 379.050 177.450 ;
        RECT 370.950 175.800 373.050 176.250 ;
        RECT 376.950 175.800 379.050 176.250 ;
        RECT 412.950 177.450 415.050 177.900 ;
        RECT 424.950 177.450 427.050 177.900 ;
        RECT 412.950 176.250 427.050 177.450 ;
        RECT 437.400 177.600 438.600 182.100 ;
        RECT 509.400 181.950 514.050 183.600 ;
        RECT 529.950 183.600 532.050 184.200 ;
        RECT 586.950 183.600 589.050 184.500 ;
        RECT 758.400 184.200 759.600 185.400 ;
        RECT 790.950 185.400 805.050 186.600 ;
        RECT 790.950 185.100 793.050 185.400 ;
        RECT 802.950 184.950 805.050 185.400 ;
        RECT 806.400 185.400 814.050 186.600 ;
        RECT 529.950 182.400 589.050 183.600 ;
        RECT 598.950 183.750 601.050 184.200 ;
        RECT 607.950 183.750 610.050 184.200 ;
        RECT 598.950 182.550 610.050 183.750 ;
        RECT 529.950 182.100 532.050 182.400 ;
        RECT 454.950 177.600 457.050 177.900 ;
        RECT 437.400 176.400 457.050 177.600 ;
        RECT 412.950 175.800 415.050 176.250 ;
        RECT 424.950 175.800 427.050 176.250 ;
        RECT 454.950 175.800 457.050 176.400 ;
        RECT 463.950 177.600 466.050 178.050 ;
        RECT 472.950 177.600 475.050 177.900 ;
        RECT 509.400 177.600 510.600 181.950 ;
        RECT 517.950 177.600 520.050 178.050 ;
        RECT 551.400 177.900 552.600 182.400 ;
        RECT 587.400 180.600 588.600 182.400 ;
        RECT 598.950 182.100 601.050 182.550 ;
        RECT 607.950 182.100 610.050 182.550 ;
        RECT 628.950 183.600 631.050 184.200 ;
        RECT 643.950 183.600 646.050 184.050 ;
        RECT 628.950 182.400 646.050 183.600 ;
        RECT 628.950 182.100 631.050 182.400 ;
        RECT 643.950 181.950 646.050 182.400 ;
        RECT 670.950 183.600 673.050 184.050 ;
        RECT 757.950 183.750 760.050 184.200 ;
        RECT 763.950 183.750 766.050 184.200 ;
        RECT 670.950 182.400 687.600 183.600 ;
        RECT 670.950 181.950 673.050 182.400 ;
        RECT 587.400 179.400 609.600 180.600 ;
        RECT 526.950 177.600 529.050 177.900 ;
        RECT 463.950 176.400 475.050 177.600 ;
        RECT 463.950 175.950 466.050 176.400 ;
        RECT 472.950 175.800 475.050 176.400 ;
        RECT 508.950 175.500 511.050 177.600 ;
        RECT 517.950 176.400 529.050 177.600 ;
        RECT 517.950 175.950 520.050 176.400 ;
        RECT 526.950 175.800 529.050 176.400 ;
        RECT 538.950 177.450 541.050 177.900 ;
        RECT 544.950 177.450 547.050 177.900 ;
        RECT 538.950 176.250 547.050 177.450 ;
        RECT 538.950 175.800 541.050 176.250 ;
        RECT 544.950 175.800 547.050 176.250 ;
        RECT 550.950 175.800 553.050 177.900 ;
        RECT 577.950 177.450 580.050 177.900 ;
        RECT 604.950 177.450 607.050 177.900 ;
        RECT 577.950 176.250 607.050 177.450 ;
        RECT 608.400 177.600 609.600 179.400 ;
        RECT 686.400 177.900 687.600 182.400 ;
        RECT 757.950 182.550 766.050 183.750 ;
        RECT 790.950 183.600 793.050 184.050 ;
        RECT 757.950 182.100 760.050 182.550 ;
        RECT 763.950 182.100 766.050 182.550 ;
        RECT 767.400 182.400 793.050 183.600 ;
        RECT 767.400 180.600 768.600 182.400 ;
        RECT 790.950 181.950 793.050 182.400 ;
        RECT 746.400 179.400 768.600 180.600 ;
        RECT 625.950 177.600 628.050 177.900 ;
        RECT 608.400 176.400 628.050 177.600 ;
        RECT 577.950 175.800 580.050 176.250 ;
        RECT 604.950 175.800 607.050 176.250 ;
        RECT 625.950 175.800 628.050 176.400 ;
        RECT 655.950 177.450 658.050 177.900 ;
        RECT 664.950 177.450 667.050 177.900 ;
        RECT 655.950 176.250 667.050 177.450 ;
        RECT 655.950 175.800 658.050 176.250 ;
        RECT 664.950 175.800 667.050 176.250 ;
        RECT 685.950 175.800 688.050 177.900 ;
        RECT 736.950 177.600 739.050 178.050 ;
        RECT 742.950 177.600 745.050 177.900 ;
        RECT 746.400 177.600 747.600 179.400 ;
        RECT 806.400 178.050 807.600 185.400 ;
        RECT 811.950 184.950 814.050 185.400 ;
        RECT 814.950 181.950 817.050 184.050 ;
        RECT 815.400 178.050 816.600 181.950 ;
        RECT 823.950 180.600 826.050 184.050 ;
        RECT 826.950 183.600 829.050 187.050 ;
        RECT 853.950 186.600 856.050 187.050 ;
        RECT 853.950 185.400 879.600 186.600 ;
        RECT 853.950 184.950 856.050 185.400 ;
        RECT 835.950 183.600 838.050 184.050 ;
        RECT 841.950 183.600 844.050 183.900 ;
        RECT 826.950 183.000 834.600 183.600 ;
        RECT 827.400 182.400 834.600 183.000 ;
        RECT 823.950 180.000 828.600 180.600 ;
        RECT 824.400 179.400 828.600 180.000 ;
        RECT 781.950 177.600 784.050 177.900 ;
        RECT 736.950 176.400 747.600 177.600 ;
        RECT 776.400 176.400 784.050 177.600 ;
        RECT 736.950 175.950 739.050 176.400 ;
        RECT 742.950 175.800 745.050 176.400 ;
        RECT 40.950 174.600 43.050 175.050 ;
        RECT 46.950 174.600 49.050 175.050 ;
        RECT 40.950 173.400 49.050 174.600 ;
        RECT 40.950 172.950 43.050 173.400 ;
        RECT 46.950 172.950 49.050 173.400 ;
        RECT 73.950 174.600 76.050 175.050 ;
        RECT 79.950 174.600 82.050 175.050 ;
        RECT 73.950 173.400 82.050 174.600 ;
        RECT 73.950 172.950 76.050 173.400 ;
        RECT 79.950 172.950 82.050 173.400 ;
        RECT 190.950 174.600 193.050 175.050 ;
        RECT 196.950 174.600 199.050 175.050 ;
        RECT 190.950 173.400 199.050 174.600 ;
        RECT 190.950 172.950 193.050 173.400 ;
        RECT 196.950 172.950 199.050 173.400 ;
        RECT 268.950 173.400 273.600 175.050 ;
        RECT 280.950 174.600 283.050 175.050 ;
        RECT 298.950 174.600 301.050 175.050 ;
        RECT 280.950 173.400 301.050 174.600 ;
        RECT 268.950 172.950 273.000 173.400 ;
        RECT 280.950 172.950 283.050 173.400 ;
        RECT 298.950 172.950 301.050 173.400 ;
        RECT 466.950 174.600 469.050 175.050 ;
        RECT 475.950 174.600 478.050 175.050 ;
        RECT 466.950 173.400 478.050 174.600 ;
        RECT 466.950 172.950 469.050 173.400 ;
        RECT 475.950 172.950 478.050 173.400 ;
        RECT 508.950 174.600 511.050 175.050 ;
        RECT 559.950 174.600 562.050 175.050 ;
        RECT 508.950 173.400 562.050 174.600 ;
        RECT 508.950 172.950 511.050 173.400 ;
        RECT 559.950 172.950 562.050 173.400 ;
        RECT 652.950 174.600 655.050 175.050 ;
        RECT 673.950 174.600 676.050 175.050 ;
        RECT 652.950 173.400 676.050 174.600 ;
        RECT 652.950 172.950 655.050 173.400 ;
        RECT 673.950 172.950 676.050 173.400 ;
        RECT 88.950 171.600 91.050 172.050 ;
        RECT 133.950 171.600 136.050 172.050 ;
        RECT 88.950 170.400 136.050 171.600 ;
        RECT 88.950 169.950 91.050 170.400 ;
        RECT 133.950 169.950 136.050 170.400 ;
        RECT 148.950 171.600 151.050 172.050 ;
        RECT 274.950 171.600 277.050 172.050 ;
        RECT 148.950 170.400 277.050 171.600 ;
        RECT 148.950 169.950 151.050 170.400 ;
        RECT 274.950 169.950 277.050 170.400 ;
        RECT 304.950 171.600 307.050 172.050 ;
        RECT 316.950 171.600 319.050 172.050 ;
        RECT 304.950 170.400 319.050 171.600 ;
        RECT 304.950 169.950 307.050 170.400 ;
        RECT 316.950 169.950 319.050 170.400 ;
        RECT 325.950 171.600 328.050 172.050 ;
        RECT 388.950 171.600 391.050 172.050 ;
        RECT 325.950 170.400 391.050 171.600 ;
        RECT 325.950 169.950 328.050 170.400 ;
        RECT 388.950 169.950 391.050 170.400 ;
        RECT 397.950 171.600 400.050 172.050 ;
        RECT 433.950 171.600 436.050 172.050 ;
        RECT 397.950 170.400 436.050 171.600 ;
        RECT 397.950 169.950 400.050 170.400 ;
        RECT 433.950 169.950 436.050 170.400 ;
        RECT 568.950 171.600 571.050 172.050 ;
        RECT 619.950 171.600 622.050 172.050 ;
        RECT 568.950 170.400 622.050 171.600 ;
        RECT 568.950 169.950 571.050 170.400 ;
        RECT 619.950 169.950 622.050 170.400 ;
        RECT 715.950 171.600 718.050 172.050 ;
        RECT 776.400 171.600 777.600 176.400 ;
        RECT 781.950 175.800 784.050 176.400 ;
        RECT 805.950 175.950 808.050 178.050 ;
        RECT 815.400 176.400 820.050 178.050 ;
        RECT 827.400 177.900 828.600 179.400 ;
        RECT 833.400 177.900 834.600 182.400 ;
        RECT 835.950 182.400 844.050 183.600 ;
        RECT 835.950 181.950 838.050 182.400 ;
        RECT 841.950 181.800 844.050 182.400 ;
        RECT 850.950 183.600 853.050 184.200 ;
        RECT 850.950 182.400 855.600 183.600 ;
        RECT 850.950 182.100 853.050 182.400 ;
        RECT 816.000 175.950 820.050 176.400 ;
        RECT 826.950 175.800 829.050 177.900 ;
        RECT 832.950 177.600 835.050 177.900 ;
        RECT 847.950 177.600 850.050 177.900 ;
        RECT 832.950 176.400 850.050 177.600 ;
        RECT 832.950 175.800 835.050 176.400 ;
        RECT 847.950 175.800 850.050 176.400 ;
        RECT 854.400 175.050 855.600 182.400 ;
        RECT 865.950 181.950 868.050 184.050 ;
        RECT 866.400 178.050 867.600 181.950 ;
        RECT 878.400 178.050 879.600 185.400 ;
        RECT 865.950 175.950 868.050 178.050 ;
        RECT 877.950 175.950 880.050 178.050 ;
        RECT 778.950 174.600 781.050 175.050 ;
        RECT 811.950 174.600 814.050 175.050 ;
        RECT 778.950 173.400 814.050 174.600 ;
        RECT 778.950 172.950 781.050 173.400 ;
        RECT 811.950 172.950 814.050 173.400 ;
        RECT 850.950 173.400 855.600 175.050 ;
        RECT 850.950 172.950 855.000 173.400 ;
        RECT 715.950 170.400 777.600 171.600 ;
        RECT 817.950 171.600 820.050 172.050 ;
        RECT 835.950 171.600 838.050 172.050 ;
        RECT 817.950 170.400 838.050 171.600 ;
        RECT 715.950 169.950 718.050 170.400 ;
        RECT 817.950 169.950 820.050 170.400 ;
        RECT 835.950 169.950 838.050 170.400 ;
        RECT 844.950 171.600 847.050 172.050 ;
        RECT 874.950 171.600 877.050 172.050 ;
        RECT 844.950 170.400 877.050 171.600 ;
        RECT 844.950 169.950 847.050 170.400 ;
        RECT 874.950 169.950 877.050 170.400 ;
        RECT 169.950 168.600 172.050 169.050 ;
        RECT 214.950 168.600 217.050 169.050 ;
        RECT 169.950 167.400 217.050 168.600 ;
        RECT 169.950 166.950 172.050 167.400 ;
        RECT 214.950 166.950 217.050 167.400 ;
        RECT 679.950 168.600 682.050 169.050 ;
        RECT 691.950 168.600 694.050 169.050 ;
        RECT 679.950 167.400 694.050 168.600 ;
        RECT 679.950 166.950 682.050 167.400 ;
        RECT 691.950 166.950 694.050 167.400 ;
        RECT 757.950 168.600 760.050 169.050 ;
        RECT 817.950 168.600 820.050 168.900 ;
        RECT 757.950 167.400 820.050 168.600 ;
        RECT 757.950 166.950 760.050 167.400 ;
        RECT 817.950 166.800 820.050 167.400 ;
        RECT 871.950 168.600 874.050 169.050 ;
        RECT 880.950 168.600 883.050 169.050 ;
        RECT 871.950 167.400 883.050 168.600 ;
        RECT 871.950 166.950 874.050 167.400 ;
        RECT 880.950 166.950 883.050 167.400 ;
        RECT 268.950 165.600 271.050 166.050 ;
        RECT 430.950 165.600 433.050 166.050 ;
        RECT 511.950 165.600 514.050 166.050 ;
        RECT 268.950 164.400 514.050 165.600 ;
        RECT 268.950 163.950 271.050 164.400 ;
        RECT 430.950 163.950 433.050 164.400 ;
        RECT 511.950 163.950 514.050 164.400 ;
        RECT 748.950 165.600 751.050 166.050 ;
        RECT 823.950 165.600 826.050 166.050 ;
        RECT 748.950 164.400 826.050 165.600 ;
        RECT 748.950 163.950 751.050 164.400 ;
        RECT 823.950 163.950 826.050 164.400 ;
        RECT 271.950 162.600 274.050 163.050 ;
        RECT 343.950 162.600 346.050 163.050 ;
        RECT 271.950 161.400 346.050 162.600 ;
        RECT 271.950 160.950 274.050 161.400 ;
        RECT 343.950 160.950 346.050 161.400 ;
        RECT 379.950 162.600 382.050 163.050 ;
        RECT 418.950 162.600 421.050 163.050 ;
        RECT 379.950 161.400 421.050 162.600 ;
        RECT 379.950 160.950 382.050 161.400 ;
        RECT 418.950 160.950 421.050 161.400 ;
        RECT 598.950 162.600 601.050 163.050 ;
        RECT 634.950 162.600 637.050 163.050 ;
        RECT 598.950 161.400 637.050 162.600 ;
        RECT 598.950 160.950 601.050 161.400 ;
        RECT 634.950 160.950 637.050 161.400 ;
        RECT 694.950 162.600 697.050 163.050 ;
        RECT 751.950 162.600 754.050 163.050 ;
        RECT 694.950 161.400 754.050 162.600 ;
        RECT 694.950 160.950 697.050 161.400 ;
        RECT 751.950 160.950 754.050 161.400 ;
        RECT 853.950 162.600 856.050 163.050 ;
        RECT 886.950 162.600 889.050 163.050 ;
        RECT 853.950 161.400 889.050 162.600 ;
        RECT 853.950 160.950 856.050 161.400 ;
        RECT 886.950 160.950 889.050 161.400 ;
        RECT 178.950 159.600 181.050 160.050 ;
        RECT 367.950 159.600 370.050 160.050 ;
        RECT 178.950 158.400 370.050 159.600 ;
        RECT 178.950 157.950 181.050 158.400 ;
        RECT 367.950 157.950 370.050 158.400 ;
        RECT 406.950 159.600 409.050 160.050 ;
        RECT 442.950 159.600 445.050 160.050 ;
        RECT 406.950 158.400 445.050 159.600 ;
        RECT 406.950 157.950 409.050 158.400 ;
        RECT 442.950 157.950 445.050 158.400 ;
        RECT 502.950 159.600 505.050 160.050 ;
        RECT 514.950 159.600 517.050 160.050 ;
        RECT 502.950 158.400 517.050 159.600 ;
        RECT 502.950 157.950 505.050 158.400 ;
        RECT 514.950 157.950 517.050 158.400 ;
        RECT 769.950 159.600 772.050 160.050 ;
        RECT 826.950 159.600 829.050 160.050 ;
        RECT 769.950 158.400 829.050 159.600 ;
        RECT 769.950 157.950 772.050 158.400 ;
        RECT 826.950 157.950 829.050 158.400 ;
        RECT 154.950 156.600 157.050 157.050 ;
        RECT 274.950 156.600 277.050 157.050 ;
        RECT 154.950 155.400 277.050 156.600 ;
        RECT 154.950 154.950 157.050 155.400 ;
        RECT 274.950 154.950 277.050 155.400 ;
        RECT 472.950 156.600 475.050 157.050 ;
        RECT 508.950 156.600 511.050 157.050 ;
        RECT 472.950 155.400 511.050 156.600 ;
        RECT 472.950 154.950 475.050 155.400 ;
        RECT 508.950 154.950 511.050 155.400 ;
        RECT 574.950 156.600 577.050 157.050 ;
        RECT 631.950 156.600 634.050 157.050 ;
        RECT 574.950 155.400 634.050 156.600 ;
        RECT 574.950 154.950 577.050 155.400 ;
        RECT 631.950 154.950 634.050 155.400 ;
        RECT 667.950 156.600 670.050 157.050 ;
        RECT 733.950 156.600 736.050 157.050 ;
        RECT 667.950 155.400 736.050 156.600 ;
        RECT 667.950 154.950 670.050 155.400 ;
        RECT 733.950 154.950 736.050 155.400 ;
        RECT 145.950 153.600 148.050 154.050 ;
        RECT 313.950 153.600 316.050 154.050 ;
        RECT 145.950 152.400 316.050 153.600 ;
        RECT 145.950 151.950 148.050 152.400 ;
        RECT 313.950 151.950 316.050 152.400 ;
        RECT 526.950 153.600 529.050 154.050 ;
        RECT 535.950 153.600 538.050 154.050 ;
        RECT 526.950 152.400 538.050 153.600 ;
        RECT 526.950 151.950 529.050 152.400 ;
        RECT 535.950 151.950 538.050 152.400 ;
        RECT 778.950 153.600 781.050 154.050 ;
        RECT 787.950 153.600 790.050 154.050 ;
        RECT 856.950 153.600 859.050 154.050 ;
        RECT 778.950 152.400 859.050 153.600 ;
        RECT 778.950 151.950 781.050 152.400 ;
        RECT 787.950 151.950 790.050 152.400 ;
        RECT 856.950 151.950 859.050 152.400 ;
        RECT 250.950 150.600 253.050 151.050 ;
        RECT 367.950 150.600 370.050 151.050 ;
        RECT 760.950 150.600 763.050 151.050 ;
        RECT 772.950 150.600 775.050 151.050 ;
        RECT 250.950 149.400 300.600 150.600 ;
        RECT 250.950 148.950 253.050 149.400 ;
        RECT 299.400 147.600 300.600 149.400 ;
        RECT 367.950 149.400 438.600 150.600 ;
        RECT 367.950 148.950 370.050 149.400 ;
        RECT 437.400 148.050 438.600 149.400 ;
        RECT 760.950 149.400 775.050 150.600 ;
        RECT 760.950 148.950 763.050 149.400 ;
        RECT 772.950 148.950 775.050 149.400 ;
        RECT 793.950 150.600 796.050 151.050 ;
        RECT 829.950 150.600 832.050 151.050 ;
        RECT 793.950 149.400 832.050 150.600 ;
        RECT 793.950 148.950 796.050 149.400 ;
        RECT 829.950 148.950 832.050 149.400 ;
        RECT 340.950 147.600 343.050 148.050 ;
        RECT 299.400 146.400 343.050 147.600 ;
        RECT 340.950 145.950 343.050 146.400 ;
        RECT 436.950 147.600 439.050 148.050 ;
        RECT 463.950 147.600 466.050 148.050 ;
        RECT 436.950 146.400 466.050 147.600 ;
        RECT 436.950 145.950 439.050 146.400 ;
        RECT 463.950 145.950 466.050 146.400 ;
        RECT 499.950 147.600 502.050 148.050 ;
        RECT 514.950 147.600 517.050 148.050 ;
        RECT 499.950 146.400 517.050 147.600 ;
        RECT 499.950 145.950 502.050 146.400 ;
        RECT 514.950 145.950 517.050 146.400 ;
        RECT 775.950 147.600 778.050 148.050 ;
        RECT 784.950 147.600 787.050 148.050 ;
        RECT 775.950 146.400 787.050 147.600 ;
        RECT 775.950 145.950 778.050 146.400 ;
        RECT 784.950 145.950 787.050 146.400 ;
        RECT 838.950 147.600 841.050 148.050 ;
        RECT 847.950 147.600 850.050 148.050 ;
        RECT 838.950 146.400 850.050 147.600 ;
        RECT 838.950 145.950 841.050 146.400 ;
        RECT 847.950 145.950 850.050 146.400 ;
        RECT 877.950 147.600 880.050 148.050 ;
        RECT 886.950 147.600 889.050 148.050 ;
        RECT 877.950 146.400 889.050 147.600 ;
        RECT 877.950 145.950 880.050 146.400 ;
        RECT 886.950 145.950 889.050 146.400 ;
        RECT 46.950 144.600 49.050 145.050 ;
        RECT 73.950 144.600 76.050 145.050 ;
        RECT 112.950 144.600 115.050 145.050 ;
        RECT 46.950 143.400 115.050 144.600 ;
        RECT 46.950 142.950 49.050 143.400 ;
        RECT 73.950 142.950 76.050 143.400 ;
        RECT 112.950 142.950 115.050 143.400 ;
        RECT 217.950 144.600 220.050 145.050 ;
        RECT 259.950 144.600 262.050 145.050 ;
        RECT 217.950 143.400 262.050 144.600 ;
        RECT 217.950 142.950 220.050 143.400 ;
        RECT 259.950 142.950 262.050 143.400 ;
        RECT 295.950 144.600 298.050 145.050 ;
        RECT 361.950 144.600 364.050 145.050 ;
        RECT 295.950 143.400 364.050 144.600 ;
        RECT 295.950 142.950 298.050 143.400 ;
        RECT 361.950 142.950 364.050 143.400 ;
        RECT 688.950 144.600 691.050 145.050 ;
        RECT 706.950 144.600 709.050 145.050 ;
        RECT 688.950 143.400 709.050 144.600 ;
        RECT 688.950 142.950 691.050 143.400 ;
        RECT 706.950 142.950 709.050 143.400 ;
        RECT 790.950 144.600 793.050 145.050 ;
        RECT 796.950 144.600 799.050 145.050 ;
        RECT 790.950 143.400 799.050 144.600 ;
        RECT 790.950 142.950 793.050 143.400 ;
        RECT 796.950 142.950 799.050 143.400 ;
        RECT 817.950 144.600 820.050 145.050 ;
        RECT 835.950 144.600 838.050 145.050 ;
        RECT 817.950 143.400 838.050 144.600 ;
        RECT 817.950 142.950 820.050 143.400 ;
        RECT 835.950 142.950 838.050 143.400 ;
        RECT 19.950 139.950 22.050 142.050 ;
        RECT 106.950 141.600 109.050 142.050 ;
        RECT 145.950 141.600 148.050 142.050 ;
        RECT 92.400 140.400 148.050 141.600 ;
        RECT 20.400 130.050 21.600 139.950 ;
        RECT 55.950 138.600 58.050 139.200 ;
        RECT 92.400 139.050 93.600 140.400 ;
        RECT 106.950 139.950 109.050 140.400 ;
        RECT 145.950 139.950 148.050 140.400 ;
        RECT 442.950 141.600 445.050 142.050 ;
        RECT 457.950 141.600 460.050 142.050 ;
        RECT 442.950 140.400 460.050 141.600 ;
        RECT 442.950 139.950 445.050 140.400 ;
        RECT 457.950 139.950 460.050 140.400 ;
        RECT 511.950 139.950 514.050 142.050 ;
        RECT 697.950 141.600 700.050 142.050 ;
        RECT 653.400 140.400 700.050 141.600 ;
        RECT 61.950 138.600 64.050 139.050 ;
        RECT 55.950 137.400 64.050 138.600 ;
        RECT 55.950 137.100 58.050 137.400 ;
        RECT 61.950 136.950 64.050 137.400 ;
        RECT 91.950 136.950 94.050 139.050 ;
        RECT 100.950 138.600 103.050 139.200 ;
        RECT 127.950 138.600 130.050 139.200 ;
        RECT 100.950 137.400 130.050 138.600 ;
        RECT 100.950 137.100 103.050 137.400 ;
        RECT 127.950 137.100 130.050 137.400 ;
        RECT 151.950 138.600 154.050 139.200 ;
        RECT 160.950 138.600 163.050 139.050 ;
        RECT 169.950 138.600 172.050 139.200 ;
        RECT 151.950 137.400 172.050 138.600 ;
        RECT 151.950 137.100 154.050 137.400 ;
        RECT 160.950 136.950 163.050 137.400 ;
        RECT 169.950 137.100 172.050 137.400 ;
        RECT 184.950 138.750 187.050 139.200 ;
        RECT 190.950 138.750 193.050 139.200 ;
        RECT 184.950 137.550 193.050 138.750 ;
        RECT 184.950 137.100 187.050 137.550 ;
        RECT 190.950 137.100 193.050 137.550 ;
        RECT 226.950 137.400 229.050 139.500 ;
        RECT 227.400 135.600 228.600 137.400 ;
        RECT 244.950 137.100 247.050 139.200 ;
        RECT 268.950 138.600 271.050 139.200 ;
        RECT 283.950 138.600 286.050 139.050 ;
        RECT 268.950 137.400 286.050 138.600 ;
        RECT 268.950 137.100 271.050 137.400 ;
        RECT 245.400 135.600 246.600 137.100 ;
        RECT 283.950 136.950 286.050 137.400 ;
        RECT 289.950 137.100 292.050 139.200 ;
        RECT 322.950 138.600 325.050 139.500 ;
        RECT 308.400 137.400 325.050 138.600 ;
        RECT 331.950 137.400 334.050 139.500 ;
        RECT 343.950 138.600 346.050 139.050 ;
        RECT 349.950 138.600 352.050 139.200 ;
        RECT 367.950 138.600 370.050 139.200 ;
        RECT 343.950 137.400 370.050 138.600 ;
        RECT 227.400 135.000 231.600 135.600 ;
        RECT 239.400 135.000 246.600 135.600 ;
        RECT 227.400 134.400 232.050 135.000 ;
        RECT 22.950 132.600 25.050 133.050 ;
        RECT 28.950 132.600 31.050 133.050 ;
        RECT 22.950 131.400 31.050 132.600 ;
        RECT 22.950 130.950 25.050 131.400 ;
        RECT 28.950 130.950 31.050 131.400 ;
        RECT 76.950 132.600 79.050 132.900 ;
        RECT 85.950 132.600 88.050 133.050 ;
        RECT 76.950 131.400 88.050 132.600 ;
        RECT 76.950 130.800 79.050 131.400 ;
        RECT 85.950 130.950 88.050 131.400 ;
        RECT 115.950 132.600 118.050 133.050 ;
        RECT 124.950 132.600 127.050 132.900 ;
        RECT 115.950 131.400 127.050 132.600 ;
        RECT 115.950 130.950 118.050 131.400 ;
        RECT 124.950 130.800 127.050 131.400 ;
        RECT 130.950 132.600 133.050 132.900 ;
        RECT 148.950 132.600 151.050 132.900 ;
        RECT 130.950 131.400 151.050 132.600 ;
        RECT 130.950 130.800 133.050 131.400 ;
        RECT 148.950 130.800 151.050 131.400 ;
        RECT 172.950 132.600 175.050 133.050 ;
        RECT 184.950 132.600 187.050 133.050 ;
        RECT 172.950 131.400 187.050 132.600 ;
        RECT 172.950 130.950 175.050 131.400 ;
        RECT 184.950 130.950 187.050 131.400 ;
        RECT 193.950 132.600 196.050 132.900 ;
        RECT 193.950 131.400 202.050 132.600 ;
        RECT 193.950 130.800 196.050 131.400 ;
        RECT 199.950 130.500 202.050 131.400 ;
        RECT 229.950 130.950 232.050 134.400 ;
        RECT 238.950 134.400 246.600 135.000 ;
        RECT 238.950 130.950 241.050 134.400 ;
        RECT 247.950 132.450 250.050 132.900 ;
        RECT 259.950 132.450 262.050 132.900 ;
        RECT 247.950 131.250 262.050 132.450 ;
        RECT 247.950 130.800 250.050 131.250 ;
        RECT 259.950 130.800 262.050 131.250 ;
        RECT 271.950 132.600 274.050 132.900 ;
        RECT 290.400 132.600 291.600 137.100 ;
        RECT 271.950 131.400 291.600 132.600 ;
        RECT 292.950 132.600 295.050 132.900 ;
        RECT 308.400 132.600 309.600 137.400 ;
        RECT 292.950 131.400 309.600 132.600 ;
        RECT 332.400 133.050 333.600 137.400 ;
        RECT 343.950 136.950 346.050 137.400 ;
        RECT 349.950 137.100 352.050 137.400 ;
        RECT 367.950 137.100 370.050 137.400 ;
        RECT 373.950 138.750 376.050 139.200 ;
        RECT 379.950 138.750 382.050 139.200 ;
        RECT 373.950 137.550 382.050 138.750 ;
        RECT 373.950 137.100 376.050 137.550 ;
        RECT 379.950 137.100 382.050 137.550 ;
        RECT 406.950 138.600 409.050 139.050 ;
        RECT 412.950 138.600 415.050 139.200 ;
        RECT 406.950 137.400 415.050 138.600 ;
        RECT 406.950 136.950 409.050 137.400 ;
        RECT 412.950 137.100 415.050 137.400 ;
        RECT 451.950 137.100 454.050 139.200 ;
        RECT 478.950 139.050 481.050 139.500 ;
        RECT 484.950 139.050 487.050 139.500 ;
        RECT 463.950 138.600 468.000 139.050 ;
        RECT 332.400 131.400 337.050 133.050 ;
        RECT 271.950 130.800 274.050 131.400 ;
        RECT 292.950 130.800 295.050 131.400 ;
        RECT 333.000 130.950 337.050 131.400 ;
        RECT 340.950 132.600 343.050 133.050 ;
        RECT 370.950 132.600 373.050 132.900 ;
        RECT 340.950 131.400 373.050 132.600 ;
        RECT 340.950 130.950 343.050 131.400 ;
        RECT 370.950 130.800 373.050 131.400 ;
        RECT 433.950 132.600 436.050 132.900 ;
        RECT 452.400 132.600 453.600 137.100 ;
        RECT 463.950 136.950 468.600 138.600 ;
        RECT 478.950 137.850 487.050 139.050 ;
        RECT 478.950 137.400 481.050 137.850 ;
        RECT 484.950 137.400 487.050 137.850 ;
        RECT 493.950 139.050 496.050 139.500 ;
        RECT 499.950 139.050 502.050 139.500 ;
        RECT 493.950 137.850 502.050 139.050 ;
        RECT 493.950 137.400 496.050 137.850 ;
        RECT 499.950 137.400 502.050 137.850 ;
        RECT 467.400 132.600 468.600 136.950 ;
        RECT 475.950 132.600 478.050 133.050 ;
        RECT 505.950 132.600 508.050 133.050 ;
        RECT 512.400 132.900 513.600 139.950 ;
        RECT 520.950 138.600 523.050 139.200 ;
        RECT 538.950 138.600 541.050 139.200 ;
        RECT 520.950 137.400 541.050 138.600 ;
        RECT 520.950 137.100 523.050 137.400 ;
        RECT 538.950 137.100 541.050 137.400 ;
        RECT 547.950 138.750 550.050 139.200 ;
        RECT 553.950 138.750 556.050 139.200 ;
        RECT 547.950 138.600 556.050 138.750 ;
        RECT 562.950 138.600 565.050 139.200 ;
        RECT 547.950 137.550 565.050 138.600 ;
        RECT 547.950 137.100 550.050 137.550 ;
        RECT 553.950 137.400 565.050 137.550 ;
        RECT 553.950 137.100 556.050 137.400 ;
        RECT 562.950 137.100 565.050 137.400 ;
        RECT 568.950 138.750 571.050 139.200 ;
        RECT 574.950 138.750 577.050 139.200 ;
        RECT 568.950 137.550 577.050 138.750 ;
        RECT 568.950 137.100 571.050 137.550 ;
        RECT 574.950 137.100 577.050 137.550 ;
        RECT 580.950 138.600 583.050 139.050 ;
        RECT 589.950 138.600 592.050 139.200 ;
        RECT 580.950 137.400 592.050 138.600 ;
        RECT 580.950 136.950 583.050 137.400 ;
        RECT 589.950 137.100 592.050 137.400 ;
        RECT 607.950 137.100 610.050 139.200 ;
        RECT 643.950 138.600 646.050 139.500 ;
        RECT 649.950 138.600 652.050 139.050 ;
        RECT 653.400 138.600 654.600 140.400 ;
        RECT 697.950 139.950 700.050 140.400 ;
        RECT 715.950 141.600 718.050 142.050 ;
        RECT 748.950 141.600 751.050 142.050 ;
        RECT 715.950 140.400 751.050 141.600 ;
        RECT 715.950 139.950 718.050 140.400 ;
        RECT 748.950 139.950 751.050 140.400 ;
        RECT 766.950 141.600 769.050 142.050 ;
        RECT 775.950 141.600 778.050 142.050 ;
        RECT 791.400 141.600 792.600 142.950 ;
        RECT 766.950 140.400 774.600 141.600 ;
        RECT 766.950 139.950 769.050 140.400 ;
        RECT 643.950 137.400 654.600 138.600 ;
        RECT 655.950 138.600 658.050 139.050 ;
        RECT 661.950 138.600 664.050 139.200 ;
        RECT 655.950 137.400 714.600 138.600 ;
        RECT 433.950 131.400 453.600 132.600 ;
        RECT 433.950 130.800 436.050 131.400 ;
        RECT 466.950 130.500 469.050 132.600 ;
        RECT 475.950 131.400 508.050 132.600 ;
        RECT 475.950 130.950 478.050 131.400 ;
        RECT 505.950 130.950 508.050 131.400 ;
        RECT 511.950 130.800 514.050 132.900 ;
        RECT 577.950 132.450 580.050 132.900 ;
        RECT 586.950 132.450 589.050 132.900 ;
        RECT 577.950 131.250 589.050 132.450 ;
        RECT 608.400 132.600 609.600 137.100 ;
        RECT 628.950 135.600 631.050 136.050 ;
        RECT 644.400 135.600 645.600 137.400 ;
        RECT 649.950 136.950 652.050 137.400 ;
        RECT 655.950 136.950 658.050 137.400 ;
        RECT 661.950 137.100 664.050 137.400 ;
        RECT 628.950 134.400 645.600 135.600 ;
        RECT 628.950 133.950 631.050 134.400 ;
        RECT 613.950 132.600 616.050 133.050 ;
        RECT 713.400 132.900 714.600 137.400 ;
        RECT 715.950 137.100 718.050 139.200 ;
        RECT 721.950 137.100 724.050 139.200 ;
        RECT 608.400 131.400 616.050 132.600 ;
        RECT 577.950 130.800 580.050 131.250 ;
        RECT 586.950 130.800 589.050 131.250 ;
        RECT 613.950 130.950 616.050 131.400 ;
        RECT 712.950 130.800 715.050 132.900 ;
        RECT 716.400 130.050 717.600 137.100 ;
        RECT 722.400 132.600 723.600 137.100 ;
        RECT 736.950 136.950 739.050 139.050 ;
        RECT 742.950 137.100 745.050 139.200 ;
        RECT 727.950 132.600 730.050 133.050 ;
        RECT 722.400 131.400 730.050 132.600 ;
        RECT 727.950 130.950 730.050 131.400 ;
        RECT 19.950 127.950 22.050 130.050 ;
        RECT 49.950 129.600 52.050 130.050 ;
        RECT 55.950 129.600 58.050 130.050 ;
        RECT 49.950 128.400 58.050 129.600 ;
        RECT 49.950 127.950 52.050 128.400 ;
        RECT 55.950 127.950 58.050 128.400 ;
        RECT 91.950 129.600 94.050 130.050 ;
        RECT 97.950 129.600 100.050 130.050 ;
        RECT 91.950 128.400 100.050 129.600 ;
        RECT 91.950 127.950 94.050 128.400 ;
        RECT 97.950 127.950 100.050 128.400 ;
        RECT 241.950 129.600 244.050 130.050 ;
        RECT 253.950 129.600 256.050 130.050 ;
        RECT 286.950 129.600 289.050 130.050 ;
        RECT 241.950 128.400 289.050 129.600 ;
        RECT 241.950 127.950 244.050 128.400 ;
        RECT 253.950 127.950 256.050 128.400 ;
        RECT 286.950 127.950 289.050 128.400 ;
        RECT 520.950 129.600 523.050 130.050 ;
        RECT 544.950 129.600 547.050 130.050 ;
        RECT 565.950 129.600 568.050 130.050 ;
        RECT 580.950 129.600 583.050 130.050 ;
        RECT 520.950 128.400 583.050 129.600 ;
        RECT 520.950 127.950 523.050 128.400 ;
        RECT 544.950 127.950 547.050 128.400 ;
        RECT 565.950 127.950 568.050 128.400 ;
        RECT 580.950 127.950 583.050 128.400 ;
        RECT 610.950 129.600 613.050 130.050 ;
        RECT 616.950 129.600 619.050 130.050 ;
        RECT 610.950 128.400 619.050 129.600 ;
        RECT 610.950 127.950 613.050 128.400 ;
        RECT 616.950 127.950 619.050 128.400 ;
        RECT 634.950 129.600 637.050 130.050 ;
        RECT 652.950 129.600 655.050 130.050 ;
        RECT 634.950 128.400 655.050 129.600 ;
        RECT 634.950 127.950 637.050 128.400 ;
        RECT 652.950 127.950 655.050 128.400 ;
        RECT 679.950 129.600 682.050 130.050 ;
        RECT 688.950 129.600 691.050 130.050 ;
        RECT 679.950 128.400 691.050 129.600 ;
        RECT 679.950 127.950 682.050 128.400 ;
        RECT 688.950 127.950 691.050 128.400 ;
        RECT 715.950 127.950 718.050 130.050 ;
        RECT 737.400 129.900 738.600 136.950 ;
        RECT 743.400 132.600 744.600 137.100 ;
        RECT 773.400 132.900 774.600 140.400 ;
        RECT 775.950 140.400 792.600 141.600 ;
        RECT 823.950 141.600 826.050 142.050 ;
        RECT 832.950 141.600 835.050 142.050 ;
        RECT 865.950 141.600 868.050 142.050 ;
        RECT 823.950 140.400 835.050 141.600 ;
        RECT 775.950 139.950 778.050 140.400 ;
        RECT 823.950 139.950 826.050 140.400 ;
        RECT 832.950 139.950 835.050 140.400 ;
        RECT 845.400 140.400 868.050 141.600 ;
        RECT 778.950 138.600 781.050 139.050 ;
        RECT 799.950 138.600 802.050 139.050 ;
        RECT 808.950 138.600 811.050 139.050 ;
        RECT 778.950 137.400 789.600 138.600 ;
        RECT 778.950 136.950 781.050 137.400 ;
        RECT 788.400 132.900 789.600 137.400 ;
        RECT 799.950 137.400 811.050 138.600 ;
        RECT 799.950 136.950 802.050 137.400 ;
        RECT 808.950 136.950 811.050 137.400 ;
        RECT 820.950 136.950 823.050 139.050 ;
        RECT 821.400 133.050 822.600 136.950 ;
        RECT 766.950 132.600 769.050 132.900 ;
        RECT 743.400 131.400 769.050 132.600 ;
        RECT 766.950 130.800 769.050 131.400 ;
        RECT 772.950 130.800 775.050 132.900 ;
        RECT 787.950 130.800 790.050 132.900 ;
        RECT 820.950 130.950 823.050 133.050 ;
        RECT 826.950 132.600 829.050 133.050 ;
        RECT 835.950 132.600 838.050 132.900 ;
        RECT 826.950 131.400 838.050 132.600 ;
        RECT 826.950 130.950 829.050 131.400 ;
        RECT 835.950 130.800 838.050 131.400 ;
        RECT 736.800 127.800 738.900 129.900 ;
        RECT 739.950 129.600 742.050 130.050 ;
        RECT 817.950 129.600 820.050 130.050 ;
        RECT 845.400 129.900 846.600 140.400 ;
        RECT 865.950 139.950 868.050 140.400 ;
        RECT 871.950 137.100 874.050 139.200 ;
        RECT 850.950 132.450 853.050 132.900 ;
        RECT 859.950 132.450 862.050 132.900 ;
        RECT 850.950 131.250 862.050 132.450 ;
        RECT 850.950 130.800 853.050 131.250 ;
        RECT 859.950 130.800 862.050 131.250 ;
        RECT 739.950 128.400 820.050 129.600 ;
        RECT 739.950 127.950 742.050 128.400 ;
        RECT 817.950 127.950 820.050 128.400 ;
        RECT 844.950 127.800 847.050 129.900 ;
        RECT 872.400 129.600 873.600 137.100 ;
        RECT 883.950 136.950 886.050 139.050 ;
        RECT 884.400 130.050 885.600 136.950 ;
        RECT 877.800 129.600 879.900 130.050 ;
        RECT 872.400 128.400 879.900 129.600 ;
        RECT 877.800 127.950 879.900 128.400 ;
        RECT 880.950 128.400 885.600 130.050 ;
        RECT 880.950 127.950 885.000 128.400 ;
        RECT 175.950 126.600 178.050 127.050 ;
        RECT 232.950 126.600 235.050 127.050 ;
        RECT 175.950 125.400 235.050 126.600 ;
        RECT 175.950 124.950 178.050 125.400 ;
        RECT 232.950 124.950 235.050 125.400 ;
        RECT 283.950 126.600 286.050 127.050 ;
        RECT 298.950 126.600 301.050 127.050 ;
        RECT 283.950 125.400 301.050 126.600 ;
        RECT 283.950 124.950 286.050 125.400 ;
        RECT 298.950 124.950 301.050 125.400 ;
        RECT 355.950 126.600 358.050 127.050 ;
        RECT 400.950 126.600 403.050 127.050 ;
        RECT 355.950 125.400 403.050 126.600 ;
        RECT 355.950 124.950 358.050 125.400 ;
        RECT 400.950 124.950 403.050 125.400 ;
        RECT 454.950 126.600 457.050 127.050 ;
        RECT 478.950 126.600 481.050 127.050 ;
        RECT 454.950 125.400 481.050 126.600 ;
        RECT 454.950 124.950 457.050 125.400 ;
        RECT 478.950 124.950 481.050 125.400 ;
        RECT 523.950 126.600 526.050 127.050 ;
        RECT 541.950 126.600 544.050 127.050 ;
        RECT 523.950 125.400 544.050 126.600 ;
        RECT 523.950 124.950 526.050 125.400 ;
        RECT 541.950 124.950 544.050 125.400 ;
        RECT 706.950 126.600 709.050 127.050 ;
        RECT 718.950 126.600 721.050 127.050 ;
        RECT 706.950 125.400 721.050 126.600 ;
        RECT 706.950 124.950 709.050 125.400 ;
        RECT 718.950 124.950 721.050 125.400 ;
        RECT 757.950 126.600 760.050 127.050 ;
        RECT 787.950 126.600 790.050 127.050 ;
        RECT 757.950 125.400 790.050 126.600 ;
        RECT 757.950 124.950 760.050 125.400 ;
        RECT 787.950 124.950 790.050 125.400 ;
        RECT 805.950 126.600 808.050 127.050 ;
        RECT 838.950 126.600 841.050 127.050 ;
        RECT 805.950 125.400 841.050 126.600 ;
        RECT 805.950 124.950 808.050 125.400 ;
        RECT 838.950 124.950 841.050 125.400 ;
        RECT 97.950 123.600 100.050 124.050 ;
        RECT 142.950 123.600 145.050 124.050 ;
        RECT 97.950 122.400 145.050 123.600 ;
        RECT 97.950 121.950 100.050 122.400 ;
        RECT 142.950 121.950 145.050 122.400 ;
        RECT 442.950 123.600 445.050 124.050 ;
        RECT 475.950 123.600 478.050 124.050 ;
        RECT 442.950 122.400 478.050 123.600 ;
        RECT 442.950 121.950 445.050 122.400 ;
        RECT 475.950 121.950 478.050 122.400 ;
        RECT 703.950 123.600 706.050 124.050 ;
        RECT 724.800 123.600 726.900 124.050 ;
        RECT 703.950 122.400 726.900 123.600 ;
        RECT 703.950 121.950 706.050 122.400 ;
        RECT 724.800 121.950 726.900 122.400 ;
        RECT 727.950 123.600 730.050 124.050 ;
        RECT 745.950 123.600 748.050 124.050 ;
        RECT 727.950 122.400 748.050 123.600 ;
        RECT 727.950 121.950 730.050 122.400 ;
        RECT 745.950 121.950 748.050 122.400 ;
        RECT 841.950 123.600 844.050 124.050 ;
        RECT 868.950 123.600 871.050 124.050 ;
        RECT 841.950 122.400 871.050 123.600 ;
        RECT 841.950 121.950 844.050 122.400 ;
        RECT 868.950 121.950 871.050 122.400 ;
        RECT 874.950 123.600 877.050 124.050 ;
        RECT 895.950 123.600 898.050 124.050 ;
        RECT 874.950 122.400 898.050 123.600 ;
        RECT 874.950 121.950 877.050 122.400 ;
        RECT 895.950 121.950 898.050 122.400 ;
        RECT 172.950 120.600 175.050 121.050 ;
        RECT 238.950 120.600 241.050 121.050 ;
        RECT 172.950 119.400 241.050 120.600 ;
        RECT 172.950 118.950 175.050 119.400 ;
        RECT 238.950 118.950 241.050 119.400 ;
        RECT 280.950 120.600 283.050 121.050 ;
        RECT 301.950 120.600 304.050 121.050 ;
        RECT 280.950 119.400 304.050 120.600 ;
        RECT 280.950 118.950 283.050 119.400 ;
        RECT 301.950 118.950 304.050 119.400 ;
        RECT 307.950 120.600 310.050 121.050 ;
        RECT 313.950 120.600 316.050 121.050 ;
        RECT 340.950 120.600 343.050 121.050 ;
        RECT 307.950 119.400 343.050 120.600 ;
        RECT 307.950 118.950 310.050 119.400 ;
        RECT 313.950 118.950 316.050 119.400 ;
        RECT 340.950 118.950 343.050 119.400 ;
        RECT 487.950 120.600 490.050 121.050 ;
        RECT 499.950 120.600 502.050 121.050 ;
        RECT 628.950 120.600 631.050 121.050 ;
        RECT 487.950 119.400 631.050 120.600 ;
        RECT 487.950 118.950 490.050 119.400 ;
        RECT 499.950 118.950 502.050 119.400 ;
        RECT 628.950 118.950 631.050 119.400 ;
        RECT 754.950 120.600 757.050 121.050 ;
        RECT 766.950 120.600 769.050 121.050 ;
        RECT 754.950 119.400 769.050 120.600 ;
        RECT 754.950 118.950 757.050 119.400 ;
        RECT 766.950 118.950 769.050 119.400 ;
        RECT 781.950 120.600 784.050 121.050 ;
        RECT 835.950 120.600 838.050 121.050 ;
        RECT 781.950 119.400 838.050 120.600 ;
        RECT 781.950 118.950 784.050 119.400 ;
        RECT 835.950 118.950 838.050 119.400 ;
        RECT 286.950 117.600 289.050 118.050 ;
        RECT 316.950 117.600 319.050 118.050 ;
        RECT 343.950 117.600 346.050 118.050 ;
        RECT 286.950 116.400 346.050 117.600 ;
        RECT 286.950 115.950 289.050 116.400 ;
        RECT 316.950 115.950 319.050 116.400 ;
        RECT 343.950 115.950 346.050 116.400 ;
        RECT 406.950 117.600 409.050 118.050 ;
        RECT 415.950 117.600 418.050 118.050 ;
        RECT 406.950 116.400 418.050 117.600 ;
        RECT 406.950 115.950 409.050 116.400 ;
        RECT 415.950 115.950 418.050 116.400 ;
        RECT 631.950 117.600 634.050 118.050 ;
        RECT 655.950 117.600 658.050 118.050 ;
        RECT 631.950 116.400 658.050 117.600 ;
        RECT 631.950 115.950 634.050 116.400 ;
        RECT 655.950 115.950 658.050 116.400 ;
        RECT 670.950 117.600 673.050 118.050 ;
        RECT 682.950 117.600 685.050 118.050 ;
        RECT 670.950 116.400 685.050 117.600 ;
        RECT 670.950 115.950 673.050 116.400 ;
        RECT 682.950 115.950 685.050 116.400 ;
        RECT 805.950 117.600 808.050 118.050 ;
        RECT 841.950 117.600 844.050 118.050 ;
        RECT 805.950 116.400 844.050 117.600 ;
        RECT 805.950 115.950 808.050 116.400 ;
        RECT 841.950 115.950 844.050 116.400 ;
        RECT 847.950 117.600 850.050 118.050 ;
        RECT 874.950 117.600 877.050 118.050 ;
        RECT 847.950 116.400 877.050 117.600 ;
        RECT 847.950 115.950 850.050 116.400 ;
        RECT 874.950 115.950 877.050 116.400 ;
        RECT 85.950 114.600 88.050 115.050 ;
        RECT 97.950 114.600 100.050 115.050 ;
        RECT 106.950 114.600 109.050 115.050 ;
        RECT 85.950 113.400 109.050 114.600 ;
        RECT 85.950 112.950 88.050 113.400 ;
        RECT 97.950 112.950 100.050 113.400 ;
        RECT 106.950 112.950 109.050 113.400 ;
        RECT 277.950 114.600 280.050 115.050 ;
        RECT 490.950 114.600 493.050 115.050 ;
        RECT 277.950 113.400 493.050 114.600 ;
        RECT 277.950 112.950 280.050 113.400 ;
        RECT 490.950 112.950 493.050 113.400 ;
        RECT 496.950 114.600 499.050 115.050 ;
        RECT 586.950 114.600 589.050 115.050 ;
        RECT 496.950 113.400 589.050 114.600 ;
        RECT 496.950 112.950 499.050 113.400 ;
        RECT 586.950 112.950 589.050 113.400 ;
        RECT 595.950 114.600 598.050 115.050 ;
        RECT 700.950 114.600 703.050 115.050 ;
        RECT 595.950 113.400 703.050 114.600 ;
        RECT 595.950 112.950 598.050 113.400 ;
        RECT 700.950 112.950 703.050 113.400 ;
        RECT 763.950 114.600 766.050 115.050 ;
        RECT 796.950 114.600 799.050 115.050 ;
        RECT 763.950 113.400 799.050 114.600 ;
        RECT 763.950 112.950 766.050 113.400 ;
        RECT 796.950 112.950 799.050 113.400 ;
        RECT 802.950 114.600 805.050 115.050 ;
        RECT 883.950 114.600 886.050 115.050 ;
        RECT 802.950 113.400 886.050 114.600 ;
        RECT 802.950 112.950 805.050 113.400 ;
        RECT 883.950 112.950 886.050 113.400 ;
        RECT 43.950 111.600 46.050 112.050 ;
        RECT 76.950 111.600 79.050 112.050 ;
        RECT 43.950 110.400 79.050 111.600 ;
        RECT 43.950 109.950 46.050 110.400 ;
        RECT 76.950 109.950 79.050 110.400 ;
        RECT 142.950 111.600 145.050 112.050 ;
        RECT 157.950 111.600 160.050 112.050 ;
        RECT 142.950 110.400 160.050 111.600 ;
        RECT 142.950 109.950 145.050 110.400 ;
        RECT 157.950 109.950 160.050 110.400 ;
        RECT 331.950 111.600 334.050 112.050 ;
        RECT 346.950 111.600 349.050 112.050 ;
        RECT 331.950 110.400 349.050 111.600 ;
        RECT 331.950 109.950 334.050 110.400 ;
        RECT 346.950 109.950 349.050 110.400 ;
        RECT 391.950 111.600 394.050 112.050 ;
        RECT 427.950 111.600 430.050 112.050 ;
        RECT 391.950 110.400 430.050 111.600 ;
        RECT 391.950 109.950 394.050 110.400 ;
        RECT 427.950 109.950 430.050 110.400 ;
        RECT 457.950 111.600 460.050 112.050 ;
        RECT 493.950 111.600 496.050 112.050 ;
        RECT 589.950 111.600 592.050 111.900 ;
        RECT 457.950 110.400 592.050 111.600 ;
        RECT 457.950 109.950 460.050 110.400 ;
        RECT 493.950 109.950 496.050 110.400 ;
        RECT 589.950 109.800 592.050 110.400 ;
        RECT 649.950 111.600 652.050 112.050 ;
        RECT 691.950 111.600 694.050 112.050 ;
        RECT 764.400 111.600 765.600 112.950 ;
        RECT 649.950 110.400 694.050 111.600 ;
        RECT 649.950 109.950 652.050 110.400 ;
        RECT 691.950 109.950 694.050 110.400 ;
        RECT 755.400 110.400 765.600 111.600 ;
        RECT 820.950 111.600 823.050 112.050 ;
        RECT 841.950 111.600 844.050 112.050 ;
        RECT 820.950 110.400 844.050 111.600 ;
        RECT 343.950 106.950 346.050 109.050 ;
        RECT 370.950 108.600 373.050 109.050 ;
        RECT 421.950 108.600 424.050 109.050 ;
        RECT 433.950 108.600 436.050 109.050 ;
        RECT 370.950 107.400 436.050 108.600 ;
        RECT 370.950 106.950 373.050 107.400 ;
        RECT 421.950 106.950 424.050 107.400 ;
        RECT 433.950 106.950 436.050 107.400 ;
        RECT 580.950 108.600 585.000 109.050 ;
        RECT 628.950 108.600 631.050 109.050 ;
        RECT 580.950 106.950 585.600 108.600 ;
        RECT 49.950 104.100 52.050 106.200 ;
        RECT 67.950 105.600 70.050 106.200 ;
        RECT 67.950 104.400 75.600 105.600 ;
        RECT 67.950 104.100 70.050 104.400 ;
        RECT 31.950 99.600 34.050 100.050 ;
        RECT 46.950 99.600 49.050 99.900 ;
        RECT 31.950 98.400 49.050 99.600 ;
        RECT 50.400 99.600 51.600 104.100 ;
        RECT 74.400 100.050 75.600 104.400 ;
        RECT 91.950 104.100 94.050 106.200 ;
        RECT 103.950 105.750 106.050 106.200 ;
        RECT 115.800 105.750 117.900 106.200 ;
        RECT 103.950 104.550 117.900 105.750 ;
        RECT 103.950 104.100 106.050 104.550 ;
        RECT 115.800 104.100 117.900 104.550 ;
        RECT 118.950 105.750 121.050 106.200 ;
        RECT 124.950 105.750 127.050 106.200 ;
        RECT 118.950 104.550 127.050 105.750 ;
        RECT 118.950 104.100 121.050 104.550 ;
        RECT 124.950 104.100 127.050 104.550 ;
        RECT 130.950 104.100 133.050 106.200 ;
        RECT 166.950 104.100 169.050 106.200 ;
        RECT 187.950 105.600 190.050 106.200 ;
        RECT 214.950 105.600 217.050 106.200 ;
        RECT 220.950 105.600 223.050 106.500 ;
        RECT 187.950 104.400 223.050 105.600 ;
        RECT 232.950 105.750 235.050 106.200 ;
        RECT 262.950 105.750 265.050 106.200 ;
        RECT 232.950 104.550 265.050 105.750 ;
        RECT 187.950 104.100 190.050 104.400 ;
        RECT 214.950 104.100 217.050 104.400 ;
        RECT 232.950 104.100 235.050 104.550 ;
        RECT 262.950 104.100 265.050 104.550 ;
        RECT 268.950 105.600 271.050 106.200 ;
        RECT 331.950 105.600 334.050 106.050 ;
        RECT 268.950 104.400 276.600 105.600 ;
        RECT 268.950 104.100 271.050 104.400 ;
        RECT 61.950 99.600 64.050 100.050 ;
        RECT 50.400 98.400 64.050 99.600 ;
        RECT 31.950 97.950 34.050 98.400 ;
        RECT 46.950 97.800 49.050 98.400 ;
        RECT 61.950 97.950 64.050 98.400 ;
        RECT 73.950 97.950 76.050 100.050 ;
        RECT 92.400 99.600 93.600 104.100 ;
        RECT 106.950 99.600 109.050 99.900 ;
        RECT 92.400 98.400 109.050 99.600 ;
        RECT 106.950 97.800 109.050 98.400 ;
        RECT 115.950 99.600 118.050 100.050 ;
        RECT 127.950 99.600 130.050 99.900 ;
        RECT 115.950 98.400 130.050 99.600 ;
        RECT 131.400 99.600 132.600 104.100 ;
        RECT 167.400 102.600 168.600 104.100 ;
        RECT 167.400 101.400 195.600 102.600 ;
        RECT 190.950 99.600 193.050 99.900 ;
        RECT 131.400 98.400 193.050 99.600 ;
        RECT 194.400 99.600 195.600 101.400 ;
        RECT 275.400 100.050 276.600 104.400 ;
        RECT 317.400 104.400 334.050 105.600 ;
        RECT 211.950 99.600 214.050 99.900 ;
        RECT 232.950 99.600 235.050 100.050 ;
        RECT 194.400 98.400 235.050 99.600 ;
        RECT 115.950 97.950 118.050 98.400 ;
        RECT 127.950 97.800 130.050 98.400 ;
        RECT 190.950 97.800 193.050 98.400 ;
        RECT 211.950 97.800 214.050 98.400 ;
        RECT 232.950 97.950 235.050 98.400 ;
        RECT 253.950 99.450 256.050 99.900 ;
        RECT 265.950 99.450 268.050 99.900 ;
        RECT 253.950 98.250 268.050 99.450 ;
        RECT 253.950 97.800 256.050 98.250 ;
        RECT 265.950 97.800 268.050 98.250 ;
        RECT 274.950 97.950 277.050 100.050 ;
        RECT 289.950 99.450 292.050 99.900 ;
        RECT 307.950 99.450 310.050 99.900 ;
        RECT 317.400 99.600 318.600 104.400 ;
        RECT 331.950 103.950 334.050 104.400 ;
        RECT 328.950 99.600 331.050 100.050 ;
        RECT 334.950 99.600 337.050 100.050 ;
        RECT 344.400 99.900 345.600 106.950 ;
        RECT 352.950 105.750 355.050 106.200 ;
        RECT 358.950 105.750 361.050 106.200 ;
        RECT 352.950 104.550 361.050 105.750 ;
        RECT 352.950 104.100 355.050 104.550 ;
        RECT 358.950 104.100 361.050 104.550 ;
        RECT 364.950 105.750 367.050 106.200 ;
        RECT 370.950 105.750 373.050 106.200 ;
        RECT 364.950 104.550 373.050 105.750 ;
        RECT 364.950 104.100 367.050 104.550 ;
        RECT 370.950 104.100 373.050 104.550 ;
        RECT 376.950 105.600 379.050 106.200 ;
        RECT 382.950 105.600 385.050 106.500 ;
        RECT 376.950 104.400 385.050 105.600 ;
        RECT 394.950 105.600 397.050 106.050 ;
        RECT 421.950 105.600 424.050 105.900 ;
        RECT 394.950 104.400 424.050 105.600 ;
        RECT 376.950 104.100 379.050 104.400 ;
        RECT 394.950 103.950 397.050 104.400 ;
        RECT 421.950 103.800 424.050 104.400 ;
        RECT 442.950 105.750 445.050 106.200 ;
        RECT 451.950 105.750 454.050 106.200 ;
        RECT 442.950 104.550 454.050 105.750 ;
        RECT 442.950 104.100 445.050 104.550 ;
        RECT 451.950 104.100 454.050 104.550 ;
        RECT 481.950 105.600 484.050 106.200 ;
        RECT 514.950 105.600 517.050 106.200 ;
        RECT 532.950 105.600 535.050 106.200 ;
        RECT 481.950 104.400 535.050 105.600 ;
        RECT 481.950 104.100 484.050 104.400 ;
        RECT 514.950 104.100 517.050 104.400 ;
        RECT 532.950 104.100 535.050 104.400 ;
        RECT 538.950 105.600 541.050 106.200 ;
        RECT 553.950 105.600 556.050 106.050 ;
        RECT 538.950 104.400 556.050 105.600 ;
        RECT 538.950 104.100 541.050 104.400 ;
        RECT 289.950 98.250 310.050 99.450 ;
        RECT 289.950 97.800 292.050 98.250 ;
        RECT 307.950 97.800 310.050 98.250 ;
        RECT 316.950 97.500 319.050 99.600 ;
        RECT 328.950 98.400 337.050 99.600 ;
        RECT 328.950 97.950 331.050 98.400 ;
        RECT 334.950 97.950 337.050 98.400 ;
        RECT 343.950 97.800 346.050 99.900 ;
        RECT 373.950 99.600 376.050 99.900 ;
        RECT 394.950 99.600 397.050 100.050 ;
        RECT 373.950 98.400 397.050 99.600 ;
        RECT 373.950 97.800 376.050 98.400 ;
        RECT 394.950 97.950 397.050 98.400 ;
        RECT 409.950 99.150 412.050 99.600 ;
        RECT 415.950 99.150 418.050 99.600 ;
        RECT 409.950 97.950 418.050 99.150 ;
        RECT 409.950 97.500 412.050 97.950 ;
        RECT 415.950 97.500 418.050 97.950 ;
        RECT 421.950 99.450 424.050 99.900 ;
        RECT 430.950 99.450 433.050 99.900 ;
        RECT 421.950 98.250 433.050 99.450 ;
        RECT 421.950 97.800 424.050 98.250 ;
        RECT 430.950 97.800 433.050 98.250 ;
        RECT 454.950 99.600 457.050 99.900 ;
        RECT 463.950 99.600 466.050 100.050 ;
        RECT 454.950 98.400 466.050 99.600 ;
        RECT 482.400 99.600 483.600 104.100 ;
        RECT 553.950 103.950 556.050 104.400 ;
        RECT 577.950 103.950 580.050 106.050 ;
        RECT 584.400 105.600 585.600 106.950 ;
        RECT 602.400 107.400 631.050 108.600 ;
        RECT 598.950 105.600 601.050 106.050 ;
        RECT 584.400 104.400 601.050 105.600 ;
        RECT 598.950 103.950 601.050 104.400 ;
        RECT 578.400 100.050 579.600 103.950 ;
        RECT 496.950 99.600 499.050 99.900 ;
        RECT 482.400 98.400 499.050 99.600 ;
        RECT 454.950 97.800 457.050 98.400 ;
        RECT 463.950 97.950 466.050 98.400 ;
        RECT 496.950 97.800 499.050 98.400 ;
        RECT 541.950 99.600 544.050 99.900 ;
        RECT 559.950 99.600 562.050 99.900 ;
        RECT 574.800 99.600 576.900 99.900 ;
        RECT 541.950 98.400 576.900 99.600 ;
        RECT 541.950 97.800 544.050 98.400 ;
        RECT 559.950 97.800 562.050 98.400 ;
        RECT 574.800 97.800 576.900 98.400 ;
        RECT 577.950 97.950 580.050 100.050 ;
        RECT 583.950 99.600 586.050 99.900 ;
        RECT 589.950 99.600 592.050 100.050 ;
        RECT 602.400 99.900 603.600 107.400 ;
        RECT 628.950 106.950 631.050 107.400 ;
        RECT 616.950 105.750 619.050 106.200 ;
        RECT 622.950 105.750 625.050 106.200 ;
        RECT 616.950 104.550 625.050 105.750 ;
        RECT 616.950 104.100 619.050 104.550 ;
        RECT 622.950 104.100 625.050 104.550 ;
        RECT 649.950 105.600 652.050 106.200 ;
        RECT 655.950 105.600 658.050 106.500 ;
        RECT 649.950 104.400 658.050 105.600 ;
        RECT 670.950 105.600 675.000 106.050 ;
        RECT 706.950 105.600 709.050 106.200 ;
        RECT 724.950 105.600 727.050 106.200 ;
        RECT 755.400 105.600 756.600 110.400 ;
        RECT 820.950 109.950 823.050 110.400 ;
        RECT 841.950 109.950 844.050 110.400 ;
        RECT 769.950 108.600 772.050 109.050 ;
        RECT 781.950 108.600 784.050 109.050 ;
        RECT 769.950 107.400 784.050 108.600 ;
        RECT 769.950 106.950 772.050 107.400 ;
        RECT 781.950 106.950 784.050 107.400 ;
        RECT 856.950 108.600 859.050 109.050 ;
        RECT 865.950 108.600 868.050 109.050 ;
        RECT 886.950 108.600 889.050 109.050 ;
        RECT 856.950 107.400 868.050 108.600 ;
        RECT 856.950 106.950 859.050 107.400 ;
        RECT 865.950 106.950 868.050 107.400 ;
        RECT 872.400 107.400 889.050 108.600 ;
        RECT 649.950 104.100 652.050 104.400 ;
        RECT 653.400 100.050 654.600 104.400 ;
        RECT 670.950 103.950 675.600 105.600 ;
        RECT 706.950 104.400 727.050 105.600 ;
        RECT 743.400 105.000 756.600 105.600 ;
        RECT 706.950 104.100 709.050 104.400 ;
        RECT 724.950 104.100 727.050 104.400 ;
        RECT 742.950 104.400 756.600 105.000 ;
        RECT 781.950 105.600 784.050 106.200 ;
        RECT 805.950 105.600 808.050 106.200 ;
        RECT 823.950 105.600 826.050 106.200 ;
        RECT 781.950 104.400 798.600 105.600 ;
        RECT 583.950 98.400 592.050 99.600 ;
        RECT 583.950 97.800 586.050 98.400 ;
        RECT 589.950 97.950 592.050 98.400 ;
        RECT 601.950 97.800 604.050 99.900 ;
        RECT 607.950 99.600 610.050 99.900 ;
        RECT 616.950 99.600 619.050 100.050 ;
        RECT 607.950 98.400 619.050 99.600 ;
        RECT 607.950 97.800 610.050 98.400 ;
        RECT 616.950 97.950 619.050 98.400 ;
        RECT 652.950 97.950 655.050 100.050 ;
        RECT 674.400 99.600 675.600 103.950 ;
        RECT 742.950 100.800 745.050 104.400 ;
        RECT 781.950 104.100 784.050 104.400 ;
        RECT 797.400 99.900 798.600 104.400 ;
        RECT 805.950 104.400 826.050 105.600 ;
        RECT 805.950 104.100 808.050 104.400 ;
        RECT 823.950 104.100 826.050 104.400 ;
        RECT 829.950 103.950 832.050 106.050 ;
        RECT 838.950 103.950 841.050 106.050 ;
        RECT 830.400 100.050 831.600 103.950 ;
        RECT 839.400 100.050 840.600 103.950 ;
        RECT 872.400 100.050 873.600 107.400 ;
        RECT 886.950 106.950 889.050 107.400 ;
        RECT 673.950 97.500 676.050 99.600 ;
        RECT 682.950 99.150 685.050 99.600 ;
        RECT 691.950 99.150 694.050 99.600 ;
        RECT 682.950 97.950 694.050 99.150 ;
        RECT 682.950 97.500 685.050 97.950 ;
        RECT 691.950 97.500 694.050 97.950 ;
        RECT 727.950 99.450 730.050 99.900 ;
        RECT 736.950 99.450 739.050 99.900 ;
        RECT 727.950 98.250 739.050 99.450 ;
        RECT 727.950 97.800 730.050 98.250 ;
        RECT 736.950 97.800 739.050 98.250 ;
        RECT 766.950 99.450 769.050 99.900 ;
        RECT 772.950 99.450 775.050 99.900 ;
        RECT 766.950 98.250 775.050 99.450 ;
        RECT 766.950 97.800 769.050 98.250 ;
        RECT 772.950 97.800 775.050 98.250 ;
        RECT 796.950 97.800 799.050 99.900 ;
        RECT 817.950 99.600 820.050 100.050 ;
        RECT 826.950 99.600 829.050 99.900 ;
        RECT 817.950 98.400 829.050 99.600 ;
        RECT 830.400 98.400 835.050 100.050 ;
        RECT 817.950 97.950 820.050 98.400 ;
        RECT 826.950 97.800 829.050 98.400 ;
        RECT 831.000 97.950 835.050 98.400 ;
        RECT 838.950 97.950 841.050 100.050 ;
        RECT 850.950 99.600 853.050 100.050 ;
        RECT 865.950 99.600 868.050 99.900 ;
        RECT 850.950 98.400 868.050 99.600 ;
        RECT 850.950 97.950 853.050 98.400 ;
        RECT 865.950 97.800 868.050 98.400 ;
        RECT 871.950 97.950 874.050 100.050 ;
        RECT 877.950 99.600 880.050 100.050 ;
        RECT 886.950 99.600 889.050 99.900 ;
        RECT 877.950 98.400 889.050 99.600 ;
        RECT 877.950 97.950 880.050 98.400 ;
        RECT 886.950 97.800 889.050 98.400 ;
        RECT 76.950 96.600 79.050 97.050 ;
        RECT 88.950 96.600 91.050 97.050 ;
        RECT 76.950 95.400 91.050 96.600 ;
        RECT 76.950 94.950 79.050 95.400 ;
        RECT 88.950 94.950 91.050 95.400 ;
        RECT 118.950 96.600 121.050 97.050 ;
        RECT 169.950 96.600 172.050 97.050 ;
        RECT 118.950 95.400 172.050 96.600 ;
        RECT 118.950 94.950 121.050 95.400 ;
        RECT 169.950 94.950 172.050 95.400 ;
        RECT 271.950 96.600 274.050 97.050 ;
        RECT 277.950 96.600 280.050 97.050 ;
        RECT 271.950 95.400 280.050 96.600 ;
        RECT 271.950 94.950 274.050 95.400 ;
        RECT 277.950 94.950 280.050 95.400 ;
        RECT 391.950 96.600 394.050 97.050 ;
        RECT 400.950 96.600 403.050 97.050 ;
        RECT 391.950 95.400 403.050 96.600 ;
        RECT 391.950 94.950 394.050 95.400 ;
        RECT 400.950 94.950 403.050 95.400 ;
        RECT 418.950 96.600 421.050 97.050 ;
        RECT 436.950 96.600 439.050 97.050 ;
        RECT 418.950 95.400 439.050 96.600 ;
        RECT 418.950 94.950 421.050 95.400 ;
        RECT 436.950 94.950 439.050 95.400 ;
        RECT 835.950 96.600 838.050 97.050 ;
        RECT 835.950 95.400 852.600 96.600 ;
        RECT 835.950 94.950 838.050 95.400 ;
        RECT 61.950 93.600 64.050 94.050 ;
        RECT 119.400 93.600 120.600 94.950 ;
        RECT 61.950 92.400 120.600 93.600 ;
        RECT 196.950 93.600 199.050 94.050 ;
        RECT 238.950 93.600 241.050 94.050 ;
        RECT 268.950 93.600 271.050 94.050 ;
        RECT 196.950 92.400 237.600 93.600 ;
        RECT 61.950 91.950 64.050 92.400 ;
        RECT 196.950 91.950 199.050 92.400 ;
        RECT 4.950 90.600 7.050 91.050 ;
        RECT 16.950 90.600 19.050 91.050 ;
        RECT 4.950 89.400 19.050 90.600 ;
        RECT 236.400 90.600 237.600 92.400 ;
        RECT 238.950 92.400 271.050 93.600 ;
        RECT 238.950 91.950 241.050 92.400 ;
        RECT 268.950 91.950 271.050 92.400 ;
        RECT 316.950 93.600 319.050 94.050 ;
        RECT 361.950 93.600 364.050 94.050 ;
        RECT 316.950 92.400 364.050 93.600 ;
        RECT 316.950 91.950 319.050 92.400 ;
        RECT 361.950 91.950 364.050 92.400 ;
        RECT 472.950 93.600 475.050 94.050 ;
        RECT 526.950 93.600 529.050 94.050 ;
        RECT 616.950 93.600 619.050 94.050 ;
        RECT 673.950 93.600 676.050 94.050 ;
        RECT 709.950 93.600 712.050 94.050 ;
        RECT 715.950 93.600 718.050 94.050 ;
        RECT 790.950 93.600 793.050 93.900 ;
        RECT 472.950 92.400 793.050 93.600 ;
        RECT 472.950 91.950 475.050 92.400 ;
        RECT 526.950 91.950 529.050 92.400 ;
        RECT 616.950 91.950 619.050 92.400 ;
        RECT 673.950 91.950 676.050 92.400 ;
        RECT 709.950 91.950 712.050 92.400 ;
        RECT 715.950 91.950 718.050 92.400 ;
        RECT 790.950 91.800 793.050 92.400 ;
        RECT 799.950 93.600 802.050 94.050 ;
        RECT 823.950 93.600 826.050 94.050 ;
        RECT 799.950 92.400 826.050 93.600 ;
        RECT 851.400 93.600 852.600 95.400 ;
        RECT 865.950 93.600 868.050 94.050 ;
        RECT 851.400 92.400 868.050 93.600 ;
        RECT 799.950 91.950 802.050 92.400 ;
        RECT 823.950 91.950 826.050 92.400 ;
        RECT 865.950 91.950 868.050 92.400 ;
        RECT 259.950 90.600 262.050 91.050 ;
        RECT 236.400 89.400 262.050 90.600 ;
        RECT 4.950 88.950 7.050 89.400 ;
        RECT 16.950 88.950 19.050 89.400 ;
        RECT 259.950 88.950 262.050 89.400 ;
        RECT 478.950 90.600 481.050 91.050 ;
        RECT 535.950 90.600 538.050 91.050 ;
        RECT 478.950 89.400 538.050 90.600 ;
        RECT 478.950 88.950 481.050 89.400 ;
        RECT 535.950 88.950 538.050 89.400 ;
        RECT 568.950 90.600 571.050 91.050 ;
        RECT 625.950 90.600 628.050 91.050 ;
        RECT 568.950 89.400 628.050 90.600 ;
        RECT 568.950 88.950 571.050 89.400 ;
        RECT 625.950 88.950 628.050 89.400 ;
        RECT 721.950 90.600 724.050 91.050 ;
        RECT 739.950 90.600 742.050 91.050 ;
        RECT 745.950 90.600 748.050 91.050 ;
        RECT 721.950 89.400 748.050 90.600 ;
        RECT 721.950 88.950 724.050 89.400 ;
        RECT 739.950 88.950 742.050 89.400 ;
        RECT 745.950 88.950 748.050 89.400 ;
        RECT 796.950 90.600 799.050 91.050 ;
        RECT 853.950 90.600 856.050 91.050 ;
        RECT 796.950 89.400 856.050 90.600 ;
        RECT 796.950 88.950 799.050 89.400 ;
        RECT 853.950 88.950 856.050 89.400 ;
        RECT 64.950 87.600 67.050 88.050 ;
        RECT 115.950 87.600 118.050 88.050 ;
        RECT 64.950 86.400 118.050 87.600 ;
        RECT 64.950 85.950 67.050 86.400 ;
        RECT 115.950 85.950 118.050 86.400 ;
        RECT 214.950 87.600 217.050 88.050 ;
        RECT 442.950 87.600 445.050 88.050 ;
        RECT 214.950 86.400 445.050 87.600 ;
        RECT 214.950 85.950 217.050 86.400 ;
        RECT 442.950 85.950 445.050 86.400 ;
        RECT 691.950 87.600 694.050 88.050 ;
        RECT 703.950 87.600 706.050 88.050 ;
        RECT 784.950 87.600 787.050 88.050 ;
        RECT 691.950 86.400 787.050 87.600 ;
        RECT 691.950 85.950 694.050 86.400 ;
        RECT 703.950 85.950 706.050 86.400 ;
        RECT 784.950 85.950 787.050 86.400 ;
        RECT 832.950 87.600 835.050 88.050 ;
        RECT 850.950 87.600 853.050 88.050 ;
        RECT 832.950 86.400 853.050 87.600 ;
        RECT 832.950 85.950 835.050 86.400 ;
        RECT 850.950 85.950 853.050 86.400 ;
        RECT 79.950 84.600 82.050 85.050 ;
        RECT 91.950 84.600 94.050 85.050 ;
        RECT 79.950 83.400 94.050 84.600 ;
        RECT 79.950 82.950 82.050 83.400 ;
        RECT 91.950 82.950 94.050 83.400 ;
        RECT 136.950 84.600 139.050 85.050 ;
        RECT 172.950 84.600 175.050 85.050 ;
        RECT 136.950 83.400 175.050 84.600 ;
        RECT 136.950 82.950 139.050 83.400 ;
        RECT 172.950 82.950 175.050 83.400 ;
        RECT 358.950 84.600 361.050 85.050 ;
        RECT 403.950 84.600 406.050 85.050 ;
        RECT 358.950 83.400 406.050 84.600 ;
        RECT 358.950 82.950 361.050 83.400 ;
        RECT 403.950 82.950 406.050 83.400 ;
        RECT 445.950 84.600 448.050 85.050 ;
        RECT 523.950 84.600 526.050 85.050 ;
        RECT 445.950 83.400 526.050 84.600 ;
        RECT 445.950 82.950 448.050 83.400 ;
        RECT 523.950 82.950 526.050 83.400 ;
        RECT 58.950 81.600 61.050 82.050 ;
        RECT 115.950 81.600 118.050 82.050 ;
        RECT 166.950 81.600 169.050 82.050 ;
        RECT 217.950 81.600 220.050 82.050 ;
        RECT 229.950 81.600 232.050 82.050 ;
        RECT 250.950 81.600 253.050 82.050 ;
        RECT 271.950 81.600 274.050 82.050 ;
        RECT 298.950 81.600 301.050 82.050 ;
        RECT 328.950 81.600 331.050 82.050 ;
        RECT 58.950 80.400 331.050 81.600 ;
        RECT 58.950 79.950 61.050 80.400 ;
        RECT 115.950 79.950 118.050 80.400 ;
        RECT 166.950 79.950 169.050 80.400 ;
        RECT 217.950 79.950 220.050 80.400 ;
        RECT 229.950 79.950 232.050 80.400 ;
        RECT 250.950 79.950 253.050 80.400 ;
        RECT 271.950 79.950 274.050 80.400 ;
        RECT 298.950 79.950 301.050 80.400 ;
        RECT 328.950 79.950 331.050 80.400 ;
        RECT 718.950 81.600 721.050 82.050 ;
        RECT 751.950 81.600 754.050 82.050 ;
        RECT 718.950 80.400 754.050 81.600 ;
        RECT 718.950 79.950 721.050 80.400 ;
        RECT 751.950 79.950 754.050 80.400 ;
        RECT 151.950 78.600 154.050 79.050 ;
        RECT 160.950 78.600 163.050 79.050 ;
        RECT 151.950 77.400 163.050 78.600 ;
        RECT 151.950 76.950 154.050 77.400 ;
        RECT 160.950 76.950 163.050 77.400 ;
        RECT 688.950 78.600 691.050 79.050 ;
        RECT 688.950 77.400 849.600 78.600 ;
        RECT 688.950 76.950 691.050 77.400 ;
        RECT 94.950 75.600 97.050 76.050 ;
        RECT 214.950 75.600 217.050 76.050 ;
        RECT 94.950 74.400 217.050 75.600 ;
        RECT 94.950 73.950 97.050 74.400 ;
        RECT 214.950 73.950 217.050 74.400 ;
        RECT 733.950 75.600 736.050 76.050 ;
        RECT 844.950 75.600 847.050 76.050 ;
        RECT 733.950 74.400 847.050 75.600 ;
        RECT 848.400 75.600 849.600 77.400 ;
        RECT 880.950 75.600 883.050 76.050 ;
        RECT 848.400 74.400 883.050 75.600 ;
        RECT 733.950 73.950 736.050 74.400 ;
        RECT 844.950 73.950 847.050 74.400 ;
        RECT 880.950 73.950 883.050 74.400 ;
        RECT 16.950 72.600 19.050 73.050 ;
        RECT 52.950 72.600 55.050 73.050 ;
        RECT 70.950 72.600 73.050 73.050 ;
        RECT 16.950 71.400 73.050 72.600 ;
        RECT 16.950 70.950 19.050 71.400 ;
        RECT 52.950 70.950 55.050 71.400 ;
        RECT 70.950 70.950 73.050 71.400 ;
        RECT 229.950 72.600 232.050 73.050 ;
        RECT 364.950 72.600 367.050 73.050 ;
        RECT 229.950 71.400 367.050 72.600 ;
        RECT 229.950 70.950 232.050 71.400 ;
        RECT 364.950 70.950 367.050 71.400 ;
        RECT 454.950 72.600 457.050 73.050 ;
        RECT 502.950 72.600 505.050 73.050 ;
        RECT 514.950 72.600 517.050 73.050 ;
        RECT 454.950 71.400 517.050 72.600 ;
        RECT 454.950 70.950 457.050 71.400 ;
        RECT 502.950 70.950 505.050 71.400 ;
        RECT 514.950 70.950 517.050 71.400 ;
        RECT 253.950 69.600 256.050 70.050 ;
        RECT 427.950 69.600 430.050 70.050 ;
        RECT 253.950 68.400 430.050 69.600 ;
        RECT 253.950 67.950 256.050 68.400 ;
        RECT 427.950 67.950 430.050 68.400 ;
        RECT 442.950 69.600 445.050 70.050 ;
        RECT 472.950 69.600 475.050 70.050 ;
        RECT 505.950 69.600 508.050 70.050 ;
        RECT 442.950 68.400 508.050 69.600 ;
        RECT 442.950 67.950 445.050 68.400 ;
        RECT 472.950 67.950 475.050 68.400 ;
        RECT 505.950 67.950 508.050 68.400 ;
        RECT 730.950 69.600 733.050 70.050 ;
        RECT 748.950 69.600 751.050 70.050 ;
        RECT 760.950 69.600 763.050 70.050 ;
        RECT 730.950 68.400 763.050 69.600 ;
        RECT 730.950 67.950 733.050 68.400 ;
        RECT 748.950 67.950 751.050 68.400 ;
        RECT 760.950 67.950 763.050 68.400 ;
        RECT 55.950 66.600 58.050 67.050 ;
        RECT 70.950 66.600 73.050 67.050 ;
        RECT 55.950 65.400 73.050 66.600 ;
        RECT 55.950 64.950 58.050 65.400 ;
        RECT 70.950 64.950 73.050 65.400 ;
        RECT 172.950 66.600 175.050 67.050 ;
        RECT 229.950 66.600 232.050 67.050 ;
        RECT 172.950 65.400 232.050 66.600 ;
        RECT 172.950 64.950 175.050 65.400 ;
        RECT 229.950 64.950 232.050 65.400 ;
        RECT 310.950 66.600 313.050 67.050 ;
        RECT 361.950 66.600 364.050 67.050 ;
        RECT 310.950 65.400 364.050 66.600 ;
        RECT 310.950 64.950 313.050 65.400 ;
        RECT 361.950 64.950 364.050 65.400 ;
        RECT 595.950 66.600 598.050 67.050 ;
        RECT 643.950 66.600 646.050 67.050 ;
        RECT 712.950 66.600 715.050 67.050 ;
        RECT 595.950 65.400 646.050 66.600 ;
        RECT 595.950 64.950 598.050 65.400 ;
        RECT 643.950 64.950 646.050 65.400 ;
        RECT 698.400 65.400 715.050 66.600 ;
        RECT 61.950 63.600 64.050 64.050 ;
        RECT 56.400 62.400 64.050 63.600 ;
        RECT 25.950 60.600 28.050 61.050 ;
        RECT 34.950 60.600 37.050 61.200 ;
        RECT 25.950 59.400 37.050 60.600 ;
        RECT 25.950 58.950 28.050 59.400 ;
        RECT 34.950 59.100 37.050 59.400 ;
        RECT 56.400 54.900 57.600 62.400 ;
        RECT 61.950 61.950 64.050 62.400 ;
        RECT 85.950 63.600 88.050 64.050 ;
        RECT 97.950 63.600 100.050 64.050 ;
        RECT 85.950 62.400 100.050 63.600 ;
        RECT 85.950 61.950 88.050 62.400 ;
        RECT 97.950 61.950 100.050 62.400 ;
        RECT 388.950 63.600 391.050 64.050 ;
        RECT 415.950 63.600 418.050 64.050 ;
        RECT 469.950 63.600 472.050 64.050 ;
        RECT 487.950 63.600 490.050 64.050 ;
        RECT 388.950 62.400 490.050 63.600 ;
        RECT 388.950 61.950 391.050 62.400 ;
        RECT 415.950 61.950 418.050 62.400 ;
        RECT 469.950 61.950 472.050 62.400 ;
        RECT 487.950 61.950 490.050 62.400 ;
        RECT 568.950 63.600 571.050 64.050 ;
        RECT 577.950 63.600 580.050 64.050 ;
        RECT 586.950 63.600 589.050 64.050 ;
        RECT 568.950 62.400 589.050 63.600 ;
        RECT 568.950 61.950 571.050 62.400 ;
        RECT 577.950 61.950 580.050 62.400 ;
        RECT 586.950 61.950 589.050 62.400 ;
        RECT 634.950 63.600 637.050 64.050 ;
        RECT 646.950 63.600 649.050 64.050 ;
        RECT 698.400 63.600 699.600 65.400 ;
        RECT 712.950 64.950 715.050 65.400 ;
        RECT 826.950 66.600 829.050 67.050 ;
        RECT 838.950 66.600 841.050 67.050 ;
        RECT 859.950 66.600 862.050 67.050 ;
        RECT 826.950 65.400 862.050 66.600 ;
        RECT 826.950 64.950 829.050 65.400 ;
        RECT 838.950 64.950 841.050 65.400 ;
        RECT 859.950 64.950 862.050 65.400 ;
        RECT 634.950 62.400 649.050 63.600 ;
        RECT 634.950 61.950 637.050 62.400 ;
        RECT 646.950 61.950 649.050 62.400 ;
        RECT 695.400 62.400 699.600 63.600 ;
        RECT 736.950 63.600 739.050 64.050 ;
        RECT 742.950 63.600 745.050 64.050 ;
        RECT 736.950 62.400 745.050 63.600 ;
        RECT 58.950 59.100 61.050 61.200 ;
        RECT 67.950 60.750 70.050 61.200 ;
        RECT 79.950 60.750 82.050 61.200 ;
        RECT 67.950 59.550 82.050 60.750 ;
        RECT 67.950 59.100 70.050 59.550 ;
        RECT 79.950 59.100 82.050 59.550 ;
        RECT 55.950 52.800 58.050 54.900 ;
        RECT 59.400 54.600 60.600 59.100 ;
        RECT 91.950 58.950 94.050 61.050 ;
        RECT 100.950 60.600 103.050 61.200 ;
        RECT 98.400 59.400 103.050 60.600 ;
        RECT 92.400 55.050 93.600 58.950 ;
        RECT 98.400 55.050 99.600 59.400 ;
        RECT 100.950 59.100 103.050 59.400 ;
        RECT 106.950 60.750 109.050 61.200 ;
        RECT 112.950 60.750 115.050 61.200 ;
        RECT 106.950 59.550 115.050 60.750 ;
        RECT 106.950 59.100 109.050 59.550 ;
        RECT 112.950 59.100 115.050 59.550 ;
        RECT 121.950 59.100 124.050 61.200 ;
        RECT 127.950 60.750 130.050 61.200 ;
        RECT 145.950 60.750 148.050 61.200 ;
        RECT 127.950 59.550 148.050 60.750 ;
        RECT 127.950 59.100 130.050 59.550 ;
        RECT 145.950 59.100 148.050 59.550 ;
        RECT 64.950 54.600 67.050 55.050 ;
        RECT 59.400 53.400 67.050 54.600 ;
        RECT 64.950 52.950 67.050 53.400 ;
        RECT 91.950 52.950 94.050 55.050 ;
        RECT 97.950 52.950 100.050 55.050 ;
        RECT 103.950 54.600 106.050 54.900 ;
        RECT 122.400 54.600 123.600 59.100 ;
        RECT 151.950 58.950 154.050 61.050 ;
        RECT 181.950 60.600 184.050 61.200 ;
        RECT 205.950 60.600 208.050 61.200 ;
        RECT 181.950 59.400 208.050 60.600 ;
        RECT 181.950 59.100 184.050 59.400 ;
        RECT 205.950 59.100 208.050 59.400 ;
        RECT 211.950 59.100 214.050 61.200 ;
        RECT 226.950 59.100 229.050 61.200 ;
        RECT 232.950 59.100 235.050 61.200 ;
        RECT 250.950 60.600 253.050 61.050 ;
        RECT 256.950 60.600 259.050 61.050 ;
        RECT 286.950 60.600 289.050 61.200 ;
        RECT 250.950 59.400 289.050 60.600 ;
        RECT 152.400 55.050 153.600 58.950 ;
        RECT 103.950 53.400 123.600 54.600 ;
        RECT 103.950 52.800 106.050 53.400 ;
        RECT 151.950 52.950 154.050 55.050 ;
        RECT 172.950 54.450 175.050 54.900 ;
        RECT 184.950 54.600 187.050 54.900 ;
        RECT 208.950 54.600 211.050 54.900 ;
        RECT 184.950 54.450 211.050 54.600 ;
        RECT 172.950 53.400 211.050 54.450 ;
        RECT 212.400 54.600 213.600 59.100 ;
        RECT 223.950 54.600 226.050 54.900 ;
        RECT 212.400 53.400 226.050 54.600 ;
        RECT 172.950 53.250 187.050 53.400 ;
        RECT 172.950 52.800 175.050 53.250 ;
        RECT 184.950 52.800 187.050 53.250 ;
        RECT 208.950 52.800 211.050 53.400 ;
        RECT 223.950 52.800 226.050 53.400 ;
        RECT 227.400 52.050 228.600 59.100 ;
        RECT 233.400 55.050 234.600 59.100 ;
        RECT 250.950 58.950 253.050 59.400 ;
        RECT 256.950 58.950 259.050 59.400 ;
        RECT 286.950 59.100 289.050 59.400 ;
        RECT 304.950 59.100 307.050 61.200 ;
        RECT 328.950 59.100 331.050 61.200 ;
        RECT 334.950 59.100 337.050 61.200 ;
        RECT 358.950 60.600 361.050 61.050 ;
        RECT 370.950 60.600 373.050 61.200 ;
        RECT 358.950 59.400 373.050 60.600 ;
        RECT 233.400 53.400 238.050 55.050 ;
        RECT 305.400 54.600 306.600 59.100 ;
        RECT 325.950 54.600 328.050 54.900 ;
        RECT 305.400 53.400 328.050 54.600 ;
        RECT 234.000 52.950 238.050 53.400 ;
        RECT 325.950 52.800 328.050 53.400 ;
        RECT 82.950 51.600 85.050 52.050 ;
        RECT 94.950 51.600 97.050 52.050 ;
        RECT 136.950 51.600 139.050 52.050 ;
        RECT 82.950 50.400 97.050 51.600 ;
        RECT 82.950 49.950 85.050 50.400 ;
        RECT 94.950 49.950 97.050 50.400 ;
        RECT 131.400 50.400 139.050 51.600 ;
        RECT 131.400 49.050 132.600 50.400 ;
        RECT 136.950 49.950 139.050 50.400 ;
        RECT 226.950 49.950 229.050 52.050 ;
        RECT 307.950 51.600 310.050 52.050 ;
        RECT 316.950 51.600 319.050 52.050 ;
        RECT 307.950 50.400 319.050 51.600 ;
        RECT 329.400 51.600 330.600 59.100 ;
        RECT 335.400 54.600 336.600 59.100 ;
        RECT 358.950 58.950 361.050 59.400 ;
        RECT 370.950 59.100 373.050 59.400 ;
        RECT 376.950 60.600 379.050 61.200 ;
        RECT 412.950 60.600 415.050 61.200 ;
        RECT 376.950 59.400 415.050 60.600 ;
        RECT 376.950 59.100 379.050 59.400 ;
        RECT 412.950 59.100 415.050 59.400 ;
        RECT 418.950 60.750 421.050 61.200 ;
        RECT 424.950 60.750 427.050 61.200 ;
        RECT 418.950 59.550 427.050 60.750 ;
        RECT 418.950 59.100 421.050 59.550 ;
        RECT 424.950 59.100 427.050 59.550 ;
        RECT 436.950 60.600 439.050 61.200 ;
        RECT 445.950 60.600 448.050 61.050 ;
        RECT 436.950 59.400 448.050 60.600 ;
        RECT 436.950 59.100 439.050 59.400 ;
        RECT 340.950 57.600 343.050 58.050 ;
        RECT 340.950 56.400 351.600 57.600 ;
        RECT 340.950 55.950 343.050 56.400 ;
        RECT 346.950 54.600 349.050 54.900 ;
        RECT 335.400 53.400 349.050 54.600 ;
        RECT 350.400 54.600 351.600 56.400 ;
        RECT 352.950 54.600 355.050 54.900 ;
        RECT 350.400 53.400 355.050 54.600 ;
        RECT 346.950 52.800 349.050 53.400 ;
        RECT 352.950 52.800 355.050 53.400 ;
        RECT 361.950 54.600 364.050 55.050 ;
        RECT 373.950 54.600 376.050 54.900 ;
        RECT 361.950 53.400 376.050 54.600 ;
        RECT 361.950 52.950 364.050 53.400 ;
        RECT 373.950 52.800 376.050 53.400 ;
        RECT 397.950 54.600 400.050 54.900 ;
        RECT 413.400 54.600 414.600 59.100 ;
        RECT 445.950 58.950 448.050 59.400 ;
        RECT 460.950 59.100 463.050 61.200 ;
        RECT 499.950 60.600 502.050 61.200 ;
        RECT 541.950 60.600 544.050 61.200 ;
        RECT 571.950 60.600 574.050 61.050 ;
        RECT 499.950 59.400 544.050 60.600 ;
        RECT 499.950 59.100 502.050 59.400 ;
        RECT 541.950 59.100 544.050 59.400 ;
        RECT 566.400 59.400 574.050 60.600 ;
        RECT 461.400 55.050 462.600 59.100 ;
        RECT 397.950 53.400 414.600 54.600 ;
        RECT 445.950 54.450 448.050 54.900 ;
        RECT 451.950 54.450 454.050 54.900 ;
        RECT 397.950 52.800 400.050 53.400 ;
        RECT 445.950 53.250 454.050 54.450 ;
        RECT 461.400 53.400 466.050 55.050 ;
        RECT 566.400 54.900 567.600 59.400 ;
        RECT 571.950 58.950 574.050 59.400 ;
        RECT 577.950 60.600 580.050 60.900 ;
        RECT 607.950 60.600 610.050 61.200 ;
        RECT 577.950 59.400 610.050 60.600 ;
        RECT 577.950 58.800 580.050 59.400 ;
        RECT 607.950 59.100 610.050 59.400 ;
        RECT 619.950 60.750 622.050 61.200 ;
        RECT 625.950 60.750 628.050 61.200 ;
        RECT 619.950 59.550 628.050 60.750 ;
        RECT 619.950 59.100 622.050 59.550 ;
        RECT 625.950 59.100 628.050 59.550 ;
        RECT 667.950 60.750 670.050 61.200 ;
        RECT 679.950 60.750 682.050 61.200 ;
        RECT 667.950 59.550 682.050 60.750 ;
        RECT 667.950 59.100 670.050 59.550 ;
        RECT 679.950 59.100 682.050 59.550 ;
        RECT 634.950 57.600 637.050 58.050 ;
        RECT 605.400 56.400 637.050 57.600 ;
        RECT 605.400 54.900 606.600 56.400 ;
        RECT 634.950 55.950 637.050 56.400 ;
        RECT 445.950 52.800 448.050 53.250 ;
        RECT 451.950 52.800 454.050 53.250 ;
        RECT 462.000 52.950 466.050 53.400 ;
        RECT 472.950 54.450 475.050 54.900 ;
        RECT 481.950 54.450 484.050 54.900 ;
        RECT 472.950 53.250 484.050 54.450 ;
        RECT 472.950 52.800 475.050 53.250 ;
        RECT 481.950 52.800 484.050 53.250 ;
        RECT 502.950 54.450 505.050 54.900 ;
        RECT 517.950 54.450 520.050 54.900 ;
        RECT 502.950 53.250 520.050 54.450 ;
        RECT 502.950 52.800 505.050 53.250 ;
        RECT 517.950 52.800 520.050 53.250 ;
        RECT 544.950 54.600 547.050 54.900 ;
        RECT 559.950 54.600 562.050 54.900 ;
        RECT 544.950 53.400 562.050 54.600 ;
        RECT 544.950 52.800 547.050 53.400 ;
        RECT 559.950 52.800 562.050 53.400 ;
        RECT 565.950 52.800 568.050 54.900 ;
        RECT 577.950 54.450 580.050 54.900 ;
        RECT 583.950 54.450 586.050 54.900 ;
        RECT 577.950 53.250 586.050 54.450 ;
        RECT 577.950 52.800 580.050 53.250 ;
        RECT 583.950 52.800 586.050 53.250 ;
        RECT 589.950 54.450 592.050 54.900 ;
        RECT 595.950 54.450 598.050 54.900 ;
        RECT 589.950 53.250 598.050 54.450 ;
        RECT 589.950 52.800 592.050 53.250 ;
        RECT 595.950 52.800 598.050 53.250 ;
        RECT 604.950 52.800 607.050 54.900 ;
        RECT 610.950 54.600 613.050 54.900 ;
        RECT 619.950 54.600 622.050 55.050 ;
        RECT 610.950 53.400 622.050 54.600 ;
        RECT 610.950 52.800 613.050 53.400 ;
        RECT 619.950 52.950 622.050 53.400 ;
        RECT 628.950 54.600 631.050 54.900 ;
        RECT 640.950 54.600 643.050 54.900 ;
        RECT 628.950 53.400 643.050 54.600 ;
        RECT 628.950 52.800 631.050 53.400 ;
        RECT 640.950 52.800 643.050 53.400 ;
        RECT 646.950 54.450 649.050 54.900 ;
        RECT 652.950 54.450 655.050 54.900 ;
        RECT 646.950 53.250 655.050 54.450 ;
        RECT 646.950 52.800 649.050 53.250 ;
        RECT 652.950 52.800 655.050 53.250 ;
        RECT 679.950 54.600 682.050 55.050 ;
        RECT 695.400 54.900 696.600 62.400 ;
        RECT 736.950 61.950 739.050 62.400 ;
        RECT 742.950 61.950 745.050 62.400 ;
        RECT 778.950 63.600 781.050 64.050 ;
        RECT 799.950 63.600 802.050 64.050 ;
        RECT 778.950 62.400 802.050 63.600 ;
        RECT 778.950 61.950 781.050 62.400 ;
        RECT 799.950 61.950 802.050 62.400 ;
        RECT 808.950 63.600 811.050 64.050 ;
        RECT 817.950 63.600 820.050 64.050 ;
        RECT 808.950 62.400 820.050 63.600 ;
        RECT 808.950 61.950 811.050 62.400 ;
        RECT 817.950 61.950 820.050 62.400 ;
        RECT 841.950 63.600 844.050 64.050 ;
        RECT 874.950 63.600 877.050 64.050 ;
        RECT 886.950 63.600 889.050 64.050 ;
        RECT 841.950 62.400 855.600 63.600 ;
        RECT 841.950 61.950 844.050 62.400 ;
        RECT 854.400 61.200 855.600 62.400 ;
        RECT 874.950 62.400 889.050 63.600 ;
        RECT 874.950 61.950 877.050 62.400 ;
        RECT 886.950 61.950 889.050 62.400 ;
        RECT 703.950 60.600 706.050 61.050 ;
        RECT 721.950 60.750 724.050 61.200 ;
        RECT 727.950 60.750 730.050 61.200 ;
        RECT 721.950 60.600 730.050 60.750 ;
        RECT 703.950 59.550 730.050 60.600 ;
        RECT 703.950 59.400 724.050 59.550 ;
        RECT 703.950 58.950 706.050 59.400 ;
        RECT 721.950 59.100 724.050 59.400 ;
        RECT 727.950 59.100 730.050 59.550 ;
        RECT 733.950 59.100 736.050 61.200 ;
        RECT 754.950 59.100 757.050 61.200 ;
        RECT 763.950 60.600 766.050 61.050 ;
        RECT 811.950 60.600 814.050 61.050 ;
        RECT 844.950 60.600 847.050 61.050 ;
        RECT 763.950 59.400 798.600 60.600 ;
        RECT 688.950 54.600 691.050 54.900 ;
        RECT 679.950 53.400 691.050 54.600 ;
        RECT 679.950 52.950 682.050 53.400 ;
        RECT 688.950 52.800 691.050 53.400 ;
        RECT 694.950 52.800 697.050 54.900 ;
        RECT 700.950 54.600 703.050 55.050 ;
        RECT 709.950 54.600 712.050 54.900 ;
        RECT 700.950 54.450 712.050 54.600 ;
        RECT 718.950 54.600 721.050 54.900 ;
        RECT 730.950 54.600 733.050 54.900 ;
        RECT 718.950 54.450 733.050 54.600 ;
        RECT 700.950 53.400 733.050 54.450 ;
        RECT 734.400 54.600 735.600 59.100 ;
        RECT 739.950 54.600 742.050 55.050 ;
        RECT 734.400 53.400 742.050 54.600 ;
        RECT 755.400 54.600 756.600 59.100 ;
        RECT 763.950 58.950 766.050 59.400 ;
        RECT 769.950 54.600 772.050 55.050 ;
        RECT 797.400 54.900 798.600 59.400 ;
        RECT 811.950 59.400 847.050 60.600 ;
        RECT 811.950 58.950 814.050 59.400 ;
        RECT 844.950 58.950 847.050 59.400 ;
        RECT 853.950 60.600 856.050 61.200 ;
        RECT 868.950 60.600 871.050 61.050 ;
        RECT 853.950 59.400 871.050 60.600 ;
        RECT 853.950 59.100 856.050 59.400 ;
        RECT 868.950 58.950 871.050 59.400 ;
        RECT 883.950 58.950 886.050 61.050 ;
        RECT 884.400 55.050 885.600 58.950 ;
        RECT 755.400 53.400 772.050 54.600 ;
        RECT 700.950 52.950 703.050 53.400 ;
        RECT 709.950 53.250 721.050 53.400 ;
        RECT 709.950 52.800 712.050 53.250 ;
        RECT 718.950 52.800 721.050 53.250 ;
        RECT 730.950 52.800 733.050 53.400 ;
        RECT 739.950 52.950 742.050 53.400 ;
        RECT 769.950 52.950 772.050 53.400 ;
        RECT 775.950 54.450 778.050 54.900 ;
        RECT 784.950 54.450 787.050 54.900 ;
        RECT 775.950 53.250 787.050 54.450 ;
        RECT 775.950 52.800 778.050 53.250 ;
        RECT 784.950 52.800 787.050 53.250 ;
        RECT 796.950 52.800 799.050 54.900 ;
        RECT 847.950 54.450 850.050 54.900 ;
        RECT 856.950 54.450 859.050 54.900 ;
        RECT 847.950 53.250 859.050 54.450 ;
        RECT 847.950 52.800 850.050 53.250 ;
        RECT 856.950 52.800 859.050 53.250 ;
        RECT 871.950 54.450 874.050 54.900 ;
        RECT 877.950 54.450 880.050 54.900 ;
        RECT 871.950 53.250 880.050 54.450 ;
        RECT 871.950 52.800 874.050 53.250 ;
        RECT 877.950 52.800 880.050 53.250 ;
        RECT 883.950 52.950 886.050 55.050 ;
        RECT 340.950 51.600 343.050 52.050 ;
        RECT 329.400 50.400 343.050 51.600 ;
        RECT 307.950 49.950 310.050 50.400 ;
        RECT 316.950 49.950 319.050 50.400 ;
        RECT 340.950 49.950 343.050 50.400 ;
        RECT 352.950 51.600 355.050 52.050 ;
        RECT 385.950 51.600 388.050 52.050 ;
        RECT 352.950 50.400 388.050 51.600 ;
        RECT 352.950 49.950 355.050 50.400 ;
        RECT 385.950 49.950 388.050 50.400 ;
        RECT 403.950 51.600 406.050 52.050 ;
        RECT 415.950 51.600 418.050 52.050 ;
        RECT 403.950 50.400 418.050 51.600 ;
        RECT 403.950 49.950 406.050 50.400 ;
        RECT 415.950 49.950 418.050 50.400 ;
        RECT 721.950 51.600 724.050 52.050 ;
        RECT 757.950 51.600 760.050 52.050 ;
        RECT 805.950 51.600 808.050 52.050 ;
        RECT 721.950 50.400 808.050 51.600 ;
        RECT 721.950 49.950 724.050 50.400 ;
        RECT 757.950 49.950 760.050 50.400 ;
        RECT 805.950 49.950 808.050 50.400 ;
        RECT 31.950 48.600 34.050 49.050 ;
        RECT 130.950 48.600 133.050 49.050 ;
        RECT 31.950 47.400 133.050 48.600 ;
        RECT 31.950 46.950 34.050 47.400 ;
        RECT 130.950 46.950 133.050 47.400 ;
        RECT 148.950 48.600 151.050 49.050 ;
        RECT 283.950 48.600 286.050 48.900 ;
        RECT 403.950 48.600 406.050 48.900 ;
        RECT 424.950 48.600 427.050 49.050 ;
        RECT 148.950 47.400 427.050 48.600 ;
        RECT 148.950 46.950 151.050 47.400 ;
        RECT 283.950 46.800 286.050 47.400 ;
        RECT 403.950 46.800 406.050 47.400 ;
        RECT 424.950 46.950 427.050 47.400 ;
        RECT 451.950 48.600 454.050 49.050 ;
        RECT 463.950 48.600 466.050 49.050 ;
        RECT 451.950 47.400 466.050 48.600 ;
        RECT 451.950 46.950 454.050 47.400 ;
        RECT 463.950 46.950 466.050 47.400 ;
        RECT 793.950 48.600 796.050 49.050 ;
        RECT 814.950 48.600 817.050 49.050 ;
        RECT 823.950 48.600 826.050 49.050 ;
        RECT 793.950 47.400 826.050 48.600 ;
        RECT 793.950 46.950 796.050 47.400 ;
        RECT 814.950 46.950 817.050 47.400 ;
        RECT 823.950 46.950 826.050 47.400 ;
        RECT 871.950 48.600 874.050 49.050 ;
        RECT 892.950 48.600 895.050 49.050 ;
        RECT 871.950 47.400 895.050 48.600 ;
        RECT 871.950 46.950 874.050 47.400 ;
        RECT 892.950 46.950 895.050 47.400 ;
        RECT 46.950 45.600 49.050 46.050 ;
        RECT 64.950 45.600 67.050 46.050 ;
        RECT 46.950 44.400 67.050 45.600 ;
        RECT 46.950 43.950 49.050 44.400 ;
        RECT 64.950 43.950 67.050 44.400 ;
        RECT 79.950 45.600 82.050 46.050 ;
        RECT 91.950 45.600 94.050 46.050 ;
        RECT 79.950 44.400 94.050 45.600 ;
        RECT 79.950 43.950 82.050 44.400 ;
        RECT 91.950 43.950 94.050 44.400 ;
        RECT 223.950 45.600 226.050 46.050 ;
        RECT 250.950 45.600 253.050 46.050 ;
        RECT 223.950 44.400 253.050 45.600 ;
        RECT 223.950 43.950 226.050 44.400 ;
        RECT 250.950 43.950 253.050 44.400 ;
        RECT 670.950 45.600 673.050 46.050 ;
        RECT 691.950 45.600 694.050 46.050 ;
        RECT 670.950 44.400 694.050 45.600 ;
        RECT 670.950 43.950 673.050 44.400 ;
        RECT 691.950 43.950 694.050 44.400 ;
        RECT 736.950 45.600 739.050 46.050 ;
        RECT 787.950 45.600 790.050 46.050 ;
        RECT 736.950 44.400 790.050 45.600 ;
        RECT 736.950 43.950 739.050 44.400 ;
        RECT 787.950 43.950 790.050 44.400 ;
        RECT 850.950 45.600 853.050 46.050 ;
        RECT 883.950 45.600 886.050 46.050 ;
        RECT 850.950 44.400 886.050 45.600 ;
        RECT 850.950 43.950 853.050 44.400 ;
        RECT 883.950 43.950 886.050 44.400 ;
        RECT 58.950 42.600 61.050 43.050 ;
        RECT 70.950 42.600 73.050 43.050 ;
        RECT 58.950 41.400 73.050 42.600 ;
        RECT 58.950 40.950 61.050 41.400 ;
        RECT 70.950 40.950 73.050 41.400 ;
        RECT 196.950 42.600 199.050 43.050 ;
        RECT 229.950 42.600 232.050 43.050 ;
        RECT 196.950 41.400 232.050 42.600 ;
        RECT 196.950 40.950 199.050 41.400 ;
        RECT 229.950 40.950 232.050 41.400 ;
        RECT 238.950 42.600 241.050 43.050 ;
        RECT 244.950 42.600 247.050 43.050 ;
        RECT 238.950 41.400 247.050 42.600 ;
        RECT 238.950 40.950 241.050 41.400 ;
        RECT 244.950 40.950 247.050 41.400 ;
        RECT 397.950 42.600 400.050 43.050 ;
        RECT 496.950 42.600 499.050 43.050 ;
        RECT 397.950 41.400 499.050 42.600 ;
        RECT 397.950 40.950 400.050 41.400 ;
        RECT 496.950 40.950 499.050 41.400 ;
        RECT 790.950 42.600 793.050 43.050 ;
        RECT 832.950 42.600 835.050 43.050 ;
        RECT 790.950 41.400 835.050 42.600 ;
        RECT 790.950 40.950 793.050 41.400 ;
        RECT 832.950 40.950 835.050 41.400 ;
        RECT 13.950 39.600 16.050 40.050 ;
        RECT 46.950 39.600 49.050 40.050 ;
        RECT 13.950 38.400 49.050 39.600 ;
        RECT 13.950 37.950 16.050 38.400 ;
        RECT 46.950 37.950 49.050 38.400 ;
        RECT 265.950 39.600 268.050 40.050 ;
        RECT 283.800 39.600 285.900 40.050 ;
        RECT 265.950 38.400 285.900 39.600 ;
        RECT 265.950 37.950 268.050 38.400 ;
        RECT 283.800 37.950 285.900 38.400 ;
        RECT 286.950 39.600 289.050 40.050 ;
        RECT 340.950 39.600 343.050 40.050 ;
        RECT 286.950 38.400 343.050 39.600 ;
        RECT 286.950 37.950 289.050 38.400 ;
        RECT 340.950 37.950 343.050 38.400 ;
        RECT 388.950 39.600 391.050 40.050 ;
        RECT 394.950 39.600 397.050 40.050 ;
        RECT 388.950 38.400 397.050 39.600 ;
        RECT 388.950 37.950 391.050 38.400 ;
        RECT 394.950 37.950 397.050 38.400 ;
        RECT 427.950 39.600 430.050 40.050 ;
        RECT 664.950 39.600 667.050 40.050 ;
        RECT 427.950 38.400 667.050 39.600 ;
        RECT 427.950 37.950 430.050 38.400 ;
        RECT 664.950 37.950 667.050 38.400 ;
        RECT 733.950 39.600 736.050 40.050 ;
        RECT 745.950 39.600 748.050 40.050 ;
        RECT 733.950 38.400 748.050 39.600 ;
        RECT 733.950 37.950 736.050 38.400 ;
        RECT 745.950 37.950 748.050 38.400 ;
        RECT 145.950 36.600 148.050 37.050 ;
        RECT 253.950 36.600 256.050 37.050 ;
        RECT 145.950 35.400 256.050 36.600 ;
        RECT 145.950 34.950 148.050 35.400 ;
        RECT 253.950 34.950 256.050 35.400 ;
        RECT 370.950 36.600 373.050 37.050 ;
        RECT 379.950 36.600 382.050 37.050 ;
        RECT 397.950 36.600 400.050 37.050 ;
        RECT 409.950 36.600 412.050 37.050 ;
        RECT 370.950 35.400 412.050 36.600 ;
        RECT 370.950 34.950 373.050 35.400 ;
        RECT 379.950 34.950 382.050 35.400 ;
        RECT 397.950 34.950 400.050 35.400 ;
        RECT 409.950 34.950 412.050 35.400 ;
        RECT 844.950 36.600 847.050 37.050 ;
        RECT 877.950 36.600 880.050 37.050 ;
        RECT 844.950 35.400 880.050 36.600 ;
        RECT 844.950 34.950 847.050 35.400 ;
        RECT 877.950 34.950 880.050 35.400 ;
        RECT 22.950 33.600 25.050 34.050 ;
        RECT 31.950 33.600 34.050 34.050 ;
        RECT 22.950 32.400 34.050 33.600 ;
        RECT 22.950 31.950 25.050 32.400 ;
        RECT 31.950 31.950 34.050 32.400 ;
        RECT 277.950 33.600 280.050 34.050 ;
        RECT 304.950 33.600 307.050 34.050 ;
        RECT 277.950 32.400 307.050 33.600 ;
        RECT 277.950 31.950 280.050 32.400 ;
        RECT 304.950 31.950 307.050 32.400 ;
        RECT 340.950 33.600 343.050 34.050 ;
        RECT 358.950 33.600 361.050 34.050 ;
        RECT 340.950 32.400 361.050 33.600 ;
        RECT 340.950 31.950 343.050 32.400 ;
        RECT 358.950 31.950 361.050 32.400 ;
        RECT 418.950 33.600 421.050 34.050 ;
        RECT 430.950 33.600 433.050 34.050 ;
        RECT 418.950 32.400 433.050 33.600 ;
        RECT 418.950 31.950 421.050 32.400 ;
        RECT 430.950 31.950 433.050 32.400 ;
        RECT 457.950 33.600 460.050 34.050 ;
        RECT 475.950 33.600 478.050 34.050 ;
        RECT 457.950 32.400 478.050 33.600 ;
        RECT 457.950 31.950 460.050 32.400 ;
        RECT 475.950 31.950 478.050 32.400 ;
        RECT 538.950 33.600 541.050 34.050 ;
        RECT 553.950 33.600 556.050 34.050 ;
        RECT 538.950 32.400 556.050 33.600 ;
        RECT 538.950 31.950 541.050 32.400 ;
        RECT 553.950 31.950 556.050 32.400 ;
        RECT 577.950 33.600 580.050 34.050 ;
        RECT 682.950 33.600 685.050 34.050 ;
        RECT 577.950 32.400 685.050 33.600 ;
        RECT 577.950 31.950 580.050 32.400 ;
        RECT 682.950 31.950 685.050 32.400 ;
        RECT 808.950 33.600 811.050 34.050 ;
        RECT 814.950 33.600 817.050 34.050 ;
        RECT 808.950 32.400 817.050 33.600 ;
        RECT 808.950 31.950 811.050 32.400 ;
        RECT 814.950 31.950 817.050 32.400 ;
        RECT 826.950 33.600 829.050 34.050 ;
        RECT 835.950 33.600 838.050 34.050 ;
        RECT 826.950 32.400 838.050 33.600 ;
        RECT 826.950 31.950 829.050 32.400 ;
        RECT 835.950 31.950 838.050 32.400 ;
        RECT 13.950 28.950 16.050 31.050 ;
        RECT 178.950 30.600 181.050 31.050 ;
        RECT 187.950 30.600 190.050 31.050 ;
        RECT 298.950 30.600 301.050 31.050 ;
        RECT 178.950 29.400 190.050 30.600 ;
        RECT 178.950 28.950 181.050 29.400 ;
        RECT 187.950 28.950 190.050 29.400 ;
        RECT 290.400 29.400 301.050 30.600 ;
        RECT 14.400 21.900 15.600 28.950 ;
        RECT 16.950 27.600 19.050 28.200 ;
        RECT 31.950 27.600 34.050 28.200 ;
        RECT 85.950 28.050 88.050 28.500 ;
        RECT 97.950 28.050 100.050 28.500 ;
        RECT 16.950 26.400 34.050 27.600 ;
        RECT 16.950 26.100 19.050 26.400 ;
        RECT 31.950 26.100 34.050 26.400 ;
        RECT 37.950 27.600 40.050 28.050 ;
        RECT 85.950 27.600 100.050 28.050 ;
        RECT 37.950 26.850 100.050 27.600 ;
        RECT 37.950 26.400 88.050 26.850 ;
        RECT 97.950 26.400 100.050 26.850 ;
        RECT 148.950 27.600 151.050 28.200 ;
        RECT 166.950 27.600 169.050 28.050 ;
        RECT 187.950 27.600 190.050 28.500 ;
        RECT 148.950 26.400 169.050 27.600 ;
        RECT 37.950 25.950 40.050 26.400 ;
        RECT 148.950 26.100 151.050 26.400 ;
        RECT 166.950 25.950 169.050 26.400 ;
        RECT 179.400 26.400 190.050 27.600 ;
        RECT 256.950 27.600 259.050 28.200 ;
        RECT 268.950 27.600 271.050 28.050 ;
        RECT 286.950 27.600 289.050 28.050 ;
        RECT 256.950 26.400 271.050 27.600 ;
        RECT 38.400 24.600 39.600 25.950 ;
        RECT 124.950 24.600 127.050 25.050 ;
        RECT 35.400 23.400 39.600 24.600 ;
        RECT 104.400 23.400 127.050 24.600 ;
        RECT 35.400 21.900 36.600 23.400 ;
        RECT 13.950 19.800 16.050 21.900 ;
        RECT 22.950 21.450 25.050 21.900 ;
        RECT 28.950 21.450 31.050 21.900 ;
        RECT 22.950 20.250 31.050 21.450 ;
        RECT 22.950 19.800 25.050 20.250 ;
        RECT 28.950 19.800 31.050 20.250 ;
        RECT 34.950 19.800 37.050 21.900 ;
        RECT 104.400 21.600 105.600 23.400 ;
        RECT 124.950 22.950 127.050 23.400 ;
        RECT 179.400 21.900 180.600 26.400 ;
        RECT 256.950 26.100 259.050 26.400 ;
        RECT 268.950 25.950 271.050 26.400 ;
        RECT 281.400 26.400 289.050 27.600 ;
        RECT 133.950 21.600 136.050 21.900 ;
        RECT 151.950 21.600 154.050 21.900 ;
        RECT 103.950 19.500 106.050 21.600 ;
        RECT 133.950 20.400 154.050 21.600 ;
        RECT 133.950 19.800 136.050 20.400 ;
        RECT 151.950 19.800 154.050 20.400 ;
        RECT 166.950 21.450 169.050 21.900 ;
        RECT 172.950 21.450 175.050 21.900 ;
        RECT 166.950 20.250 175.050 21.450 ;
        RECT 166.950 19.800 169.050 20.250 ;
        RECT 172.950 19.800 175.050 20.250 ;
        RECT 178.950 19.800 181.050 21.900 ;
        RECT 238.950 21.600 241.050 21.900 ;
        RECT 244.950 21.600 247.050 22.050 ;
        RECT 281.400 21.900 282.600 26.400 ;
        RECT 286.950 25.950 289.050 26.400 ;
        RECT 253.950 21.600 256.050 21.900 ;
        RECT 199.950 21.150 202.050 21.600 ;
        RECT 205.950 21.150 208.050 21.600 ;
        RECT 199.950 19.950 208.050 21.150 ;
        RECT 199.950 19.500 202.050 19.950 ;
        RECT 205.950 19.500 208.050 19.950 ;
        RECT 214.950 21.150 217.050 21.600 ;
        RECT 220.950 21.150 223.050 21.600 ;
        RECT 214.950 19.950 223.050 21.150 ;
        RECT 214.950 19.500 217.050 19.950 ;
        RECT 220.950 19.500 223.050 19.950 ;
        RECT 238.950 20.400 256.050 21.600 ;
        RECT 238.950 19.800 241.050 20.400 ;
        RECT 244.950 19.950 247.050 20.400 ;
        RECT 253.950 19.800 256.050 20.400 ;
        RECT 259.950 21.450 262.050 21.900 ;
        RECT 265.950 21.450 268.050 21.900 ;
        RECT 259.950 20.250 268.050 21.450 ;
        RECT 259.950 19.800 262.050 20.250 ;
        RECT 265.950 19.800 268.050 20.250 ;
        RECT 280.950 19.800 283.050 21.900 ;
        RECT 290.400 21.600 291.600 29.400 ;
        RECT 298.950 28.950 301.050 29.400 ;
        RECT 766.950 30.600 769.050 31.050 ;
        RECT 823.950 30.600 826.050 31.050 ;
        RECT 766.950 29.400 826.050 30.600 ;
        RECT 766.950 28.950 769.050 29.400 ;
        RECT 823.950 28.950 826.050 29.400 ;
        RECT 856.950 30.600 859.050 31.050 ;
        RECT 868.950 30.600 871.050 31.050 ;
        RECT 856.950 29.400 871.050 30.600 ;
        RECT 856.950 28.950 859.050 29.400 ;
        RECT 868.950 28.950 871.050 29.400 ;
        RECT 316.950 27.600 319.050 28.500 ;
        RECT 331.950 27.600 334.050 28.200 ;
        RECT 316.950 26.400 334.050 27.600 ;
        RECT 331.950 26.100 334.050 26.400 ;
        RECT 346.950 27.750 349.050 28.200 ;
        RECT 355.950 27.750 358.050 28.200 ;
        RECT 346.950 27.600 358.050 27.750 ;
        RECT 361.950 27.600 364.050 28.500 ;
        RECT 409.950 27.600 412.050 28.200 ;
        RECT 442.950 28.050 445.050 28.500 ;
        RECT 463.950 28.050 466.050 28.500 ;
        RECT 346.950 26.550 364.050 27.600 ;
        RECT 346.950 26.100 349.050 26.550 ;
        RECT 355.950 26.400 364.050 26.550 ;
        RECT 395.400 26.400 412.050 27.600 ;
        RECT 355.950 26.100 358.050 26.400 ;
        RECT 304.950 21.600 307.050 22.050 ;
        RECT 289.950 19.500 292.050 21.600 ;
        RECT 298.950 20.400 307.050 21.600 ;
        RECT 298.950 19.500 301.050 20.400 ;
        RECT 304.950 19.950 307.050 20.400 ;
        RECT 352.950 21.450 355.050 21.900 ;
        RECT 370.950 21.450 373.050 21.900 ;
        RECT 395.400 21.600 396.600 26.400 ;
        RECT 409.950 26.100 412.050 26.400 ;
        RECT 424.950 27.600 429.000 28.050 ;
        RECT 424.950 25.950 429.600 27.600 ;
        RECT 442.950 26.850 466.050 28.050 ;
        RECT 442.950 26.400 445.050 26.850 ;
        RECT 463.950 26.400 466.050 26.850 ;
        RECT 472.950 27.600 475.050 28.050 ;
        RECT 511.950 27.600 514.050 28.050 ;
        RECT 523.950 27.600 526.050 28.200 ;
        RECT 472.950 26.400 492.600 27.600 ;
        RECT 472.950 25.950 475.050 26.400 ;
        RECT 428.400 21.900 429.600 25.950 ;
        RECT 352.950 20.250 373.050 21.450 ;
        RECT 352.950 19.800 355.050 20.250 ;
        RECT 370.950 19.800 373.050 20.250 ;
        RECT 379.950 20.400 396.600 21.600 ;
        RECT 397.950 21.450 400.050 21.900 ;
        RECT 406.950 21.450 409.050 21.900 ;
        RECT 379.950 19.500 382.050 20.400 ;
        RECT 397.950 20.250 409.050 21.450 ;
        RECT 397.950 19.800 400.050 20.250 ;
        RECT 406.950 19.800 409.050 20.250 ;
        RECT 412.950 21.450 415.050 21.900 ;
        RECT 418.950 21.450 421.050 21.900 ;
        RECT 412.950 20.250 421.050 21.450 ;
        RECT 412.950 19.800 415.050 20.250 ;
        RECT 418.950 19.800 421.050 20.250 ;
        RECT 427.950 19.800 430.050 21.900 ;
        RECT 433.950 21.600 436.050 21.900 ;
        RECT 442.950 21.600 445.050 22.050 ;
        RECT 448.950 21.600 451.050 21.900 ;
        RECT 491.400 21.600 492.600 26.400 ;
        RECT 511.950 26.400 526.050 27.600 ;
        RECT 511.950 25.950 514.050 26.400 ;
        RECT 523.950 26.100 526.050 26.400 ;
        RECT 529.950 27.600 532.050 28.200 ;
        RECT 580.950 28.050 583.050 28.500 ;
        RECT 589.950 28.050 592.050 28.500 ;
        RECT 544.950 27.600 547.050 28.050 ;
        RECT 529.950 26.400 547.050 27.600 ;
        RECT 580.950 26.850 592.050 28.050 ;
        RECT 616.950 27.750 619.050 28.200 ;
        RECT 625.950 27.750 628.050 28.200 ;
        RECT 616.950 27.600 628.050 27.750 ;
        RECT 580.950 26.400 583.050 26.850 ;
        RECT 589.950 26.400 592.050 26.850 ;
        RECT 614.400 26.550 628.050 27.600 ;
        RECT 614.400 26.400 619.050 26.550 ;
        RECT 529.950 26.100 532.050 26.400 ;
        RECT 508.950 21.600 511.050 21.900 ;
        RECT 524.400 21.600 525.600 26.100 ;
        RECT 544.950 25.950 547.050 26.400 ;
        RECT 577.950 24.600 580.050 25.050 ;
        RECT 563.400 23.400 580.050 24.600 ;
        RECT 433.950 20.400 451.050 21.600 ;
        RECT 433.950 19.800 436.050 20.400 ;
        RECT 442.950 19.950 445.050 20.400 ;
        RECT 448.950 19.800 451.050 20.400 ;
        RECT 475.950 21.150 478.050 21.600 ;
        RECT 481.950 21.150 484.050 21.600 ;
        RECT 475.950 19.950 484.050 21.150 ;
        RECT 475.950 19.500 478.050 19.950 ;
        RECT 481.950 19.500 484.050 19.950 ;
        RECT 490.950 19.500 493.050 21.600 ;
        RECT 508.950 20.400 525.600 21.600 ;
        RECT 532.950 21.450 535.050 21.900 ;
        RECT 538.950 21.450 541.050 21.900 ;
        RECT 563.400 21.600 564.600 23.400 ;
        RECT 577.950 22.950 580.050 23.400 ;
        RECT 614.400 21.900 615.600 26.400 ;
        RECT 616.950 26.100 619.050 26.400 ;
        RECT 625.950 26.100 628.050 26.550 ;
        RECT 631.950 27.750 634.050 28.200 ;
        RECT 652.950 27.750 655.050 28.200 ;
        RECT 631.950 26.550 655.050 27.750 ;
        RECT 712.950 27.600 715.050 28.200 ;
        RECT 631.950 26.100 634.050 26.550 ;
        RECT 652.950 26.100 655.050 26.550 ;
        RECT 689.400 26.400 715.050 27.600 ;
        RECT 682.950 24.600 685.050 25.050 ;
        RECT 671.400 23.400 685.050 24.600 ;
        RECT 508.950 19.800 511.050 20.400 ;
        RECT 532.950 20.250 541.050 21.450 ;
        RECT 532.950 19.800 535.050 20.250 ;
        RECT 538.950 19.800 541.050 20.250 ;
        RECT 562.950 19.500 565.050 21.600 ;
        RECT 613.950 19.800 616.050 21.900 ;
        RECT 619.950 21.450 622.050 21.900 ;
        RECT 628.950 21.450 631.050 21.900 ;
        RECT 619.950 20.250 631.050 21.450 ;
        RECT 619.950 19.800 622.050 20.250 ;
        RECT 628.950 19.800 631.050 20.250 ;
        RECT 652.950 21.600 655.050 22.050 ;
        RECT 671.400 21.600 672.600 23.400 ;
        RECT 682.950 22.950 685.050 23.400 ;
        RECT 689.400 21.900 690.600 26.400 ;
        RECT 712.950 26.100 715.050 26.400 ;
        RECT 718.950 27.600 721.050 28.200 ;
        RECT 733.950 27.600 736.050 28.200 ;
        RECT 718.950 26.400 736.050 27.600 ;
        RECT 718.950 26.100 721.050 26.400 ;
        RECT 733.950 26.100 736.050 26.400 ;
        RECT 748.950 27.750 751.050 28.200 ;
        RECT 760.950 27.750 763.050 28.200 ;
        RECT 748.950 26.550 763.050 27.750 ;
        RECT 748.950 26.100 751.050 26.550 ;
        RECT 760.950 26.100 763.050 26.550 ;
        RECT 793.950 27.600 796.050 28.050 ;
        RECT 805.950 27.600 808.050 28.200 ;
        RECT 793.950 26.400 808.050 27.600 ;
        RECT 793.950 25.950 796.050 26.400 ;
        RECT 805.950 26.100 808.050 26.400 ;
        RECT 814.950 24.600 817.050 25.050 ;
        RECT 803.400 23.400 817.050 24.600 ;
        RECT 652.950 20.400 664.050 21.600 ;
        RECT 652.950 19.950 655.050 20.400 ;
        RECT 661.950 19.500 664.050 20.400 ;
        RECT 670.950 19.500 673.050 21.600 ;
        RECT 688.950 19.800 691.050 21.900 ;
        RECT 694.950 21.450 697.050 21.900 ;
        RECT 700.950 21.450 703.050 21.900 ;
        RECT 694.950 20.250 703.050 21.450 ;
        RECT 694.950 19.800 697.050 20.250 ;
        RECT 700.950 19.800 703.050 20.250 ;
        RECT 736.950 21.600 739.050 21.900 ;
        RECT 745.950 21.600 748.050 22.050 ;
        RECT 754.950 21.600 757.050 21.900 ;
        RECT 736.950 20.400 757.050 21.600 ;
        RECT 736.950 19.800 739.050 20.400 ;
        RECT 745.950 19.950 748.050 20.400 ;
        RECT 754.950 19.800 757.050 20.400 ;
        RECT 763.950 21.600 766.050 21.900 ;
        RECT 769.950 21.600 772.050 22.050 ;
        RECT 803.400 21.900 804.600 23.400 ;
        RECT 814.950 22.950 817.050 23.400 ;
        RECT 778.950 21.600 781.050 21.900 ;
        RECT 763.950 20.400 781.050 21.600 ;
        RECT 763.950 19.800 766.050 20.400 ;
        RECT 769.950 19.950 772.050 20.400 ;
        RECT 778.950 19.800 781.050 20.400 ;
        RECT 787.950 21.450 790.050 21.900 ;
        RECT 793.950 21.450 796.050 21.900 ;
        RECT 787.950 20.250 796.050 21.450 ;
        RECT 787.950 19.800 790.050 20.250 ;
        RECT 793.950 19.800 796.050 20.250 ;
        RECT 802.950 19.800 805.050 21.900 ;
        RECT 808.950 21.600 811.050 21.900 ;
        RECT 826.950 21.600 829.050 21.900 ;
        RECT 808.950 20.400 829.050 21.600 ;
        RECT 808.950 19.800 811.050 20.400 ;
        RECT 826.950 19.800 829.050 20.400 ;
        RECT 835.950 21.450 838.050 21.900 ;
        RECT 841.950 21.450 844.050 21.900 ;
        RECT 835.950 20.250 844.050 21.450 ;
        RECT 835.950 19.800 838.050 20.250 ;
        RECT 841.950 19.800 844.050 20.250 ;
        RECT 847.950 21.450 850.050 21.900 ;
        RECT 856.950 21.450 859.050 21.900 ;
        RECT 847.950 20.250 859.050 21.450 ;
        RECT 847.950 19.800 850.050 20.250 ;
        RECT 856.950 19.800 859.050 20.250 ;
        RECT 868.950 21.450 871.050 21.900 ;
        RECT 886.950 21.450 889.050 21.900 ;
        RECT 868.950 20.250 889.050 21.450 ;
        RECT 868.950 19.800 871.050 20.250 ;
        RECT 886.950 19.800 889.050 20.250 ;
        RECT 514.950 18.600 517.050 19.050 ;
        RECT 526.950 18.600 529.050 19.050 ;
        RECT 550.950 18.600 553.050 19.050 ;
        RECT 514.950 17.400 553.050 18.600 ;
        RECT 514.950 16.950 517.050 17.400 ;
        RECT 526.950 16.950 529.050 17.400 ;
        RECT 550.950 16.950 553.050 17.400 ;
        RECT 709.950 18.600 712.050 19.050 ;
        RECT 727.950 18.600 730.050 19.050 ;
        RECT 709.950 17.400 730.050 18.600 ;
        RECT 709.950 16.950 712.050 17.400 ;
        RECT 727.950 16.950 730.050 17.400 ;
        RECT 454.950 15.600 457.050 16.050 ;
        RECT 515.400 15.600 516.600 16.950 ;
        RECT 454.950 14.400 516.600 15.600 ;
        RECT 556.950 15.600 559.050 16.050 ;
        RECT 580.950 15.600 583.050 16.050 ;
        RECT 607.950 15.600 610.050 16.050 ;
        RECT 556.950 14.400 610.050 15.600 ;
        RECT 454.950 13.950 457.050 14.400 ;
        RECT 556.950 13.950 559.050 14.400 ;
        RECT 580.950 13.950 583.050 14.400 ;
        RECT 607.950 13.950 610.050 14.400 ;
        RECT 622.950 15.600 625.050 16.050 ;
        RECT 634.950 15.600 637.050 16.050 ;
        RECT 622.950 14.400 637.050 15.600 ;
        RECT 622.950 13.950 625.050 14.400 ;
        RECT 634.950 13.950 637.050 14.400 ;
        RECT 715.950 15.600 718.050 16.050 ;
        RECT 742.950 15.600 745.050 16.050 ;
        RECT 715.950 14.400 745.050 15.600 ;
        RECT 715.950 13.950 718.050 14.400 ;
        RECT 742.950 13.950 745.050 14.400 ;
        RECT 544.950 12.600 547.050 13.050 ;
        RECT 553.950 12.600 556.050 13.050 ;
        RECT 544.950 11.400 556.050 12.600 ;
        RECT 544.950 10.950 547.050 11.400 ;
        RECT 553.950 10.950 556.050 11.400 ;
        RECT 559.950 12.600 562.050 13.050 ;
        RECT 571.950 12.600 574.050 13.050 ;
        RECT 559.950 11.400 574.050 12.600 ;
        RECT 559.950 10.950 562.050 11.400 ;
        RECT 571.950 10.950 574.050 11.400 ;
        RECT 226.950 6.600 229.050 7.050 ;
        RECT 232.950 6.600 235.050 7.050 ;
        RECT 454.950 6.600 457.050 7.050 ;
        RECT 226.950 5.400 457.050 6.600 ;
        RECT 226.950 4.950 229.050 5.400 ;
        RECT 232.950 4.950 235.050 5.400 ;
        RECT 454.950 4.950 457.050 5.400 ;
        RECT 598.950 6.600 601.050 7.050 ;
        RECT 874.950 6.600 877.050 7.050 ;
        RECT 598.950 5.400 877.050 6.600 ;
        RECT 598.950 4.950 601.050 5.400 ;
        RECT 874.950 4.950 877.050 5.400 ;
  END
END fir_pe
END LIBRARY

