* NGSPICE file created from pong_pt1.ext - technology: scmos

.subckt INVX1 A Y vdd gnd
M1000 Y A gnd gnd nfet w=3u l=0.6u
+  ad=6.3p pd=10.2u as=6.3p ps=10.2u
M1001 Y A vdd vdd pfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=12.6p ps=16.2u
.ends

.subckt OAI21X1 A B C Y vdd gnd
M1000 Y C a_7_14# gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.4u
M1001 a_30_146# A vdd vdd pfet w=12u l=0.6u
+  ad=3.6p pd=12.6u as=25.2p ps=28.2u
M1002 vdd C Y vdd pfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=14.4p ps=14.7u
M1003 gnd A a_7_14# gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=12.6p ps=16.2u
M1004 Y B a_30_146# vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.7u as=3.6p ps=12.6u
M1005 a_7_14# B gnd gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
.ends

.subckt NAND2X1 A B Y vdd gnd
M1000 a_27_14# A gnd gnd nfet w=6u l=0.6u
+  ad=2.7p pd=6.9u as=12.6p ps=16.2u
M1001 Y B a_27_14# gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=2.7p ps=6.9u
M1002 vdd B Y vdd pfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.4u
M1003 Y A vdd vdd pfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=12.6p ps=16.2u
.ends

.subckt AOI21X1 A B C Y vdd gnd
M1000 vdd A a_7_146# vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=25.2p ps=28.2u
M1001 Y C a_7_146# vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=14.4p ps=14.4u
M1002 a_28_14# A gnd gnd nfet w=6u l=0.6u
+  ad=1.8p pd=6.6u as=12.6p ps=16.2u
M1003 Y B a_28_14# gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.7u as=1.8p ps=6.6u
M1004 a_7_146# B vdd vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
M1005 gnd C Y gnd nfet w=3u l=0.6u
+  ad=6.3p pd=10.2u as=7.2p ps=8.7u
.ends

.subckt NOR2X1 A B Y vdd gnd
M1000 a_25_146# A vdd vdd pfet w=12u l=0.6u
+  ad=3.6p pd=12.6u as=25.2p ps=28.2u
M1001 Y A gnd gnd nfet w=3u l=0.6u
+  ad=3.6p pd=5.4u as=6.3p ps=10.2u
M1002 Y B a_25_146# vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=3.6p ps=12.6u
M1003 gnd B Y gnd nfet w=3u l=0.6u
+  ad=6.3p pd=10.2u as=3.6p ps=5.4u
.ends

.subckt DFFSR R S D CLK Q vdd gnd
M1000 a_146_14# a_122_10# a_60_10# vdd pfet w=3u l=0.6u
+  ad=6.3p pd=8.4u as=3.6p ps=5.4u
M1001 a_64_14# a_60_10# gnd gnd nfet w=6u l=0.6u
+  ad=3.6p pd=7.2u as=9p ps=9u
M1002 vdd S a_301_14# vdd pfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.4u
M1003 a_146_14# a_115_95# a_60_10# gnd nfet w=3u l=0.6u
+  ad=3.6p pd=5.4u as=3.6p ps=5.4u
M1004 a_36_10# a_60_10# vdd vdd pfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1005 a_391_14# a_334_14# gnd gnd nfet w=6u l=0.6u
+  ad=3.6p pd=7.2u as=9.45p ps=9.15u
M1006 a_8_14# R vdd vdd pfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=12.6p ps=16.2u
M1007 a_36_10# S a_64_14# gnd nfet w=6u l=0.6u
+  ad=14.4p pd=16.8u as=3.6p ps=7.2u
M1008 gnd a_334_14# Q gnd nfet w=3u l=0.6u
+  ad=6.3p pd=10.2u as=6.3p ps=10.2u
M1009 a_281_14# a_122_10# a_36_10# gnd nfet w=3u l=0.6u
+  ad=3.6p pd=5.4u as=6.3p ps=10.2u
M1010 a_28_14# R a_8_14# gnd nfet w=6u l=0.6u
+  ad=3.6p pd=7.2u as=14.4p ps=16.8u
M1011 a_301_14# S a_391_14# gnd nfet w=6u l=0.6u
+  ad=14.4p pd=16.8u as=3.6p ps=7.2u
M1012 gnd a_36_10# a_28_14# gnd nfet w=6u l=0.6u
+  ad=9p pd=9u as=3.6p ps=7.2u
M1013 gnd a_115_95# a_122_10# gnd nfet w=3u l=0.6u
+  ad=3.6p pd=5.4u as=6.3p ps=10.2u
M1014 a_301_14# a_334_14# vdd vdd pfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1015 vdd D a_146_14# vdd pfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=6.3p ps=8.4u
M1016 a_334_14# a_281_14# vdd vdd pfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=12.6p ps=16.2u
M1017 vdd a_115_95# a_122_10# vdd pfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=12.6p ps=16.2u
M1018 a_301_14# a_122_10# a_281_14# vdd pfet w=3u l=0.6u
+  ad=6.3p pd=10.2u as=3.6p ps=5.4u
M1019 gnd D a_146_14# gnd nfet w=3u l=0.6u
+  ad=6.3p pd=10.2u as=3.6p ps=5.4u
M1020 a_60_10# a_115_95# a_8_14# vdd pfet w=3u l=0.6u
+  ad=3.6p pd=5.4u as=6.3p ps=10.2u
M1021 a_301_14# a_115_95# a_281_14# gnd nfet w=3u l=0.6u
+  ad=6.3p pd=10.2u as=3.6p ps=5.4u
M1022 vdd S a_36_10# vdd pfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.4u
M1023 vdd a_36_10# a_8_14# vdd pfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1024 a_115_95# CLK gnd gnd nfet w=3u l=0.6u
+  ad=6.3p pd=10.2u as=3.6p ps=5.4u
M1025 a_60_10# a_122_10# a_8_14# gnd nfet w=3u l=0.6u
+  ad=3.6p pd=5.4u as=6.3p ps=10.2u
M1026 a_354_14# a_281_14# a_334_14# gnd nfet w=6u l=0.6u
+  ad=3.6p pd=7.2u as=14.4p ps=16.8u
M1027 vdd R a_334_14# vdd pfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1028 a_115_95# CLK vdd vdd pfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.4u
M1029 a_281_14# a_115_95# a_36_10# vdd pfet w=3u l=0.6u
+  ad=3.6p pd=5.4u as=6.3p ps=10.2u
M1030 gnd R a_354_14# gnd nfet w=6u l=0.6u
+  ad=9.45p pd=9.15u as=3.6p ps=7.2u
M1031 vdd a_334_14# Q vdd pfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=12.6p ps=16.2u
.ends

.subckt BUFX2 A Y vdd gnd
M1000 Y a_7_14# vdd vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=14.4p ps=14.7u
M1001 gnd A a_7_14# gnd nfet w=3u l=0.6u
+  ad=7.2p pd=8.7u as=6.3p ps=10.2u
M1002 Y a_7_14# gnd gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.7u
M1003 vdd A a_7_14# vdd pfet w=6u l=0.6u
+  ad=14.4p pd=14.7u as=12.6p ps=16.2u
.ends

.subckt NAND3X1 A B C Y vdd gnd
M1000 Y C a_34_14# gnd nfet w=9u l=0.6u
+  ad=18.9p pd=22.2u as=2.7p ps=9.6u
M1001 a_26_14# A gnd gnd nfet w=9u l=0.6u
+  ad=2.7p pd=9.6u as=18.9p ps=22.2u
M1002 vdd B Y vdd pfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1003 a_34_14# B a_26_14# gnd nfet w=9u l=0.6u
+  ad=2.7p pd=9.6u as=2.7p ps=9.6u
M1004 Y C vdd vdd pfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.4u
M1005 Y A vdd vdd pfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=12.6p ps=16.2u
.ends

.subckt NOR3X1 A B C Y vdd gnd
M1000 gnd B Y gnd nfet w=3u l=0.6u
+  ad=3.6p pd=5.4u as=3.6p ps=5.4u
M1001 a_7_166# A vdd vdd pfet w=9u l=0.6u
+  ad=10.8p pd=11.4u as=10.8p ps=11.4u
M1002 a_7_166# B a_65_166# vdd pfet w=9u l=0.6u
+  ad=18.9p pd=22.2u as=10.8p ps=11.4u
M1003 a_65_166# C Y vdd pfet w=9u l=0.6u
+  ad=18.9p pd=22.2u as=10.8p ps=11.4u
M1004 Y C gnd gnd nfet w=3u l=0.6u
+  ad=6.3p pd=10.2u as=3.6p ps=5.4u
M1005 a_65_166# B a_7_166# vdd pfet w=9u l=0.6u
+  ad=10.8p pd=11.4u as=10.8p ps=11.4u
M1006 vdd A a_7_166# vdd pfet w=9u l=0.6u
+  ad=10.8p pd=11.4u as=18.9p ps=22.2u
M1007 Y C a_65_166# vdd pfet w=9u l=0.6u
+  ad=10.8p pd=11.4u as=18.9p ps=22.2u
M1008 Y A gnd gnd nfet w=3u l=0.6u
+  ad=3.6p pd=5.4u as=7.2p ps=10.8u
.ends

.subckt AND2X2 A B Y vdd gnd
M1000 a_25_14# A a_7_14# gnd nfet w=6u l=0.6u
+  ad=2.7p pd=6.9u as=12.6p ps=16.2u
M1001 gnd B a_25_14# gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=2.7p ps=6.9u
M1002 vdd B a_7_14# vdd pfet w=6u l=0.6u
+  ad=14.4p pd=14.7u as=8.1p ps=8.7u
M1003 Y a_7_14# gnd gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.4u
M1004 Y a_7_14# vdd vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=14.4p ps=14.7u
M1005 a_7_14# A vdd vdd pfet w=6u l=0.6u
+  ad=8.1p pd=8.7u as=12.6p ps=16.2u
.ends

.subckt INVX2 A Y vdd gnd
M1000 Y A vdd vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=25.2p ps=28.2u
M1001 Y A gnd gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=12.6p ps=16.2u
.ends

.subckt OR2X2 A B Y vdd gnd
M1000 Y a_7_146# gnd gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=6.3p ps=8.4u
M1001 a_25_146# A a_7_146# vdd pfet w=12u l=0.6u
+  ad=5.4p pd=12.9u as=25.2p ps=28.2u
M1002 a_7_146# A gnd gnd nfet w=3u l=0.6u
+  ad=3.6p pd=5.4u as=6.3p ps=10.2u
M1003 Y a_7_146# vdd vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=14.4p ps=14.4u
M1004 gnd B a_7_146# gnd nfet w=3u l=0.6u
+  ad=6.3p pd=8.4u as=3.6p ps=5.4u
M1005 vdd B a_25_146# vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=5.4p ps=12.9u
.ends

.subckt AOI22X1 A B C D Y vdd gnd
M1000 gnd C a_56_14# gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=1.8p ps=6.6u
M1001 vdd A a_7_146# vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=25.2p ps=28.2u
M1002 Y D a_7_146# vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
M1003 a_28_14# A gnd gnd nfet w=6u l=0.6u
+  ad=1.8p pd=6.6u as=12.6p ps=16.2u
M1004 Y B a_28_14# gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=1.8p ps=6.6u
M1005 a_7_146# C Y vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=14.4p ps=14.4u
M1006 a_7_146# B vdd vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
M1007 a_56_14# D Y gnd nfet w=6u l=0.6u
+  ad=1.8p pd=6.6u as=7.2p ps=8.4u
.ends

.subckt CLKBUF1 A Y vdd gnd
M1000 Y a_105_14# vdd vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
M1001 a_65_14# a_25_14# gnd gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1002 a_105_14# a_65_14# vdd vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
M1003 Y a_105_14# gnd gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1004 a_25_14# A vdd vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=25.2p ps=28.2u
M1005 a_65_14# a_25_14# vdd vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
M1006 a_25_14# A gnd gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=12.6p ps=16.2u
M1007 gnd a_25_14# a_65_14# gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1008 a_105_14# a_65_14# gnd gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1009 gnd a_105_14# Y gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.4u
M1010 vdd a_65_14# a_105_14# vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
M1011 vdd a_105_14# Y vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=14.4p ps=14.4u
M1012 vdd a_25_14# a_65_14# vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
M1013 gnd A a_25_14# gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1014 vdd A a_25_14# vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
M1015 gnd a_65_14# a_105_14# gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
.ends

.subckt OAI22X1 A B C D Y vdd gnd
M1000 Y D a_7_14# gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1001 a_25_146# A vdd vdd pfet w=12u l=0.6u
+  ad=5.4p pd=12.9u as=25.2p ps=28.2u
M1002 a_65_146# D Y vdd pfet w=12u l=0.6u
+  ad=5.4p pd=12.9u as=23.4p ps=15.9u
M1003 gnd A a_7_14# gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=12.6p ps=16.2u
M1004 a_7_14# C Y gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.4u
M1005 a_7_14# B gnd gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1006 Y B a_25_146# vdd pfet w=12u l=0.6u
+  ad=23.4p pd=15.9u as=5.4p ps=12.9u
M1007 vdd C a_65_146# vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=5.4p ps=12.9u
.ends

.subckt INVX8 A Y vdd gnd
M1000 Y A gnd gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1001 Y A vdd vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=25.2p ps=28.2u
M1002 Y A vdd vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
M1003 Y A gnd gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=12.6p ps=16.2u
M1004 gnd A Y gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.4u
M1005 vdd A Y vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=14.4p ps=14.4u
M1006 gnd A Y gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1007 vdd A Y vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
.ends

.subckt INVX4 A Y vdd gnd
M1000 Y A vdd vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=25.2p ps=28.2u
M1001 Y A gnd gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=12.6p ps=16.2u
M1002 gnd A Y gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.4u
M1003 vdd A Y vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=14.4p ps=14.4u
.ends

.subckt pong_pt1 gnd vdd clk down enable hsync p_tick reset rgb up vsync
X_1270_ _1916_/Q _1757_/C vdd gnd INVX1
X_1606_ _1606_/A _1606_/B _1651_/A _1607_/C vdd gnd OAI21X1
X_1399_ _1442_/B _1718_/B _1400_/A vdd gnd NAND2X1
X_1468_ _972_/A _975_/A _1469_/C vdd gnd NAND2X1
X_1537_ _1743_/A _1904_/B _1537_/C _1911_/D vdd gnd OAI21X1
X_981_ _981_/A _998_/B _981_/C _981_/Y vdd gnd OAI21X1
X_1322_ _1322_/A _1911_/Q _1912_/Q _1675_/A vdd gnd AOI21X1
X_1253_ _1253_/A _1253_/B _1254_/C vdd gnd NOR2X1
X_1184_ _1909_/Q _1487_/A _1300_/A vdd gnd NAND2X1
X_964_ _967_/B _964_/Y vdd gnd INVX1
X_1871_ _1871_/A _1871_/B _1871_/C _1872_/B vdd gnd OAI21X1
X_1940_ _1940_/R vdd _1940_/D _1940_/CLK _1940_/Q vdd gnd DFFSR
X_1236_ _950_/A _1787_/A _1236_/C _1262_/B vdd gnd AOI21X1
X_1305_ _1489_/B _1684_/B _1306_/B vdd gnd NAND2X1
X_1098_ _1845_/A _1111_/B _1101_/A vdd gnd NOR2X1
X_1167_ _949_/A _1167_/B _1210_/B vdd gnd NOR2X1
XBUFX2_insert0 _969_/Y _1074_/R vdd gnd BUFX2
X_947_ _947_/A _971_/C _947_/C _948_/A vdd gnd NAND3X1
X_1021_ _1021_/A _1063_/C _1072_/D vdd gnd NOR2X1
X_1854_ _1876_/A _1855_/B vdd gnd INVX1
X_1785_ _1785_/A _1785_/B _1786_/C vdd gnd NOR2X1
X_1923_ _1924_/R vdd _1923_/D _1940_/CLK _1923_/Q vdd gnd DFFSR
X_1219_ _1911_/Q _1487_/B _1226_/B vdd gnd NOR2X1
X_1570_ _1940_/Q _1787_/C _1583_/A vdd gnd NOR2X1
X_1004_ _1004_/A _998_/B _999_/Y _1069_/D vdd gnd OAI21X1
X_1768_ _1768_/A _1768_/B _1768_/C _1770_/A vdd gnd NOR3X1
X_1837_ _1937_/Q _1837_/B _1838_/A vdd gnd NAND2X1
X_1906_ _1906_/A _1907_/B _1907_/C _1939_/D vdd gnd OAI21X1
X_1699_ _1699_/A _1699_/B _1771_/B vdd gnd NAND2X1
X_1622_ _1635_/A _1622_/B _1627_/C vdd gnd NOR2X1
X_1553_ _1554_/B _1557_/A _1555_/B vdd gnd AND2X2
X_1484_ _973_/A _949_/A _1501_/B vdd gnd NOR2X1
X_1536_ _1602_/B _1536_/B _1536_/C _1537_/C vdd gnd NAND3X1
X_1605_ _1605_/A _1635_/A _1606_/B vdd gnd NOR2X1
X_1467_ _1467_/A _1467_/B _1476_/A vdd gnd AND2X2
X_1398_ _1398_/A _1398_/B _1718_/B vdd gnd NAND2X1
X_980_ _999_/A _999_/B _989_/B _981_/C vdd gnd OAI21X1
X_1321_ _1735_/C _1743_/A _1321_/C _1675_/B vdd gnd NOR3X1
X_1252_ _1482_/B _1914_/Q _1252_/C _1257_/B vdd gnd OAI21X1
X_1183_ _989_/A _1487_/A vdd gnd INVX2
X_1519_ _1543_/C _1543_/A _1520_/C vdd gnd OR2X2
X_963_ _963_/A _997_/C _999_/B _967_/B vdd gnd NAND3X1
X_1870_ _1870_/A _1870_/B _1872_/A vdd gnd NAND2X1
X_1304_ _1304_/A _1322_/A _1684_/B vdd gnd NAND2X1
X_1166_ _1166_/A _1166_/B _1166_/C _1339_/C vdd gnd OAI21X1
X_1235_ _950_/A _1787_/A _1251_/A _1236_/C vdd gnd OAI21X1
XBUFX2_insert1 _969_/Y _1071_/S vdd gnd BUFX2
X_1097_ _1932_/Q _1753_/B _1127_/B _1111_/B vdd gnd NAND3X1
X_1020_ _1020_/A _971_/B _999_/A _1063_/C vdd gnd AOI21X1
X_946_ _973_/B _972_/B _947_/C vdd gnd NOR2X1
X_1922_ _1924_/R vdd _1922_/D _1925_/CLK _1922_/Q vdd gnd DFFSR
X_1853_ _1853_/A _1853_/B _1876_/A _1856_/A vdd gnd NAND3X1
X_1784_ _1784_/A _1784_/B _1784_/C _1788_/A vdd gnd OAI21X1
X_1218_ _994_/A _1487_/B vdd gnd INVX1
X_1149_ _1287_/A _1208_/A _1289_/A vdd gnd NOR2X1
X_1003_ _1015_/B _1003_/B _997_/C _1004_/A vdd gnd NAND3X1
X_1905_ _1905_/A _1905_/B _1938_/D vdd gnd NAND2X1
X_1836_ _1837_/B _1937_/Q _1838_/B vdd gnd OR2X2
X_1767_ _1767_/A _1767_/B _1767_/C _1768_/C vdd gnd NAND3X1
X_1698_ _1698_/A _1705_/B _1699_/B vdd gnd NAND2X1
X_1621_ _1700_/C _1621_/B _1622_/B vdd gnd NOR2X1
X_1552_ _1552_/A _1552_/B _1557_/A vdd gnd NAND2X1
X_1483_ _1525_/C _1522_/A _1500_/B vdd gnd AND2X2
X_1819_ _1932_/Q _1928_/Q _1820_/A vdd gnd NOR2X1
X_1604_ _1650_/B _1635_/A vdd gnd INVX1
X_1535_ _1543_/B _1535_/B _1536_/B vdd gnd NAND2X1
X_1397_ _1921_/Q _1589_/C _1727_/A _1398_/A vdd gnd NAND3X1
X_1466_ _951_/B _1790_/A _1467_/B vdd gnd NAND2X1
X_1320_ _1677_/C _1677_/B _1702_/B vdd gnd AND2X2
X_1251_ _1251_/A _1255_/A _1252_/C vdd gnd AND2X2
X_1182_ _1182_/A _1261_/A _1199_/A vdd gnd NAND2X1
X_1449_ _1449_/A _1449_/B _1454_/C vdd gnd NAND2X1
X_1518_ _1543_/A _1543_/C _1530_/C vdd gnd NAND2X1
X_962_ _962_/A _962_/B _966_/A _997_/C vdd gnd OAI21X1
X_1303_ _1909_/Q _1908_/Q _1910_/Q _1304_/A vdd gnd OAI21X1
X_1096_ _1935_/Q _1845_/A vdd gnd INVX1
X_1165_ _1524_/B _1791_/A _1165_/C _1343_/A _1166_/C vdd gnd AOI22X1
X_1234_ _1256_/A _1255_/B _1251_/A vdd gnd NOR2X1
XBUFX2_insert2 _969_/Y _1082_/R vdd gnd BUFX2
X_945_ _975_/A _975_/B _971_/C vdd gnd NOR2X1
X_1852_ _1875_/B _1875_/A _1876_/A vdd gnd NAND2X1
X_1921_ _1925_/R vdd _1921_/D _1925_/CLK _1921_/Q vdd gnd DFFSR
X_1783_ _1783_/A _1783_/B _1783_/C _1784_/B vdd gnd AOI21X1
X_1217_ _1217_/A _1217_/B _1217_/C _1281_/B vdd gnd AOI21X1
X_1148_ _1930_/Q _1525_/B _1208_/A vdd gnd NOR2X1
X_1079_ _1083_/R vdd _1079_/D _1083_/CLK _975_/A vdd gnd DFFSR
X_1002_ _996_/C _991_/A _1013_/B _1003_/B vdd gnd OAI21X1
X_1904_ _1904_/A _1904_/B _1937_/D vdd gnd NOR2X1
X_1835_ _1928_/Q _1835_/B _1835_/C _1837_/B vdd gnd OAI21X1
X_1766_ _1766_/A _1766_/B _1767_/C vdd gnd AND2X2
X_1697_ _1924_/Q _1697_/B _1697_/C _1699_/A vdd gnd NAND3X1
X_1482_ _951_/A _1482_/B _1525_/C vdd gnd NOR2X1
X_1551_ _1913_/Q _1940_/Q _1552_/A vdd gnd NAND2X1
X_1620_ _1682_/A _1648_/B _1620_/C _1920_/D vdd gnd OAI21X1
X_1818_ _1818_/A _1845_/B _1820_/B vdd gnd NOR2X1
X_1749_ _1915_/Q _1749_/B _1749_/C _1914_/Q _1750_/C vdd gnd AOI22X1
X_1465_ _1465_/A _1465_/B _1465_/C _1467_/A vdd gnd NAND3X1
X_1534_ _1535_/B _1543_/B _1536_/C vdd gnd OR2X2
X_1603_ _1603_/A _1650_/B _1606_/A vdd gnd NOR2X1
X_1396_ _1920_/Q _1720_/C _1700_/C _1398_/B vdd gnd OAI21X1
X_1181_ _1261_/A _1182_/A _1199_/C vdd gnd OR2X2
X_1250_ _1914_/Q _1482_/B _1255_/A vdd gnd NAND2X1
X_1517_ _1517_/A _1517_/B _1543_/A vdd gnd NOR2X1
X_1448_ _994_/A _1920_/Q _1449_/A vdd gnd NAND2X1
X_1379_ _1919_/Q _1691_/C _1920_/Q _1781_/A vdd gnd OAI21X1
X_961_ _990_/A _990_/B _961_/C _962_/B vdd gnd NAND3X1
X_1302_ _1723_/A _1727_/C _1708_/B _1322_/A vdd gnd NAND3X1
X_1233_ _1915_/Q _1434_/A _1255_/B vdd gnd NOR2X1
X_1095_ _1161_/A _1161_/B _1163_/B vdd gnd NOR2X1
X_1164_ _1276_/B _1276_/C _1791_/A vdd gnd NAND2X1
XBUFX2_insert3 _969_/Y _1083_/R vdd gnd BUFX2
X_944_ _973_/A _972_/A _947_/A vdd gnd NOR2X1
X_1851_ _1851_/A _1851_/B _1898_/B vdd gnd NAND2X1
X_1920_ _1925_/R vdd _1920_/D _1925_/CLK _1920_/Q vdd gnd DFFSR
X_1782_ _1782_/A _1782_/B _1782_/C _1783_/C vdd gnd OAI21X1
X_1216_ _1216_/A _1216_/B _1217_/C vdd gnd OR2X2
X_1147_ _973_/A _1525_/B vdd gnd INVX1
X_1078_ _1083_/R vdd _1078_/D _1083_/CLK _972_/B vdd gnd DFFSR
X_1001_ _999_/C _1013_/B vdd gnd INVX1
XCLKBUF1_insert10 clk _1936_/CLK vdd gnd CLKBUF1
X_1834_ _1928_/Q _1834_/B _1835_/B _1835_/C vdd gnd NAND3X1
X_1765_ _1922_/Q _1765_/B _1767_/A vdd gnd NAND2X1
X_1903_ _1903_/A _1903_/B _1903_/C _1936_/D vdd gnd OAI21X1
X_1696_ _1696_/A _1696_/B _1771_/A vdd gnd AND2X2
X_1481_ _957_/A _999_/C _1522_/A vdd gnd NOR2X1
X_1550_ _1734_/C _1907_/A _1552_/B vdd gnd NAND2X1
X_1748_ _1914_/Q _1749_/C _1748_/C _1784_/A _1750_/A vdd gnd OAI22X1
X_1817_ _1871_/B _1871_/A _1870_/B vdd gnd NOR2X1
X_1679_ _1922_/Q _1765_/B _1679_/C _1771_/C vdd gnd AOI21X1
X_1602_ _1602_/A _1602_/B _1651_/A vdd gnd AND2X2
X_1464_ _1464_/A _1464_/B _1465_/C vdd gnd NOR2X1
X_1533_ _1533_/A _1533_/B _1543_/B vdd gnd NOR2X1
X_1395_ _1395_/A _1395_/B _1395_/C _1401_/C vdd gnd OAI21X1
X_1180_ _1191_/C _1191_/A _1190_/A _1182_/A vdd gnd OAI21X1
X_1516_ _1723_/A _1907_/A _1517_/B vdd gnd NOR2X1
X_1378_ _989_/A _989_/B _1378_/C _1691_/C _1395_/A vdd gnd AOI22X1
X_1447_ _1487_/B _1682_/A _1449_/B vdd gnd NAND2X1
X_960_ _989_/B _990_/B vdd gnd INVX1
X_1232_ _951_/A _1434_/A vdd gnd INVX1
X_1301_ _1487_/A _1497_/B _1301_/C _1306_/A vdd gnd OAI21X1
X_1094_ _1936_/Q _1935_/Q _1753_/B _1161_/A vdd gnd NAND3X1
X_1163_ _1904_/A _1163_/B _1276_/C vdd gnd NAND2X1
X_1781_ _1781_/A _1781_/B _1911_/Q _1782_/B vdd gnd AOI21X1
X_1850_ _1850_/A _1850_/B _1850_/C _1851_/A vdd gnd NAND3X1
X_1215_ _1215_/A _1215_/B _1215_/C _1217_/B vdd gnd NAND3X1
X_1146_ _1146_/A _1161_/B _1755_/B vdd gnd AND2X2
X_1077_ _1082_/R vdd _1077_/D _1083_/CLK _972_/A vdd gnd DFFSR
X_1000_ _999_/C _995_/A _995_/B _1015_/B vdd gnd NAND3X1
X_1902_ _1902_/A _1902_/B _1936_/Q _1903_/C vdd gnd OAI21X1
X_1833_ _1833_/A _1834_/B vdd gnd INVX1
X_1764_ _1764_/A _1797_/B vdd gnd INVX1
X_1695_ _1771_/C _1770_/B _1713_/C _1707_/C vdd gnd NAND3X1
X_1129_ _1141_/B _972_/A _1129_/C _1157_/A vdd gnd AOI21X1
X_1480_ _1938_/Q _1905_/A vdd gnd INVX1
X_1678_ _1766_/B _1766_/A _1767_/B _1679_/C vdd gnd NAND3X1
X_1816_ _1931_/Q _1928_/Q _1871_/B vdd gnd NOR2X1
X_1747_ _1747_/A _1783_/B _1748_/C vdd gnd NAND2X1
X_1532_ _1743_/A _1907_/A _1533_/B vdd gnd NOR2X1
X_1601_ _1601_/A _1601_/B _1917_/D vdd gnd NAND2X1
X_1394_ _1416_/B _1394_/B _1394_/C _1395_/C vdd gnd AOI21X1
X_1463_ _989_/A _1722_/C _1463_/C _1464_/B vdd gnd OAI21X1
X_1515_ _1940_/Q _1907_/A vdd gnd INVX2
X_1377_ _1453_/A _1453_/B _1378_/C vdd gnd OR2X2
X_1446_ _1446_/A _1460_/A _1464_/A vdd gnd NAND2X1
X_1162_ _1937_/Q _1904_/A vdd gnd INVX1
X_1231_ _951_/A _1787_/C _1256_/A vdd gnd NOR2X1
X_1300_ _1300_/A _1300_/B _1687_/B _1301_/C vdd gnd OAI21X1
X_1093_ _1109_/B _1753_/B vdd gnd INVX1
X_1429_ _1924_/Q _1925_/Q _1429_/C _1757_/A vdd gnd NAND3X1
X_1780_ _1780_/A _1780_/B _1780_/C _1783_/A vdd gnd OAI21X1
X_1214_ _1289_/B _1214_/B _1214_/C _1217_/A vdd gnd NAND3X1
X_1145_ _972_/A _1345_/C vdd gnd INVX1
X_1076_ _1082_/R vdd _1076_/D _1083_/CLK _973_/B vdd gnd DFFSR
X_1832_ _1832_/A _1841_/A _1875_/A _1835_/B vdd gnd NAND3X1
X_1901_ _1901_/A _1901_/B _1901_/C _1903_/B vdd gnd NAND3X1
X_1694_ _1694_/A _1694_/B _1694_/C _1712_/B _1770_/B vdd gnd OAI22X1
X_1763_ _1927_/Q _1798_/A vdd gnd INVX1
X_1128_ _1524_/A _1137_/B _1129_/C vdd gnd NOR2X1
X_1059_ _1059_/A _1059_/B _1059_/C _1060_/A vdd gnd OAI21X1
X_1815_ _1815_/A _1845_/B _1871_/A vdd gnd NOR2X1
X_1746_ _1785_/A _1747_/A vdd gnd INVX1
X_1677_ _1702_/A _1677_/B _1677_/C _1767_/B vdd gnd NAND3X1
X_1462_ _1462_/A _1465_/B vdd gnd INVX1
X_1531_ _1911_/Q _1940_/Q _1533_/A vdd gnd NOR2X1
X_1600_ _1722_/B _1648_/B _1601_/B vdd gnd NAND2X1
X_1393_ _1487_/B _1593_/A _1394_/C vdd gnd NOR2X1
X_1729_ _1782_/A _1731_/B vdd gnd INVX1
X_1445_ _1457_/B _1445_/B _1446_/A vdd gnd NOR2X1
X_1514_ _1910_/Q _1940_/Q _1517_/A vdd gnd NOR2X1
X_1376_ _1918_/Q _1487_/A _1453_/B vdd gnd NAND2X1
X_1230_ _1915_/Q _1787_/C vdd gnd INVX2
X_1092_ _1934_/Q _1933_/Q _1109_/B vdd gnd NAND2X1
X_1161_ _1161_/A _1161_/B _1937_/Q _1276_/B vdd gnd OAI21X1
X_1428_ _1649_/B _1733_/B _1790_/A _1757_/B vdd gnd OAI21X1
X_1359_ _1700_/C _1589_/C _1727_/A _1736_/B vdd gnd NAND3X1
X_1213_ _1213_/A _1213_/B _1213_/C _1281_/A vdd gnd AOI21X1
X_1144_ _1144_/A _1144_/B _1144_/C _1158_/C vdd gnd NAND3X1
X_1075_ _1082_/R vdd _1075_/D _1082_/CLK _973_/A vdd gnd DFFSR
X_1831_ _1853_/A _1875_/B _1841_/A vdd gnd AND2X2
X_1900_ _1900_/A _1900_/B _1901_/B vdd gnd NAND2X1
X_1693_ _1728_/A _1728_/B _1710_/A _1694_/C vdd gnd OAI21X1
X_1762_ _1907_/B _1762_/B _1762_/C _1926_/D vdd gnd OAI21X1
X_1058_ _975_/B _1059_/C vdd gnd INVX1
X_1127_ _1127_/A _1127_/B _1137_/B vdd gnd NAND2X1
X_1745_ _1780_/C _1779_/B _1745_/C _1785_/A vdd gnd NAND3X1
X_1814_ _1868_/C _1868_/A _1867_/A _1870_/A vdd gnd OAI21X1
X_1676_ _1700_/C _1700_/B _1700_/A _1766_/B vdd gnd NAND3X1
X_1392_ _1416_/B _1416_/A _1417_/B _1395_/B vdd gnd NAND3X1
X_1461_ _1464_/A _1461_/B _1461_/C _1476_/B vdd gnd OAI21X1
X_1530_ _1723_/A _1907_/A _1530_/C _1535_/B vdd gnd OAI21X1
X_1728_ _1728_/A _1728_/B _1779_/B _1732_/A vdd gnd OAI21X1
X_1659_ _1936_/Q _1935_/Q _1660_/B vdd gnd NOR2X1
X_1375_ _1375_/A _1453_/A vdd gnd INVX1
X_1444_ _1457_/A _1444_/B _1445_/B vdd gnd NAND2X1
X_1513_ _1727_/C _1906_/A _1513_/C _1543_/C vdd gnd OAI21X1
X_1160_ _976_/C _1524_/B vdd gnd INVX1
X_1091_ _1932_/Q _1127_/B _1161_/B vdd gnd NAND2X1
X_1358_ _1406_/A _1371_/C vdd gnd INVX1
X_1427_ _1925_/Q _1790_/A vdd gnd INVX2
X_1289_ _1289_/A _1289_/B _1290_/B vdd gnd NAND2X1
X_1212_ _1216_/B _1216_/A _1213_/C vdd gnd NAND2X1
X_1143_ _1144_/C _1143_/B _1143_/C _1159_/B vdd gnd NAND3X1
X_1074_ _1074_/R vdd _1074_/D _1082_/CLK _949_/A vdd gnd DFFSR
X_1761_ _1761_/A _1774_/C _1764_/A _1762_/B vdd gnd AOI21X1
X_1830_ _1830_/A _1855_/A _1875_/B vdd gnd NOR2X1
X_1692_ _1780_/C _1728_/B vdd gnd INVX1
X_1126_ _1930_/Q _1929_/Q _1931_/Q _1127_/A vdd gnd OAI21X1
X_1057_ _975_/B _1057_/B _1057_/C _1063_/B vdd gnd NAND3X1
X_1744_ _1744_/A _1744_/B _1744_/C _1783_/B vdd gnd AOI21X1
X_1813_ _1930_/Q _1927_/Q _1868_/A vdd gnd NOR2X1
X_1675_ _1675_/A _1675_/B _1921_/Q _1766_/A vdd gnd OAI21X1
X_1109_ _1161_/B _1109_/B _1111_/A _1121_/B vdd gnd OAI21X1
X_1460_ _1460_/A _1460_/B _1460_/C _1461_/C vdd gnd AOI21X1
X_1391_ _1391_/A _1394_/B _1417_/B vdd gnd NOR2X1
X_1658_ _1934_/Q _1933_/Q _1842_/B vdd gnd NOR2X1
X_1727_ _1727_/A _1727_/B _1727_/C _1779_/B vdd gnd OAI21X1
X_1589_ _1722_/C _1790_/A _1589_/C _1590_/B vdd gnd NAND3X1
X_1512_ _1727_/C _1904_/B _1512_/C _1909_/D vdd gnd OAI21X1
X_1374_ _989_/B _1722_/B _1375_/A vdd gnd NAND2X1
X_1443_ _999_/C _1700_/C _1444_/B vdd gnd NAND2X1
X_1090_ _1815_/A _1884_/A _1167_/B _1127_/B vdd gnd NAND3X1
X_1426_ _1482_/B _1787_/B _1434_/A _1787_/D _1433_/A vdd gnd OAI22X1
X_1288_ _1288_/A _1288_/B _1290_/A _1288_/D _1290_/C vdd gnd OAI22X1
X_1357_ _1734_/A _1734_/B _957_/A _1406_/A vdd gnd OAI21X1
X_1142_ _1157_/A _1142_/B _1142_/C _1143_/C vdd gnd AOI21X1
X_1211_ _1211_/A _1211_/B _1216_/B vdd gnd NOR2X1
X_999_ _999_/A _999_/B _999_/C _999_/Y vdd gnd OAI21X1
X_1073_ _1074_/R vdd _1073_/D _1082_/CLK _951_/B vdd gnd DFFSR
X_1409_ _1917_/Q _1918_/Q _1691_/B vdd gnd NAND2X1
X_1760_ _1760_/A _1789_/A _1760_/C _1774_/C vdd gnd AOI21X1
X_1691_ _1909_/Q _1691_/B _1691_/C _1780_/C vdd gnd NAND3X1
X_1125_ _973_/B _1524_/A vdd gnd INVX1
X_1056_ _1059_/A _1057_/B vdd gnd INVX1
X_1889_ _1898_/A _1889_/B _1889_/C _1890_/A vdd gnd NAND3X1
X_1743_ _1743_/A _1781_/B _1781_/A _1744_/B vdd gnd NAND3X1
X_1812_ _1929_/Q _1926_/Q _1868_/C vdd gnd NAND2X1
X_1674_ _1674_/A _1674_/B _1677_/C _1765_/B vdd gnd OAI21X1
X_1039_ _1047_/B _1047_/C _1047_/A _1043_/A vdd gnd OAI21X1
X_1108_ _1291_/B _1161_/B _1824_/A _1111_/A vdd gnd OAI21X1
X_1390_ _1489_/B _1611_/A _1394_/B vdd gnd NOR2X1
X_1588_ _1702_/A _1700_/C _1588_/C _1640_/B vdd gnd NAND3X1
X_1726_ _1731_/A _1782_/C _1726_/C _1785_/B vdd gnd NAND3X1
X_1657_ _1657_/A _1907_/C _1907_/B vdd gnd NAND2X1
X_1511_ _1513_/C _1511_/B _1904_/B _1512_/C vdd gnd NAND3X1
X_1442_ _1921_/Q _1442_/B _1457_/A vdd gnd NAND2X1
X_1373_ _1722_/B _1722_/C _1691_/C vdd gnd NAND2X1
X_1709_ _1780_/A _1709_/B _1745_/C vdd gnd NOR2X1
X_1425_ _1749_/B _1787_/D vdd gnd INVX1
X_1356_ _1922_/Q _1735_/A _1734_/B vdd gnd NOR2X1
X_1287_ _1287_/A _1287_/B _1287_/C _1288_/D vdd gnd OAI21X1
X_1210_ _1210_/A _1210_/B _1211_/B vdd gnd AND2X2
X_998_ _998_/A _998_/B _998_/C _998_/Y vdd gnd OAI21X1
X_1141_ _972_/A _1141_/B _1157_/B _1142_/C vdd gnd OAI21X1
X_1072_ _1074_/R vdd _1072_/D _1082_/CLK _951_/A vdd gnd DFFSR
X_1408_ _1408_/A _1453_/A _1465_/A vdd gnd NOR2X1
X_1339_ _1339_/A _1339_/B _1339_/C _1478_/A vdd gnd NAND3X1
X_1690_ _1780_/A _1728_/A vdd gnd INVX1
X_1055_ _1055_/A _1063_/C _1079_/D vdd gnd NOR2X1
X_1124_ _1161_/B _1146_/A _1141_/B vdd gnd NAND2X1
X_1888_ _1902_/A _1902_/B _1932_/Q _1890_/C vdd gnd OAI21X1
X_1811_ _1930_/Q _1927_/Q _1867_/A vdd gnd NAND2X1
X_1742_ _1911_/Q _1742_/B _1742_/C _1744_/A vdd gnd NAND3X1
X_1673_ _1768_/A _1768_/B _1713_/C vdd gnd NOR2X1
X_1107_ _1933_/Q _1291_/B vdd gnd INVX1
X_1038_ _972_/A _1047_/A vdd gnd INVX1
X_1725_ _1911_/Q _1781_/B _1781_/A _1782_/C vdd gnd NAND3X1
X_1656_ _1757_/C _1656_/B _1656_/C _1657_/A vdd gnd NAND3X1
X_1587_ _1924_/Q _1923_/Q _1588_/C vdd gnd NOR2X1
X_1510_ _1510_/A _1510_/B _1511_/B vdd gnd OR2X2
X_1441_ _1441_/A _1457_/C _1457_/B vdd gnd NAND2X1
X_1372_ _1406_/B _1406_/A _1401_/B vdd gnd AND2X2
X_1708_ _1722_/B _1708_/B _1709_/B vdd gnd NOR2X1
X_1639_ _1639_/A _1639_/B _1923_/D vdd gnd NOR2X1
X_1355_ _1589_/C _1727_/A _1700_/C _1735_/A vdd gnd AOI21X1
X_1424_ _1733_/B _1649_/B _1424_/C _1749_/B vdd gnd OAI21X1
X_1286_ _1932_/Q _1345_/C _1288_/B vdd gnd NOR2X1
X_997_ _997_/A _997_/B _997_/C _998_/A vdd gnd NAND3X1
X_1140_ _1471_/B _1140_/B _1140_/C _1157_/B vdd gnd NAND3X1
X_1071_ vdd _1071_/S _1071_/D _1937_/CLK _950_/A vdd gnd DFFSR
X_1338_ _1338_/A _1338_/B _1338_/C _1338_/D _1339_/B vdd gnd AOI22X1
X_1407_ _989_/B _1722_/B _1408_/A vdd gnd NOR2X1
X_1269_ _1787_/C _1704_/B _1916_/Q _1335_/A vdd gnd OAI21X1
X_1123_ _1818_/A _1123_/B _1146_/A vdd gnd NAND2X1
X_1054_ _1059_/B _1059_/A _1054_/C _1055_/A vdd gnd OAI21X1
X_1887_ _1887_/A _1899_/B _1887_/C _1931_/D vdd gnd OAI21X1
X_1741_ _1741_/A _1782_/A _1744_/C vdd gnd NAND2X1
X_1810_ _1932_/Q _1931_/Q _1928_/Q _1822_/A vdd gnd OAI21X1
X_1672_ _1672_/A _1706_/B _1768_/B vdd gnd NAND2X1
X_1106_ _1934_/Q _1824_/A vdd gnd INVX1
X_1037_ _1037_/A _1063_/C _1076_/D vdd gnd NOR2X1
X_1939_ vdd _1939_/S _1939_/D _1939_/CLK _1939_/Q vdd gnd DFFSR
X_1724_ _1782_/A _1741_/A _1726_/C vdd gnd AND2X2
X_1655_ _1655_/A _1656_/B vdd gnd INVX1
X_1586_ _1586_/A _1586_/B _1916_/D vdd gnd NAND2X1
X_1371_ _1371_/A _1406_/B _1371_/C _1419_/B vdd gnd AOI21X1
X_1440_ _1922_/Q _1440_/B _1457_/C vdd gnd NAND2X1
X_1638_ _1651_/A _1638_/B _1923_/Q _1639_/A vdd gnd AOI21X1
X_1707_ _1769_/B _1769_/A _1707_/C _1796_/B vdd gnd NAND3X1
X_1569_ _1787_/A _1907_/A _1569_/C _1575_/C vdd gnd OAI21X1
X_1354_ _1781_/B _1632_/A _1734_/A vdd gnd AND2X2
X_1285_ _1345_/C _1932_/Q _1285_/C _1290_/A vdd gnd OAI21X1
X_1423_ _1704_/C _1733_/B _1698_/A _1424_/C vdd gnd OAI21X1
X_996_ _996_/A _996_/B _996_/C _997_/B vdd gnd OAI21X1
X_1070_ _1071_/S vdd _1070_/D _1937_/CLK _957_/A vdd gnd DFFSR
X_1406_ _1406_/A _1406_/B _1406_/C _1418_/D vdd gnd NAND3X1
X_1268_ _1914_/Q _1326_/B _1326_/A _1704_/B vdd gnd NAND3X1
X_1337_ _1434_/A _1337_/B _1790_/B _1525_/A _1338_/B vdd gnd AOI22X1
X_1199_ _1199_/A _1199_/B _1199_/C _1214_/B vdd gnd NAND3X1
X_1122_ _1144_/B _1144_/A _1143_/B vdd gnd AND2X2
X_979_ _990_/B _997_/C _981_/A vdd gnd NAND2X1
X_1053_ _972_/B _975_/A _1059_/A vdd gnd NAND2X1
X_1886_ _1892_/B _1886_/B _1887_/A vdd gnd OR2X2
X_1740_ _1740_/A _1778_/A _1740_/C _1784_/A vdd gnd NAND3X1
X_1671_ _1924_/Q _1705_/B _1706_/B vdd gnd NAND2X1
X_1105_ _1343_/A _1165_/C _1472_/B _1793_/B _1166_/A vdd gnd OAI22X1
X_1036_ _1036_/A _1036_/B _1037_/A vdd gnd NAND2X1
X_1869_ _1869_/A _1869_/B _1883_/B vdd gnd NAND2X1
X_1938_ _1939_/S vdd _1938_/D _1939_/CLK _1938_/Q vdd gnd DFFSR
X_1723_ _1723_/A _1723_/B _1723_/C _1741_/A vdd gnd NAND3X1
X_1654_ _1654_/A _1790_/B _1907_/C vdd gnd NOR2X1
X_1585_ _1916_/Q _1585_/B _1586_/A vdd gnd NAND2X1
X_1019_ _976_/B _948_/A _1020_/A vdd gnd NAND2X1
X_1370_ _1440_/B _1733_/B _1733_/C _1406_/B vdd gnd NAND3X1
X_1706_ _1706_/A _1706_/B _1769_/A vdd gnd AND2X2
X_1637_ _1704_/C _1637_/B _1639_/B vdd gnd NOR2X1
X_1499_ _1522_/C _1522_/B _1500_/C vdd gnd AND2X2
X_1568_ _1787_/A _1904_/B _1568_/C _1914_/D vdd gnd OAI21X1
X_1422_ _1924_/Q _1698_/A vdd gnd INVX2
X_1284_ _1284_/A _1291_/D vdd gnd INVX1
X_1353_ _1702_/A _1700_/C _1632_/A vdd gnd NOR2X1
X_995_ _995_/A _995_/B _997_/A vdd gnd NAND2X1
X_1405_ _1420_/B _1429_/C _1749_/C vdd gnd OR2X2
X_1336_ _1705_/B _1337_/B vdd gnd INVX1
X_1267_ _1674_/B _1326_/B vdd gnd INVX1
X_1198_ _1200_/B _1260_/B _1199_/B vdd gnd NAND2X1
XCLKBUF1_insert4 clk _1925_/CLK vdd gnd CLKBUF1
X_978_ _978_/A _978_/B _998_/B vdd gnd NAND2X1
X_1121_ _975_/A _1121_/B _1144_/A vdd gnd NAND2X1
X_1052_ _1052_/A _1059_/B _1052_/C _1054_/C vdd gnd OAI21X1
X_1885_ _1902_/A _1902_/B _1931_/Q _1887_/C vdd gnd OAI21X1
X_1319_ _1734_/C _1700_/B _1677_/C vdd gnd NAND2X1
X_1670_ _1698_/A _1697_/B _1697_/C _1672_/A vdd gnd NAND3X1
X_1035_ _1047_/C _1047_/B _1036_/B vdd gnd OR2X2
X_1104_ _1756_/B _1793_/B vdd gnd INVX1
X_1937_ _1940_/R vdd _1937_/D _1937_/CLK _1937_/Q vdd gnd DFFSR
X_1799_ _1928_/Q _1845_/B vdd gnd INVX2
X_1868_ _1868_/A _1868_/B _1868_/C _1869_/A vdd gnd OAI21X1
X_1584_ _1585_/B _1916_/Q _1586_/B vdd gnd OR2X2
X_1722_ _1919_/Q _1722_/B _1722_/C _1723_/C vdd gnd NAND3X1
X_1653_ _1666_/B _1666_/A _1705_/B _1654_/A vdd gnd OAI21X1
X_1018_ _951_/A _1021_/A vdd gnd INVX1
X_1705_ _1924_/Q _1705_/B _1705_/C _1706_/A vdd gnd OAI21X1
X_1567_ _1904_/B _1567_/B _1569_/C _1568_/C vdd gnd NAND3X1
X_1636_ _1638_/B _1651_/A _1637_/B vdd gnd NAND2X1
X_1498_ _994_/A _994_/B _1522_/B vdd gnd NOR2X1
X_1421_ _1924_/Q _1923_/Q _1649_/B vdd gnd NAND2X1
X_1352_ _1921_/Q _1700_/C vdd gnd INVX2
X_1283_ _972_/A _1818_/A _1284_/A vdd gnd NOR2X1
X_1619_ _1619_/A _1648_/B _1620_/C vdd gnd NAND2X1
X_994_ _994_/A _994_/B _995_/B vdd gnd AND2X2
X_1404_ _1923_/Q _1734_/A _1420_/B vdd gnd NOR2X1
X_1335_ _1335_/A _1335_/B _1790_/B vdd gnd NAND2X1
X_1197_ _1289_/B _1215_/A vdd gnd INVX1
X_1266_ _1913_/Q _1912_/Q _1674_/B vdd gnd NAND2X1
XCLKBUF1_insert5 clk _1939_/CLK vdd gnd CLKBUF1
X_977_ _977_/A _977_/B _977_/C _978_/B vdd gnd OAI21X1
X_1051_ _975_/A _1052_/C vdd gnd INVX1
X_1120_ _1120_/A _1120_/B _1144_/C vdd gnd NAND2X1
X_1884_ _1884_/A _1904_/B _1884_/C _1884_/D _1930_/D vdd gnd OAI22X1
X_1318_ _1911_/Q _1326_/B _1322_/A _1677_/B vdd gnd NAND3X1
X_1249_ _950_/A _1482_/B vdd gnd INVX2
X_1034_ _1047_/B _1047_/C _1036_/A vdd gnd NAND2X1
X_1103_ _1103_/A _1103_/B _1756_/B vdd gnd NAND2X1
X_1867_ _1867_/A _1868_/B vdd gnd INVX1
X_1936_ _1936_/R vdd _1936_/D _1936_/CLK _1936_/Q vdd gnd DFFSR
X_1798_ _1798_/A _1800_/B _1800_/C _1927_/D vdd gnd OAI21X1
X_1721_ _1917_/Q _1918_/Q _1721_/C _1723_/B vdd gnd OAI21X1
X_1652_ _1926_/Q _1762_/C vdd gnd INVX1
X_1583_ _1583_/A _1583_/B _1583_/C _1585_/B vdd gnd OAI21X1
X_1017_ _998_/B _1017_/B _1017_/C _1071_/D vdd gnd OAI21X1
X_1919_ _1925_/R vdd _1919_/D _1925_/CLK _1919_/Q vdd gnd DFFSR
X_1704_ _1704_/A _1704_/B _1704_/C _1705_/C vdd gnd AOI21X1
X_1497_ _989_/A _1497_/B _1522_/C vdd gnd NOR2X1
X_1566_ _1566_/A _1566_/B _1566_/C _1567_/B vdd gnd OAI21X1
X_1635_ _1635_/A _1649_/A _1635_/C _1638_/B vdd gnd OAI21X1
X_1351_ _1922_/Q _1702_/A vdd gnd INVX2
X_1420_ _1429_/C _1420_/B _1787_/B vdd gnd NOR2X1
X_1282_ _975_/A _1824_/A _972_/B _1291_/B _1293_/A vdd gnd OAI22X1
X_1618_ _1618_/A _1650_/B _1618_/C _1619_/A vdd gnd OAI21X1
X_1549_ _1735_/C _1907_/A _1549_/C _1554_/B vdd gnd OAI21X1
X_993_ _999_/A _999_/B _994_/A _998_/C vdd gnd OAI21X1
X_1265_ _1309_/C _1723_/A _1743_/A _1326_/A vdd gnd AOI21X1
X_1403_ _1704_/C _1733_/B _1429_/C vdd gnd NOR2X1
X_1334_ _1334_/A _1334_/B _1338_/A vdd gnd NAND2X1
X_1196_ _1289_/B _1215_/B _1215_/C _1213_/B vdd gnd NAND3X1
XCLKBUF1_insert6 clk _1082_/CLK vdd gnd CLKBUF1
X_976_ _976_/A _976_/B _976_/C _977_/C vdd gnd AOI21X1
X_1050_ _1050_/A _1063_/C _1078_/D vdd gnd NOR2X1
X_1883_ _1903_/A _1883_/B _1884_/C vdd gnd OR2X2
X_1317_ _1317_/A _1317_/B _1317_/C _1329_/B vdd gnd AOI21X1
X_1248_ _1262_/B _1262_/A _1258_/A vdd gnd AND2X2
X_1179_ _989_/A _1727_/C _1191_/A vdd gnd NOR2X1
X_959_ _989_/A _990_/A vdd gnd INVX1
X_1102_ _1109_/B _1161_/B _1845_/A _1103_/A vdd gnd OAI21X1
X_1033_ _973_/B _1047_/B vdd gnd INVX1
X_1797_ _1905_/B _1797_/B _1797_/C _1800_/C vdd gnd NAND3X1
X_1866_ _1867_/A _1866_/B _1866_/C _1869_/B vdd gnd NAND3X1
X_1935_ _1936_/R vdd _1935_/D _1936_/CLK _1935_/Q vdd gnd DFFSR
X_1651_ _1651_/A _1651_/B _1790_/A _1925_/D vdd gnd AOI21X1
X_1720_ _1910_/Q _1720_/B _1720_/C _1782_/A vdd gnd NAND3X1
X_1582_ _1583_/B _1582_/B _1903_/A _1583_/C vdd gnd AOI21X1
X_1016_ _997_/C _1016_/B _1016_/C _1017_/B vdd gnd NAND3X1
X_1849_ _1934_/Q _1933_/Q _1928_/Q _1850_/B vdd gnd OAI21X1
X_1918_ _1925_/R vdd _1918_/D _1925_/CLK _1918_/Q vdd gnd DFFSR
X_1703_ _1703_/A _1771_/A _1771_/B _1769_/B vdd gnd NAND3X1
X_1634_ _1642_/A _1635_/A _1635_/C vdd gnd NAND2X1
X_1565_ _1566_/C _1565_/B _1569_/C vdd gnd OR2X2
X_1496_ _1496_/A _1496_/B _1908_/D vdd gnd NAND2X1
X_1281_ _1281_/A _1281_/B _1281_/C _1339_/A vdd gnd NOR3X1
X_1350_ _1589_/C _1727_/A _1781_/B vdd gnd NAND2X1
X_1617_ _1650_/B _1617_/B _1621_/B _1618_/C vdd gnd NAND3X1
X_1479_ reset _1479_/Y vdd gnd INVX8
X_1548_ _1735_/C _1904_/B _1548_/C _1912_/D vdd gnd OAI21X1
XBUFX2_insert11 _1479_/Y _1936_/R vdd gnd BUFX2
X_992_ _992_/A _998_/B _992_/C _992_/Y vdd gnd OAI21X1
X_1402_ _1923_/Q _1704_/C vdd gnd INVX2
X_1333_ _951_/A _1705_/B _1333_/C _950_/A _1334_/A vdd gnd AOI22X1
X_1264_ _1909_/Q _1908_/Q _1309_/C vdd gnd NOR2X1
X_1195_ _1260_/B _1300_/B _1200_/C _1215_/C vdd gnd OAI21X1
XCLKBUF1_insert7 clk _1083_/CLK vdd gnd CLKBUF1
X_975_ _975_/A _975_/B _976_/A vdd gnd OR2X2
X_1882_ _1901_/A _1882_/B _1884_/D vdd gnd NAND2X1
X_1316_ _994_/A _1681_/A _999_/C _1316_/D _1317_/C vdd gnd OAI22X1
X_1178_ _989_/B _1708_/B _1191_/C vdd gnd NOR2X1
X_1247_ _1253_/B _1247_/B _1262_/A vdd gnd NOR2X1
X_958_ _996_/C _996_/A _958_/C _962_/A vdd gnd NAND3X1
X_1101_ _1101_/A _1103_/B vdd gnd INVX1
X_1032_ _1032_/A _1063_/C _1075_/D vdd gnd NOR2X1
X_1934_ _1936_/R vdd _1934_/D _1936_/CLK _1934_/Q vdd gnd DFFSR
X_1796_ _1796_/A _1796_/B _1796_/C _1797_/C vdd gnd AOI21X1
X_1865_ _1868_/A _1866_/B vdd gnd INVX1
X_1650_ _1650_/A _1650_/B _1650_/C _1651_/B vdd gnd AOI21X1
X_1581_ _1940_/Q _1656_/C _1582_/B vdd gnd NAND2X1
X_1015_ _1015_/A _1015_/B _952_/A _1016_/B vdd gnd OAI21X1
X_1917_ _1925_/R vdd _1917_/D _1925_/CLK _1917_/Q vdd gnd DFFSR
X_1779_ _1780_/C _1779_/B _1780_/B vdd gnd NAND2X1
X_1848_ _1848_/A _1848_/B _1848_/C _1851_/B vdd gnd OAI21X1
X_1564_ _1578_/B _1565_/B vdd gnd INVX1
X_1633_ _1922_/Q _1736_/B _1642_/A vdd gnd NOR2X1
X_1702_ _1702_/A _1702_/B _1702_/C _1703_/A vdd gnd OAI21X1
X_1495_ _1708_/B _1938_/Q _1898_/A _1496_/A vdd gnd NAND3X1
X_1280_ _1280_/A _1280_/B _1280_/C _1281_/C vdd gnd OAI21X1
X_1547_ _1904_/B _1549_/C _1547_/C _1548_/C vdd gnd NAND3X1
X_1616_ _1721_/C _1691_/B _1682_/A _1617_/B vdd gnd OAI21X1
X_1478_ _1478_/A _1478_/B _1478_/C _1943_/A vdd gnd AOI21X1
XBUFX2_insert12 _1479_/Y _1939_/S vdd gnd BUFX2
X_991_ _991_/A _991_/B _997_/C _992_/A vdd gnd NAND3X1
X_1401_ _1406_/C _1401_/B _1401_/C _1419_/A vdd gnd NAND3X1
X_1263_ _1525_/A _1916_/Q _1263_/C _1263_/D _1280_/A vdd gnd OAI22X1
X_1194_ _1199_/A _1199_/C _1200_/C vdd gnd NAND2X1
X_1332_ _1697_/B _1697_/C _1705_/B vdd gnd NAND2X1
XCLKBUF1_insert8 clk _1937_/CLK vdd gnd CLKBUF1
X_974_ _974_/A _974_/B _977_/B vdd gnd AND2X2
X_1881_ _1881_/A _1899_/B _1881_/C _1929_/D vdd gnd OAI21X1
X_1315_ _1700_/B _1700_/A _1316_/D vdd gnd NAND2X1
X_1177_ _1908_/Q _1708_/B vdd gnd INVX2
X_1246_ _1253_/A _1246_/B _1247_/B vdd gnd NAND2X1
X_957_ _957_/A _999_/C _958_/C vdd gnd NOR2X1
X_1100_ _1163_/B _1100_/B _1165_/C vdd gnd NOR2X1
X_1031_ _1047_/C _1031_/B _1032_/A vdd gnd NAND2X1
X_1933_ _1936_/R vdd _1933_/D _1936_/CLK _1933_/Q vdd gnd DFFSR
X_1864_ _1866_/C _1864_/B _1880_/B vdd gnd OR2X2
X_1795_ _1795_/A _1795_/B _1795_/C _1796_/C vdd gnd OAI21X1
X_1229_ _1914_/Q _1787_/A vdd gnd INVX4
X_1580_ _1580_/A _1580_/B _1656_/C vdd gnd NOR2X1
X_1014_ _950_/A _957_/A _1014_/C _1016_/C vdd gnd NAND3X1
X_1847_ _1900_/B _1900_/A _1882_/B vdd gnd AND2X2
X_1916_ _1940_/R vdd _1916_/D _1937_/CLK _1916_/Q vdd gnd DFFSR
X_1778_ _1778_/A _1778_/B _1784_/C vdd gnd NAND2X1
X_1701_ _1701_/A _1767_/B _1702_/C vdd gnd NAND2X1
X_1563_ _1566_/A _1566_/B _1578_/B vdd gnd NOR2X1
X_1632_ _1632_/A _1632_/B _1649_/A vdd gnd NAND2X1
X_1494_ _1905_/A _1892_/B _1908_/Q _1496_/B vdd gnd OAI21X1
X_1546_ _1578_/C _1546_/B _1547_/C vdd gnd OR2X2
X_1477_ _1477_/A _1477_/B _1477_/C _1478_/B vdd gnd AOI21X1
X_1615_ _1632_/B _1621_/B vdd gnd INVX1
XBUFX2_insert13 _1479_/Y _1924_/R vdd gnd BUFX2
X_990_ _990_/A _990_/B _996_/A _991_/B vdd gnd OAI21X1
X_1400_ _1400_/A _1400_/B _1406_/C vdd gnd AND2X2
X_1331_ _1787_/A _1677_/B _1787_/C _1697_/C vdd gnd OAI21X1
X_1193_ _1199_/A _1199_/C _1306_/C _1215_/B vdd gnd NAND3X1
X_1262_ _1262_/A _1262_/B _1263_/D vdd gnd NAND2X1
X_1529_ _1903_/A _1602_/B vdd gnd INVX1
X_973_ _973_/A _973_/B _974_/B vdd gnd NOR2X1
XCLKBUF1_insert9 clk _1940_/CLK vdd gnd CLKBUF1
X_1880_ _1892_/B _1880_/B _1881_/A vdd gnd OR2X2
X_1314_ _1743_/A _1321_/C _1735_/C _1700_/A vdd gnd OAI21X1
X_1176_ _989_/A _1727_/C _1190_/A vdd gnd NAND2X1
X_1245_ _999_/C _1735_/C _1246_/B vdd gnd NAND2X1
X_956_ _994_/B _996_/A vdd gnd INVX1
X_1030_ _949_/A _973_/A _978_/A _1047_/C vdd gnd NAND3X1
X_1863_ _1929_/Q _1926_/Q _1864_/B vdd gnd NOR2X1
X_1932_ _1936_/R vdd _1932_/D _1936_/CLK _1932_/Q vdd gnd DFFSR
X_1794_ _1794_/A _1794_/B _1794_/C _1795_/C vdd gnd NOR3X1
X_1228_ _1228_/A _1228_/B _1228_/C _1258_/B vdd gnd OAI21X1
X_1159_ _1159_/A _1159_/B _1159_/C _1166_/B vdd gnd AOI21X1
X_1013_ _996_/C _1013_/B _991_/A _1014_/C vdd gnd NOR3X1
X_1777_ _1777_/A _1777_/B _1796_/A vdd gnd AND2X2
X_1846_ _1846_/A _1846_/B _1900_/B vdd gnd NAND2X1
X_1915_ _1940_/R vdd _1915_/D _1940_/CLK _1915_/Q vdd gnd DFFSR
X_1700_ _1700_/A _1700_/B _1700_/C _1701_/A vdd gnd AOI21X1
X_1631_ _1631_/A _1631_/B _1922_/D vdd gnd NAND2X1
X_1493_ _1898_/A _1892_/B vdd gnd INVX1
X_1562_ _1787_/A _1907_/A _1566_/B vdd gnd NOR2X1
X_1829_ _1933_/Q _1928_/Q _1830_/A vdd gnd NOR2X1
X_1614_ _1682_/A _1614_/B _1632_/B vdd gnd NOR2X1
X_1476_ _1476_/A _1476_/B _1476_/C _1477_/B vdd gnd AOI21X1
X_1545_ _1546_/B _1578_/C _1549_/C vdd gnd NAND2X1
XBUFX2_insert14 _1479_/Y _1940_/R vdd gnd BUFX2
X_1261_ _1261_/A _1261_/B _1261_/C _1263_/C vdd gnd NAND3X1
X_1330_ _1330_/A _1333_/C vdd gnd INVX1
X_1192_ _1192_/A _1200_/B _1260_/B _1306_/C vdd gnd NAND3X1
X_1528_ _1528_/A _1528_/B _1903_/A vdd gnd OR2X2
X_1459_ _951_/A _1698_/A _1459_/C _1460_/C vdd gnd OAI21X1
X_972_ _972_/A _972_/B _974_/A vdd gnd NOR2X1
X_1313_ _1910_/Q _1909_/Q _1908_/Q _1321_/C vdd gnd NOR3X1
X_1244_ _1912_/Q _1735_/C vdd gnd INVX2
X_1175_ _1909_/Q _1727_/C vdd gnd INVX2
X_955_ _994_/A _996_/C vdd gnd INVX1
X_1862_ _1868_/C _1866_/C vdd gnd INVX1
X_1793_ _1793_/A _1793_/B _1793_/C _1794_/C vdd gnd NAND3X1
X_1931_ _1936_/R vdd _1931_/D _1936_/CLK _1931_/Q vdd gnd DFFSR
X_1158_ _975_/B _1756_/B _1158_/C _1158_/D _1159_/C vdd gnd OAI22X1
X_1227_ _1227_/A _1227_/B _1228_/C vdd gnd NOR2X1
X_1089_ _1929_/Q _1167_/B vdd gnd INVX1
X_1012_ _999_/A _999_/B _950_/A _1017_/C vdd gnd OAI21X1
X_1914_ _1924_/R vdd _1914_/D _1940_/CLK _1914_/Q vdd gnd DFFSR
X_1776_ _1907_/B _1905_/B vdd gnd INVX1
X_1845_ _1845_/A _1845_/B _1845_/C _1846_/B vdd gnd OAI21X1
X_1630_ _1702_/A _1630_/B _1651_/A _1631_/A vdd gnd NAND3X1
X_1492_ _1492_/A _1492_/B _1898_/A vdd gnd NOR2X1
X_1561_ _1914_/Q _1940_/Q _1566_/A vdd gnd NOR2X1
X_1828_ _1853_/B _1855_/A vdd gnd INVX1
X_1759_ _1759_/A _1759_/B _1759_/C _1760_/C vdd gnd NAND3X1
X_1544_ _1544_/A _1544_/B _1578_/C vdd gnd NAND2X1
X_1613_ _1613_/A _1613_/B _1613_/C _1919_/D vdd gnd OAI21X1
X_1475_ _1525_/A _1751_/C _1475_/C _1476_/C vdd gnd OAI21X1
XBUFX2_insert15 _1479_/Y _1925_/R vdd gnd BUFX2
X_1260_ _1300_/B _1260_/B _1261_/C vdd gnd NOR2X1
X_1191_ _1191_/A _1191_/B _1191_/C _1200_/B vdd gnd OAI21X1
X_1527_ _1527_/A _1527_/B _1528_/A vdd gnd NAND2X1
X_1458_ _1482_/B _1923_/Q _1458_/C _1459_/C vdd gnd NAND3X1
X_1389_ _1720_/B _1720_/C _1611_/A vdd gnd NAND2X1
X_971_ _976_/B _971_/B _971_/C _977_/A vdd gnd NAND3X1
X_1312_ _1912_/Q _1911_/Q _1322_/A _1700_/B vdd gnd NAND3X1
X_1174_ _1174_/A _1261_/A vdd gnd INVX1
X_1243_ _1912_/Q _1442_/B _1253_/A vdd gnd NAND2X1
X_954_ _999_/B _954_/B _954_/Y vdd gnd AND2X2
X_1930_ _1936_/R vdd _1930_/D _1936_/CLK _1930_/Q vdd gnd DFFSR
X_1792_ _1792_/A _1793_/A vdd gnd INVX1
X_1861_ _1861_/A _1861_/B _1889_/B vdd gnd NAND2X1
X_1157_ _1157_/A _1157_/B _1157_/C _1158_/D vdd gnd NAND3X1
X_1226_ _1226_/A _1226_/B _1227_/B vdd gnd NOR2X1
X_1088_ _1930_/Q _1884_/A vdd gnd INVX1
X_1011_ _1011_/A _998_/B _1011_/C _1070_/D vdd gnd OAI21X1
X_1913_ _1924_/R vdd _1913_/D _1940_/CLK _1913_/Q vdd gnd DFFSR
X_1775_ _1775_/A _1797_/B _1907_/B _1800_/B vdd gnd AOI21X1
X_1844_ _1844_/A _1844_/B _1845_/C _1900_/A vdd gnd NAND3X1
X_1209_ _1209_/A _1209_/B _1216_/A vdd gnd NAND2X1
X_1560_ _1940_/Q _1580_/B _1578_/C _1578_/A _1566_/C vdd gnd AOI22X1
X_1491_ _1527_/A _1491_/B _1492_/B vdd gnd NAND2X1
X_1827_ _1933_/Q _1928_/Q _1853_/B vdd gnd NAND2X1
X_1758_ _1794_/B _1759_/A vdd gnd INVX1
X_1689_ _1917_/Q _1908_/Q _1780_/A vdd gnd NOR2X1
X_1543_ _1543_/A _1543_/B _1543_/C _1544_/B vdd gnd NAND3X1
X_1474_ _1474_/A _1474_/B _1475_/C vdd gnd NOR2X1
X_1612_ _1919_/Q _1613_/A _1613_/C vdd gnd NAND2X1
X_1190_ _1190_/A _1191_/B vdd gnd INVX1
X_1526_ _1526_/A _1526_/B _1527_/B vdd gnd NOR2X1
X_1457_ _1457_/A _1457_/B _1457_/C _1460_/B vdd gnd OAI21X1
X_1388_ _1720_/C _1720_/B _994_/B _1391_/A vdd gnd AOI21X1
X_970_ _976_/C _971_/B vdd gnd INVX1
X_1311_ _994_/B _1680_/B _1681_/A _994_/A _1317_/B vdd gnd AOI22X1
X_1242_ _999_/C _1442_/B vdd gnd INVX1
X_1173_ _1173_/A _1226_/A _1174_/A vdd gnd NAND2X1
X_1509_ _1510_/B _1510_/A _1513_/C vdd gnd NAND2X1
X_953_ _963_/A _966_/A _954_/B vdd gnd NOR2X1
X_1860_ _1861_/B _1861_/A _1889_/C vdd gnd OR2X2
X_1791_ _1791_/A _1793_/C vdd gnd INVX1
X_1156_ _1345_/C _1755_/B _1156_/C _1157_/C vdd gnd AOI21X1
X_1087_ _1931_/Q _1815_/A vdd gnd INVX1
X_1225_ _1487_/A _1909_/Q _1225_/C _1228_/A vdd gnd OAI21X1
X_1010_ _1010_/A _1010_/B _997_/C _1011_/A vdd gnd NAND3X1
X_1843_ _1850_/A _1848_/C _1845_/C vdd gnd NAND2X1
X_1912_ _1924_/R vdd _1912_/D _1940_/CLK _1912_/Q vdd gnd DFFSR
X_1774_ _1774_/A _1774_/B _1774_/C _1775_/A vdd gnd OAI21X1
X_1208_ _1208_/A _1211_/A _1208_/C _1209_/A vdd gnd OAI21X1
X_1139_ _972_/B _1471_/B vdd gnd INVX1
X_1490_ _1490_/A _1490_/B _1491_/B vdd gnd NOR2X1
X_1826_ _1855_/C _1853_/A vdd gnd INVX1
X_1757_ _1757_/A _1757_/B _1757_/C _1794_/B vdd gnd AOI21X1
X_1688_ _1722_/C _1711_/B _1710_/A vdd gnd NAND2X1
X_1611_ _1611_/A _1650_/B _1611_/C _1613_/B vdd gnd OAI21X1
X_1473_ _1473_/A _1473_/B _1473_/C _1474_/B vdd gnd NAND3X1
X_1542_ _1911_/Q _1910_/Q _1940_/Q _1544_/A vdd gnd OAI21X1
X_1809_ _1846_/A _1840_/A _1832_/A vdd gnd NOR2X1
X_1525_ _1525_/A _1525_/B _1525_/C _1526_/B vdd gnd NAND3X1
X_1456_ _1463_/C _1456_/B _1456_/C _1461_/B vdd gnd AOI21X1
X_1387_ _1917_/Q _1918_/Q _1919_/Q _1720_/B vdd gnd OAI21X1
X_1241_ _1241_/A _1241_/B _1253_/B vdd gnd NAND2X1
X_1310_ _1655_/A _1674_/A _1681_/A vdd gnd NAND2X1
X_1172_ _1910_/Q _1489_/B _1226_/A vdd gnd NAND2X1
X_1439_ _957_/A _1702_/A _1441_/A vdd gnd NAND2X1
X_1508_ _1508_/A _1508_/B _1510_/A vdd gnd NAND2X1
X_952_ _952_/A _961_/C _966_/A vdd gnd NAND2X1
X_1790_ _1790_/A _1790_/B _1794_/A vdd gnd NOR2X1
X_1224_ _989_/A _1727_/C _1300_/B _1225_/C vdd gnd OAI21X1
X_1155_ _1155_/A _1155_/B _1206_/C _1156_/C vdd gnd NAND3X1
X_1086_ _975_/B _1472_/B vdd gnd INVX1
X_1773_ _1773_/A _1773_/B _1777_/B _1774_/A vdd gnd OAI21X1
X_1842_ _1845_/B _1842_/B _1850_/C _1848_/C vdd gnd OAI21X1
X_1911_ _1924_/R vdd _1911_/D _1940_/CLK _1911_/Q vdd gnd DFFSR
X_1207_ _1210_/B _1210_/A _1211_/A vdd gnd NOR2X1
X_1138_ _1340_/B _1138_/B _1155_/A _1142_/B vdd gnd OAI21X1
X_1069_ _1074_/R vdd _1069_/D _1082_/CLK _999_/C vdd gnd DFFSR
X_1756_ _1792_/A _1756_/B _1791_/A _1759_/C vdd gnd NOR3X1
X_1825_ _1825_/A _1825_/B _1855_/C vdd gnd NAND2X1
X_1687_ _1687_/A _1687_/B _1711_/B vdd gnd NAND2X1
X_1610_ _1610_/A _1610_/B _1650_/B _1611_/C vdd gnd OAI21X1
X_1541_ _1557_/B _1546_/B vdd gnd INVX1
X_1472_ _976_/C _1472_/B _1473_/B vdd gnd NOR2X1
X_1808_ _1848_/A _1848_/B _1840_/A vdd gnd OR2X2
X_1739_ _1739_/A _1739_/B _1740_/C vdd gnd NAND2X1
X_1524_ _1524_/A _1524_/B _1524_/C _1526_/A vdd gnd NAND3X1
X_1386_ _994_/A _1618_/A _1416_/A vdd gnd NAND2X1
X_1455_ _994_/A _1682_/A _1455_/C _1456_/C vdd gnd OAI21X1
X_1171_ _994_/B _1489_/B vdd gnd INVX1
X_1240_ _957_/A _1734_/C _1241_/B vdd gnd NAND2X1
X_1507_ _1939_/Q _1727_/C _1508_/B vdd gnd NAND2X1
X_1438_ _950_/A _1704_/C _1438_/C _1460_/A vdd gnd AOI21X1
X_1369_ _1702_/A _1736_/C _1733_/C vdd gnd NAND2X1
X_951_ _951_/A _951_/B _961_/C vdd gnd NOR2X1
X_1223_ _1261_/B _1261_/A _1228_/B vdd gnd NAND2X1
X_1154_ _1154_/A _1929_/Q _1210_/A _1155_/B vdd gnd OAI21X1
X_1085_ _976_/B _1343_/A vdd gnd INVX1
X_1910_ _1940_/R vdd _1910_/D _1939_/CLK _1910_/Q vdd gnd DFFSR
X_1772_ _1772_/A _1773_/B vdd gnd INVX1
X_1841_ _1841_/A _1875_/A _1850_/C vdd gnd NAND2X1
X_1206_ _1287_/C _1285_/C _1206_/C _1209_/B vdd gnd NAND3X1
X_1137_ _1524_/A _1137_/B _1155_/A vdd gnd NAND2X1
X_1068_ _1071_/S vdd _998_/Y _1937_/CLK _994_/A vdd gnd DFFSR
X_1686_ _1909_/Q _1908_/Q _1687_/A vdd gnd NAND2X1
X_1755_ _1755_/A _1755_/B _1792_/A vdd gnd NAND2X1
X_1824_ _1824_/A _1845_/B _1825_/B vdd gnd NAND2X1
X_1540_ _1540_/A _1540_/B _1557_/B vdd gnd OR2X2
X_1471_ _976_/B _1471_/B _1473_/A vdd gnd NOR2X1
X_1807_ _1935_/Q _1928_/Q _1848_/B vdd gnd NOR2X1
X_1738_ _1778_/A _1778_/B _1786_/D _1738_/D _1750_/B vdd gnd AOI22X1
X_1669_ _1696_/B _1696_/A _1768_/A vdd gnd NAND2X1
X_1454_ _1489_/B _1919_/Q _1454_/C _1455_/C vdd gnd NAND3X1
X_1523_ _949_/A _972_/A _1524_/C vdd gnd NOR2X1
X_1385_ _1742_/B _1742_/C _1618_/A vdd gnd NAND2X1
X_1170_ _994_/B _1723_/A _1173_/A vdd gnd NAND2X1
X_1506_ _1909_/Q _1906_/A _1508_/A vdd gnd NAND2X1
X_1437_ _950_/A _1704_/C _1458_/C _1438_/C vdd gnd OAI21X1
X_1368_ _1735_/A _1736_/C vdd gnd INVX1
X_1299_ _1727_/C _1708_/B _1687_/B vdd gnd NAND2X1
X_950_ _950_/A _952_/A vdd gnd INVX1
X_1084_ _964_/Y _1478_/C vdd gnd INVX1
X_1222_ _1226_/B _1227_/A _1261_/B vdd gnd NOR2X1
X_1153_ _1153_/A _1287_/C _1210_/A vdd gnd NAND2X1
X_1840_ _1840_/A _1850_/A vdd gnd INVX1
X_1771_ _1771_/A _1771_/B _1771_/C _1773_/A vdd gnd NAND3X1
X_1205_ _1208_/C _1285_/C vdd gnd INVX1
X_1136_ _1884_/A _1167_/B _1287_/B _1287_/A _1138_/B vdd gnd AOI22X1
X_1067_ _1071_/S vdd _992_/Y _1082_/CLK _994_/B vdd gnd DFFSR
X_1823_ _1934_/Q _1928_/Q _1825_/A vdd gnd NAND2X1
X_1754_ _1815_/A _1754_/B _1754_/C _1755_/A vdd gnd AOI21X1
X_1685_ _1694_/A _1685_/B _1685_/C _1712_/B vdd gnd NAND3X1
X_1119_ _975_/A _1121_/B _1119_/C _1159_/A vdd gnd AOI21X1
X_1470_ _973_/A _973_/B _1470_/C _1474_/A vdd gnd OAI21X1
X_1806_ _1844_/B _1848_/A vdd gnd INVX1
X_1737_ _1739_/B _1739_/A _1737_/C _1737_/D _1786_/D vdd gnd AOI22X1
X_1599_ _1613_/A _1648_/B vdd gnd INVX2
X_1668_ _1704_/C _1704_/B _1704_/A _1696_/B vdd gnd NAND3X1
X_1522_ _1522_/A _1522_/B _1522_/C _1528_/B vdd gnd NAND3X1
X_1453_ _1453_/A _1453_/B _1462_/A _1456_/B vdd gnd AOI21X1
X_1384_ _1920_/Q _1721_/C _1727_/A _1742_/B vdd gnd NAND3X1
X_1505_ _1939_/Q _1906_/A vdd gnd INVX1
X_1436_ _1436_/A _1436_/B _1458_/C vdd gnd NAND2X1
X_1367_ _1920_/Q _1720_/C _1632_/A _1733_/B vdd gnd OAI21X1
X_1298_ _1803_/A _976_/B _976_/C _1904_/A _1338_/D vdd gnd AOI22X1
X_1221_ _994_/A _1743_/A _1227_/A vdd gnd NOR2X1
X_1152_ _973_/A _1884_/A _1287_/C vdd gnd NAND2X1
X_1083_ _1083_/R vdd _968_/Y _1083_/CLK _978_/A vdd gnd DFFSR
X_1419_ _1419_/A _1419_/B _1419_/C _1433_/B vdd gnd AOI21X1
X_1770_ _1770_/A _1770_/B _1770_/C _1774_/B vdd gnd AOI21X1
X_1204_ _1288_/A _1204_/B _1208_/C vdd gnd NAND2X1
X_1135_ _1168_/A _1287_/B vdd gnd INVX1
X_1066_ _1074_/R vdd _987_/Y _1082_/CLK _989_/A vdd gnd DFFSR
X_1899_ _1899_/A _1899_/B _1899_/C _1935_/D vdd gnd OAI21X1
X_1753_ _1803_/A _1753_/B _1754_/C vdd gnd NAND2X1
X_1822_ _1822_/A _1822_/B _1875_/A vdd gnd NAND2X1
X_1684_ _1721_/C _1684_/B _1685_/B vdd gnd NAND2X1
X_1118_ _1120_/A _1120_/B _1144_/B _1119_/C vdd gnd AOI21X1
X_1049_ _1049_/A _1049_/B _1050_/A vdd gnd NAND2X1
X_1736_ _1912_/Q _1736_/B _1736_/C _1739_/A vdd gnd NAND3X1
X_1805_ _1935_/Q _1928_/Q _1844_/B vdd gnd NAND2X1
X_1598_ _1917_/Q _1613_/A _1601_/A vdd gnd NAND2X1
X_1667_ _1674_/B _1674_/A _1787_/A _1704_/A vdd gnd OAI21X1
X_1452_ _1918_/Q _1487_/A _1462_/A vdd gnd NOR2X1
X_1383_ _1919_/Q _1691_/C _1682_/A _1742_/C vdd gnd OAI21X1
X_1521_ _1723_/A _1904_/B _1521_/C _1910_/D vdd gnd OAI21X1
X_1719_ _1743_/A _1742_/B _1742_/C _1731_/A vdd gnd NAND3X1
X_1504_ _1708_/B _1905_/A _1510_/B vdd gnd NOR2X1
X_1366_ _1721_/C _1722_/B _1722_/C _1720_/C vdd gnd NAND3X1
X_1435_ _951_/A _1924_/Q _1436_/A vdd gnd NAND2X1
X_1297_ _1297_/A _1297_/B _1338_/C vdd gnd NAND2X1
X_1220_ _1911_/Q _1743_/A vdd gnd INVX2
X_1151_ _1930_/Q _1525_/B _1153_/A vdd gnd NAND2X1
X_1082_ _1082_/R vdd _1082_/D _1082_/CLK _976_/C vdd gnd DFFSR
X_1418_ _950_/A _1749_/C _1418_/C _1418_/D _1419_/C vdd gnd OAI22X1
X_1349_ _1917_/Q _1918_/Q _1727_/A vdd gnd NOR2X1
X_1134_ _1929_/Q _1154_/A _1168_/A vdd gnd NOR2X1
X_1203_ _973_/B _1815_/A _1204_/B vdd gnd NAND2X1
X_1065_ _1071_/S vdd _981_/Y _1937_/CLK _989_/B vdd gnd DFFSR
X_1898_ _1898_/A _1898_/B _1899_/A vdd gnd NAND2X1
X_1752_ _1790_/B _1790_/A _1759_/B vdd gnd OR2X2
X_1683_ _1685_/C _1694_/B vdd gnd INVX1
X_1821_ _1870_/A _1870_/B _1861_/A _1822_/B vdd gnd NAND3X1
X_1117_ _972_/B _1117_/B _1144_/B vdd gnd NAND2X1
X_1048_ _972_/B _1057_/C _1049_/B vdd gnd NAND2X1
X_1804_ _1804_/A _1804_/B _1846_/A vdd gnd NAND2X1
X_1666_ _1666_/A _1666_/B _1923_/Q _1696_/A vdd gnd OAI21X1
X_1735_ _1735_/A _1735_/B _1735_/C _1739_/B vdd gnd OAI21X1
X_1597_ _1904_/B _1602_/A _1613_/A vdd gnd NAND2X1
X_1520_ _1904_/B _1530_/C _1520_/C _1521_/C vdd gnd NAND3X1
X_1451_ _994_/B _1721_/C _1451_/C _1463_/C vdd gnd AOI21X1
X_1382_ _1920_/Q _1682_/A vdd gnd INVX2
X_1649_ _1649_/A _1649_/B _1650_/A vdd gnd OR2X2
X_1718_ _1735_/C _1718_/B _1740_/A _1778_/B vdd gnd OAI21X1
X_1503_ _1902_/A _1902_/B _1904_/B vdd gnd NOR2X1
X_1296_ _1472_/B _1935_/Q _1296_/C _1297_/A vdd gnd AOI21X1
X_1365_ _1918_/Q _1722_/C vdd gnd INVX2
X_1434_ _1434_/A _1698_/A _1436_/B vdd gnd NAND2X1
X_1150_ _949_/A _1167_/B _1289_/A _1206_/C vdd gnd OAI21X1
X_1081_ vdd _1083_/R _1081_/D _1083_/CLK _976_/B vdd gnd DFFSR
X_1417_ _1417_/A _1417_/B _1417_/C _1418_/C vdd gnd NAND3X1
X_1279_ _1279_/A _1280_/C vdd gnd INVX1
X_1348_ _1920_/Q _1919_/Q _1589_/C vdd gnd NOR2X1
X_1133_ _949_/A _1154_/A vdd gnd INVX1
X_1064_ _978_/A _971_/B _1082_/D vdd gnd NOR2X1
X_1202_ _1931_/Q _1524_/A _1288_/A vdd gnd NAND2X1
X_1897_ _1902_/A _1902_/B _1935_/Q _1899_/C vdd gnd OAI21X1
X_1820_ _1820_/A _1820_/B _1861_/A vdd gnd NOR2X1
X_1751_ _1787_/C _1787_/D _1751_/C _1757_/C _1789_/A vdd gnd AOI22X1
X_1682_ _1682_/A _1682_/B _1685_/C vdd gnd NAND2X1
X_1047_ _1047_/A _1047_/B _1047_/C _1057_/C vdd gnd NOR3X1
X_1116_ _1140_/B _1140_/C _1117_/B vdd gnd NAND2X1
X_1803_ _1803_/A _1845_/B _1804_/B vdd gnd NAND2X1
X_1665_ _1833_/A _1665_/B _1764_/A vdd gnd NOR2X1
X_1596_ _1751_/C _1596_/B _1650_/B _1602_/A vdd gnd OAI21X1
X_1734_ _1734_/A _1734_/B _1734_/C _1737_/D vdd gnd OAI21X1
X_1450_ _994_/B _1721_/C _1454_/C _1451_/C vdd gnd OAI21X1
X_1381_ _1487_/B _1593_/A _1416_/B vdd gnd NAND2X1
X_1579_ _1787_/C _1787_/A _1580_/A vdd gnd NAND2X1
X_1648_ _1698_/A _1648_/B _1648_/C _1924_/D vdd gnd OAI21X1
X_1717_ _1734_/A _1734_/B _1913_/Q _1740_/A vdd gnd OAI21X1
X_1502_ _1524_/B _1502_/B _1527_/A _1902_/A vdd gnd NAND3X1
X_1433_ _1433_/A _1433_/B _1433_/C _1477_/A vdd gnd OAI21X1
X_1364_ _1917_/Q _1722_/B vdd gnd INVX2
X_1295_ _976_/B _1803_/A _1296_/C vdd gnd NOR2X1
X_1080_ _1082_/R vdd _1080_/D _1083_/CLK _975_/B vdd gnd DFFSR
X_1416_ _1416_/A _1416_/B _1417_/C vdd gnd AND2X2
X_1347_ _1347_/A _1347_/B _1477_/C vdd gnd NOR2X1
X_1278_ _1278_/A _1278_/B _1278_/C _1279_/A vdd gnd NAND3X1
X_1201_ _1215_/A _1214_/B _1214_/C _1213_/A vdd gnd NAND3X1
X_989_ _989_/A _989_/B _994_/B _991_/A vdd gnd NAND3X1
X_1063_ _1063_/A _1063_/B _1063_/C _1081_/D vdd gnd AOI21X1
X_1132_ _973_/A _1884_/A _1287_/A vdd gnd NOR2X1
X_1896_ _1896_/A _1899_/B _1896_/C _1934_/D vdd gnd OAI21X1
X_1750_ _1750_/A _1750_/B _1750_/C _1760_/A vdd gnd OAI21X1
X_1681_ _1681_/A _1682_/B vdd gnd INVX1
X_1046_ _1052_/A _1059_/B _1049_/A vdd gnd NAND2X1
X_1115_ _1818_/A _1123_/B _1291_/B _1140_/B vdd gnd OAI21X1
X_1879_ _1901_/C _1882_/B _1901_/A _1899_/B vdd gnd OAI21X1
X_1733_ _1913_/Q _1733_/B _1733_/C _1737_/C vdd gnd NAND3X1
X_1802_ _1936_/Q _1928_/Q _1804_/A vdd gnd NAND2X1
X_1595_ down _1749_/C _1595_/C _1596_/B vdd gnd NAND3X1
X_1664_ _1754_/B _1664_/B _1904_/A _1665_/B vdd gnd OAI21X1
X_1029_ _1029_/A _999_/A _1029_/C _1031_/B vdd gnd OAI21X1
X_1380_ _1781_/B _1781_/A _1593_/A vdd gnd NAND2X1
X_1716_ _1734_/C _1733_/B _1733_/C _1778_/A vdd gnd NAND3X1
X_1578_ _1578_/A _1578_/B _1578_/C _1583_/B vdd gnd NAND3X1
X_1647_ _1647_/A _1648_/B _1648_/C vdd gnd NAND2X1
X_1432_ _1434_/A _1787_/D _1751_/C _1525_/A _1433_/C vdd gnd AOI22X1
X_1363_ _1919_/Q _1721_/C vdd gnd INVX2
X_1501_ _1501_/A _1501_/B _1502_/B vdd gnd AND2X2
X_1294_ _1936_/Q _1803_/A vdd gnd INVX1
X_1415_ _1415_/A _1415_/B _1465_/A _1417_/A vdd gnd AOI21X1
X_1346_ _1346_/A _1527_/A _1347_/B vdd gnd NAND2X1
X_1277_ _1525_/A _1916_/Q _1524_/B _1937_/Q _1278_/B vdd gnd AOI22X1
X_1200_ _1260_/B _1200_/B _1200_/C _1214_/C vdd gnd NAND3X1
X_988_ _999_/A _999_/B _994_/B _992_/C vdd gnd OAI21X1
X_1131_ _1131_/A _1340_/B vdd gnd INVX1
X_1062_ _976_/B _1063_/A vdd gnd INVX1
X_1895_ _1898_/A _1895_/B _1896_/A vdd gnd NAND2X1
X_1329_ _1329_/A _1329_/B _1329_/C _1334_/B vdd gnd OAI21X1
X_1680_ _1919_/Q _1680_/B _1681_/A _1920_/Q _1694_/A vdd gnd AOI22X1
X_1114_ _1127_/B _1123_/B vdd gnd INVX1
X_1045_ _972_/B _1052_/A vdd gnd INVX1
X_1878_ _1878_/A _1898_/B _1895_/B _1901_/C vdd gnd NOR3X1
X_1663_ _1930_/Q _1929_/Q _1754_/B vdd gnd NAND2X1
X_1732_ _1732_/A _1785_/B _1732_/C _1738_/D vdd gnd OAI21X1
X_1801_ _1902_/A _1902_/B _1929_/Q _1881_/C vdd gnd OAI21X1
X_1594_ _1749_/B _1594_/B _1595_/C vdd gnd AND2X2
X_1028_ _973_/A _1029_/C vdd gnd INVX1
X_1646_ _1650_/C _1646_/B _1646_/C _1650_/B _1647_/A vdd gnd AOI22X1
X_1715_ _1777_/A _1777_/B _1796_/B _1761_/A vdd gnd NAND3X1
X_1577_ _1787_/C _1904_/B _1577_/C _1915_/D vdd gnd OAI21X1
X_1500_ _1525_/A _1500_/B _1500_/C _1902_/B vdd gnd NAND3X1
X_1431_ _1431_/A _1751_/C vdd gnd INVX1
X_1362_ _1400_/B _1371_/A vdd gnd INVX1
X_1293_ _1293_/A _1293_/B _1293_/C _1297_/B vdd gnd OAI21X1
X_1629_ _1922_/Q _1629_/B _1631_/B vdd gnd NAND2X1
X_1276_ _976_/C _1276_/B _1276_/C _1278_/A vdd gnd NAND3X1
X_1414_ _1487_/A _1603_/A _1415_/A vdd gnd NAND2X1
X_1345_ _1525_/B _1524_/A _1345_/C _1346_/A vdd gnd OAI21X1
X_1130_ _973_/A _949_/A _1131_/A vdd gnd NAND2X1
X_987_ _987_/A _998_/B _987_/C _987_/Y vdd gnd OAI21X1
X_1061_ _1063_/C _1061_/B _1080_/D vdd gnd NOR2X1
X_1894_ _1902_/A _1902_/B _1934_/Q _1896_/C vdd gnd OAI21X1
X_1328_ _1440_/B _1702_/B _1330_/A _1482_/B _1329_/C vdd gnd AOI22X1
X_1259_ _951_/B _1525_/A vdd gnd INVX2
X_1113_ _1932_/Q _1818_/A vdd gnd INVX1
X_1044_ _1044_/A _1063_/C _1077_/D vdd gnd NOR2X1
X_1877_ _1877_/A _1892_/A _1878_/A vdd gnd NAND2X1
X_1800_ _1845_/B _1800_/B _1800_/C _1928_/D vdd gnd OAI21X1
X_1731_ _1731_/A _1731_/B _1731_/C _1732_/C vdd gnd AOI21X1
X_1662_ _1662_/A _1664_/B vdd gnd INVX1
X_1593_ _1593_/A _1593_/B _1718_/B _1594_/B vdd gnd NAND3X1
X_1027_ _1027_/A _978_/B _1027_/C _1074_/D vdd gnd OAI21X1
X_1929_ _1939_/S vdd _1929_/D _1939_/CLK _1929_/Q vdd gnd DFFSR
X_1576_ _1904_/B _1576_/B _1576_/C _1577_/C vdd gnd NAND3X1
X_1714_ _1790_/A _1790_/B _1777_/B vdd gnd NAND2X1
X_1645_ _1649_/B _1649_/A _1645_/C _1646_/C vdd gnd OAI21X1
X_1430_ _1757_/B _1757_/A _1431_/A vdd gnd NAND2X1
X_1292_ _1845_/A _975_/B _975_/A _1824_/A _1293_/C vdd gnd AOI22X1
X_1361_ _1735_/A _1735_/B _999_/C _1400_/B vdd gnd OAI21X1
X_1559_ _1559_/A _1580_/B vdd gnd INVX1
X_1628_ _1630_/B _1651_/A _1629_/B vdd gnd NAND2X1
X_1413_ _1605_/A _1603_/A vdd gnd INVX1
X_1275_ _951_/B _1335_/A _1335_/B _1278_/C vdd gnd NAND3X1
X_1344_ _1344_/A _1527_/A vdd gnd INVX1
X_1060_ _1060_/A _1063_/B _1061_/B vdd gnd NAND2X1
X_986_ _999_/A _999_/B _989_/A _987_/C vdd gnd OAI21X1
X_1893_ _1893_/A _1899_/B _1893_/C _1933_/D vdd gnd OAI21X1
X_1189_ _1191_/C _1300_/B _1192_/A vdd gnd OR2X2
X_1258_ _1258_/A _1258_/B _1258_/C _1280_/B vdd gnd AOI21X1
X_1327_ _1666_/A _1666_/B _1330_/A vdd gnd NOR2X1
X_1112_ _1161_/B _1291_/B _1140_/C vdd gnd OR2X2
X_969_ reset _969_/Y vdd gnd INVX8
X_1043_ _1043_/A _1059_/B _1044_/A vdd gnd NAND2X1
X_1876_ _1876_/A _1876_/B _1892_/A vdd gnd NAND2X1
X_1730_ _1742_/C _1742_/B _1743_/A _1731_/C vdd gnd AOI21X1
X_1592_ _1614_/B _1720_/C _1702_/A _1593_/B vdd gnd AOI21X1
X_1661_ _1818_/A _1815_/A _1662_/A vdd gnd NOR2X1
X_1026_ _978_/A _1029_/A _1027_/A vdd gnd NAND2X1
X_1859_ _1871_/B _1871_/C _1859_/C _1861_/B vdd gnd OAI21X1
X_1928_ _1939_/S vdd _1928_/D _1939_/CLK _1928_/Q vdd gnd DFFSR
X_1713_ _1771_/C _1772_/A _1713_/C _1777_/A vdd gnd NAND3X1
X_1575_ _1583_/A _1575_/B _1575_/C _1576_/B vdd gnd OAI21X1
X_1644_ _1704_/C _1649_/A _1698_/A _1645_/C vdd gnd OAI21X1
X_1009_ _1013_/B _997_/A _1015_/A _1010_/B vdd gnd OAI21X1
X_1360_ _1736_/B _1735_/B vdd gnd INVX1
X_1291_ _972_/B _1291_/B _1291_/C _1291_/D _1293_/B vdd gnd AOI22X1
X_1489_ _989_/B _1489_/B _1501_/A _1490_/B vdd gnd NAND3X1
X_1627_ _1736_/B _1635_/A _1627_/C _1630_/B vdd gnd AOI21X1
X_1558_ _1913_/Q _1912_/Q _1559_/A vdd gnd NOR2X1
X_1343_ _1343_/A _1472_/B _1343_/C _1344_/A vdd gnd NAND3X1
X_1412_ _1691_/B _1691_/C _1605_/A vdd gnd NAND2X1
X_1274_ _1757_/C _1274_/B _1335_/B vdd gnd NAND2X1
X_985_ _985_/A _996_/B _997_/C _987_/A vdd gnd NAND3X1
X_1892_ _1892_/A _1892_/B _1893_/A vdd gnd OR2X2
X_1326_ _1326_/A _1326_/B _1914_/Q _1666_/A vdd gnd AOI21X1
X_1188_ _1908_/Q _1497_/B _1300_/B vdd gnd NOR2X1
X_1257_ _1257_/A _1257_/B _1257_/C _1258_/C vdd gnd OAI21X1
X_968_ _999_/A enable _968_/Y vdd gnd AND2X2
X_1042_ _978_/A _1042_/B _1042_/C _1059_/B vdd gnd NAND3X1
X_1111_ _1111_/A _1111_/B _1120_/B vdd gnd AND2X2
X_1875_ _1875_/A _1875_/B _1876_/B vdd gnd OR2X2
X_1944_ _966_/A vsync vdd gnd BUFX2
X_1309_ _1743_/A _1723_/A _1309_/C _1655_/A vdd gnd NAND3X1
X_1591_ _1919_/Q _1727_/B _1614_/B vdd gnd NAND2X1
X_1660_ _1842_/B _1660_/B _1833_/A vdd gnd NAND2X1
X_1025_ _949_/A _1029_/A vdd gnd INVX1
X_1858_ _1870_/A _1871_/C vdd gnd INVX1
X_1927_ vdd _1940_/R _1927_/D _1937_/CLK _1927_/Q vdd gnd DFFSR
X_1789_ _1789_/A _1795_/B vdd gnd INVX1
X_1712_ _1712_/A _1712_/B _1772_/A vdd gnd NOR2X1
X_1643_ _1923_/Q _1643_/B _1924_/Q _1646_/B vdd gnd OAI21X1
X_1574_ _1575_/C _1574_/B _1576_/C vdd gnd OR2X2
X_1008_ _957_/A _1015_/A vdd gnd INVX1
X_1290_ _1290_/A _1290_/B _1290_/C _1291_/C vdd gnd OAI21X1
X_1626_ _1700_/C _1648_/B _1626_/C _1921_/D vdd gnd OAI21X1
X_1488_ _972_/A _973_/B _1501_/A vdd gnd NOR2X1
X_1557_ _1557_/A _1557_/B _1578_/A vdd gnd NOR2X1
X_1273_ _1697_/B _1274_/B vdd gnd INVX1
X_1342_ _975_/A _972_/B _1343_/C vdd gnd NOR2X1
X_1411_ _1727_/A _1727_/B _989_/A _1415_/B vdd gnd OAI21X1
X_1609_ _1919_/Q _1727_/B _1610_/A vdd gnd NOR2X1
X_984_ _995_/A _996_/B vdd gnd INVX1
X_1891_ _1902_/A _1902_/B _1933_/Q _1893_/C vdd gnd OAI21X1
X_1256_ _1256_/A _1256_/B _1257_/C vdd gnd NOR2X1
X_1325_ _1787_/A _1677_/B _1666_/B vdd gnd NOR2X1
X_1187_ _989_/B _1497_/B vdd gnd INVX1
X_1110_ _975_/A _1120_/A vdd gnd INVX1
X_967_ _967_/A _967_/B _967_/Y vdd gnd NOR2X1
X_1041_ _973_/A _972_/A _1042_/C vdd gnd AND2X2
X_1874_ _1889_/C _1889_/B _1874_/C _1877_/A vdd gnd AOI21X1
X_1943_ _1943_/A rgb vdd gnd BUFX2
X_1239_ _1913_/Q _1734_/C vdd gnd INVX1
X_1308_ _1910_/Q _1687_/B _1911_/Q _1674_/A vdd gnd OAI21X1
X_1590_ _1640_/B _1590_/B up _1650_/B vdd gnd OAI21X1
X_1024_ _949_/A _999_/A _1027_/C vdd gnd NAND2X1
X_1788_ _1788_/A _1788_/B _1788_/C _1795_/A vdd gnd AOI21X1
X_1857_ _1871_/A _1859_/C vdd gnd INVX1
X_1926_ _1939_/S vdd _1926_/D _1939_/CLK _1926_/Q vdd gnd DFFSR
X_1642_ _1642_/A _1643_/B vdd gnd INVX1
X_1711_ _1722_/C _1711_/B _1711_/C _1712_/A vdd gnd OAI21X1
X_1573_ _1573_/A _1574_/B vdd gnd INVX1
X_1007_ _957_/A _999_/C _1007_/C _1010_/A vdd gnd NAND3X1
X_1909_ _1939_/S vdd _1909_/D _1939_/CLK _1909_/Q vdd gnd DFFSR
X_1625_ _1625_/A _1651_/A _1626_/C vdd gnd NAND2X1
X_1556_ _1734_/C _1904_/B _1556_/C _1913_/D vdd gnd OAI21X1
X_1487_ _1487_/A _1487_/B _1490_/A vdd gnd NAND2X1
X_1410_ _1691_/B _1727_/B vdd gnd INVX1
X_1272_ _1326_/B _1272_/B _1326_/A _1697_/B vdd gnd NAND3X1
X_1341_ _1345_/C _1473_/C _1524_/B _1347_/A vdd gnd OAI21X1
X_1608_ _1614_/B _1610_/B vdd gnd INVX1
X_1539_ _1735_/C _1907_/A _1540_/A vdd gnd NOR2X1
X_983_ _989_/A _989_/B _995_/A vdd gnd AND2X2
X_1890_ _1890_/A _1899_/B _1890_/C _1932_/D vdd gnd OAI21X1
X_1255_ _1255_/A _1255_/B _1256_/B vdd gnd NOR2X1
X_1186_ _989_/B _1708_/B _1186_/C _1260_/B vdd gnd OAI21X1
X_1324_ _1440_/B _1702_/B _1324_/C _1329_/A vdd gnd OAI21X1
X_966_ _966_/A _999_/A _967_/A vdd gnd OR2X2
X_1040_ _949_/A _973_/B _1042_/B vdd gnd AND2X2
X_1942_ _967_/Y p_tick vdd gnd BUFX2
X_1873_ _1880_/B _1883_/B _1886_/B _1874_/C vdd gnd NAND3X1
X_1307_ _1684_/B _1680_/B vdd gnd INVX1
X_1169_ _1910_/Q _1723_/A vdd gnd INVX2
X_1238_ _1913_/Q _1440_/B _1241_/A vdd gnd NAND2X1
X_1023_ _1023_/A _1063_/C _1073_/D vdd gnd NOR2X1
X_949_ _949_/A _976_/B _963_/A vdd gnd NAND2X1
X_1925_ _1925_/R vdd _1925_/D _1925_/CLK _1925_/Q vdd gnd DFFSR
X_1787_ _1787_/A _1787_/B _1787_/C _1787_/D _1788_/C vdd gnd OAI22X1
X_1856_ _1856_/A _1856_/B _1895_/B vdd gnd NAND2X1
X_1710_ _1710_/A _1745_/C _1711_/C vdd gnd AND2X2
X_1572_ _1583_/A _1575_/B _1573_/A vdd gnd NOR2X1
X_1641_ _1641_/A _1650_/B _1650_/C vdd gnd NOR2X1
X_1006_ _996_/C _991_/A _1007_/C vdd gnd NOR2X1
X_1839_ _1846_/A _1844_/A vdd gnd INVX1
X_1908_ _1939_/S vdd _1908_/D _1939_/CLK _1908_/Q vdd gnd DFFSR
X_1555_ _1555_/A _1555_/B _1904_/B _1556_/C vdd gnd OAI21X1
X_1624_ _1718_/B _1650_/B _1624_/C _1625_/A vdd gnd OAI21X1
X_1486_ _1501_/B _1486_/B _1500_/B _1492_/A vdd gnd NAND3X1
X_1340_ _973_/B _1340_/B _1473_/C vdd gnd NAND2X1
X_1271_ _1787_/C _1787_/A _1272_/B vdd gnd NOR2X1
X_1469_ _1525_/A _1925_/Q _1469_/C _1470_/C vdd gnd AOI21X1
X_1538_ _1912_/Q _1940_/Q _1540_/B vdd gnd NOR2X1
X_1607_ _1722_/C _1648_/B _1607_/C _1918_/D vdd gnd OAI21X1
X_982_ _990_/A _990_/B _985_/A vdd gnd NAND2X1
X_1323_ _1675_/A _1675_/B _999_/C _1324_/C vdd gnd OAI21X1
X_1254_ _1440_/B _1913_/Q _1254_/C _1257_/A vdd gnd AOI21X1
X_1185_ _1190_/A _1300_/A _1186_/C vdd gnd AND2X2
X_965_ _978_/A _999_/A vdd gnd INVX4
X_1872_ _1872_/A _1872_/B _1886_/B vdd gnd NAND2X1
X_1941_ _954_/Y hsync vdd gnd BUFX2
X_1306_ _1306_/A _1306_/B _1306_/C _1317_/A vdd gnd NAND3X1
X_1237_ _957_/A _1440_/B vdd gnd INVX2
X_1099_ _1936_/Q _1101_/A _1100_/B vdd gnd NOR2X1
X_1168_ _1168_/A _1210_/B _1289_/B vdd gnd NOR2X1
X_948_ _948_/A _976_/B _976_/C _999_/B vdd gnd AOI21X1
X_1022_ _951_/B _1023_/A vdd gnd INVX1
X_1855_ _1855_/A _1855_/B _1855_/C _1856_/B vdd gnd OAI21X1
X_1924_ _1924_/R vdd _1924_/D _1925_/CLK _1924_/Q vdd gnd DFFSR
X_1786_ _1787_/A _1787_/B _1786_/C _1786_/D _1788_/B vdd gnd AOI22X1
X_1571_ _1915_/Q _1907_/A _1575_/B vdd gnd NOR2X1
X_1640_ _1781_/B _1640_/B _1641_/A vdd gnd NOR2X1
X_1005_ _999_/A _999_/B _957_/A _1011_/C vdd gnd OAI21X1
X_1838_ _1838_/A _1838_/B _1901_/A vdd gnd NAND2X1
X_1907_ _1907_/A _1907_/B _1907_/C _1940_/D vdd gnd OAI21X1
X_1769_ _1769_/A _1769_/B _1770_/C vdd gnd NAND2X1
X_1485_ _951_/B _976_/C _1486_/B vdd gnd NOR2X1
X_1554_ _1557_/A _1554_/B _1555_/A vdd gnd NOR2X1
X_1623_ _1921_/Q _1632_/B _1627_/C _1624_/C vdd gnd OAI21X1
.ends

