magic
tech scmos
magscale 1 2
timestamp 1702310163
<< nwell >>
rect -13 154 93 272
<< ntransistor >>
rect 18 14 22 34
rect 38 14 42 34
rect 58 14 62 54
<< ptransistor >>
rect 18 166 22 246
rect 28 166 32 246
rect 48 166 52 246
<< ndiffusion >>
rect 48 50 58 54
rect 16 14 18 34
rect 22 14 24 34
rect 36 14 38 34
rect 42 14 44 34
rect 56 14 58 50
rect 62 14 64 54
<< pdiffusion >>
rect 16 166 18 246
rect 22 166 28 246
rect 32 166 34 246
rect 46 166 48 246
rect 52 166 54 246
<< ndcontact >>
rect 4 14 16 34
rect 24 14 36 34
rect 44 14 56 50
rect 64 14 76 54
<< pdcontact >>
rect 4 166 16 246
rect 34 166 46 246
rect 54 166 66 246
<< psubstratepcontact >>
rect -7 -6 87 6
<< nsubstratencontact >>
rect -7 254 87 266
<< polysilicon >>
rect 18 246 22 250
rect 28 246 32 250
rect 48 246 52 250
rect 18 117 22 166
rect 17 105 22 117
rect 18 34 22 105
rect 28 97 32 166
rect 48 156 52 166
rect 28 85 30 97
rect 28 47 33 85
rect 60 60 62 72
rect 58 54 62 60
rect 28 43 42 47
rect 38 34 42 43
rect 18 10 22 14
rect 38 10 42 14
rect 58 10 62 14
<< polycontact >>
rect 5 105 17 117
rect 48 144 60 156
rect 30 85 42 97
rect 48 60 60 72
<< metal1 >>
rect -7 266 87 268
rect -7 252 87 254
rect 34 246 46 252
rect 4 156 12 166
rect 4 148 48 156
rect 3 123 17 137
rect 5 117 17 123
rect 23 103 37 117
rect 26 97 37 103
rect 26 85 30 97
rect 48 72 57 144
rect 66 137 74 182
rect 63 123 77 137
rect 26 60 48 67
rect 26 34 32 60
rect 66 54 74 123
rect 4 8 12 14
rect 44 8 56 14
rect -7 6 87 8
rect -7 -8 87 -6
<< m1p >>
rect -7 252 87 268
rect 3 123 17 137
rect 63 123 77 137
rect 23 103 37 117
rect -7 -8 87 8
<< labels >>
rlabel nsubstratencontact 40 260 40 260 0 vdd
port 4 nsew power bidirectional abutment
rlabel psubstratepcontact 40 0 40 0 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal1 10 127 10 127 0 A
port 1 nsew signal input
rlabel metal1 30 106 30 106 0 B
port 2 nsew signal input
rlabel metal1 70 131 70 131 0 Y
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 80 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
