magic
tech scmos
magscale 1 3
timestamp 1554524574
<< checkpaint >>
rect -56 -56 82 164
<< genericcontact >>
rect 10 79 16 85
rect 10 51 16 57
rect 10 23 16 29
<< metal1 >>
rect 4 4 22 104
<< end >>
