magic
tech scmos
magscale 1 3
timestamp 1554524574
<< checkpaint >>
rect -60 -60 78 78
<< polysilicon >>
rect 1 12 17 17
rect 1 6 6 12
rect 12 6 17 12
rect 1 1 17 6
<< polycontact >>
rect 6 6 12 12
<< metal1 >>
rect 0 12 18 18
rect 0 6 6 12
rect 12 6 18 12
rect 0 0 18 6
<< end >>
