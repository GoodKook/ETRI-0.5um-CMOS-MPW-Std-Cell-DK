magic
tech scmos
magscale 1 3
timestamp 1725342160
<< nwell >>
rect 110 110 380 380
<< diffusion >>
rect 76 426 414 444
rect 46 76 64 414
rect 151 341 339 359
rect 131 151 149 339
rect 196 196 294 294
rect 341 151 359 339
rect 151 131 339 149
rect 426 76 444 414
rect 76 46 414 64
<< pdiffusion >>
rect 195 294 295 295
rect 195 196 196 294
rect 294 196 295 294
rect 195 195 295 196
<< psubstratepdiff >>
rect 45 444 445 445
rect 45 426 76 444
rect 414 426 445 444
rect 45 425 445 426
rect 45 414 65 425
rect 45 76 46 414
rect 64 76 65 414
rect 425 414 445 425
rect 45 65 65 76
rect 425 76 426 414
rect 444 76 445 414
rect 425 65 445 76
rect 45 64 445 65
rect 45 46 76 64
rect 414 46 445 64
rect 45 45 445 46
<< nsubstratendiff >>
rect 130 359 360 360
rect 130 341 151 359
rect 339 341 360 359
rect 130 340 360 341
rect 130 339 150 340
rect 130 151 131 339
rect 149 151 150 339
rect 340 339 360 340
rect 130 150 150 151
rect 340 151 341 339
rect 359 151 360 339
rect 340 150 360 151
rect 130 149 360 150
rect 130 131 151 149
rect 339 131 360 149
rect 130 130 360 131
<< metal1 >>
rect 45 425 445 445
rect 45 65 65 425
rect 130 340 360 360
rect 130 150 150 340
rect 195 195 295 295
rect 340 150 360 340
rect 130 130 360 150
rect 425 65 445 425
rect 45 45 445 65
<< end >>
