magic
tech scmos
magscale 1 3
timestamp 1723010381
<< checkpaint >>
rect -15 -15 425 425
use pnp2_CDNS_7230122529112  pnp2_CDNS_7230122529112_0
timestamp 1723012252
transform 1 0 0 0 1 0
box 45 45 365 365
<< end >>
