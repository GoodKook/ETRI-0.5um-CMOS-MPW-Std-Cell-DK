VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pong_pt1
  CLASS BLOCK ;
  FOREIGN pong_pt1 ;
  ORIGIN 0.000 6.000 ;
  SIZE 864.000 BY 843.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 828.300 873.300 830.700 ;
        RECT 864.300 758.700 873.300 828.300 ;
        RECT 0.600 756.300 873.300 758.700 ;
        RECT 864.300 686.700 873.300 756.300 ;
        RECT 0.600 684.300 873.300 686.700 ;
        RECT 864.300 614.700 873.300 684.300 ;
        RECT 0.600 612.300 873.300 614.700 ;
        RECT 864.300 542.700 873.300 612.300 ;
        RECT 0.600 540.300 873.300 542.700 ;
        RECT 864.300 470.700 873.300 540.300 ;
        RECT 0.600 468.300 873.300 470.700 ;
        RECT 864.300 398.700 873.300 468.300 ;
        RECT 0.600 396.300 873.300 398.700 ;
        RECT 864.300 326.700 873.300 396.300 ;
        RECT 0.600 324.300 873.300 326.700 ;
        RECT 864.300 254.700 873.300 324.300 ;
        RECT 0.600 252.300 873.300 254.700 ;
        RECT 864.300 182.700 873.300 252.300 ;
        RECT 0.600 180.300 873.300 182.700 ;
        RECT 864.300 110.700 873.300 180.300 ;
        RECT 0.600 108.300 873.300 110.700 ;
        RECT 864.300 38.700 873.300 108.300 ;
        RECT 0.600 36.300 873.300 38.700 ;
        RECT 864.300 0.300 873.300 36.300 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -9.300 794.700 -0.300 830.700 ;
        RECT -9.300 792.300 863.400 794.700 ;
        RECT -9.300 722.700 -0.300 792.300 ;
        RECT 61.950 790.950 64.050 792.300 ;
        RECT 271.950 722.700 274.050 724.050 ;
        RECT -9.300 720.300 863.400 722.700 ;
        RECT -9.300 650.700 -0.300 720.300 ;
        RECT 16.950 718.950 19.050 720.300 ;
        RECT 199.950 718.950 202.050 720.300 ;
        RECT 691.950 718.950 694.050 720.300 ;
        RECT 859.950 718.950 862.050 720.300 ;
        RECT 766.950 650.700 769.050 652.050 ;
        RECT -9.300 648.300 863.400 650.700 ;
        RECT -9.300 578.700 -0.300 648.300 ;
        RECT 76.950 646.950 79.050 648.300 ;
        RECT 859.950 646.950 862.050 648.300 ;
        RECT -9.300 576.300 863.400 578.700 ;
        RECT -9.300 506.700 -0.300 576.300 ;
        RECT 13.950 574.950 16.050 576.300 ;
        RECT 469.950 574.950 472.050 576.300 ;
        RECT 607.950 574.950 610.050 576.300 ;
        RECT 754.950 574.950 757.050 576.300 ;
        RECT 859.950 574.950 862.050 576.300 ;
        RECT 859.950 506.700 862.050 508.050 ;
        RECT -9.300 504.300 863.400 506.700 ;
        RECT -9.300 434.700 -0.300 504.300 ;
        RECT 460.950 502.950 463.050 504.300 ;
        RECT 721.950 502.950 724.050 504.300 ;
        RECT 745.950 502.950 748.050 504.300 ;
        RECT 856.950 438.450 859.050 439.050 ;
        RECT 856.950 437.550 861.450 438.450 ;
        RECT 856.950 436.950 859.050 437.550 ;
        RECT 220.950 434.700 223.050 436.050 ;
        RECT 860.550 434.700 861.450 437.550 ;
        RECT -9.300 432.300 863.400 434.700 ;
        RECT -9.300 362.700 -0.300 432.300 ;
        RECT 148.950 430.950 151.050 432.300 ;
        RECT 613.950 430.950 616.050 432.300 ;
        RECT 688.950 362.700 691.050 364.050 ;
        RECT -9.300 360.300 863.400 362.700 ;
        RECT -9.300 290.700 -0.300 360.300 ;
        RECT 466.950 358.950 469.050 360.300 ;
        RECT -9.300 288.300 863.400 290.700 ;
        RECT -9.300 218.700 -0.300 288.300 ;
        RECT 763.950 286.950 766.050 288.300 ;
        RECT -9.300 216.300 863.400 218.700 ;
        RECT -9.300 146.700 -0.300 216.300 ;
        RECT 13.950 213.450 16.050 214.050 ;
        RECT 20.550 213.450 21.450 216.300 ;
        RECT 334.950 214.950 337.050 216.300 ;
        RECT 835.950 214.950 838.050 216.300 ;
        RECT 13.950 212.550 21.450 213.450 ;
        RECT 13.950 211.950 16.050 212.550 ;
        RECT -9.300 144.300 863.400 146.700 ;
        RECT -9.300 74.700 -0.300 144.300 ;
        RECT 76.950 142.950 79.050 144.300 ;
        RECT -9.300 72.300 863.400 74.700 ;
        RECT -9.300 2.700 -0.300 72.300 ;
        RECT 73.950 70.950 76.050 72.300 ;
        RECT 190.950 70.950 193.050 72.300 ;
        RECT 502.950 70.950 505.050 72.300 ;
        RECT 691.950 70.950 694.050 72.300 ;
        RECT 859.950 70.950 862.050 72.300 ;
        RECT 100.950 2.700 103.050 4.050 ;
        RECT 859.950 2.700 862.050 4.050 ;
        RECT -9.300 0.300 863.400 2.700 ;
      LAYER metal2 ;
        RECT 58.950 813.450 61.050 814.050 ;
        RECT 277.950 813.450 280.050 814.050 ;
        RECT 58.950 812.400 63.450 813.450 ;
        RECT 58.950 811.950 61.050 812.400 ;
        RECT 62.400 793.050 63.450 812.400 ;
        RECT 277.950 812.400 282.450 813.450 ;
        RECT 277.950 811.950 280.050 812.400 ;
        RECT 61.950 792.450 64.050 793.050 ;
        RECT 61.950 791.400 66.450 792.450 ;
        RECT 61.950 790.950 64.050 791.400 ;
        RECT 65.400 775.050 66.450 791.400 ;
        RECT 281.400 775.050 282.450 812.400 ;
        RECT 64.950 772.950 67.050 775.050 ;
        RECT 73.950 772.950 76.050 775.050 ;
        RECT 220.950 772.950 223.050 775.050 ;
        RECT 280.950 772.950 283.050 775.050 ;
        RECT 343.950 772.950 346.050 775.050 ;
        RECT 281.400 760.050 282.450 772.950 ;
        RECT 271.950 757.950 274.050 760.050 ;
        RECT 280.950 757.950 283.050 760.050 ;
        RECT 10.950 741.450 13.050 742.050 ;
        RECT 10.950 740.400 15.450 741.450 ;
        RECT 10.950 739.950 13.050 740.400 ;
        RECT 14.400 720.450 15.450 740.400 ;
        RECT 272.400 739.050 273.450 757.950 ;
        RECT 832.950 739.950 835.050 742.050 ;
        RECT 859.950 739.950 862.050 742.050 ;
        RECT 229.950 736.950 232.050 739.050 ;
        RECT 271.950 736.950 274.050 739.050 ;
        RECT 272.400 724.050 273.450 736.950 ;
        RECT 271.950 721.950 274.050 724.050 ;
        RECT 860.400 721.050 861.450 739.950 ;
        RECT 16.950 720.450 19.050 721.050 ;
        RECT 14.400 719.400 19.050 720.450 ;
        RECT 16.950 718.950 19.050 719.400 ;
        RECT 199.950 718.950 202.050 721.050 ;
        RECT 691.950 720.450 694.050 721.050 ;
        RECT 694.950 720.450 697.050 721.050 ;
        RECT 691.950 719.400 697.050 720.450 ;
        RECT 691.950 718.950 694.050 719.400 ;
        RECT 694.950 718.950 697.050 719.400 ;
        RECT 706.950 718.950 709.050 721.050 ;
        RECT 859.950 718.950 862.050 721.050 ;
        RECT 17.400 700.050 18.450 718.950 ;
        RECT 200.400 703.050 201.450 718.950 ;
        RECT 40.950 700.950 43.050 703.050 ;
        RECT 199.950 700.950 202.050 703.050 ;
        RECT 223.950 700.950 226.050 703.050 ;
        RECT 41.400 700.050 42.450 700.950 ;
        RECT 10.950 697.950 13.050 700.050 ;
        RECT 16.950 697.950 19.050 700.050 ;
        RECT 40.950 697.950 43.050 700.050 ;
        RECT 11.400 670.050 12.450 697.950 ;
        RECT 707.400 670.050 708.450 718.950 ;
        RECT 829.950 700.950 832.050 703.050 ;
        RECT 830.400 700.050 831.450 700.950 ;
        RECT 860.400 700.050 861.450 718.950 ;
        RECT 829.950 697.950 832.050 700.050 ;
        RECT 859.950 697.950 862.050 700.050 ;
        RECT 10.950 667.950 13.050 670.050 ;
        RECT 706.950 667.950 709.050 670.050 ;
        RECT 766.950 649.950 769.050 652.050 ;
        RECT 76.950 646.950 79.050 649.050 ;
        RECT 77.400 631.050 78.450 646.950 ;
        RECT 767.400 631.050 768.450 649.950 ;
        RECT 826.950 646.950 829.050 649.050 ;
        RECT 859.950 646.950 862.050 649.050 ;
        RECT 10.950 628.950 13.050 631.050 ;
        RECT 76.950 628.950 79.050 631.050 ;
        RECT 757.950 628.950 760.050 631.050 ;
        RECT 766.950 628.950 769.050 631.050 ;
        RECT 827.400 630.450 828.450 646.950 ;
        RECT 860.400 646.050 861.450 646.950 ;
        RECT 859.950 643.950 862.050 646.050 ;
        RECT 829.950 630.450 832.050 631.050 ;
        RECT 827.400 629.400 832.050 630.450 ;
        RECT 829.950 628.950 832.050 629.400 ;
        RECT 10.950 597.450 13.050 598.050 ;
        RECT 751.950 597.450 754.050 598.050 ;
        RECT 10.950 596.400 15.450 597.450 ;
        RECT 10.950 595.950 13.050 596.400 ;
        RECT 14.400 577.050 15.450 596.400 ;
        RECT 751.950 596.400 756.450 597.450 ;
        RECT 751.950 595.950 754.050 596.400 ;
        RECT 755.400 577.050 756.450 596.400 ;
        RECT 13.950 574.950 16.050 577.050 ;
        RECT 469.950 574.950 472.050 577.050 ;
        RECT 607.950 574.950 610.050 577.050 ;
        RECT 754.950 574.950 757.050 577.050 ;
        RECT 859.950 574.950 862.050 577.050 ;
        RECT 470.400 559.050 471.450 574.950 ;
        RECT 448.950 556.950 451.050 559.050 ;
        RECT 469.950 556.950 472.050 559.050 ;
        RECT 608.400 531.450 609.450 574.950 ;
        RECT 860.400 559.050 861.450 574.950 ;
        RECT 835.950 556.950 838.050 559.050 ;
        RECT 859.950 556.950 862.050 559.050 ;
        RECT 608.400 530.400 612.450 531.450 ;
        RECT 472.950 523.950 475.050 526.050 ;
        RECT 490.950 523.950 493.050 526.050 ;
        RECT 473.400 505.050 474.450 523.950 ;
        RECT 611.400 523.050 612.450 530.400 ;
        RECT 742.950 525.450 745.050 526.050 ;
        RECT 742.950 524.400 747.450 525.450 ;
        RECT 742.950 523.950 745.050 524.400 ;
        RECT 610.950 520.950 613.050 523.050 ;
        RECT 619.950 520.950 622.050 523.050 ;
        RECT 460.950 504.450 463.050 505.050 ;
        RECT 463.950 504.450 466.050 505.050 ;
        RECT 460.950 503.400 466.050 504.450 ;
        RECT 460.950 502.950 463.050 503.400 ;
        RECT 463.950 502.950 466.050 503.400 ;
        RECT 472.950 502.950 475.050 505.050 ;
        RECT 481.950 502.950 484.050 505.050 ;
        RECT 130.950 484.950 133.050 487.050 ;
        RECT 145.950 484.950 148.050 487.050 ;
        RECT 482.400 486.450 483.450 502.950 ;
        RECT 484.950 486.450 487.050 487.050 ;
        RECT 482.400 485.400 487.050 486.450 ;
        RECT 620.400 486.450 621.450 520.950 ;
        RECT 746.400 505.050 747.450 524.400 ;
        RECT 847.950 523.950 850.050 526.050 ;
        RECT 859.950 523.950 862.050 526.050 ;
        RECT 860.400 508.050 861.450 523.950 ;
        RECT 859.950 505.950 862.050 508.050 ;
        RECT 721.950 502.950 724.050 505.050 ;
        RECT 745.950 502.950 748.050 505.050 ;
        RECT 722.400 487.050 723.450 502.950 ;
        RECT 622.950 486.450 625.050 487.050 ;
        RECT 620.400 485.400 625.050 486.450 ;
        RECT 484.950 484.950 487.050 485.400 ;
        RECT 622.950 484.950 625.050 485.400 ;
        RECT 709.950 484.950 712.050 487.050 ;
        RECT 721.950 484.950 724.050 487.050 ;
        RECT 838.950 484.950 841.050 487.050 ;
        RECT 146.400 456.450 147.450 484.950 ;
        RECT 146.400 455.400 150.450 456.450 ;
        RECT 149.400 453.450 150.450 455.400 ;
        RECT 151.950 453.450 154.050 454.050 ;
        RECT 149.400 452.400 154.050 453.450 ;
        RECT 149.400 433.050 150.450 452.400 ;
        RECT 151.950 451.950 154.050 452.400 ;
        RECT 835.950 453.450 838.050 454.050 ;
        RECT 839.400 453.450 840.450 484.950 ;
        RECT 835.950 452.400 840.450 453.450 ;
        RECT 835.950 451.950 838.050 452.400 ;
        RECT 622.950 448.950 625.050 451.050 ;
        RECT 220.950 433.950 223.050 436.050 ;
        RECT 148.950 430.950 151.050 433.050 ;
        RECT 221.400 415.050 222.450 433.950 ;
        RECT 623.400 433.050 624.450 448.950 ;
        RECT 839.400 439.050 840.450 452.400 ;
        RECT 856.950 439.950 859.050 442.050 ;
        RECT 857.400 439.050 858.450 439.950 ;
        RECT 838.950 436.950 841.050 439.050 ;
        RECT 844.950 436.950 847.050 439.050 ;
        RECT 856.950 436.950 859.050 439.050 ;
        RECT 604.950 430.950 607.050 433.050 ;
        RECT 610.950 432.450 613.050 433.050 ;
        RECT 613.950 432.450 616.050 433.050 ;
        RECT 610.950 431.400 616.050 432.450 ;
        RECT 610.950 430.950 613.050 431.400 ;
        RECT 613.950 430.950 616.050 431.400 ;
        RECT 622.950 430.950 625.050 433.050 ;
        RECT 220.950 412.950 223.050 415.050 ;
        RECT 238.950 412.950 241.050 415.050 ;
        RECT 605.400 382.050 606.450 430.950 ;
        RECT 845.400 418.050 846.450 436.950 ;
        RECT 844.950 415.950 847.050 418.050 ;
        RECT 691.950 412.950 694.050 415.050 ;
        RECT 692.400 387.450 693.450 412.950 ;
        RECT 689.400 386.400 693.450 387.450 ;
        RECT 689.400 382.050 690.450 386.400 ;
        RECT 604.950 379.950 607.050 382.050 ;
        RECT 688.950 379.950 691.050 382.050 ;
        RECT 712.950 379.950 715.050 382.050 ;
        RECT 466.950 376.950 469.050 379.050 ;
        RECT 467.400 361.050 468.450 376.950 ;
        RECT 689.400 364.050 690.450 379.950 ;
        RECT 688.950 361.950 691.050 364.050 ;
        RECT 466.950 358.950 469.050 361.050 ;
        RECT 689.400 343.050 690.450 361.950 ;
        RECT 664.950 340.950 667.050 343.050 ;
        RECT 685.950 340.950 688.050 343.050 ;
        RECT 688.950 340.950 691.050 343.050 ;
        RECT 763.950 286.950 766.050 289.050 ;
        RECT 764.400 277.050 765.450 286.950 ;
        RECT 763.950 274.950 766.050 277.050 ;
        RECT 10.950 268.950 13.050 271.050 ;
        RECT 790.950 268.950 793.050 271.050 ;
        RECT 11.400 243.450 12.450 268.950 ;
        RECT 11.400 242.400 15.450 243.450 ;
        RECT 14.400 214.050 15.450 242.400 ;
        RECT 319.950 235.950 322.050 238.050 ;
        RECT 334.950 235.950 337.050 238.050 ;
        RECT 335.400 217.050 336.450 235.950 ;
        RECT 334.950 214.950 337.050 217.050 ;
        RECT 835.950 214.950 838.050 217.050 ;
        RECT 13.950 211.950 16.050 214.050 ;
        RECT 836.400 166.050 837.450 214.950 ;
        RECT 835.950 163.950 838.050 166.050 ;
        RECT 76.950 142.950 79.050 145.050 ;
        RECT 77.400 127.050 78.450 142.950 ;
        RECT 10.950 124.950 13.050 127.050 ;
        RECT 76.950 124.950 79.050 127.050 ;
        RECT 73.950 70.950 76.050 73.050 ;
        RECT 190.950 70.950 193.050 73.050 ;
        RECT 502.950 72.450 505.050 73.050 ;
        RECT 505.950 72.450 508.050 73.050 ;
        RECT 502.950 71.400 508.050 72.450 ;
        RECT 502.950 70.950 505.050 71.400 ;
        RECT 505.950 70.950 508.050 71.400 ;
        RECT 544.950 70.950 547.050 73.050 ;
        RECT 691.950 70.950 694.050 73.050 ;
        RECT 859.950 70.950 862.050 73.050 ;
        RECT 74.400 55.050 75.450 70.950 ;
        RECT 10.950 52.950 13.050 55.050 ;
        RECT 73.950 52.950 76.050 55.050 ;
        RECT 191.400 22.050 192.450 70.950 ;
        RECT 545.400 46.050 546.450 70.950 ;
        RECT 604.950 52.950 607.050 55.050 ;
        RECT 676.950 52.950 679.050 55.050 ;
        RECT 605.400 46.050 606.450 52.950 ;
        RECT 544.950 43.950 547.050 46.050 ;
        RECT 604.950 43.950 607.050 46.050 ;
        RECT 677.400 25.050 678.450 52.950 ;
        RECT 692.400 25.050 693.450 70.950 ;
        RECT 860.400 55.050 861.450 70.950 ;
        RECT 835.950 52.950 838.050 55.050 ;
        RECT 859.950 52.950 862.050 55.050 ;
        RECT 646.950 22.950 649.050 25.050 ;
        RECT 676.950 22.950 679.050 25.050 ;
        RECT 691.950 22.950 694.050 25.050 ;
        RECT 647.400 22.050 648.450 22.950 ;
        RECT 10.950 19.950 13.050 22.050 ;
        RECT 100.950 19.950 103.050 22.050 ;
        RECT 190.950 19.950 193.050 22.050 ;
        RECT 646.950 19.950 649.050 22.050 ;
        RECT 841.950 19.950 844.050 22.050 ;
        RECT 859.950 19.950 862.050 22.050 ;
        RECT 101.400 4.050 102.450 19.950 ;
        RECT 860.400 4.050 861.450 19.950 ;
        RECT 100.950 1.950 103.050 4.050 ;
        RECT 859.950 1.950 862.050 4.050 ;
      LAYER metal3 ;
        RECT 64.950 774.600 67.050 775.050 ;
        RECT 73.950 774.600 76.050 775.050 ;
        RECT 64.950 773.400 76.050 774.600 ;
        RECT 64.950 772.950 67.050 773.400 ;
        RECT 73.950 772.950 76.050 773.400 ;
        RECT 220.950 774.600 223.050 775.050 ;
        RECT 280.950 774.600 283.050 775.050 ;
        RECT 343.950 774.600 346.050 775.050 ;
        RECT 220.950 773.400 346.050 774.600 ;
        RECT 220.950 772.950 223.050 773.400 ;
        RECT 280.950 772.950 283.050 773.400 ;
        RECT 343.950 772.950 346.050 773.400 ;
        RECT 271.950 759.600 274.050 760.050 ;
        RECT 280.950 759.600 283.050 760.050 ;
        RECT 271.950 758.400 283.050 759.600 ;
        RECT 271.950 757.950 274.050 758.400 ;
        RECT 280.950 757.950 283.050 758.400 ;
        RECT 832.950 741.600 835.050 742.050 ;
        RECT 859.950 741.600 862.050 742.050 ;
        RECT 832.950 740.400 862.050 741.600 ;
        RECT 832.950 739.950 835.050 740.400 ;
        RECT 859.950 739.950 862.050 740.400 ;
        RECT 229.950 738.600 232.050 739.050 ;
        RECT 271.950 738.600 274.050 739.050 ;
        RECT 229.950 737.400 274.050 738.600 ;
        RECT 229.950 736.950 232.050 737.400 ;
        RECT 271.950 736.950 274.050 737.400 ;
        RECT 694.950 720.600 697.050 721.050 ;
        RECT 706.950 720.600 709.050 721.050 ;
        RECT 694.950 719.400 709.050 720.600 ;
        RECT 694.950 718.950 697.050 719.400 ;
        RECT 706.950 718.950 709.050 719.400 ;
        RECT 199.950 702.600 202.050 703.050 ;
        RECT 223.950 702.600 226.050 703.050 ;
        RECT 199.950 701.400 226.050 702.600 ;
        RECT 199.950 700.950 202.050 701.400 ;
        RECT 223.950 700.950 226.050 701.400 ;
        RECT 10.950 699.600 13.050 700.050 ;
        RECT 16.950 699.600 19.050 700.050 ;
        RECT 40.950 699.600 43.050 700.050 ;
        RECT 10.950 698.400 43.050 699.600 ;
        RECT 10.950 697.950 13.050 698.400 ;
        RECT 16.950 697.950 19.050 698.400 ;
        RECT 40.950 697.950 43.050 698.400 ;
        RECT 829.950 699.600 832.050 700.050 ;
        RECT 859.950 699.600 862.050 700.050 ;
        RECT 829.950 698.400 862.050 699.600 ;
        RECT 829.950 697.950 832.050 698.400 ;
        RECT 859.950 697.950 862.050 698.400 ;
        RECT 826.950 648.600 829.050 649.050 ;
        RECT 826.950 647.400 861.600 648.600 ;
        RECT 826.950 646.950 829.050 647.400 ;
        RECT 860.400 646.050 861.600 647.400 ;
        RECT 859.950 643.950 862.050 646.050 ;
        RECT 10.950 630.600 13.050 631.050 ;
        RECT 76.950 630.600 79.050 631.050 ;
        RECT 10.950 629.400 79.050 630.600 ;
        RECT 10.950 628.950 13.050 629.400 ;
        RECT 76.950 628.950 79.050 629.400 ;
        RECT 757.950 630.600 760.050 631.050 ;
        RECT 766.950 630.600 769.050 631.050 ;
        RECT 757.950 629.400 769.050 630.600 ;
        RECT 757.950 628.950 760.050 629.400 ;
        RECT 766.950 628.950 769.050 629.400 ;
        RECT 448.950 558.600 451.050 559.050 ;
        RECT 469.950 558.600 472.050 559.050 ;
        RECT 448.950 557.400 472.050 558.600 ;
        RECT 448.950 556.950 451.050 557.400 ;
        RECT 469.950 556.950 472.050 557.400 ;
        RECT 835.950 558.600 838.050 559.050 ;
        RECT 859.950 558.600 862.050 559.050 ;
        RECT 835.950 557.400 862.050 558.600 ;
        RECT 835.950 556.950 838.050 557.400 ;
        RECT 859.950 556.950 862.050 557.400 ;
        RECT 472.950 525.600 475.050 526.050 ;
        RECT 490.950 525.600 493.050 526.050 ;
        RECT 472.950 524.400 493.050 525.600 ;
        RECT 472.950 523.950 475.050 524.400 ;
        RECT 490.950 523.950 493.050 524.400 ;
        RECT 847.950 525.600 850.050 526.050 ;
        RECT 859.950 525.600 862.050 526.050 ;
        RECT 847.950 524.400 862.050 525.600 ;
        RECT 847.950 523.950 850.050 524.400 ;
        RECT 859.950 523.950 862.050 524.400 ;
        RECT 610.950 522.600 613.050 523.050 ;
        RECT 619.950 522.600 622.050 523.050 ;
        RECT 610.950 521.400 622.050 522.600 ;
        RECT 610.950 520.950 613.050 521.400 ;
        RECT 619.950 520.950 622.050 521.400 ;
        RECT 463.950 504.600 466.050 505.050 ;
        RECT 472.950 504.600 475.050 505.050 ;
        RECT 481.950 504.600 484.050 505.050 ;
        RECT 463.950 503.400 484.050 504.600 ;
        RECT 463.950 502.950 466.050 503.400 ;
        RECT 472.950 502.950 475.050 503.400 ;
        RECT 481.950 502.950 484.050 503.400 ;
        RECT 130.950 486.600 133.050 487.050 ;
        RECT 145.950 486.600 148.050 487.050 ;
        RECT 130.950 485.400 148.050 486.600 ;
        RECT 130.950 484.950 133.050 485.400 ;
        RECT 145.950 484.950 148.050 485.400 ;
        RECT 709.950 486.600 712.050 487.050 ;
        RECT 721.950 486.600 724.050 487.050 ;
        RECT 709.950 485.400 724.050 486.600 ;
        RECT 709.950 484.950 712.050 485.400 ;
        RECT 721.950 484.950 724.050 485.400 ;
        RECT 856.950 439.950 859.050 442.050 ;
        RECT 838.950 438.600 841.050 439.050 ;
        RECT 844.950 438.600 847.050 439.050 ;
        RECT 857.400 438.600 858.600 439.950 ;
        RECT 838.950 437.400 858.600 438.600 ;
        RECT 838.950 436.950 841.050 437.400 ;
        RECT 844.950 436.950 847.050 437.400 ;
        RECT 604.950 432.600 607.050 433.050 ;
        RECT 610.950 432.600 613.050 433.050 ;
        RECT 622.950 432.600 625.050 433.050 ;
        RECT 604.950 431.400 625.050 432.600 ;
        RECT 604.950 430.950 607.050 431.400 ;
        RECT 610.950 430.950 613.050 431.400 ;
        RECT 622.950 430.950 625.050 431.400 ;
        RECT 220.950 414.600 223.050 415.050 ;
        RECT 238.950 414.600 241.050 415.050 ;
        RECT 220.950 413.400 241.050 414.600 ;
        RECT 220.950 412.950 223.050 413.400 ;
        RECT 238.950 412.950 241.050 413.400 ;
        RECT 688.950 381.600 691.050 382.050 ;
        RECT 712.950 381.600 715.050 382.050 ;
        RECT 688.950 380.400 715.050 381.600 ;
        RECT 688.950 379.950 691.050 380.400 ;
        RECT 712.950 379.950 715.050 380.400 ;
        RECT 664.950 342.600 667.050 343.050 ;
        RECT 685.950 342.600 688.050 343.050 ;
        RECT 688.950 342.600 691.050 343.050 ;
        RECT 664.950 341.400 691.050 342.600 ;
        RECT 664.950 340.950 667.050 341.400 ;
        RECT 685.950 340.950 688.050 341.400 ;
        RECT 688.950 340.950 691.050 341.400 ;
        RECT 763.950 276.600 766.050 277.050 ;
        RECT 763.950 275.400 792.600 276.600 ;
        RECT 763.950 274.950 766.050 275.400 ;
        RECT 791.400 271.050 792.600 275.400 ;
        RECT 790.950 268.950 793.050 271.050 ;
        RECT 319.950 237.600 322.050 238.050 ;
        RECT 334.950 237.600 337.050 238.050 ;
        RECT 319.950 236.400 337.050 237.600 ;
        RECT 319.950 235.950 322.050 236.400 ;
        RECT 334.950 235.950 337.050 236.400 ;
        RECT 10.950 126.600 13.050 127.050 ;
        RECT 76.950 126.600 79.050 127.050 ;
        RECT 10.950 125.400 79.050 126.600 ;
        RECT 10.950 124.950 13.050 125.400 ;
        RECT 76.950 124.950 79.050 125.400 ;
        RECT 505.950 72.600 508.050 73.050 ;
        RECT 544.950 72.600 547.050 73.050 ;
        RECT 505.950 71.400 547.050 72.600 ;
        RECT 505.950 70.950 508.050 71.400 ;
        RECT 544.950 70.950 547.050 71.400 ;
        RECT 10.950 54.600 13.050 55.050 ;
        RECT 73.950 54.600 76.050 55.050 ;
        RECT 10.950 53.400 76.050 54.600 ;
        RECT 10.950 52.950 13.050 53.400 ;
        RECT 73.950 52.950 76.050 53.400 ;
        RECT 835.950 54.600 838.050 55.050 ;
        RECT 859.950 54.600 862.050 55.050 ;
        RECT 835.950 53.400 862.050 54.600 ;
        RECT 835.950 52.950 838.050 53.400 ;
        RECT 859.950 52.950 862.050 53.400 ;
        RECT 544.950 45.600 547.050 46.050 ;
        RECT 604.950 45.600 607.050 46.050 ;
        RECT 544.950 44.400 607.050 45.600 ;
        RECT 544.950 43.950 547.050 44.400 ;
        RECT 604.950 43.950 607.050 44.400 ;
        RECT 646.950 24.600 649.050 25.050 ;
        RECT 676.950 24.600 679.050 25.050 ;
        RECT 691.950 24.600 694.050 25.050 ;
        RECT 646.950 23.400 694.050 24.600 ;
        RECT 646.950 22.950 649.050 23.400 ;
        RECT 676.950 22.950 679.050 23.400 ;
        RECT 691.950 22.950 694.050 23.400 ;
        RECT 10.950 21.600 13.050 22.050 ;
        RECT 100.950 21.600 103.050 22.050 ;
        RECT 10.950 20.400 103.050 21.600 ;
        RECT 10.950 19.950 13.050 20.400 ;
        RECT 100.950 19.950 103.050 20.400 ;
        RECT 841.950 21.600 844.050 22.050 ;
        RECT 859.950 21.600 862.050 22.050 ;
        RECT 841.950 20.400 862.050 21.600 ;
        RECT 841.950 19.950 844.050 20.400 ;
        RECT 859.950 19.950 862.050 20.400 ;
    END
  END vdd
  PIN clk
    PORT
      LAYER metal2 ;
        RECT 410.400 813.450 411.450 837.450 ;
        RECT 412.950 813.450 415.050 814.050 ;
        RECT 410.400 812.400 415.050 813.450 ;
        RECT 412.950 811.950 415.050 812.400 ;
        RECT 413.400 793.050 414.450 811.950 ;
        RECT 262.950 790.950 265.050 793.050 ;
        RECT 412.950 790.950 415.050 793.050 ;
        RECT 718.950 790.950 721.050 793.050 ;
        RECT 263.400 747.450 264.450 790.950 ;
        RECT 263.400 746.400 267.450 747.450 ;
        RECT 266.400 640.050 267.450 746.400 ;
        RECT 719.400 646.050 720.450 790.950 ;
        RECT 736.950 667.950 739.050 670.050 ;
        RECT 737.400 646.050 738.450 667.950 ;
        RECT 703.950 643.950 706.050 646.050 ;
        RECT 718.950 643.950 721.050 646.050 ;
        RECT 736.950 643.950 739.050 646.050 ;
        RECT 211.950 637.950 214.050 640.050 ;
        RECT 265.950 637.950 268.050 640.050 ;
        RECT 212.400 607.050 213.450 637.950 ;
        RECT 704.400 615.450 705.450 643.950 ;
        RECT 701.400 614.400 705.450 615.450 ;
        RECT 169.950 604.950 172.050 607.050 ;
        RECT 211.950 604.950 214.050 607.050 ;
        RECT 170.400 562.050 171.450 604.950 ;
        RECT 157.950 559.950 160.050 562.050 ;
        RECT 169.950 559.950 172.050 562.050 ;
        RECT 158.400 559.050 159.450 559.950 ;
        RECT 701.400 559.050 702.450 614.400 ;
        RECT 157.950 556.950 160.050 559.050 ;
        RECT 700.950 556.950 703.050 559.050 ;
        RECT 718.950 556.950 721.050 559.050 ;
        RECT 701.400 502.050 702.450 556.950 ;
        RECT 625.950 499.950 628.050 502.050 ;
        RECT 700.950 499.950 703.050 502.050 ;
        RECT 626.400 418.050 627.450 499.950 ;
        RECT 607.950 415.950 610.050 418.050 ;
        RECT 613.950 415.950 616.050 418.050 ;
        RECT 625.950 415.950 628.050 418.050 ;
        RECT 608.400 415.050 609.450 415.950 ;
        RECT 607.950 412.950 610.050 415.050 ;
        RECT 614.400 328.050 615.450 415.950 ;
        RECT 592.950 325.950 595.050 328.050 ;
        RECT 613.950 325.950 616.050 328.050 ;
        RECT 593.400 274.050 594.450 325.950 ;
        RECT 592.950 271.950 595.050 274.050 ;
        RECT 580.950 268.950 583.050 271.050 ;
        RECT 581.400 249.450 582.450 268.950 ;
        RECT 578.400 248.400 582.450 249.450 ;
        RECT 578.400 244.050 579.450 248.400 ;
        RECT 577.950 241.950 580.050 244.050 ;
        RECT 565.950 229.950 568.050 232.050 ;
        RECT 566.400 208.050 567.450 229.950 ;
        RECT 553.950 205.950 556.050 208.050 ;
        RECT 565.950 205.950 568.050 208.050 ;
        RECT 554.400 160.050 555.450 205.950 ;
        RECT 544.950 157.950 547.050 160.050 ;
        RECT 553.950 157.950 556.050 160.050 ;
        RECT 545.400 130.050 546.450 157.950 ;
        RECT 544.950 127.950 547.050 130.050 ;
        RECT 517.950 121.950 520.050 124.050 ;
        RECT 518.400 64.050 519.450 121.950 ;
        RECT 517.950 61.950 520.050 64.050 ;
        RECT 736.950 61.950 739.050 64.050 ;
        RECT 518.400 55.050 519.450 61.950 ;
        RECT 737.400 55.050 738.450 61.950 ;
        RECT 517.950 52.950 520.050 55.050 ;
        RECT 736.950 52.950 739.050 55.050 ;
      LAYER metal3 ;
        RECT 262.950 792.600 265.050 793.050 ;
        RECT 412.950 792.600 415.050 793.050 ;
        RECT 718.950 792.600 721.050 793.050 ;
        RECT 262.950 791.400 721.050 792.600 ;
        RECT 262.950 790.950 265.050 791.400 ;
        RECT 412.950 790.950 415.050 791.400 ;
        RECT 718.950 790.950 721.050 791.400 ;
        RECT 703.950 645.600 706.050 646.050 ;
        RECT 718.950 645.600 721.050 646.050 ;
        RECT 736.950 645.600 739.050 646.050 ;
        RECT 703.950 644.400 739.050 645.600 ;
        RECT 703.950 643.950 706.050 644.400 ;
        RECT 718.950 643.950 721.050 644.400 ;
        RECT 736.950 643.950 739.050 644.400 ;
        RECT 211.950 639.600 214.050 640.050 ;
        RECT 265.950 639.600 268.050 640.050 ;
        RECT 211.950 638.400 268.050 639.600 ;
        RECT 211.950 637.950 214.050 638.400 ;
        RECT 265.950 637.950 268.050 638.400 ;
        RECT 169.950 606.600 172.050 607.050 ;
        RECT 211.950 606.600 214.050 607.050 ;
        RECT 169.950 605.400 214.050 606.600 ;
        RECT 169.950 604.950 172.050 605.400 ;
        RECT 211.950 604.950 214.050 605.400 ;
        RECT 157.950 561.600 160.050 562.050 ;
        RECT 169.950 561.600 172.050 562.050 ;
        RECT 157.950 560.400 172.050 561.600 ;
        RECT 157.950 559.950 160.050 560.400 ;
        RECT 169.950 559.950 172.050 560.400 ;
        RECT 700.950 558.600 703.050 559.050 ;
        RECT 718.950 558.600 721.050 559.050 ;
        RECT 700.950 557.400 721.050 558.600 ;
        RECT 700.950 556.950 703.050 557.400 ;
        RECT 718.950 556.950 721.050 557.400 ;
        RECT 625.950 501.600 628.050 502.050 ;
        RECT 700.950 501.600 703.050 502.050 ;
        RECT 625.950 500.400 703.050 501.600 ;
        RECT 625.950 499.950 628.050 500.400 ;
        RECT 700.950 499.950 703.050 500.400 ;
        RECT 607.950 417.600 610.050 418.050 ;
        RECT 613.950 417.600 616.050 418.050 ;
        RECT 625.950 417.600 628.050 418.050 ;
        RECT 607.950 416.400 628.050 417.600 ;
        RECT 607.950 415.950 610.050 416.400 ;
        RECT 613.950 415.950 616.050 416.400 ;
        RECT 625.950 415.950 628.050 416.400 ;
        RECT 592.950 327.600 595.050 328.050 ;
        RECT 613.950 327.600 616.050 328.050 ;
        RECT 592.950 326.400 616.050 327.600 ;
        RECT 592.950 325.950 595.050 326.400 ;
        RECT 613.950 325.950 616.050 326.400 ;
        RECT 592.950 273.600 595.050 274.050 ;
        RECT 581.400 272.400 595.050 273.600 ;
        RECT 581.400 271.050 582.600 272.400 ;
        RECT 592.950 271.950 595.050 272.400 ;
        RECT 580.950 268.950 583.050 271.050 ;
        RECT 577.950 243.600 580.050 244.050 ;
        RECT 572.400 242.400 580.050 243.600 ;
        RECT 572.400 240.600 573.600 242.400 ;
        RECT 577.950 241.950 580.050 242.400 ;
        RECT 566.400 239.400 573.600 240.600 ;
        RECT 566.400 232.050 567.600 239.400 ;
        RECT 565.950 229.950 568.050 232.050 ;
        RECT 553.950 207.600 556.050 208.050 ;
        RECT 565.950 207.600 568.050 208.050 ;
        RECT 553.950 206.400 568.050 207.600 ;
        RECT 553.950 205.950 556.050 206.400 ;
        RECT 565.950 205.950 568.050 206.400 ;
        RECT 544.950 159.600 547.050 160.050 ;
        RECT 553.950 159.600 556.050 160.050 ;
        RECT 544.950 158.400 556.050 159.600 ;
        RECT 544.950 157.950 547.050 158.400 ;
        RECT 553.950 157.950 556.050 158.400 ;
        RECT 544.950 129.600 547.050 130.050 ;
        RECT 542.400 128.400 547.050 129.600 ;
        RECT 542.400 126.600 543.600 128.400 ;
        RECT 544.950 127.950 547.050 128.400 ;
        RECT 539.400 125.400 543.600 126.600 ;
        RECT 517.950 123.600 520.050 124.050 ;
        RECT 539.400 123.600 540.600 125.400 ;
        RECT 517.950 122.400 540.600 123.600 ;
        RECT 517.950 121.950 520.050 122.400 ;
        RECT 517.950 63.600 520.050 64.050 ;
        RECT 736.950 63.600 739.050 64.050 ;
        RECT 517.950 62.400 739.050 63.600 ;
        RECT 517.950 61.950 520.050 62.400 ;
        RECT 736.950 61.950 739.050 62.400 ;
    END
  END clk
  PIN down
    PORT
      LAYER metal1 ;
        RECT 478.950 201.450 481.050 202.050 ;
        RECT 470.550 200.550 481.050 201.450 ;
        RECT 466.950 192.450 469.050 193.050 ;
        RECT 470.550 192.450 471.450 200.550 ;
        RECT 478.950 199.950 481.050 200.550 ;
        RECT 466.950 191.550 471.450 192.450 ;
        RECT 466.950 190.950 469.050 191.550 ;
      LAYER metal2 ;
        RECT 464.400 807.450 465.450 837.450 ;
        RECT 461.400 806.400 465.450 807.450 ;
        RECT 461.400 802.050 462.450 806.400 ;
        RECT 460.950 799.950 463.050 802.050 ;
        RECT 490.950 799.950 493.050 802.050 ;
        RECT 491.400 676.050 492.450 799.950 ;
        RECT 490.950 673.950 493.050 676.050 ;
        RECT 487.950 664.950 490.050 667.050 ;
        RECT 488.400 601.050 489.450 664.950 ;
        RECT 463.950 598.950 466.050 601.050 ;
        RECT 487.950 598.950 490.050 601.050 ;
        RECT 464.400 592.050 465.450 598.950 ;
        RECT 457.950 589.950 460.050 592.050 ;
        RECT 463.950 589.950 466.050 592.050 ;
        RECT 458.400 544.050 459.450 589.950 ;
        RECT 439.950 541.950 442.050 544.050 ;
        RECT 457.950 541.950 460.050 544.050 ;
        RECT 440.400 510.450 441.450 541.950 ;
        RECT 440.400 509.400 444.450 510.450 ;
        RECT 443.400 481.050 444.450 509.400 ;
        RECT 442.950 478.950 445.050 481.050 ;
        RECT 469.950 478.950 472.050 481.050 ;
        RECT 470.400 445.050 471.450 478.950 ;
        RECT 442.950 442.950 445.050 445.050 ;
        RECT 469.950 442.950 472.050 445.050 ;
        RECT 443.400 393.450 444.450 442.950 ;
        RECT 443.400 392.400 447.450 393.450 ;
        RECT 446.400 367.050 447.450 392.400 ;
        RECT 439.950 364.950 442.050 367.050 ;
        RECT 445.950 364.950 448.050 367.050 ;
        RECT 440.400 319.050 441.450 364.950 ;
        RECT 439.950 316.950 442.050 319.050 ;
        RECT 445.950 316.950 448.050 319.050 ;
        RECT 446.400 306.450 447.450 316.950 ;
        RECT 443.400 305.400 447.450 306.450 ;
        RECT 443.400 294.450 444.450 305.400 ;
        RECT 440.400 293.400 444.450 294.450 ;
        RECT 440.400 277.050 441.450 293.400 ;
        RECT 439.950 274.950 442.050 277.050 ;
        RECT 433.950 271.950 436.050 274.050 ;
        RECT 434.400 247.050 435.450 271.950 ;
        RECT 433.950 244.950 436.050 247.050 ;
        RECT 478.950 235.950 481.050 238.050 ;
        RECT 479.400 202.050 480.450 235.950 ;
        RECT 478.950 199.950 481.050 202.050 ;
        RECT 466.950 190.950 469.050 193.050 ;
        RECT 467.400 166.050 468.450 190.950 ;
        RECT 466.950 163.950 469.050 166.050 ;
      LAYER metal3 ;
        RECT 460.950 801.600 463.050 802.050 ;
        RECT 490.950 801.600 493.050 802.050 ;
        RECT 460.950 800.400 493.050 801.600 ;
        RECT 460.950 799.950 463.050 800.400 ;
        RECT 490.950 799.950 493.050 800.400 ;
        RECT 490.950 673.950 493.050 676.050 ;
        RECT 491.400 672.600 492.600 673.950 ;
        RECT 488.400 671.400 492.600 672.600 ;
        RECT 488.400 667.050 489.600 671.400 ;
        RECT 487.950 664.950 490.050 667.050 ;
        RECT 463.950 600.600 466.050 601.050 ;
        RECT 487.950 600.600 490.050 601.050 ;
        RECT 463.950 599.400 490.050 600.600 ;
        RECT 463.950 598.950 466.050 599.400 ;
        RECT 487.950 598.950 490.050 599.400 ;
        RECT 457.950 591.600 460.050 592.050 ;
        RECT 463.950 591.600 466.050 592.050 ;
        RECT 457.950 590.400 466.050 591.600 ;
        RECT 457.950 589.950 460.050 590.400 ;
        RECT 463.950 589.950 466.050 590.400 ;
        RECT 439.950 543.600 442.050 544.050 ;
        RECT 457.950 543.600 460.050 544.050 ;
        RECT 439.950 542.400 460.050 543.600 ;
        RECT 439.950 541.950 442.050 542.400 ;
        RECT 457.950 541.950 460.050 542.400 ;
        RECT 442.950 480.600 445.050 481.050 ;
        RECT 469.950 480.600 472.050 481.050 ;
        RECT 442.950 479.400 472.050 480.600 ;
        RECT 442.950 478.950 445.050 479.400 ;
        RECT 469.950 478.950 472.050 479.400 ;
        RECT 442.950 444.600 445.050 445.050 ;
        RECT 469.950 444.600 472.050 445.050 ;
        RECT 442.950 443.400 472.050 444.600 ;
        RECT 442.950 442.950 445.050 443.400 ;
        RECT 469.950 442.950 472.050 443.400 ;
        RECT 439.950 366.600 442.050 367.050 ;
        RECT 445.950 366.600 448.050 367.050 ;
        RECT 439.950 365.400 448.050 366.600 ;
        RECT 439.950 364.950 442.050 365.400 ;
        RECT 445.950 364.950 448.050 365.400 ;
        RECT 439.950 318.600 442.050 319.050 ;
        RECT 445.950 318.600 448.050 319.050 ;
        RECT 439.950 317.400 448.050 318.600 ;
        RECT 439.950 316.950 442.050 317.400 ;
        RECT 445.950 316.950 448.050 317.400 ;
        RECT 439.950 274.950 442.050 277.050 ;
        RECT 433.950 273.600 436.050 274.050 ;
        RECT 440.400 273.600 441.600 274.950 ;
        RECT 433.950 272.400 441.600 273.600 ;
        RECT 433.950 271.950 436.050 272.400 ;
        RECT 433.950 246.600 436.050 247.050 ;
        RECT 433.950 245.400 474.600 246.600 ;
        RECT 433.950 244.950 436.050 245.400 ;
        RECT 473.400 237.600 474.600 245.400 ;
        RECT 478.950 237.600 481.050 238.050 ;
        RECT 473.400 236.400 481.050 237.600 ;
        RECT 478.950 235.950 481.050 236.400 ;
    END
  END down
  PIN enable
    PORT
      LAYER metal2 ;
        RECT 416.400 829.050 417.450 837.450 ;
        RECT 361.950 826.950 364.050 829.050 ;
        RECT 415.950 826.950 418.050 829.050 ;
        RECT 362.400 778.050 363.450 826.950 ;
        RECT 361.950 775.950 364.050 778.050 ;
      LAYER metal3 ;
        RECT 361.950 828.600 364.050 829.050 ;
        RECT 415.950 828.600 418.050 829.050 ;
        RECT 361.950 827.400 418.050 828.600 ;
        RECT 361.950 826.950 364.050 827.400 ;
        RECT 415.950 826.950 418.050 827.400 ;
    END
  END enable
  PIN hsync
    PORT
      LAYER metal2 ;
        RECT 547.950 337.950 550.050 340.050 ;
        RECT 548.400 315.450 549.450 337.950 ;
        RECT 545.400 314.400 549.450 315.450 ;
        RECT 545.400 202.050 546.450 314.400 ;
        RECT 544.950 199.950 547.050 202.050 ;
        RECT 550.950 199.950 553.050 202.050 ;
        RECT 551.400 172.050 552.450 199.950 ;
        RECT 502.950 169.950 505.050 172.050 ;
        RECT 550.950 169.950 553.050 172.050 ;
        RECT 503.400 151.050 504.450 169.950 ;
        RECT 502.950 148.950 505.050 151.050 ;
        RECT 514.950 148.950 517.050 151.050 ;
        RECT 515.400 100.050 516.450 148.950 ;
        RECT 514.950 97.950 517.050 100.050 ;
        RECT 520.950 97.950 523.050 100.050 ;
        RECT 521.400 4.050 522.450 97.950 ;
        RECT 520.950 1.950 523.050 4.050 ;
        RECT 544.950 1.950 547.050 4.050 ;
        RECT 545.400 -3.600 546.450 1.950 ;
      LAYER metal3 ;
        RECT 544.950 201.600 547.050 202.050 ;
        RECT 550.950 201.600 553.050 202.050 ;
        RECT 544.950 200.400 553.050 201.600 ;
        RECT 544.950 199.950 547.050 200.400 ;
        RECT 550.950 199.950 553.050 200.400 ;
        RECT 502.950 171.600 505.050 172.050 ;
        RECT 550.950 171.600 553.050 172.050 ;
        RECT 502.950 170.400 553.050 171.600 ;
        RECT 502.950 169.950 505.050 170.400 ;
        RECT 550.950 169.950 553.050 170.400 ;
        RECT 502.950 150.600 505.050 151.050 ;
        RECT 514.950 150.600 517.050 151.050 ;
        RECT 502.950 149.400 517.050 150.600 ;
        RECT 502.950 148.950 505.050 149.400 ;
        RECT 514.950 148.950 517.050 149.400 ;
        RECT 514.950 99.600 517.050 100.050 ;
        RECT 520.950 99.600 523.050 100.050 ;
        RECT 514.950 98.400 523.050 99.600 ;
        RECT 514.950 97.950 517.050 98.400 ;
        RECT 520.950 97.950 523.050 98.400 ;
        RECT 520.950 3.600 523.050 4.050 ;
        RECT 544.950 3.600 547.050 4.050 ;
        RECT 520.950 2.400 547.050 3.600 ;
        RECT 520.950 1.950 523.050 2.400 ;
        RECT 544.950 1.950 547.050 2.400 ;
    END
  END hsync
  PIN p_tick
    PORT
      LAYER metal1 ;
        RECT 580.950 273.450 583.050 274.050 ;
        RECT 580.950 272.550 585.450 273.450 ;
        RECT 580.950 271.950 583.050 272.550 ;
        RECT 584.550 265.050 585.450 272.550 ;
        RECT 583.950 262.950 586.050 265.050 ;
      LAYER metal2 ;
        RECT 577.950 409.950 580.050 412.050 ;
        RECT 578.400 397.050 579.450 409.950 ;
        RECT 550.950 394.950 553.050 397.050 ;
        RECT 577.950 394.950 580.050 397.050 ;
        RECT 551.400 280.050 552.450 394.950 ;
        RECT 550.950 277.950 553.050 280.050 ;
        RECT 580.950 277.950 583.050 280.050 ;
        RECT 581.400 274.050 582.450 277.950 ;
        RECT 580.950 271.950 583.050 274.050 ;
        RECT 583.950 262.950 586.050 265.050 ;
        RECT 584.400 249.450 585.450 262.950 ;
        RECT 584.400 248.400 588.450 249.450 ;
        RECT 587.400 193.050 588.450 248.400 ;
        RECT 556.950 190.950 559.050 193.050 ;
        RECT 586.950 190.950 589.050 193.050 ;
        RECT 557.400 151.050 558.450 190.950 ;
        RECT 556.950 148.950 559.050 151.050 ;
        RECT 583.950 148.950 586.050 151.050 ;
        RECT 584.400 103.050 585.450 148.950 ;
        RECT 556.950 100.950 559.050 103.050 ;
        RECT 583.950 100.950 586.050 103.050 ;
        RECT 557.400 4.050 558.450 100.950 ;
        RECT 556.950 1.950 559.050 4.050 ;
        RECT 574.950 1.950 577.050 4.050 ;
        RECT 575.400 -3.600 576.450 1.950 ;
      LAYER metal3 ;
        RECT 550.950 396.600 553.050 397.050 ;
        RECT 577.950 396.600 580.050 397.050 ;
        RECT 550.950 395.400 580.050 396.600 ;
        RECT 550.950 394.950 553.050 395.400 ;
        RECT 577.950 394.950 580.050 395.400 ;
        RECT 550.950 279.600 553.050 280.050 ;
        RECT 580.950 279.600 583.050 280.050 ;
        RECT 550.950 278.400 583.050 279.600 ;
        RECT 550.950 277.950 553.050 278.400 ;
        RECT 580.950 277.950 583.050 278.400 ;
        RECT 556.950 192.600 559.050 193.050 ;
        RECT 586.950 192.600 589.050 193.050 ;
        RECT 556.950 191.400 589.050 192.600 ;
        RECT 556.950 190.950 559.050 191.400 ;
        RECT 586.950 190.950 589.050 191.400 ;
        RECT 556.950 150.600 559.050 151.050 ;
        RECT 583.950 150.600 586.050 151.050 ;
        RECT 556.950 149.400 586.050 150.600 ;
        RECT 556.950 148.950 559.050 149.400 ;
        RECT 583.950 148.950 586.050 149.400 ;
        RECT 556.950 102.600 559.050 103.050 ;
        RECT 583.950 102.600 586.050 103.050 ;
        RECT 556.950 101.400 586.050 102.600 ;
        RECT 556.950 100.950 559.050 101.400 ;
        RECT 583.950 100.950 586.050 101.400 ;
        RECT 556.950 3.600 559.050 4.050 ;
        RECT 574.950 3.600 577.050 4.050 ;
        RECT 556.950 2.400 577.050 3.600 ;
        RECT 556.950 1.950 559.050 2.400 ;
        RECT 574.950 1.950 577.050 2.400 ;
    END
  END p_tick
  PIN reset
    PORT
      LAYER metal2 ;
        RECT 422.400 832.050 423.450 837.450 ;
        RECT 379.950 829.950 382.050 832.050 ;
        RECT 421.950 829.950 424.050 832.050 ;
        RECT 376.950 816.450 379.050 817.050 ;
        RECT 380.400 816.450 381.450 829.950 ;
        RECT 376.950 815.400 381.450 816.450 ;
        RECT 376.950 814.950 379.050 815.400 ;
        RECT 380.400 807.450 381.450 815.400 ;
        RECT 377.400 806.400 381.450 807.450 ;
        RECT 377.400 771.450 378.450 806.400 ;
        RECT 379.950 771.450 382.050 772.050 ;
        RECT 377.400 770.400 382.050 771.450 ;
        RECT 379.950 769.950 382.050 770.400 ;
      LAYER metal3 ;
        RECT 379.950 831.600 382.050 832.050 ;
        RECT 421.950 831.600 424.050 832.050 ;
        RECT 379.950 830.400 424.050 831.600 ;
        RECT 379.950 829.950 382.050 830.400 ;
        RECT 421.950 829.950 424.050 830.400 ;
    END
  END reset
  PIN rgb
    PORT
      LAYER metal1 ;
        RECT 514.950 276.450 517.050 277.050 ;
        RECT 512.550 275.550 517.050 276.450 ;
        RECT 512.550 273.450 513.450 275.550 ;
        RECT 514.950 274.950 517.050 275.550 ;
        RECT 509.550 272.550 513.450 273.450 ;
        RECT 505.950 264.450 508.050 265.050 ;
        RECT 509.550 264.450 510.450 272.550 ;
        RECT 505.950 263.550 510.450 264.450 ;
        RECT 505.950 262.950 508.050 263.550 ;
        RECT 520.950 240.450 523.050 241.050 ;
        RECT 520.950 239.550 525.450 240.450 ;
        RECT 520.950 238.950 523.050 239.550 ;
        RECT 524.550 234.450 525.450 239.550 ;
        RECT 532.950 234.450 535.050 235.050 ;
        RECT 524.550 233.550 535.050 234.450 ;
        RECT 532.950 232.950 535.050 233.550 ;
      LAYER metal2 ;
        RECT 535.950 337.950 538.050 340.050 ;
        RECT 536.400 325.050 537.450 337.950 ;
        RECT 511.950 322.950 514.050 325.050 ;
        RECT 535.950 322.950 538.050 325.050 ;
        RECT 512.400 300.450 513.450 322.950 ;
        RECT 512.400 299.400 516.450 300.450 ;
        RECT 515.400 277.050 516.450 299.400 ;
        RECT 514.950 274.950 517.050 277.050 ;
        RECT 505.950 262.950 508.050 265.050 ;
        RECT 506.400 259.050 507.450 262.950 ;
        RECT 505.950 256.950 508.050 259.050 ;
        RECT 520.950 256.950 523.050 259.050 ;
        RECT 521.400 241.050 522.450 256.950 ;
        RECT 520.950 238.950 523.050 241.050 ;
        RECT 532.950 232.950 535.050 235.050 ;
        RECT 533.400 187.050 534.450 232.950 ;
        RECT 517.950 184.950 520.050 187.050 ;
        RECT 532.950 184.950 535.050 187.050 ;
        RECT 518.400 145.050 519.450 184.950 ;
        RECT 517.950 142.950 520.050 145.050 ;
        RECT 565.950 142.950 568.050 145.050 ;
        RECT 566.400 99.450 567.450 142.950 ;
        RECT 566.400 98.400 570.450 99.450 ;
        RECT 569.400 73.050 570.450 98.400 ;
        RECT 562.950 70.950 565.050 73.050 ;
        RECT 568.950 70.950 571.050 73.050 ;
        RECT 563.400 31.050 564.450 70.950 ;
        RECT 538.950 28.950 541.050 31.050 ;
        RECT 562.950 28.950 565.050 31.050 ;
        RECT 539.400 13.050 540.450 28.950 ;
        RECT 532.950 10.950 535.050 13.050 ;
        RECT 538.950 10.950 541.050 13.050 ;
        RECT 533.400 -3.600 534.450 10.950 ;
      LAYER metal3 ;
        RECT 511.950 324.600 514.050 325.050 ;
        RECT 535.950 324.600 538.050 325.050 ;
        RECT 511.950 323.400 538.050 324.600 ;
        RECT 511.950 322.950 514.050 323.400 ;
        RECT 535.950 322.950 538.050 323.400 ;
        RECT 505.950 258.600 508.050 259.050 ;
        RECT 520.950 258.600 523.050 259.050 ;
        RECT 505.950 257.400 523.050 258.600 ;
        RECT 505.950 256.950 508.050 257.400 ;
        RECT 520.950 256.950 523.050 257.400 ;
        RECT 517.950 186.600 520.050 187.050 ;
        RECT 532.950 186.600 535.050 187.050 ;
        RECT 517.950 185.400 535.050 186.600 ;
        RECT 517.950 184.950 520.050 185.400 ;
        RECT 532.950 184.950 535.050 185.400 ;
        RECT 517.950 144.600 520.050 145.050 ;
        RECT 565.950 144.600 568.050 145.050 ;
        RECT 517.950 143.400 568.050 144.600 ;
        RECT 517.950 142.950 520.050 143.400 ;
        RECT 565.950 142.950 568.050 143.400 ;
        RECT 562.950 72.600 565.050 73.050 ;
        RECT 568.950 72.600 571.050 73.050 ;
        RECT 562.950 71.400 571.050 72.600 ;
        RECT 562.950 70.950 565.050 71.400 ;
        RECT 568.950 70.950 571.050 71.400 ;
        RECT 538.950 30.600 541.050 31.050 ;
        RECT 562.950 30.600 565.050 31.050 ;
        RECT 538.950 29.400 565.050 30.600 ;
        RECT 538.950 28.950 541.050 29.400 ;
        RECT 562.950 28.950 565.050 29.400 ;
        RECT 532.950 12.600 535.050 13.050 ;
        RECT 538.950 12.600 541.050 13.050 ;
        RECT 532.950 11.400 541.050 12.600 ;
        RECT 532.950 10.950 535.050 11.400 ;
        RECT 538.950 10.950 541.050 11.400 ;
    END
  END rgb
  PIN up
    PORT
      LAYER metal2 ;
        RECT 470.400 829.050 471.450 837.450 ;
        RECT 469.950 826.950 472.050 829.050 ;
        RECT 496.950 826.950 499.050 829.050 ;
        RECT 497.400 799.050 498.450 826.950 ;
        RECT 496.950 796.950 499.050 799.050 ;
        RECT 703.950 796.950 706.050 799.050 ;
        RECT 704.400 742.050 705.450 796.950 ;
        RECT 703.950 739.950 706.050 742.050 ;
        RECT 709.950 739.950 712.050 742.050 ;
        RECT 710.400 544.050 711.450 739.950 ;
        RECT 667.950 541.950 670.050 544.050 ;
        RECT 709.950 541.950 712.050 544.050 ;
        RECT 668.400 483.450 669.450 541.950 ;
        RECT 665.400 482.400 669.450 483.450 ;
        RECT 665.400 451.050 666.450 482.400 ;
        RECT 664.950 448.950 667.050 451.050 ;
        RECT 688.950 448.950 691.050 451.050 ;
        RECT 689.400 409.050 690.450 448.950 ;
        RECT 688.950 406.950 691.050 409.050 ;
        RECT 709.950 406.950 712.050 409.050 ;
        RECT 710.400 367.050 711.450 406.950 ;
        RECT 709.950 364.950 712.050 367.050 ;
        RECT 733.950 364.950 736.050 367.050 ;
        RECT 734.400 328.050 735.450 364.950 ;
        RECT 721.950 325.950 724.050 328.050 ;
        RECT 733.950 325.950 736.050 328.050 ;
        RECT 722.400 277.050 723.450 325.950 ;
        RECT 721.950 274.950 724.050 277.050 ;
        RECT 718.950 268.950 721.050 271.050 ;
        RECT 719.400 253.050 720.450 268.950 ;
        RECT 703.950 250.950 706.050 253.050 ;
        RECT 718.950 250.950 721.050 253.050 ;
        RECT 704.400 226.050 705.450 250.950 ;
        RECT 688.950 223.950 691.050 226.050 ;
        RECT 703.950 223.950 706.050 226.050 ;
        RECT 689.400 193.050 690.450 223.950 ;
        RECT 667.950 190.950 670.050 193.050 ;
        RECT 688.950 190.950 691.050 193.050 ;
        RECT 668.400 112.050 669.450 190.950 ;
        RECT 655.950 109.950 658.050 112.050 ;
        RECT 667.950 109.950 670.050 112.050 ;
        RECT 457.950 94.950 460.050 97.050 ;
        RECT 458.400 94.050 459.450 94.950 ;
        RECT 457.950 91.950 460.050 94.050 ;
        RECT 481.950 88.950 484.050 91.050 ;
        RECT 482.400 70.050 483.450 88.950 ;
        RECT 656.400 70.050 657.450 109.950 ;
        RECT 481.950 67.950 484.050 70.050 ;
        RECT 655.950 67.950 658.050 70.050 ;
      LAYER metal3 ;
        RECT 469.950 828.600 472.050 829.050 ;
        RECT 496.950 828.600 499.050 829.050 ;
        RECT 469.950 827.400 499.050 828.600 ;
        RECT 469.950 826.950 472.050 827.400 ;
        RECT 496.950 826.950 499.050 827.400 ;
        RECT 496.950 798.600 499.050 799.050 ;
        RECT 703.950 798.600 706.050 799.050 ;
        RECT 496.950 797.400 706.050 798.600 ;
        RECT 496.950 796.950 499.050 797.400 ;
        RECT 703.950 796.950 706.050 797.400 ;
        RECT 703.950 741.600 706.050 742.050 ;
        RECT 709.950 741.600 712.050 742.050 ;
        RECT 703.950 740.400 712.050 741.600 ;
        RECT 703.950 739.950 706.050 740.400 ;
        RECT 709.950 739.950 712.050 740.400 ;
        RECT 667.950 543.600 670.050 544.050 ;
        RECT 709.950 543.600 712.050 544.050 ;
        RECT 667.950 542.400 712.050 543.600 ;
        RECT 667.950 541.950 670.050 542.400 ;
        RECT 709.950 541.950 712.050 542.400 ;
        RECT 664.950 450.600 667.050 451.050 ;
        RECT 688.950 450.600 691.050 451.050 ;
        RECT 664.950 449.400 691.050 450.600 ;
        RECT 664.950 448.950 667.050 449.400 ;
        RECT 688.950 448.950 691.050 449.400 ;
        RECT 688.950 408.600 691.050 409.050 ;
        RECT 709.950 408.600 712.050 409.050 ;
        RECT 688.950 407.400 712.050 408.600 ;
        RECT 688.950 406.950 691.050 407.400 ;
        RECT 709.950 406.950 712.050 407.400 ;
        RECT 709.950 366.600 712.050 367.050 ;
        RECT 733.950 366.600 736.050 367.050 ;
        RECT 709.950 365.400 736.050 366.600 ;
        RECT 709.950 364.950 712.050 365.400 ;
        RECT 733.950 364.950 736.050 365.400 ;
        RECT 721.950 327.600 724.050 328.050 ;
        RECT 733.950 327.600 736.050 328.050 ;
        RECT 721.950 326.400 736.050 327.600 ;
        RECT 721.950 325.950 724.050 326.400 ;
        RECT 733.950 325.950 736.050 326.400 ;
        RECT 721.950 274.950 724.050 277.050 ;
        RECT 718.950 270.600 721.050 271.050 ;
        RECT 722.400 270.600 723.600 274.950 ;
        RECT 718.950 269.400 723.600 270.600 ;
        RECT 718.950 268.950 721.050 269.400 ;
        RECT 703.950 252.600 706.050 253.050 ;
        RECT 718.950 252.600 721.050 253.050 ;
        RECT 703.950 251.400 721.050 252.600 ;
        RECT 703.950 250.950 706.050 251.400 ;
        RECT 718.950 250.950 721.050 251.400 ;
        RECT 688.950 225.600 691.050 226.050 ;
        RECT 703.950 225.600 706.050 226.050 ;
        RECT 688.950 224.400 706.050 225.600 ;
        RECT 688.950 223.950 691.050 224.400 ;
        RECT 703.950 223.950 706.050 224.400 ;
        RECT 667.950 192.600 670.050 193.050 ;
        RECT 688.950 192.600 691.050 193.050 ;
        RECT 667.950 191.400 691.050 192.600 ;
        RECT 667.950 190.950 670.050 191.400 ;
        RECT 688.950 190.950 691.050 191.400 ;
        RECT 655.950 111.600 658.050 112.050 ;
        RECT 667.950 111.600 670.050 112.050 ;
        RECT 655.950 110.400 670.050 111.600 ;
        RECT 655.950 109.950 658.050 110.400 ;
        RECT 667.950 109.950 670.050 110.400 ;
        RECT 457.950 96.600 460.050 97.050 ;
        RECT 457.950 95.400 474.600 96.600 ;
        RECT 457.950 94.950 460.050 95.400 ;
        RECT 473.400 93.600 474.600 95.400 ;
        RECT 473.400 92.400 480.600 93.600 ;
        RECT 479.400 90.600 480.600 92.400 ;
        RECT 481.950 90.600 484.050 91.050 ;
        RECT 479.400 89.400 484.050 90.600 ;
        RECT 481.950 88.950 484.050 89.400 ;
        RECT 481.950 69.600 484.050 70.050 ;
        RECT 655.950 69.600 658.050 70.050 ;
        RECT 481.950 68.400 658.050 69.600 ;
        RECT 481.950 67.950 484.050 68.400 ;
        RECT 655.950 67.950 658.050 68.400 ;
    END
  END up
  PIN vsync
    PORT
      LAYER metal2 ;
        RECT 517.950 388.950 520.050 391.050 ;
        RECT 553.950 388.950 556.050 391.050 ;
        RECT 518.400 385.050 519.450 388.950 ;
        RECT 517.950 382.950 520.050 385.050 ;
        RECT 554.400 373.050 555.450 388.950 ;
        RECT 544.950 370.950 547.050 373.050 ;
        RECT 553.950 370.950 556.050 373.050 ;
        RECT 545.400 319.050 546.450 370.950 ;
        RECT 544.950 316.950 547.050 319.050 ;
        RECT 559.950 316.950 562.050 319.050 ;
        RECT 560.400 301.050 561.450 316.950 ;
        RECT 559.950 298.950 562.050 301.050 ;
        RECT 625.950 298.950 628.050 301.050 ;
        RECT 626.400 246.450 627.450 298.950 ;
        RECT 626.400 245.400 630.450 246.450 ;
        RECT 629.400 244.050 630.450 245.400 ;
        RECT 628.950 241.950 631.050 244.050 ;
        RECT 646.950 232.950 649.050 235.050 ;
        RECT 647.400 205.050 648.450 232.950 ;
        RECT 646.950 202.950 649.050 205.050 ;
        RECT 658.950 202.950 661.050 205.050 ;
        RECT 659.400 193.050 660.450 202.950 ;
        RECT 646.950 190.950 649.050 193.050 ;
        RECT 658.950 190.950 661.050 193.050 ;
        RECT 647.400 142.050 648.450 190.950 ;
        RECT 637.950 139.950 640.050 142.050 ;
        RECT 646.950 139.950 649.050 142.050 ;
        RECT 638.400 69.450 639.450 139.950 ;
        RECT 635.400 68.400 639.450 69.450 ;
        RECT 635.400 33.450 636.450 68.400 ;
        RECT 632.400 32.400 636.450 33.450 ;
        RECT 632.400 7.050 633.450 32.400 ;
        RECT 538.950 4.950 541.050 7.050 ;
        RECT 631.950 4.950 634.050 7.050 ;
        RECT 539.400 -3.600 540.450 4.950 ;
      LAYER metal3 ;
        RECT 517.950 390.600 520.050 391.050 ;
        RECT 553.950 390.600 556.050 391.050 ;
        RECT 517.950 389.400 556.050 390.600 ;
        RECT 517.950 388.950 520.050 389.400 ;
        RECT 553.950 388.950 556.050 389.400 ;
        RECT 544.950 372.600 547.050 373.050 ;
        RECT 553.950 372.600 556.050 373.050 ;
        RECT 544.950 371.400 556.050 372.600 ;
        RECT 544.950 370.950 547.050 371.400 ;
        RECT 553.950 370.950 556.050 371.400 ;
        RECT 544.950 318.600 547.050 319.050 ;
        RECT 559.950 318.600 562.050 319.050 ;
        RECT 544.950 317.400 562.050 318.600 ;
        RECT 544.950 316.950 547.050 317.400 ;
        RECT 559.950 316.950 562.050 317.400 ;
        RECT 559.950 300.600 562.050 301.050 ;
        RECT 625.950 300.600 628.050 301.050 ;
        RECT 559.950 299.400 628.050 300.600 ;
        RECT 559.950 298.950 562.050 299.400 ;
        RECT 625.950 298.950 628.050 299.400 ;
        RECT 628.950 243.600 631.050 244.050 ;
        RECT 628.950 242.400 633.600 243.600 ;
        RECT 628.950 241.950 631.050 242.400 ;
        RECT 632.400 237.600 633.600 242.400 ;
        RECT 632.400 236.400 648.600 237.600 ;
        RECT 647.400 235.050 648.600 236.400 ;
        RECT 646.950 232.950 649.050 235.050 ;
        RECT 646.950 204.600 649.050 205.050 ;
        RECT 658.950 204.600 661.050 205.050 ;
        RECT 646.950 203.400 661.050 204.600 ;
        RECT 646.950 202.950 649.050 203.400 ;
        RECT 658.950 202.950 661.050 203.400 ;
        RECT 646.950 192.600 649.050 193.050 ;
        RECT 658.950 192.600 661.050 193.050 ;
        RECT 646.950 191.400 661.050 192.600 ;
        RECT 646.950 190.950 649.050 191.400 ;
        RECT 658.950 190.950 661.050 191.400 ;
        RECT 637.950 141.600 640.050 142.050 ;
        RECT 646.950 141.600 649.050 142.050 ;
        RECT 637.950 140.400 649.050 141.600 ;
        RECT 637.950 139.950 640.050 140.400 ;
        RECT 646.950 139.950 649.050 140.400 ;
        RECT 538.950 6.600 541.050 7.050 ;
        RECT 631.950 6.600 634.050 7.050 ;
        RECT 538.950 5.400 634.050 6.600 ;
        RECT 538.950 4.950 541.050 5.400 ;
        RECT 631.950 4.950 634.050 5.400 ;
    END
  END vsync
  OBS
      LAYER metal1 ;
        RECT 7.650 821.400 9.450 827.250 ;
        RECT 8.250 819.300 9.450 821.400 ;
        RECT 10.650 822.300 12.450 827.250 ;
        RECT 13.650 823.200 15.450 827.250 ;
        RECT 16.650 822.300 18.450 827.250 ;
        RECT 10.650 820.950 18.450 822.300 ;
        RECT 26.850 820.200 28.650 827.250 ;
        RECT 31.350 821.400 33.150 827.250 ;
        RECT 38.550 824.400 40.350 827.250 ;
        RECT 41.550 824.400 43.350 827.250 ;
        RECT 44.550 824.400 46.350 827.250 ;
        RECT 26.850 819.300 30.450 820.200 ;
        RECT 8.250 818.250 12.000 819.300 ;
        RECT 10.950 814.950 12.150 818.250 ;
        RECT 14.100 816.150 15.900 817.950 ;
        RECT 10.950 812.850 13.050 814.950 ;
        RECT 13.950 814.050 16.050 816.150 ;
        RECT 16.950 812.850 19.050 814.950 ;
        RECT 26.100 813.150 27.900 814.950 ;
        RECT 7.950 809.850 10.050 811.950 ;
        RECT 8.250 808.050 10.050 809.850 ;
        RECT 11.850 807.600 13.050 812.850 ;
        RECT 17.100 811.050 18.900 812.850 ;
        RECT 25.950 811.050 28.050 813.150 ;
        RECT 29.250 811.950 30.450 819.300 ;
        RECT 42.000 817.950 43.050 824.400 ;
        RECT 40.950 815.850 43.050 817.950 ;
        RECT 32.100 813.150 33.900 814.950 ;
        RECT 28.950 809.850 31.050 811.950 ;
        RECT 31.950 811.050 34.050 813.150 ;
        RECT 37.950 812.850 40.050 814.950 ;
        RECT 38.100 811.050 39.900 812.850 ;
        RECT 8.400 795.750 10.200 801.600 ;
        RECT 11.700 795.750 13.500 807.600 ;
        RECT 15.900 795.750 17.700 807.600 ;
        RECT 29.250 801.600 30.450 809.850 ;
        RECT 42.000 808.650 43.050 815.850 ;
        RECT 50.700 821.400 52.500 827.250 ;
        RECT 56.100 821.400 57.900 827.250 ;
        RECT 61.500 821.400 63.300 827.250 ;
        RECT 65.700 824.400 67.500 827.250 ;
        RECT 68.700 824.400 70.500 827.250 ;
        RECT 71.700 824.400 73.500 827.250 ;
        RECT 74.700 824.400 76.500 827.250 ;
        RECT 65.700 823.050 67.050 824.400 ;
        RECT 68.700 823.050 70.050 824.400 ;
        RECT 71.700 823.050 73.050 824.400 ;
        RECT 79.200 823.500 81.000 827.250 ;
        RECT 82.200 824.400 84.000 827.250 ;
        RECT 85.200 823.500 87.000 827.250 ;
        RECT 50.700 817.800 51.900 821.400 ;
        RECT 61.800 820.500 63.300 821.400 ;
        RECT 54.900 819.300 63.300 820.500 ;
        RECT 64.950 820.950 67.050 823.050 ;
        RECT 67.950 820.950 70.050 823.050 ;
        RECT 70.950 820.950 73.050 823.050 ;
        RECT 76.500 822.750 78.300 823.200 ;
        RECT 74.250 821.400 78.300 822.750 ;
        RECT 79.200 821.700 82.050 823.500 ;
        RECT 79.950 821.400 82.050 821.700 ;
        RECT 84.150 821.700 87.000 823.500 ;
        RECT 88.950 823.500 90.750 827.250 ;
        RECT 91.950 823.500 93.750 827.250 ;
        RECT 94.950 823.500 96.750 827.250 ;
        RECT 84.150 821.400 86.250 821.700 ;
        RECT 88.950 821.400 91.050 823.500 ;
        RECT 91.950 821.400 94.050 823.500 ;
        RECT 94.950 821.400 97.050 823.500 ;
        RECT 99.600 822.600 101.400 827.250 ;
        RECT 99.600 821.400 103.800 822.600 ;
        RECT 105.150 821.400 106.950 827.250 ;
        RECT 110.550 821.400 112.350 827.250 ;
        RECT 54.900 818.700 56.700 819.300 ;
        RECT 64.950 817.800 66.000 820.950 ;
        RECT 74.250 820.050 75.150 821.400 ;
        RECT 70.050 819.900 75.150 820.050 ;
        RECT 50.700 816.900 66.000 817.800 ;
        RECT 67.500 819.150 75.150 819.900 ;
        RECT 67.500 818.700 71.850 819.150 ;
        RECT 83.100 818.700 90.000 820.500 ;
        RECT 90.900 818.700 97.650 820.500 ;
        RECT 43.950 812.850 46.050 814.950 ;
        RECT 44.100 811.050 45.900 812.850 ;
        RECT 42.000 807.600 44.550 808.650 ;
        RECT 25.650 795.750 27.450 801.600 ;
        RECT 28.650 795.750 30.450 801.600 ;
        RECT 31.650 795.750 33.450 801.600 ;
        RECT 38.550 795.750 40.350 807.600 ;
        RECT 42.750 795.750 44.550 807.600 ;
        RECT 50.700 803.400 51.900 816.900 ;
        RECT 53.100 814.950 64.950 816.000 ;
        RECT 67.500 815.250 68.550 818.700 ;
        RECT 70.050 818.250 71.850 818.700 ;
        RECT 76.950 817.650 79.050 817.950 ;
        RECT 88.950 817.800 90.000 818.700 ;
        RECT 102.300 817.800 103.800 821.400 ;
        RECT 75.150 815.850 79.050 817.650 ;
        RECT 80.400 816.450 88.050 817.800 ;
        RECT 88.950 816.750 98.850 817.800 ;
        RECT 53.100 813.150 54.900 814.950 ;
        RECT 52.950 811.050 55.050 813.150 ;
        RECT 63.750 812.550 64.950 814.950 ;
        RECT 66.750 813.450 68.550 815.250 ;
        RECT 80.400 814.950 81.450 816.450 ;
        RECT 87.150 815.700 88.050 816.450 ;
        RECT 69.450 814.050 81.450 814.950 ;
        RECT 69.450 812.550 70.500 814.050 ;
        RECT 82.350 813.750 86.250 815.550 ;
        RECT 87.150 814.650 96.750 815.700 ;
        RECT 84.150 813.450 86.250 813.750 ;
        RECT 58.950 811.650 61.050 811.950 ;
        RECT 63.750 811.650 70.500 812.550 ;
        RECT 71.400 812.550 73.200 813.150 ;
        RECT 79.950 812.550 82.050 812.850 ;
        RECT 71.400 811.950 82.050 812.550 ;
        RECT 92.700 811.950 94.500 813.750 ;
        RECT 58.950 810.450 62.850 811.650 ;
        RECT 71.400 811.350 94.500 811.950 ;
        RECT 79.950 810.750 94.500 811.350 ;
        RECT 95.850 813.000 96.750 814.650 ;
        RECT 97.800 814.950 98.850 816.750 ;
        RECT 102.300 816.000 110.100 817.800 ;
        RECT 97.800 813.900 106.050 814.950 ;
        RECT 95.850 811.200 102.900 813.000 ;
        RECT 58.950 809.850 72.900 810.450 ;
        RECT 103.950 809.850 106.050 813.900 ;
        RECT 59.250 809.550 99.000 809.850 ;
        RECT 70.950 808.650 99.000 809.550 ;
        RECT 108.450 808.650 110.250 809.250 ;
        RECT 58.500 808.050 60.300 808.650 ;
        RECT 67.950 808.050 70.050 808.350 ;
        RECT 58.500 806.850 70.050 808.050 ;
        RECT 67.950 806.250 70.050 806.850 ;
        RECT 70.950 806.400 91.050 807.750 ;
        RECT 55.200 805.350 57.000 806.100 ;
        RECT 70.950 805.350 72.900 806.400 ;
        RECT 88.950 805.650 91.050 806.400 ;
        RECT 94.950 806.550 97.050 807.750 ;
        RECT 97.950 807.450 110.250 808.650 ;
        RECT 111.150 806.550 112.350 821.400 ;
        RECT 94.950 805.650 112.350 806.550 ;
        RECT 114.450 824.400 116.250 827.250 ;
        RECT 117.450 824.400 119.250 827.250 ;
        RECT 127.650 824.400 129.450 827.250 ;
        RECT 130.650 824.400 132.450 827.250 ;
        RECT 140.250 824.400 142.350 827.250 ;
        RECT 143.550 824.400 145.350 827.250 ;
        RECT 146.550 824.400 148.350 827.250 ;
        RECT 149.550 824.400 151.350 827.250 ;
        RECT 114.450 816.150 115.950 824.400 ;
        RECT 128.400 816.150 129.600 824.400 ;
        RECT 144.300 823.500 145.350 824.400 ;
        RECT 150.300 823.500 151.350 824.400 ;
        RECT 144.300 822.600 155.100 823.500 ;
        RECT 114.450 814.050 118.050 816.150 ;
        RECT 127.950 814.050 130.050 816.150 ;
        RECT 130.950 815.850 133.050 817.950 ;
        RECT 146.100 816.150 147.900 817.950 ;
        RECT 153.900 816.150 155.100 822.600 ;
        RECT 173.850 820.200 175.650 827.250 ;
        RECT 178.350 821.400 180.150 827.250 ;
        RECT 185.850 820.200 187.650 827.250 ;
        RECT 190.350 821.400 192.150 827.250 ;
        RECT 197.850 821.400 199.650 827.250 ;
        RECT 202.350 820.200 204.150 827.250 ;
        RECT 215.550 822.300 217.350 827.250 ;
        RECT 218.550 823.200 220.350 827.250 ;
        RECT 221.550 822.300 223.350 827.250 ;
        RECT 215.550 820.950 223.350 822.300 ;
        RECT 224.550 821.400 226.350 827.250 ;
        RECT 230.550 824.400 232.350 827.250 ;
        RECT 233.550 824.400 235.350 827.250 ;
        RECT 242.550 824.400 244.350 827.250 ;
        RECT 245.550 824.400 247.350 827.250 ;
        RECT 257.550 824.400 259.350 827.250 ;
        RECT 260.550 824.400 262.350 827.250 ;
        RECT 263.550 824.400 265.350 827.250 ;
        RECT 173.850 819.300 177.450 820.200 ;
        RECT 185.850 819.300 189.450 820.200 ;
        RECT 131.100 814.050 132.900 815.850 ;
        RECT 55.200 804.300 72.900 805.350 ;
        RECT 50.700 802.500 54.750 803.400 ;
        RECT 53.700 801.600 54.750 802.500 ;
        RECT 50.700 795.750 52.500 801.600 ;
        RECT 53.700 795.750 55.500 801.600 ;
        RECT 56.700 795.750 58.500 801.600 ;
        RECT 59.700 795.750 61.500 804.300 ;
        RECT 79.950 804.150 82.050 804.600 ;
        RECT 79.650 802.500 82.050 804.150 ;
        RECT 84.000 802.800 87.900 804.600 ;
        RECT 84.000 802.500 87.000 802.800 ;
        RECT 64.950 799.950 67.050 802.050 ;
        RECT 67.950 799.950 70.050 802.050 ;
        RECT 70.950 801.600 73.050 802.050 ;
        RECT 79.650 801.600 81.000 802.500 ;
        RECT 70.950 799.950 73.500 801.600 ;
        RECT 62.700 795.750 64.500 799.050 ;
        RECT 65.850 798.600 67.050 799.950 ;
        RECT 69.150 798.600 70.050 799.950 ;
        RECT 72.300 798.600 73.500 799.950 ;
        RECT 65.850 795.750 68.250 798.600 ;
        RECT 69.150 795.750 71.250 798.600 ;
        RECT 72.300 795.750 74.250 798.600 ;
        RECT 75.450 795.750 77.250 801.600 ;
        RECT 79.200 795.750 81.000 801.600 ;
        RECT 82.200 795.750 84.000 801.600 ;
        RECT 85.200 795.750 87.000 802.500 ;
        RECT 89.100 798.600 90.450 805.650 ;
        RECT 98.850 804.150 100.650 804.300 ;
        RECT 91.950 802.950 100.650 804.150 ;
        RECT 105.600 803.700 107.400 804.300 ;
        RECT 91.950 802.050 94.050 802.950 ;
        RECT 98.850 802.500 100.650 802.950 ;
        RECT 101.700 802.500 107.400 803.700 ;
        RECT 88.950 795.750 90.750 798.600 ;
        RECT 91.950 795.750 93.750 802.050 ;
        RECT 95.100 799.800 97.200 801.900 ;
        RECT 95.100 798.600 96.600 799.800 ;
        RECT 94.950 795.750 96.750 798.600 ;
        RECT 98.700 795.750 100.500 801.600 ;
        RECT 101.700 795.750 103.500 802.500 ;
        RECT 108.300 801.600 109.500 805.650 ;
        RECT 114.450 801.600 115.950 814.050 ;
        RECT 128.400 801.600 129.600 814.050 ;
        RECT 139.950 812.850 142.050 814.950 ;
        RECT 145.950 814.050 148.050 816.150 ;
        RECT 148.950 812.850 151.050 814.950 ;
        RECT 153.900 814.050 157.050 816.150 ;
        RECT 140.100 811.050 141.900 812.850 ;
        RECT 149.100 811.050 150.900 812.850 ;
        RECT 153.900 808.800 155.100 814.050 ;
        RECT 173.100 813.150 174.900 814.950 ;
        RECT 172.950 811.050 175.050 813.150 ;
        RECT 176.250 811.950 177.450 819.300 ;
        RECT 179.100 813.150 180.900 814.950 ;
        RECT 185.100 813.150 186.900 814.950 ;
        RECT 175.950 809.850 178.050 811.950 ;
        RECT 178.950 811.050 181.050 813.150 ;
        RECT 184.950 811.050 187.050 813.150 ;
        RECT 188.250 811.950 189.450 819.300 ;
        RECT 200.550 819.300 204.150 820.200 ;
        RECT 224.550 819.300 225.750 821.400 ;
        RECT 191.100 813.150 192.900 814.950 ;
        RECT 197.100 813.150 198.900 814.950 ;
        RECT 187.950 809.850 190.050 811.950 ;
        RECT 190.950 811.050 193.050 813.150 ;
        RECT 196.950 811.050 199.050 813.150 ;
        RECT 200.550 811.950 201.750 819.300 ;
        RECT 222.000 818.250 225.750 819.300 ;
        RECT 218.100 816.150 219.900 817.950 ;
        RECT 203.100 813.150 204.900 814.950 ;
        RECT 199.950 809.850 202.050 811.950 ;
        RECT 202.950 811.050 205.050 813.150 ;
        RECT 214.950 812.850 217.050 814.950 ;
        RECT 217.950 814.050 220.050 816.150 ;
        RECT 221.850 814.950 223.050 818.250 ;
        RECT 229.950 815.850 232.050 817.950 ;
        RECT 233.400 816.150 234.600 824.400 ;
        RECT 220.950 812.850 223.050 814.950 ;
        RECT 230.100 814.050 231.900 815.850 ;
        RECT 232.950 814.050 235.050 816.150 ;
        RECT 241.950 815.850 244.050 817.950 ;
        RECT 245.400 816.150 246.600 824.400 ;
        RECT 261.000 817.950 262.050 824.400 ;
        RECT 242.100 814.050 243.900 815.850 ;
        RECT 244.950 814.050 247.050 816.150 ;
        RECT 259.950 815.850 262.050 817.950 ;
        RECT 215.100 811.050 216.900 812.850 ;
        RECT 153.900 807.600 157.350 808.800 ;
        RECT 137.550 805.500 145.350 806.400 ;
        RECT 104.700 795.750 106.500 801.600 ;
        RECT 107.700 795.750 109.500 801.600 ;
        RECT 110.700 795.750 112.500 801.600 ;
        RECT 114.450 795.750 116.250 801.600 ;
        RECT 117.450 795.750 119.250 801.600 ;
        RECT 127.650 795.750 129.450 801.600 ;
        RECT 130.650 795.750 132.450 801.600 ;
        RECT 137.550 795.750 139.350 805.500 ;
        RECT 140.550 795.750 142.350 804.600 ;
        RECT 143.550 796.500 145.350 805.500 ;
        RECT 146.550 805.200 154.950 806.100 ;
        RECT 146.550 797.400 148.350 805.200 ;
        RECT 149.550 796.500 151.350 804.300 ;
        RECT 143.550 795.750 151.350 796.500 ;
        RECT 153.150 796.500 154.950 805.200 ;
        RECT 156.150 805.200 157.350 807.600 ;
        RECT 156.150 797.400 157.950 805.200 ;
        RECT 159.150 796.500 160.950 805.800 ;
        RECT 176.250 801.600 177.450 809.850 ;
        RECT 188.250 801.600 189.450 809.850 ;
        RECT 200.550 801.600 201.750 809.850 ;
        RECT 220.950 807.600 222.150 812.850 ;
        RECT 223.950 809.850 226.050 811.950 ;
        RECT 223.950 808.050 225.750 809.850 ;
        RECT 153.150 795.750 160.950 796.500 ;
        RECT 172.650 795.750 174.450 801.600 ;
        RECT 175.650 795.750 177.450 801.600 ;
        RECT 178.650 795.750 180.450 801.600 ;
        RECT 184.650 795.750 186.450 801.600 ;
        RECT 187.650 795.750 189.450 801.600 ;
        RECT 190.650 795.750 192.450 801.600 ;
        RECT 197.550 795.750 199.350 801.600 ;
        RECT 200.550 795.750 202.350 801.600 ;
        RECT 203.550 795.750 205.350 801.600 ;
        RECT 216.300 795.750 218.100 807.600 ;
        RECT 220.500 795.750 222.300 807.600 ;
        RECT 233.400 801.600 234.600 814.050 ;
        RECT 245.400 801.600 246.600 814.050 ;
        RECT 256.950 812.850 259.050 814.950 ;
        RECT 257.100 811.050 258.900 812.850 ;
        RECT 261.000 808.650 262.050 815.850 ;
        RECT 269.700 821.400 271.500 827.250 ;
        RECT 275.100 821.400 276.900 827.250 ;
        RECT 280.500 821.400 282.300 827.250 ;
        RECT 284.700 824.400 286.500 827.250 ;
        RECT 287.700 824.400 289.500 827.250 ;
        RECT 290.700 824.400 292.500 827.250 ;
        RECT 293.700 824.400 295.500 827.250 ;
        RECT 284.700 823.050 286.050 824.400 ;
        RECT 287.700 823.050 289.050 824.400 ;
        RECT 290.700 823.050 292.050 824.400 ;
        RECT 298.200 823.500 300.000 827.250 ;
        RECT 301.200 824.400 303.000 827.250 ;
        RECT 304.200 823.500 306.000 827.250 ;
        RECT 269.700 817.800 270.900 821.400 ;
        RECT 280.800 820.500 282.300 821.400 ;
        RECT 273.900 819.300 282.300 820.500 ;
        RECT 283.950 820.950 286.050 823.050 ;
        RECT 286.950 820.950 289.050 823.050 ;
        RECT 289.950 820.950 292.050 823.050 ;
        RECT 295.500 822.750 297.300 823.200 ;
        RECT 293.250 821.400 297.300 822.750 ;
        RECT 298.200 821.700 301.050 823.500 ;
        RECT 298.950 821.400 301.050 821.700 ;
        RECT 303.150 821.700 306.000 823.500 ;
        RECT 307.950 823.500 309.750 827.250 ;
        RECT 310.950 823.500 312.750 827.250 ;
        RECT 313.950 823.500 315.750 827.250 ;
        RECT 303.150 821.400 305.250 821.700 ;
        RECT 307.950 821.400 310.050 823.500 ;
        RECT 310.950 821.400 313.050 823.500 ;
        RECT 313.950 821.400 316.050 823.500 ;
        RECT 318.600 822.600 320.400 827.250 ;
        RECT 318.600 821.400 322.800 822.600 ;
        RECT 324.150 821.400 325.950 827.250 ;
        RECT 329.550 821.400 331.350 827.250 ;
        RECT 273.900 818.700 275.700 819.300 ;
        RECT 283.950 817.800 285.000 820.950 ;
        RECT 293.250 820.050 294.150 821.400 ;
        RECT 289.050 819.900 294.150 820.050 ;
        RECT 269.700 816.900 285.000 817.800 ;
        RECT 286.500 819.150 294.150 819.900 ;
        RECT 286.500 818.700 290.850 819.150 ;
        RECT 302.100 818.700 309.000 820.500 ;
        RECT 309.900 818.700 316.650 820.500 ;
        RECT 262.950 812.850 265.050 814.950 ;
        RECT 263.100 811.050 264.900 812.850 ;
        RECT 261.000 807.600 263.550 808.650 ;
        RECT 223.800 795.750 225.600 801.600 ;
        RECT 230.550 795.750 232.350 801.600 ;
        RECT 233.550 795.750 235.350 801.600 ;
        RECT 242.550 795.750 244.350 801.600 ;
        RECT 245.550 795.750 247.350 801.600 ;
        RECT 257.550 795.750 259.350 807.600 ;
        RECT 261.750 795.750 263.550 807.600 ;
        RECT 269.700 803.400 270.900 816.900 ;
        RECT 272.100 814.950 283.950 816.000 ;
        RECT 286.500 815.250 287.550 818.700 ;
        RECT 289.050 818.250 290.850 818.700 ;
        RECT 295.950 817.650 298.050 817.950 ;
        RECT 307.950 817.800 309.000 818.700 ;
        RECT 321.300 817.800 322.800 821.400 ;
        RECT 294.150 815.850 298.050 817.650 ;
        RECT 299.400 816.450 307.050 817.800 ;
        RECT 307.950 816.750 317.850 817.800 ;
        RECT 272.100 813.150 273.900 814.950 ;
        RECT 271.950 811.050 274.050 813.150 ;
        RECT 282.750 812.550 283.950 814.950 ;
        RECT 285.750 813.450 287.550 815.250 ;
        RECT 299.400 814.950 300.450 816.450 ;
        RECT 306.150 815.700 307.050 816.450 ;
        RECT 288.450 814.050 300.450 814.950 ;
        RECT 288.450 812.550 289.500 814.050 ;
        RECT 301.350 813.750 305.250 815.550 ;
        RECT 306.150 814.650 315.750 815.700 ;
        RECT 303.150 813.450 305.250 813.750 ;
        RECT 277.950 811.650 280.050 811.950 ;
        RECT 282.750 811.650 289.500 812.550 ;
        RECT 290.400 812.550 292.200 813.150 ;
        RECT 298.950 812.550 301.050 812.850 ;
        RECT 290.400 811.950 301.050 812.550 ;
        RECT 311.700 811.950 313.500 813.750 ;
        RECT 277.950 810.450 281.850 811.650 ;
        RECT 290.400 811.350 313.500 811.950 ;
        RECT 298.950 810.750 313.500 811.350 ;
        RECT 314.850 813.000 315.750 814.650 ;
        RECT 316.800 814.950 317.850 816.750 ;
        RECT 321.300 816.000 329.100 817.800 ;
        RECT 316.800 813.900 325.050 814.950 ;
        RECT 314.850 811.200 321.900 813.000 ;
        RECT 277.950 809.850 291.900 810.450 ;
        RECT 322.950 809.850 325.050 813.900 ;
        RECT 278.250 809.550 318.000 809.850 ;
        RECT 289.950 808.650 318.000 809.550 ;
        RECT 327.450 808.650 329.250 809.250 ;
        RECT 277.500 808.050 279.300 808.650 ;
        RECT 286.950 808.050 289.050 808.350 ;
        RECT 277.500 806.850 289.050 808.050 ;
        RECT 286.950 806.250 289.050 806.850 ;
        RECT 289.950 806.400 310.050 807.750 ;
        RECT 274.200 805.350 276.000 806.100 ;
        RECT 289.950 805.350 291.900 806.400 ;
        RECT 307.950 805.650 310.050 806.400 ;
        RECT 313.950 806.550 316.050 807.750 ;
        RECT 316.950 807.450 329.250 808.650 ;
        RECT 330.150 806.550 331.350 821.400 ;
        RECT 313.950 805.650 331.350 806.550 ;
        RECT 333.450 824.400 335.250 827.250 ;
        RECT 336.450 824.400 338.250 827.250 ;
        RECT 347.550 824.400 349.350 827.250 ;
        RECT 333.450 816.150 334.950 824.400 ;
        RECT 348.150 820.500 349.350 824.400 ;
        RECT 350.850 821.400 352.650 827.250 ;
        RECT 353.850 821.400 355.650 827.250 ;
        RECT 367.650 821.400 369.450 827.250 ;
        RECT 370.650 821.400 372.450 827.250 ;
        RECT 373.650 821.400 375.450 827.250 ;
        RECT 376.650 821.400 378.450 827.250 ;
        RECT 379.650 821.400 381.450 827.250 ;
        RECT 391.650 821.400 393.450 827.250 ;
        RECT 394.650 821.400 396.450 827.250 ;
        RECT 397.650 821.400 399.450 827.250 ;
        RECT 400.650 821.400 402.450 827.250 ;
        RECT 403.650 821.400 405.450 827.250 ;
        RECT 348.150 819.600 353.250 820.500 ;
        RECT 351.000 818.700 353.250 819.600 ;
        RECT 333.450 814.050 337.050 816.150 ;
        RECT 274.200 804.300 291.900 805.350 ;
        RECT 269.700 802.500 273.750 803.400 ;
        RECT 272.700 801.600 273.750 802.500 ;
        RECT 269.700 795.750 271.500 801.600 ;
        RECT 272.700 795.750 274.500 801.600 ;
        RECT 275.700 795.750 277.500 801.600 ;
        RECT 278.700 795.750 280.500 804.300 ;
        RECT 298.950 804.150 301.050 804.600 ;
        RECT 298.650 802.500 301.050 804.150 ;
        RECT 303.000 802.800 306.900 804.600 ;
        RECT 303.000 802.500 306.000 802.800 ;
        RECT 283.950 799.950 286.050 802.050 ;
        RECT 286.950 799.950 289.050 802.050 ;
        RECT 289.950 801.600 292.050 802.050 ;
        RECT 298.650 801.600 300.000 802.500 ;
        RECT 289.950 799.950 292.500 801.600 ;
        RECT 281.700 795.750 283.500 799.050 ;
        RECT 284.850 798.600 286.050 799.950 ;
        RECT 288.150 798.600 289.050 799.950 ;
        RECT 291.300 798.600 292.500 799.950 ;
        RECT 284.850 795.750 287.250 798.600 ;
        RECT 288.150 795.750 290.250 798.600 ;
        RECT 291.300 795.750 293.250 798.600 ;
        RECT 294.450 795.750 296.250 801.600 ;
        RECT 298.200 795.750 300.000 801.600 ;
        RECT 301.200 795.750 303.000 801.600 ;
        RECT 304.200 795.750 306.000 802.500 ;
        RECT 308.100 798.600 309.450 805.650 ;
        RECT 317.850 804.150 319.650 804.300 ;
        RECT 310.950 802.950 319.650 804.150 ;
        RECT 324.600 803.700 326.400 804.300 ;
        RECT 310.950 802.050 313.050 802.950 ;
        RECT 317.850 802.500 319.650 802.950 ;
        RECT 320.700 802.500 326.400 803.700 ;
        RECT 307.950 795.750 309.750 798.600 ;
        RECT 310.950 795.750 312.750 802.050 ;
        RECT 314.100 799.800 316.200 801.900 ;
        RECT 314.100 798.600 315.600 799.800 ;
        RECT 313.950 795.750 315.750 798.600 ;
        RECT 317.700 795.750 319.500 801.600 ;
        RECT 320.700 795.750 322.500 802.500 ;
        RECT 327.300 801.600 328.500 805.650 ;
        RECT 333.450 801.600 334.950 814.050 ;
        RECT 346.950 812.850 349.050 814.950 ;
        RECT 347.100 811.050 348.900 812.850 ;
        RECT 351.000 810.300 352.050 818.700 ;
        RECT 354.150 814.950 355.350 821.400 ;
        RECT 371.250 820.500 372.450 821.400 ;
        RECT 377.250 820.500 378.450 821.400 ;
        RECT 394.800 820.500 396.600 821.400 ;
        RECT 400.800 820.500 402.600 821.400 ;
        RECT 406.650 820.500 408.450 827.250 ;
        RECT 409.650 821.400 411.450 827.250 ;
        RECT 412.650 821.400 414.450 827.250 ;
        RECT 415.650 821.400 417.450 827.250 ;
        RECT 422.550 824.400 424.350 827.250 ;
        RECT 425.550 824.400 427.350 827.250 ;
        RECT 412.800 820.500 414.600 821.400 ;
        RECT 371.250 819.300 378.450 820.500 ;
        RECT 393.900 820.350 396.600 820.500 ;
        RECT 393.750 819.300 396.600 820.350 ;
        RECT 398.700 819.300 402.600 820.500 ;
        RECT 404.700 819.300 408.450 820.500 ;
        RECT 410.550 819.300 414.600 820.500 ;
        RECT 371.250 814.950 372.450 819.300 ;
        RECT 393.750 816.150 394.800 819.300 ;
        RECT 398.700 818.400 399.900 819.300 ;
        RECT 404.700 818.400 405.900 819.300 ;
        RECT 410.550 818.400 411.750 819.300 ;
        RECT 395.700 816.600 399.900 818.400 ;
        RECT 401.700 816.600 405.900 818.400 ;
        RECT 407.700 816.600 411.750 818.400 ;
        RECT 352.950 812.850 355.350 814.950 ;
        RECT 370.950 812.850 373.050 814.950 ;
        RECT 376.950 812.850 379.050 814.950 ;
        RECT 391.950 814.050 394.800 816.150 ;
        RECT 351.000 809.400 353.250 810.300 ;
        RECT 347.550 808.500 353.250 809.400 ;
        RECT 347.550 801.600 348.750 808.500 ;
        RECT 354.150 807.600 355.350 812.850 ;
        RECT 371.250 809.400 372.450 812.850 ;
        RECT 377.100 811.050 378.900 812.850 ;
        RECT 393.750 809.700 394.800 814.050 ;
        RECT 398.700 809.700 399.900 816.600 ;
        RECT 404.700 809.700 405.900 816.600 ;
        RECT 410.550 809.700 411.750 816.600 ;
        RECT 413.100 816.150 414.900 817.950 ;
        RECT 412.950 814.050 415.050 816.150 ;
        RECT 421.950 815.850 424.050 817.950 ;
        RECT 425.400 816.150 426.600 824.400 ;
        RECT 434.850 821.400 436.650 827.250 ;
        RECT 439.350 820.200 441.150 827.250 ;
        RECT 450.000 821.400 451.800 827.250 ;
        RECT 454.200 823.050 456.000 827.250 ;
        RECT 457.500 824.400 459.300 827.250 ;
        RECT 470.700 824.400 472.500 827.250 ;
        RECT 474.000 823.050 475.800 827.250 ;
        RECT 454.200 821.400 459.900 823.050 ;
        RECT 437.550 819.300 441.150 820.200 ;
        RECT 422.100 814.050 423.900 815.850 ;
        RECT 424.950 814.050 427.050 816.150 ;
        RECT 371.250 808.500 378.450 809.400 ;
        RECT 393.750 808.500 396.450 809.700 ;
        RECT 398.700 808.500 402.450 809.700 ;
        RECT 404.700 808.500 408.450 809.700 ;
        RECT 410.550 808.500 414.450 809.700 ;
        RECT 371.250 807.600 372.450 808.500 ;
        RECT 323.700 795.750 325.500 801.600 ;
        RECT 326.700 795.750 328.500 801.600 ;
        RECT 329.700 795.750 331.500 801.600 ;
        RECT 333.450 795.750 335.250 801.600 ;
        RECT 336.450 795.750 338.250 801.600 ;
        RECT 347.550 795.750 349.350 801.600 ;
        RECT 350.850 795.750 352.650 807.600 ;
        RECT 353.850 795.750 355.650 807.600 ;
        RECT 367.650 795.750 369.450 807.600 ;
        RECT 370.650 795.750 372.450 807.600 ;
        RECT 373.650 795.750 375.450 807.600 ;
        RECT 376.650 795.750 378.450 808.500 ;
        RECT 379.650 795.750 381.450 807.600 ;
        RECT 391.650 795.750 393.450 807.600 ;
        RECT 394.650 795.750 396.450 808.500 ;
        RECT 397.650 795.750 399.450 807.600 ;
        RECT 400.650 795.750 402.450 808.500 ;
        RECT 403.650 795.750 405.450 807.600 ;
        RECT 406.650 795.750 408.450 808.500 ;
        RECT 409.650 795.750 411.450 807.600 ;
        RECT 412.650 795.750 414.450 808.500 ;
        RECT 415.650 795.750 417.450 807.600 ;
        RECT 425.400 801.600 426.600 814.050 ;
        RECT 434.100 813.150 435.900 814.950 ;
        RECT 433.950 811.050 436.050 813.150 ;
        RECT 437.550 811.950 438.750 819.300 ;
        RECT 449.100 816.150 450.900 817.950 ;
        RECT 440.100 813.150 441.900 814.950 ;
        RECT 448.950 814.050 451.050 816.150 ;
        RECT 451.950 815.850 454.050 817.950 ;
        RECT 455.100 816.150 456.900 817.950 ;
        RECT 452.100 814.050 453.900 815.850 ;
        RECT 454.950 814.050 457.050 816.150 ;
        RECT 458.700 814.950 459.900 821.400 ;
        RECT 470.100 821.400 475.800 823.050 ;
        RECT 478.200 821.400 480.000 827.250 ;
        RECT 470.100 814.950 471.300 821.400 ;
        RECT 488.850 820.200 490.650 827.250 ;
        RECT 493.350 821.400 495.150 827.250 ;
        RECT 504.150 822.900 505.950 827.250 ;
        RECT 502.650 821.400 505.950 822.900 ;
        RECT 507.150 821.400 508.950 827.250 ;
        RECT 488.850 819.300 492.450 820.200 ;
        RECT 473.100 816.150 474.900 817.950 ;
        RECT 436.950 809.850 439.050 811.950 ;
        RECT 439.950 811.050 442.050 813.150 ;
        RECT 457.950 812.850 460.050 814.950 ;
        RECT 469.950 812.850 472.050 814.950 ;
        RECT 472.950 814.050 475.050 816.150 ;
        RECT 475.950 815.850 478.050 817.950 ;
        RECT 479.100 816.150 480.900 817.950 ;
        RECT 476.100 814.050 477.900 815.850 ;
        RECT 478.950 814.050 481.050 816.150 ;
        RECT 488.100 813.150 489.900 814.950 ;
        RECT 437.550 801.600 438.750 809.850 ;
        RECT 458.700 807.600 459.900 812.850 ;
        RECT 470.100 807.600 471.300 812.850 ;
        RECT 487.950 811.050 490.050 813.150 ;
        RECT 491.250 811.950 492.450 819.300 ;
        RECT 502.650 814.950 503.850 821.400 ;
        RECT 505.950 819.900 507.750 820.500 ;
        RECT 511.650 819.900 513.450 827.250 ;
        RECT 517.650 826.500 525.450 827.250 ;
        RECT 517.650 821.400 519.450 826.500 ;
        RECT 520.650 821.400 522.450 825.600 ;
        RECT 523.650 822.000 525.450 826.500 ;
        RECT 526.650 822.900 528.450 827.250 ;
        RECT 529.650 822.000 531.450 827.250 ;
        RECT 505.950 818.700 513.450 819.900 ;
        RECT 521.250 819.900 522.150 821.400 ;
        RECT 523.650 821.100 531.450 822.000 ;
        RECT 538.650 821.400 540.450 827.250 ;
        RECT 521.250 818.850 525.600 819.900 ;
        RECT 494.100 813.150 495.900 814.950 ;
        RECT 490.950 809.850 493.050 811.950 ;
        RECT 493.950 811.050 496.050 813.150 ;
        RECT 502.650 812.850 505.050 814.950 ;
        RECT 506.100 813.150 507.900 814.950 ;
        RECT 449.550 806.700 457.350 807.600 ;
        RECT 422.550 795.750 424.350 801.600 ;
        RECT 425.550 795.750 427.350 801.600 ;
        RECT 434.550 795.750 436.350 801.600 ;
        RECT 437.550 795.750 439.350 801.600 ;
        RECT 440.550 795.750 442.350 801.600 ;
        RECT 449.550 795.750 451.350 806.700 ;
        RECT 452.550 795.750 454.350 805.800 ;
        RECT 455.550 795.750 457.350 806.700 ;
        RECT 458.550 795.750 460.350 807.600 ;
        RECT 469.650 795.750 471.450 807.600 ;
        RECT 472.650 806.700 480.450 807.600 ;
        RECT 472.650 795.750 474.450 806.700 ;
        RECT 475.650 795.750 477.450 805.800 ;
        RECT 478.650 795.750 480.450 806.700 ;
        RECT 491.250 801.600 492.450 809.850 ;
        RECT 502.650 807.600 503.850 812.850 ;
        RECT 505.950 811.050 508.050 813.150 ;
        RECT 487.650 795.750 489.450 801.600 ;
        RECT 490.650 795.750 492.450 801.600 ;
        RECT 493.650 795.750 495.450 801.600 ;
        RECT 502.050 795.750 503.850 807.600 ;
        RECT 505.050 795.750 506.850 807.600 ;
        RECT 509.100 801.600 510.300 818.700 ;
        RECT 521.700 816.150 523.500 817.950 ;
        RECT 511.950 812.850 514.050 814.950 ;
        RECT 517.950 812.850 520.050 814.950 ;
        RECT 520.950 814.050 523.050 816.150 ;
        RECT 524.400 814.950 525.600 818.850 ;
        RECT 539.250 819.300 540.450 821.400 ;
        RECT 541.650 822.300 543.450 827.250 ;
        RECT 544.650 823.200 546.450 827.250 ;
        RECT 547.650 822.300 549.450 827.250 ;
        RECT 541.650 820.950 549.450 822.300 ;
        RECT 554.550 822.300 556.350 827.250 ;
        RECT 557.550 823.200 559.350 827.250 ;
        RECT 560.550 822.300 562.350 827.250 ;
        RECT 554.550 820.950 562.350 822.300 ;
        RECT 563.550 821.400 565.350 827.250 ;
        RECT 574.650 824.400 576.450 827.250 ;
        RECT 577.650 824.400 579.450 827.250 ;
        RECT 563.550 819.300 564.750 821.400 ;
        RECT 539.250 818.250 543.000 819.300 ;
        RECT 561.000 818.250 564.750 819.300 ;
        RECT 527.100 816.150 528.900 817.950 ;
        RECT 523.950 812.850 526.050 814.950 ;
        RECT 526.950 814.050 529.050 816.150 ;
        RECT 541.950 814.950 543.150 818.250 ;
        RECT 545.100 816.150 546.900 817.950 ;
        RECT 557.100 816.150 558.900 817.950 ;
        RECT 529.950 812.850 532.050 814.950 ;
        RECT 541.950 812.850 544.050 814.950 ;
        RECT 544.950 814.050 547.050 816.150 ;
        RECT 547.950 812.850 550.050 814.950 ;
        RECT 553.950 812.850 556.050 814.950 ;
        RECT 556.950 814.050 559.050 816.150 ;
        RECT 560.850 814.950 562.050 818.250 ;
        RECT 575.400 816.150 576.600 824.400 ;
        RECT 584.850 820.200 586.650 827.250 ;
        RECT 589.350 821.400 591.150 827.250 ;
        RECT 596.550 824.400 598.350 827.250 ;
        RECT 599.550 824.400 601.350 827.250 ;
        RECT 584.850 819.300 588.450 820.200 ;
        RECT 559.950 812.850 562.050 814.950 ;
        RECT 574.950 814.050 577.050 816.150 ;
        RECT 577.950 815.850 580.050 817.950 ;
        RECT 578.100 814.050 579.900 815.850 ;
        RECT 512.100 811.050 513.900 812.850 ;
        RECT 518.250 811.050 520.050 812.850 ;
        RECT 524.250 807.600 525.450 812.850 ;
        RECT 530.100 811.050 531.900 812.850 ;
        RECT 538.950 809.850 541.050 811.950 ;
        RECT 539.250 808.050 541.050 809.850 ;
        RECT 542.850 807.600 544.050 812.850 ;
        RECT 548.100 811.050 549.900 812.850 ;
        RECT 554.100 811.050 555.900 812.850 ;
        RECT 559.950 807.600 561.150 812.850 ;
        RECT 562.950 809.850 565.050 811.950 ;
        RECT 562.950 808.050 564.750 809.850 ;
        RECT 508.650 795.750 510.450 801.600 ;
        RECT 511.650 795.750 513.450 801.600 ;
        RECT 519.150 795.750 520.950 807.600 ;
        RECT 523.650 795.750 526.950 807.600 ;
        RECT 529.650 795.750 531.450 807.600 ;
        RECT 539.400 795.750 541.200 801.600 ;
        RECT 542.700 795.750 544.500 807.600 ;
        RECT 546.900 795.750 548.700 807.600 ;
        RECT 555.300 795.750 557.100 807.600 ;
        RECT 559.500 795.750 561.300 807.600 ;
        RECT 575.400 801.600 576.600 814.050 ;
        RECT 584.100 813.150 585.900 814.950 ;
        RECT 583.950 811.050 586.050 813.150 ;
        RECT 587.250 811.950 588.450 819.300 ;
        RECT 595.950 815.850 598.050 817.950 ;
        RECT 599.400 816.150 600.600 824.400 ;
        RECT 610.650 821.400 612.450 827.250 ;
        RECT 611.250 819.300 612.450 821.400 ;
        RECT 613.650 822.300 615.450 827.250 ;
        RECT 616.650 823.200 618.450 827.250 ;
        RECT 619.650 822.300 621.450 827.250 ;
        RECT 613.650 820.950 621.450 822.300 ;
        RECT 611.250 818.250 615.000 819.300 ;
        RECT 632.100 819.000 633.900 827.250 ;
        RECT 590.100 813.150 591.900 814.950 ;
        RECT 596.100 814.050 597.900 815.850 ;
        RECT 598.950 814.050 601.050 816.150 ;
        RECT 613.950 814.950 615.150 818.250 ;
        RECT 617.100 816.150 618.900 817.950 ;
        RECT 629.400 817.350 633.900 819.000 ;
        RECT 637.500 818.400 639.300 827.250 ;
        RECT 641.550 821.400 643.350 827.250 ;
        RECT 644.550 821.400 646.350 827.250 ;
        RECT 586.950 809.850 589.050 811.950 ;
        RECT 589.950 811.050 592.050 813.150 ;
        RECT 587.250 801.600 588.450 809.850 ;
        RECT 599.400 801.600 600.600 814.050 ;
        RECT 613.950 812.850 616.050 814.950 ;
        RECT 616.950 814.050 619.050 816.150 ;
        RECT 619.950 812.850 622.050 814.950 ;
        RECT 629.400 813.150 630.600 817.350 ;
        RECT 641.100 816.150 642.900 817.950 ;
        RECT 640.950 814.050 643.050 816.150 ;
        RECT 644.400 814.950 645.600 821.400 ;
        RECT 656.850 820.200 658.650 827.250 ;
        RECT 661.350 821.400 663.150 827.250 ;
        RECT 656.850 819.300 660.450 820.200 ;
        RECT 610.950 809.850 613.050 811.950 ;
        RECT 611.250 808.050 613.050 809.850 ;
        RECT 614.850 807.600 616.050 812.850 ;
        RECT 620.100 811.050 621.900 812.850 ;
        RECT 628.950 811.050 631.050 813.150 ;
        RECT 643.950 812.850 646.050 814.950 ;
        RECT 656.100 813.150 657.900 814.950 ;
        RECT 562.800 795.750 564.600 801.600 ;
        RECT 574.650 795.750 576.450 801.600 ;
        RECT 577.650 795.750 579.450 801.600 ;
        RECT 583.650 795.750 585.450 801.600 ;
        RECT 586.650 795.750 588.450 801.600 ;
        RECT 589.650 795.750 591.450 801.600 ;
        RECT 596.550 795.750 598.350 801.600 ;
        RECT 599.550 795.750 601.350 801.600 ;
        RECT 611.400 795.750 613.200 801.600 ;
        RECT 614.700 795.750 616.500 807.600 ;
        RECT 618.900 795.750 620.700 807.600 ;
        RECT 629.250 802.800 630.300 811.050 ;
        RECT 631.950 809.850 634.050 811.950 ;
        RECT 637.950 809.850 640.050 811.950 ;
        RECT 631.950 808.050 633.750 809.850 ;
        RECT 634.950 806.850 637.050 808.950 ;
        RECT 638.100 808.050 639.900 809.850 ;
        RECT 644.400 807.600 645.600 812.850 ;
        RECT 655.950 811.050 658.050 813.150 ;
        RECT 659.250 811.950 660.450 819.300 ;
        RECT 674.100 819.000 675.900 827.250 ;
        RECT 671.400 817.350 675.900 819.000 ;
        RECT 679.500 818.400 681.300 827.250 ;
        RECT 689.850 820.200 691.650 827.250 ;
        RECT 694.350 821.400 696.150 827.250 ;
        RECT 701.850 821.400 703.650 827.250 ;
        RECT 706.350 820.200 708.150 827.250 ;
        RECT 716.850 821.400 718.650 827.250 ;
        RECT 721.350 820.200 723.150 827.250 ;
        RECT 735.150 822.900 736.950 827.250 ;
        RECT 689.850 819.300 693.450 820.200 ;
        RECT 662.100 813.150 663.900 814.950 ;
        RECT 671.400 813.150 672.600 817.350 ;
        RECT 689.100 813.150 690.900 814.950 ;
        RECT 658.950 809.850 661.050 811.950 ;
        RECT 661.950 811.050 664.050 813.150 ;
        RECT 670.950 811.050 673.050 813.150 ;
        RECT 635.100 805.050 636.900 806.850 ;
        RECT 629.250 801.900 636.300 802.800 ;
        RECT 629.250 801.600 630.450 801.900 ;
        RECT 628.650 795.750 630.450 801.600 ;
        RECT 634.650 801.600 636.300 801.900 ;
        RECT 631.650 795.750 633.450 801.000 ;
        RECT 634.650 795.750 636.450 801.600 ;
        RECT 637.650 795.750 639.450 801.600 ;
        RECT 641.550 795.750 643.350 807.600 ;
        RECT 644.550 795.750 646.350 807.600 ;
        RECT 659.250 801.600 660.450 809.850 ;
        RECT 671.250 802.800 672.300 811.050 ;
        RECT 673.950 809.850 676.050 811.950 ;
        RECT 679.950 809.850 682.050 811.950 ;
        RECT 688.950 811.050 691.050 813.150 ;
        RECT 692.250 811.950 693.450 819.300 ;
        RECT 704.550 819.300 708.150 820.200 ;
        RECT 719.550 819.300 723.150 820.200 ;
        RECT 733.650 821.400 736.950 822.900 ;
        RECT 738.150 821.400 739.950 827.250 ;
        RECT 695.100 813.150 696.900 814.950 ;
        RECT 701.100 813.150 702.900 814.950 ;
        RECT 691.950 809.850 694.050 811.950 ;
        RECT 694.950 811.050 697.050 813.150 ;
        RECT 700.950 811.050 703.050 813.150 ;
        RECT 704.550 811.950 705.750 819.300 ;
        RECT 707.100 813.150 708.900 814.950 ;
        RECT 716.100 813.150 717.900 814.950 ;
        RECT 703.950 809.850 706.050 811.950 ;
        RECT 706.950 811.050 709.050 813.150 ;
        RECT 715.950 811.050 718.050 813.150 ;
        RECT 719.550 811.950 720.750 819.300 ;
        RECT 733.650 814.950 734.850 821.400 ;
        RECT 736.950 819.900 738.750 820.500 ;
        RECT 742.650 819.900 744.450 827.250 ;
        RECT 751.650 824.400 753.450 827.250 ;
        RECT 754.650 824.400 756.450 827.250 ;
        RECT 736.950 818.700 744.450 819.900 ;
        RECT 722.100 813.150 723.900 814.950 ;
        RECT 718.950 809.850 721.050 811.950 ;
        RECT 721.950 811.050 724.050 813.150 ;
        RECT 733.650 812.850 736.050 814.950 ;
        RECT 737.100 813.150 738.900 814.950 ;
        RECT 673.950 808.050 675.750 809.850 ;
        RECT 676.950 806.850 679.050 808.950 ;
        RECT 680.100 808.050 681.900 809.850 ;
        RECT 677.100 805.050 678.900 806.850 ;
        RECT 671.250 801.900 678.300 802.800 ;
        RECT 671.250 801.600 672.450 801.900 ;
        RECT 655.650 795.750 657.450 801.600 ;
        RECT 658.650 795.750 660.450 801.600 ;
        RECT 661.650 795.750 663.450 801.600 ;
        RECT 670.650 795.750 672.450 801.600 ;
        RECT 676.650 801.600 678.300 801.900 ;
        RECT 692.250 801.600 693.450 809.850 ;
        RECT 704.550 801.600 705.750 809.850 ;
        RECT 719.550 801.600 720.750 809.850 ;
        RECT 733.650 807.600 734.850 812.850 ;
        RECT 736.950 811.050 739.050 813.150 ;
        RECT 673.650 795.750 675.450 801.000 ;
        RECT 676.650 795.750 678.450 801.600 ;
        RECT 679.650 795.750 681.450 801.600 ;
        RECT 688.650 795.750 690.450 801.600 ;
        RECT 691.650 795.750 693.450 801.600 ;
        RECT 694.650 795.750 696.450 801.600 ;
        RECT 701.550 795.750 703.350 801.600 ;
        RECT 704.550 795.750 706.350 801.600 ;
        RECT 707.550 795.750 709.350 801.600 ;
        RECT 716.550 795.750 718.350 801.600 ;
        RECT 719.550 795.750 721.350 801.600 ;
        RECT 722.550 795.750 724.350 801.600 ;
        RECT 733.050 795.750 734.850 807.600 ;
        RECT 736.050 795.750 737.850 807.600 ;
        RECT 740.100 801.600 741.300 818.700 ;
        RECT 752.400 816.150 753.600 824.400 ;
        RECT 767.850 820.200 769.650 827.250 ;
        RECT 772.350 821.400 774.150 827.250 ;
        RECT 767.850 819.300 771.450 820.200 ;
        RECT 742.950 812.850 745.050 814.950 ;
        RECT 751.950 814.050 754.050 816.150 ;
        RECT 754.950 815.850 757.050 817.950 ;
        RECT 755.100 814.050 756.900 815.850 ;
        RECT 743.100 811.050 744.900 812.850 ;
        RECT 752.400 801.600 753.600 814.050 ;
        RECT 767.100 813.150 768.900 814.950 ;
        RECT 766.950 811.050 769.050 813.150 ;
        RECT 770.250 811.950 771.450 819.300 ;
        RECT 776.700 818.400 778.500 827.250 ;
        RECT 782.100 819.000 783.900 827.250 ;
        RECT 793.650 821.400 795.450 827.250 ;
        RECT 782.100 817.350 786.600 819.000 ;
        RECT 787.950 817.950 790.050 820.050 ;
        RECT 794.250 819.300 795.450 821.400 ;
        RECT 796.650 822.300 798.450 827.250 ;
        RECT 799.650 823.200 801.450 827.250 ;
        RECT 802.650 822.300 804.450 827.250 ;
        RECT 812.550 824.400 814.350 827.250 ;
        RECT 815.550 824.400 817.350 827.250 ;
        RECT 826.650 824.400 828.450 827.250 ;
        RECT 829.650 824.400 831.450 827.250 ;
        RECT 796.650 820.950 804.450 822.300 ;
        RECT 794.250 818.250 798.000 819.300 ;
        RECT 773.100 813.150 774.900 814.950 ;
        RECT 785.400 813.150 786.600 817.350 ;
        RECT 769.950 809.850 772.050 811.950 ;
        RECT 772.950 811.050 775.050 813.150 ;
        RECT 775.950 809.850 778.050 811.950 ;
        RECT 781.950 809.850 784.050 811.950 ;
        RECT 784.950 811.050 787.050 813.150 ;
        RECT 770.250 801.600 771.450 809.850 ;
        RECT 776.100 808.050 777.900 809.850 ;
        RECT 778.950 806.850 781.050 808.950 ;
        RECT 782.250 808.050 784.050 809.850 ;
        RECT 779.100 805.050 780.900 806.850 ;
        RECT 785.700 802.800 786.750 811.050 ;
        RECT 788.550 807.450 789.450 817.950 ;
        RECT 796.950 814.950 798.150 818.250 ;
        RECT 800.100 816.150 801.900 817.950 ;
        RECT 796.950 812.850 799.050 814.950 ;
        RECT 799.950 814.050 802.050 816.150 ;
        RECT 811.950 815.850 814.050 817.950 ;
        RECT 815.400 816.150 816.600 824.400 ;
        RECT 827.400 816.150 828.600 824.400 ;
        RECT 836.850 821.400 838.650 827.250 ;
        RECT 841.350 820.200 843.150 827.250 ;
        RECT 839.550 819.300 843.150 820.200 ;
        RECT 802.950 812.850 805.050 814.950 ;
        RECT 812.100 814.050 813.900 815.850 ;
        RECT 814.950 814.050 817.050 816.150 ;
        RECT 826.950 814.050 829.050 816.150 ;
        RECT 829.950 815.850 832.050 817.950 ;
        RECT 830.100 814.050 831.900 815.850 ;
        RECT 793.950 809.850 796.050 811.950 ;
        RECT 794.250 808.050 796.050 809.850 ;
        RECT 797.850 807.600 799.050 812.850 ;
        RECT 803.100 811.050 804.900 812.850 ;
        RECT 788.550 806.550 792.450 807.450 ;
        RECT 791.550 804.450 792.450 806.550 ;
        RECT 793.950 804.450 796.050 805.050 ;
        RECT 791.550 803.550 796.050 804.450 ;
        RECT 793.950 802.950 796.050 803.550 ;
        RECT 779.700 801.900 786.750 802.800 ;
        RECT 779.700 801.600 781.350 801.900 ;
        RECT 739.650 795.750 741.450 801.600 ;
        RECT 742.650 795.750 744.450 801.600 ;
        RECT 751.650 795.750 753.450 801.600 ;
        RECT 754.650 795.750 756.450 801.600 ;
        RECT 766.650 795.750 768.450 801.600 ;
        RECT 769.650 795.750 771.450 801.600 ;
        RECT 772.650 795.750 774.450 801.600 ;
        RECT 776.550 795.750 778.350 801.600 ;
        RECT 779.550 795.750 781.350 801.600 ;
        RECT 785.550 801.600 786.750 801.900 ;
        RECT 782.550 795.750 784.350 801.000 ;
        RECT 785.550 795.750 787.350 801.600 ;
        RECT 794.400 795.750 796.200 801.600 ;
        RECT 797.700 795.750 799.500 807.600 ;
        RECT 801.900 795.750 803.700 807.600 ;
        RECT 815.400 801.600 816.600 814.050 ;
        RECT 827.400 801.600 828.600 814.050 ;
        RECT 836.100 813.150 837.900 814.950 ;
        RECT 835.950 811.050 838.050 813.150 ;
        RECT 839.550 811.950 840.750 819.300 ;
        RECT 842.100 813.150 843.900 814.950 ;
        RECT 838.950 809.850 841.050 811.950 ;
        RECT 841.950 811.050 844.050 813.150 ;
        RECT 839.550 801.600 840.750 809.850 ;
        RECT 812.550 795.750 814.350 801.600 ;
        RECT 815.550 795.750 817.350 801.600 ;
        RECT 826.650 795.750 828.450 801.600 ;
        RECT 829.650 795.750 831.450 801.600 ;
        RECT 836.550 795.750 838.350 801.600 ;
        RECT 839.550 795.750 841.350 801.600 ;
        RECT 842.550 795.750 844.350 801.600 ;
        RECT 7.650 785.400 9.450 791.250 ;
        RECT 10.650 785.400 12.450 791.250 ;
        RECT 13.650 785.400 15.450 791.250 ;
        RECT 11.250 777.150 12.450 785.400 ;
        RECT 20.550 779.400 22.350 791.250 ;
        RECT 25.050 779.550 26.850 791.250 ;
        RECT 28.050 780.900 29.850 791.250 ;
        RECT 40.650 785.400 42.450 791.250 ;
        RECT 43.650 785.400 45.450 791.250 ;
        RECT 46.650 785.400 48.450 791.250 ;
        RECT 28.050 779.550 30.450 780.900 ;
        RECT 20.550 778.200 21.750 779.400 ;
        RECT 25.950 778.200 27.750 778.650 ;
        RECT 7.950 773.850 10.050 775.950 ;
        RECT 10.950 775.050 13.050 777.150 ;
        RECT 20.550 777.000 27.750 778.200 ;
        RECT 25.950 776.850 27.750 777.000 ;
        RECT 8.100 772.050 9.900 773.850 ;
        RECT 11.250 767.700 12.450 775.050 ;
        RECT 13.950 773.850 16.050 775.950 ;
        RECT 23.100 774.150 24.900 775.950 ;
        RECT 14.100 772.050 15.900 773.850 ;
        RECT 20.100 771.150 21.900 772.950 ;
        RECT 22.950 772.050 25.050 774.150 ;
        RECT 19.950 769.050 22.050 771.150 ;
        RECT 26.700 768.600 27.600 776.850 ;
        RECT 29.100 772.950 30.450 779.550 ;
        RECT 44.250 777.150 45.450 785.400 ;
        RECT 53.550 779.400 55.350 791.250 ;
        RECT 57.750 779.400 59.550 791.250 ;
        RECT 65.700 785.400 67.500 791.250 ;
        RECT 68.700 785.400 70.500 791.250 ;
        RECT 71.700 785.400 73.500 791.250 ;
        RECT 68.700 784.500 69.750 785.400 ;
        RECT 57.000 778.350 59.550 779.400 ;
        RECT 65.700 783.600 69.750 784.500 ;
        RECT 40.950 773.850 43.050 775.950 ;
        RECT 43.950 775.050 46.050 777.150 ;
        RECT 28.950 770.850 31.050 772.950 ;
        RECT 41.100 772.050 42.900 773.850 ;
        RECT 25.950 767.700 27.750 768.600 ;
        RECT 8.850 766.800 12.450 767.700 ;
        RECT 24.450 766.800 27.750 767.700 ;
        RECT 8.850 759.750 10.650 766.800 ;
        RECT 13.350 759.750 15.150 765.600 ;
        RECT 24.450 762.600 25.350 766.800 ;
        RECT 30.000 765.600 31.050 770.850 ;
        RECT 44.250 767.700 45.450 775.050 ;
        RECT 46.950 773.850 49.050 775.950 ;
        RECT 53.100 774.150 54.900 775.950 ;
        RECT 47.100 772.050 48.900 773.850 ;
        RECT 52.950 772.050 55.050 774.150 ;
        RECT 57.000 771.150 58.050 778.350 ;
        RECT 59.100 774.150 60.900 775.950 ;
        RECT 58.950 772.050 61.050 774.150 ;
        RECT 55.950 769.050 58.050 771.150 ;
        RECT 41.850 766.800 45.450 767.700 ;
        RECT 20.550 759.750 22.350 762.600 ;
        RECT 23.550 759.750 25.350 762.600 ;
        RECT 26.550 759.750 28.350 762.600 ;
        RECT 29.550 759.750 31.350 765.600 ;
        RECT 41.850 759.750 43.650 766.800 ;
        RECT 46.350 759.750 48.150 765.600 ;
        RECT 57.000 762.600 58.050 769.050 ;
        RECT 65.700 770.100 66.900 783.600 ;
        RECT 74.700 782.700 76.500 791.250 ;
        RECT 77.700 787.950 79.500 791.250 ;
        RECT 80.850 788.400 83.250 791.250 ;
        RECT 84.150 788.400 86.250 791.250 ;
        RECT 87.300 788.400 89.250 791.250 ;
        RECT 80.850 787.050 82.050 788.400 ;
        RECT 84.150 787.050 85.050 788.400 ;
        RECT 87.300 787.050 88.500 788.400 ;
        RECT 79.950 784.950 82.050 787.050 ;
        RECT 82.950 784.950 85.050 787.050 ;
        RECT 85.950 785.400 88.500 787.050 ;
        RECT 90.450 785.400 92.250 791.250 ;
        RECT 94.200 785.400 96.000 791.250 ;
        RECT 97.200 785.400 99.000 791.250 ;
        RECT 85.950 784.950 88.050 785.400 ;
        RECT 94.650 784.500 96.000 785.400 ;
        RECT 100.200 784.500 102.000 791.250 ;
        RECT 103.950 788.400 105.750 791.250 ;
        RECT 94.650 782.850 97.050 784.500 ;
        RECT 70.200 781.650 87.900 782.700 ;
        RECT 94.950 782.400 97.050 782.850 ;
        RECT 99.000 784.200 102.000 784.500 ;
        RECT 99.000 782.400 102.900 784.200 ;
        RECT 70.200 780.900 72.000 781.650 ;
        RECT 82.950 780.150 85.050 780.750 ;
        RECT 73.500 778.950 85.050 780.150 ;
        RECT 85.950 780.600 87.900 781.650 ;
        RECT 104.100 781.350 105.450 788.400 ;
        RECT 106.950 784.950 108.750 791.250 ;
        RECT 109.950 788.400 111.750 791.250 ;
        RECT 110.100 787.200 111.600 788.400 ;
        RECT 110.100 785.100 112.200 787.200 ;
        RECT 113.700 785.400 115.500 791.250 ;
        RECT 106.950 784.050 109.050 784.950 ;
        RECT 116.700 784.500 118.500 791.250 ;
        RECT 119.700 785.400 121.500 791.250 ;
        RECT 122.700 785.400 124.500 791.250 ;
        RECT 125.700 785.400 127.500 791.250 ;
        RECT 129.450 785.400 131.250 791.250 ;
        RECT 132.450 785.400 134.250 791.250 ;
        RECT 143.550 785.400 145.350 791.250 ;
        RECT 146.550 785.400 148.350 791.250 ;
        RECT 152.550 785.400 154.350 791.250 ;
        RECT 155.550 785.400 157.350 791.250 ;
        RECT 158.550 786.000 160.350 791.250 ;
        RECT 113.850 784.050 115.650 784.500 ;
        RECT 106.950 782.850 115.650 784.050 ;
        RECT 116.700 783.300 122.400 784.500 ;
        RECT 113.850 782.700 115.650 782.850 ;
        RECT 120.600 782.700 122.400 783.300 ;
        RECT 123.300 781.350 124.500 785.400 ;
        RECT 103.950 780.600 106.050 781.350 ;
        RECT 85.950 779.250 106.050 780.600 ;
        RECT 109.950 780.450 127.350 781.350 ;
        RECT 109.950 779.250 112.050 780.450 ;
        RECT 73.500 778.350 75.300 778.950 ;
        RECT 82.950 778.650 85.050 778.950 ;
        RECT 112.950 778.350 125.250 779.550 ;
        RECT 85.950 777.450 114.000 778.350 ;
        RECT 123.450 777.750 125.250 778.350 ;
        RECT 74.250 777.150 114.000 777.450 ;
        RECT 73.950 776.550 87.900 777.150 ;
        RECT 67.950 773.850 70.050 775.950 ;
        RECT 73.950 775.350 77.850 776.550 ;
        RECT 94.950 775.650 109.500 776.250 ;
        RECT 73.950 775.050 76.050 775.350 ;
        RECT 78.750 774.450 85.500 775.350 ;
        RECT 68.100 772.050 69.900 773.850 ;
        RECT 78.750 772.050 79.950 774.450 ;
        RECT 68.100 771.000 79.950 772.050 ;
        RECT 81.750 771.750 83.550 773.550 ;
        RECT 84.450 772.950 85.500 774.450 ;
        RECT 86.400 775.050 109.500 775.650 ;
        RECT 86.400 774.450 97.050 775.050 ;
        RECT 86.400 773.850 88.200 774.450 ;
        RECT 94.950 774.150 97.050 774.450 ;
        RECT 99.150 773.250 101.250 773.550 ;
        RECT 107.700 773.250 109.500 775.050 ;
        RECT 110.850 774.000 117.900 775.800 ;
        RECT 84.450 772.050 96.450 772.950 ;
        RECT 65.700 769.200 81.000 770.100 ;
        RECT 65.700 765.600 66.900 769.200 ;
        RECT 69.900 767.700 71.700 768.300 ;
        RECT 69.900 766.500 78.300 767.700 ;
        RECT 76.800 765.600 78.300 766.500 ;
        RECT 53.550 759.750 55.350 762.600 ;
        RECT 56.550 759.750 58.350 762.600 ;
        RECT 59.550 759.750 61.350 762.600 ;
        RECT 65.700 759.750 67.500 765.600 ;
        RECT 71.100 759.750 72.900 765.600 ;
        RECT 76.500 759.750 78.300 765.600 ;
        RECT 79.950 766.050 81.000 769.200 ;
        RECT 82.500 768.300 83.550 771.750 ;
        RECT 90.150 769.350 94.050 771.150 ;
        RECT 91.950 769.050 94.050 769.350 ;
        RECT 95.400 770.550 96.450 772.050 ;
        RECT 97.350 771.450 101.250 773.250 ;
        RECT 110.850 772.350 111.750 774.000 ;
        RECT 118.950 773.100 121.050 777.150 ;
        RECT 102.150 771.300 111.750 772.350 ;
        RECT 112.800 772.050 121.050 773.100 ;
        RECT 102.150 770.550 103.050 771.300 ;
        RECT 95.400 769.200 103.050 770.550 ;
        RECT 112.800 770.250 113.850 772.050 ;
        RECT 103.950 769.200 113.850 770.250 ;
        RECT 117.300 769.200 125.100 771.000 ;
        RECT 85.050 768.300 86.850 768.750 ;
        RECT 103.950 768.300 105.000 769.200 ;
        RECT 82.500 767.850 86.850 768.300 ;
        RECT 82.500 767.100 90.150 767.850 ;
        RECT 85.050 766.950 90.150 767.100 ;
        RECT 79.950 763.950 82.050 766.050 ;
        RECT 82.950 763.950 85.050 766.050 ;
        RECT 85.950 763.950 88.050 766.050 ;
        RECT 89.250 765.600 90.150 766.950 ;
        RECT 98.100 766.500 105.000 768.300 ;
        RECT 105.900 766.500 112.650 768.300 ;
        RECT 117.300 765.600 118.800 769.200 ;
        RECT 126.150 765.600 127.350 780.450 ;
        RECT 89.250 764.250 93.300 765.600 ;
        RECT 94.950 765.300 97.050 765.600 ;
        RECT 80.700 762.600 82.050 763.950 ;
        RECT 83.700 762.600 85.050 763.950 ;
        RECT 86.700 762.600 88.050 763.950 ;
        RECT 91.500 763.800 93.300 764.250 ;
        RECT 94.200 763.500 97.050 765.300 ;
        RECT 99.150 765.300 101.250 765.600 ;
        RECT 99.150 763.500 102.000 765.300 ;
        RECT 80.700 759.750 82.500 762.600 ;
        RECT 83.700 759.750 85.500 762.600 ;
        RECT 86.700 759.750 88.500 762.600 ;
        RECT 89.700 759.750 91.500 762.600 ;
        RECT 94.200 759.750 96.000 763.500 ;
        RECT 97.200 759.750 99.000 762.600 ;
        RECT 100.200 759.750 102.000 763.500 ;
        RECT 103.950 763.500 106.050 765.600 ;
        RECT 106.950 763.500 109.050 765.600 ;
        RECT 109.950 763.500 112.050 765.600 ;
        RECT 114.600 764.400 118.800 765.600 ;
        RECT 103.950 759.750 105.750 763.500 ;
        RECT 106.950 759.750 108.750 763.500 ;
        RECT 109.950 759.750 111.750 763.500 ;
        RECT 114.600 759.750 116.400 764.400 ;
        RECT 120.150 759.750 121.950 765.600 ;
        RECT 125.550 759.750 127.350 765.600 ;
        RECT 129.450 772.950 130.950 785.400 ;
        RECT 146.400 772.950 147.600 785.400 ;
        RECT 155.700 785.100 157.350 785.400 ;
        RECT 161.550 785.400 163.350 791.250 ;
        RECT 169.650 785.400 171.450 791.250 ;
        RECT 172.650 785.400 174.450 791.250 ;
        RECT 175.650 785.400 177.450 791.250 ;
        RECT 161.550 785.100 162.750 785.400 ;
        RECT 155.700 784.200 162.750 785.100 ;
        RECT 155.100 780.150 156.900 781.950 ;
        RECT 152.100 777.150 153.900 778.950 ;
        RECT 154.950 778.050 157.050 780.150 ;
        RECT 158.250 777.150 160.050 778.950 ;
        RECT 151.950 775.050 154.050 777.150 ;
        RECT 157.950 775.050 160.050 777.150 ;
        RECT 161.700 775.950 162.750 784.200 ;
        RECT 173.250 777.150 174.450 785.400 ;
        RECT 186.300 779.400 188.100 791.250 ;
        RECT 190.500 779.400 192.300 791.250 ;
        RECT 193.800 785.400 195.600 791.250 ;
        RECT 200.550 779.400 202.350 791.250 ;
        RECT 204.750 779.400 206.550 791.250 ;
        RECT 212.700 785.400 214.500 791.250 ;
        RECT 215.700 785.400 217.500 791.250 ;
        RECT 218.700 785.400 220.500 791.250 ;
        RECT 215.700 784.500 216.750 785.400 ;
        RECT 160.950 773.850 163.050 775.950 ;
        RECT 169.950 773.850 172.050 775.950 ;
        RECT 172.950 775.050 175.050 777.150 ;
        RECT 129.450 770.850 133.050 772.950 ;
        RECT 143.100 771.150 144.900 772.950 ;
        RECT 129.450 762.600 130.950 770.850 ;
        RECT 142.950 769.050 145.050 771.150 ;
        RECT 145.950 770.850 148.050 772.950 ;
        RECT 146.400 762.600 147.600 770.850 ;
        RECT 161.400 769.650 162.600 773.850 ;
        RECT 170.100 772.050 171.900 773.850 ;
        RECT 129.450 759.750 131.250 762.600 ;
        RECT 132.450 759.750 134.250 762.600 ;
        RECT 143.550 759.750 145.350 762.600 ;
        RECT 146.550 759.750 148.350 762.600 ;
        RECT 152.700 759.750 154.500 768.600 ;
        RECT 158.100 768.000 162.600 769.650 ;
        RECT 158.100 759.750 159.900 768.000 ;
        RECT 173.250 767.700 174.450 775.050 ;
        RECT 175.950 773.850 178.050 775.950 ;
        RECT 185.100 774.150 186.900 775.950 ;
        RECT 190.950 774.150 192.150 779.400 ;
        RECT 193.950 777.150 195.750 778.950 ;
        RECT 204.000 778.350 206.550 779.400 ;
        RECT 212.700 783.600 216.750 784.500 ;
        RECT 193.950 775.050 196.050 777.150 ;
        RECT 200.100 774.150 201.900 775.950 ;
        RECT 176.100 772.050 177.900 773.850 ;
        RECT 184.950 772.050 187.050 774.150 ;
        RECT 187.950 770.850 190.050 772.950 ;
        RECT 190.950 772.050 193.050 774.150 ;
        RECT 199.950 772.050 202.050 774.150 ;
        RECT 188.100 769.050 189.900 770.850 ;
        RECT 191.850 768.750 193.050 772.050 ;
        RECT 204.000 771.150 205.050 778.350 ;
        RECT 206.100 774.150 207.900 775.950 ;
        RECT 205.950 772.050 208.050 774.150 ;
        RECT 202.950 769.050 205.050 771.150 ;
        RECT 192.000 767.700 195.750 768.750 ;
        RECT 170.850 766.800 174.450 767.700 ;
        RECT 170.850 759.750 172.650 766.800 ;
        RECT 175.350 759.750 177.150 765.600 ;
        RECT 185.550 764.700 193.350 766.050 ;
        RECT 185.550 759.750 187.350 764.700 ;
        RECT 188.550 759.750 190.350 763.800 ;
        RECT 191.550 759.750 193.350 764.700 ;
        RECT 194.550 765.600 195.750 767.700 ;
        RECT 194.550 759.750 196.350 765.600 ;
        RECT 204.000 762.600 205.050 769.050 ;
        RECT 212.700 770.100 213.900 783.600 ;
        RECT 221.700 782.700 223.500 791.250 ;
        RECT 224.700 787.950 226.500 791.250 ;
        RECT 227.850 788.400 230.250 791.250 ;
        RECT 231.150 788.400 233.250 791.250 ;
        RECT 234.300 788.400 236.250 791.250 ;
        RECT 227.850 787.050 229.050 788.400 ;
        RECT 231.150 787.050 232.050 788.400 ;
        RECT 234.300 787.050 235.500 788.400 ;
        RECT 226.950 784.950 229.050 787.050 ;
        RECT 229.950 784.950 232.050 787.050 ;
        RECT 232.950 785.400 235.500 787.050 ;
        RECT 237.450 785.400 239.250 791.250 ;
        RECT 241.200 785.400 243.000 791.250 ;
        RECT 244.200 785.400 246.000 791.250 ;
        RECT 232.950 784.950 235.050 785.400 ;
        RECT 241.650 784.500 243.000 785.400 ;
        RECT 247.200 784.500 249.000 791.250 ;
        RECT 250.950 788.400 252.750 791.250 ;
        RECT 241.650 782.850 244.050 784.500 ;
        RECT 217.200 781.650 234.900 782.700 ;
        RECT 241.950 782.400 244.050 782.850 ;
        RECT 246.000 784.200 249.000 784.500 ;
        RECT 246.000 782.400 249.900 784.200 ;
        RECT 217.200 780.900 219.000 781.650 ;
        RECT 229.950 780.150 232.050 780.750 ;
        RECT 220.500 778.950 232.050 780.150 ;
        RECT 232.950 780.600 234.900 781.650 ;
        RECT 251.100 781.350 252.450 788.400 ;
        RECT 253.950 784.950 255.750 791.250 ;
        RECT 256.950 788.400 258.750 791.250 ;
        RECT 257.100 787.200 258.600 788.400 ;
        RECT 257.100 785.100 259.200 787.200 ;
        RECT 260.700 785.400 262.500 791.250 ;
        RECT 253.950 784.050 256.050 784.950 ;
        RECT 263.700 784.500 265.500 791.250 ;
        RECT 266.700 785.400 268.500 791.250 ;
        RECT 269.700 785.400 271.500 791.250 ;
        RECT 272.700 785.400 274.500 791.250 ;
        RECT 276.450 785.400 278.250 791.250 ;
        RECT 279.450 785.400 281.250 791.250 ;
        RECT 285.750 785.400 287.550 791.250 ;
        RECT 288.750 785.400 290.550 791.250 ;
        RECT 292.500 785.400 294.300 791.250 ;
        RECT 295.500 785.400 297.300 791.250 ;
        RECT 298.500 785.400 300.300 791.250 ;
        RECT 260.850 784.050 262.650 784.500 ;
        RECT 253.950 782.850 262.650 784.050 ;
        RECT 263.700 783.300 269.400 784.500 ;
        RECT 260.850 782.700 262.650 782.850 ;
        RECT 267.600 782.700 269.400 783.300 ;
        RECT 270.300 781.350 271.500 785.400 ;
        RECT 250.950 780.600 253.050 781.350 ;
        RECT 232.950 779.250 253.050 780.600 ;
        RECT 256.950 780.450 274.350 781.350 ;
        RECT 256.950 779.250 259.050 780.450 ;
        RECT 220.500 778.350 222.300 778.950 ;
        RECT 229.950 778.650 232.050 778.950 ;
        RECT 259.950 778.350 272.250 779.550 ;
        RECT 232.950 777.450 261.000 778.350 ;
        RECT 270.450 777.750 272.250 778.350 ;
        RECT 221.250 777.150 261.000 777.450 ;
        RECT 220.950 776.550 234.900 777.150 ;
        RECT 214.950 773.850 217.050 775.950 ;
        RECT 220.950 775.350 224.850 776.550 ;
        RECT 241.950 775.650 256.500 776.250 ;
        RECT 220.950 775.050 223.050 775.350 ;
        RECT 225.750 774.450 232.500 775.350 ;
        RECT 215.100 772.050 216.900 773.850 ;
        RECT 225.750 772.050 226.950 774.450 ;
        RECT 215.100 771.000 226.950 772.050 ;
        RECT 228.750 771.750 230.550 773.550 ;
        RECT 231.450 772.950 232.500 774.450 ;
        RECT 233.400 775.050 256.500 775.650 ;
        RECT 233.400 774.450 244.050 775.050 ;
        RECT 233.400 773.850 235.200 774.450 ;
        RECT 241.950 774.150 244.050 774.450 ;
        RECT 246.150 773.250 248.250 773.550 ;
        RECT 254.700 773.250 256.500 775.050 ;
        RECT 257.850 774.000 264.900 775.800 ;
        RECT 231.450 772.050 243.450 772.950 ;
        RECT 212.700 769.200 228.000 770.100 ;
        RECT 212.700 765.600 213.900 769.200 ;
        RECT 216.900 767.700 218.700 768.300 ;
        RECT 216.900 766.500 225.300 767.700 ;
        RECT 223.800 765.600 225.300 766.500 ;
        RECT 200.550 759.750 202.350 762.600 ;
        RECT 203.550 759.750 205.350 762.600 ;
        RECT 206.550 759.750 208.350 762.600 ;
        RECT 212.700 759.750 214.500 765.600 ;
        RECT 218.100 759.750 219.900 765.600 ;
        RECT 223.500 759.750 225.300 765.600 ;
        RECT 226.950 766.050 228.000 769.200 ;
        RECT 229.500 768.300 230.550 771.750 ;
        RECT 237.150 769.350 241.050 771.150 ;
        RECT 238.950 769.050 241.050 769.350 ;
        RECT 242.400 770.550 243.450 772.050 ;
        RECT 244.350 771.450 248.250 773.250 ;
        RECT 257.850 772.350 258.750 774.000 ;
        RECT 265.950 773.100 268.050 777.150 ;
        RECT 249.150 771.300 258.750 772.350 ;
        RECT 259.800 772.050 268.050 773.100 ;
        RECT 249.150 770.550 250.050 771.300 ;
        RECT 242.400 769.200 250.050 770.550 ;
        RECT 259.800 770.250 260.850 772.050 ;
        RECT 250.950 769.200 260.850 770.250 ;
        RECT 264.300 769.200 272.100 771.000 ;
        RECT 232.050 768.300 233.850 768.750 ;
        RECT 250.950 768.300 252.000 769.200 ;
        RECT 229.500 767.850 233.850 768.300 ;
        RECT 229.500 767.100 237.150 767.850 ;
        RECT 232.050 766.950 237.150 767.100 ;
        RECT 226.950 763.950 229.050 766.050 ;
        RECT 229.950 763.950 232.050 766.050 ;
        RECT 232.950 763.950 235.050 766.050 ;
        RECT 236.250 765.600 237.150 766.950 ;
        RECT 245.100 766.500 252.000 768.300 ;
        RECT 252.900 766.500 259.650 768.300 ;
        RECT 264.300 765.600 265.800 769.200 ;
        RECT 273.150 765.600 274.350 780.450 ;
        RECT 236.250 764.250 240.300 765.600 ;
        RECT 241.950 765.300 244.050 765.600 ;
        RECT 227.700 762.600 229.050 763.950 ;
        RECT 230.700 762.600 232.050 763.950 ;
        RECT 233.700 762.600 235.050 763.950 ;
        RECT 238.500 763.800 240.300 764.250 ;
        RECT 241.200 763.500 244.050 765.300 ;
        RECT 246.150 765.300 248.250 765.600 ;
        RECT 246.150 763.500 249.000 765.300 ;
        RECT 227.700 759.750 229.500 762.600 ;
        RECT 230.700 759.750 232.500 762.600 ;
        RECT 233.700 759.750 235.500 762.600 ;
        RECT 236.700 759.750 238.500 762.600 ;
        RECT 241.200 759.750 243.000 763.500 ;
        RECT 244.200 759.750 246.000 762.600 ;
        RECT 247.200 759.750 249.000 763.500 ;
        RECT 250.950 763.500 253.050 765.600 ;
        RECT 253.950 763.500 256.050 765.600 ;
        RECT 256.950 763.500 259.050 765.600 ;
        RECT 261.600 764.400 265.800 765.600 ;
        RECT 250.950 759.750 252.750 763.500 ;
        RECT 253.950 759.750 255.750 763.500 ;
        RECT 256.950 759.750 258.750 763.500 ;
        RECT 261.600 759.750 263.400 764.400 ;
        RECT 267.150 759.750 268.950 765.600 ;
        RECT 272.550 759.750 274.350 765.600 ;
        RECT 276.450 772.950 277.950 785.400 ;
        RECT 289.050 772.950 290.550 785.400 ;
        RECT 295.500 781.350 296.700 785.400 ;
        RECT 301.500 784.500 303.300 791.250 ;
        RECT 304.500 785.400 306.300 791.250 ;
        RECT 308.250 788.400 310.050 791.250 ;
        RECT 308.400 787.200 309.900 788.400 ;
        RECT 307.800 785.100 309.900 787.200 ;
        RECT 311.250 784.950 313.050 791.250 ;
        RECT 314.250 788.400 316.050 791.250 ;
        RECT 297.600 783.300 303.300 784.500 ;
        RECT 304.350 784.050 306.150 784.500 ;
        RECT 310.950 784.050 313.050 784.950 ;
        RECT 297.600 782.700 299.400 783.300 ;
        RECT 304.350 782.850 313.050 784.050 ;
        RECT 304.350 782.700 306.150 782.850 ;
        RECT 314.550 781.350 315.900 788.400 ;
        RECT 318.000 784.500 319.800 791.250 ;
        RECT 321.000 785.400 322.800 791.250 ;
        RECT 324.000 785.400 325.800 791.250 ;
        RECT 327.750 785.400 329.550 791.250 ;
        RECT 330.750 788.400 332.700 791.250 ;
        RECT 333.750 788.400 335.850 791.250 ;
        RECT 336.750 788.400 339.150 791.250 ;
        RECT 331.500 787.050 332.700 788.400 ;
        RECT 334.950 787.050 335.850 788.400 ;
        RECT 337.950 787.050 339.150 788.400 ;
        RECT 340.500 787.950 342.300 791.250 ;
        RECT 331.500 785.400 334.050 787.050 ;
        RECT 324.000 784.500 325.350 785.400 ;
        RECT 331.950 784.950 334.050 785.400 ;
        RECT 334.950 784.950 337.050 787.050 ;
        RECT 337.950 784.950 340.050 787.050 ;
        RECT 318.000 784.200 321.000 784.500 ;
        RECT 317.100 782.400 321.000 784.200 ;
        RECT 322.950 782.850 325.350 784.500 ;
        RECT 322.950 782.400 325.050 782.850 ;
        RECT 343.500 782.700 345.300 791.250 ;
        RECT 346.500 785.400 348.300 791.250 ;
        RECT 349.500 785.400 351.300 791.250 ;
        RECT 352.500 785.400 354.300 791.250 ;
        RECT 350.250 784.500 351.300 785.400 ;
        RECT 350.250 783.600 354.300 784.500 ;
        RECT 332.100 781.650 349.800 782.700 ;
        RECT 276.450 770.850 280.050 772.950 ;
        RECT 286.950 770.850 290.550 772.950 ;
        RECT 276.450 762.600 277.950 770.850 ;
        RECT 289.050 762.600 290.550 770.850 ;
        RECT 276.450 759.750 278.250 762.600 ;
        RECT 279.450 759.750 281.250 762.600 ;
        RECT 285.750 759.750 287.550 762.600 ;
        RECT 288.750 759.750 290.550 762.600 ;
        RECT 292.650 780.450 310.050 781.350 ;
        RECT 292.650 765.600 293.850 780.450 ;
        RECT 294.750 778.350 307.050 779.550 ;
        RECT 307.950 779.250 310.050 780.450 ;
        RECT 313.950 780.600 316.050 781.350 ;
        RECT 332.100 780.600 334.050 781.650 ;
        RECT 348.000 780.900 349.800 781.650 ;
        RECT 313.950 779.250 334.050 780.600 ;
        RECT 334.950 780.150 337.050 780.750 ;
        RECT 334.950 778.950 346.500 780.150 ;
        RECT 334.950 778.650 337.050 778.950 ;
        RECT 344.700 778.350 346.500 778.950 ;
        RECT 294.750 777.750 296.550 778.350 ;
        RECT 306.000 777.450 334.050 778.350 ;
        RECT 306.000 777.150 345.750 777.450 ;
        RECT 298.950 773.100 301.050 777.150 ;
        RECT 332.100 776.550 346.050 777.150 ;
        RECT 302.100 774.000 309.150 775.800 ;
        RECT 298.950 772.050 307.200 773.100 ;
        RECT 294.900 769.200 302.700 771.000 ;
        RECT 306.150 770.250 307.200 772.050 ;
        RECT 308.250 772.350 309.150 774.000 ;
        RECT 310.500 775.650 325.050 776.250 ;
        RECT 310.500 775.050 333.600 775.650 ;
        RECT 342.150 775.350 346.050 776.550 ;
        RECT 310.500 773.250 312.300 775.050 ;
        RECT 322.950 774.450 333.600 775.050 ;
        RECT 322.950 774.150 325.050 774.450 ;
        RECT 331.800 773.850 333.600 774.450 ;
        RECT 334.500 774.450 341.250 775.350 ;
        RECT 343.950 775.050 346.050 775.350 ;
        RECT 318.750 773.250 320.850 773.550 ;
        RECT 308.250 771.300 317.850 772.350 ;
        RECT 318.750 771.450 322.650 773.250 ;
        RECT 334.500 772.950 335.550 774.450 ;
        RECT 323.550 772.050 335.550 772.950 ;
        RECT 316.950 770.550 317.850 771.300 ;
        RECT 323.550 770.550 324.600 772.050 ;
        RECT 336.450 771.750 338.250 773.550 ;
        RECT 340.050 772.050 341.250 774.450 ;
        RECT 349.950 773.850 352.050 775.950 ;
        RECT 350.100 772.050 351.900 773.850 ;
        RECT 306.150 769.200 316.050 770.250 ;
        RECT 316.950 769.200 324.600 770.550 ;
        RECT 325.950 769.350 329.850 771.150 ;
        RECT 301.200 765.600 302.700 769.200 ;
        RECT 315.000 768.300 316.050 769.200 ;
        RECT 325.950 769.050 328.050 769.350 ;
        RECT 333.150 768.300 334.950 768.750 ;
        RECT 336.450 768.300 337.500 771.750 ;
        RECT 340.050 771.000 351.900 772.050 ;
        RECT 353.100 770.100 354.300 783.600 ;
        RECT 358.050 779.400 359.850 791.250 ;
        RECT 361.050 779.400 362.850 791.250 ;
        RECT 364.650 785.400 366.450 791.250 ;
        RECT 367.650 785.400 369.450 791.250 ;
        RECT 307.350 766.500 314.100 768.300 ;
        RECT 315.000 766.500 321.900 768.300 ;
        RECT 333.150 767.850 337.500 768.300 ;
        RECT 329.850 767.100 337.500 767.850 ;
        RECT 339.000 769.200 354.300 770.100 ;
        RECT 329.850 766.950 334.950 767.100 ;
        RECT 329.850 765.600 330.750 766.950 ;
        RECT 339.000 766.050 340.050 769.200 ;
        RECT 348.300 767.700 350.100 768.300 ;
        RECT 292.650 759.750 294.450 765.600 ;
        RECT 298.050 759.750 299.850 765.600 ;
        RECT 301.200 764.400 305.400 765.600 ;
        RECT 303.600 759.750 305.400 764.400 ;
        RECT 307.950 763.500 310.050 765.600 ;
        RECT 310.950 763.500 313.050 765.600 ;
        RECT 313.950 763.500 316.050 765.600 ;
        RECT 318.750 765.300 320.850 765.600 ;
        RECT 308.250 759.750 310.050 763.500 ;
        RECT 311.250 759.750 313.050 763.500 ;
        RECT 314.250 759.750 316.050 763.500 ;
        RECT 318.000 763.500 320.850 765.300 ;
        RECT 322.950 765.300 325.050 765.600 ;
        RECT 322.950 763.500 325.800 765.300 ;
        RECT 326.700 764.250 330.750 765.600 ;
        RECT 326.700 763.800 328.500 764.250 ;
        RECT 331.950 763.950 334.050 766.050 ;
        RECT 334.950 763.950 337.050 766.050 ;
        RECT 337.950 763.950 340.050 766.050 ;
        RECT 341.700 766.500 350.100 767.700 ;
        RECT 341.700 765.600 343.200 766.500 ;
        RECT 353.100 765.600 354.300 769.200 ;
        RECT 318.000 759.750 319.800 763.500 ;
        RECT 321.000 759.750 322.800 762.600 ;
        RECT 324.000 759.750 325.800 763.500 ;
        RECT 331.950 762.600 333.300 763.950 ;
        RECT 334.950 762.600 336.300 763.950 ;
        RECT 337.950 762.600 339.300 763.950 ;
        RECT 328.500 759.750 330.300 762.600 ;
        RECT 331.500 759.750 333.300 762.600 ;
        RECT 334.500 759.750 336.300 762.600 ;
        RECT 337.500 759.750 339.300 762.600 ;
        RECT 341.700 759.750 343.500 765.600 ;
        RECT 347.100 759.750 348.900 765.600 ;
        RECT 352.500 759.750 354.300 765.600 ;
        RECT 358.650 774.150 359.850 779.400 ;
        RECT 358.650 772.050 361.050 774.150 ;
        RECT 361.950 773.850 364.050 775.950 ;
        RECT 362.100 772.050 363.900 773.850 ;
        RECT 358.650 765.600 359.850 772.050 ;
        RECT 365.100 768.300 366.300 785.400 ;
        RECT 377.550 779.400 379.350 791.250 ;
        RECT 380.550 778.500 382.350 791.250 ;
        RECT 383.550 779.400 385.350 791.250 ;
        RECT 386.550 779.400 388.350 791.250 ;
        RECT 389.550 779.400 391.350 791.250 ;
        RECT 403.650 785.400 405.450 791.250 ;
        RECT 406.650 786.000 408.450 791.250 ;
        RECT 404.250 785.100 405.450 785.400 ;
        RECT 409.650 785.400 411.450 791.250 ;
        RECT 412.650 785.400 414.450 791.250 ;
        RECT 409.650 785.100 411.300 785.400 ;
        RECT 404.250 784.200 411.300 785.100 ;
        RECT 386.550 778.500 387.750 779.400 ;
        RECT 380.550 777.600 387.750 778.500 ;
        RECT 368.100 774.150 369.900 775.950 ;
        RECT 380.100 774.150 381.900 775.950 ;
        RECT 386.550 774.150 387.750 777.600 ;
        RECT 404.250 775.950 405.300 784.200 ;
        RECT 412.950 783.450 415.050 784.050 ;
        RECT 412.950 782.550 417.450 783.450 ;
        RECT 412.950 781.950 415.050 782.550 ;
        RECT 410.100 780.150 411.900 781.950 ;
        RECT 406.950 777.150 408.750 778.950 ;
        RECT 409.950 778.050 412.050 780.150 ;
        RECT 413.100 777.150 414.900 778.950 ;
        RECT 367.950 772.050 370.050 774.150 ;
        RECT 379.950 772.050 382.050 774.150 ;
        RECT 385.950 772.050 388.050 774.150 ;
        RECT 403.950 773.850 406.050 775.950 ;
        RECT 406.950 775.050 409.050 777.150 ;
        RECT 412.950 775.050 415.050 777.150 ;
        RECT 361.950 767.100 369.450 768.300 ;
        RECT 386.550 767.700 387.750 772.050 ;
        RECT 404.400 769.650 405.600 773.850 ;
        RECT 412.950 771.450 415.050 772.050 ;
        RECT 416.550 771.450 417.450 782.550 ;
        RECT 421.050 779.400 422.850 791.250 ;
        RECT 424.050 779.400 425.850 791.250 ;
        RECT 427.650 785.400 429.450 791.250 ;
        RECT 430.650 785.400 432.450 791.250 ;
        RECT 439.650 785.400 441.450 791.250 ;
        RECT 442.650 785.400 444.450 791.250 ;
        RECT 445.650 785.400 447.450 791.250 ;
        RECT 454.650 785.400 456.450 791.250 ;
        RECT 457.650 785.400 459.450 791.250 ;
        RECT 460.650 785.400 462.450 791.250 ;
        RECT 412.950 770.550 417.450 771.450 ;
        RECT 421.650 774.150 422.850 779.400 ;
        RECT 421.650 772.050 424.050 774.150 ;
        RECT 424.950 773.850 427.050 775.950 ;
        RECT 425.100 772.050 426.900 773.850 ;
        RECT 412.950 769.950 415.050 770.550 ;
        RECT 404.400 768.000 408.900 769.650 ;
        RECT 361.950 766.500 363.750 767.100 ;
        RECT 358.650 764.100 361.950 765.600 ;
        RECT 360.150 759.750 361.950 764.100 ;
        RECT 363.150 759.750 364.950 765.600 ;
        RECT 367.650 759.750 369.450 767.100 ;
        RECT 380.550 766.500 387.750 767.700 ;
        RECT 380.550 765.600 381.750 766.500 ;
        RECT 386.550 765.600 387.750 766.500 ;
        RECT 377.550 759.750 379.350 765.600 ;
        RECT 380.550 759.750 382.350 765.600 ;
        RECT 383.550 759.750 385.350 765.600 ;
        RECT 386.550 759.750 388.350 765.600 ;
        RECT 389.550 759.750 391.350 765.600 ;
        RECT 407.100 759.750 408.900 768.000 ;
        RECT 412.500 759.750 414.300 768.600 ;
        RECT 421.650 765.600 422.850 772.050 ;
        RECT 428.100 768.300 429.300 785.400 ;
        RECT 443.250 777.150 444.450 785.400 ;
        RECT 454.950 780.450 457.050 781.050 ;
        RECT 452.550 779.550 457.050 780.450 ;
        RECT 431.100 774.150 432.900 775.950 ;
        RECT 430.950 772.050 433.050 774.150 ;
        RECT 439.950 773.850 442.050 775.950 ;
        RECT 442.950 775.050 445.050 777.150 ;
        RECT 440.100 772.050 441.900 773.850 ;
        RECT 424.950 767.100 432.450 768.300 ;
        RECT 443.250 767.700 444.450 775.050 ;
        RECT 445.950 773.850 448.050 775.950 ;
        RECT 446.100 772.050 447.900 773.850 ;
        RECT 424.950 766.500 426.750 767.100 ;
        RECT 421.650 764.100 424.950 765.600 ;
        RECT 423.150 759.750 424.950 764.100 ;
        RECT 426.150 759.750 427.950 765.600 ;
        RECT 430.650 759.750 432.450 767.100 ;
        RECT 440.850 766.800 444.450 767.700 ;
        RECT 445.950 768.450 448.050 769.050 ;
        RECT 452.550 768.450 453.450 779.550 ;
        RECT 454.950 778.950 457.050 779.550 ;
        RECT 458.250 777.150 459.450 785.400 ;
        RECT 470.550 779.400 472.350 791.250 ;
        RECT 474.750 779.400 476.550 791.250 ;
        RECT 482.550 785.400 484.350 791.250 ;
        RECT 485.550 785.400 487.350 791.250 ;
        RECT 499.650 790.500 507.450 791.250 ;
        RECT 474.000 778.350 476.550 779.400 ;
        RECT 454.950 773.850 457.050 775.950 ;
        RECT 457.950 775.050 460.050 777.150 ;
        RECT 455.100 772.050 456.900 773.850 ;
        RECT 445.950 767.550 453.450 768.450 ;
        RECT 458.250 767.700 459.450 775.050 ;
        RECT 460.950 773.850 463.050 775.950 ;
        RECT 470.100 774.150 471.900 775.950 ;
        RECT 461.100 772.050 462.900 773.850 ;
        RECT 469.950 772.050 472.050 774.150 ;
        RECT 474.000 771.150 475.050 778.350 ;
        RECT 476.100 774.150 477.900 775.950 ;
        RECT 475.950 772.050 478.050 774.150 ;
        RECT 485.400 772.950 486.600 785.400 ;
        RECT 499.650 779.400 501.450 790.500 ;
        RECT 502.650 779.400 504.450 789.600 ;
        RECT 505.650 780.600 507.450 790.500 ;
        RECT 508.650 781.500 510.450 791.250 ;
        RECT 511.650 780.600 513.450 791.250 ;
        RECT 505.650 779.700 513.450 780.600 ;
        RECT 522.300 779.400 524.100 791.250 ;
        RECT 526.500 779.400 528.300 791.250 ;
        RECT 529.800 785.400 531.600 791.250 ;
        RECT 538.650 790.500 546.450 791.250 ;
        RECT 538.650 779.400 540.450 790.500 ;
        RECT 541.650 779.400 543.450 789.600 ;
        RECT 544.650 780.600 546.450 790.500 ;
        RECT 547.650 781.500 549.450 791.250 ;
        RECT 550.650 780.600 552.450 791.250 ;
        RECT 544.650 779.700 552.450 780.600 ;
        RECT 558.450 779.400 560.250 791.250 ;
        RECT 562.650 779.400 564.450 791.250 ;
        RECT 569.550 785.400 571.350 791.250 ;
        RECT 572.550 785.400 574.350 791.250 ;
        RECT 583.650 785.400 585.450 791.250 ;
        RECT 586.650 785.400 588.450 791.250 ;
        RECT 589.650 785.400 591.450 791.250 ;
        RECT 502.800 778.500 504.600 779.400 ;
        RECT 502.800 777.600 506.850 778.500 ;
        RECT 500.100 774.150 501.900 775.950 ;
        RECT 505.950 774.150 506.850 777.600 ;
        RECT 511.950 774.150 513.750 775.950 ;
        RECT 521.100 774.150 522.900 775.950 ;
        RECT 526.950 774.150 528.150 779.400 ;
        RECT 529.950 777.150 531.750 778.950 ;
        RECT 541.800 778.500 543.600 779.400 ;
        RECT 541.800 777.600 545.850 778.500 ;
        RECT 558.450 778.350 561.000 779.400 ;
        RECT 529.950 775.050 532.050 777.150 ;
        RECT 539.100 774.150 540.900 775.950 ;
        RECT 544.950 774.150 545.850 777.600 ;
        RECT 550.950 774.150 552.750 775.950 ;
        RECT 557.100 774.150 558.900 775.950 ;
        RECT 482.100 771.150 483.900 772.950 ;
        RECT 472.950 769.050 475.050 771.150 ;
        RECT 481.950 769.050 484.050 771.150 ;
        RECT 484.950 770.850 487.050 772.950 ;
        RECT 499.950 772.050 502.050 774.150 ;
        RECT 502.950 770.850 505.050 772.950 ;
        RECT 505.950 772.050 508.050 774.150 ;
        RECT 445.950 766.950 448.050 767.550 ;
        RECT 455.850 766.800 459.450 767.700 ;
        RECT 440.850 759.750 442.650 766.800 ;
        RECT 445.350 759.750 447.150 765.600 ;
        RECT 455.850 759.750 457.650 766.800 ;
        RECT 460.350 759.750 462.150 765.600 ;
        RECT 474.000 762.600 475.050 769.050 ;
        RECT 485.400 762.600 486.600 770.850 ;
        RECT 503.250 769.050 505.050 770.850 ;
        RECT 507.000 765.600 508.050 772.050 ;
        RECT 508.950 770.850 511.050 772.950 ;
        RECT 511.950 772.050 514.050 774.150 ;
        RECT 520.950 772.050 523.050 774.150 ;
        RECT 523.950 770.850 526.050 772.950 ;
        RECT 526.950 772.050 529.050 774.150 ;
        RECT 538.950 772.050 541.050 774.150 ;
        RECT 508.950 769.050 510.750 770.850 ;
        RECT 524.100 769.050 525.900 770.850 ;
        RECT 527.850 768.750 529.050 772.050 ;
        RECT 541.950 770.850 544.050 772.950 ;
        RECT 544.950 772.050 547.050 774.150 ;
        RECT 542.250 769.050 544.050 770.850 ;
        RECT 528.000 767.700 531.750 768.750 ;
        RECT 470.550 759.750 472.350 762.600 ;
        RECT 473.550 759.750 475.350 762.600 ;
        RECT 476.550 759.750 478.350 762.600 ;
        RECT 482.550 759.750 484.350 762.600 ;
        RECT 485.550 759.750 487.350 762.600 ;
        RECT 502.800 759.750 504.600 765.600 ;
        RECT 507.000 759.750 508.800 765.600 ;
        RECT 511.200 759.750 513.000 765.600 ;
        RECT 521.550 764.700 529.350 766.050 ;
        RECT 521.550 759.750 523.350 764.700 ;
        RECT 524.550 759.750 526.350 763.800 ;
        RECT 527.550 759.750 529.350 764.700 ;
        RECT 530.550 765.600 531.750 767.700 ;
        RECT 546.000 765.600 547.050 772.050 ;
        RECT 547.950 770.850 550.050 772.950 ;
        RECT 550.950 772.050 553.050 774.150 ;
        RECT 556.950 772.050 559.050 774.150 ;
        RECT 559.950 771.150 561.000 778.350 ;
        RECT 563.100 774.150 564.900 775.950 ;
        RECT 562.950 772.050 565.050 774.150 ;
        RECT 572.400 772.950 573.600 785.400 ;
        RECT 587.250 777.150 588.450 785.400 ;
        RECT 597.300 779.400 599.100 791.250 ;
        RECT 601.500 779.400 603.300 791.250 ;
        RECT 604.800 785.400 606.600 791.250 ;
        RECT 619.650 785.400 621.450 791.250 ;
        RECT 622.650 785.400 624.450 791.250 ;
        RECT 625.650 785.400 627.450 791.250 ;
        RECT 632.550 785.400 634.350 791.250 ;
        RECT 635.550 785.400 637.350 791.250 ;
        RECT 583.950 773.850 586.050 775.950 ;
        RECT 586.950 775.050 589.050 777.150 ;
        RECT 569.100 771.150 570.900 772.950 ;
        RECT 547.950 769.050 549.750 770.850 ;
        RECT 559.950 769.050 562.050 771.150 ;
        RECT 568.950 769.050 571.050 771.150 ;
        RECT 571.950 770.850 574.050 772.950 ;
        RECT 584.100 772.050 585.900 773.850 ;
        RECT 530.550 759.750 532.350 765.600 ;
        RECT 541.800 759.750 543.600 765.600 ;
        RECT 546.000 759.750 547.800 765.600 ;
        RECT 550.200 759.750 552.000 765.600 ;
        RECT 559.950 762.600 561.000 769.050 ;
        RECT 572.400 762.600 573.600 770.850 ;
        RECT 587.250 767.700 588.450 775.050 ;
        RECT 589.950 773.850 592.050 775.950 ;
        RECT 596.100 774.150 597.900 775.950 ;
        RECT 601.950 774.150 603.150 779.400 ;
        RECT 604.950 777.150 606.750 778.950 ;
        RECT 623.250 777.150 624.450 785.400 ;
        RECT 604.950 775.050 607.050 777.150 ;
        RECT 590.100 772.050 591.900 773.850 ;
        RECT 595.950 772.050 598.050 774.150 ;
        RECT 598.950 770.850 601.050 772.950 ;
        RECT 601.950 772.050 604.050 774.150 ;
        RECT 619.950 773.850 622.050 775.950 ;
        RECT 622.950 775.050 625.050 777.150 ;
        RECT 620.100 772.050 621.900 773.850 ;
        RECT 599.100 769.050 600.900 770.850 ;
        RECT 602.850 768.750 604.050 772.050 ;
        RECT 603.000 767.700 606.750 768.750 ;
        RECT 623.250 767.700 624.450 775.050 ;
        RECT 625.950 773.850 628.050 775.950 ;
        RECT 626.100 772.050 627.900 773.850 ;
        RECT 635.400 772.950 636.600 785.400 ;
        RECT 651.450 779.400 653.250 791.250 ;
        RECT 655.650 779.400 657.450 791.250 ;
        RECT 666.300 779.400 668.100 791.250 ;
        RECT 670.500 779.400 672.300 791.250 ;
        RECT 673.800 785.400 675.600 791.250 ;
        RECT 680.550 779.400 682.350 791.250 ;
        RECT 684.750 779.400 686.550 791.250 ;
        RECT 692.550 785.400 694.350 791.250 ;
        RECT 695.550 785.400 697.350 791.250 ;
        RECT 698.550 785.400 700.350 791.250 ;
        RECT 709.650 785.400 711.450 791.250 ;
        RECT 712.650 785.400 714.450 791.250 ;
        RECT 722.550 785.400 724.350 791.250 ;
        RECT 725.550 785.400 727.350 791.250 ;
        RECT 728.550 786.000 730.350 791.250 ;
        RECT 651.450 778.350 654.000 779.400 ;
        RECT 650.100 774.150 651.900 775.950 ;
        RECT 632.100 771.150 633.900 772.950 ;
        RECT 631.950 769.050 634.050 771.150 ;
        RECT 634.950 770.850 637.050 772.950 ;
        RECT 649.950 772.050 652.050 774.150 ;
        RECT 652.950 771.150 654.000 778.350 ;
        RECT 656.100 774.150 657.900 775.950 ;
        RECT 665.100 774.150 666.900 775.950 ;
        RECT 670.950 774.150 672.150 779.400 ;
        RECT 673.950 777.150 675.750 778.950 ;
        RECT 684.000 778.350 686.550 779.400 ;
        RECT 673.950 775.050 676.050 777.150 ;
        RECT 680.100 774.150 681.900 775.950 ;
        RECT 655.950 772.050 658.050 774.150 ;
        RECT 664.950 772.050 667.050 774.150 ;
        RECT 584.850 766.800 588.450 767.700 ;
        RECT 556.650 759.750 558.450 762.600 ;
        RECT 559.650 759.750 561.450 762.600 ;
        RECT 562.650 759.750 564.450 762.600 ;
        RECT 569.550 759.750 571.350 762.600 ;
        RECT 572.550 759.750 574.350 762.600 ;
        RECT 584.850 759.750 586.650 766.800 ;
        RECT 589.350 759.750 591.150 765.600 ;
        RECT 596.550 764.700 604.350 766.050 ;
        RECT 596.550 759.750 598.350 764.700 ;
        RECT 599.550 759.750 601.350 763.800 ;
        RECT 602.550 759.750 604.350 764.700 ;
        RECT 605.550 765.600 606.750 767.700 ;
        RECT 620.850 766.800 624.450 767.700 ;
        RECT 605.550 759.750 607.350 765.600 ;
        RECT 620.850 759.750 622.650 766.800 ;
        RECT 625.350 759.750 627.150 765.600 ;
        RECT 635.400 762.600 636.600 770.850 ;
        RECT 652.950 769.050 655.050 771.150 ;
        RECT 667.950 770.850 670.050 772.950 ;
        RECT 670.950 772.050 673.050 774.150 ;
        RECT 679.950 772.050 682.050 774.150 ;
        RECT 668.100 769.050 669.900 770.850 ;
        RECT 652.950 762.600 654.000 769.050 ;
        RECT 671.850 768.750 673.050 772.050 ;
        RECT 684.000 771.150 685.050 778.350 ;
        RECT 695.550 777.150 696.750 785.400 ;
        RECT 700.950 783.450 703.050 784.050 ;
        RECT 706.950 783.450 709.050 784.050 ;
        RECT 700.950 782.550 709.050 783.450 ;
        RECT 700.950 781.950 703.050 782.550 ;
        RECT 706.950 781.950 709.050 782.550 ;
        RECT 686.100 774.150 687.900 775.950 ;
        RECT 685.950 772.050 688.050 774.150 ;
        RECT 691.950 773.850 694.050 775.950 ;
        RECT 694.950 775.050 697.050 777.150 ;
        RECT 692.100 772.050 693.900 773.850 ;
        RECT 682.950 769.050 685.050 771.150 ;
        RECT 672.000 767.700 675.750 768.750 ;
        RECT 665.550 764.700 673.350 766.050 ;
        RECT 632.550 759.750 634.350 762.600 ;
        RECT 635.550 759.750 637.350 762.600 ;
        RECT 649.650 759.750 651.450 762.600 ;
        RECT 652.650 759.750 654.450 762.600 ;
        RECT 655.650 759.750 657.450 762.600 ;
        RECT 665.550 759.750 667.350 764.700 ;
        RECT 668.550 759.750 670.350 763.800 ;
        RECT 671.550 759.750 673.350 764.700 ;
        RECT 674.550 765.600 675.750 767.700 ;
        RECT 674.550 759.750 676.350 765.600 ;
        RECT 684.000 762.600 685.050 769.050 ;
        RECT 695.550 767.700 696.750 775.050 ;
        RECT 697.950 773.850 700.050 775.950 ;
        RECT 698.100 772.050 699.900 773.850 ;
        RECT 710.400 772.950 711.600 785.400 ;
        RECT 725.700 785.100 727.350 785.400 ;
        RECT 731.550 785.400 733.350 791.250 ;
        RECT 737.550 785.400 739.350 791.250 ;
        RECT 740.550 785.400 742.350 791.250 ;
        RECT 743.550 785.400 745.350 791.250 ;
        RECT 752.400 785.400 754.200 791.250 ;
        RECT 731.550 785.100 732.750 785.400 ;
        RECT 725.700 784.200 732.750 785.100 ;
        RECT 725.100 780.150 726.900 781.950 ;
        RECT 722.100 777.150 723.900 778.950 ;
        RECT 724.950 778.050 727.050 780.150 ;
        RECT 728.250 777.150 730.050 778.950 ;
        RECT 721.950 775.050 724.050 777.150 ;
        RECT 727.950 775.050 730.050 777.150 ;
        RECT 731.700 775.950 732.750 784.200 ;
        RECT 740.550 777.150 741.750 785.400 ;
        RECT 755.700 779.400 757.500 791.250 ;
        RECT 759.900 779.400 761.700 791.250 ;
        RECT 767.550 779.400 769.350 791.250 ;
        RECT 772.050 779.550 773.850 791.250 ;
        RECT 775.050 780.900 776.850 791.250 ;
        RECT 788.550 785.400 790.350 791.250 ;
        RECT 791.550 785.400 793.350 791.250 ;
        RECT 794.550 785.400 796.350 791.250 ;
        RECT 803.550 785.400 805.350 791.250 ;
        RECT 806.550 785.400 808.350 791.250 ;
        RECT 809.550 785.400 811.350 791.250 ;
        RECT 775.050 779.550 777.450 780.900 ;
        RECT 752.250 777.150 754.050 778.950 ;
        RECT 730.950 773.850 733.050 775.950 ;
        RECT 736.950 773.850 739.050 775.950 ;
        RECT 739.950 775.050 742.050 777.150 ;
        RECT 709.950 770.850 712.050 772.950 ;
        RECT 713.100 771.150 714.900 772.950 ;
        RECT 695.550 766.800 699.150 767.700 ;
        RECT 680.550 759.750 682.350 762.600 ;
        RECT 683.550 759.750 685.350 762.600 ;
        RECT 686.550 759.750 688.350 762.600 ;
        RECT 692.850 759.750 694.650 765.600 ;
        RECT 697.350 759.750 699.150 766.800 ;
        RECT 710.400 762.600 711.600 770.850 ;
        RECT 712.950 769.050 715.050 771.150 ;
        RECT 731.400 769.650 732.600 773.850 ;
        RECT 737.100 772.050 738.900 773.850 ;
        RECT 709.650 759.750 711.450 762.600 ;
        RECT 712.650 759.750 714.450 762.600 ;
        RECT 722.700 759.750 724.500 768.600 ;
        RECT 728.100 768.000 732.600 769.650 ;
        RECT 728.100 759.750 729.900 768.000 ;
        RECT 740.550 767.700 741.750 775.050 ;
        RECT 742.950 773.850 745.050 775.950 ;
        RECT 751.950 775.050 754.050 777.150 ;
        RECT 755.850 774.150 757.050 779.400 ;
        RECT 767.550 778.200 768.750 779.400 ;
        RECT 772.950 778.200 774.750 778.650 ;
        RECT 767.550 777.000 774.750 778.200 ;
        RECT 772.950 776.850 774.750 777.000 ;
        RECT 761.100 774.150 762.900 775.950 ;
        RECT 770.100 774.150 771.900 775.950 ;
        RECT 743.100 772.050 744.900 773.850 ;
        RECT 754.950 772.050 757.050 774.150 ;
        RECT 754.950 768.750 756.150 772.050 ;
        RECT 757.950 770.850 760.050 772.950 ;
        RECT 760.950 772.050 763.050 774.150 ;
        RECT 767.100 771.150 768.900 772.950 ;
        RECT 769.950 772.050 772.050 774.150 ;
        RECT 758.100 769.050 759.900 770.850 ;
        RECT 766.950 769.050 769.050 771.150 ;
        RECT 752.250 767.700 756.000 768.750 ;
        RECT 773.700 768.600 774.600 776.850 ;
        RECT 776.100 772.950 777.450 779.550 ;
        RECT 791.550 777.150 792.750 785.400 ;
        RECT 806.550 777.150 807.750 785.400 ;
        RECT 822.450 779.400 824.250 791.250 ;
        RECT 826.650 779.400 828.450 791.250 ;
        RECT 833.550 779.400 835.350 791.250 ;
        RECT 837.750 779.400 839.550 791.250 ;
        RECT 848.550 779.400 850.350 791.250 ;
        RECT 851.550 779.400 853.350 791.250 ;
        RECT 822.450 778.350 825.000 779.400 ;
        RECT 787.950 773.850 790.050 775.950 ;
        RECT 790.950 775.050 793.050 777.150 ;
        RECT 775.950 770.850 778.050 772.950 ;
        RECT 788.100 772.050 789.900 773.850 ;
        RECT 772.950 767.700 774.750 768.600 ;
        RECT 740.550 766.800 744.150 767.700 ;
        RECT 737.850 759.750 739.650 765.600 ;
        RECT 742.350 759.750 744.150 766.800 ;
        RECT 752.250 765.600 753.450 767.700 ;
        RECT 771.450 766.800 774.750 767.700 ;
        RECT 751.650 759.750 753.450 765.600 ;
        RECT 754.650 764.700 762.450 766.050 ;
        RECT 754.650 759.750 756.450 764.700 ;
        RECT 757.650 759.750 759.450 763.800 ;
        RECT 760.650 759.750 762.450 764.700 ;
        RECT 771.450 762.600 772.350 766.800 ;
        RECT 777.000 765.600 778.050 770.850 ;
        RECT 791.550 767.700 792.750 775.050 ;
        RECT 793.950 773.850 796.050 775.950 ;
        RECT 802.950 773.850 805.050 775.950 ;
        RECT 805.950 775.050 808.050 777.150 ;
        RECT 794.100 772.050 795.900 773.850 ;
        RECT 803.100 772.050 804.900 773.850 ;
        RECT 806.550 767.700 807.750 775.050 ;
        RECT 808.950 773.850 811.050 775.950 ;
        RECT 821.100 774.150 822.900 775.950 ;
        RECT 809.100 772.050 810.900 773.850 ;
        RECT 820.950 772.050 823.050 774.150 ;
        RECT 823.950 771.150 825.000 778.350 ;
        RECT 837.000 778.350 839.550 779.400 ;
        RECT 827.100 774.150 828.900 775.950 ;
        RECT 833.100 774.150 834.900 775.950 ;
        RECT 826.950 772.050 829.050 774.150 ;
        RECT 832.950 772.050 835.050 774.150 ;
        RECT 837.000 771.150 838.050 778.350 ;
        RECT 839.100 774.150 840.900 775.950 ;
        RECT 851.400 774.150 852.600 779.400 ;
        RECT 838.950 772.050 841.050 774.150 ;
        RECT 823.950 769.050 826.050 771.150 ;
        RECT 835.950 769.050 838.050 771.150 ;
        RECT 847.950 770.850 850.050 772.950 ;
        RECT 850.950 772.050 853.050 774.150 ;
        RECT 848.100 769.050 849.900 770.850 ;
        RECT 791.550 766.800 795.150 767.700 ;
        RECT 806.550 766.800 810.150 767.700 ;
        RECT 767.550 759.750 769.350 762.600 ;
        RECT 770.550 759.750 772.350 762.600 ;
        RECT 773.550 759.750 775.350 762.600 ;
        RECT 776.550 759.750 778.350 765.600 ;
        RECT 788.850 759.750 790.650 765.600 ;
        RECT 793.350 759.750 795.150 766.800 ;
        RECT 803.850 759.750 805.650 765.600 ;
        RECT 808.350 759.750 810.150 766.800 ;
        RECT 823.950 762.600 825.000 769.050 ;
        RECT 837.000 762.600 838.050 769.050 ;
        RECT 851.400 765.600 852.600 772.050 ;
        RECT 820.650 759.750 822.450 762.600 ;
        RECT 823.650 759.750 825.450 762.600 ;
        RECT 826.650 759.750 828.450 762.600 ;
        RECT 833.550 759.750 835.350 762.600 ;
        RECT 836.550 759.750 838.350 762.600 ;
        RECT 839.550 759.750 841.350 762.600 ;
        RECT 848.550 759.750 850.350 765.600 ;
        RECT 851.550 759.750 853.350 765.600 ;
        RECT 2.700 749.400 4.500 755.250 ;
        RECT 8.100 749.400 9.900 755.250 ;
        RECT 13.500 749.400 15.300 755.250 ;
        RECT 17.700 752.400 19.500 755.250 ;
        RECT 20.700 752.400 22.500 755.250 ;
        RECT 23.700 752.400 25.500 755.250 ;
        RECT 26.700 752.400 28.500 755.250 ;
        RECT 17.700 751.050 19.050 752.400 ;
        RECT 20.700 751.050 22.050 752.400 ;
        RECT 23.700 751.050 25.050 752.400 ;
        RECT 31.200 751.500 33.000 755.250 ;
        RECT 34.200 752.400 36.000 755.250 ;
        RECT 37.200 751.500 39.000 755.250 ;
        RECT 2.700 745.800 3.900 749.400 ;
        RECT 13.800 748.500 15.300 749.400 ;
        RECT 6.900 747.300 15.300 748.500 ;
        RECT 16.950 748.950 19.050 751.050 ;
        RECT 19.950 748.950 22.050 751.050 ;
        RECT 22.950 748.950 25.050 751.050 ;
        RECT 28.500 750.750 30.300 751.200 ;
        RECT 26.250 749.400 30.300 750.750 ;
        RECT 31.200 749.700 34.050 751.500 ;
        RECT 31.950 749.400 34.050 749.700 ;
        RECT 36.150 749.700 39.000 751.500 ;
        RECT 40.950 751.500 42.750 755.250 ;
        RECT 43.950 751.500 45.750 755.250 ;
        RECT 46.950 751.500 48.750 755.250 ;
        RECT 36.150 749.400 38.250 749.700 ;
        RECT 40.950 749.400 43.050 751.500 ;
        RECT 43.950 749.400 46.050 751.500 ;
        RECT 46.950 749.400 49.050 751.500 ;
        RECT 51.600 750.600 53.400 755.250 ;
        RECT 51.600 749.400 55.800 750.600 ;
        RECT 57.150 749.400 58.950 755.250 ;
        RECT 62.550 749.400 64.350 755.250 ;
        RECT 6.900 746.700 8.700 747.300 ;
        RECT 16.950 745.800 18.000 748.950 ;
        RECT 26.250 748.050 27.150 749.400 ;
        RECT 22.050 747.900 27.150 748.050 ;
        RECT 2.700 744.900 18.000 745.800 ;
        RECT 19.500 747.150 27.150 747.900 ;
        RECT 19.500 746.700 23.850 747.150 ;
        RECT 35.100 746.700 42.000 748.500 ;
        RECT 42.900 746.700 49.650 748.500 ;
        RECT 2.700 731.400 3.900 744.900 ;
        RECT 5.100 742.950 16.950 744.000 ;
        RECT 19.500 743.250 20.550 746.700 ;
        RECT 22.050 746.250 23.850 746.700 ;
        RECT 28.950 745.650 31.050 745.950 ;
        RECT 40.950 745.800 42.000 746.700 ;
        RECT 54.300 745.800 55.800 749.400 ;
        RECT 27.150 743.850 31.050 745.650 ;
        RECT 32.400 744.450 40.050 745.800 ;
        RECT 40.950 744.750 50.850 745.800 ;
        RECT 5.100 741.150 6.900 742.950 ;
        RECT 4.950 739.050 7.050 741.150 ;
        RECT 15.750 740.550 16.950 742.950 ;
        RECT 18.750 741.450 20.550 743.250 ;
        RECT 32.400 742.950 33.450 744.450 ;
        RECT 39.150 743.700 40.050 744.450 ;
        RECT 21.450 742.050 33.450 742.950 ;
        RECT 21.450 740.550 22.500 742.050 ;
        RECT 34.350 741.750 38.250 743.550 ;
        RECT 39.150 742.650 48.750 743.700 ;
        RECT 36.150 741.450 38.250 741.750 ;
        RECT 10.950 739.650 13.050 739.950 ;
        RECT 15.750 739.650 22.500 740.550 ;
        RECT 23.400 740.550 25.200 741.150 ;
        RECT 31.950 740.550 34.050 740.850 ;
        RECT 23.400 739.950 34.050 740.550 ;
        RECT 44.700 739.950 46.500 741.750 ;
        RECT 10.950 738.450 14.850 739.650 ;
        RECT 23.400 739.350 46.500 739.950 ;
        RECT 31.950 738.750 46.500 739.350 ;
        RECT 47.850 741.000 48.750 742.650 ;
        RECT 49.800 742.950 50.850 744.750 ;
        RECT 54.300 744.000 62.100 745.800 ;
        RECT 49.800 741.900 58.050 742.950 ;
        RECT 47.850 739.200 54.900 741.000 ;
        RECT 10.950 737.850 24.900 738.450 ;
        RECT 55.950 737.850 58.050 741.900 ;
        RECT 11.250 737.550 51.000 737.850 ;
        RECT 22.950 736.650 51.000 737.550 ;
        RECT 60.450 736.650 62.250 737.250 ;
        RECT 10.500 736.050 12.300 736.650 ;
        RECT 19.950 736.050 22.050 736.350 ;
        RECT 10.500 734.850 22.050 736.050 ;
        RECT 19.950 734.250 22.050 734.850 ;
        RECT 22.950 734.400 43.050 735.750 ;
        RECT 7.200 733.350 9.000 734.100 ;
        RECT 22.950 733.350 24.900 734.400 ;
        RECT 40.950 733.650 43.050 734.400 ;
        RECT 46.950 734.550 49.050 735.750 ;
        RECT 49.950 735.450 62.250 736.650 ;
        RECT 63.150 734.550 64.350 749.400 ;
        RECT 46.950 733.650 64.350 734.550 ;
        RECT 66.450 752.400 68.250 755.250 ;
        RECT 69.450 752.400 71.250 755.250 ;
        RECT 74.550 752.400 76.350 755.250 ;
        RECT 77.550 752.400 79.350 755.250 ;
        RECT 80.550 752.400 82.350 755.250 ;
        RECT 66.450 744.150 67.950 752.400 ;
        RECT 78.000 745.950 79.050 752.400 ;
        RECT 95.850 748.200 97.650 755.250 ;
        RECT 100.350 749.400 102.150 755.250 ;
        RECT 106.650 749.400 108.450 755.250 ;
        RECT 95.850 747.300 99.450 748.200 ;
        RECT 66.450 742.050 70.050 744.150 ;
        RECT 76.950 743.850 79.050 745.950 ;
        RECT 7.200 732.300 24.900 733.350 ;
        RECT 2.700 730.500 6.750 731.400 ;
        RECT 5.700 729.600 6.750 730.500 ;
        RECT 2.700 723.750 4.500 729.600 ;
        RECT 5.700 723.750 7.500 729.600 ;
        RECT 8.700 723.750 10.500 729.600 ;
        RECT 11.700 723.750 13.500 732.300 ;
        RECT 31.950 732.150 34.050 732.600 ;
        RECT 31.650 730.500 34.050 732.150 ;
        RECT 36.000 730.800 39.900 732.600 ;
        RECT 36.000 730.500 39.000 730.800 ;
        RECT 16.950 727.950 19.050 730.050 ;
        RECT 19.950 727.950 22.050 730.050 ;
        RECT 22.950 729.600 25.050 730.050 ;
        RECT 31.650 729.600 33.000 730.500 ;
        RECT 22.950 727.950 25.500 729.600 ;
        RECT 14.700 723.750 16.500 727.050 ;
        RECT 17.850 726.600 19.050 727.950 ;
        RECT 21.150 726.600 22.050 727.950 ;
        RECT 24.300 726.600 25.500 727.950 ;
        RECT 17.850 723.750 20.250 726.600 ;
        RECT 21.150 723.750 23.250 726.600 ;
        RECT 24.300 723.750 26.250 726.600 ;
        RECT 27.450 723.750 29.250 729.600 ;
        RECT 31.200 723.750 33.000 729.600 ;
        RECT 34.200 723.750 36.000 729.600 ;
        RECT 37.200 723.750 39.000 730.500 ;
        RECT 41.100 726.600 42.450 733.650 ;
        RECT 50.850 732.150 52.650 732.300 ;
        RECT 43.950 730.950 52.650 732.150 ;
        RECT 57.600 731.700 59.400 732.300 ;
        RECT 43.950 730.050 46.050 730.950 ;
        RECT 50.850 730.500 52.650 730.950 ;
        RECT 53.700 730.500 59.400 731.700 ;
        RECT 40.950 723.750 42.750 726.600 ;
        RECT 43.950 723.750 45.750 730.050 ;
        RECT 47.100 727.800 49.200 729.900 ;
        RECT 47.100 726.600 48.600 727.800 ;
        RECT 46.950 723.750 48.750 726.600 ;
        RECT 50.700 723.750 52.500 729.600 ;
        RECT 53.700 723.750 55.500 730.500 ;
        RECT 60.300 729.600 61.500 733.650 ;
        RECT 66.450 729.600 67.950 742.050 ;
        RECT 73.950 740.850 76.050 742.950 ;
        RECT 74.100 739.050 75.900 740.850 ;
        RECT 78.000 736.650 79.050 743.850 ;
        RECT 79.950 740.850 82.050 742.950 ;
        RECT 95.100 741.150 96.900 742.950 ;
        RECT 80.100 739.050 81.900 740.850 ;
        RECT 94.950 739.050 97.050 741.150 ;
        RECT 98.250 739.950 99.450 747.300 ;
        RECT 107.250 747.300 108.450 749.400 ;
        RECT 109.650 750.300 111.450 755.250 ;
        RECT 112.650 751.200 114.450 755.250 ;
        RECT 115.650 750.300 117.450 755.250 ;
        RECT 127.650 752.400 129.450 755.250 ;
        RECT 130.650 752.400 132.450 755.250 ;
        RECT 142.650 752.400 144.450 755.250 ;
        RECT 145.650 752.400 147.450 755.250 ;
        RECT 109.650 748.950 117.450 750.300 ;
        RECT 107.250 746.250 111.000 747.300 ;
        RECT 109.950 742.950 111.150 746.250 ;
        RECT 113.100 744.150 114.900 745.950 ;
        RECT 128.400 744.150 129.600 752.400 ;
        RECT 101.100 741.150 102.900 742.950 ;
        RECT 97.950 737.850 100.050 739.950 ;
        RECT 100.950 739.050 103.050 741.150 ;
        RECT 109.950 740.850 112.050 742.950 ;
        RECT 112.950 742.050 115.050 744.150 ;
        RECT 115.950 740.850 118.050 742.950 ;
        RECT 127.950 742.050 130.050 744.150 ;
        RECT 130.950 743.850 133.050 745.950 ;
        RECT 143.400 744.150 144.600 752.400 ;
        RECT 150.000 749.400 151.800 755.250 ;
        RECT 154.200 751.050 156.000 755.250 ;
        RECT 157.500 752.400 159.300 755.250 ;
        RECT 165.750 752.400 167.550 755.250 ;
        RECT 168.750 752.400 170.550 755.250 ;
        RECT 154.200 749.400 159.900 751.050 ;
        RECT 131.100 742.050 132.900 743.850 ;
        RECT 142.950 742.050 145.050 744.150 ;
        RECT 145.950 743.850 148.050 745.950 ;
        RECT 149.100 744.150 150.900 745.950 ;
        RECT 146.100 742.050 147.900 743.850 ;
        RECT 148.950 742.050 151.050 744.150 ;
        RECT 151.950 743.850 154.050 745.950 ;
        RECT 155.100 744.150 156.900 745.950 ;
        RECT 152.100 742.050 153.900 743.850 ;
        RECT 154.950 742.050 157.050 744.150 ;
        RECT 158.700 742.950 159.900 749.400 ;
        RECT 169.050 744.150 170.550 752.400 ;
        RECT 106.950 737.850 109.050 739.950 ;
        RECT 78.000 735.600 80.550 736.650 ;
        RECT 56.700 723.750 58.500 729.600 ;
        RECT 59.700 723.750 61.500 729.600 ;
        RECT 62.700 723.750 64.500 729.600 ;
        RECT 66.450 723.750 68.250 729.600 ;
        RECT 69.450 723.750 71.250 729.600 ;
        RECT 74.550 723.750 76.350 735.600 ;
        RECT 78.750 723.750 80.550 735.600 ;
        RECT 98.250 729.600 99.450 737.850 ;
        RECT 107.250 736.050 109.050 737.850 ;
        RECT 110.850 735.600 112.050 740.850 ;
        RECT 116.100 739.050 117.900 740.850 ;
        RECT 94.650 723.750 96.450 729.600 ;
        RECT 97.650 723.750 99.450 729.600 ;
        RECT 100.650 723.750 102.450 729.600 ;
        RECT 107.400 723.750 109.200 729.600 ;
        RECT 110.700 723.750 112.500 735.600 ;
        RECT 114.900 723.750 116.700 735.600 ;
        RECT 128.400 729.600 129.600 742.050 ;
        RECT 143.400 729.600 144.600 742.050 ;
        RECT 157.950 740.850 160.050 742.950 ;
        RECT 166.950 742.050 170.550 744.150 ;
        RECT 158.700 735.600 159.900 740.850 ;
        RECT 149.550 734.700 157.350 735.600 ;
        RECT 127.650 723.750 129.450 729.600 ;
        RECT 130.650 723.750 132.450 729.600 ;
        RECT 142.650 723.750 144.450 729.600 ;
        RECT 145.650 723.750 147.450 729.600 ;
        RECT 149.550 723.750 151.350 734.700 ;
        RECT 152.550 723.750 154.350 733.800 ;
        RECT 155.550 723.750 157.350 734.700 ;
        RECT 158.550 723.750 160.350 735.600 ;
        RECT 169.050 729.600 170.550 742.050 ;
        RECT 172.650 749.400 174.450 755.250 ;
        RECT 178.050 749.400 179.850 755.250 ;
        RECT 183.600 750.600 185.400 755.250 ;
        RECT 188.250 751.500 190.050 755.250 ;
        RECT 191.250 751.500 193.050 755.250 ;
        RECT 194.250 751.500 196.050 755.250 ;
        RECT 181.200 749.400 185.400 750.600 ;
        RECT 187.950 749.400 190.050 751.500 ;
        RECT 190.950 749.400 193.050 751.500 ;
        RECT 193.950 749.400 196.050 751.500 ;
        RECT 198.000 751.500 199.800 755.250 ;
        RECT 201.000 752.400 202.800 755.250 ;
        RECT 204.000 751.500 205.800 755.250 ;
        RECT 208.500 752.400 210.300 755.250 ;
        RECT 211.500 752.400 213.300 755.250 ;
        RECT 214.500 752.400 216.300 755.250 ;
        RECT 217.500 752.400 219.300 755.250 ;
        RECT 198.000 749.700 200.850 751.500 ;
        RECT 198.750 749.400 200.850 749.700 ;
        RECT 202.950 749.700 205.800 751.500 ;
        RECT 206.700 750.750 208.500 751.200 ;
        RECT 211.950 751.050 213.300 752.400 ;
        RECT 214.950 751.050 216.300 752.400 ;
        RECT 217.950 751.050 219.300 752.400 ;
        RECT 202.950 749.400 205.050 749.700 ;
        RECT 206.700 749.400 210.750 750.750 ;
        RECT 172.650 734.550 173.850 749.400 ;
        RECT 181.200 745.800 182.700 749.400 ;
        RECT 187.350 746.700 194.100 748.500 ;
        RECT 195.000 746.700 201.900 748.500 ;
        RECT 209.850 748.050 210.750 749.400 ;
        RECT 211.950 748.950 214.050 751.050 ;
        RECT 214.950 748.950 217.050 751.050 ;
        RECT 217.950 748.950 220.050 751.050 ;
        RECT 209.850 747.900 214.950 748.050 ;
        RECT 209.850 747.150 217.500 747.900 ;
        RECT 213.150 746.700 217.500 747.150 ;
        RECT 195.000 745.800 196.050 746.700 ;
        RECT 213.150 746.250 214.950 746.700 ;
        RECT 174.900 744.000 182.700 745.800 ;
        RECT 186.150 744.750 196.050 745.800 ;
        RECT 186.150 742.950 187.200 744.750 ;
        RECT 196.950 744.450 204.600 745.800 ;
        RECT 196.950 743.700 197.850 744.450 ;
        RECT 178.950 741.900 187.200 742.950 ;
        RECT 188.250 742.650 197.850 743.700 ;
        RECT 178.950 737.850 181.050 741.900 ;
        RECT 188.250 741.000 189.150 742.650 ;
        RECT 198.750 741.750 202.650 743.550 ;
        RECT 203.550 742.950 204.600 744.450 ;
        RECT 205.950 745.650 208.050 745.950 ;
        RECT 205.950 743.850 209.850 745.650 ;
        RECT 216.450 743.250 217.500 746.700 ;
        RECT 219.000 745.800 220.050 748.950 ;
        RECT 221.700 749.400 223.500 755.250 ;
        RECT 227.100 749.400 228.900 755.250 ;
        RECT 232.500 749.400 234.300 755.250 ;
        RECT 242.550 752.400 244.350 755.250 ;
        RECT 245.550 752.400 247.350 755.250 ;
        RECT 248.550 752.400 250.350 755.250 ;
        RECT 221.700 748.500 223.200 749.400 ;
        RECT 221.700 747.300 230.100 748.500 ;
        RECT 228.300 746.700 230.100 747.300 ;
        RECT 233.100 745.800 234.300 749.400 ;
        RECT 246.000 745.950 247.050 752.400 ;
        RECT 262.650 749.400 264.450 755.250 ;
        RECT 265.650 749.400 267.450 755.250 ;
        RECT 268.650 749.400 270.450 755.250 ;
        RECT 274.650 752.400 276.450 755.250 ;
        RECT 277.650 752.400 279.450 755.250 ;
        RECT 280.650 752.400 282.450 755.250 ;
        RECT 219.000 744.900 234.300 745.800 ;
        RECT 203.550 742.050 215.550 742.950 ;
        RECT 182.100 739.200 189.150 741.000 ;
        RECT 190.500 739.950 192.300 741.750 ;
        RECT 198.750 741.450 200.850 741.750 ;
        RECT 202.950 740.550 205.050 740.850 ;
        RECT 211.800 740.550 213.600 741.150 ;
        RECT 202.950 739.950 213.600 740.550 ;
        RECT 190.500 739.350 213.600 739.950 ;
        RECT 214.500 740.550 215.550 742.050 ;
        RECT 216.450 741.450 218.250 743.250 ;
        RECT 220.050 742.950 231.900 744.000 ;
        RECT 220.050 740.550 221.250 742.950 ;
        RECT 230.100 741.150 231.900 742.950 ;
        RECT 214.500 739.650 221.250 740.550 ;
        RECT 223.950 739.650 226.050 739.950 ;
        RECT 190.500 738.750 205.050 739.350 ;
        RECT 222.150 738.450 226.050 739.650 ;
        RECT 229.950 739.050 232.050 741.150 ;
        RECT 212.100 737.850 226.050 738.450 ;
        RECT 186.000 737.550 225.750 737.850 ;
        RECT 174.750 736.650 176.550 737.250 ;
        RECT 186.000 736.650 214.050 737.550 ;
        RECT 174.750 735.450 187.050 736.650 ;
        RECT 214.950 736.050 217.050 736.350 ;
        RECT 224.700 736.050 226.500 736.650 ;
        RECT 187.950 734.550 190.050 735.750 ;
        RECT 172.650 733.650 190.050 734.550 ;
        RECT 193.950 734.400 214.050 735.750 ;
        RECT 193.950 733.650 196.050 734.400 ;
        RECT 175.500 729.600 176.700 733.650 ;
        RECT 177.600 731.700 179.400 732.300 ;
        RECT 184.350 732.150 186.150 732.300 ;
        RECT 177.600 730.500 183.300 731.700 ;
        RECT 184.350 730.950 193.050 732.150 ;
        RECT 184.350 730.500 186.150 730.950 ;
        RECT 165.750 723.750 167.550 729.600 ;
        RECT 168.750 723.750 170.550 729.600 ;
        RECT 172.500 723.750 174.300 729.600 ;
        RECT 175.500 723.750 177.300 729.600 ;
        RECT 178.500 723.750 180.300 729.600 ;
        RECT 181.500 723.750 183.300 730.500 ;
        RECT 190.950 730.050 193.050 730.950 ;
        RECT 184.500 723.750 186.300 729.600 ;
        RECT 187.800 727.800 189.900 729.900 ;
        RECT 188.400 726.600 189.900 727.800 ;
        RECT 188.250 723.750 190.050 726.600 ;
        RECT 191.250 723.750 193.050 730.050 ;
        RECT 194.550 726.600 195.900 733.650 ;
        RECT 212.100 733.350 214.050 734.400 ;
        RECT 214.950 734.850 226.500 736.050 ;
        RECT 214.950 734.250 217.050 734.850 ;
        RECT 228.000 733.350 229.800 734.100 ;
        RECT 197.100 730.800 201.000 732.600 ;
        RECT 198.000 730.500 201.000 730.800 ;
        RECT 202.950 732.150 205.050 732.600 ;
        RECT 212.100 732.300 229.800 733.350 ;
        RECT 202.950 730.500 205.350 732.150 ;
        RECT 194.250 723.750 196.050 726.600 ;
        RECT 198.000 723.750 199.800 730.500 ;
        RECT 204.000 729.600 205.350 730.500 ;
        RECT 211.950 729.600 214.050 730.050 ;
        RECT 201.000 723.750 202.800 729.600 ;
        RECT 204.000 723.750 205.800 729.600 ;
        RECT 207.750 723.750 209.550 729.600 ;
        RECT 211.500 727.950 214.050 729.600 ;
        RECT 214.950 727.950 217.050 730.050 ;
        RECT 217.950 727.950 220.050 730.050 ;
        RECT 211.500 726.600 212.700 727.950 ;
        RECT 214.950 726.600 215.850 727.950 ;
        RECT 217.950 726.600 219.150 727.950 ;
        RECT 210.750 723.750 212.700 726.600 ;
        RECT 213.750 723.750 215.850 726.600 ;
        RECT 216.750 723.750 219.150 726.600 ;
        RECT 220.500 723.750 222.300 727.050 ;
        RECT 223.500 723.750 225.300 732.300 ;
        RECT 233.100 731.400 234.300 744.900 ;
        RECT 244.950 743.850 247.050 745.950 ;
        RECT 265.800 744.150 267.150 749.400 ;
        RECT 277.950 745.950 279.000 752.400 ;
        RECT 280.950 747.450 283.050 748.050 ;
        RECT 280.950 746.550 285.450 747.450 ;
        RECT 280.950 745.950 283.050 746.550 ;
        RECT 269.100 744.150 270.900 745.950 ;
        RECT 241.950 740.850 244.050 742.950 ;
        RECT 242.100 739.050 243.900 740.850 ;
        RECT 246.000 736.650 247.050 743.850 ;
        RECT 247.950 740.850 250.050 742.950 ;
        RECT 262.950 742.050 267.150 744.150 ;
        RECT 268.950 742.050 271.050 744.150 ;
        RECT 277.950 743.850 280.050 745.950 ;
        RECT 248.100 739.050 249.900 740.850 ;
        RECT 246.000 735.600 248.550 736.650 ;
        RECT 265.800 735.600 267.150 742.050 ;
        RECT 274.950 740.850 277.050 742.950 ;
        RECT 275.100 739.050 276.900 740.850 ;
        RECT 277.950 736.650 279.000 743.850 ;
        RECT 280.950 740.850 283.050 742.950 ;
        RECT 281.100 739.050 282.900 740.850 ;
        RECT 284.550 738.450 285.450 746.550 ;
        RECT 290.700 746.400 292.500 755.250 ;
        RECT 296.100 747.000 297.900 755.250 ;
        RECT 305.550 752.400 307.350 755.250 ;
        RECT 308.550 752.400 310.350 755.250 ;
        RECT 311.550 752.400 313.350 755.250 ;
        RECT 320.550 752.400 322.350 755.250 ;
        RECT 323.550 752.400 325.350 755.250 ;
        RECT 326.550 752.400 328.350 755.250 ;
        RECT 296.100 745.350 300.600 747.000 ;
        RECT 309.000 745.950 310.050 752.400 ;
        RECT 324.450 748.200 325.350 752.400 ;
        RECT 329.550 749.400 331.350 755.250 ;
        RECT 337.650 752.400 339.450 755.250 ;
        RECT 340.650 752.400 342.450 755.250 ;
        RECT 343.650 752.400 345.450 755.250 ;
        RECT 347.550 752.400 349.350 755.250 ;
        RECT 350.550 752.400 352.350 755.250 ;
        RECT 324.450 747.300 327.750 748.200 ;
        RECT 325.950 746.400 327.750 747.300 ;
        RECT 299.400 741.150 300.600 745.350 ;
        RECT 307.950 743.850 310.050 745.950 ;
        RECT 319.950 743.850 322.050 745.950 ;
        RECT 286.950 738.450 289.050 739.050 ;
        RECT 284.550 737.550 289.050 738.450 ;
        RECT 289.950 737.850 292.050 739.950 ;
        RECT 295.950 737.850 298.050 739.950 ;
        RECT 298.950 739.050 301.050 741.150 ;
        RECT 304.950 740.850 307.050 742.950 ;
        RECT 305.100 739.050 306.900 740.850 ;
        RECT 286.950 736.950 289.050 737.550 ;
        RECT 276.450 735.600 279.000 736.650 ;
        RECT 290.100 736.050 291.900 737.850 ;
        RECT 230.250 730.500 234.300 731.400 ;
        RECT 230.250 729.600 231.300 730.500 ;
        RECT 226.500 723.750 228.300 729.600 ;
        RECT 229.500 723.750 231.300 729.600 ;
        RECT 232.500 723.750 234.300 729.600 ;
        RECT 242.550 723.750 244.350 735.600 ;
        RECT 246.750 723.750 248.550 735.600 ;
        RECT 262.650 723.750 264.450 735.600 ;
        RECT 265.650 723.750 267.450 735.600 ;
        RECT 268.650 723.750 270.450 735.600 ;
        RECT 276.450 723.750 278.250 735.600 ;
        RECT 280.650 723.750 282.450 735.600 ;
        RECT 292.950 734.850 295.050 736.950 ;
        RECT 296.250 736.050 298.050 737.850 ;
        RECT 293.100 733.050 294.900 734.850 ;
        RECT 299.700 730.800 300.750 739.050 ;
        RECT 309.000 736.650 310.050 743.850 ;
        RECT 310.950 740.850 313.050 742.950 ;
        RECT 320.100 742.050 321.900 743.850 ;
        RECT 322.950 740.850 325.050 742.950 ;
        RECT 311.100 739.050 312.900 740.850 ;
        RECT 323.100 739.050 324.900 740.850 ;
        RECT 326.700 738.150 327.600 746.400 ;
        RECT 330.000 744.150 331.050 749.400 ;
        RECT 328.950 742.050 331.050 744.150 ;
        RECT 340.950 745.950 342.000 752.400 ;
        RECT 340.950 743.850 343.050 745.950 ;
        RECT 346.950 743.850 349.050 745.950 ;
        RECT 350.400 744.150 351.600 752.400 ;
        RECT 362.700 746.400 364.500 755.250 ;
        RECT 368.100 747.000 369.900 755.250 ;
        RECT 385.650 754.500 393.450 755.250 ;
        RECT 385.650 749.400 387.450 754.500 ;
        RECT 388.650 749.400 390.450 753.600 ;
        RECT 391.650 750.000 393.450 754.500 ;
        RECT 394.650 750.900 396.450 755.250 ;
        RECT 397.650 750.000 399.450 755.250 ;
        RECT 389.250 747.900 390.150 749.400 ;
        RECT 391.650 749.100 399.450 750.000 ;
        RECT 368.100 745.350 372.600 747.000 ;
        RECT 389.250 746.850 393.600 747.900 ;
        RECT 407.100 747.000 408.900 755.250 ;
        RECT 325.950 738.000 327.750 738.150 ;
        RECT 320.550 736.800 327.750 738.000 ;
        RECT 309.000 735.600 311.550 736.650 ;
        RECT 293.700 729.900 300.750 730.800 ;
        RECT 293.700 729.600 295.350 729.900 ;
        RECT 290.550 723.750 292.350 729.600 ;
        RECT 293.550 723.750 295.350 729.600 ;
        RECT 299.550 729.600 300.750 729.900 ;
        RECT 296.550 723.750 298.350 729.000 ;
        RECT 299.550 723.750 301.350 729.600 ;
        RECT 305.550 723.750 307.350 735.600 ;
        RECT 309.750 723.750 311.550 735.600 ;
        RECT 320.550 735.600 321.750 736.800 ;
        RECT 325.950 736.350 327.750 736.800 ;
        RECT 320.550 723.750 322.350 735.600 ;
        RECT 329.100 735.450 330.450 742.050 ;
        RECT 337.950 740.850 340.050 742.950 ;
        RECT 338.100 739.050 339.900 740.850 ;
        RECT 340.950 736.650 342.000 743.850 ;
        RECT 343.950 740.850 346.050 742.950 ;
        RECT 347.100 742.050 348.900 743.850 ;
        RECT 349.950 742.050 352.050 744.150 ;
        RECT 344.100 739.050 345.900 740.850 ;
        RECT 325.050 723.750 326.850 735.450 ;
        RECT 328.050 734.100 330.450 735.450 ;
        RECT 339.450 735.600 342.000 736.650 ;
        RECT 328.050 723.750 329.850 734.100 ;
        RECT 339.450 723.750 341.250 735.600 ;
        RECT 343.650 723.750 345.450 735.600 ;
        RECT 350.400 729.600 351.600 742.050 ;
        RECT 371.400 741.150 372.600 745.350 ;
        RECT 389.700 744.150 391.500 745.950 ;
        RECT 361.950 737.850 364.050 739.950 ;
        RECT 367.950 737.850 370.050 739.950 ;
        RECT 370.950 739.050 373.050 741.150 ;
        RECT 385.950 740.850 388.050 742.950 ;
        RECT 388.950 742.050 391.050 744.150 ;
        RECT 392.400 742.950 393.600 746.850 ;
        RECT 395.100 744.150 396.900 745.950 ;
        RECT 404.400 745.350 408.900 747.000 ;
        RECT 412.500 746.400 414.300 755.250 ;
        RECT 417.000 749.400 418.800 755.250 ;
        RECT 421.200 751.050 423.000 755.250 ;
        RECT 424.500 752.400 426.300 755.250 ;
        RECT 421.200 749.400 426.900 751.050 ;
        RECT 436.650 749.400 438.450 755.250 ;
        RECT 439.650 752.400 441.450 755.250 ;
        RECT 442.650 752.400 444.450 755.250 ;
        RECT 445.650 752.400 447.450 755.250 ;
        RECT 391.950 740.850 394.050 742.950 ;
        RECT 394.950 742.050 397.050 744.150 ;
        RECT 397.950 740.850 400.050 742.950 ;
        RECT 404.400 741.150 405.600 745.350 ;
        RECT 416.100 744.150 417.900 745.950 ;
        RECT 415.950 742.050 418.050 744.150 ;
        RECT 418.950 743.850 421.050 745.950 ;
        RECT 422.100 744.150 423.900 745.950 ;
        RECT 419.100 742.050 420.900 743.850 ;
        RECT 421.950 742.050 424.050 744.150 ;
        RECT 425.700 742.950 426.900 749.400 ;
        RECT 436.950 744.150 438.000 749.400 ;
        RECT 442.650 748.200 443.550 752.400 ;
        RECT 454.650 749.400 456.450 755.250 ;
        RECT 440.250 747.300 443.550 748.200 ;
        RECT 455.250 747.300 456.450 749.400 ;
        RECT 457.650 750.300 459.450 755.250 ;
        RECT 460.650 751.200 462.450 755.250 ;
        RECT 463.650 750.300 465.450 755.250 ;
        RECT 467.550 752.400 469.350 755.250 ;
        RECT 470.550 752.400 472.350 755.250 ;
        RECT 457.650 748.950 465.450 750.300 ;
        RECT 440.250 746.400 442.050 747.300 ;
        RECT 386.250 739.050 388.050 740.850 ;
        RECT 362.100 736.050 363.900 737.850 ;
        RECT 364.950 734.850 367.050 736.950 ;
        RECT 368.250 736.050 370.050 737.850 ;
        RECT 365.100 733.050 366.900 734.850 ;
        RECT 371.700 730.800 372.750 739.050 ;
        RECT 392.250 735.600 393.450 740.850 ;
        RECT 398.100 739.050 399.900 740.850 ;
        RECT 403.950 739.050 406.050 741.150 ;
        RECT 424.950 740.850 427.050 742.950 ;
        RECT 436.950 742.050 439.050 744.150 ;
        RECT 365.700 729.900 372.750 730.800 ;
        RECT 365.700 729.600 367.350 729.900 ;
        RECT 347.550 723.750 349.350 729.600 ;
        RECT 350.550 723.750 352.350 729.600 ;
        RECT 362.550 723.750 364.350 729.600 ;
        RECT 365.550 723.750 367.350 729.600 ;
        RECT 371.550 729.600 372.750 729.900 ;
        RECT 368.550 723.750 370.350 729.000 ;
        RECT 371.550 723.750 373.350 729.600 ;
        RECT 387.150 723.750 388.950 735.600 ;
        RECT 391.650 723.750 394.950 735.600 ;
        RECT 397.650 723.750 399.450 735.600 ;
        RECT 404.250 730.800 405.300 739.050 ;
        RECT 406.950 737.850 409.050 739.950 ;
        RECT 412.950 737.850 415.050 739.950 ;
        RECT 406.950 736.050 408.750 737.850 ;
        RECT 409.950 734.850 412.050 736.950 ;
        RECT 413.100 736.050 414.900 737.850 ;
        RECT 425.700 735.600 426.900 740.850 ;
        RECT 410.100 733.050 411.900 734.850 ;
        RECT 416.550 734.700 424.350 735.600 ;
        RECT 404.250 729.900 411.300 730.800 ;
        RECT 404.250 729.600 405.450 729.900 ;
        RECT 403.650 723.750 405.450 729.600 ;
        RECT 409.650 729.600 411.300 729.900 ;
        RECT 406.650 723.750 408.450 729.000 ;
        RECT 409.650 723.750 411.450 729.600 ;
        RECT 412.650 723.750 414.450 729.600 ;
        RECT 416.550 723.750 418.350 734.700 ;
        RECT 419.550 723.750 421.350 733.800 ;
        RECT 422.550 723.750 424.350 734.700 ;
        RECT 425.550 723.750 427.350 735.600 ;
        RECT 437.550 735.450 438.900 742.050 ;
        RECT 440.400 738.150 441.300 746.400 ;
        RECT 455.250 746.250 459.000 747.300 ;
        RECT 445.950 743.850 448.050 745.950 ;
        RECT 442.950 740.850 445.050 742.950 ;
        RECT 446.100 742.050 447.900 743.850 ;
        RECT 457.950 742.950 459.150 746.250 ;
        RECT 461.100 744.150 462.900 745.950 ;
        RECT 457.950 740.850 460.050 742.950 ;
        RECT 460.950 742.050 463.050 744.150 ;
        RECT 466.950 743.850 469.050 745.950 ;
        RECT 470.400 744.150 471.600 752.400 ;
        RECT 482.850 748.200 484.650 755.250 ;
        RECT 487.350 749.400 489.150 755.250 ;
        RECT 497.700 752.400 499.500 755.250 ;
        RECT 501.000 751.050 502.800 755.250 ;
        RECT 497.100 749.400 502.800 751.050 ;
        RECT 505.200 749.400 507.000 755.250 ;
        RECT 512.550 752.400 514.350 755.250 ;
        RECT 515.550 752.400 517.350 755.250 ;
        RECT 518.550 752.400 520.350 755.250 ;
        RECT 532.650 752.400 534.450 755.250 ;
        RECT 535.650 752.400 537.450 755.250 ;
        RECT 482.850 747.300 486.450 748.200 ;
        RECT 463.950 740.850 466.050 742.950 ;
        RECT 467.100 742.050 468.900 743.850 ;
        RECT 469.950 742.050 472.050 744.150 ;
        RECT 443.100 739.050 444.900 740.850 ;
        RECT 440.250 738.000 442.050 738.150 ;
        RECT 440.250 736.800 447.450 738.000 ;
        RECT 454.950 737.850 457.050 739.950 ;
        RECT 440.250 736.350 442.050 736.800 ;
        RECT 446.250 735.600 447.450 736.800 ;
        RECT 455.250 736.050 457.050 737.850 ;
        RECT 458.850 735.600 460.050 740.850 ;
        RECT 464.100 739.050 465.900 740.850 ;
        RECT 437.550 734.100 439.950 735.450 ;
        RECT 438.150 723.750 439.950 734.100 ;
        RECT 441.150 723.750 442.950 735.450 ;
        RECT 445.650 723.750 447.450 735.600 ;
        RECT 455.400 723.750 457.200 729.600 ;
        RECT 458.700 723.750 460.500 735.600 ;
        RECT 462.900 723.750 464.700 735.600 ;
        RECT 470.400 729.600 471.600 742.050 ;
        RECT 482.100 741.150 483.900 742.950 ;
        RECT 481.950 739.050 484.050 741.150 ;
        RECT 485.250 739.950 486.450 747.300 ;
        RECT 497.100 742.950 498.300 749.400 ;
        RECT 516.000 745.950 517.050 752.400 ;
        RECT 500.100 744.150 501.900 745.950 ;
        RECT 488.100 741.150 489.900 742.950 ;
        RECT 484.950 737.850 487.050 739.950 ;
        RECT 487.950 739.050 490.050 741.150 ;
        RECT 496.950 740.850 499.050 742.950 ;
        RECT 499.950 742.050 502.050 744.150 ;
        RECT 502.950 743.850 505.050 745.950 ;
        RECT 506.100 744.150 507.900 745.950 ;
        RECT 503.100 742.050 504.900 743.850 ;
        RECT 505.950 742.050 508.050 744.150 ;
        RECT 514.950 743.850 517.050 745.950 ;
        RECT 533.400 744.150 534.600 752.400 ;
        RECT 539.850 749.400 541.650 755.250 ;
        RECT 544.350 748.200 546.150 755.250 ;
        RECT 542.550 747.300 546.150 748.200 ;
        RECT 560.850 748.200 562.650 755.250 ;
        RECT 565.350 749.400 567.150 755.250 ;
        RECT 575.850 749.400 577.650 755.250 ;
        RECT 580.350 748.200 582.150 755.250 ;
        RECT 589.650 752.400 591.450 755.250 ;
        RECT 592.650 752.400 594.450 755.250 ;
        RECT 598.650 752.400 600.450 755.250 ;
        RECT 601.650 752.400 603.450 755.250 ;
        RECT 604.650 752.400 606.450 755.250 ;
        RECT 560.850 747.300 564.450 748.200 ;
        RECT 511.950 740.850 514.050 742.950 ;
        RECT 485.250 729.600 486.450 737.850 ;
        RECT 497.100 735.600 498.300 740.850 ;
        RECT 512.100 739.050 513.900 740.850 ;
        RECT 516.000 736.650 517.050 743.850 ;
        RECT 517.950 740.850 520.050 742.950 ;
        RECT 532.950 742.050 535.050 744.150 ;
        RECT 535.950 743.850 538.050 745.950 ;
        RECT 536.100 742.050 537.900 743.850 ;
        RECT 518.100 739.050 519.900 740.850 ;
        RECT 516.000 735.600 518.550 736.650 ;
        RECT 467.550 723.750 469.350 729.600 ;
        RECT 470.550 723.750 472.350 729.600 ;
        RECT 481.650 723.750 483.450 729.600 ;
        RECT 484.650 723.750 486.450 729.600 ;
        RECT 487.650 723.750 489.450 729.600 ;
        RECT 496.650 723.750 498.450 735.600 ;
        RECT 499.650 734.700 507.450 735.600 ;
        RECT 499.650 723.750 501.450 734.700 ;
        RECT 502.650 723.750 504.450 733.800 ;
        RECT 505.650 723.750 507.450 734.700 ;
        RECT 512.550 723.750 514.350 735.600 ;
        RECT 516.750 723.750 518.550 735.600 ;
        RECT 533.400 729.600 534.600 742.050 ;
        RECT 539.100 741.150 540.900 742.950 ;
        RECT 538.950 739.050 541.050 741.150 ;
        RECT 542.550 739.950 543.750 747.300 ;
        RECT 545.100 741.150 546.900 742.950 ;
        RECT 560.100 741.150 561.900 742.950 ;
        RECT 541.950 737.850 544.050 739.950 ;
        RECT 544.950 739.050 547.050 741.150 ;
        RECT 559.950 739.050 562.050 741.150 ;
        RECT 563.250 739.950 564.450 747.300 ;
        RECT 578.550 747.300 582.150 748.200 ;
        RECT 566.100 741.150 567.900 742.950 ;
        RECT 575.100 741.150 576.900 742.950 ;
        RECT 562.950 737.850 565.050 739.950 ;
        RECT 565.950 739.050 568.050 741.150 ;
        RECT 574.950 739.050 577.050 741.150 ;
        RECT 578.550 739.950 579.750 747.300 ;
        RECT 590.400 744.150 591.600 752.400 ;
        RECT 601.950 745.950 603.000 752.400 ;
        RECT 608.550 750.300 610.350 755.250 ;
        RECT 611.550 751.200 613.350 755.250 ;
        RECT 614.550 750.300 616.350 755.250 ;
        RECT 608.550 748.950 616.350 750.300 ;
        RECT 617.550 749.400 619.350 755.250 ;
        RECT 617.550 747.300 618.750 749.400 ;
        RECT 632.850 748.200 634.650 755.250 ;
        RECT 637.350 749.400 639.150 755.250 ;
        RECT 644.550 752.400 646.350 755.250 ;
        RECT 647.550 752.400 649.350 755.250 ;
        RECT 632.850 747.300 636.450 748.200 ;
        RECT 615.000 746.250 618.750 747.300 ;
        RECT 581.100 741.150 582.900 742.950 ;
        RECT 589.950 742.050 592.050 744.150 ;
        RECT 592.950 743.850 595.050 745.950 ;
        RECT 601.950 743.850 604.050 745.950 ;
        RECT 611.100 744.150 612.900 745.950 ;
        RECT 593.100 742.050 594.900 743.850 ;
        RECT 577.950 737.850 580.050 739.950 ;
        RECT 580.950 739.050 583.050 741.150 ;
        RECT 542.550 729.600 543.750 737.850 ;
        RECT 563.250 729.600 564.450 737.850 ;
        RECT 578.550 729.600 579.750 737.850 ;
        RECT 590.400 729.600 591.600 742.050 ;
        RECT 598.950 740.850 601.050 742.950 ;
        RECT 599.100 739.050 600.900 740.850 ;
        RECT 601.950 736.650 603.000 743.850 ;
        RECT 604.950 740.850 607.050 742.950 ;
        RECT 607.950 740.850 610.050 742.950 ;
        RECT 610.950 742.050 613.050 744.150 ;
        RECT 614.850 742.950 616.050 746.250 ;
        RECT 613.950 740.850 616.050 742.950 ;
        RECT 632.100 741.150 633.900 742.950 ;
        RECT 605.100 739.050 606.900 740.850 ;
        RECT 608.100 739.050 609.900 740.850 ;
        RECT 600.450 735.600 603.000 736.650 ;
        RECT 613.950 735.600 615.150 740.850 ;
        RECT 616.950 737.850 619.050 739.950 ;
        RECT 631.950 739.050 634.050 741.150 ;
        RECT 635.250 739.950 636.450 747.300 ;
        RECT 643.950 743.850 646.050 745.950 ;
        RECT 647.400 744.150 648.600 752.400 ;
        RECT 659.700 746.400 661.500 755.250 ;
        RECT 665.100 747.000 666.900 755.250 ;
        RECT 677.850 749.400 679.650 755.250 ;
        RECT 682.350 748.200 684.150 755.250 ;
        RECT 680.550 747.300 684.150 748.200 ;
        RECT 689.550 747.900 691.350 755.250 ;
        RECT 694.050 749.400 695.850 755.250 ;
        RECT 697.050 750.900 698.850 755.250 ;
        RECT 710.550 752.400 712.350 755.250 ;
        RECT 713.550 752.400 715.350 755.250 ;
        RECT 697.050 749.400 700.350 750.900 ;
        RECT 695.250 747.900 697.050 748.500 ;
        RECT 665.100 745.350 669.600 747.000 ;
        RECT 649.950 744.450 652.050 745.050 ;
        RECT 658.950 744.450 661.050 745.050 ;
        RECT 638.100 741.150 639.900 742.950 ;
        RECT 644.100 742.050 645.900 743.850 ;
        RECT 646.950 742.050 649.050 744.150 ;
        RECT 649.950 743.550 661.050 744.450 ;
        RECT 649.950 742.950 652.050 743.550 ;
        RECT 658.950 742.950 661.050 743.550 ;
        RECT 634.950 737.850 637.050 739.950 ;
        RECT 637.950 739.050 640.050 741.150 ;
        RECT 616.950 736.050 618.750 737.850 ;
        RECT 532.650 723.750 534.450 729.600 ;
        RECT 535.650 723.750 537.450 729.600 ;
        RECT 539.550 723.750 541.350 729.600 ;
        RECT 542.550 723.750 544.350 729.600 ;
        RECT 545.550 723.750 547.350 729.600 ;
        RECT 559.650 723.750 561.450 729.600 ;
        RECT 562.650 723.750 564.450 729.600 ;
        RECT 565.650 723.750 567.450 729.600 ;
        RECT 575.550 723.750 577.350 729.600 ;
        RECT 578.550 723.750 580.350 729.600 ;
        RECT 581.550 723.750 583.350 729.600 ;
        RECT 589.650 723.750 591.450 729.600 ;
        RECT 592.650 723.750 594.450 729.600 ;
        RECT 600.450 723.750 602.250 735.600 ;
        RECT 604.650 723.750 606.450 735.600 ;
        RECT 609.300 723.750 611.100 735.600 ;
        RECT 613.500 723.750 615.300 735.600 ;
        RECT 635.250 729.600 636.450 737.850 ;
        RECT 647.400 729.600 648.600 742.050 ;
        RECT 668.400 741.150 669.600 745.350 ;
        RECT 677.100 741.150 678.900 742.950 ;
        RECT 658.950 737.850 661.050 739.950 ;
        RECT 664.950 737.850 667.050 739.950 ;
        RECT 667.950 739.050 670.050 741.150 ;
        RECT 676.950 739.050 679.050 741.150 ;
        RECT 680.550 739.950 681.750 747.300 ;
        RECT 689.550 746.700 697.050 747.900 ;
        RECT 683.100 741.150 684.900 742.950 ;
        RECT 659.100 736.050 660.900 737.850 ;
        RECT 661.950 734.850 664.050 736.950 ;
        RECT 665.250 736.050 667.050 737.850 ;
        RECT 662.100 733.050 663.900 734.850 ;
        RECT 668.700 730.800 669.750 739.050 ;
        RECT 679.950 737.850 682.050 739.950 ;
        RECT 682.950 739.050 685.050 741.150 ;
        RECT 688.950 740.850 691.050 742.950 ;
        RECT 689.100 739.050 690.900 740.850 ;
        RECT 662.700 729.900 669.750 730.800 ;
        RECT 662.700 729.600 664.350 729.900 ;
        RECT 616.800 723.750 618.600 729.600 ;
        RECT 631.650 723.750 633.450 729.600 ;
        RECT 634.650 723.750 636.450 729.600 ;
        RECT 637.650 723.750 639.450 729.600 ;
        RECT 644.550 723.750 646.350 729.600 ;
        RECT 647.550 723.750 649.350 729.600 ;
        RECT 659.550 723.750 661.350 729.600 ;
        RECT 662.550 723.750 664.350 729.600 ;
        RECT 668.550 729.600 669.750 729.900 ;
        RECT 680.550 729.600 681.750 737.850 ;
        RECT 692.700 729.600 693.900 746.700 ;
        RECT 699.150 742.950 700.350 749.400 ;
        RECT 709.950 743.850 712.050 745.950 ;
        RECT 713.400 744.150 714.600 752.400 ;
        RECT 727.650 749.400 729.450 755.250 ;
        RECT 730.650 752.400 732.450 755.250 ;
        RECT 733.650 752.400 735.450 755.250 ;
        RECT 736.650 752.400 738.450 755.250 ;
        RECT 727.950 744.150 729.000 749.400 ;
        RECT 733.650 748.200 734.550 752.400 ;
        RECT 746.550 750.300 748.350 755.250 ;
        RECT 749.550 751.200 751.350 755.250 ;
        RECT 752.550 750.300 754.350 755.250 ;
        RECT 746.550 748.950 754.350 750.300 ;
        RECT 755.550 749.400 757.350 755.250 ;
        RECT 761.550 752.400 763.350 755.250 ;
        RECT 764.550 752.400 766.350 755.250 ;
        RECT 767.550 752.400 769.350 755.250 ;
        RECT 774.750 752.400 776.550 755.250 ;
        RECT 777.750 752.400 779.550 755.250 ;
        RECT 731.250 747.300 734.550 748.200 ;
        RECT 755.550 747.300 756.750 749.400 ;
        RECT 731.250 746.400 733.050 747.300 ;
        RECT 695.100 741.150 696.900 742.950 ;
        RECT 694.950 739.050 697.050 741.150 ;
        RECT 697.950 740.850 700.350 742.950 ;
        RECT 710.100 742.050 711.900 743.850 ;
        RECT 712.950 742.050 715.050 744.150 ;
        RECT 727.950 742.050 730.050 744.150 ;
        RECT 699.150 735.600 700.350 740.850 ;
        RECT 665.550 723.750 667.350 729.000 ;
        RECT 668.550 723.750 670.350 729.600 ;
        RECT 677.550 723.750 679.350 729.600 ;
        RECT 680.550 723.750 682.350 729.600 ;
        RECT 683.550 723.750 685.350 729.600 ;
        RECT 689.550 723.750 691.350 729.600 ;
        RECT 692.550 723.750 694.350 729.600 ;
        RECT 696.150 723.750 697.950 735.600 ;
        RECT 699.150 723.750 700.950 735.600 ;
        RECT 713.400 729.600 714.600 742.050 ;
        RECT 728.550 735.450 729.900 742.050 ;
        RECT 731.400 738.150 732.300 746.400 ;
        RECT 753.000 746.250 756.750 747.300 ;
        RECT 736.950 743.850 739.050 745.950 ;
        RECT 749.100 744.150 750.900 745.950 ;
        RECT 733.950 740.850 736.050 742.950 ;
        RECT 737.100 742.050 738.900 743.850 ;
        RECT 745.950 740.850 748.050 742.950 ;
        RECT 748.950 742.050 751.050 744.150 ;
        RECT 752.850 742.950 754.050 746.250 ;
        RECT 765.000 745.950 766.050 752.400 ;
        RECT 763.950 743.850 766.050 745.950 ;
        RECT 778.050 744.150 779.550 752.400 ;
        RECT 751.950 740.850 754.050 742.950 ;
        RECT 760.950 740.850 763.050 742.950 ;
        RECT 734.100 739.050 735.900 740.850 ;
        RECT 746.100 739.050 747.900 740.850 ;
        RECT 731.250 738.000 733.050 738.150 ;
        RECT 731.250 736.800 738.450 738.000 ;
        RECT 731.250 736.350 733.050 736.800 ;
        RECT 737.250 735.600 738.450 736.800 ;
        RECT 751.950 735.600 753.150 740.850 ;
        RECT 754.950 737.850 757.050 739.950 ;
        RECT 761.100 739.050 762.900 740.850 ;
        RECT 754.950 736.050 756.750 737.850 ;
        RECT 765.000 736.650 766.050 743.850 ;
        RECT 766.950 740.850 769.050 742.950 ;
        RECT 775.950 742.050 779.550 744.150 ;
        RECT 767.100 739.050 768.900 740.850 ;
        RECT 765.000 735.600 767.550 736.650 ;
        RECT 728.550 734.100 730.950 735.450 ;
        RECT 710.550 723.750 712.350 729.600 ;
        RECT 713.550 723.750 715.350 729.600 ;
        RECT 729.150 723.750 730.950 734.100 ;
        RECT 732.150 723.750 733.950 735.450 ;
        RECT 736.650 723.750 738.450 735.600 ;
        RECT 747.300 723.750 749.100 735.600 ;
        RECT 751.500 723.750 753.300 735.600 ;
        RECT 754.800 723.750 756.600 729.600 ;
        RECT 761.550 723.750 763.350 735.600 ;
        RECT 765.750 723.750 767.550 735.600 ;
        RECT 778.050 729.600 779.550 742.050 ;
        RECT 781.650 749.400 783.450 755.250 ;
        RECT 787.050 749.400 788.850 755.250 ;
        RECT 792.600 750.600 794.400 755.250 ;
        RECT 797.250 751.500 799.050 755.250 ;
        RECT 800.250 751.500 802.050 755.250 ;
        RECT 803.250 751.500 805.050 755.250 ;
        RECT 790.200 749.400 794.400 750.600 ;
        RECT 796.950 749.400 799.050 751.500 ;
        RECT 799.950 749.400 802.050 751.500 ;
        RECT 802.950 749.400 805.050 751.500 ;
        RECT 807.000 751.500 808.800 755.250 ;
        RECT 810.000 752.400 811.800 755.250 ;
        RECT 813.000 751.500 814.800 755.250 ;
        RECT 817.500 752.400 819.300 755.250 ;
        RECT 820.500 752.400 822.300 755.250 ;
        RECT 823.500 752.400 825.300 755.250 ;
        RECT 826.500 752.400 828.300 755.250 ;
        RECT 807.000 749.700 809.850 751.500 ;
        RECT 807.750 749.400 809.850 749.700 ;
        RECT 811.950 749.700 814.800 751.500 ;
        RECT 815.700 750.750 817.500 751.200 ;
        RECT 820.950 751.050 822.300 752.400 ;
        RECT 823.950 751.050 825.300 752.400 ;
        RECT 826.950 751.050 828.300 752.400 ;
        RECT 811.950 749.400 814.050 749.700 ;
        RECT 815.700 749.400 819.750 750.750 ;
        RECT 781.650 734.550 782.850 749.400 ;
        RECT 790.200 745.800 791.700 749.400 ;
        RECT 796.350 746.700 803.100 748.500 ;
        RECT 804.000 746.700 810.900 748.500 ;
        RECT 818.850 748.050 819.750 749.400 ;
        RECT 820.950 748.950 823.050 751.050 ;
        RECT 823.950 748.950 826.050 751.050 ;
        RECT 826.950 748.950 829.050 751.050 ;
        RECT 818.850 747.900 823.950 748.050 ;
        RECT 818.850 747.150 826.500 747.900 ;
        RECT 822.150 746.700 826.500 747.150 ;
        RECT 804.000 745.800 805.050 746.700 ;
        RECT 822.150 746.250 823.950 746.700 ;
        RECT 783.900 744.000 791.700 745.800 ;
        RECT 795.150 744.750 805.050 745.800 ;
        RECT 795.150 742.950 796.200 744.750 ;
        RECT 805.950 744.450 813.600 745.800 ;
        RECT 805.950 743.700 806.850 744.450 ;
        RECT 787.950 741.900 796.200 742.950 ;
        RECT 797.250 742.650 806.850 743.700 ;
        RECT 787.950 737.850 790.050 741.900 ;
        RECT 797.250 741.000 798.150 742.650 ;
        RECT 807.750 741.750 811.650 743.550 ;
        RECT 812.550 742.950 813.600 744.450 ;
        RECT 814.950 745.650 817.050 745.950 ;
        RECT 814.950 743.850 818.850 745.650 ;
        RECT 825.450 743.250 826.500 746.700 ;
        RECT 828.000 745.800 829.050 748.950 ;
        RECT 830.700 749.400 832.500 755.250 ;
        RECT 836.100 749.400 837.900 755.250 ;
        RECT 841.500 749.400 843.300 755.250 ;
        RECT 830.700 748.500 832.200 749.400 ;
        RECT 830.700 747.300 839.100 748.500 ;
        RECT 837.300 746.700 839.100 747.300 ;
        RECT 842.100 745.800 843.300 749.400 ;
        RECT 845.550 750.300 847.350 755.250 ;
        RECT 848.550 751.200 850.350 755.250 ;
        RECT 851.550 750.300 853.350 755.250 ;
        RECT 845.550 748.950 853.350 750.300 ;
        RECT 854.550 749.400 856.350 755.250 ;
        RECT 854.550 747.300 855.750 749.400 ;
        RECT 852.000 746.250 855.750 747.300 ;
        RECT 828.000 744.900 843.300 745.800 ;
        RECT 812.550 742.050 824.550 742.950 ;
        RECT 791.100 739.200 798.150 741.000 ;
        RECT 799.500 739.950 801.300 741.750 ;
        RECT 807.750 741.450 809.850 741.750 ;
        RECT 811.950 740.550 814.050 740.850 ;
        RECT 820.800 740.550 822.600 741.150 ;
        RECT 811.950 739.950 822.600 740.550 ;
        RECT 799.500 739.350 822.600 739.950 ;
        RECT 823.500 740.550 824.550 742.050 ;
        RECT 825.450 741.450 827.250 743.250 ;
        RECT 829.050 742.950 840.900 744.000 ;
        RECT 829.050 740.550 830.250 742.950 ;
        RECT 839.100 741.150 840.900 742.950 ;
        RECT 823.500 739.650 830.250 740.550 ;
        RECT 832.950 739.650 835.050 739.950 ;
        RECT 799.500 738.750 814.050 739.350 ;
        RECT 831.150 738.450 835.050 739.650 ;
        RECT 838.950 739.050 841.050 741.150 ;
        RECT 821.100 737.850 835.050 738.450 ;
        RECT 795.000 737.550 834.750 737.850 ;
        RECT 783.750 736.650 785.550 737.250 ;
        RECT 795.000 736.650 823.050 737.550 ;
        RECT 783.750 735.450 796.050 736.650 ;
        RECT 823.950 736.050 826.050 736.350 ;
        RECT 833.700 736.050 835.500 736.650 ;
        RECT 796.950 734.550 799.050 735.750 ;
        RECT 781.650 733.650 799.050 734.550 ;
        RECT 802.950 734.400 823.050 735.750 ;
        RECT 802.950 733.650 805.050 734.400 ;
        RECT 784.500 729.600 785.700 733.650 ;
        RECT 786.600 731.700 788.400 732.300 ;
        RECT 793.350 732.150 795.150 732.300 ;
        RECT 786.600 730.500 792.300 731.700 ;
        RECT 793.350 730.950 802.050 732.150 ;
        RECT 793.350 730.500 795.150 730.950 ;
        RECT 774.750 723.750 776.550 729.600 ;
        RECT 777.750 723.750 779.550 729.600 ;
        RECT 781.500 723.750 783.300 729.600 ;
        RECT 784.500 723.750 786.300 729.600 ;
        RECT 787.500 723.750 789.300 729.600 ;
        RECT 790.500 723.750 792.300 730.500 ;
        RECT 799.950 730.050 802.050 730.950 ;
        RECT 793.500 723.750 795.300 729.600 ;
        RECT 796.800 727.800 798.900 729.900 ;
        RECT 797.400 726.600 798.900 727.800 ;
        RECT 797.250 723.750 799.050 726.600 ;
        RECT 800.250 723.750 802.050 730.050 ;
        RECT 803.550 726.600 804.900 733.650 ;
        RECT 821.100 733.350 823.050 734.400 ;
        RECT 823.950 734.850 835.500 736.050 ;
        RECT 823.950 734.250 826.050 734.850 ;
        RECT 837.000 733.350 838.800 734.100 ;
        RECT 806.100 730.800 810.000 732.600 ;
        RECT 807.000 730.500 810.000 730.800 ;
        RECT 811.950 732.150 814.050 732.600 ;
        RECT 821.100 732.300 838.800 733.350 ;
        RECT 811.950 730.500 814.350 732.150 ;
        RECT 803.250 723.750 805.050 726.600 ;
        RECT 807.000 723.750 808.800 730.500 ;
        RECT 813.000 729.600 814.350 730.500 ;
        RECT 820.950 729.600 823.050 730.050 ;
        RECT 810.000 723.750 811.800 729.600 ;
        RECT 813.000 723.750 814.800 729.600 ;
        RECT 816.750 723.750 818.550 729.600 ;
        RECT 820.500 727.950 823.050 729.600 ;
        RECT 823.950 727.950 826.050 730.050 ;
        RECT 826.950 727.950 829.050 730.050 ;
        RECT 820.500 726.600 821.700 727.950 ;
        RECT 823.950 726.600 824.850 727.950 ;
        RECT 826.950 726.600 828.150 727.950 ;
        RECT 819.750 723.750 821.700 726.600 ;
        RECT 822.750 723.750 824.850 726.600 ;
        RECT 825.750 723.750 828.150 726.600 ;
        RECT 829.500 723.750 831.300 727.050 ;
        RECT 832.500 723.750 834.300 732.300 ;
        RECT 842.100 731.400 843.300 744.900 ;
        RECT 848.100 744.150 849.900 745.950 ;
        RECT 844.950 740.850 847.050 742.950 ;
        RECT 847.950 742.050 850.050 744.150 ;
        RECT 851.850 742.950 853.050 746.250 ;
        RECT 850.950 740.850 853.050 742.950 ;
        RECT 845.100 739.050 846.900 740.850 ;
        RECT 850.950 735.600 852.150 740.850 ;
        RECT 853.950 737.850 856.050 739.950 ;
        RECT 853.950 736.050 855.750 737.850 ;
        RECT 839.250 730.500 843.300 731.400 ;
        RECT 839.250 729.600 840.300 730.500 ;
        RECT 835.500 723.750 837.300 729.600 ;
        RECT 838.500 723.750 840.300 729.600 ;
        RECT 841.500 723.750 843.300 729.600 ;
        RECT 846.300 723.750 848.100 735.600 ;
        RECT 850.500 723.750 852.300 735.600 ;
        RECT 853.800 723.750 855.600 729.600 ;
        RECT 7.650 713.400 9.450 719.250 ;
        RECT 10.650 713.400 12.450 719.250 ;
        RECT 13.650 713.400 15.450 719.250 ;
        RECT 11.250 705.150 12.450 713.400 ;
        RECT 20.550 707.400 22.350 719.250 ;
        RECT 24.750 707.400 26.550 719.250 ;
        RECT 32.700 713.400 34.500 719.250 ;
        RECT 35.700 713.400 37.500 719.250 ;
        RECT 38.700 713.400 40.500 719.250 ;
        RECT 35.700 712.500 36.750 713.400 ;
        RECT 24.000 706.350 26.550 707.400 ;
        RECT 32.700 711.600 36.750 712.500 ;
        RECT 7.950 701.850 10.050 703.950 ;
        RECT 10.950 703.050 13.050 705.150 ;
        RECT 8.100 700.050 9.900 701.850 ;
        RECT 11.250 695.700 12.450 703.050 ;
        RECT 13.950 701.850 16.050 703.950 ;
        RECT 20.100 702.150 21.900 703.950 ;
        RECT 14.100 700.050 15.900 701.850 ;
        RECT 19.950 700.050 22.050 702.150 ;
        RECT 24.000 699.150 25.050 706.350 ;
        RECT 26.100 702.150 27.900 703.950 ;
        RECT 25.950 700.050 28.050 702.150 ;
        RECT 22.950 697.050 25.050 699.150 ;
        RECT 8.850 694.800 12.450 695.700 ;
        RECT 8.850 687.750 10.650 694.800 ;
        RECT 13.350 687.750 15.150 693.600 ;
        RECT 24.000 690.600 25.050 697.050 ;
        RECT 32.700 698.100 33.900 711.600 ;
        RECT 41.700 710.700 43.500 719.250 ;
        RECT 44.700 715.950 46.500 719.250 ;
        RECT 47.850 716.400 50.250 719.250 ;
        RECT 51.150 716.400 53.250 719.250 ;
        RECT 54.300 716.400 56.250 719.250 ;
        RECT 47.850 715.050 49.050 716.400 ;
        RECT 51.150 715.050 52.050 716.400 ;
        RECT 54.300 715.050 55.500 716.400 ;
        RECT 46.950 712.950 49.050 715.050 ;
        RECT 49.950 712.950 52.050 715.050 ;
        RECT 52.950 713.400 55.500 715.050 ;
        RECT 57.450 713.400 59.250 719.250 ;
        RECT 61.200 713.400 63.000 719.250 ;
        RECT 64.200 713.400 66.000 719.250 ;
        RECT 52.950 712.950 55.050 713.400 ;
        RECT 61.650 712.500 63.000 713.400 ;
        RECT 67.200 712.500 69.000 719.250 ;
        RECT 70.950 716.400 72.750 719.250 ;
        RECT 61.650 710.850 64.050 712.500 ;
        RECT 37.200 709.650 54.900 710.700 ;
        RECT 61.950 710.400 64.050 710.850 ;
        RECT 66.000 712.200 69.000 712.500 ;
        RECT 66.000 710.400 69.900 712.200 ;
        RECT 37.200 708.900 39.000 709.650 ;
        RECT 49.950 708.150 52.050 708.750 ;
        RECT 40.500 706.950 52.050 708.150 ;
        RECT 52.950 708.600 54.900 709.650 ;
        RECT 71.100 709.350 72.450 716.400 ;
        RECT 73.950 712.950 75.750 719.250 ;
        RECT 76.950 716.400 78.750 719.250 ;
        RECT 77.100 715.200 78.600 716.400 ;
        RECT 77.100 713.100 79.200 715.200 ;
        RECT 80.700 713.400 82.500 719.250 ;
        RECT 73.950 712.050 76.050 712.950 ;
        RECT 83.700 712.500 85.500 719.250 ;
        RECT 86.700 713.400 88.500 719.250 ;
        RECT 89.700 713.400 91.500 719.250 ;
        RECT 92.700 713.400 94.500 719.250 ;
        RECT 96.450 713.400 98.250 719.250 ;
        RECT 99.450 713.400 101.250 719.250 ;
        RECT 109.650 713.400 111.450 719.250 ;
        RECT 112.650 713.400 114.450 719.250 ;
        RECT 121.650 713.400 123.450 719.250 ;
        RECT 124.650 714.000 126.450 719.250 ;
        RECT 80.850 712.050 82.650 712.500 ;
        RECT 73.950 710.850 82.650 712.050 ;
        RECT 83.700 711.300 89.400 712.500 ;
        RECT 80.850 710.700 82.650 710.850 ;
        RECT 87.600 710.700 89.400 711.300 ;
        RECT 90.300 709.350 91.500 713.400 ;
        RECT 70.950 708.600 73.050 709.350 ;
        RECT 52.950 707.250 73.050 708.600 ;
        RECT 76.950 708.450 94.350 709.350 ;
        RECT 76.950 707.250 79.050 708.450 ;
        RECT 40.500 706.350 42.300 706.950 ;
        RECT 49.950 706.650 52.050 706.950 ;
        RECT 79.950 706.350 92.250 707.550 ;
        RECT 52.950 705.450 81.000 706.350 ;
        RECT 90.450 705.750 92.250 706.350 ;
        RECT 41.250 705.150 81.000 705.450 ;
        RECT 40.950 704.550 54.900 705.150 ;
        RECT 34.950 701.850 37.050 703.950 ;
        RECT 40.950 703.350 44.850 704.550 ;
        RECT 61.950 703.650 76.500 704.250 ;
        RECT 40.950 703.050 43.050 703.350 ;
        RECT 45.750 702.450 52.500 703.350 ;
        RECT 35.100 700.050 36.900 701.850 ;
        RECT 45.750 700.050 46.950 702.450 ;
        RECT 35.100 699.000 46.950 700.050 ;
        RECT 48.750 699.750 50.550 701.550 ;
        RECT 51.450 700.950 52.500 702.450 ;
        RECT 53.400 703.050 76.500 703.650 ;
        RECT 53.400 702.450 64.050 703.050 ;
        RECT 53.400 701.850 55.200 702.450 ;
        RECT 61.950 702.150 64.050 702.450 ;
        RECT 66.150 701.250 68.250 701.550 ;
        RECT 74.700 701.250 76.500 703.050 ;
        RECT 77.850 702.000 84.900 703.800 ;
        RECT 51.450 700.050 63.450 700.950 ;
        RECT 32.700 697.200 48.000 698.100 ;
        RECT 32.700 693.600 33.900 697.200 ;
        RECT 36.900 695.700 38.700 696.300 ;
        RECT 36.900 694.500 45.300 695.700 ;
        RECT 43.800 693.600 45.300 694.500 ;
        RECT 20.550 687.750 22.350 690.600 ;
        RECT 23.550 687.750 25.350 690.600 ;
        RECT 26.550 687.750 28.350 690.600 ;
        RECT 32.700 687.750 34.500 693.600 ;
        RECT 38.100 687.750 39.900 693.600 ;
        RECT 43.500 687.750 45.300 693.600 ;
        RECT 46.950 694.050 48.000 697.200 ;
        RECT 49.500 696.300 50.550 699.750 ;
        RECT 57.150 697.350 61.050 699.150 ;
        RECT 58.950 697.050 61.050 697.350 ;
        RECT 62.400 698.550 63.450 700.050 ;
        RECT 64.350 699.450 68.250 701.250 ;
        RECT 77.850 700.350 78.750 702.000 ;
        RECT 85.950 701.100 88.050 705.150 ;
        RECT 69.150 699.300 78.750 700.350 ;
        RECT 79.800 700.050 88.050 701.100 ;
        RECT 69.150 698.550 70.050 699.300 ;
        RECT 62.400 697.200 70.050 698.550 ;
        RECT 79.800 698.250 80.850 700.050 ;
        RECT 70.950 697.200 80.850 698.250 ;
        RECT 84.300 697.200 92.100 699.000 ;
        RECT 52.050 696.300 53.850 696.750 ;
        RECT 70.950 696.300 72.000 697.200 ;
        RECT 49.500 695.850 53.850 696.300 ;
        RECT 49.500 695.100 57.150 695.850 ;
        RECT 52.050 694.950 57.150 695.100 ;
        RECT 46.950 691.950 49.050 694.050 ;
        RECT 49.950 691.950 52.050 694.050 ;
        RECT 52.950 691.950 55.050 694.050 ;
        RECT 56.250 693.600 57.150 694.950 ;
        RECT 65.100 694.500 72.000 696.300 ;
        RECT 72.900 694.500 79.650 696.300 ;
        RECT 84.300 693.600 85.800 697.200 ;
        RECT 93.150 693.600 94.350 708.450 ;
        RECT 56.250 692.250 60.300 693.600 ;
        RECT 61.950 693.300 64.050 693.600 ;
        RECT 47.700 690.600 49.050 691.950 ;
        RECT 50.700 690.600 52.050 691.950 ;
        RECT 53.700 690.600 55.050 691.950 ;
        RECT 58.500 691.800 60.300 692.250 ;
        RECT 61.200 691.500 64.050 693.300 ;
        RECT 66.150 693.300 68.250 693.600 ;
        RECT 66.150 691.500 69.000 693.300 ;
        RECT 47.700 687.750 49.500 690.600 ;
        RECT 50.700 687.750 52.500 690.600 ;
        RECT 53.700 687.750 55.500 690.600 ;
        RECT 56.700 687.750 58.500 690.600 ;
        RECT 61.200 687.750 63.000 691.500 ;
        RECT 64.200 687.750 66.000 690.600 ;
        RECT 67.200 687.750 69.000 691.500 ;
        RECT 70.950 691.500 73.050 693.600 ;
        RECT 73.950 691.500 76.050 693.600 ;
        RECT 76.950 691.500 79.050 693.600 ;
        RECT 81.600 692.400 85.800 693.600 ;
        RECT 70.950 687.750 72.750 691.500 ;
        RECT 73.950 687.750 75.750 691.500 ;
        RECT 76.950 687.750 78.750 691.500 ;
        RECT 81.600 687.750 83.400 692.400 ;
        RECT 87.150 687.750 88.950 693.600 ;
        RECT 92.550 687.750 94.350 693.600 ;
        RECT 96.450 700.950 97.950 713.400 ;
        RECT 110.400 700.950 111.600 713.400 ;
        RECT 122.250 713.100 123.450 713.400 ;
        RECT 127.650 713.400 129.450 719.250 ;
        RECT 130.650 713.400 132.450 719.250 ;
        RECT 137.550 713.400 139.350 719.250 ;
        RECT 140.550 713.400 142.350 719.250 ;
        RECT 127.650 713.100 129.300 713.400 ;
        RECT 122.250 712.200 129.300 713.100 ;
        RECT 122.250 703.950 123.300 712.200 ;
        RECT 128.100 708.150 129.900 709.950 ;
        RECT 124.950 705.150 126.750 706.950 ;
        RECT 127.950 706.050 130.050 708.150 ;
        RECT 131.100 705.150 132.900 706.950 ;
        RECT 121.950 701.850 124.050 703.950 ;
        RECT 124.950 703.050 127.050 705.150 ;
        RECT 130.950 703.050 133.050 705.150 ;
        RECT 137.100 702.150 138.900 703.950 ;
        RECT 96.450 698.850 100.050 700.950 ;
        RECT 109.950 698.850 112.050 700.950 ;
        RECT 113.100 699.150 114.900 700.950 ;
        RECT 96.450 690.600 97.950 698.850 ;
        RECT 110.400 690.600 111.600 698.850 ;
        RECT 112.950 697.050 115.050 699.150 ;
        RECT 122.400 697.650 123.600 701.850 ;
        RECT 136.950 700.050 139.050 702.150 ;
        RECT 122.400 696.000 126.900 697.650 ;
        RECT 96.450 687.750 98.250 690.600 ;
        RECT 99.450 687.750 101.250 690.600 ;
        RECT 109.650 687.750 111.450 690.600 ;
        RECT 112.650 687.750 114.450 690.600 ;
        RECT 125.100 687.750 126.900 696.000 ;
        RECT 130.500 687.750 132.300 696.600 ;
        RECT 140.700 696.300 141.900 713.400 ;
        RECT 144.150 707.400 145.950 719.250 ;
        RECT 147.150 707.400 148.950 719.250 ;
        RECT 157.650 713.400 159.450 719.250 ;
        RECT 160.650 714.000 162.450 719.250 ;
        RECT 158.250 713.100 159.450 713.400 ;
        RECT 163.650 713.400 165.450 719.250 ;
        RECT 166.650 713.400 168.450 719.250 ;
        RECT 163.650 713.100 165.300 713.400 ;
        RECT 158.250 712.200 165.300 713.100 ;
        RECT 142.950 701.850 145.050 703.950 ;
        RECT 147.150 702.150 148.350 707.400 ;
        RECT 158.250 703.950 159.300 712.200 ;
        RECT 164.100 708.150 165.900 709.950 ;
        RECT 160.950 705.150 162.750 706.950 ;
        RECT 163.950 706.050 166.050 708.150 ;
        RECT 175.050 707.400 176.850 719.250 ;
        RECT 178.050 707.400 179.850 719.250 ;
        RECT 181.650 713.400 183.450 719.250 ;
        RECT 184.650 713.400 186.450 719.250 ;
        RECT 167.100 705.150 168.900 706.950 ;
        RECT 143.100 700.050 144.900 701.850 ;
        RECT 145.950 700.050 148.350 702.150 ;
        RECT 157.950 701.850 160.050 703.950 ;
        RECT 160.950 703.050 163.050 705.150 ;
        RECT 166.950 703.050 169.050 705.150 ;
        RECT 175.650 702.150 176.850 707.400 ;
        RECT 137.550 695.100 145.050 696.300 ;
        RECT 137.550 687.750 139.350 695.100 ;
        RECT 143.250 694.500 145.050 695.100 ;
        RECT 147.150 693.600 148.350 700.050 ;
        RECT 158.400 697.650 159.600 701.850 ;
        RECT 175.650 700.050 178.050 702.150 ;
        RECT 178.950 701.850 181.050 703.950 ;
        RECT 179.100 700.050 180.900 701.850 ;
        RECT 158.400 696.000 162.900 697.650 ;
        RECT 142.050 687.750 143.850 693.600 ;
        RECT 145.050 692.100 148.350 693.600 ;
        RECT 145.050 687.750 146.850 692.100 ;
        RECT 161.100 687.750 162.900 696.000 ;
        RECT 166.500 687.750 168.300 696.600 ;
        RECT 175.650 693.600 176.850 700.050 ;
        RECT 182.100 696.300 183.300 713.400 ;
        RECT 191.550 707.400 193.350 719.250 ;
        RECT 195.750 707.400 197.550 719.250 ;
        RECT 205.350 707.400 207.150 719.250 ;
        RECT 208.350 707.400 210.150 719.250 ;
        RECT 211.650 713.400 213.450 719.250 ;
        RECT 215.700 713.400 217.500 719.250 ;
        RECT 218.700 713.400 220.500 719.250 ;
        RECT 221.700 713.400 223.500 719.250 ;
        RECT 195.000 706.350 197.550 707.400 ;
        RECT 185.100 702.150 186.900 703.950 ;
        RECT 191.100 702.150 192.900 703.950 ;
        RECT 184.950 700.050 187.050 702.150 ;
        RECT 190.950 700.050 193.050 702.150 ;
        RECT 195.000 699.150 196.050 706.350 ;
        RECT 197.100 702.150 198.900 703.950 ;
        RECT 205.650 702.150 206.850 707.400 ;
        RECT 212.250 706.500 213.450 713.400 ;
        RECT 218.700 712.500 219.750 713.400 ;
        RECT 207.750 705.600 213.450 706.500 ;
        RECT 215.700 711.600 219.750 712.500 ;
        RECT 207.750 704.700 210.000 705.600 ;
        RECT 196.950 700.050 199.050 702.150 ;
        RECT 205.650 700.050 208.050 702.150 ;
        RECT 193.950 697.050 196.050 699.150 ;
        RECT 178.950 695.100 186.450 696.300 ;
        RECT 178.950 694.500 180.750 695.100 ;
        RECT 175.650 692.100 178.950 693.600 ;
        RECT 177.150 687.750 178.950 692.100 ;
        RECT 180.150 687.750 181.950 693.600 ;
        RECT 184.650 687.750 186.450 695.100 ;
        RECT 195.000 690.600 196.050 697.050 ;
        RECT 205.650 693.600 206.850 700.050 ;
        RECT 208.950 696.300 210.000 704.700 ;
        RECT 212.100 702.150 213.900 703.950 ;
        RECT 211.950 700.050 214.050 702.150 ;
        RECT 207.750 695.400 210.000 696.300 ;
        RECT 215.700 698.100 216.900 711.600 ;
        RECT 224.700 710.700 226.500 719.250 ;
        RECT 227.700 715.950 229.500 719.250 ;
        RECT 230.850 716.400 233.250 719.250 ;
        RECT 234.150 716.400 236.250 719.250 ;
        RECT 237.300 716.400 239.250 719.250 ;
        RECT 230.850 715.050 232.050 716.400 ;
        RECT 234.150 715.050 235.050 716.400 ;
        RECT 237.300 715.050 238.500 716.400 ;
        RECT 229.950 712.950 232.050 715.050 ;
        RECT 232.950 712.950 235.050 715.050 ;
        RECT 235.950 713.400 238.500 715.050 ;
        RECT 240.450 713.400 242.250 719.250 ;
        RECT 244.200 713.400 246.000 719.250 ;
        RECT 247.200 713.400 249.000 719.250 ;
        RECT 235.950 712.950 238.050 713.400 ;
        RECT 244.650 712.500 246.000 713.400 ;
        RECT 250.200 712.500 252.000 719.250 ;
        RECT 253.950 716.400 255.750 719.250 ;
        RECT 244.650 710.850 247.050 712.500 ;
        RECT 220.200 709.650 237.900 710.700 ;
        RECT 244.950 710.400 247.050 710.850 ;
        RECT 249.000 712.200 252.000 712.500 ;
        RECT 249.000 710.400 252.900 712.200 ;
        RECT 220.200 708.900 222.000 709.650 ;
        RECT 232.950 708.150 235.050 708.750 ;
        RECT 223.500 706.950 235.050 708.150 ;
        RECT 235.950 708.600 237.900 709.650 ;
        RECT 254.100 709.350 255.450 716.400 ;
        RECT 256.950 712.950 258.750 719.250 ;
        RECT 259.950 716.400 261.750 719.250 ;
        RECT 260.100 715.200 261.600 716.400 ;
        RECT 260.100 713.100 262.200 715.200 ;
        RECT 263.700 713.400 265.500 719.250 ;
        RECT 256.950 712.050 259.050 712.950 ;
        RECT 266.700 712.500 268.500 719.250 ;
        RECT 269.700 713.400 271.500 719.250 ;
        RECT 272.700 713.400 274.500 719.250 ;
        RECT 275.700 713.400 277.500 719.250 ;
        RECT 279.450 713.400 281.250 719.250 ;
        RECT 282.450 713.400 284.250 719.250 ;
        RECT 263.850 712.050 265.650 712.500 ;
        RECT 256.950 710.850 265.650 712.050 ;
        RECT 266.700 711.300 272.400 712.500 ;
        RECT 263.850 710.700 265.650 710.850 ;
        RECT 270.600 710.700 272.400 711.300 ;
        RECT 273.300 709.350 274.500 713.400 ;
        RECT 253.950 708.600 256.050 709.350 ;
        RECT 235.950 707.250 256.050 708.600 ;
        RECT 259.950 708.450 277.350 709.350 ;
        RECT 259.950 707.250 262.050 708.450 ;
        RECT 223.500 706.350 225.300 706.950 ;
        RECT 232.950 706.650 235.050 706.950 ;
        RECT 262.950 706.350 275.250 707.550 ;
        RECT 235.950 705.450 264.000 706.350 ;
        RECT 273.450 705.750 275.250 706.350 ;
        RECT 224.250 705.150 264.000 705.450 ;
        RECT 223.950 704.550 237.900 705.150 ;
        RECT 217.950 701.850 220.050 703.950 ;
        RECT 223.950 703.350 227.850 704.550 ;
        RECT 244.950 703.650 259.500 704.250 ;
        RECT 223.950 703.050 226.050 703.350 ;
        RECT 228.750 702.450 235.500 703.350 ;
        RECT 218.100 700.050 219.900 701.850 ;
        RECT 228.750 700.050 229.950 702.450 ;
        RECT 218.100 699.000 229.950 700.050 ;
        RECT 231.750 699.750 233.550 701.550 ;
        RECT 234.450 700.950 235.500 702.450 ;
        RECT 236.400 703.050 259.500 703.650 ;
        RECT 236.400 702.450 247.050 703.050 ;
        RECT 236.400 701.850 238.200 702.450 ;
        RECT 244.950 702.150 247.050 702.450 ;
        RECT 249.150 701.250 251.250 701.550 ;
        RECT 257.700 701.250 259.500 703.050 ;
        RECT 260.850 702.000 267.900 703.800 ;
        RECT 234.450 700.050 246.450 700.950 ;
        RECT 215.700 697.200 231.000 698.100 ;
        RECT 207.750 694.500 212.850 695.400 ;
        RECT 191.550 687.750 193.350 690.600 ;
        RECT 194.550 687.750 196.350 690.600 ;
        RECT 197.550 687.750 199.350 690.600 ;
        RECT 205.350 687.750 207.150 693.600 ;
        RECT 208.350 687.750 210.150 693.600 ;
        RECT 211.650 690.600 212.850 694.500 ;
        RECT 215.700 693.600 216.900 697.200 ;
        RECT 219.900 695.700 221.700 696.300 ;
        RECT 219.900 694.500 228.300 695.700 ;
        RECT 226.800 693.600 228.300 694.500 ;
        RECT 211.650 687.750 213.450 690.600 ;
        RECT 215.700 687.750 217.500 693.600 ;
        RECT 221.100 687.750 222.900 693.600 ;
        RECT 226.500 687.750 228.300 693.600 ;
        RECT 229.950 694.050 231.000 697.200 ;
        RECT 232.500 696.300 233.550 699.750 ;
        RECT 240.150 697.350 244.050 699.150 ;
        RECT 241.950 697.050 244.050 697.350 ;
        RECT 245.400 698.550 246.450 700.050 ;
        RECT 247.350 699.450 251.250 701.250 ;
        RECT 260.850 700.350 261.750 702.000 ;
        RECT 268.950 701.100 271.050 705.150 ;
        RECT 252.150 699.300 261.750 700.350 ;
        RECT 262.800 700.050 271.050 701.100 ;
        RECT 252.150 698.550 253.050 699.300 ;
        RECT 245.400 697.200 253.050 698.550 ;
        RECT 262.800 698.250 263.850 700.050 ;
        RECT 253.950 697.200 263.850 698.250 ;
        RECT 267.300 697.200 275.100 699.000 ;
        RECT 235.050 696.300 236.850 696.750 ;
        RECT 253.950 696.300 255.000 697.200 ;
        RECT 232.500 695.850 236.850 696.300 ;
        RECT 232.500 695.100 240.150 695.850 ;
        RECT 235.050 694.950 240.150 695.100 ;
        RECT 229.950 691.950 232.050 694.050 ;
        RECT 232.950 691.950 235.050 694.050 ;
        RECT 235.950 691.950 238.050 694.050 ;
        RECT 239.250 693.600 240.150 694.950 ;
        RECT 248.100 694.500 255.000 696.300 ;
        RECT 255.900 694.500 262.650 696.300 ;
        RECT 267.300 693.600 268.800 697.200 ;
        RECT 276.150 693.600 277.350 708.450 ;
        RECT 239.250 692.250 243.300 693.600 ;
        RECT 244.950 693.300 247.050 693.600 ;
        RECT 230.700 690.600 232.050 691.950 ;
        RECT 233.700 690.600 235.050 691.950 ;
        RECT 236.700 690.600 238.050 691.950 ;
        RECT 241.500 691.800 243.300 692.250 ;
        RECT 244.200 691.500 247.050 693.300 ;
        RECT 249.150 693.300 251.250 693.600 ;
        RECT 249.150 691.500 252.000 693.300 ;
        RECT 230.700 687.750 232.500 690.600 ;
        RECT 233.700 687.750 235.500 690.600 ;
        RECT 236.700 687.750 238.500 690.600 ;
        RECT 239.700 687.750 241.500 690.600 ;
        RECT 244.200 687.750 246.000 691.500 ;
        RECT 247.200 687.750 249.000 690.600 ;
        RECT 250.200 687.750 252.000 691.500 ;
        RECT 253.950 691.500 256.050 693.600 ;
        RECT 256.950 691.500 259.050 693.600 ;
        RECT 259.950 691.500 262.050 693.600 ;
        RECT 264.600 692.400 268.800 693.600 ;
        RECT 253.950 687.750 255.750 691.500 ;
        RECT 256.950 687.750 258.750 691.500 ;
        RECT 259.950 687.750 261.750 691.500 ;
        RECT 264.600 687.750 266.400 692.400 ;
        RECT 270.150 687.750 271.950 693.600 ;
        RECT 275.550 687.750 277.350 693.600 ;
        RECT 279.450 700.950 280.950 713.400 ;
        RECT 292.650 707.400 294.450 719.250 ;
        RECT 295.650 708.300 297.450 719.250 ;
        RECT 298.650 709.200 300.450 719.250 ;
        RECT 301.650 708.300 303.450 719.250 ;
        RECT 308.550 713.400 310.350 719.250 ;
        RECT 311.550 713.400 313.350 719.250 ;
        RECT 314.550 713.400 316.350 719.250 ;
        RECT 295.650 707.400 303.450 708.300 ;
        RECT 293.100 702.150 294.300 707.400 ;
        RECT 311.550 705.150 312.750 713.400 ;
        RECT 325.650 707.400 327.450 719.250 ;
        RECT 328.650 708.300 330.450 719.250 ;
        RECT 331.650 709.200 333.450 719.250 ;
        RECT 334.650 708.300 336.450 719.250 ;
        RECT 328.650 707.400 336.450 708.300 ;
        RECT 338.550 708.300 340.350 719.250 ;
        RECT 341.550 709.200 343.350 719.250 ;
        RECT 344.550 708.300 346.350 719.250 ;
        RECT 338.550 707.400 346.350 708.300 ;
        RECT 347.550 707.400 349.350 719.250 ;
        RECT 359.550 707.400 361.350 719.250 ;
        RECT 363.750 707.400 365.550 719.250 ;
        RECT 373.650 713.400 375.450 719.250 ;
        RECT 376.650 713.400 378.450 719.250 ;
        RECT 379.650 713.400 381.450 719.250 ;
        RECT 385.650 713.400 387.450 719.250 ;
        RECT 388.650 714.000 390.450 719.250 ;
        RECT 279.450 698.850 283.050 700.950 ;
        RECT 292.950 700.050 295.050 702.150 ;
        RECT 307.950 701.850 310.050 703.950 ;
        RECT 310.950 703.050 313.050 705.150 ;
        RECT 279.450 690.600 280.950 698.850 ;
        RECT 293.100 693.600 294.300 700.050 ;
        RECT 295.950 698.850 298.050 700.950 ;
        RECT 299.100 699.150 300.900 700.950 ;
        RECT 296.100 697.050 297.900 698.850 ;
        RECT 298.950 697.050 301.050 699.150 ;
        RECT 301.950 698.850 304.050 700.950 ;
        RECT 308.100 700.050 309.900 701.850 ;
        RECT 302.100 697.050 303.900 698.850 ;
        RECT 311.550 695.700 312.750 703.050 ;
        RECT 313.950 701.850 316.050 703.950 ;
        RECT 326.100 702.150 327.300 707.400 ;
        RECT 347.700 702.150 348.900 707.400 ;
        RECT 363.000 706.350 365.550 707.400 ;
        RECT 359.100 702.150 360.900 703.950 ;
        RECT 314.100 700.050 315.900 701.850 ;
        RECT 325.950 700.050 328.050 702.150 ;
        RECT 311.550 694.800 315.150 695.700 ;
        RECT 293.100 691.950 298.800 693.600 ;
        RECT 279.450 687.750 281.250 690.600 ;
        RECT 282.450 687.750 284.250 690.600 ;
        RECT 293.700 687.750 295.500 690.600 ;
        RECT 297.000 687.750 298.800 691.950 ;
        RECT 301.200 687.750 303.000 693.600 ;
        RECT 308.850 687.750 310.650 693.600 ;
        RECT 313.350 687.750 315.150 694.800 ;
        RECT 326.100 693.600 327.300 700.050 ;
        RECT 328.950 698.850 331.050 700.950 ;
        RECT 332.100 699.150 333.900 700.950 ;
        RECT 329.100 697.050 330.900 698.850 ;
        RECT 331.950 697.050 334.050 699.150 ;
        RECT 334.950 698.850 337.050 700.950 ;
        RECT 337.950 698.850 340.050 700.950 ;
        RECT 341.100 699.150 342.900 700.950 ;
        RECT 335.100 697.050 336.900 698.850 ;
        RECT 338.100 697.050 339.900 698.850 ;
        RECT 340.950 697.050 343.050 699.150 ;
        RECT 343.950 698.850 346.050 700.950 ;
        RECT 346.950 700.050 349.050 702.150 ;
        RECT 358.950 700.050 361.050 702.150 ;
        RECT 344.100 697.050 345.900 698.850 ;
        RECT 347.700 693.600 348.900 700.050 ;
        RECT 363.000 699.150 364.050 706.350 ;
        RECT 377.250 705.150 378.450 713.400 ;
        RECT 386.250 713.100 387.450 713.400 ;
        RECT 391.650 713.400 393.450 719.250 ;
        RECT 394.650 713.400 396.450 719.250 ;
        RECT 391.650 713.100 393.300 713.400 ;
        RECT 386.250 712.200 393.300 713.100 ;
        RECT 365.100 702.150 366.900 703.950 ;
        RECT 364.950 700.050 367.050 702.150 ;
        RECT 373.950 701.850 376.050 703.950 ;
        RECT 376.950 703.050 379.050 705.150 ;
        RECT 386.250 703.950 387.300 712.200 ;
        RECT 392.100 708.150 393.900 709.950 ;
        RECT 404.550 708.300 406.350 719.250 ;
        RECT 407.550 709.200 409.350 719.250 ;
        RECT 410.550 708.300 412.350 719.250 ;
        RECT 388.950 705.150 390.750 706.950 ;
        RECT 391.950 706.050 394.050 708.150 ;
        RECT 404.550 707.400 412.350 708.300 ;
        RECT 413.550 707.400 415.350 719.250 ;
        RECT 422.400 713.400 424.200 719.250 ;
        RECT 425.700 707.400 427.500 719.250 ;
        RECT 429.900 707.400 431.700 719.250 ;
        RECT 437.550 713.400 439.350 719.250 ;
        RECT 440.550 713.400 442.350 719.250 ;
        RECT 443.550 713.400 445.350 719.250 ;
        RECT 452.550 713.400 454.350 719.250 ;
        RECT 455.550 713.400 457.350 719.250 ;
        RECT 458.550 713.400 460.350 719.250 ;
        RECT 467.550 713.400 469.350 719.250 ;
        RECT 470.550 713.400 472.350 719.250 ;
        RECT 482.550 713.400 484.350 719.250 ;
        RECT 485.550 713.400 487.350 719.250 ;
        RECT 488.550 713.400 490.350 719.250 ;
        RECT 502.650 713.400 504.450 719.250 ;
        RECT 505.650 714.000 507.450 719.250 ;
        RECT 395.100 705.150 396.900 706.950 ;
        RECT 374.100 700.050 375.900 701.850 ;
        RECT 361.950 697.050 364.050 699.150 ;
        RECT 349.950 694.950 352.050 697.050 ;
        RECT 326.100 691.950 331.800 693.600 ;
        RECT 326.700 687.750 328.500 690.600 ;
        RECT 330.000 687.750 331.800 691.950 ;
        RECT 334.200 687.750 336.000 693.600 ;
        RECT 339.000 687.750 340.800 693.600 ;
        RECT 343.200 691.950 348.900 693.600 ;
        RECT 350.550 693.450 351.450 694.950 ;
        RECT 358.950 693.450 361.050 694.050 ;
        RECT 350.550 692.550 361.050 693.450 ;
        RECT 358.950 691.950 361.050 692.550 ;
        RECT 343.200 687.750 345.000 691.950 ;
        RECT 363.000 690.600 364.050 697.050 ;
        RECT 377.250 695.700 378.450 703.050 ;
        RECT 379.950 701.850 382.050 703.950 ;
        RECT 385.950 701.850 388.050 703.950 ;
        RECT 388.950 703.050 391.050 705.150 ;
        RECT 394.950 703.050 397.050 705.150 ;
        RECT 413.700 702.150 414.900 707.400 ;
        RECT 422.250 705.150 424.050 706.950 ;
        RECT 421.950 703.050 424.050 705.150 ;
        RECT 425.850 702.150 427.050 707.400 ;
        RECT 440.550 705.150 441.750 713.400 ;
        RECT 455.550 705.150 456.750 713.400 ;
        RECT 431.100 702.150 432.900 703.950 ;
        RECT 380.100 700.050 381.900 701.850 ;
        RECT 386.400 697.650 387.600 701.850 ;
        RECT 403.950 698.850 406.050 700.950 ;
        RECT 407.100 699.150 408.900 700.950 ;
        RECT 386.400 696.000 390.900 697.650 ;
        RECT 404.100 697.050 405.900 698.850 ;
        RECT 406.950 697.050 409.050 699.150 ;
        RECT 409.950 698.850 412.050 700.950 ;
        RECT 412.950 700.050 415.050 702.150 ;
        RECT 424.950 700.050 427.050 702.150 ;
        RECT 410.100 697.050 411.900 698.850 ;
        RECT 374.850 694.800 378.450 695.700 ;
        RECT 346.500 687.750 348.300 690.600 ;
        RECT 359.550 687.750 361.350 690.600 ;
        RECT 362.550 687.750 364.350 690.600 ;
        RECT 365.550 687.750 367.350 690.600 ;
        RECT 374.850 687.750 376.650 694.800 ;
        RECT 379.350 687.750 381.150 693.600 ;
        RECT 389.100 687.750 390.900 696.000 ;
        RECT 394.500 687.750 396.300 696.600 ;
        RECT 413.700 693.600 414.900 700.050 ;
        RECT 424.950 696.750 426.150 700.050 ;
        RECT 427.950 698.850 430.050 700.950 ;
        RECT 430.950 700.050 433.050 702.150 ;
        RECT 436.950 701.850 439.050 703.950 ;
        RECT 439.950 703.050 442.050 705.150 ;
        RECT 437.100 700.050 438.900 701.850 ;
        RECT 428.100 697.050 429.900 698.850 ;
        RECT 422.250 695.700 426.000 696.750 ;
        RECT 440.550 695.700 441.750 703.050 ;
        RECT 442.950 701.850 445.050 703.950 ;
        RECT 451.950 701.850 454.050 703.950 ;
        RECT 454.950 703.050 457.050 705.150 ;
        RECT 443.100 700.050 444.900 701.850 ;
        RECT 452.100 700.050 453.900 701.850 ;
        RECT 455.550 695.700 456.750 703.050 ;
        RECT 457.950 701.850 460.050 703.950 ;
        RECT 458.100 700.050 459.900 701.850 ;
        RECT 470.400 700.950 471.600 713.400 ;
        RECT 485.550 705.150 486.750 713.400 ;
        RECT 503.250 713.100 504.450 713.400 ;
        RECT 508.650 713.400 510.450 719.250 ;
        RECT 511.650 713.400 513.450 719.250 ;
        RECT 508.650 713.100 510.300 713.400 ;
        RECT 503.250 712.200 510.300 713.100 ;
        RECT 481.950 701.850 484.050 703.950 ;
        RECT 484.950 703.050 487.050 705.150 ;
        RECT 503.250 703.950 504.300 712.200 ;
        RECT 509.100 708.150 510.900 709.950 ;
        RECT 505.950 705.150 507.750 706.950 ;
        RECT 508.950 706.050 511.050 708.150 ;
        RECT 525.450 707.400 527.250 719.250 ;
        RECT 529.650 707.400 531.450 719.250 ;
        RECT 538.650 713.400 540.450 719.250 ;
        RECT 541.650 713.400 543.450 719.250 ;
        RECT 547.650 713.400 549.450 719.250 ;
        RECT 550.650 714.000 552.450 719.250 ;
        RECT 512.100 705.150 513.900 706.950 ;
        RECT 525.450 706.350 528.000 707.400 ;
        RECT 467.100 699.150 468.900 700.950 ;
        RECT 466.950 697.050 469.050 699.150 ;
        RECT 469.950 698.850 472.050 700.950 ;
        RECT 482.100 700.050 483.900 701.850 ;
        RECT 422.250 693.600 423.450 695.700 ;
        RECT 440.550 694.800 444.150 695.700 ;
        RECT 455.550 694.800 459.150 695.700 ;
        RECT 405.000 687.750 406.800 693.600 ;
        RECT 409.200 691.950 414.900 693.600 ;
        RECT 409.200 687.750 411.000 691.950 ;
        RECT 412.500 687.750 414.300 690.600 ;
        RECT 421.650 687.750 423.450 693.600 ;
        RECT 424.650 692.700 432.450 694.050 ;
        RECT 424.650 687.750 426.450 692.700 ;
        RECT 427.650 687.750 429.450 691.800 ;
        RECT 430.650 687.750 432.450 692.700 ;
        RECT 437.850 687.750 439.650 693.600 ;
        RECT 442.350 687.750 444.150 694.800 ;
        RECT 452.850 687.750 454.650 693.600 ;
        RECT 457.350 687.750 459.150 694.800 ;
        RECT 470.400 690.600 471.600 698.850 ;
        RECT 485.550 695.700 486.750 703.050 ;
        RECT 487.950 701.850 490.050 703.950 ;
        RECT 502.950 701.850 505.050 703.950 ;
        RECT 505.950 703.050 508.050 705.150 ;
        RECT 511.950 703.050 514.050 705.150 ;
        RECT 524.100 702.150 525.900 703.950 ;
        RECT 488.100 700.050 489.900 701.850 ;
        RECT 503.400 697.650 504.600 701.850 ;
        RECT 523.950 700.050 526.050 702.150 ;
        RECT 526.950 699.150 528.000 706.350 ;
        RECT 530.100 702.150 531.900 703.950 ;
        RECT 529.950 700.050 532.050 702.150 ;
        RECT 539.400 700.950 540.600 713.400 ;
        RECT 548.250 713.100 549.450 713.400 ;
        RECT 553.650 713.400 555.450 719.250 ;
        RECT 556.650 713.400 558.450 719.250 ;
        RECT 563.550 713.400 565.350 719.250 ;
        RECT 566.550 713.400 568.350 719.250 ;
        RECT 569.550 713.400 571.350 719.250 ;
        RECT 553.650 713.100 555.300 713.400 ;
        RECT 548.250 712.200 555.300 713.100 ;
        RECT 541.950 705.450 544.050 706.050 ;
        RECT 541.950 704.550 546.450 705.450 ;
        RECT 541.950 703.950 544.050 704.550 ;
        RECT 503.400 696.000 507.900 697.650 ;
        RECT 526.950 697.050 529.050 699.150 ;
        RECT 538.950 698.850 541.050 700.950 ;
        RECT 542.100 699.150 543.900 700.950 ;
        RECT 485.550 694.800 489.150 695.700 ;
        RECT 467.550 687.750 469.350 690.600 ;
        RECT 470.550 687.750 472.350 690.600 ;
        RECT 482.850 687.750 484.650 693.600 ;
        RECT 487.350 687.750 489.150 694.800 ;
        RECT 506.100 687.750 507.900 696.000 ;
        RECT 511.500 687.750 513.300 696.600 ;
        RECT 526.950 690.600 528.000 697.050 ;
        RECT 539.400 690.600 540.600 698.850 ;
        RECT 541.950 697.050 544.050 699.150 ;
        RECT 545.550 694.050 546.450 704.550 ;
        RECT 548.250 703.950 549.300 712.200 ;
        RECT 556.950 711.450 559.050 712.050 ;
        RECT 556.950 710.550 561.450 711.450 ;
        RECT 556.950 709.950 559.050 710.550 ;
        RECT 554.100 708.150 555.900 709.950 ;
        RECT 550.950 705.150 552.750 706.950 ;
        RECT 553.950 706.050 556.050 708.150 ;
        RECT 557.100 705.150 558.900 706.950 ;
        RECT 547.950 701.850 550.050 703.950 ;
        RECT 550.950 703.050 553.050 705.150 ;
        RECT 556.950 703.050 559.050 705.150 ;
        RECT 548.400 697.650 549.600 701.850 ;
        RECT 556.950 699.450 559.050 700.050 ;
        RECT 560.550 699.450 561.450 710.550 ;
        RECT 566.550 705.150 567.750 713.400 ;
        RECT 578.550 707.400 580.350 719.250 ;
        RECT 583.050 707.550 584.850 719.250 ;
        RECT 586.050 708.900 587.850 719.250 ;
        RECT 596.550 713.400 598.350 719.250 ;
        RECT 599.550 713.400 601.350 719.250 ;
        RECT 602.550 713.400 604.350 719.250 ;
        RECT 586.050 707.550 588.450 708.900 ;
        RECT 578.550 706.200 579.750 707.400 ;
        RECT 583.950 706.200 585.750 706.650 ;
        RECT 562.950 701.850 565.050 703.950 ;
        RECT 565.950 703.050 568.050 705.150 ;
        RECT 578.550 705.000 585.750 706.200 ;
        RECT 583.950 704.850 585.750 705.000 ;
        RECT 563.100 700.050 564.900 701.850 ;
        RECT 556.950 698.550 561.450 699.450 ;
        RECT 556.950 697.950 559.050 698.550 ;
        RECT 548.400 696.000 552.900 697.650 ;
        RECT 544.950 691.950 547.050 694.050 ;
        RECT 523.650 687.750 525.450 690.600 ;
        RECT 526.650 687.750 528.450 690.600 ;
        RECT 529.650 687.750 531.450 690.600 ;
        RECT 538.650 687.750 540.450 690.600 ;
        RECT 541.650 687.750 543.450 690.600 ;
        RECT 551.100 687.750 552.900 696.000 ;
        RECT 556.500 687.750 558.300 696.600 ;
        RECT 566.550 695.700 567.750 703.050 ;
        RECT 568.950 701.850 571.050 703.950 ;
        RECT 581.100 702.150 582.900 703.950 ;
        RECT 569.100 700.050 570.900 701.850 ;
        RECT 578.100 699.150 579.900 700.950 ;
        RECT 580.950 700.050 583.050 702.150 ;
        RECT 577.950 697.050 580.050 699.150 ;
        RECT 584.700 696.600 585.600 704.850 ;
        RECT 587.100 700.950 588.450 707.550 ;
        RECT 599.550 705.150 600.750 713.400 ;
        RECT 615.300 707.400 617.100 719.250 ;
        RECT 619.500 707.400 621.300 719.250 ;
        RECT 622.800 713.400 624.600 719.250 ;
        RECT 632.550 713.400 634.350 719.250 ;
        RECT 635.550 713.400 637.350 719.250 ;
        RECT 638.550 713.400 640.350 719.250 ;
        RECT 646.650 713.400 648.450 719.250 ;
        RECT 649.650 713.400 651.450 719.250 ;
        RECT 652.650 713.400 654.450 719.250 ;
        RECT 661.650 713.400 663.450 719.250 ;
        RECT 664.650 714.000 666.450 719.250 ;
        RECT 631.950 711.450 634.050 712.050 ;
        RECT 626.550 710.550 634.050 711.450 ;
        RECT 595.950 701.850 598.050 703.950 ;
        RECT 598.950 703.050 601.050 705.150 ;
        RECT 586.950 698.850 589.050 700.950 ;
        RECT 596.100 700.050 597.900 701.850 ;
        RECT 583.950 695.700 585.750 696.600 ;
        RECT 566.550 694.800 570.150 695.700 ;
        RECT 563.850 687.750 565.650 693.600 ;
        RECT 568.350 687.750 570.150 694.800 ;
        RECT 582.450 694.800 585.750 695.700 ;
        RECT 582.450 690.600 583.350 694.800 ;
        RECT 588.000 693.600 589.050 698.850 ;
        RECT 599.550 695.700 600.750 703.050 ;
        RECT 601.950 701.850 604.050 703.950 ;
        RECT 614.100 702.150 615.900 703.950 ;
        RECT 619.950 702.150 621.150 707.400 ;
        RECT 622.950 705.150 624.750 706.950 ;
        RECT 622.950 703.050 625.050 705.150 ;
        RECT 602.100 700.050 603.900 701.850 ;
        RECT 613.950 700.050 616.050 702.150 ;
        RECT 616.950 698.850 619.050 700.950 ;
        RECT 619.950 700.050 622.050 702.150 ;
        RECT 617.100 697.050 618.900 698.850 ;
        RECT 620.850 696.750 622.050 700.050 ;
        RECT 621.000 695.700 624.750 696.750 ;
        RECT 599.550 694.800 603.150 695.700 ;
        RECT 578.550 687.750 580.350 690.600 ;
        RECT 581.550 687.750 583.350 690.600 ;
        RECT 584.550 687.750 586.350 690.600 ;
        RECT 587.550 687.750 589.350 693.600 ;
        RECT 596.850 687.750 598.650 693.600 ;
        RECT 601.350 687.750 603.150 694.800 ;
        RECT 614.550 692.700 622.350 694.050 ;
        RECT 614.550 687.750 616.350 692.700 ;
        RECT 617.550 687.750 619.350 691.800 ;
        RECT 620.550 687.750 622.350 692.700 ;
        RECT 623.550 693.600 624.750 695.700 ;
        RECT 626.550 696.450 627.450 710.550 ;
        RECT 631.950 709.950 634.050 710.550 ;
        RECT 631.950 708.450 634.050 709.050 ;
        RECT 629.550 707.550 634.050 708.450 ;
        RECT 629.550 700.050 630.450 707.550 ;
        RECT 631.950 706.950 634.050 707.550 ;
        RECT 635.550 705.150 636.750 713.400 ;
        RECT 650.250 705.150 651.450 713.400 ;
        RECT 662.250 713.100 663.450 713.400 ;
        RECT 667.650 713.400 669.450 719.250 ;
        RECT 670.650 713.400 672.450 719.250 ;
        RECT 679.650 713.400 681.450 719.250 ;
        RECT 682.650 713.400 684.450 719.250 ;
        RECT 685.650 713.400 687.450 719.250 ;
        RECT 695.400 713.400 697.200 719.250 ;
        RECT 667.650 713.100 669.300 713.400 ;
        RECT 662.250 712.200 669.300 713.100 ;
        RECT 631.950 701.850 634.050 703.950 ;
        RECT 634.950 703.050 637.050 705.150 ;
        RECT 632.100 700.050 633.900 701.850 ;
        RECT 628.950 697.950 631.050 700.050 ;
        RECT 631.950 696.450 634.050 697.050 ;
        RECT 626.550 695.550 634.050 696.450 ;
        RECT 631.950 694.950 634.050 695.550 ;
        RECT 635.550 695.700 636.750 703.050 ;
        RECT 637.950 701.850 640.050 703.950 ;
        RECT 646.950 701.850 649.050 703.950 ;
        RECT 649.950 703.050 652.050 705.150 ;
        RECT 662.250 703.950 663.300 712.200 ;
        RECT 668.100 708.150 669.900 709.950 ;
        RECT 664.950 705.150 666.750 706.950 ;
        RECT 667.950 706.050 670.050 708.150 ;
        RECT 671.100 705.150 672.900 706.950 ;
        RECT 683.250 705.150 684.450 713.400 ;
        RECT 698.700 707.400 700.500 719.250 ;
        RECT 702.900 707.400 704.700 719.250 ;
        RECT 712.050 718.500 719.850 719.250 ;
        RECT 712.050 709.200 713.850 718.500 ;
        RECT 715.050 709.800 716.850 717.600 ;
        RECT 715.650 707.400 716.850 709.800 ;
        RECT 718.050 709.800 719.850 718.500 ;
        RECT 721.650 718.500 729.450 719.250 ;
        RECT 721.650 710.700 723.450 718.500 ;
        RECT 724.650 709.800 726.450 717.600 ;
        RECT 718.050 708.900 726.450 709.800 ;
        RECT 727.650 709.500 729.450 718.500 ;
        RECT 730.650 710.400 732.450 719.250 ;
        RECT 733.650 709.500 735.450 719.250 ;
        RECT 742.650 713.400 744.450 719.250 ;
        RECT 745.650 713.400 747.450 719.250 ;
        RECT 748.650 713.400 750.450 719.250 ;
        RECT 727.650 708.600 735.450 709.500 ;
        RECT 695.250 705.150 697.050 706.950 ;
        RECT 638.100 700.050 639.900 701.850 ;
        RECT 647.100 700.050 648.900 701.850 ;
        RECT 650.250 695.700 651.450 703.050 ;
        RECT 652.950 701.850 655.050 703.950 ;
        RECT 661.950 701.850 664.050 703.950 ;
        RECT 664.950 703.050 667.050 705.150 ;
        RECT 670.950 703.050 673.050 705.150 ;
        RECT 679.950 701.850 682.050 703.950 ;
        RECT 682.950 703.050 685.050 705.150 ;
        RECT 653.100 700.050 654.900 701.850 ;
        RECT 662.400 697.650 663.600 701.850 ;
        RECT 680.100 700.050 681.900 701.850 ;
        RECT 662.400 696.000 666.900 697.650 ;
        RECT 635.550 694.800 639.150 695.700 ;
        RECT 623.550 687.750 625.350 693.600 ;
        RECT 632.850 687.750 634.650 693.600 ;
        RECT 637.350 687.750 639.150 694.800 ;
        RECT 647.850 694.800 651.450 695.700 ;
        RECT 647.850 687.750 649.650 694.800 ;
        RECT 652.350 687.750 654.150 693.600 ;
        RECT 665.100 687.750 666.900 696.000 ;
        RECT 670.500 687.750 672.300 696.600 ;
        RECT 683.250 695.700 684.450 703.050 ;
        RECT 685.950 701.850 688.050 703.950 ;
        RECT 694.950 703.050 697.050 705.150 ;
        RECT 698.850 702.150 700.050 707.400 ;
        RECT 715.650 706.200 719.100 707.400 ;
        RECT 704.100 702.150 705.900 703.950 ;
        RECT 686.100 700.050 687.900 701.850 ;
        RECT 697.950 700.050 700.050 702.150 ;
        RECT 697.950 696.750 699.150 700.050 ;
        RECT 700.950 698.850 703.050 700.950 ;
        RECT 703.950 700.050 706.050 702.150 ;
        RECT 717.900 700.950 719.100 706.200 ;
        RECT 746.250 705.150 747.450 713.400 ;
        RECT 756.300 707.400 758.100 719.250 ;
        RECT 760.500 707.400 762.300 719.250 ;
        RECT 763.800 713.400 765.600 719.250 ;
        RECT 771.750 713.400 773.550 719.250 ;
        RECT 774.750 713.400 776.550 719.250 ;
        RECT 778.500 713.400 780.300 719.250 ;
        RECT 781.500 713.400 783.300 719.250 ;
        RECT 784.500 713.400 786.300 719.250 ;
        RECT 722.100 702.150 723.900 703.950 ;
        RECT 731.100 702.150 732.900 703.950 ;
        RECT 715.950 698.850 719.100 700.950 ;
        RECT 721.950 700.050 724.050 702.150 ;
        RECT 724.950 698.850 727.050 700.950 ;
        RECT 730.950 700.050 733.050 702.150 ;
        RECT 742.950 701.850 745.050 703.950 ;
        RECT 745.950 703.050 748.050 705.150 ;
        RECT 743.100 700.050 744.900 701.850 ;
        RECT 701.100 697.050 702.900 698.850 ;
        RECT 680.850 694.800 684.450 695.700 ;
        RECT 695.250 695.700 699.000 696.750 ;
        RECT 680.850 687.750 682.650 694.800 ;
        RECT 695.250 693.600 696.450 695.700 ;
        RECT 685.350 687.750 687.150 693.600 ;
        RECT 694.650 687.750 696.450 693.600 ;
        RECT 697.650 692.700 705.450 694.050 ;
        RECT 697.650 687.750 699.450 692.700 ;
        RECT 700.650 687.750 702.450 691.800 ;
        RECT 703.650 687.750 705.450 692.700 ;
        RECT 717.900 692.400 719.100 698.850 ;
        RECT 725.100 697.050 726.900 698.850 ;
        RECT 746.250 695.700 747.450 703.050 ;
        RECT 748.950 701.850 751.050 703.950 ;
        RECT 755.100 702.150 756.900 703.950 ;
        RECT 760.950 702.150 762.150 707.400 ;
        RECT 763.950 705.150 765.750 706.950 ;
        RECT 763.950 703.050 766.050 705.150 ;
        RECT 749.100 700.050 750.900 701.850 ;
        RECT 754.950 700.050 757.050 702.150 ;
        RECT 757.950 698.850 760.050 700.950 ;
        RECT 760.950 700.050 763.050 702.150 ;
        RECT 775.050 700.950 776.550 713.400 ;
        RECT 781.500 709.350 782.700 713.400 ;
        RECT 787.500 712.500 789.300 719.250 ;
        RECT 790.500 713.400 792.300 719.250 ;
        RECT 794.250 716.400 796.050 719.250 ;
        RECT 794.400 715.200 795.900 716.400 ;
        RECT 793.800 713.100 795.900 715.200 ;
        RECT 797.250 712.950 799.050 719.250 ;
        RECT 800.250 716.400 802.050 719.250 ;
        RECT 783.600 711.300 789.300 712.500 ;
        RECT 790.350 712.050 792.150 712.500 ;
        RECT 796.950 712.050 799.050 712.950 ;
        RECT 783.600 710.700 785.400 711.300 ;
        RECT 790.350 710.850 799.050 712.050 ;
        RECT 790.350 710.700 792.150 710.850 ;
        RECT 800.550 709.350 801.900 716.400 ;
        RECT 804.000 712.500 805.800 719.250 ;
        RECT 807.000 713.400 808.800 719.250 ;
        RECT 810.000 713.400 811.800 719.250 ;
        RECT 813.750 713.400 815.550 719.250 ;
        RECT 816.750 716.400 818.700 719.250 ;
        RECT 819.750 716.400 821.850 719.250 ;
        RECT 822.750 716.400 825.150 719.250 ;
        RECT 817.500 715.050 818.700 716.400 ;
        RECT 820.950 715.050 821.850 716.400 ;
        RECT 823.950 715.050 825.150 716.400 ;
        RECT 826.500 715.950 828.300 719.250 ;
        RECT 817.500 713.400 820.050 715.050 ;
        RECT 810.000 712.500 811.350 713.400 ;
        RECT 817.950 712.950 820.050 713.400 ;
        RECT 820.950 712.950 823.050 715.050 ;
        RECT 823.950 712.950 826.050 715.050 ;
        RECT 804.000 712.200 807.000 712.500 ;
        RECT 803.100 710.400 807.000 712.200 ;
        RECT 808.950 710.850 811.350 712.500 ;
        RECT 808.950 710.400 811.050 710.850 ;
        RECT 829.500 710.700 831.300 719.250 ;
        RECT 832.500 713.400 834.300 719.250 ;
        RECT 835.500 713.400 837.300 719.250 ;
        RECT 838.500 713.400 840.300 719.250 ;
        RECT 847.650 713.400 849.450 719.250 ;
        RECT 850.650 713.400 852.450 719.250 ;
        RECT 836.250 712.500 837.300 713.400 ;
        RECT 836.250 711.600 840.300 712.500 ;
        RECT 818.100 709.650 835.800 710.700 ;
        RECT 758.100 697.050 759.900 698.850 ;
        RECT 761.850 696.750 763.050 700.050 ;
        RECT 772.950 698.850 776.550 700.950 ;
        RECT 762.000 695.700 765.750 696.750 ;
        RECT 743.850 694.800 747.450 695.700 ;
        RECT 717.900 691.500 728.700 692.400 ;
        RECT 721.650 690.600 722.700 691.500 ;
        RECT 727.650 690.600 728.700 691.500 ;
        RECT 721.650 687.750 723.450 690.600 ;
        RECT 724.650 687.750 726.450 690.600 ;
        RECT 727.650 687.750 729.450 690.600 ;
        RECT 730.650 687.750 732.750 690.600 ;
        RECT 743.850 687.750 745.650 694.800 ;
        RECT 748.350 687.750 750.150 693.600 ;
        RECT 755.550 692.700 763.350 694.050 ;
        RECT 755.550 687.750 757.350 692.700 ;
        RECT 758.550 687.750 760.350 691.800 ;
        RECT 761.550 687.750 763.350 692.700 ;
        RECT 764.550 693.600 765.750 695.700 ;
        RECT 764.550 687.750 766.350 693.600 ;
        RECT 775.050 690.600 776.550 698.850 ;
        RECT 771.750 687.750 773.550 690.600 ;
        RECT 774.750 687.750 776.550 690.600 ;
        RECT 778.650 708.450 796.050 709.350 ;
        RECT 778.650 693.600 779.850 708.450 ;
        RECT 780.750 706.350 793.050 707.550 ;
        RECT 793.950 707.250 796.050 708.450 ;
        RECT 799.950 708.600 802.050 709.350 ;
        RECT 818.100 708.600 820.050 709.650 ;
        RECT 834.000 708.900 835.800 709.650 ;
        RECT 799.950 707.250 820.050 708.600 ;
        RECT 820.950 708.150 823.050 708.750 ;
        RECT 820.950 706.950 832.500 708.150 ;
        RECT 820.950 706.650 823.050 706.950 ;
        RECT 830.700 706.350 832.500 706.950 ;
        RECT 780.750 705.750 782.550 706.350 ;
        RECT 792.000 705.450 820.050 706.350 ;
        RECT 792.000 705.150 831.750 705.450 ;
        RECT 784.950 701.100 787.050 705.150 ;
        RECT 818.100 704.550 832.050 705.150 ;
        RECT 788.100 702.000 795.150 703.800 ;
        RECT 784.950 700.050 793.200 701.100 ;
        RECT 780.900 697.200 788.700 699.000 ;
        RECT 792.150 698.250 793.200 700.050 ;
        RECT 794.250 700.350 795.150 702.000 ;
        RECT 796.500 703.650 811.050 704.250 ;
        RECT 796.500 703.050 819.600 703.650 ;
        RECT 828.150 703.350 832.050 704.550 ;
        RECT 796.500 701.250 798.300 703.050 ;
        RECT 808.950 702.450 819.600 703.050 ;
        RECT 808.950 702.150 811.050 702.450 ;
        RECT 817.800 701.850 819.600 702.450 ;
        RECT 820.500 702.450 827.250 703.350 ;
        RECT 829.950 703.050 832.050 703.350 ;
        RECT 804.750 701.250 806.850 701.550 ;
        RECT 794.250 699.300 803.850 700.350 ;
        RECT 804.750 699.450 808.650 701.250 ;
        RECT 820.500 700.950 821.550 702.450 ;
        RECT 809.550 700.050 821.550 700.950 ;
        RECT 802.950 698.550 803.850 699.300 ;
        RECT 809.550 698.550 810.600 700.050 ;
        RECT 822.450 699.750 824.250 701.550 ;
        RECT 826.050 700.050 827.250 702.450 ;
        RECT 835.950 701.850 838.050 703.950 ;
        RECT 836.100 700.050 837.900 701.850 ;
        RECT 792.150 697.200 802.050 698.250 ;
        RECT 802.950 697.200 810.600 698.550 ;
        RECT 811.950 697.350 815.850 699.150 ;
        RECT 787.200 693.600 788.700 697.200 ;
        RECT 801.000 696.300 802.050 697.200 ;
        RECT 811.950 697.050 814.050 697.350 ;
        RECT 819.150 696.300 820.950 696.750 ;
        RECT 822.450 696.300 823.500 699.750 ;
        RECT 826.050 699.000 837.900 700.050 ;
        RECT 839.100 698.100 840.300 711.600 ;
        RECT 848.400 700.950 849.600 713.400 ;
        RECT 847.950 698.850 850.050 700.950 ;
        RECT 851.100 699.150 852.900 700.950 ;
        RECT 793.350 694.500 800.100 696.300 ;
        RECT 801.000 694.500 807.900 696.300 ;
        RECT 819.150 695.850 823.500 696.300 ;
        RECT 815.850 695.100 823.500 695.850 ;
        RECT 825.000 697.200 840.300 698.100 ;
        RECT 815.850 694.950 820.950 695.100 ;
        RECT 815.850 693.600 816.750 694.950 ;
        RECT 825.000 694.050 826.050 697.200 ;
        RECT 834.300 695.700 836.100 696.300 ;
        RECT 778.650 687.750 780.450 693.600 ;
        RECT 784.050 687.750 785.850 693.600 ;
        RECT 787.200 692.400 791.400 693.600 ;
        RECT 789.600 687.750 791.400 692.400 ;
        RECT 793.950 691.500 796.050 693.600 ;
        RECT 796.950 691.500 799.050 693.600 ;
        RECT 799.950 691.500 802.050 693.600 ;
        RECT 804.750 693.300 806.850 693.600 ;
        RECT 794.250 687.750 796.050 691.500 ;
        RECT 797.250 687.750 799.050 691.500 ;
        RECT 800.250 687.750 802.050 691.500 ;
        RECT 804.000 691.500 806.850 693.300 ;
        RECT 808.950 693.300 811.050 693.600 ;
        RECT 808.950 691.500 811.800 693.300 ;
        RECT 812.700 692.250 816.750 693.600 ;
        RECT 812.700 691.800 814.500 692.250 ;
        RECT 817.950 691.950 820.050 694.050 ;
        RECT 820.950 691.950 823.050 694.050 ;
        RECT 823.950 691.950 826.050 694.050 ;
        RECT 827.700 694.500 836.100 695.700 ;
        RECT 827.700 693.600 829.200 694.500 ;
        RECT 839.100 693.600 840.300 697.200 ;
        RECT 804.000 687.750 805.800 691.500 ;
        RECT 807.000 687.750 808.800 690.600 ;
        RECT 810.000 687.750 811.800 691.500 ;
        RECT 817.950 690.600 819.300 691.950 ;
        RECT 820.950 690.600 822.300 691.950 ;
        RECT 823.950 690.600 825.300 691.950 ;
        RECT 814.500 687.750 816.300 690.600 ;
        RECT 817.500 687.750 819.300 690.600 ;
        RECT 820.500 687.750 822.300 690.600 ;
        RECT 823.500 687.750 825.300 690.600 ;
        RECT 827.700 687.750 829.500 693.600 ;
        RECT 833.100 687.750 834.900 693.600 ;
        RECT 838.500 687.750 840.300 693.600 ;
        RECT 848.400 690.600 849.600 698.850 ;
        RECT 850.950 697.050 853.050 699.150 ;
        RECT 847.650 687.750 849.450 690.600 ;
        RECT 850.650 687.750 852.450 690.600 ;
        RECT 2.700 677.400 4.500 683.250 ;
        RECT 8.100 677.400 9.900 683.250 ;
        RECT 13.500 677.400 15.300 683.250 ;
        RECT 17.700 680.400 19.500 683.250 ;
        RECT 20.700 680.400 22.500 683.250 ;
        RECT 23.700 680.400 25.500 683.250 ;
        RECT 26.700 680.400 28.500 683.250 ;
        RECT 17.700 679.050 19.050 680.400 ;
        RECT 20.700 679.050 22.050 680.400 ;
        RECT 23.700 679.050 25.050 680.400 ;
        RECT 31.200 679.500 33.000 683.250 ;
        RECT 34.200 680.400 36.000 683.250 ;
        RECT 37.200 679.500 39.000 683.250 ;
        RECT 2.700 673.800 3.900 677.400 ;
        RECT 13.800 676.500 15.300 677.400 ;
        RECT 6.900 675.300 15.300 676.500 ;
        RECT 16.950 676.950 19.050 679.050 ;
        RECT 19.950 676.950 22.050 679.050 ;
        RECT 22.950 676.950 25.050 679.050 ;
        RECT 28.500 678.750 30.300 679.200 ;
        RECT 26.250 677.400 30.300 678.750 ;
        RECT 31.200 677.700 34.050 679.500 ;
        RECT 31.950 677.400 34.050 677.700 ;
        RECT 36.150 677.700 39.000 679.500 ;
        RECT 40.950 679.500 42.750 683.250 ;
        RECT 43.950 679.500 45.750 683.250 ;
        RECT 46.950 679.500 48.750 683.250 ;
        RECT 36.150 677.400 38.250 677.700 ;
        RECT 40.950 677.400 43.050 679.500 ;
        RECT 43.950 677.400 46.050 679.500 ;
        RECT 46.950 677.400 49.050 679.500 ;
        RECT 51.600 678.600 53.400 683.250 ;
        RECT 51.600 677.400 55.800 678.600 ;
        RECT 57.150 677.400 58.950 683.250 ;
        RECT 62.550 677.400 64.350 683.250 ;
        RECT 6.900 674.700 8.700 675.300 ;
        RECT 16.950 673.800 18.000 676.950 ;
        RECT 26.250 676.050 27.150 677.400 ;
        RECT 22.050 675.900 27.150 676.050 ;
        RECT 2.700 672.900 18.000 673.800 ;
        RECT 19.500 675.150 27.150 675.900 ;
        RECT 19.500 674.700 23.850 675.150 ;
        RECT 35.100 674.700 42.000 676.500 ;
        RECT 42.900 674.700 49.650 676.500 ;
        RECT 2.700 659.400 3.900 672.900 ;
        RECT 5.100 670.950 16.950 672.000 ;
        RECT 19.500 671.250 20.550 674.700 ;
        RECT 22.050 674.250 23.850 674.700 ;
        RECT 28.950 673.650 31.050 673.950 ;
        RECT 40.950 673.800 42.000 674.700 ;
        RECT 54.300 673.800 55.800 677.400 ;
        RECT 27.150 671.850 31.050 673.650 ;
        RECT 32.400 672.450 40.050 673.800 ;
        RECT 40.950 672.750 50.850 673.800 ;
        RECT 5.100 669.150 6.900 670.950 ;
        RECT 4.950 667.050 7.050 669.150 ;
        RECT 15.750 668.550 16.950 670.950 ;
        RECT 18.750 669.450 20.550 671.250 ;
        RECT 32.400 670.950 33.450 672.450 ;
        RECT 39.150 671.700 40.050 672.450 ;
        RECT 21.450 670.050 33.450 670.950 ;
        RECT 21.450 668.550 22.500 670.050 ;
        RECT 34.350 669.750 38.250 671.550 ;
        RECT 39.150 670.650 48.750 671.700 ;
        RECT 36.150 669.450 38.250 669.750 ;
        RECT 10.950 667.650 13.050 667.950 ;
        RECT 15.750 667.650 22.500 668.550 ;
        RECT 23.400 668.550 25.200 669.150 ;
        RECT 31.950 668.550 34.050 668.850 ;
        RECT 23.400 667.950 34.050 668.550 ;
        RECT 44.700 667.950 46.500 669.750 ;
        RECT 10.950 666.450 14.850 667.650 ;
        RECT 23.400 667.350 46.500 667.950 ;
        RECT 31.950 666.750 46.500 667.350 ;
        RECT 47.850 669.000 48.750 670.650 ;
        RECT 49.800 670.950 50.850 672.750 ;
        RECT 54.300 672.000 62.100 673.800 ;
        RECT 49.800 669.900 58.050 670.950 ;
        RECT 47.850 667.200 54.900 669.000 ;
        RECT 10.950 665.850 24.900 666.450 ;
        RECT 55.950 665.850 58.050 669.900 ;
        RECT 11.250 665.550 51.000 665.850 ;
        RECT 22.950 664.650 51.000 665.550 ;
        RECT 60.450 664.650 62.250 665.250 ;
        RECT 10.500 664.050 12.300 664.650 ;
        RECT 19.950 664.050 22.050 664.350 ;
        RECT 10.500 662.850 22.050 664.050 ;
        RECT 19.950 662.250 22.050 662.850 ;
        RECT 22.950 662.400 43.050 663.750 ;
        RECT 7.200 661.350 9.000 662.100 ;
        RECT 22.950 661.350 24.900 662.400 ;
        RECT 40.950 661.650 43.050 662.400 ;
        RECT 46.950 662.550 49.050 663.750 ;
        RECT 49.950 663.450 62.250 664.650 ;
        RECT 63.150 662.550 64.350 677.400 ;
        RECT 46.950 661.650 64.350 662.550 ;
        RECT 66.450 680.400 68.250 683.250 ;
        RECT 69.450 680.400 71.250 683.250 ;
        RECT 79.650 680.400 81.450 683.250 ;
        RECT 82.650 680.400 84.450 683.250 ;
        RECT 66.450 672.150 67.950 680.400 ;
        RECT 80.400 672.150 81.600 680.400 ;
        RECT 91.650 677.400 93.450 683.250 ;
        RECT 92.250 675.300 93.450 677.400 ;
        RECT 94.650 678.300 96.450 683.250 ;
        RECT 97.650 679.200 99.450 683.250 ;
        RECT 100.650 678.300 102.450 683.250 ;
        RECT 94.650 676.950 102.450 678.300 ;
        RECT 110.850 676.200 112.650 683.250 ;
        RECT 115.350 677.400 117.150 683.250 ;
        RECT 122.550 678.300 124.350 683.250 ;
        RECT 125.550 679.200 127.350 683.250 ;
        RECT 128.550 678.300 130.350 683.250 ;
        RECT 122.550 676.950 130.350 678.300 ;
        RECT 131.550 677.400 133.350 683.250 ;
        RECT 140.850 677.400 142.650 683.250 ;
        RECT 110.850 675.300 114.450 676.200 ;
        RECT 131.550 675.300 132.750 677.400 ;
        RECT 145.350 676.200 147.150 683.250 ;
        RECT 157.650 680.400 159.450 683.250 ;
        RECT 160.650 680.400 162.450 683.250 ;
        RECT 163.650 680.400 165.450 683.250 ;
        RECT 92.250 674.250 96.000 675.300 ;
        RECT 66.450 670.050 70.050 672.150 ;
        RECT 79.950 670.050 82.050 672.150 ;
        RECT 82.950 671.850 85.050 673.950 ;
        RECT 83.100 670.050 84.900 671.850 ;
        RECT 94.950 670.950 96.150 674.250 ;
        RECT 98.100 672.150 99.900 673.950 ;
        RECT 7.200 660.300 24.900 661.350 ;
        RECT 2.700 658.500 6.750 659.400 ;
        RECT 5.700 657.600 6.750 658.500 ;
        RECT 2.700 651.750 4.500 657.600 ;
        RECT 5.700 651.750 7.500 657.600 ;
        RECT 8.700 651.750 10.500 657.600 ;
        RECT 11.700 651.750 13.500 660.300 ;
        RECT 31.950 660.150 34.050 660.600 ;
        RECT 31.650 658.500 34.050 660.150 ;
        RECT 36.000 658.800 39.900 660.600 ;
        RECT 36.000 658.500 39.000 658.800 ;
        RECT 16.950 655.950 19.050 658.050 ;
        RECT 19.950 655.950 22.050 658.050 ;
        RECT 22.950 657.600 25.050 658.050 ;
        RECT 31.650 657.600 33.000 658.500 ;
        RECT 22.950 655.950 25.500 657.600 ;
        RECT 14.700 651.750 16.500 655.050 ;
        RECT 17.850 654.600 19.050 655.950 ;
        RECT 21.150 654.600 22.050 655.950 ;
        RECT 24.300 654.600 25.500 655.950 ;
        RECT 17.850 651.750 20.250 654.600 ;
        RECT 21.150 651.750 23.250 654.600 ;
        RECT 24.300 651.750 26.250 654.600 ;
        RECT 27.450 651.750 29.250 657.600 ;
        RECT 31.200 651.750 33.000 657.600 ;
        RECT 34.200 651.750 36.000 657.600 ;
        RECT 37.200 651.750 39.000 658.500 ;
        RECT 41.100 654.600 42.450 661.650 ;
        RECT 50.850 660.150 52.650 660.300 ;
        RECT 43.950 658.950 52.650 660.150 ;
        RECT 57.600 659.700 59.400 660.300 ;
        RECT 43.950 658.050 46.050 658.950 ;
        RECT 50.850 658.500 52.650 658.950 ;
        RECT 53.700 658.500 59.400 659.700 ;
        RECT 40.950 651.750 42.750 654.600 ;
        RECT 43.950 651.750 45.750 658.050 ;
        RECT 47.100 655.800 49.200 657.900 ;
        RECT 47.100 654.600 48.600 655.800 ;
        RECT 46.950 651.750 48.750 654.600 ;
        RECT 50.700 651.750 52.500 657.600 ;
        RECT 53.700 651.750 55.500 658.500 ;
        RECT 60.300 657.600 61.500 661.650 ;
        RECT 66.450 657.600 67.950 670.050 ;
        RECT 80.400 657.600 81.600 670.050 ;
        RECT 94.950 668.850 97.050 670.950 ;
        RECT 97.950 670.050 100.050 672.150 ;
        RECT 100.950 668.850 103.050 670.950 ;
        RECT 110.100 669.150 111.900 670.950 ;
        RECT 91.950 665.850 94.050 667.950 ;
        RECT 92.250 664.050 94.050 665.850 ;
        RECT 95.850 663.600 97.050 668.850 ;
        RECT 101.100 667.050 102.900 668.850 ;
        RECT 109.950 667.050 112.050 669.150 ;
        RECT 113.250 667.950 114.450 675.300 ;
        RECT 129.000 674.250 132.750 675.300 ;
        RECT 143.550 675.300 147.150 676.200 ;
        RECT 125.100 672.150 126.900 673.950 ;
        RECT 116.100 669.150 117.900 670.950 ;
        RECT 112.950 665.850 115.050 667.950 ;
        RECT 115.950 667.050 118.050 669.150 ;
        RECT 121.950 668.850 124.050 670.950 ;
        RECT 124.950 670.050 127.050 672.150 ;
        RECT 128.850 670.950 130.050 674.250 ;
        RECT 127.950 668.850 130.050 670.950 ;
        RECT 140.100 669.150 141.900 670.950 ;
        RECT 122.100 667.050 123.900 668.850 ;
        RECT 56.700 651.750 58.500 657.600 ;
        RECT 59.700 651.750 61.500 657.600 ;
        RECT 62.700 651.750 64.500 657.600 ;
        RECT 66.450 651.750 68.250 657.600 ;
        RECT 69.450 651.750 71.250 657.600 ;
        RECT 79.650 651.750 81.450 657.600 ;
        RECT 82.650 651.750 84.450 657.600 ;
        RECT 92.400 651.750 94.200 657.600 ;
        RECT 95.700 651.750 97.500 663.600 ;
        RECT 99.900 651.750 101.700 663.600 ;
        RECT 113.250 657.600 114.450 665.850 ;
        RECT 127.950 663.600 129.150 668.850 ;
        RECT 130.950 665.850 133.050 667.950 ;
        RECT 139.950 667.050 142.050 669.150 ;
        RECT 143.550 667.950 144.750 675.300 ;
        RECT 160.950 673.950 162.000 680.400 ;
        RECT 174.150 678.900 175.950 683.250 ;
        RECT 172.650 677.400 175.950 678.900 ;
        RECT 177.150 677.400 178.950 683.250 ;
        RECT 160.950 671.850 163.050 673.950 ;
        RECT 146.100 669.150 147.900 670.950 ;
        RECT 142.950 665.850 145.050 667.950 ;
        RECT 145.950 667.050 148.050 669.150 ;
        RECT 157.950 668.850 160.050 670.950 ;
        RECT 158.100 667.050 159.900 668.850 ;
        RECT 130.950 664.050 132.750 665.850 ;
        RECT 109.650 651.750 111.450 657.600 ;
        RECT 112.650 651.750 114.450 657.600 ;
        RECT 115.650 651.750 117.450 657.600 ;
        RECT 123.300 651.750 125.100 663.600 ;
        RECT 127.500 651.750 129.300 663.600 ;
        RECT 143.550 657.600 144.750 665.850 ;
        RECT 160.950 664.650 162.000 671.850 ;
        RECT 172.650 670.950 173.850 677.400 ;
        RECT 175.950 675.900 177.750 676.500 ;
        RECT 181.650 675.900 183.450 683.250 ;
        RECT 190.650 677.400 192.450 683.250 ;
        RECT 175.950 674.700 183.450 675.900 ;
        RECT 191.250 675.300 192.450 677.400 ;
        RECT 193.650 678.300 195.450 683.250 ;
        RECT 196.650 679.200 198.450 683.250 ;
        RECT 199.650 678.300 201.450 683.250 ;
        RECT 193.650 676.950 201.450 678.300 ;
        RECT 163.950 668.850 166.050 670.950 ;
        RECT 172.650 668.850 175.050 670.950 ;
        RECT 176.100 669.150 177.900 670.950 ;
        RECT 164.100 667.050 165.900 668.850 ;
        RECT 159.450 663.600 162.000 664.650 ;
        RECT 172.650 663.600 173.850 668.850 ;
        RECT 175.950 667.050 178.050 669.150 ;
        RECT 130.800 651.750 132.600 657.600 ;
        RECT 140.550 651.750 142.350 657.600 ;
        RECT 143.550 651.750 145.350 657.600 ;
        RECT 146.550 651.750 148.350 657.600 ;
        RECT 159.450 651.750 161.250 663.600 ;
        RECT 163.650 651.750 165.450 663.600 ;
        RECT 172.050 651.750 173.850 663.600 ;
        RECT 175.050 651.750 176.850 663.600 ;
        RECT 179.100 657.600 180.300 674.700 ;
        RECT 191.250 674.250 195.000 675.300 ;
        RECT 215.100 675.000 216.900 683.250 ;
        RECT 193.950 670.950 195.150 674.250 ;
        RECT 197.100 672.150 198.900 673.950 ;
        RECT 212.400 673.350 216.900 675.000 ;
        RECT 220.500 674.400 222.300 683.250 ;
        RECT 232.650 680.400 234.450 683.250 ;
        RECT 235.650 680.400 237.450 683.250 ;
        RECT 238.650 680.400 240.450 683.250 ;
        RECT 244.650 680.400 246.450 683.250 ;
        RECT 247.650 680.400 249.450 683.250 ;
        RECT 235.950 673.950 237.000 680.400 ;
        RECT 181.950 668.850 184.050 670.950 ;
        RECT 193.950 668.850 196.050 670.950 ;
        RECT 196.950 670.050 199.050 672.150 ;
        RECT 199.950 668.850 202.050 670.950 ;
        RECT 212.400 669.150 213.600 673.350 ;
        RECT 235.950 671.850 238.050 673.950 ;
        RECT 245.400 672.150 246.600 680.400 ;
        RECT 251.550 678.300 253.350 683.250 ;
        RECT 254.550 679.200 256.350 683.250 ;
        RECT 257.550 678.300 259.350 683.250 ;
        RECT 251.550 676.950 259.350 678.300 ;
        RECT 260.550 677.400 262.350 683.250 ;
        RECT 268.650 682.500 276.450 683.250 ;
        RECT 268.650 677.400 270.450 682.500 ;
        RECT 271.650 677.400 273.450 681.600 ;
        RECT 274.650 678.000 276.450 682.500 ;
        RECT 277.650 678.900 279.450 683.250 ;
        RECT 280.650 678.000 282.450 683.250 ;
        RECT 260.550 675.300 261.750 677.400 ;
        RECT 258.000 674.250 261.750 675.300 ;
        RECT 262.950 675.450 265.050 676.050 ;
        RECT 268.950 675.450 271.050 676.050 ;
        RECT 262.950 674.550 271.050 675.450 ;
        RECT 272.250 675.900 273.150 677.400 ;
        RECT 274.650 677.100 282.450 678.000 ;
        RECT 292.650 677.400 294.450 683.250 ;
        RECT 272.250 674.850 276.600 675.900 ;
        RECT 182.100 667.050 183.900 668.850 ;
        RECT 190.950 665.850 193.050 667.950 ;
        RECT 191.250 664.050 193.050 665.850 ;
        RECT 194.850 663.600 196.050 668.850 ;
        RECT 200.100 667.050 201.900 668.850 ;
        RECT 211.950 667.050 214.050 669.150 ;
        RECT 232.950 668.850 235.050 670.950 ;
        RECT 178.650 651.750 180.450 657.600 ;
        RECT 181.650 651.750 183.450 657.600 ;
        RECT 191.400 651.750 193.200 657.600 ;
        RECT 194.700 651.750 196.500 663.600 ;
        RECT 198.900 651.750 200.700 663.600 ;
        RECT 212.250 658.800 213.300 667.050 ;
        RECT 214.950 665.850 217.050 667.950 ;
        RECT 220.950 665.850 223.050 667.950 ;
        RECT 233.100 667.050 234.900 668.850 ;
        RECT 214.950 664.050 216.750 665.850 ;
        RECT 217.950 662.850 220.050 664.950 ;
        RECT 221.100 664.050 222.900 665.850 ;
        RECT 235.950 664.650 237.000 671.850 ;
        RECT 238.950 668.850 241.050 670.950 ;
        RECT 244.950 670.050 247.050 672.150 ;
        RECT 247.950 671.850 250.050 673.950 ;
        RECT 254.100 672.150 255.900 673.950 ;
        RECT 248.100 670.050 249.900 671.850 ;
        RECT 239.100 667.050 240.900 668.850 ;
        RECT 234.450 663.600 237.000 664.650 ;
        RECT 218.100 661.050 219.900 662.850 ;
        RECT 212.250 657.900 219.300 658.800 ;
        RECT 212.250 657.600 213.450 657.900 ;
        RECT 211.650 651.750 213.450 657.600 ;
        RECT 217.650 657.600 219.300 657.900 ;
        RECT 214.650 651.750 216.450 657.000 ;
        RECT 217.650 651.750 219.450 657.600 ;
        RECT 220.650 651.750 222.450 657.600 ;
        RECT 234.450 651.750 236.250 663.600 ;
        RECT 238.650 651.750 240.450 663.600 ;
        RECT 245.400 657.600 246.600 670.050 ;
        RECT 250.950 668.850 253.050 670.950 ;
        RECT 253.950 670.050 256.050 672.150 ;
        RECT 257.850 670.950 259.050 674.250 ;
        RECT 262.950 673.950 265.050 674.550 ;
        RECT 268.950 673.950 271.050 674.550 ;
        RECT 272.700 672.150 274.500 673.950 ;
        RECT 256.950 668.850 259.050 670.950 ;
        RECT 268.950 668.850 271.050 670.950 ;
        RECT 271.950 670.050 274.050 672.150 ;
        RECT 275.400 670.950 276.600 674.850 ;
        RECT 280.950 675.450 283.050 676.050 ;
        RECT 286.950 675.450 289.050 676.050 ;
        RECT 280.950 674.550 289.050 675.450 ;
        RECT 280.950 673.950 283.050 674.550 ;
        RECT 286.950 673.950 289.050 674.550 ;
        RECT 293.250 675.300 294.450 677.400 ;
        RECT 295.650 678.300 297.450 683.250 ;
        RECT 298.650 679.200 300.450 683.250 ;
        RECT 301.650 678.300 303.450 683.250 ;
        RECT 305.550 680.400 307.350 683.250 ;
        RECT 308.550 680.400 310.350 683.250 ;
        RECT 311.550 680.400 313.350 683.250 ;
        RECT 295.650 676.950 303.450 678.300 ;
        RECT 293.250 674.250 297.000 675.300 ;
        RECT 278.100 672.150 279.900 673.950 ;
        RECT 274.950 668.850 277.050 670.950 ;
        RECT 277.950 670.050 280.050 672.150 ;
        RECT 295.950 670.950 297.150 674.250 ;
        RECT 309.000 673.950 310.050 680.400 ;
        RECT 329.100 675.000 330.900 683.250 ;
        RECT 299.100 672.150 300.900 673.950 ;
        RECT 280.950 668.850 283.050 670.950 ;
        RECT 295.950 668.850 298.050 670.950 ;
        RECT 298.950 670.050 301.050 672.150 ;
        RECT 307.950 671.850 310.050 673.950 ;
        RECT 301.950 668.850 304.050 670.950 ;
        RECT 304.950 668.850 307.050 670.950 ;
        RECT 251.100 667.050 252.900 668.850 ;
        RECT 256.950 663.600 258.150 668.850 ;
        RECT 259.950 665.850 262.050 667.950 ;
        RECT 269.250 667.050 271.050 668.850 ;
        RECT 259.950 664.050 261.750 665.850 ;
        RECT 275.250 663.600 276.450 668.850 ;
        RECT 281.100 667.050 282.900 668.850 ;
        RECT 292.950 665.850 295.050 667.950 ;
        RECT 293.250 664.050 295.050 665.850 ;
        RECT 296.850 663.600 298.050 668.850 ;
        RECT 302.100 667.050 303.900 668.850 ;
        RECT 305.100 667.050 306.900 668.850 ;
        RECT 309.000 664.650 310.050 671.850 ;
        RECT 326.400 673.350 330.900 675.000 ;
        RECT 334.500 674.400 336.300 683.250 ;
        RECT 345.000 677.400 346.800 683.250 ;
        RECT 349.200 679.050 351.000 683.250 ;
        RECT 352.500 680.400 354.300 683.250 ;
        RECT 359.550 680.400 361.350 683.250 ;
        RECT 362.550 680.400 364.350 683.250 ;
        RECT 365.550 680.400 367.350 683.250 ;
        RECT 349.200 677.400 354.900 679.050 ;
        RECT 310.950 668.850 313.050 670.950 ;
        RECT 326.400 669.150 327.600 673.350 ;
        RECT 344.100 672.150 345.900 673.950 ;
        RECT 343.950 670.050 346.050 672.150 ;
        RECT 346.950 671.850 349.050 673.950 ;
        RECT 350.100 672.150 351.900 673.950 ;
        RECT 347.100 670.050 348.900 671.850 ;
        RECT 349.950 670.050 352.050 672.150 ;
        RECT 353.700 670.950 354.900 677.400 ;
        RECT 363.000 673.950 364.050 680.400 ;
        RECT 383.100 675.000 384.900 683.250 ;
        RECT 361.950 671.850 364.050 673.950 ;
        RECT 311.100 667.050 312.900 668.850 ;
        RECT 325.950 667.050 328.050 669.150 ;
        RECT 352.950 668.850 355.050 670.950 ;
        RECT 358.950 668.850 361.050 670.950 ;
        RECT 309.000 663.600 311.550 664.650 ;
        RECT 244.650 651.750 246.450 657.600 ;
        RECT 247.650 651.750 249.450 657.600 ;
        RECT 252.300 651.750 254.100 663.600 ;
        RECT 256.500 651.750 258.300 663.600 ;
        RECT 259.800 651.750 261.600 657.600 ;
        RECT 270.150 651.750 271.950 663.600 ;
        RECT 274.650 651.750 277.950 663.600 ;
        RECT 280.650 651.750 282.450 663.600 ;
        RECT 293.400 651.750 295.200 657.600 ;
        RECT 296.700 651.750 298.500 663.600 ;
        RECT 300.900 651.750 302.700 663.600 ;
        RECT 305.550 651.750 307.350 663.600 ;
        RECT 309.750 651.750 311.550 663.600 ;
        RECT 326.250 658.800 327.300 667.050 ;
        RECT 328.950 665.850 331.050 667.950 ;
        RECT 334.950 665.850 337.050 667.950 ;
        RECT 328.950 664.050 330.750 665.850 ;
        RECT 331.950 662.850 334.050 664.950 ;
        RECT 335.100 664.050 336.900 665.850 ;
        RECT 353.700 663.600 354.900 668.850 ;
        RECT 359.100 667.050 360.900 668.850 ;
        RECT 363.000 664.650 364.050 671.850 ;
        RECT 380.400 673.350 384.900 675.000 ;
        RECT 388.500 674.400 390.300 683.250 ;
        RECT 398.700 680.400 400.500 683.250 ;
        RECT 402.000 679.050 403.800 683.250 ;
        RECT 398.100 677.400 403.800 679.050 ;
        RECT 406.200 677.400 408.000 683.250 ;
        RECT 418.650 680.400 420.450 683.250 ;
        RECT 421.650 680.400 423.450 683.250 ;
        RECT 364.950 668.850 367.050 670.950 ;
        RECT 380.400 669.150 381.600 673.350 ;
        RECT 398.100 670.950 399.300 677.400 ;
        RECT 401.100 672.150 402.900 673.950 ;
        RECT 365.100 667.050 366.900 668.850 ;
        RECT 379.950 667.050 382.050 669.150 ;
        RECT 397.950 668.850 400.050 670.950 ;
        RECT 400.950 670.050 403.050 672.150 ;
        RECT 403.950 671.850 406.050 673.950 ;
        RECT 407.100 672.150 408.900 673.950 ;
        RECT 419.400 672.150 420.600 680.400 ;
        RECT 435.150 678.900 436.950 683.250 ;
        RECT 433.650 677.400 436.950 678.900 ;
        RECT 438.150 677.400 439.950 683.250 ;
        RECT 404.100 670.050 405.900 671.850 ;
        RECT 406.950 670.050 409.050 672.150 ;
        RECT 418.950 670.050 421.050 672.150 ;
        RECT 421.950 671.850 424.050 673.950 ;
        RECT 422.100 670.050 423.900 671.850 ;
        RECT 433.650 670.950 434.850 677.400 ;
        RECT 436.950 675.900 438.750 676.500 ;
        RECT 442.650 675.900 444.450 683.250 ;
        RECT 451.650 677.400 453.450 683.250 ;
        RECT 436.950 674.700 444.450 675.900 ;
        RECT 452.250 675.300 453.450 677.400 ;
        RECT 454.650 678.300 456.450 683.250 ;
        RECT 457.650 679.200 459.450 683.250 ;
        RECT 460.650 678.300 462.450 683.250 ;
        RECT 454.650 676.950 462.450 678.300 ;
        RECT 468.000 677.400 469.800 683.250 ;
        RECT 472.200 677.400 474.000 683.250 ;
        RECT 476.400 677.400 478.200 683.250 ;
        RECT 488.550 678.000 490.350 683.250 ;
        RECT 491.550 678.900 493.350 683.250 ;
        RECT 494.550 682.500 502.350 683.250 ;
        RECT 494.550 678.000 496.350 682.500 ;
        RECT 363.000 663.600 365.550 664.650 ;
        RECT 332.100 661.050 333.900 662.850 ;
        RECT 344.550 662.700 352.350 663.600 ;
        RECT 326.250 657.900 333.300 658.800 ;
        RECT 326.250 657.600 327.450 657.900 ;
        RECT 325.650 651.750 327.450 657.600 ;
        RECT 331.650 657.600 333.300 657.900 ;
        RECT 328.650 651.750 330.450 657.000 ;
        RECT 331.650 651.750 333.450 657.600 ;
        RECT 334.650 651.750 336.450 657.600 ;
        RECT 344.550 651.750 346.350 662.700 ;
        RECT 347.550 651.750 349.350 661.800 ;
        RECT 350.550 651.750 352.350 662.700 ;
        RECT 353.550 651.750 355.350 663.600 ;
        RECT 359.550 651.750 361.350 663.600 ;
        RECT 363.750 651.750 365.550 663.600 ;
        RECT 380.250 658.800 381.300 667.050 ;
        RECT 382.950 665.850 385.050 667.950 ;
        RECT 388.950 665.850 391.050 667.950 ;
        RECT 382.950 664.050 384.750 665.850 ;
        RECT 385.950 662.850 388.050 664.950 ;
        RECT 389.100 664.050 390.900 665.850 ;
        RECT 398.100 663.600 399.300 668.850 ;
        RECT 386.100 661.050 387.900 662.850 ;
        RECT 380.250 657.900 387.300 658.800 ;
        RECT 380.250 657.600 381.450 657.900 ;
        RECT 379.650 651.750 381.450 657.600 ;
        RECT 385.650 657.600 387.300 657.900 ;
        RECT 382.650 651.750 384.450 657.000 ;
        RECT 385.650 651.750 387.450 657.600 ;
        RECT 388.650 651.750 390.450 657.600 ;
        RECT 397.650 651.750 399.450 663.600 ;
        RECT 400.650 662.700 408.450 663.600 ;
        RECT 400.650 651.750 402.450 662.700 ;
        RECT 403.650 651.750 405.450 661.800 ;
        RECT 406.650 651.750 408.450 662.700 ;
        RECT 419.400 657.600 420.600 670.050 ;
        RECT 433.650 668.850 436.050 670.950 ;
        RECT 437.100 669.150 438.900 670.950 ;
        RECT 433.650 663.600 434.850 668.850 ;
        RECT 436.950 667.050 439.050 669.150 ;
        RECT 418.650 651.750 420.450 657.600 ;
        RECT 421.650 651.750 423.450 657.600 ;
        RECT 433.050 651.750 434.850 663.600 ;
        RECT 436.050 651.750 437.850 663.600 ;
        RECT 440.100 657.600 441.300 674.700 ;
        RECT 452.250 674.250 456.000 675.300 ;
        RECT 454.950 670.950 456.150 674.250 ;
        RECT 458.100 672.150 459.900 673.950 ;
        RECT 470.250 672.150 472.050 673.950 ;
        RECT 442.950 668.850 445.050 670.950 ;
        RECT 454.950 668.850 457.050 670.950 ;
        RECT 457.950 670.050 460.050 672.150 ;
        RECT 460.950 668.850 463.050 670.950 ;
        RECT 466.950 668.850 469.050 670.950 ;
        RECT 469.950 670.050 472.050 672.150 ;
        RECT 472.950 670.950 474.000 677.400 ;
        RECT 488.550 677.100 496.350 678.000 ;
        RECT 497.550 677.400 499.350 681.600 ;
        RECT 500.550 677.400 502.350 682.500 ;
        RECT 511.650 680.400 513.450 683.250 ;
        RECT 514.650 680.400 516.450 683.250 ;
        RECT 523.650 680.400 525.450 683.250 ;
        RECT 526.650 680.400 528.450 683.250 ;
        RECT 529.650 680.400 531.450 683.250 ;
        RECT 497.850 675.900 498.750 677.400 ;
        RECT 494.400 674.850 498.750 675.900 ;
        RECT 475.950 672.150 477.750 673.950 ;
        RECT 491.100 672.150 492.900 673.950 ;
        RECT 472.950 668.850 475.050 670.950 ;
        RECT 475.950 670.050 478.050 672.150 ;
        RECT 478.950 668.850 481.050 670.950 ;
        RECT 487.950 668.850 490.050 670.950 ;
        RECT 490.950 670.050 493.050 672.150 ;
        RECT 494.400 670.950 495.600 674.850 ;
        RECT 496.500 672.150 498.300 673.950 ;
        RECT 512.400 672.150 513.600 680.400 ;
        RECT 523.950 675.450 526.050 676.050 ;
        RECT 518.550 674.550 526.050 675.450 ;
        RECT 493.950 668.850 496.050 670.950 ;
        RECT 496.950 670.050 499.050 672.150 ;
        RECT 499.950 668.850 502.050 670.950 ;
        RECT 511.950 670.050 514.050 672.150 ;
        RECT 514.950 671.850 517.050 673.950 ;
        RECT 515.100 670.050 516.900 671.850 ;
        RECT 443.100 667.050 444.900 668.850 ;
        RECT 451.950 665.850 454.050 667.950 ;
        RECT 452.250 664.050 454.050 665.850 ;
        RECT 455.850 663.600 457.050 668.850 ;
        RECT 461.100 667.050 462.900 668.850 ;
        RECT 467.250 667.050 469.050 668.850 ;
        RECT 474.150 665.400 475.050 668.850 ;
        RECT 479.100 667.050 480.900 668.850 ;
        RECT 488.100 667.050 489.900 668.850 ;
        RECT 474.150 664.500 478.200 665.400 ;
        RECT 476.400 663.600 478.200 664.500 ;
        RECT 494.550 663.600 495.750 668.850 ;
        RECT 499.950 667.050 501.750 668.850 ;
        RECT 439.650 651.750 441.450 657.600 ;
        RECT 442.650 651.750 444.450 657.600 ;
        RECT 452.400 651.750 454.200 657.600 ;
        RECT 455.700 651.750 457.500 663.600 ;
        RECT 459.900 651.750 461.700 663.600 ;
        RECT 467.550 662.400 475.350 663.300 ;
        RECT 467.550 651.750 469.350 662.400 ;
        RECT 470.550 651.750 472.350 661.500 ;
        RECT 473.550 652.500 475.350 662.400 ;
        RECT 476.550 653.400 478.350 663.600 ;
        RECT 479.550 652.500 481.350 663.600 ;
        RECT 473.550 651.750 481.350 652.500 ;
        RECT 488.550 651.750 490.350 663.600 ;
        RECT 493.050 651.750 496.350 663.600 ;
        RECT 499.050 651.750 500.850 663.600 ;
        RECT 512.400 657.600 513.600 670.050 ;
        RECT 514.950 666.450 517.050 667.050 ;
        RECT 518.550 666.450 519.450 674.550 ;
        RECT 523.950 673.950 526.050 674.550 ;
        RECT 526.950 673.950 528.000 680.400 ;
        RECT 535.650 677.400 537.450 683.250 ;
        RECT 529.950 675.450 532.050 676.050 ;
        RECT 529.950 674.550 534.450 675.450 ;
        RECT 529.950 673.950 532.050 674.550 ;
        RECT 526.950 671.850 529.050 673.950 ;
        RECT 523.950 668.850 526.050 670.950 ;
        RECT 524.100 667.050 525.900 668.850 ;
        RECT 514.950 665.550 519.450 666.450 ;
        RECT 514.950 664.950 517.050 665.550 ;
        RECT 526.950 664.650 528.000 671.850 ;
        RECT 529.950 668.850 532.050 670.950 ;
        RECT 530.100 667.050 531.900 668.850 ;
        RECT 525.450 663.600 528.000 664.650 ;
        RECT 511.650 651.750 513.450 657.600 ;
        RECT 514.650 651.750 516.450 657.600 ;
        RECT 525.450 651.750 527.250 663.600 ;
        RECT 529.650 651.750 531.450 663.600 ;
        RECT 533.550 661.050 534.450 674.550 ;
        RECT 536.250 675.300 537.450 677.400 ;
        RECT 538.650 678.300 540.450 683.250 ;
        RECT 541.650 679.200 543.450 683.250 ;
        RECT 544.650 678.300 546.450 683.250 ;
        RECT 554.550 680.400 556.350 683.250 ;
        RECT 557.550 680.400 559.350 683.250 ;
        RECT 560.550 680.400 562.350 683.250 ;
        RECT 569.550 680.400 571.350 683.250 ;
        RECT 572.550 680.400 574.350 683.250 ;
        RECT 575.550 680.400 577.350 683.250 ;
        RECT 586.650 680.400 588.450 683.250 ;
        RECT 589.650 680.400 591.450 683.250 ;
        RECT 592.650 680.400 594.450 683.250 ;
        RECT 599.550 680.400 601.350 683.250 ;
        RECT 602.550 680.400 604.350 683.250 ;
        RECT 605.550 680.400 607.350 683.250 ;
        RECT 538.650 676.950 546.450 678.300 ;
        RECT 544.950 675.450 547.050 676.050 ;
        RECT 553.950 675.450 556.050 676.050 ;
        RECT 536.250 674.250 540.000 675.300 ;
        RECT 544.950 674.550 556.050 675.450 ;
        RECT 538.950 670.950 540.150 674.250 ;
        RECT 544.950 673.950 547.050 674.550 ;
        RECT 553.950 673.950 556.050 674.550 ;
        RECT 558.000 673.950 559.050 680.400 ;
        RECT 573.000 673.950 574.050 680.400 ;
        RECT 542.100 672.150 543.900 673.950 ;
        RECT 538.950 668.850 541.050 670.950 ;
        RECT 541.950 670.050 544.050 672.150 ;
        RECT 556.950 671.850 559.050 673.950 ;
        RECT 571.950 671.850 574.050 673.950 ;
        RECT 544.950 668.850 547.050 670.950 ;
        RECT 553.950 668.850 556.050 670.950 ;
        RECT 535.950 665.850 538.050 667.950 ;
        RECT 536.250 664.050 538.050 665.850 ;
        RECT 539.850 663.600 541.050 668.850 ;
        RECT 545.100 667.050 546.900 668.850 ;
        RECT 554.100 667.050 555.900 668.850 ;
        RECT 558.000 664.650 559.050 671.850 ;
        RECT 559.950 668.850 562.050 670.950 ;
        RECT 568.950 668.850 571.050 670.950 ;
        RECT 560.100 667.050 561.900 668.850 ;
        RECT 569.100 667.050 570.900 668.850 ;
        RECT 573.000 664.650 574.050 671.850 ;
        RECT 589.950 673.950 591.000 680.400 ;
        RECT 603.000 673.950 604.050 680.400 ;
        RECT 616.650 677.400 618.450 683.250 ;
        RECT 617.250 675.300 618.450 677.400 ;
        RECT 619.650 678.300 621.450 683.250 ;
        RECT 622.650 679.200 624.450 683.250 ;
        RECT 625.650 678.300 627.450 683.250 ;
        RECT 619.650 676.950 627.450 678.300 ;
        RECT 634.650 677.400 636.450 683.250 ;
        RECT 635.250 675.300 636.450 677.400 ;
        RECT 637.650 678.300 639.450 683.250 ;
        RECT 640.650 679.200 642.450 683.250 ;
        RECT 643.650 678.300 645.450 683.250 ;
        RECT 648.750 680.400 650.550 683.250 ;
        RECT 651.750 680.400 653.550 683.250 ;
        RECT 637.650 676.950 645.450 678.300 ;
        RECT 617.250 674.250 621.000 675.300 ;
        RECT 635.250 674.250 639.000 675.300 ;
        RECT 589.950 671.850 592.050 673.950 ;
        RECT 601.950 671.850 604.050 673.950 ;
        RECT 574.950 668.850 577.050 670.950 ;
        RECT 586.950 668.850 589.050 670.950 ;
        RECT 575.100 667.050 576.900 668.850 ;
        RECT 587.100 667.050 588.900 668.850 ;
        RECT 589.950 664.650 591.000 671.850 ;
        RECT 592.950 668.850 595.050 670.950 ;
        RECT 598.950 668.850 601.050 670.950 ;
        RECT 593.100 667.050 594.900 668.850 ;
        RECT 599.100 667.050 600.900 668.850 ;
        RECT 558.000 663.600 560.550 664.650 ;
        RECT 573.000 663.600 575.550 664.650 ;
        RECT 532.950 658.950 535.050 661.050 ;
        RECT 536.400 651.750 538.200 657.600 ;
        RECT 539.700 651.750 541.500 663.600 ;
        RECT 543.900 651.750 545.700 663.600 ;
        RECT 554.550 651.750 556.350 663.600 ;
        RECT 558.750 651.750 560.550 663.600 ;
        RECT 569.550 651.750 571.350 663.600 ;
        RECT 573.750 651.750 575.550 663.600 ;
        RECT 588.450 663.600 591.000 664.650 ;
        RECT 603.000 664.650 604.050 671.850 ;
        RECT 619.950 670.950 621.150 674.250 ;
        RECT 623.100 672.150 624.900 673.950 ;
        RECT 604.950 668.850 607.050 670.950 ;
        RECT 619.950 668.850 622.050 670.950 ;
        RECT 622.950 670.050 625.050 672.150 ;
        RECT 637.950 670.950 639.150 674.250 ;
        RECT 641.100 672.150 642.900 673.950 ;
        RECT 652.050 672.150 653.550 680.400 ;
        RECT 625.950 668.850 628.050 670.950 ;
        RECT 637.950 668.850 640.050 670.950 ;
        RECT 640.950 670.050 643.050 672.150 ;
        RECT 643.950 668.850 646.050 670.950 ;
        RECT 649.950 670.050 653.550 672.150 ;
        RECT 605.100 667.050 606.900 668.850 ;
        RECT 616.950 665.850 619.050 667.950 ;
        RECT 603.000 663.600 605.550 664.650 ;
        RECT 617.250 664.050 619.050 665.850 ;
        RECT 620.850 663.600 622.050 668.850 ;
        RECT 626.100 667.050 627.900 668.850 ;
        RECT 634.950 665.850 637.050 667.950 ;
        RECT 635.250 664.050 637.050 665.850 ;
        RECT 638.850 663.600 640.050 668.850 ;
        RECT 644.100 667.050 645.900 668.850 ;
        RECT 588.450 651.750 590.250 663.600 ;
        RECT 592.650 651.750 594.450 663.600 ;
        RECT 599.550 651.750 601.350 663.600 ;
        RECT 603.750 651.750 605.550 663.600 ;
        RECT 617.400 651.750 619.200 657.600 ;
        RECT 620.700 651.750 622.500 663.600 ;
        RECT 624.900 651.750 626.700 663.600 ;
        RECT 635.400 651.750 637.200 657.600 ;
        RECT 638.700 651.750 640.500 663.600 ;
        RECT 642.900 651.750 644.700 663.600 ;
        RECT 652.050 657.600 653.550 670.050 ;
        RECT 655.650 677.400 657.450 683.250 ;
        RECT 661.050 677.400 662.850 683.250 ;
        RECT 666.600 678.600 668.400 683.250 ;
        RECT 671.250 679.500 673.050 683.250 ;
        RECT 674.250 679.500 676.050 683.250 ;
        RECT 677.250 679.500 679.050 683.250 ;
        RECT 664.200 677.400 668.400 678.600 ;
        RECT 670.950 677.400 673.050 679.500 ;
        RECT 673.950 677.400 676.050 679.500 ;
        RECT 676.950 677.400 679.050 679.500 ;
        RECT 681.000 679.500 682.800 683.250 ;
        RECT 684.000 680.400 685.800 683.250 ;
        RECT 687.000 679.500 688.800 683.250 ;
        RECT 691.500 680.400 693.300 683.250 ;
        RECT 694.500 680.400 696.300 683.250 ;
        RECT 697.500 680.400 699.300 683.250 ;
        RECT 700.500 680.400 702.300 683.250 ;
        RECT 681.000 677.700 683.850 679.500 ;
        RECT 681.750 677.400 683.850 677.700 ;
        RECT 685.950 677.700 688.800 679.500 ;
        RECT 689.700 678.750 691.500 679.200 ;
        RECT 694.950 679.050 696.300 680.400 ;
        RECT 697.950 679.050 699.300 680.400 ;
        RECT 700.950 679.050 702.300 680.400 ;
        RECT 685.950 677.400 688.050 677.700 ;
        RECT 689.700 677.400 693.750 678.750 ;
        RECT 655.650 662.550 656.850 677.400 ;
        RECT 664.200 673.800 665.700 677.400 ;
        RECT 670.350 674.700 677.100 676.500 ;
        RECT 678.000 674.700 684.900 676.500 ;
        RECT 692.850 676.050 693.750 677.400 ;
        RECT 694.950 676.950 697.050 679.050 ;
        RECT 697.950 676.950 700.050 679.050 ;
        RECT 700.950 676.950 703.050 679.050 ;
        RECT 692.850 675.900 697.950 676.050 ;
        RECT 692.850 675.150 700.500 675.900 ;
        RECT 696.150 674.700 700.500 675.150 ;
        RECT 678.000 673.800 679.050 674.700 ;
        RECT 696.150 674.250 697.950 674.700 ;
        RECT 657.900 672.000 665.700 673.800 ;
        RECT 669.150 672.750 679.050 673.800 ;
        RECT 669.150 670.950 670.200 672.750 ;
        RECT 679.950 672.450 687.600 673.800 ;
        RECT 679.950 671.700 680.850 672.450 ;
        RECT 661.950 669.900 670.200 670.950 ;
        RECT 671.250 670.650 680.850 671.700 ;
        RECT 661.950 665.850 664.050 669.900 ;
        RECT 671.250 669.000 672.150 670.650 ;
        RECT 681.750 669.750 685.650 671.550 ;
        RECT 686.550 670.950 687.600 672.450 ;
        RECT 688.950 673.650 691.050 673.950 ;
        RECT 688.950 671.850 692.850 673.650 ;
        RECT 699.450 671.250 700.500 674.700 ;
        RECT 702.000 673.800 703.050 676.950 ;
        RECT 704.700 677.400 706.500 683.250 ;
        RECT 710.100 677.400 711.900 683.250 ;
        RECT 715.500 677.400 717.300 683.250 ;
        RECT 722.850 677.400 724.650 683.250 ;
        RECT 704.700 676.500 706.200 677.400 ;
        RECT 704.700 675.300 713.100 676.500 ;
        RECT 711.300 674.700 713.100 675.300 ;
        RECT 716.100 673.800 717.300 677.400 ;
        RECT 727.350 676.200 729.150 683.250 ;
        RECT 734.550 677.400 736.350 683.250 ;
        RECT 737.550 677.400 739.350 683.250 ;
        RECT 740.550 677.400 742.350 683.250 ;
        RECT 702.000 672.900 717.300 673.800 ;
        RECT 686.550 670.050 698.550 670.950 ;
        RECT 665.100 667.200 672.150 669.000 ;
        RECT 673.500 667.950 675.300 669.750 ;
        RECT 681.750 669.450 683.850 669.750 ;
        RECT 685.950 668.550 688.050 668.850 ;
        RECT 694.800 668.550 696.600 669.150 ;
        RECT 685.950 667.950 696.600 668.550 ;
        RECT 673.500 667.350 696.600 667.950 ;
        RECT 697.500 668.550 698.550 670.050 ;
        RECT 699.450 669.450 701.250 671.250 ;
        RECT 703.050 670.950 714.900 672.000 ;
        RECT 703.050 668.550 704.250 670.950 ;
        RECT 713.100 669.150 714.900 670.950 ;
        RECT 697.500 667.650 704.250 668.550 ;
        RECT 706.950 667.650 709.050 667.950 ;
        RECT 673.500 666.750 688.050 667.350 ;
        RECT 705.150 666.450 709.050 667.650 ;
        RECT 712.950 667.050 715.050 669.150 ;
        RECT 695.100 665.850 709.050 666.450 ;
        RECT 669.000 665.550 708.750 665.850 ;
        RECT 657.750 664.650 659.550 665.250 ;
        RECT 669.000 664.650 697.050 665.550 ;
        RECT 657.750 663.450 670.050 664.650 ;
        RECT 697.950 664.050 700.050 664.350 ;
        RECT 707.700 664.050 709.500 664.650 ;
        RECT 670.950 662.550 673.050 663.750 ;
        RECT 655.650 661.650 673.050 662.550 ;
        RECT 676.950 662.400 697.050 663.750 ;
        RECT 676.950 661.650 679.050 662.400 ;
        RECT 658.500 657.600 659.700 661.650 ;
        RECT 660.600 659.700 662.400 660.300 ;
        RECT 667.350 660.150 669.150 660.300 ;
        RECT 660.600 658.500 666.300 659.700 ;
        RECT 667.350 658.950 676.050 660.150 ;
        RECT 667.350 658.500 669.150 658.950 ;
        RECT 648.750 651.750 650.550 657.600 ;
        RECT 651.750 651.750 653.550 657.600 ;
        RECT 655.500 651.750 657.300 657.600 ;
        RECT 658.500 651.750 660.300 657.600 ;
        RECT 661.500 651.750 663.300 657.600 ;
        RECT 664.500 651.750 666.300 658.500 ;
        RECT 673.950 658.050 676.050 658.950 ;
        RECT 667.500 651.750 669.300 657.600 ;
        RECT 670.800 655.800 672.900 657.900 ;
        RECT 671.400 654.600 672.900 655.800 ;
        RECT 671.250 651.750 673.050 654.600 ;
        RECT 674.250 651.750 676.050 658.050 ;
        RECT 677.550 654.600 678.900 661.650 ;
        RECT 695.100 661.350 697.050 662.400 ;
        RECT 697.950 662.850 709.500 664.050 ;
        RECT 697.950 662.250 700.050 662.850 ;
        RECT 711.000 661.350 712.800 662.100 ;
        RECT 680.100 658.800 684.000 660.600 ;
        RECT 681.000 658.500 684.000 658.800 ;
        RECT 685.950 660.150 688.050 660.600 ;
        RECT 695.100 660.300 712.800 661.350 ;
        RECT 685.950 658.500 688.350 660.150 ;
        RECT 677.250 651.750 679.050 654.600 ;
        RECT 681.000 651.750 682.800 658.500 ;
        RECT 687.000 657.600 688.350 658.500 ;
        RECT 694.950 657.600 697.050 658.050 ;
        RECT 684.000 651.750 685.800 657.600 ;
        RECT 687.000 651.750 688.800 657.600 ;
        RECT 690.750 651.750 692.550 657.600 ;
        RECT 694.500 655.950 697.050 657.600 ;
        RECT 697.950 655.950 700.050 658.050 ;
        RECT 700.950 655.950 703.050 658.050 ;
        RECT 694.500 654.600 695.700 655.950 ;
        RECT 697.950 654.600 698.850 655.950 ;
        RECT 700.950 654.600 702.150 655.950 ;
        RECT 693.750 651.750 695.700 654.600 ;
        RECT 696.750 651.750 698.850 654.600 ;
        RECT 699.750 651.750 702.150 654.600 ;
        RECT 703.500 651.750 705.300 655.050 ;
        RECT 706.500 651.750 708.300 660.300 ;
        RECT 716.100 659.400 717.300 672.900 ;
        RECT 725.550 675.300 729.150 676.200 ;
        RECT 737.400 676.500 739.200 677.400 ;
        RECT 743.550 676.500 745.350 683.250 ;
        RECT 746.550 677.400 748.350 683.250 ;
        RECT 749.550 677.400 751.350 683.250 ;
        RECT 752.550 677.400 754.350 683.250 ;
        RECT 755.550 677.400 757.350 683.250 ;
        RECT 758.550 677.400 760.350 683.250 ;
        RECT 769.650 677.400 771.450 683.250 ;
        RECT 749.400 676.500 751.200 677.400 ;
        RECT 755.400 676.500 757.200 677.400 ;
        RECT 737.400 675.300 741.450 676.500 ;
        RECT 743.550 675.300 747.300 676.500 ;
        RECT 749.400 675.300 753.300 676.500 ;
        RECT 755.400 676.350 758.100 676.500 ;
        RECT 755.400 675.300 758.250 676.350 ;
        RECT 722.100 669.150 723.900 670.950 ;
        RECT 721.950 667.050 724.050 669.150 ;
        RECT 725.550 667.950 726.750 675.300 ;
        RECT 740.250 674.400 741.450 675.300 ;
        RECT 746.100 674.400 747.300 675.300 ;
        RECT 752.100 674.400 753.300 675.300 ;
        RECT 737.100 672.150 738.900 673.950 ;
        RECT 740.250 672.600 744.300 674.400 ;
        RECT 746.100 672.600 750.300 674.400 ;
        RECT 752.100 672.600 756.300 674.400 ;
        RECT 728.100 669.150 729.900 670.950 ;
        RECT 736.950 670.050 739.050 672.150 ;
        RECT 724.950 665.850 727.050 667.950 ;
        RECT 727.950 667.050 730.050 669.150 ;
        RECT 713.250 658.500 717.300 659.400 ;
        RECT 713.250 657.600 714.300 658.500 ;
        RECT 725.550 657.600 726.750 665.850 ;
        RECT 740.250 665.700 741.450 672.600 ;
        RECT 746.100 665.700 747.300 672.600 ;
        RECT 752.100 665.700 753.300 672.600 ;
        RECT 757.200 672.150 758.250 675.300 ;
        RECT 770.250 675.300 771.450 677.400 ;
        RECT 772.650 678.300 774.450 683.250 ;
        RECT 775.650 679.200 777.450 683.250 ;
        RECT 778.650 678.300 780.450 683.250 ;
        RECT 785.550 680.400 787.350 683.250 ;
        RECT 788.550 680.400 790.350 683.250 ;
        RECT 797.550 680.400 799.350 683.250 ;
        RECT 800.550 680.400 802.350 683.250 ;
        RECT 803.550 680.400 805.350 683.250 ;
        RECT 772.650 676.950 780.450 678.300 ;
        RECT 770.250 674.250 774.000 675.300 ;
        RECT 757.200 670.050 760.050 672.150 ;
        RECT 772.950 670.950 774.150 674.250 ;
        RECT 776.100 672.150 777.900 673.950 ;
        RECT 757.200 665.700 758.250 670.050 ;
        RECT 772.950 668.850 775.050 670.950 ;
        RECT 775.950 670.050 778.050 672.150 ;
        RECT 784.950 671.850 787.050 673.950 ;
        RECT 788.400 672.150 789.600 680.400 ;
        RECT 801.450 676.200 802.350 680.400 ;
        RECT 806.550 677.400 808.350 683.250 ;
        RECT 815.550 678.300 817.350 683.250 ;
        RECT 818.550 679.200 820.350 683.250 ;
        RECT 821.550 678.300 823.350 683.250 ;
        RECT 801.450 675.300 804.750 676.200 ;
        RECT 802.950 674.400 804.750 675.300 ;
        RECT 778.950 668.850 781.050 670.950 ;
        RECT 785.100 670.050 786.900 671.850 ;
        RECT 787.950 670.050 790.050 672.150 ;
        RECT 796.950 671.850 799.050 673.950 ;
        RECT 797.100 670.050 798.900 671.850 ;
        RECT 769.950 665.850 772.050 667.950 ;
        RECT 737.550 664.500 741.450 665.700 ;
        RECT 743.550 664.500 747.300 665.700 ;
        RECT 749.550 664.500 753.300 665.700 ;
        RECT 755.550 664.500 758.250 665.700 ;
        RECT 709.500 651.750 711.300 657.600 ;
        RECT 712.500 651.750 714.300 657.600 ;
        RECT 715.500 651.750 717.300 657.600 ;
        RECT 722.550 651.750 724.350 657.600 ;
        RECT 725.550 651.750 727.350 657.600 ;
        RECT 728.550 651.750 730.350 657.600 ;
        RECT 734.550 651.750 736.350 663.600 ;
        RECT 737.550 651.750 739.350 664.500 ;
        RECT 740.550 651.750 742.350 663.600 ;
        RECT 743.550 651.750 745.350 664.500 ;
        RECT 746.550 651.750 748.350 663.600 ;
        RECT 749.550 651.750 751.350 664.500 ;
        RECT 752.550 651.750 754.350 663.600 ;
        RECT 755.550 651.750 757.350 664.500 ;
        RECT 770.250 664.050 772.050 665.850 ;
        RECT 773.850 663.600 775.050 668.850 ;
        RECT 779.100 667.050 780.900 668.850 ;
        RECT 758.550 651.750 760.350 663.600 ;
        RECT 770.400 651.750 772.200 657.600 ;
        RECT 773.700 651.750 775.500 663.600 ;
        RECT 777.900 651.750 779.700 663.600 ;
        RECT 788.400 657.600 789.600 670.050 ;
        RECT 799.950 668.850 802.050 670.950 ;
        RECT 800.100 667.050 801.900 668.850 ;
        RECT 803.700 666.150 804.600 674.400 ;
        RECT 807.000 672.150 808.050 677.400 ;
        RECT 815.550 676.950 823.350 678.300 ;
        RECT 824.550 677.400 826.350 683.250 ;
        RECT 833.550 678.300 835.350 683.250 ;
        RECT 836.550 679.200 838.350 683.250 ;
        RECT 839.550 678.300 841.350 683.250 ;
        RECT 808.950 675.450 811.050 676.050 ;
        RECT 814.950 675.450 817.050 676.050 ;
        RECT 808.950 674.550 817.050 675.450 ;
        RECT 824.550 675.300 825.750 677.400 ;
        RECT 833.550 676.950 841.350 678.300 ;
        RECT 842.550 677.400 844.350 683.250 ;
        RECT 842.550 675.300 843.750 677.400 ;
        RECT 808.950 673.950 811.050 674.550 ;
        RECT 814.950 673.950 817.050 674.550 ;
        RECT 822.000 674.250 825.750 675.300 ;
        RECT 840.000 674.250 843.750 675.300 ;
        RECT 818.100 672.150 819.900 673.950 ;
        RECT 805.950 670.050 808.050 672.150 ;
        RECT 802.950 666.000 804.750 666.150 ;
        RECT 797.550 664.800 804.750 666.000 ;
        RECT 797.550 663.600 798.750 664.800 ;
        RECT 802.950 664.350 804.750 664.800 ;
        RECT 785.550 651.750 787.350 657.600 ;
        RECT 788.550 651.750 790.350 657.600 ;
        RECT 797.550 651.750 799.350 663.600 ;
        RECT 806.100 663.450 807.450 670.050 ;
        RECT 814.950 668.850 817.050 670.950 ;
        RECT 817.950 670.050 820.050 672.150 ;
        RECT 821.850 670.950 823.050 674.250 ;
        RECT 836.100 672.150 837.900 673.950 ;
        RECT 820.950 668.850 823.050 670.950 ;
        RECT 832.950 668.850 835.050 670.950 ;
        RECT 835.950 670.050 838.050 672.150 ;
        RECT 839.850 670.950 841.050 674.250 ;
        RECT 838.950 668.850 841.050 670.950 ;
        RECT 815.100 667.050 816.900 668.850 ;
        RECT 820.950 663.600 822.150 668.850 ;
        RECT 823.950 665.850 826.050 667.950 ;
        RECT 833.100 667.050 834.900 668.850 ;
        RECT 823.950 664.050 825.750 665.850 ;
        RECT 838.950 663.600 840.150 668.850 ;
        RECT 841.950 665.850 844.050 667.950 ;
        RECT 841.950 664.050 843.750 665.850 ;
        RECT 802.050 651.750 803.850 663.450 ;
        RECT 805.050 662.100 807.450 663.450 ;
        RECT 805.050 651.750 806.850 662.100 ;
        RECT 816.300 651.750 818.100 663.600 ;
        RECT 820.500 651.750 822.300 663.600 ;
        RECT 823.800 651.750 825.600 657.600 ;
        RECT 834.300 651.750 836.100 663.600 ;
        RECT 838.500 651.750 840.300 663.600 ;
        RECT 841.800 651.750 843.600 657.600 ;
        RECT 2.700 641.400 4.500 647.250 ;
        RECT 5.700 641.400 7.500 647.250 ;
        RECT 8.700 641.400 10.500 647.250 ;
        RECT 5.700 640.500 6.750 641.400 ;
        RECT 2.700 639.600 6.750 640.500 ;
        RECT 2.700 626.100 3.900 639.600 ;
        RECT 11.700 638.700 13.500 647.250 ;
        RECT 14.700 643.950 16.500 647.250 ;
        RECT 17.850 644.400 20.250 647.250 ;
        RECT 21.150 644.400 23.250 647.250 ;
        RECT 24.300 644.400 26.250 647.250 ;
        RECT 17.850 643.050 19.050 644.400 ;
        RECT 21.150 643.050 22.050 644.400 ;
        RECT 24.300 643.050 25.500 644.400 ;
        RECT 16.950 640.950 19.050 643.050 ;
        RECT 19.950 640.950 22.050 643.050 ;
        RECT 22.950 641.400 25.500 643.050 ;
        RECT 27.450 641.400 29.250 647.250 ;
        RECT 31.200 641.400 33.000 647.250 ;
        RECT 34.200 641.400 36.000 647.250 ;
        RECT 22.950 640.950 25.050 641.400 ;
        RECT 31.650 640.500 33.000 641.400 ;
        RECT 37.200 640.500 39.000 647.250 ;
        RECT 40.950 644.400 42.750 647.250 ;
        RECT 31.650 638.850 34.050 640.500 ;
        RECT 7.200 637.650 24.900 638.700 ;
        RECT 31.950 638.400 34.050 638.850 ;
        RECT 36.000 640.200 39.000 640.500 ;
        RECT 36.000 638.400 39.900 640.200 ;
        RECT 7.200 636.900 9.000 637.650 ;
        RECT 19.950 636.150 22.050 636.750 ;
        RECT 10.500 634.950 22.050 636.150 ;
        RECT 22.950 636.600 24.900 637.650 ;
        RECT 41.100 637.350 42.450 644.400 ;
        RECT 43.950 640.950 45.750 647.250 ;
        RECT 46.950 644.400 48.750 647.250 ;
        RECT 47.100 643.200 48.600 644.400 ;
        RECT 47.100 641.100 49.200 643.200 ;
        RECT 50.700 641.400 52.500 647.250 ;
        RECT 43.950 640.050 46.050 640.950 ;
        RECT 53.700 640.500 55.500 647.250 ;
        RECT 56.700 641.400 58.500 647.250 ;
        RECT 59.700 641.400 61.500 647.250 ;
        RECT 62.700 641.400 64.500 647.250 ;
        RECT 66.450 641.400 68.250 647.250 ;
        RECT 69.450 641.400 71.250 647.250 ;
        RECT 50.850 640.050 52.650 640.500 ;
        RECT 43.950 638.850 52.650 640.050 ;
        RECT 53.700 639.300 59.400 640.500 ;
        RECT 50.850 638.700 52.650 638.850 ;
        RECT 57.600 638.700 59.400 639.300 ;
        RECT 60.300 637.350 61.500 641.400 ;
        RECT 40.950 636.600 43.050 637.350 ;
        RECT 22.950 635.250 43.050 636.600 ;
        RECT 46.950 636.450 64.350 637.350 ;
        RECT 46.950 635.250 49.050 636.450 ;
        RECT 10.500 634.350 12.300 634.950 ;
        RECT 19.950 634.650 22.050 634.950 ;
        RECT 49.950 634.350 62.250 635.550 ;
        RECT 22.950 633.450 51.000 634.350 ;
        RECT 60.450 633.750 62.250 634.350 ;
        RECT 11.250 633.150 51.000 633.450 ;
        RECT 10.950 632.550 24.900 633.150 ;
        RECT 4.950 629.850 7.050 631.950 ;
        RECT 10.950 631.350 14.850 632.550 ;
        RECT 31.950 631.650 46.500 632.250 ;
        RECT 10.950 631.050 13.050 631.350 ;
        RECT 15.750 630.450 22.500 631.350 ;
        RECT 5.100 628.050 6.900 629.850 ;
        RECT 15.750 628.050 16.950 630.450 ;
        RECT 5.100 627.000 16.950 628.050 ;
        RECT 18.750 627.750 20.550 629.550 ;
        RECT 21.450 628.950 22.500 630.450 ;
        RECT 23.400 631.050 46.500 631.650 ;
        RECT 23.400 630.450 34.050 631.050 ;
        RECT 23.400 629.850 25.200 630.450 ;
        RECT 31.950 630.150 34.050 630.450 ;
        RECT 36.150 629.250 38.250 629.550 ;
        RECT 44.700 629.250 46.500 631.050 ;
        RECT 47.850 630.000 54.900 631.800 ;
        RECT 21.450 628.050 33.450 628.950 ;
        RECT 2.700 625.200 18.000 626.100 ;
        RECT 2.700 621.600 3.900 625.200 ;
        RECT 6.900 623.700 8.700 624.300 ;
        RECT 6.900 622.500 15.300 623.700 ;
        RECT 13.800 621.600 15.300 622.500 ;
        RECT 2.700 615.750 4.500 621.600 ;
        RECT 8.100 615.750 9.900 621.600 ;
        RECT 13.500 615.750 15.300 621.600 ;
        RECT 16.950 622.050 18.000 625.200 ;
        RECT 19.500 624.300 20.550 627.750 ;
        RECT 27.150 625.350 31.050 627.150 ;
        RECT 28.950 625.050 31.050 625.350 ;
        RECT 32.400 626.550 33.450 628.050 ;
        RECT 34.350 627.450 38.250 629.250 ;
        RECT 47.850 628.350 48.750 630.000 ;
        RECT 55.950 629.100 58.050 633.150 ;
        RECT 39.150 627.300 48.750 628.350 ;
        RECT 49.800 628.050 58.050 629.100 ;
        RECT 39.150 626.550 40.050 627.300 ;
        RECT 32.400 625.200 40.050 626.550 ;
        RECT 49.800 626.250 50.850 628.050 ;
        RECT 40.950 625.200 50.850 626.250 ;
        RECT 54.300 625.200 62.100 627.000 ;
        RECT 22.050 624.300 23.850 624.750 ;
        RECT 40.950 624.300 42.000 625.200 ;
        RECT 19.500 623.850 23.850 624.300 ;
        RECT 19.500 623.100 27.150 623.850 ;
        RECT 22.050 622.950 27.150 623.100 ;
        RECT 16.950 619.950 19.050 622.050 ;
        RECT 19.950 619.950 22.050 622.050 ;
        RECT 22.950 619.950 25.050 622.050 ;
        RECT 26.250 621.600 27.150 622.950 ;
        RECT 35.100 622.500 42.000 624.300 ;
        RECT 42.900 622.500 49.650 624.300 ;
        RECT 54.300 621.600 55.800 625.200 ;
        RECT 63.150 621.600 64.350 636.450 ;
        RECT 26.250 620.250 30.300 621.600 ;
        RECT 31.950 621.300 34.050 621.600 ;
        RECT 17.700 618.600 19.050 619.950 ;
        RECT 20.700 618.600 22.050 619.950 ;
        RECT 23.700 618.600 25.050 619.950 ;
        RECT 28.500 619.800 30.300 620.250 ;
        RECT 31.200 619.500 34.050 621.300 ;
        RECT 36.150 621.300 38.250 621.600 ;
        RECT 36.150 619.500 39.000 621.300 ;
        RECT 17.700 615.750 19.500 618.600 ;
        RECT 20.700 615.750 22.500 618.600 ;
        RECT 23.700 615.750 25.500 618.600 ;
        RECT 26.700 615.750 28.500 618.600 ;
        RECT 31.200 615.750 33.000 619.500 ;
        RECT 34.200 615.750 36.000 618.600 ;
        RECT 37.200 615.750 39.000 619.500 ;
        RECT 40.950 619.500 43.050 621.600 ;
        RECT 43.950 619.500 46.050 621.600 ;
        RECT 46.950 619.500 49.050 621.600 ;
        RECT 51.600 620.400 55.800 621.600 ;
        RECT 40.950 615.750 42.750 619.500 ;
        RECT 43.950 615.750 45.750 619.500 ;
        RECT 46.950 615.750 48.750 619.500 ;
        RECT 51.600 615.750 53.400 620.400 ;
        RECT 57.150 615.750 58.950 621.600 ;
        RECT 62.550 615.750 64.350 621.600 ;
        RECT 66.450 628.950 67.950 641.400 ;
        RECT 81.450 635.400 83.250 647.250 ;
        RECT 85.650 635.400 87.450 647.250 ;
        RECT 94.650 641.400 96.450 647.250 ;
        RECT 97.650 641.400 99.450 647.250 ;
        RECT 106.650 641.400 108.450 647.250 ;
        RECT 109.650 641.400 111.450 647.250 ;
        RECT 113.550 641.400 115.350 647.250 ;
        RECT 116.550 641.400 118.350 647.250 ;
        RECT 81.450 634.350 84.000 635.400 ;
        RECT 80.100 630.150 81.900 631.950 ;
        RECT 66.450 626.850 70.050 628.950 ;
        RECT 79.950 628.050 82.050 630.150 ;
        RECT 82.950 627.150 84.000 634.350 ;
        RECT 86.100 630.150 87.900 631.950 ;
        RECT 85.950 628.050 88.050 630.150 ;
        RECT 95.400 628.950 96.600 641.400 ;
        RECT 107.400 628.950 108.600 641.400 ;
        RECT 116.400 628.950 117.600 641.400 ;
        RECT 132.450 635.400 134.250 647.250 ;
        RECT 136.650 635.400 138.450 647.250 ;
        RECT 147.300 635.400 149.100 647.250 ;
        RECT 151.500 635.400 153.300 647.250 ;
        RECT 154.800 641.400 156.600 647.250 ;
        RECT 166.650 641.400 168.450 647.250 ;
        RECT 169.650 641.400 171.450 647.250 ;
        RECT 172.650 641.400 174.450 647.250 ;
        RECT 178.650 641.400 180.450 647.250 ;
        RECT 181.650 641.400 183.450 647.250 ;
        RECT 184.650 641.400 186.450 647.250 ;
        RECT 132.450 634.350 135.000 635.400 ;
        RECT 131.100 630.150 132.900 631.950 ;
        RECT 66.450 618.600 67.950 626.850 ;
        RECT 82.950 625.050 85.050 627.150 ;
        RECT 94.950 626.850 97.050 628.950 ;
        RECT 98.100 627.150 99.900 628.950 ;
        RECT 82.950 618.600 84.000 625.050 ;
        RECT 95.400 618.600 96.600 626.850 ;
        RECT 97.950 625.050 100.050 627.150 ;
        RECT 106.950 626.850 109.050 628.950 ;
        RECT 110.100 627.150 111.900 628.950 ;
        RECT 113.100 627.150 114.900 628.950 ;
        RECT 107.400 618.600 108.600 626.850 ;
        RECT 109.950 625.050 112.050 627.150 ;
        RECT 112.950 625.050 115.050 627.150 ;
        RECT 115.950 626.850 118.050 628.950 ;
        RECT 130.950 628.050 133.050 630.150 ;
        RECT 133.950 627.150 135.000 634.350 ;
        RECT 137.100 630.150 138.900 631.950 ;
        RECT 146.100 630.150 147.900 631.950 ;
        RECT 151.950 630.150 153.150 635.400 ;
        RECT 154.950 633.150 156.750 634.950 ;
        RECT 170.250 633.150 171.450 641.400 ;
        RECT 182.250 633.150 183.450 641.400 ;
        RECT 184.950 636.450 187.050 637.050 ;
        RECT 184.950 635.550 189.450 636.450 ;
        RECT 184.950 634.950 187.050 635.550 ;
        RECT 154.950 631.050 157.050 633.150 ;
        RECT 136.950 628.050 139.050 630.150 ;
        RECT 145.950 628.050 148.050 630.150 ;
        RECT 116.400 618.600 117.600 626.850 ;
        RECT 133.950 625.050 136.050 627.150 ;
        RECT 148.950 626.850 151.050 628.950 ;
        RECT 151.950 628.050 154.050 630.150 ;
        RECT 166.950 629.850 169.050 631.950 ;
        RECT 169.950 631.050 172.050 633.150 ;
        RECT 167.100 628.050 168.900 629.850 ;
        RECT 149.100 625.050 150.900 626.850 ;
        RECT 133.950 618.600 135.000 625.050 ;
        RECT 152.850 624.750 154.050 628.050 ;
        RECT 153.000 623.700 156.750 624.750 ;
        RECT 170.250 623.700 171.450 631.050 ;
        RECT 172.950 629.850 175.050 631.950 ;
        RECT 178.950 629.850 181.050 631.950 ;
        RECT 181.950 631.050 184.050 633.150 ;
        RECT 173.100 628.050 174.900 629.850 ;
        RECT 179.100 628.050 180.900 629.850 ;
        RECT 182.250 623.700 183.450 631.050 ;
        RECT 184.950 629.850 187.050 631.950 ;
        RECT 185.100 628.050 186.900 629.850 ;
        RECT 146.550 620.700 154.350 622.050 ;
        RECT 66.450 615.750 68.250 618.600 ;
        RECT 69.450 615.750 71.250 618.600 ;
        RECT 79.650 615.750 81.450 618.600 ;
        RECT 82.650 615.750 84.450 618.600 ;
        RECT 85.650 615.750 87.450 618.600 ;
        RECT 94.650 615.750 96.450 618.600 ;
        RECT 97.650 615.750 99.450 618.600 ;
        RECT 106.650 615.750 108.450 618.600 ;
        RECT 109.650 615.750 111.450 618.600 ;
        RECT 113.550 615.750 115.350 618.600 ;
        RECT 116.550 615.750 118.350 618.600 ;
        RECT 130.650 615.750 132.450 618.600 ;
        RECT 133.650 615.750 135.450 618.600 ;
        RECT 136.650 615.750 138.450 618.600 ;
        RECT 146.550 615.750 148.350 620.700 ;
        RECT 149.550 615.750 151.350 619.800 ;
        RECT 152.550 615.750 154.350 620.700 ;
        RECT 155.550 621.600 156.750 623.700 ;
        RECT 167.850 622.800 171.450 623.700 ;
        RECT 179.850 622.800 183.450 623.700 ;
        RECT 188.550 624.450 189.450 635.550 ;
        RECT 195.300 635.400 197.100 647.250 ;
        RECT 199.500 635.400 201.300 647.250 ;
        RECT 202.800 641.400 204.600 647.250 ;
        RECT 217.650 641.400 219.450 647.250 ;
        RECT 220.650 642.000 222.450 647.250 ;
        RECT 218.250 641.100 219.450 641.400 ;
        RECT 223.650 641.400 225.450 647.250 ;
        RECT 226.650 641.400 228.450 647.250 ;
        RECT 232.650 641.400 234.450 647.250 ;
        RECT 235.650 641.400 237.450 647.250 ;
        RECT 239.550 641.400 241.350 647.250 ;
        RECT 242.550 641.400 244.350 647.250 ;
        RECT 245.550 642.000 247.350 647.250 ;
        RECT 223.650 641.100 225.300 641.400 ;
        RECT 218.250 640.200 225.300 641.100 ;
        RECT 194.100 630.150 195.900 631.950 ;
        RECT 199.950 630.150 201.150 635.400 ;
        RECT 202.950 633.150 204.750 634.950 ;
        RECT 202.950 631.050 205.050 633.150 ;
        RECT 218.250 631.950 219.300 640.200 ;
        RECT 224.100 636.150 225.900 637.950 ;
        RECT 220.950 633.150 222.750 634.950 ;
        RECT 223.950 634.050 226.050 636.150 ;
        RECT 227.100 633.150 228.900 634.950 ;
        RECT 193.950 628.050 196.050 630.150 ;
        RECT 196.950 626.850 199.050 628.950 ;
        RECT 199.950 628.050 202.050 630.150 ;
        RECT 217.950 629.850 220.050 631.950 ;
        RECT 220.950 631.050 223.050 633.150 ;
        RECT 226.950 631.050 229.050 633.150 ;
        RECT 197.100 625.050 198.900 626.850 ;
        RECT 193.950 624.450 196.050 625.050 ;
        RECT 200.850 624.750 202.050 628.050 ;
        RECT 218.400 625.650 219.600 629.850 ;
        RECT 233.400 628.950 234.600 641.400 ;
        RECT 242.700 641.100 244.350 641.400 ;
        RECT 248.550 641.400 250.350 647.250 ;
        RECT 262.650 641.400 264.450 647.250 ;
        RECT 265.650 641.400 267.450 647.250 ;
        RECT 268.650 641.400 270.450 647.250 ;
        RECT 281.400 641.400 283.200 647.250 ;
        RECT 248.550 641.100 249.750 641.400 ;
        RECT 242.700 640.200 249.750 641.100 ;
        RECT 242.100 636.150 243.900 637.950 ;
        RECT 239.100 633.150 240.900 634.950 ;
        RECT 241.950 634.050 244.050 636.150 ;
        RECT 245.250 633.150 247.050 634.950 ;
        RECT 238.950 631.050 241.050 633.150 ;
        RECT 244.950 631.050 247.050 633.150 ;
        RECT 248.700 631.950 249.750 640.200 ;
        RECT 266.250 633.150 267.450 641.400 ;
        RECT 284.700 635.400 286.500 647.250 ;
        RECT 288.900 635.400 290.700 647.250 ;
        RECT 298.650 641.400 300.450 647.250 ;
        RECT 301.650 641.400 303.450 647.250 ;
        RECT 307.650 641.400 309.450 647.250 ;
        RECT 310.650 641.400 312.450 647.250 ;
        RECT 313.650 641.400 315.450 647.250 ;
        RECT 317.550 641.400 319.350 647.250 ;
        RECT 320.550 641.400 322.350 647.250 ;
        RECT 323.550 641.400 325.350 647.250 ;
        RECT 281.250 633.150 283.050 634.950 ;
        RECT 247.950 629.850 250.050 631.950 ;
        RECT 262.950 629.850 265.050 631.950 ;
        RECT 265.950 631.050 268.050 633.150 ;
        RECT 232.950 626.850 235.050 628.950 ;
        RECT 236.100 627.150 237.900 628.950 ;
        RECT 188.550 623.550 196.050 624.450 ;
        RECT 201.000 623.700 204.750 624.750 ;
        RECT 218.400 624.000 222.900 625.650 ;
        RECT 193.950 622.950 196.050 623.550 ;
        RECT 155.550 615.750 157.350 621.600 ;
        RECT 167.850 615.750 169.650 622.800 ;
        RECT 172.350 615.750 174.150 621.600 ;
        RECT 179.850 615.750 181.650 622.800 ;
        RECT 184.350 615.750 186.150 621.600 ;
        RECT 194.550 620.700 202.350 622.050 ;
        RECT 194.550 615.750 196.350 620.700 ;
        RECT 197.550 615.750 199.350 619.800 ;
        RECT 200.550 615.750 202.350 620.700 ;
        RECT 203.550 621.600 204.750 623.700 ;
        RECT 203.550 615.750 205.350 621.600 ;
        RECT 221.100 615.750 222.900 624.000 ;
        RECT 226.500 615.750 228.300 624.600 ;
        RECT 233.400 618.600 234.600 626.850 ;
        RECT 235.950 625.050 238.050 627.150 ;
        RECT 248.400 625.650 249.600 629.850 ;
        RECT 263.100 628.050 264.900 629.850 ;
        RECT 232.650 615.750 234.450 618.600 ;
        RECT 235.650 615.750 237.450 618.600 ;
        RECT 239.700 615.750 241.500 624.600 ;
        RECT 245.100 624.000 249.600 625.650 ;
        RECT 245.100 615.750 246.900 624.000 ;
        RECT 266.250 623.700 267.450 631.050 ;
        RECT 268.950 629.850 271.050 631.950 ;
        RECT 280.950 631.050 283.050 633.150 ;
        RECT 284.850 630.150 286.050 635.400 ;
        RECT 290.100 630.150 291.900 631.950 ;
        RECT 269.100 628.050 270.900 629.850 ;
        RECT 283.950 628.050 286.050 630.150 ;
        RECT 283.950 624.750 285.150 628.050 ;
        RECT 286.950 626.850 289.050 628.950 ;
        RECT 289.950 628.050 292.050 630.150 ;
        RECT 299.400 628.950 300.600 641.400 ;
        RECT 311.250 633.150 312.450 641.400 ;
        RECT 320.550 633.150 321.750 641.400 ;
        RECT 336.300 635.400 338.100 647.250 ;
        RECT 340.500 635.400 342.300 647.250 ;
        RECT 343.800 641.400 345.600 647.250 ;
        RECT 350.550 641.400 352.350 647.250 ;
        RECT 353.550 641.400 355.350 647.250 ;
        RECT 356.550 641.400 358.350 647.250 ;
        RECT 370.650 641.400 372.450 647.250 ;
        RECT 373.650 641.400 375.450 647.250 ;
        RECT 376.650 641.400 378.450 647.250 ;
        RECT 307.950 629.850 310.050 631.950 ;
        RECT 310.950 631.050 313.050 633.150 ;
        RECT 298.950 626.850 301.050 628.950 ;
        RECT 302.100 627.150 303.900 628.950 ;
        RECT 308.100 628.050 309.900 629.850 ;
        RECT 287.100 625.050 288.900 626.850 ;
        RECT 263.850 622.800 267.450 623.700 ;
        RECT 281.250 623.700 285.000 624.750 ;
        RECT 263.850 615.750 265.650 622.800 ;
        RECT 281.250 621.600 282.450 623.700 ;
        RECT 268.350 615.750 270.150 621.600 ;
        RECT 280.650 615.750 282.450 621.600 ;
        RECT 283.650 620.700 291.450 622.050 ;
        RECT 283.650 615.750 285.450 620.700 ;
        RECT 286.650 615.750 288.450 619.800 ;
        RECT 289.650 615.750 291.450 620.700 ;
        RECT 299.400 618.600 300.600 626.850 ;
        RECT 301.950 625.050 304.050 627.150 ;
        RECT 311.250 623.700 312.450 631.050 ;
        RECT 313.950 629.850 316.050 631.950 ;
        RECT 316.950 629.850 319.050 631.950 ;
        RECT 319.950 631.050 322.050 633.150 ;
        RECT 314.100 628.050 315.900 629.850 ;
        RECT 317.100 628.050 318.900 629.850 ;
        RECT 308.850 622.800 312.450 623.700 ;
        RECT 320.550 623.700 321.750 631.050 ;
        RECT 322.950 629.850 325.050 631.950 ;
        RECT 335.100 630.150 336.900 631.950 ;
        RECT 340.950 630.150 342.150 635.400 ;
        RECT 343.950 633.150 345.750 634.950 ;
        RECT 353.550 633.150 354.750 641.400 ;
        RECT 374.250 633.150 375.450 641.400 ;
        RECT 383.550 635.400 385.350 647.250 ;
        RECT 387.750 635.400 389.550 647.250 ;
        RECT 400.650 641.400 402.450 647.250 ;
        RECT 403.650 641.400 405.450 647.250 ;
        RECT 406.650 641.400 408.450 647.250 ;
        RECT 415.650 641.400 417.450 647.250 ;
        RECT 418.650 641.400 420.450 647.250 ;
        RECT 427.650 641.400 429.450 647.250 ;
        RECT 430.650 641.400 432.450 647.250 ;
        RECT 433.650 641.400 435.450 647.250 ;
        RECT 400.950 636.450 403.050 637.050 ;
        RECT 387.000 634.350 389.550 635.400 ;
        RECT 398.550 635.550 403.050 636.450 ;
        RECT 343.950 631.050 346.050 633.150 ;
        RECT 323.100 628.050 324.900 629.850 ;
        RECT 334.950 628.050 337.050 630.150 ;
        RECT 337.950 626.850 340.050 628.950 ;
        RECT 340.950 628.050 343.050 630.150 ;
        RECT 349.950 629.850 352.050 631.950 ;
        RECT 352.950 631.050 355.050 633.150 ;
        RECT 350.100 628.050 351.900 629.850 ;
        RECT 338.100 625.050 339.900 626.850 ;
        RECT 341.850 624.750 343.050 628.050 ;
        RECT 342.000 623.700 345.750 624.750 ;
        RECT 320.550 622.800 324.150 623.700 ;
        RECT 298.650 615.750 300.450 618.600 ;
        RECT 301.650 615.750 303.450 618.600 ;
        RECT 308.850 615.750 310.650 622.800 ;
        RECT 313.350 615.750 315.150 621.600 ;
        RECT 317.850 615.750 319.650 621.600 ;
        RECT 322.350 615.750 324.150 622.800 ;
        RECT 335.550 620.700 343.350 622.050 ;
        RECT 335.550 615.750 337.350 620.700 ;
        RECT 338.550 615.750 340.350 619.800 ;
        RECT 341.550 615.750 343.350 620.700 ;
        RECT 344.550 621.600 345.750 623.700 ;
        RECT 353.550 623.700 354.750 631.050 ;
        RECT 355.950 629.850 358.050 631.950 ;
        RECT 370.950 629.850 373.050 631.950 ;
        RECT 373.950 631.050 376.050 633.150 ;
        RECT 356.100 628.050 357.900 629.850 ;
        RECT 371.100 628.050 372.900 629.850 ;
        RECT 374.250 623.700 375.450 631.050 ;
        RECT 376.950 629.850 379.050 631.950 ;
        RECT 383.100 630.150 384.900 631.950 ;
        RECT 377.100 628.050 378.900 629.850 ;
        RECT 382.950 628.050 385.050 630.150 ;
        RECT 387.000 627.150 388.050 634.350 ;
        RECT 389.100 630.150 390.900 631.950 ;
        RECT 388.950 628.050 391.050 630.150 ;
        RECT 385.950 625.050 388.050 627.150 ;
        RECT 353.550 622.800 357.150 623.700 ;
        RECT 344.550 615.750 346.350 621.600 ;
        RECT 350.850 615.750 352.650 621.600 ;
        RECT 355.350 615.750 357.150 622.800 ;
        RECT 371.850 622.800 375.450 623.700 ;
        RECT 371.850 615.750 373.650 622.800 ;
        RECT 376.350 615.750 378.150 621.600 ;
        RECT 387.000 618.600 388.050 625.050 ;
        RECT 388.950 624.450 391.050 625.050 ;
        RECT 398.550 624.450 399.450 635.550 ;
        RECT 400.950 634.950 403.050 635.550 ;
        RECT 404.250 633.150 405.450 641.400 ;
        RECT 406.950 636.450 409.050 637.050 ;
        RECT 412.950 636.450 415.050 637.050 ;
        RECT 406.950 635.550 415.050 636.450 ;
        RECT 406.950 634.950 409.050 635.550 ;
        RECT 412.950 634.950 415.050 635.550 ;
        RECT 400.950 629.850 403.050 631.950 ;
        RECT 403.950 631.050 406.050 633.150 ;
        RECT 401.100 628.050 402.900 629.850 ;
        RECT 388.950 623.550 399.450 624.450 ;
        RECT 404.250 623.700 405.450 631.050 ;
        RECT 406.950 629.850 409.050 631.950 ;
        RECT 407.100 628.050 408.900 629.850 ;
        RECT 416.400 628.950 417.600 641.400 ;
        RECT 431.250 633.150 432.450 641.400 ;
        RECT 442.650 635.400 444.450 647.250 ;
        RECT 445.650 636.300 447.450 647.250 ;
        RECT 448.650 637.200 450.450 647.250 ;
        RECT 451.650 636.300 453.450 647.250 ;
        RECT 458.550 637.500 460.350 647.250 ;
        RECT 461.550 638.400 463.350 647.250 ;
        RECT 464.550 646.500 472.350 647.250 ;
        RECT 464.550 637.500 466.350 646.500 ;
        RECT 458.550 636.600 466.350 637.500 ;
        RECT 467.550 637.800 469.350 645.600 ;
        RECT 470.550 638.700 472.350 646.500 ;
        RECT 474.150 646.500 481.950 647.250 ;
        RECT 474.150 637.800 475.950 646.500 ;
        RECT 467.550 636.900 475.950 637.800 ;
        RECT 477.150 637.800 478.950 645.600 ;
        RECT 445.650 635.400 453.450 636.300 ;
        RECT 477.150 635.400 478.350 637.800 ;
        RECT 480.150 637.200 481.950 646.500 ;
        RECT 493.650 641.400 495.450 647.250 ;
        RECT 496.650 641.400 498.450 647.250 ;
        RECT 499.650 641.400 501.450 647.250 ;
        RECT 506.550 641.400 508.350 647.250 ;
        RECT 509.550 641.400 511.350 647.250 ;
        RECT 512.550 641.400 514.350 647.250 ;
        RECT 427.950 629.850 430.050 631.950 ;
        RECT 430.950 631.050 433.050 633.150 ;
        RECT 415.950 626.850 418.050 628.950 ;
        RECT 419.100 627.150 420.900 628.950 ;
        RECT 428.100 628.050 429.900 629.850 ;
        RECT 388.950 622.950 391.050 623.550 ;
        RECT 401.850 622.800 405.450 623.700 ;
        RECT 383.550 615.750 385.350 618.600 ;
        RECT 386.550 615.750 388.350 618.600 ;
        RECT 389.550 615.750 391.350 618.600 ;
        RECT 401.850 615.750 403.650 622.800 ;
        RECT 406.350 615.750 408.150 621.600 ;
        RECT 416.400 618.600 417.600 626.850 ;
        RECT 418.950 625.050 421.050 627.150 ;
        RECT 431.250 623.700 432.450 631.050 ;
        RECT 433.950 629.850 436.050 631.950 ;
        RECT 443.100 630.150 444.300 635.400 ;
        RECT 474.900 634.200 478.350 635.400 ;
        RECT 484.950 636.450 487.050 637.050 ;
        RECT 493.950 636.450 496.050 637.050 ;
        RECT 484.950 635.550 496.050 636.450 ;
        RECT 484.950 634.950 487.050 635.550 ;
        RECT 493.950 634.950 496.050 635.550 ;
        RECT 461.100 630.150 462.900 631.950 ;
        RECT 470.100 630.150 471.900 631.950 ;
        RECT 434.100 628.050 435.900 629.850 ;
        RECT 442.950 628.050 445.050 630.150 ;
        RECT 428.850 622.800 432.450 623.700 ;
        RECT 415.650 615.750 417.450 618.600 ;
        RECT 418.650 615.750 420.450 618.600 ;
        RECT 428.850 615.750 430.650 622.800 ;
        RECT 443.100 621.600 444.300 628.050 ;
        RECT 445.950 626.850 448.050 628.950 ;
        RECT 449.100 627.150 450.900 628.950 ;
        RECT 446.100 625.050 447.900 626.850 ;
        RECT 448.950 625.050 451.050 627.150 ;
        RECT 451.950 626.850 454.050 628.950 ;
        RECT 460.950 628.050 463.050 630.150 ;
        RECT 466.950 626.850 469.050 628.950 ;
        RECT 469.950 628.050 472.050 630.150 ;
        RECT 474.900 628.950 476.100 634.200 ;
        RECT 497.250 633.150 498.450 641.400 ;
        RECT 499.950 636.450 502.050 637.050 ;
        RECT 499.950 635.550 504.450 636.450 ;
        RECT 499.950 634.950 502.050 635.550 ;
        RECT 493.950 629.850 496.050 631.950 ;
        RECT 496.950 631.050 499.050 633.150 ;
        RECT 474.900 626.850 478.050 628.950 ;
        RECT 494.100 628.050 495.900 629.850 ;
        RECT 452.100 625.050 453.900 626.850 ;
        RECT 467.100 625.050 468.900 626.850 ;
        RECT 433.350 615.750 435.150 621.600 ;
        RECT 443.100 619.950 448.800 621.600 ;
        RECT 443.700 615.750 445.500 618.600 ;
        RECT 447.000 615.750 448.800 619.950 ;
        RECT 451.200 615.750 453.000 621.600 ;
        RECT 474.900 620.400 476.100 626.850 ;
        RECT 497.250 623.700 498.450 631.050 ;
        RECT 499.950 629.850 502.050 631.950 ;
        RECT 500.100 628.050 501.900 629.850 ;
        RECT 465.300 619.500 476.100 620.400 ;
        RECT 494.850 622.800 498.450 623.700 ;
        RECT 503.550 624.450 504.450 635.550 ;
        RECT 509.550 633.150 510.750 641.400 ;
        RECT 521.550 635.400 523.350 647.250 ;
        RECT 525.750 635.400 527.550 647.250 ;
        RECT 535.650 641.400 537.450 647.250 ;
        RECT 538.650 641.400 540.450 647.250 ;
        RECT 545.400 641.400 547.200 647.250 ;
        RECT 525.000 634.350 527.550 635.400 ;
        RECT 505.950 629.850 508.050 631.950 ;
        RECT 508.950 631.050 511.050 633.150 ;
        RECT 506.100 628.050 507.900 629.850 ;
        RECT 505.950 624.450 508.050 625.050 ;
        RECT 503.550 623.550 508.050 624.450 ;
        RECT 505.950 622.950 508.050 623.550 ;
        RECT 509.550 623.700 510.750 631.050 ;
        RECT 511.950 629.850 514.050 631.950 ;
        RECT 521.100 630.150 522.900 631.950 ;
        RECT 512.100 628.050 513.900 629.850 ;
        RECT 520.950 628.050 523.050 630.150 ;
        RECT 525.000 627.150 526.050 634.350 ;
        RECT 527.100 630.150 528.900 631.950 ;
        RECT 526.950 628.050 529.050 630.150 ;
        RECT 536.400 628.950 537.600 641.400 ;
        RECT 548.700 635.400 550.500 647.250 ;
        RECT 552.900 635.400 554.700 647.250 ;
        RECT 560.550 635.400 562.350 647.250 ;
        RECT 564.750 635.400 566.550 647.250 ;
        RECT 574.650 641.400 576.450 647.250 ;
        RECT 577.650 641.400 579.450 647.250 ;
        RECT 580.650 641.400 582.450 647.250 ;
        RECT 545.250 633.150 547.050 634.950 ;
        RECT 544.950 631.050 547.050 633.150 ;
        RECT 548.850 630.150 550.050 635.400 ;
        RECT 564.000 634.350 566.550 635.400 ;
        RECT 554.100 630.150 555.900 631.950 ;
        RECT 560.100 630.150 561.900 631.950 ;
        RECT 523.950 625.050 526.050 627.150 ;
        RECT 535.950 626.850 538.050 628.950 ;
        RECT 539.100 627.150 540.900 628.950 ;
        RECT 547.950 628.050 550.050 630.150 ;
        RECT 509.550 622.800 513.150 623.700 ;
        RECT 465.300 618.600 466.350 619.500 ;
        RECT 471.300 618.600 472.350 619.500 ;
        RECT 461.250 615.750 463.350 618.600 ;
        RECT 464.550 615.750 466.350 618.600 ;
        RECT 467.550 615.750 469.350 618.600 ;
        RECT 470.550 615.750 472.350 618.600 ;
        RECT 494.850 615.750 496.650 622.800 ;
        RECT 499.350 615.750 501.150 621.600 ;
        RECT 506.850 615.750 508.650 621.600 ;
        RECT 511.350 615.750 513.150 622.800 ;
        RECT 525.000 618.600 526.050 625.050 ;
        RECT 536.400 618.600 537.600 626.850 ;
        RECT 538.950 625.050 541.050 627.150 ;
        RECT 547.950 624.750 549.150 628.050 ;
        RECT 550.950 626.850 553.050 628.950 ;
        RECT 553.950 628.050 556.050 630.150 ;
        RECT 559.950 628.050 562.050 630.150 ;
        RECT 564.000 627.150 565.050 634.350 ;
        RECT 578.250 633.150 579.450 641.400 ;
        RECT 590.550 635.400 592.350 647.250 ;
        RECT 595.050 635.550 596.850 647.250 ;
        RECT 598.050 636.900 599.850 647.250 ;
        RECT 608.550 641.400 610.350 647.250 ;
        RECT 611.550 641.400 613.350 647.250 ;
        RECT 614.550 642.000 616.350 647.250 ;
        RECT 611.700 641.100 613.350 641.400 ;
        RECT 617.550 641.400 619.350 647.250 ;
        RECT 628.650 641.400 630.450 647.250 ;
        RECT 631.650 642.000 633.450 647.250 ;
        RECT 617.550 641.100 618.750 641.400 ;
        RECT 611.700 640.200 618.750 641.100 ;
        RECT 598.050 635.550 600.450 636.900 ;
        RECT 611.100 636.150 612.900 637.950 ;
        RECT 590.550 634.200 591.750 635.400 ;
        RECT 595.950 634.200 597.750 634.650 ;
        RECT 566.100 630.150 567.900 631.950 ;
        RECT 565.950 628.050 568.050 630.150 ;
        RECT 574.950 629.850 577.050 631.950 ;
        RECT 577.950 631.050 580.050 633.150 ;
        RECT 590.550 633.000 597.750 634.200 ;
        RECT 595.950 632.850 597.750 633.000 ;
        RECT 575.100 628.050 576.900 629.850 ;
        RECT 551.100 625.050 552.900 626.850 ;
        RECT 562.950 625.050 565.050 627.150 ;
        RECT 545.250 623.700 549.000 624.750 ;
        RECT 545.250 621.600 546.450 623.700 ;
        RECT 521.550 615.750 523.350 618.600 ;
        RECT 524.550 615.750 526.350 618.600 ;
        RECT 527.550 615.750 529.350 618.600 ;
        RECT 535.650 615.750 537.450 618.600 ;
        RECT 538.650 615.750 540.450 618.600 ;
        RECT 544.650 615.750 546.450 621.600 ;
        RECT 547.650 620.700 555.450 622.050 ;
        RECT 547.650 615.750 549.450 620.700 ;
        RECT 550.650 615.750 552.450 619.800 ;
        RECT 553.650 615.750 555.450 620.700 ;
        RECT 564.000 618.600 565.050 625.050 ;
        RECT 578.250 623.700 579.450 631.050 ;
        RECT 580.950 629.850 583.050 631.950 ;
        RECT 593.100 630.150 594.900 631.950 ;
        RECT 581.100 628.050 582.900 629.850 ;
        RECT 590.100 627.150 591.900 628.950 ;
        RECT 592.950 628.050 595.050 630.150 ;
        RECT 589.950 625.050 592.050 627.150 ;
        RECT 596.700 624.600 597.600 632.850 ;
        RECT 599.100 628.950 600.450 635.550 ;
        RECT 608.100 633.150 609.900 634.950 ;
        RECT 610.950 634.050 613.050 636.150 ;
        RECT 614.250 633.150 616.050 634.950 ;
        RECT 607.950 631.050 610.050 633.150 ;
        RECT 613.950 631.050 616.050 633.150 ;
        RECT 617.700 631.950 618.750 640.200 ;
        RECT 629.250 641.100 630.450 641.400 ;
        RECT 634.650 641.400 636.450 647.250 ;
        RECT 637.650 641.400 639.450 647.250 ;
        RECT 634.650 641.100 636.300 641.400 ;
        RECT 629.250 640.200 636.300 641.100 ;
        RECT 629.250 631.950 630.300 640.200 ;
        RECT 635.100 636.150 636.900 637.950 ;
        RECT 647.550 636.300 649.350 647.250 ;
        RECT 650.550 637.200 652.350 647.250 ;
        RECT 653.550 636.300 655.350 647.250 ;
        RECT 631.950 633.150 633.750 634.950 ;
        RECT 634.950 634.050 637.050 636.150 ;
        RECT 647.550 635.400 655.350 636.300 ;
        RECT 656.550 635.400 658.350 647.250 ;
        RECT 666.300 635.400 668.100 647.250 ;
        RECT 670.500 635.400 672.300 647.250 ;
        RECT 673.800 641.400 675.600 647.250 ;
        RECT 686.400 641.400 688.200 647.250 ;
        RECT 689.700 635.400 691.500 647.250 ;
        RECT 693.900 635.400 695.700 647.250 ;
        RECT 699.750 641.400 701.550 647.250 ;
        RECT 702.750 641.400 704.550 647.250 ;
        RECT 706.500 641.400 708.300 647.250 ;
        RECT 709.500 641.400 711.300 647.250 ;
        RECT 712.500 641.400 714.300 647.250 ;
        RECT 638.100 633.150 639.900 634.950 ;
        RECT 616.950 629.850 619.050 631.950 ;
        RECT 628.950 629.850 631.050 631.950 ;
        RECT 631.950 631.050 634.050 633.150 ;
        RECT 637.950 631.050 640.050 633.150 ;
        RECT 656.700 630.150 657.900 635.400 ;
        RECT 665.100 630.150 666.900 631.950 ;
        RECT 670.950 630.150 672.150 635.400 ;
        RECT 673.950 633.150 675.750 634.950 ;
        RECT 686.250 633.150 688.050 634.950 ;
        RECT 673.950 631.050 676.050 633.150 ;
        RECT 685.950 631.050 688.050 633.150 ;
        RECT 689.850 630.150 691.050 635.400 ;
        RECT 695.100 630.150 696.900 631.950 ;
        RECT 598.950 626.850 601.050 628.950 ;
        RECT 595.950 623.700 597.750 624.600 ;
        RECT 575.850 622.800 579.450 623.700 ;
        RECT 594.450 622.800 597.750 623.700 ;
        RECT 560.550 615.750 562.350 618.600 ;
        RECT 563.550 615.750 565.350 618.600 ;
        RECT 566.550 615.750 568.350 618.600 ;
        RECT 575.850 615.750 577.650 622.800 ;
        RECT 580.350 615.750 582.150 621.600 ;
        RECT 594.450 618.600 595.350 622.800 ;
        RECT 600.000 621.600 601.050 626.850 ;
        RECT 617.400 625.650 618.600 629.850 ;
        RECT 590.550 615.750 592.350 618.600 ;
        RECT 593.550 615.750 595.350 618.600 ;
        RECT 596.550 615.750 598.350 618.600 ;
        RECT 599.550 615.750 601.350 621.600 ;
        RECT 608.700 615.750 610.500 624.600 ;
        RECT 614.100 624.000 618.600 625.650 ;
        RECT 629.400 625.650 630.600 629.850 ;
        RECT 646.950 626.850 649.050 628.950 ;
        RECT 650.100 627.150 651.900 628.950 ;
        RECT 629.400 624.000 633.900 625.650 ;
        RECT 647.100 625.050 648.900 626.850 ;
        RECT 649.950 625.050 652.050 627.150 ;
        RECT 652.950 626.850 655.050 628.950 ;
        RECT 655.950 628.050 658.050 630.150 ;
        RECT 664.950 628.050 667.050 630.150 ;
        RECT 653.100 625.050 654.900 626.850 ;
        RECT 614.100 615.750 615.900 624.000 ;
        RECT 632.100 615.750 633.900 624.000 ;
        RECT 637.500 615.750 639.300 624.600 ;
        RECT 656.700 621.600 657.900 628.050 ;
        RECT 667.950 626.850 670.050 628.950 ;
        RECT 670.950 628.050 673.050 630.150 ;
        RECT 668.100 625.050 669.900 626.850 ;
        RECT 671.850 624.750 673.050 628.050 ;
        RECT 688.950 628.050 691.050 630.150 ;
        RECT 688.950 624.750 690.150 628.050 ;
        RECT 691.950 626.850 694.050 628.950 ;
        RECT 694.950 628.050 697.050 630.150 ;
        RECT 703.050 628.950 704.550 641.400 ;
        RECT 709.500 637.350 710.700 641.400 ;
        RECT 715.500 640.500 717.300 647.250 ;
        RECT 718.500 641.400 720.300 647.250 ;
        RECT 722.250 644.400 724.050 647.250 ;
        RECT 722.400 643.200 723.900 644.400 ;
        RECT 721.800 641.100 723.900 643.200 ;
        RECT 725.250 640.950 727.050 647.250 ;
        RECT 728.250 644.400 730.050 647.250 ;
        RECT 711.600 639.300 717.300 640.500 ;
        RECT 718.350 640.050 720.150 640.500 ;
        RECT 724.950 640.050 727.050 640.950 ;
        RECT 711.600 638.700 713.400 639.300 ;
        RECT 718.350 638.850 727.050 640.050 ;
        RECT 718.350 638.700 720.150 638.850 ;
        RECT 728.550 637.350 729.900 644.400 ;
        RECT 732.000 640.500 733.800 647.250 ;
        RECT 735.000 641.400 736.800 647.250 ;
        RECT 738.000 641.400 739.800 647.250 ;
        RECT 741.750 641.400 743.550 647.250 ;
        RECT 744.750 644.400 746.700 647.250 ;
        RECT 747.750 644.400 749.850 647.250 ;
        RECT 750.750 644.400 753.150 647.250 ;
        RECT 745.500 643.050 746.700 644.400 ;
        RECT 748.950 643.050 749.850 644.400 ;
        RECT 751.950 643.050 753.150 644.400 ;
        RECT 754.500 643.950 756.300 647.250 ;
        RECT 745.500 641.400 748.050 643.050 ;
        RECT 738.000 640.500 739.350 641.400 ;
        RECT 745.950 640.950 748.050 641.400 ;
        RECT 748.950 640.950 751.050 643.050 ;
        RECT 751.950 640.950 754.050 643.050 ;
        RECT 732.000 640.200 735.000 640.500 ;
        RECT 731.100 638.400 735.000 640.200 ;
        RECT 736.950 638.850 739.350 640.500 ;
        RECT 736.950 638.400 739.050 638.850 ;
        RECT 757.500 638.700 759.300 647.250 ;
        RECT 760.500 641.400 762.300 647.250 ;
        RECT 763.500 641.400 765.300 647.250 ;
        RECT 766.500 641.400 768.300 647.250 ;
        RECT 771.750 641.400 773.550 647.250 ;
        RECT 774.750 641.400 776.550 647.250 ;
        RECT 778.500 641.400 780.300 647.250 ;
        RECT 781.500 641.400 783.300 647.250 ;
        RECT 784.500 641.400 786.300 647.250 ;
        RECT 764.250 640.500 765.300 641.400 ;
        RECT 764.250 639.600 768.300 640.500 ;
        RECT 746.100 637.650 763.800 638.700 ;
        RECT 700.950 626.850 704.550 628.950 ;
        RECT 692.100 625.050 693.900 626.850 ;
        RECT 672.000 623.700 675.750 624.750 ;
        RECT 648.000 615.750 649.800 621.600 ;
        RECT 652.200 619.950 657.900 621.600 ;
        RECT 665.550 620.700 673.350 622.050 ;
        RECT 652.200 615.750 654.000 619.950 ;
        RECT 655.500 615.750 657.300 618.600 ;
        RECT 665.550 615.750 667.350 620.700 ;
        RECT 668.550 615.750 670.350 619.800 ;
        RECT 671.550 615.750 673.350 620.700 ;
        RECT 674.550 621.600 675.750 623.700 ;
        RECT 686.250 623.700 690.000 624.750 ;
        RECT 686.250 621.600 687.450 623.700 ;
        RECT 674.550 615.750 676.350 621.600 ;
        RECT 685.650 615.750 687.450 621.600 ;
        RECT 688.650 620.700 696.450 622.050 ;
        RECT 688.650 615.750 690.450 620.700 ;
        RECT 691.650 615.750 693.450 619.800 ;
        RECT 694.650 615.750 696.450 620.700 ;
        RECT 703.050 618.600 704.550 626.850 ;
        RECT 699.750 615.750 701.550 618.600 ;
        RECT 702.750 615.750 704.550 618.600 ;
        RECT 706.650 636.450 724.050 637.350 ;
        RECT 706.650 621.600 707.850 636.450 ;
        RECT 708.750 634.350 721.050 635.550 ;
        RECT 721.950 635.250 724.050 636.450 ;
        RECT 727.950 636.600 730.050 637.350 ;
        RECT 746.100 636.600 748.050 637.650 ;
        RECT 762.000 636.900 763.800 637.650 ;
        RECT 727.950 635.250 748.050 636.600 ;
        RECT 748.950 636.150 751.050 636.750 ;
        RECT 748.950 634.950 760.500 636.150 ;
        RECT 748.950 634.650 751.050 634.950 ;
        RECT 758.700 634.350 760.500 634.950 ;
        RECT 708.750 633.750 710.550 634.350 ;
        RECT 720.000 633.450 748.050 634.350 ;
        RECT 720.000 633.150 759.750 633.450 ;
        RECT 712.950 629.100 715.050 633.150 ;
        RECT 746.100 632.550 760.050 633.150 ;
        RECT 716.100 630.000 723.150 631.800 ;
        RECT 712.950 628.050 721.200 629.100 ;
        RECT 708.900 625.200 716.700 627.000 ;
        RECT 720.150 626.250 721.200 628.050 ;
        RECT 722.250 628.350 723.150 630.000 ;
        RECT 724.500 631.650 739.050 632.250 ;
        RECT 724.500 631.050 747.600 631.650 ;
        RECT 756.150 631.350 760.050 632.550 ;
        RECT 724.500 629.250 726.300 631.050 ;
        RECT 736.950 630.450 747.600 631.050 ;
        RECT 736.950 630.150 739.050 630.450 ;
        RECT 745.800 629.850 747.600 630.450 ;
        RECT 748.500 630.450 755.250 631.350 ;
        RECT 757.950 631.050 760.050 631.350 ;
        RECT 732.750 629.250 734.850 629.550 ;
        RECT 722.250 627.300 731.850 628.350 ;
        RECT 732.750 627.450 736.650 629.250 ;
        RECT 748.500 628.950 749.550 630.450 ;
        RECT 737.550 628.050 749.550 628.950 ;
        RECT 730.950 626.550 731.850 627.300 ;
        RECT 737.550 626.550 738.600 628.050 ;
        RECT 750.450 627.750 752.250 629.550 ;
        RECT 754.050 628.050 755.250 630.450 ;
        RECT 763.950 629.850 766.050 631.950 ;
        RECT 764.100 628.050 765.900 629.850 ;
        RECT 720.150 625.200 730.050 626.250 ;
        RECT 730.950 625.200 738.600 626.550 ;
        RECT 739.950 625.350 743.850 627.150 ;
        RECT 715.200 621.600 716.700 625.200 ;
        RECT 729.000 624.300 730.050 625.200 ;
        RECT 739.950 625.050 742.050 625.350 ;
        RECT 747.150 624.300 748.950 624.750 ;
        RECT 750.450 624.300 751.500 627.750 ;
        RECT 754.050 627.000 765.900 628.050 ;
        RECT 767.100 626.100 768.300 639.600 ;
        RECT 775.050 628.950 776.550 641.400 ;
        RECT 781.500 637.350 782.700 641.400 ;
        RECT 787.500 640.500 789.300 647.250 ;
        RECT 790.500 641.400 792.300 647.250 ;
        RECT 794.250 644.400 796.050 647.250 ;
        RECT 794.400 643.200 795.900 644.400 ;
        RECT 793.800 641.100 795.900 643.200 ;
        RECT 797.250 640.950 799.050 647.250 ;
        RECT 800.250 644.400 802.050 647.250 ;
        RECT 783.600 639.300 789.300 640.500 ;
        RECT 790.350 640.050 792.150 640.500 ;
        RECT 796.950 640.050 799.050 640.950 ;
        RECT 783.600 638.700 785.400 639.300 ;
        RECT 790.350 638.850 799.050 640.050 ;
        RECT 790.350 638.700 792.150 638.850 ;
        RECT 800.550 637.350 801.900 644.400 ;
        RECT 804.000 640.500 805.800 647.250 ;
        RECT 807.000 641.400 808.800 647.250 ;
        RECT 810.000 641.400 811.800 647.250 ;
        RECT 813.750 641.400 815.550 647.250 ;
        RECT 816.750 644.400 818.700 647.250 ;
        RECT 819.750 644.400 821.850 647.250 ;
        RECT 822.750 644.400 825.150 647.250 ;
        RECT 817.500 643.050 818.700 644.400 ;
        RECT 820.950 643.050 821.850 644.400 ;
        RECT 823.950 643.050 825.150 644.400 ;
        RECT 826.500 643.950 828.300 647.250 ;
        RECT 817.500 641.400 820.050 643.050 ;
        RECT 810.000 640.500 811.350 641.400 ;
        RECT 817.950 640.950 820.050 641.400 ;
        RECT 820.950 640.950 823.050 643.050 ;
        RECT 823.950 640.950 826.050 643.050 ;
        RECT 804.000 640.200 807.000 640.500 ;
        RECT 803.100 638.400 807.000 640.200 ;
        RECT 808.950 638.850 811.350 640.500 ;
        RECT 808.950 638.400 811.050 638.850 ;
        RECT 829.500 638.700 831.300 647.250 ;
        RECT 832.500 641.400 834.300 647.250 ;
        RECT 835.500 641.400 837.300 647.250 ;
        RECT 838.500 641.400 840.300 647.250 ;
        RECT 848.550 641.400 850.350 647.250 ;
        RECT 851.550 641.400 853.350 647.250 ;
        RECT 854.550 641.400 856.350 647.250 ;
        RECT 836.250 640.500 837.300 641.400 ;
        RECT 836.250 639.600 840.300 640.500 ;
        RECT 818.100 637.650 835.800 638.700 ;
        RECT 772.950 626.850 776.550 628.950 ;
        RECT 721.350 622.500 728.100 624.300 ;
        RECT 729.000 622.500 735.900 624.300 ;
        RECT 747.150 623.850 751.500 624.300 ;
        RECT 743.850 623.100 751.500 623.850 ;
        RECT 753.000 625.200 768.300 626.100 ;
        RECT 743.850 622.950 748.950 623.100 ;
        RECT 743.850 621.600 744.750 622.950 ;
        RECT 753.000 622.050 754.050 625.200 ;
        RECT 762.300 623.700 764.100 624.300 ;
        RECT 706.650 615.750 708.450 621.600 ;
        RECT 712.050 615.750 713.850 621.600 ;
        RECT 715.200 620.400 719.400 621.600 ;
        RECT 717.600 615.750 719.400 620.400 ;
        RECT 721.950 619.500 724.050 621.600 ;
        RECT 724.950 619.500 727.050 621.600 ;
        RECT 727.950 619.500 730.050 621.600 ;
        RECT 732.750 621.300 734.850 621.600 ;
        RECT 722.250 615.750 724.050 619.500 ;
        RECT 725.250 615.750 727.050 619.500 ;
        RECT 728.250 615.750 730.050 619.500 ;
        RECT 732.000 619.500 734.850 621.300 ;
        RECT 736.950 621.300 739.050 621.600 ;
        RECT 736.950 619.500 739.800 621.300 ;
        RECT 740.700 620.250 744.750 621.600 ;
        RECT 740.700 619.800 742.500 620.250 ;
        RECT 745.950 619.950 748.050 622.050 ;
        RECT 748.950 619.950 751.050 622.050 ;
        RECT 751.950 619.950 754.050 622.050 ;
        RECT 755.700 622.500 764.100 623.700 ;
        RECT 755.700 621.600 757.200 622.500 ;
        RECT 767.100 621.600 768.300 625.200 ;
        RECT 732.000 615.750 733.800 619.500 ;
        RECT 735.000 615.750 736.800 618.600 ;
        RECT 738.000 615.750 739.800 619.500 ;
        RECT 745.950 618.600 747.300 619.950 ;
        RECT 748.950 618.600 750.300 619.950 ;
        RECT 751.950 618.600 753.300 619.950 ;
        RECT 742.500 615.750 744.300 618.600 ;
        RECT 745.500 615.750 747.300 618.600 ;
        RECT 748.500 615.750 750.300 618.600 ;
        RECT 751.500 615.750 753.300 618.600 ;
        RECT 755.700 615.750 757.500 621.600 ;
        RECT 761.100 615.750 762.900 621.600 ;
        RECT 766.500 615.750 768.300 621.600 ;
        RECT 775.050 618.600 776.550 626.850 ;
        RECT 771.750 615.750 773.550 618.600 ;
        RECT 774.750 615.750 776.550 618.600 ;
        RECT 778.650 636.450 796.050 637.350 ;
        RECT 778.650 621.600 779.850 636.450 ;
        RECT 780.750 634.350 793.050 635.550 ;
        RECT 793.950 635.250 796.050 636.450 ;
        RECT 799.950 636.600 802.050 637.350 ;
        RECT 818.100 636.600 820.050 637.650 ;
        RECT 834.000 636.900 835.800 637.650 ;
        RECT 799.950 635.250 820.050 636.600 ;
        RECT 820.950 636.150 823.050 636.750 ;
        RECT 820.950 634.950 832.500 636.150 ;
        RECT 820.950 634.650 823.050 634.950 ;
        RECT 830.700 634.350 832.500 634.950 ;
        RECT 780.750 633.750 782.550 634.350 ;
        RECT 792.000 633.450 820.050 634.350 ;
        RECT 792.000 633.150 831.750 633.450 ;
        RECT 784.950 629.100 787.050 633.150 ;
        RECT 818.100 632.550 832.050 633.150 ;
        RECT 788.100 630.000 795.150 631.800 ;
        RECT 784.950 628.050 793.200 629.100 ;
        RECT 780.900 625.200 788.700 627.000 ;
        RECT 792.150 626.250 793.200 628.050 ;
        RECT 794.250 628.350 795.150 630.000 ;
        RECT 796.500 631.650 811.050 632.250 ;
        RECT 796.500 631.050 819.600 631.650 ;
        RECT 828.150 631.350 832.050 632.550 ;
        RECT 796.500 629.250 798.300 631.050 ;
        RECT 808.950 630.450 819.600 631.050 ;
        RECT 808.950 630.150 811.050 630.450 ;
        RECT 817.800 629.850 819.600 630.450 ;
        RECT 820.500 630.450 827.250 631.350 ;
        RECT 829.950 631.050 832.050 631.350 ;
        RECT 804.750 629.250 806.850 629.550 ;
        RECT 794.250 627.300 803.850 628.350 ;
        RECT 804.750 627.450 808.650 629.250 ;
        RECT 820.500 628.950 821.550 630.450 ;
        RECT 809.550 628.050 821.550 628.950 ;
        RECT 802.950 626.550 803.850 627.300 ;
        RECT 809.550 626.550 810.600 628.050 ;
        RECT 822.450 627.750 824.250 629.550 ;
        RECT 826.050 628.050 827.250 630.450 ;
        RECT 835.950 629.850 838.050 631.950 ;
        RECT 836.100 628.050 837.900 629.850 ;
        RECT 792.150 625.200 802.050 626.250 ;
        RECT 802.950 625.200 810.600 626.550 ;
        RECT 811.950 625.350 815.850 627.150 ;
        RECT 787.200 621.600 788.700 625.200 ;
        RECT 801.000 624.300 802.050 625.200 ;
        RECT 811.950 625.050 814.050 625.350 ;
        RECT 819.150 624.300 820.950 624.750 ;
        RECT 822.450 624.300 823.500 627.750 ;
        RECT 826.050 627.000 837.900 628.050 ;
        RECT 839.100 626.100 840.300 639.600 ;
        RECT 851.550 633.150 852.750 641.400 ;
        RECT 847.950 629.850 850.050 631.950 ;
        RECT 850.950 631.050 853.050 633.150 ;
        RECT 848.100 628.050 849.900 629.850 ;
        RECT 793.350 622.500 800.100 624.300 ;
        RECT 801.000 622.500 807.900 624.300 ;
        RECT 819.150 623.850 823.500 624.300 ;
        RECT 815.850 623.100 823.500 623.850 ;
        RECT 825.000 625.200 840.300 626.100 ;
        RECT 815.850 622.950 820.950 623.100 ;
        RECT 815.850 621.600 816.750 622.950 ;
        RECT 825.000 622.050 826.050 625.200 ;
        RECT 834.300 623.700 836.100 624.300 ;
        RECT 778.650 615.750 780.450 621.600 ;
        RECT 784.050 615.750 785.850 621.600 ;
        RECT 787.200 620.400 791.400 621.600 ;
        RECT 789.600 615.750 791.400 620.400 ;
        RECT 793.950 619.500 796.050 621.600 ;
        RECT 796.950 619.500 799.050 621.600 ;
        RECT 799.950 619.500 802.050 621.600 ;
        RECT 804.750 621.300 806.850 621.600 ;
        RECT 794.250 615.750 796.050 619.500 ;
        RECT 797.250 615.750 799.050 619.500 ;
        RECT 800.250 615.750 802.050 619.500 ;
        RECT 804.000 619.500 806.850 621.300 ;
        RECT 808.950 621.300 811.050 621.600 ;
        RECT 808.950 619.500 811.800 621.300 ;
        RECT 812.700 620.250 816.750 621.600 ;
        RECT 812.700 619.800 814.500 620.250 ;
        RECT 817.950 619.950 820.050 622.050 ;
        RECT 820.950 619.950 823.050 622.050 ;
        RECT 823.950 619.950 826.050 622.050 ;
        RECT 827.700 622.500 836.100 623.700 ;
        RECT 827.700 621.600 829.200 622.500 ;
        RECT 839.100 621.600 840.300 625.200 ;
        RECT 851.550 623.700 852.750 631.050 ;
        RECT 853.950 629.850 856.050 631.950 ;
        RECT 854.100 628.050 855.900 629.850 ;
        RECT 851.550 622.800 855.150 623.700 ;
        RECT 804.000 615.750 805.800 619.500 ;
        RECT 807.000 615.750 808.800 618.600 ;
        RECT 810.000 615.750 811.800 619.500 ;
        RECT 817.950 618.600 819.300 619.950 ;
        RECT 820.950 618.600 822.300 619.950 ;
        RECT 823.950 618.600 825.300 619.950 ;
        RECT 814.500 615.750 816.300 618.600 ;
        RECT 817.500 615.750 819.300 618.600 ;
        RECT 820.500 615.750 822.300 618.600 ;
        RECT 823.500 615.750 825.300 618.600 ;
        RECT 827.700 615.750 829.500 621.600 ;
        RECT 833.100 615.750 834.900 621.600 ;
        RECT 838.500 615.750 840.300 621.600 ;
        RECT 848.850 615.750 850.650 621.600 ;
        RECT 853.350 615.750 855.150 622.800 ;
        RECT 2.700 605.400 4.500 611.250 ;
        RECT 8.100 605.400 9.900 611.250 ;
        RECT 13.500 605.400 15.300 611.250 ;
        RECT 17.700 608.400 19.500 611.250 ;
        RECT 20.700 608.400 22.500 611.250 ;
        RECT 23.700 608.400 25.500 611.250 ;
        RECT 26.700 608.400 28.500 611.250 ;
        RECT 17.700 607.050 19.050 608.400 ;
        RECT 20.700 607.050 22.050 608.400 ;
        RECT 23.700 607.050 25.050 608.400 ;
        RECT 31.200 607.500 33.000 611.250 ;
        RECT 34.200 608.400 36.000 611.250 ;
        RECT 37.200 607.500 39.000 611.250 ;
        RECT 2.700 601.800 3.900 605.400 ;
        RECT 13.800 604.500 15.300 605.400 ;
        RECT 6.900 603.300 15.300 604.500 ;
        RECT 16.950 604.950 19.050 607.050 ;
        RECT 19.950 604.950 22.050 607.050 ;
        RECT 22.950 604.950 25.050 607.050 ;
        RECT 28.500 606.750 30.300 607.200 ;
        RECT 26.250 605.400 30.300 606.750 ;
        RECT 31.200 605.700 34.050 607.500 ;
        RECT 31.950 605.400 34.050 605.700 ;
        RECT 36.150 605.700 39.000 607.500 ;
        RECT 40.950 607.500 42.750 611.250 ;
        RECT 43.950 607.500 45.750 611.250 ;
        RECT 46.950 607.500 48.750 611.250 ;
        RECT 36.150 605.400 38.250 605.700 ;
        RECT 40.950 605.400 43.050 607.500 ;
        RECT 43.950 605.400 46.050 607.500 ;
        RECT 46.950 605.400 49.050 607.500 ;
        RECT 51.600 606.600 53.400 611.250 ;
        RECT 51.600 605.400 55.800 606.600 ;
        RECT 57.150 605.400 58.950 611.250 ;
        RECT 62.550 605.400 64.350 611.250 ;
        RECT 6.900 602.700 8.700 603.300 ;
        RECT 16.950 601.800 18.000 604.950 ;
        RECT 26.250 604.050 27.150 605.400 ;
        RECT 22.050 603.900 27.150 604.050 ;
        RECT 2.700 600.900 18.000 601.800 ;
        RECT 19.500 603.150 27.150 603.900 ;
        RECT 19.500 602.700 23.850 603.150 ;
        RECT 35.100 602.700 42.000 604.500 ;
        RECT 42.900 602.700 49.650 604.500 ;
        RECT 2.700 587.400 3.900 600.900 ;
        RECT 5.100 598.950 16.950 600.000 ;
        RECT 19.500 599.250 20.550 602.700 ;
        RECT 22.050 602.250 23.850 602.700 ;
        RECT 28.950 601.650 31.050 601.950 ;
        RECT 40.950 601.800 42.000 602.700 ;
        RECT 54.300 601.800 55.800 605.400 ;
        RECT 27.150 599.850 31.050 601.650 ;
        RECT 32.400 600.450 40.050 601.800 ;
        RECT 40.950 600.750 50.850 601.800 ;
        RECT 5.100 597.150 6.900 598.950 ;
        RECT 4.950 595.050 7.050 597.150 ;
        RECT 15.750 596.550 16.950 598.950 ;
        RECT 18.750 597.450 20.550 599.250 ;
        RECT 32.400 598.950 33.450 600.450 ;
        RECT 39.150 599.700 40.050 600.450 ;
        RECT 21.450 598.050 33.450 598.950 ;
        RECT 21.450 596.550 22.500 598.050 ;
        RECT 34.350 597.750 38.250 599.550 ;
        RECT 39.150 598.650 48.750 599.700 ;
        RECT 36.150 597.450 38.250 597.750 ;
        RECT 10.950 595.650 13.050 595.950 ;
        RECT 15.750 595.650 22.500 596.550 ;
        RECT 23.400 596.550 25.200 597.150 ;
        RECT 31.950 596.550 34.050 596.850 ;
        RECT 23.400 595.950 34.050 596.550 ;
        RECT 44.700 595.950 46.500 597.750 ;
        RECT 10.950 594.450 14.850 595.650 ;
        RECT 23.400 595.350 46.500 595.950 ;
        RECT 31.950 594.750 46.500 595.350 ;
        RECT 47.850 597.000 48.750 598.650 ;
        RECT 49.800 598.950 50.850 600.750 ;
        RECT 54.300 600.000 62.100 601.800 ;
        RECT 49.800 597.900 58.050 598.950 ;
        RECT 47.850 595.200 54.900 597.000 ;
        RECT 10.950 593.850 24.900 594.450 ;
        RECT 55.950 593.850 58.050 597.900 ;
        RECT 11.250 593.550 51.000 593.850 ;
        RECT 22.950 592.650 51.000 593.550 ;
        RECT 60.450 592.650 62.250 593.250 ;
        RECT 10.500 592.050 12.300 592.650 ;
        RECT 19.950 592.050 22.050 592.350 ;
        RECT 10.500 590.850 22.050 592.050 ;
        RECT 19.950 590.250 22.050 590.850 ;
        RECT 22.950 590.400 43.050 591.750 ;
        RECT 7.200 589.350 9.000 590.100 ;
        RECT 22.950 589.350 24.900 590.400 ;
        RECT 40.950 589.650 43.050 590.400 ;
        RECT 46.950 590.550 49.050 591.750 ;
        RECT 49.950 591.450 62.250 592.650 ;
        RECT 63.150 590.550 64.350 605.400 ;
        RECT 46.950 589.650 64.350 590.550 ;
        RECT 66.450 608.400 68.250 611.250 ;
        RECT 69.450 608.400 71.250 611.250 ;
        RECT 79.650 608.400 81.450 611.250 ;
        RECT 82.650 608.400 84.450 611.250 ;
        RECT 85.650 608.400 87.450 611.250 ;
        RECT 92.550 608.400 94.350 611.250 ;
        RECT 95.550 608.400 97.350 611.250 ;
        RECT 66.450 600.150 67.950 608.400 ;
        RECT 82.950 601.950 84.000 608.400 ;
        RECT 85.950 603.450 88.050 604.050 ;
        RECT 85.950 602.550 90.450 603.450 ;
        RECT 85.950 601.950 88.050 602.550 ;
        RECT 66.450 598.050 70.050 600.150 ;
        RECT 82.950 599.850 85.050 601.950 ;
        RECT 7.200 588.300 24.900 589.350 ;
        RECT 2.700 586.500 6.750 587.400 ;
        RECT 5.700 585.600 6.750 586.500 ;
        RECT 2.700 579.750 4.500 585.600 ;
        RECT 5.700 579.750 7.500 585.600 ;
        RECT 8.700 579.750 10.500 585.600 ;
        RECT 11.700 579.750 13.500 588.300 ;
        RECT 31.950 588.150 34.050 588.600 ;
        RECT 31.650 586.500 34.050 588.150 ;
        RECT 36.000 586.800 39.900 588.600 ;
        RECT 36.000 586.500 39.000 586.800 ;
        RECT 16.950 583.950 19.050 586.050 ;
        RECT 19.950 583.950 22.050 586.050 ;
        RECT 22.950 585.600 25.050 586.050 ;
        RECT 31.650 585.600 33.000 586.500 ;
        RECT 22.950 583.950 25.500 585.600 ;
        RECT 14.700 579.750 16.500 583.050 ;
        RECT 17.850 582.600 19.050 583.950 ;
        RECT 21.150 582.600 22.050 583.950 ;
        RECT 24.300 582.600 25.500 583.950 ;
        RECT 17.850 579.750 20.250 582.600 ;
        RECT 21.150 579.750 23.250 582.600 ;
        RECT 24.300 579.750 26.250 582.600 ;
        RECT 27.450 579.750 29.250 585.600 ;
        RECT 31.200 579.750 33.000 585.600 ;
        RECT 34.200 579.750 36.000 585.600 ;
        RECT 37.200 579.750 39.000 586.500 ;
        RECT 41.100 582.600 42.450 589.650 ;
        RECT 50.850 588.150 52.650 588.300 ;
        RECT 43.950 586.950 52.650 588.150 ;
        RECT 57.600 587.700 59.400 588.300 ;
        RECT 43.950 586.050 46.050 586.950 ;
        RECT 50.850 586.500 52.650 586.950 ;
        RECT 53.700 586.500 59.400 587.700 ;
        RECT 40.950 579.750 42.750 582.600 ;
        RECT 43.950 579.750 45.750 586.050 ;
        RECT 47.100 583.800 49.200 585.900 ;
        RECT 47.100 582.600 48.600 583.800 ;
        RECT 46.950 579.750 48.750 582.600 ;
        RECT 50.700 579.750 52.500 585.600 ;
        RECT 53.700 579.750 55.500 586.500 ;
        RECT 60.300 585.600 61.500 589.650 ;
        RECT 66.450 585.600 67.950 598.050 ;
        RECT 79.950 596.850 82.050 598.950 ;
        RECT 80.100 595.050 81.900 596.850 ;
        RECT 82.950 592.650 84.000 599.850 ;
        RECT 85.950 596.850 88.050 598.950 ;
        RECT 86.100 595.050 87.900 596.850 ;
        RECT 89.550 594.450 90.450 602.550 ;
        RECT 91.950 599.850 94.050 601.950 ;
        RECT 95.400 600.150 96.600 608.400 ;
        RECT 103.350 605.400 105.150 611.250 ;
        RECT 106.350 605.400 108.150 611.250 ;
        RECT 109.650 608.400 111.450 611.250 ;
        RECT 118.650 608.400 120.450 611.250 ;
        RECT 121.650 608.400 123.450 611.250 ;
        RECT 124.650 608.400 126.450 611.250 ;
        RECT 130.650 608.400 132.450 611.250 ;
        RECT 133.650 608.400 135.450 611.250 ;
        RECT 136.650 608.400 138.450 611.250 ;
        RECT 140.550 608.400 142.350 611.250 ;
        RECT 143.550 608.400 145.350 611.250 ;
        RECT 152.550 608.400 154.350 611.250 ;
        RECT 155.550 608.400 157.350 611.250 ;
        RECT 158.550 608.400 160.350 611.250 ;
        RECT 92.100 598.050 93.900 599.850 ;
        RECT 94.950 598.050 97.050 600.150 ;
        RECT 103.650 598.950 104.850 605.400 ;
        RECT 109.650 604.500 110.850 608.400 ;
        RECT 105.750 603.600 110.850 604.500 ;
        RECT 105.750 602.700 108.000 603.600 ;
        RECT 91.950 594.450 94.050 595.050 ;
        RECT 89.550 593.550 94.050 594.450 ;
        RECT 91.950 592.950 94.050 593.550 ;
        RECT 81.450 591.600 84.000 592.650 ;
        RECT 56.700 579.750 58.500 585.600 ;
        RECT 59.700 579.750 61.500 585.600 ;
        RECT 62.700 579.750 64.500 585.600 ;
        RECT 66.450 579.750 68.250 585.600 ;
        RECT 69.450 579.750 71.250 585.600 ;
        RECT 81.450 579.750 83.250 591.600 ;
        RECT 85.650 579.750 87.450 591.600 ;
        RECT 95.400 585.600 96.600 598.050 ;
        RECT 103.650 596.850 106.050 598.950 ;
        RECT 103.650 591.600 104.850 596.850 ;
        RECT 106.950 594.300 108.000 602.700 ;
        RECT 121.950 601.950 123.000 608.400 ;
        RECT 133.950 601.950 135.000 608.400 ;
        RECT 121.950 599.850 124.050 601.950 ;
        RECT 133.950 599.850 136.050 601.950 ;
        RECT 139.950 599.850 142.050 601.950 ;
        RECT 143.400 600.150 144.600 608.400 ;
        RECT 156.000 601.950 157.050 608.400 ;
        RECT 173.850 604.200 175.650 611.250 ;
        RECT 178.350 605.400 180.150 611.250 ;
        RECT 182.550 608.400 184.350 611.250 ;
        RECT 185.550 608.400 187.350 611.250 ;
        RECT 199.650 608.400 201.450 611.250 ;
        RECT 202.650 608.400 204.450 611.250 ;
        RECT 205.650 608.400 207.450 611.250 ;
        RECT 211.650 608.400 213.450 611.250 ;
        RECT 214.650 608.400 216.450 611.250 ;
        RECT 217.650 608.400 219.450 611.250 ;
        RECT 173.850 603.300 177.450 604.200 ;
        RECT 109.950 596.850 112.050 598.950 ;
        RECT 118.950 596.850 121.050 598.950 ;
        RECT 110.100 595.050 111.900 596.850 ;
        RECT 119.100 595.050 120.900 596.850 ;
        RECT 105.750 593.400 108.000 594.300 ;
        RECT 105.750 592.500 111.450 593.400 ;
        RECT 121.950 592.650 123.000 599.850 ;
        RECT 124.950 596.850 127.050 598.950 ;
        RECT 130.950 596.850 133.050 598.950 ;
        RECT 125.100 595.050 126.900 596.850 ;
        RECT 131.100 595.050 132.900 596.850 ;
        RECT 133.950 592.650 135.000 599.850 ;
        RECT 136.950 596.850 139.050 598.950 ;
        RECT 140.100 598.050 141.900 599.850 ;
        RECT 142.950 598.050 145.050 600.150 ;
        RECT 154.950 599.850 157.050 601.950 ;
        RECT 137.100 595.050 138.900 596.850 ;
        RECT 92.550 579.750 94.350 585.600 ;
        RECT 95.550 579.750 97.350 585.600 ;
        RECT 103.350 579.750 105.150 591.600 ;
        RECT 106.350 579.750 108.150 591.600 ;
        RECT 110.250 585.600 111.450 592.500 ;
        RECT 109.650 579.750 111.450 585.600 ;
        RECT 120.450 591.600 123.000 592.650 ;
        RECT 132.450 591.600 135.000 592.650 ;
        RECT 120.450 579.750 122.250 591.600 ;
        RECT 124.650 579.750 126.450 591.600 ;
        RECT 132.450 579.750 134.250 591.600 ;
        RECT 136.650 579.750 138.450 591.600 ;
        RECT 143.400 585.600 144.600 598.050 ;
        RECT 151.950 596.850 154.050 598.950 ;
        RECT 152.100 595.050 153.900 596.850 ;
        RECT 156.000 592.650 157.050 599.850 ;
        RECT 157.950 596.850 160.050 598.950 ;
        RECT 173.100 597.150 174.900 598.950 ;
        RECT 158.100 595.050 159.900 596.850 ;
        RECT 172.950 595.050 175.050 597.150 ;
        RECT 176.250 595.950 177.450 603.300 ;
        RECT 181.950 599.850 184.050 601.950 ;
        RECT 185.400 600.150 186.600 608.400 ;
        RECT 202.950 601.950 204.000 608.400 ;
        RECT 214.950 601.950 216.000 608.400 ;
        RECT 229.650 605.400 231.450 611.250 ;
        RECT 230.250 603.300 231.450 605.400 ;
        RECT 232.650 606.300 234.450 611.250 ;
        RECT 235.650 607.200 237.450 611.250 ;
        RECT 238.650 606.300 240.450 611.250 ;
        RECT 232.650 604.950 240.450 606.300 ;
        RECT 250.650 605.400 252.450 611.250 ;
        RECT 251.250 603.300 252.450 605.400 ;
        RECT 253.650 606.300 255.450 611.250 ;
        RECT 256.650 607.200 258.450 611.250 ;
        RECT 259.650 606.300 261.450 611.250 ;
        RECT 253.650 604.950 261.450 606.300 ;
        RECT 274.800 605.400 276.600 611.250 ;
        RECT 279.000 605.400 280.800 611.250 ;
        RECT 283.200 605.400 285.000 611.250 ;
        RECT 293.550 608.400 295.350 611.250 ;
        RECT 296.550 608.400 298.350 611.250 ;
        RECT 299.550 608.400 301.350 611.250 ;
        RECT 230.250 602.250 234.000 603.300 ;
        RECT 251.250 602.250 255.000 603.300 ;
        RECT 179.100 597.150 180.900 598.950 ;
        RECT 182.100 598.050 183.900 599.850 ;
        RECT 184.950 598.050 187.050 600.150 ;
        RECT 202.950 599.850 205.050 601.950 ;
        RECT 214.950 599.850 217.050 601.950 ;
        RECT 175.950 593.850 178.050 595.950 ;
        RECT 178.950 595.050 181.050 597.150 ;
        RECT 156.000 591.600 158.550 592.650 ;
        RECT 140.550 579.750 142.350 585.600 ;
        RECT 143.550 579.750 145.350 585.600 ;
        RECT 152.550 579.750 154.350 591.600 ;
        RECT 156.750 579.750 158.550 591.600 ;
        RECT 176.250 585.600 177.450 593.850 ;
        RECT 185.400 585.600 186.600 598.050 ;
        RECT 199.950 596.850 202.050 598.950 ;
        RECT 200.100 595.050 201.900 596.850 ;
        RECT 202.950 592.650 204.000 599.850 ;
        RECT 205.950 596.850 208.050 598.950 ;
        RECT 211.950 596.850 214.050 598.950 ;
        RECT 206.100 595.050 207.900 596.850 ;
        RECT 212.100 595.050 213.900 596.850 ;
        RECT 214.950 592.650 216.000 599.850 ;
        RECT 232.950 598.950 234.150 602.250 ;
        RECT 236.100 600.150 237.900 601.950 ;
        RECT 217.950 596.850 220.050 598.950 ;
        RECT 232.950 596.850 235.050 598.950 ;
        RECT 235.950 598.050 238.050 600.150 ;
        RECT 253.950 598.950 255.150 602.250 ;
        RECT 257.100 600.150 258.900 601.950 ;
        RECT 275.250 600.150 277.050 601.950 ;
        RECT 238.950 596.850 241.050 598.950 ;
        RECT 253.950 596.850 256.050 598.950 ;
        RECT 256.950 598.050 259.050 600.150 ;
        RECT 259.950 596.850 262.050 598.950 ;
        RECT 271.950 596.850 274.050 598.950 ;
        RECT 274.950 598.050 277.050 600.150 ;
        RECT 279.000 598.950 280.050 605.400 ;
        RECT 297.000 601.950 298.050 608.400 ;
        RECT 308.850 605.400 310.650 611.250 ;
        RECT 313.350 604.200 315.150 611.250 ;
        RECT 320.550 608.400 322.350 611.250 ;
        RECT 323.550 608.400 325.350 611.250 ;
        RECT 277.950 596.850 280.050 598.950 ;
        RECT 280.950 600.150 282.750 601.950 ;
        RECT 280.950 598.050 283.050 600.150 ;
        RECT 295.950 599.850 298.050 601.950 ;
        RECT 283.950 596.850 286.050 598.950 ;
        RECT 292.950 596.850 295.050 598.950 ;
        RECT 218.100 595.050 219.900 596.850 ;
        RECT 229.950 593.850 232.050 595.950 ;
        RECT 201.450 591.600 204.000 592.650 ;
        RECT 213.450 591.600 216.000 592.650 ;
        RECT 230.250 592.050 232.050 593.850 ;
        RECT 233.850 591.600 235.050 596.850 ;
        RECT 239.100 595.050 240.900 596.850 ;
        RECT 250.950 593.850 253.050 595.950 ;
        RECT 251.250 592.050 253.050 593.850 ;
        RECT 254.850 591.600 256.050 596.850 ;
        RECT 260.100 595.050 261.900 596.850 ;
        RECT 272.100 595.050 273.900 596.850 ;
        RECT 277.950 593.400 278.850 596.850 ;
        RECT 283.950 595.050 285.750 596.850 ;
        RECT 293.100 595.050 294.900 596.850 ;
        RECT 274.800 592.500 278.850 593.400 ;
        RECT 297.000 592.650 298.050 599.850 ;
        RECT 311.550 603.300 315.150 604.200 ;
        RECT 298.950 596.850 301.050 598.950 ;
        RECT 308.100 597.150 309.900 598.950 ;
        RECT 299.100 595.050 300.900 596.850 ;
        RECT 307.950 595.050 310.050 597.150 ;
        RECT 311.550 595.950 312.750 603.300 ;
        RECT 319.950 599.850 322.050 601.950 ;
        RECT 323.400 600.150 324.600 608.400 ;
        RECT 335.550 606.300 337.350 611.250 ;
        RECT 338.550 607.200 340.350 611.250 ;
        RECT 341.550 606.300 343.350 611.250 ;
        RECT 335.550 604.950 343.350 606.300 ;
        RECT 344.550 605.400 346.350 611.250 ;
        RECT 350.850 605.400 352.650 611.250 ;
        RECT 344.550 603.300 345.750 605.400 ;
        RECT 355.350 604.200 357.150 611.250 ;
        RECT 368.550 608.400 370.350 611.250 ;
        RECT 371.550 608.400 373.350 611.250 ;
        RECT 374.550 608.400 376.350 611.250 ;
        RECT 380.550 608.400 382.350 611.250 ;
        RECT 383.550 608.400 385.350 611.250 ;
        RECT 397.650 608.400 399.450 611.250 ;
        RECT 400.650 608.400 402.450 611.250 ;
        RECT 342.000 602.250 345.750 603.300 ;
        RECT 353.550 603.300 357.150 604.200 ;
        RECT 338.100 600.150 339.900 601.950 ;
        RECT 314.100 597.150 315.900 598.950 ;
        RECT 320.100 598.050 321.900 599.850 ;
        RECT 322.950 598.050 325.050 600.150 ;
        RECT 310.950 593.850 313.050 595.950 ;
        RECT 313.950 595.050 316.050 597.150 ;
        RECT 274.800 591.600 276.600 592.500 ;
        RECT 297.000 591.600 299.550 592.650 ;
        RECT 172.650 579.750 174.450 585.600 ;
        RECT 175.650 579.750 177.450 585.600 ;
        RECT 178.650 579.750 180.450 585.600 ;
        RECT 182.550 579.750 184.350 585.600 ;
        RECT 185.550 579.750 187.350 585.600 ;
        RECT 201.450 579.750 203.250 591.600 ;
        RECT 205.650 579.750 207.450 591.600 ;
        RECT 213.450 579.750 215.250 591.600 ;
        RECT 217.650 579.750 219.450 591.600 ;
        RECT 230.400 579.750 232.200 585.600 ;
        RECT 233.700 579.750 235.500 591.600 ;
        RECT 237.900 579.750 239.700 591.600 ;
        RECT 251.400 579.750 253.200 585.600 ;
        RECT 254.700 579.750 256.500 591.600 ;
        RECT 258.900 579.750 260.700 591.600 ;
        RECT 271.650 580.500 273.450 591.600 ;
        RECT 274.650 581.400 276.450 591.600 ;
        RECT 277.650 590.400 285.450 591.300 ;
        RECT 277.650 580.500 279.450 590.400 ;
        RECT 271.650 579.750 279.450 580.500 ;
        RECT 280.650 579.750 282.450 589.500 ;
        RECT 283.650 579.750 285.450 590.400 ;
        RECT 293.550 579.750 295.350 591.600 ;
        RECT 297.750 579.750 299.550 591.600 ;
        RECT 311.550 585.600 312.750 593.850 ;
        RECT 323.400 585.600 324.600 598.050 ;
        RECT 334.950 596.850 337.050 598.950 ;
        RECT 337.950 598.050 340.050 600.150 ;
        RECT 341.850 598.950 343.050 602.250 ;
        RECT 340.950 596.850 343.050 598.950 ;
        RECT 350.100 597.150 351.900 598.950 ;
        RECT 335.100 595.050 336.900 596.850 ;
        RECT 340.950 591.600 342.150 596.850 ;
        RECT 343.950 593.850 346.050 595.950 ;
        RECT 349.950 595.050 352.050 597.150 ;
        RECT 353.550 595.950 354.750 603.300 ;
        RECT 372.000 601.950 373.050 608.400 ;
        RECT 370.950 599.850 373.050 601.950 ;
        RECT 379.950 599.850 382.050 601.950 ;
        RECT 383.400 600.150 384.600 608.400 ;
        RECT 398.400 600.150 399.600 608.400 ;
        RECT 410.100 603.000 411.900 611.250 ;
        RECT 356.100 597.150 357.900 598.950 ;
        RECT 352.950 593.850 355.050 595.950 ;
        RECT 355.950 595.050 358.050 597.150 ;
        RECT 367.950 596.850 370.050 598.950 ;
        RECT 368.100 595.050 369.900 596.850 ;
        RECT 343.950 592.050 345.750 593.850 ;
        RECT 308.550 579.750 310.350 585.600 ;
        RECT 311.550 579.750 313.350 585.600 ;
        RECT 314.550 579.750 316.350 585.600 ;
        RECT 320.550 579.750 322.350 585.600 ;
        RECT 323.550 579.750 325.350 585.600 ;
        RECT 336.300 579.750 338.100 591.600 ;
        RECT 340.500 579.750 342.300 591.600 ;
        RECT 353.550 585.600 354.750 593.850 ;
        RECT 372.000 592.650 373.050 599.850 ;
        RECT 373.950 596.850 376.050 598.950 ;
        RECT 380.100 598.050 381.900 599.850 ;
        RECT 382.950 598.050 385.050 600.150 ;
        RECT 397.950 598.050 400.050 600.150 ;
        RECT 400.950 599.850 403.050 601.950 ;
        RECT 407.400 601.350 411.900 603.000 ;
        RECT 415.500 602.400 417.300 611.250 ;
        RECT 422.550 606.300 424.350 611.250 ;
        RECT 425.550 607.200 427.350 611.250 ;
        RECT 428.550 606.300 430.350 611.250 ;
        RECT 422.550 604.950 430.350 606.300 ;
        RECT 431.550 605.400 433.350 611.250 ;
        RECT 445.650 608.400 447.450 611.250 ;
        RECT 448.650 608.400 450.450 611.250 ;
        RECT 431.550 603.300 432.750 605.400 ;
        RECT 429.000 602.250 432.750 603.300 ;
        RECT 401.100 598.050 402.900 599.850 ;
        RECT 374.100 595.050 375.900 596.850 ;
        RECT 372.000 591.600 374.550 592.650 ;
        RECT 343.800 579.750 345.600 585.600 ;
        RECT 350.550 579.750 352.350 585.600 ;
        RECT 353.550 579.750 355.350 585.600 ;
        RECT 356.550 579.750 358.350 585.600 ;
        RECT 368.550 579.750 370.350 591.600 ;
        RECT 372.750 579.750 374.550 591.600 ;
        RECT 383.400 585.600 384.600 598.050 ;
        RECT 398.400 585.600 399.600 598.050 ;
        RECT 407.400 597.150 408.600 601.350 ;
        RECT 412.950 600.450 415.050 601.050 ;
        RECT 418.950 600.450 421.050 601.050 ;
        RECT 412.950 599.550 421.050 600.450 ;
        RECT 425.100 600.150 426.900 601.950 ;
        RECT 412.950 598.950 415.050 599.550 ;
        RECT 418.950 598.950 421.050 599.550 ;
        RECT 406.950 595.050 409.050 597.150 ;
        RECT 421.950 596.850 424.050 598.950 ;
        RECT 424.950 598.050 427.050 600.150 ;
        RECT 428.850 598.950 430.050 602.250 ;
        RECT 446.400 600.150 447.600 608.400 ;
        RECT 452.850 605.400 454.650 611.250 ;
        RECT 457.350 604.200 459.150 611.250 ;
        RECT 470.550 608.400 472.350 611.250 ;
        RECT 473.550 608.400 475.350 611.250 ;
        RECT 481.650 608.400 483.450 611.250 ;
        RECT 484.650 608.400 486.450 611.250 ;
        RECT 455.550 603.300 459.150 604.200 ;
        RECT 427.950 596.850 430.050 598.950 ;
        RECT 445.950 598.050 448.050 600.150 ;
        RECT 448.950 599.850 451.050 601.950 ;
        RECT 449.100 598.050 450.900 599.850 ;
        RECT 407.250 586.800 408.300 595.050 ;
        RECT 409.950 593.850 412.050 595.950 ;
        RECT 415.950 593.850 418.050 595.950 ;
        RECT 422.100 595.050 423.900 596.850 ;
        RECT 409.950 592.050 411.750 593.850 ;
        RECT 412.950 590.850 415.050 592.950 ;
        RECT 416.100 592.050 417.900 593.850 ;
        RECT 427.950 591.600 429.150 596.850 ;
        RECT 430.950 593.850 433.050 595.950 ;
        RECT 430.950 592.050 432.750 593.850 ;
        RECT 413.100 589.050 414.900 590.850 ;
        RECT 407.250 585.900 414.300 586.800 ;
        RECT 407.250 585.600 408.450 585.900 ;
        RECT 380.550 579.750 382.350 585.600 ;
        RECT 383.550 579.750 385.350 585.600 ;
        RECT 397.650 579.750 399.450 585.600 ;
        RECT 400.650 579.750 402.450 585.600 ;
        RECT 406.650 579.750 408.450 585.600 ;
        RECT 412.650 585.600 414.300 585.900 ;
        RECT 409.650 579.750 411.450 585.000 ;
        RECT 412.650 579.750 414.450 585.600 ;
        RECT 415.650 579.750 417.450 585.600 ;
        RECT 423.300 579.750 425.100 591.600 ;
        RECT 427.500 579.750 429.300 591.600 ;
        RECT 446.400 585.600 447.600 598.050 ;
        RECT 452.100 597.150 453.900 598.950 ;
        RECT 451.950 595.050 454.050 597.150 ;
        RECT 455.550 595.950 456.750 603.300 ;
        RECT 469.950 599.850 472.050 601.950 ;
        RECT 473.400 600.150 474.600 608.400 ;
        RECT 482.400 600.150 483.600 608.400 ;
        RECT 488.700 602.400 490.500 611.250 ;
        RECT 494.100 603.000 495.900 611.250 ;
        RECT 458.100 597.150 459.900 598.950 ;
        RECT 470.100 598.050 471.900 599.850 ;
        RECT 472.950 598.050 475.050 600.150 ;
        RECT 481.950 598.050 484.050 600.150 ;
        RECT 484.950 599.850 487.050 601.950 ;
        RECT 494.100 601.350 498.600 603.000 ;
        RECT 503.700 602.400 505.500 611.250 ;
        RECT 509.100 603.000 510.900 611.250 ;
        RECT 518.850 605.400 520.650 611.250 ;
        RECT 523.350 604.200 525.150 611.250 ;
        RECT 532.650 608.400 534.450 611.250 ;
        RECT 535.650 608.400 537.450 611.250 ;
        RECT 538.650 608.400 540.450 611.250 ;
        RECT 548.550 608.400 550.350 611.250 ;
        RECT 551.550 608.400 553.350 611.250 ;
        RECT 562.650 608.400 564.450 611.250 ;
        RECT 565.650 608.400 567.450 611.250 ;
        RECT 568.650 608.400 570.450 611.250 ;
        RECT 521.550 603.300 525.150 604.200 ;
        RECT 509.100 601.350 513.600 603.000 ;
        RECT 485.100 598.050 486.900 599.850 ;
        RECT 454.950 593.850 457.050 595.950 ;
        RECT 457.950 595.050 460.050 597.150 ;
        RECT 455.550 585.600 456.750 593.850 ;
        RECT 473.400 585.600 474.600 598.050 ;
        RECT 482.400 585.600 483.600 598.050 ;
        RECT 497.400 597.150 498.600 601.350 ;
        RECT 512.400 597.150 513.600 601.350 ;
        RECT 518.100 597.150 519.900 598.950 ;
        RECT 487.950 593.850 490.050 595.950 ;
        RECT 493.950 593.850 496.050 595.950 ;
        RECT 496.950 595.050 499.050 597.150 ;
        RECT 488.100 592.050 489.900 593.850 ;
        RECT 490.950 590.850 493.050 592.950 ;
        RECT 494.250 592.050 496.050 593.850 ;
        RECT 491.100 589.050 492.900 590.850 ;
        RECT 497.700 586.800 498.750 595.050 ;
        RECT 502.950 593.850 505.050 595.950 ;
        RECT 508.950 593.850 511.050 595.950 ;
        RECT 511.950 595.050 514.050 597.150 ;
        RECT 517.950 595.050 520.050 597.150 ;
        RECT 521.550 595.950 522.750 603.300 ;
        RECT 535.950 601.950 537.000 608.400 ;
        RECT 535.950 599.850 538.050 601.950 ;
        RECT 547.950 599.850 550.050 601.950 ;
        RECT 551.400 600.150 552.600 608.400 ;
        RECT 565.950 601.950 567.000 608.400 ;
        RECT 572.550 606.300 574.350 611.250 ;
        RECT 575.550 607.200 577.350 611.250 ;
        RECT 578.550 606.300 580.350 611.250 ;
        RECT 572.550 604.950 580.350 606.300 ;
        RECT 581.550 605.400 583.350 611.250 ;
        RECT 595.650 608.400 597.450 611.250 ;
        RECT 598.650 608.400 600.450 611.250 ;
        RECT 581.550 603.300 582.750 605.400 ;
        RECT 579.000 602.250 582.750 603.300 ;
        RECT 524.100 597.150 525.900 598.950 ;
        RECT 503.100 592.050 504.900 593.850 ;
        RECT 505.950 590.850 508.050 592.950 ;
        RECT 509.250 592.050 511.050 593.850 ;
        RECT 506.100 589.050 507.900 590.850 ;
        RECT 512.700 586.800 513.750 595.050 ;
        RECT 520.950 593.850 523.050 595.950 ;
        RECT 523.950 595.050 526.050 597.150 ;
        RECT 532.950 596.850 535.050 598.950 ;
        RECT 533.100 595.050 534.900 596.850 ;
        RECT 491.700 585.900 498.750 586.800 ;
        RECT 491.700 585.600 493.350 585.900 ;
        RECT 430.800 579.750 432.600 585.600 ;
        RECT 445.650 579.750 447.450 585.600 ;
        RECT 448.650 579.750 450.450 585.600 ;
        RECT 452.550 579.750 454.350 585.600 ;
        RECT 455.550 579.750 457.350 585.600 ;
        RECT 458.550 579.750 460.350 585.600 ;
        RECT 470.550 579.750 472.350 585.600 ;
        RECT 473.550 579.750 475.350 585.600 ;
        RECT 481.650 579.750 483.450 585.600 ;
        RECT 484.650 579.750 486.450 585.600 ;
        RECT 488.550 579.750 490.350 585.600 ;
        RECT 491.550 579.750 493.350 585.600 ;
        RECT 497.550 585.600 498.750 585.900 ;
        RECT 506.700 585.900 513.750 586.800 ;
        RECT 506.700 585.600 508.350 585.900 ;
        RECT 494.550 579.750 496.350 585.000 ;
        RECT 497.550 579.750 499.350 585.600 ;
        RECT 503.550 579.750 505.350 585.600 ;
        RECT 506.550 579.750 508.350 585.600 ;
        RECT 512.550 585.600 513.750 585.900 ;
        RECT 521.550 585.600 522.750 593.850 ;
        RECT 535.950 592.650 537.000 599.850 ;
        RECT 538.950 596.850 541.050 598.950 ;
        RECT 548.100 598.050 549.900 599.850 ;
        RECT 550.950 598.050 553.050 600.150 ;
        RECT 565.950 599.850 568.050 601.950 ;
        RECT 575.100 600.150 576.900 601.950 ;
        RECT 539.100 595.050 540.900 596.850 ;
        RECT 534.450 591.600 537.000 592.650 ;
        RECT 509.550 579.750 511.350 585.000 ;
        RECT 512.550 579.750 514.350 585.600 ;
        RECT 518.550 579.750 520.350 585.600 ;
        RECT 521.550 579.750 523.350 585.600 ;
        RECT 524.550 579.750 526.350 585.600 ;
        RECT 534.450 579.750 536.250 591.600 ;
        RECT 538.650 579.750 540.450 591.600 ;
        RECT 551.400 585.600 552.600 598.050 ;
        RECT 562.950 596.850 565.050 598.950 ;
        RECT 563.100 595.050 564.900 596.850 ;
        RECT 565.950 592.650 567.000 599.850 ;
        RECT 568.950 596.850 571.050 598.950 ;
        RECT 571.950 596.850 574.050 598.950 ;
        RECT 574.950 598.050 577.050 600.150 ;
        RECT 578.850 598.950 580.050 602.250 ;
        RECT 596.400 600.150 597.600 608.400 ;
        RECT 608.850 605.400 610.650 611.250 ;
        RECT 613.350 604.200 615.150 611.250 ;
        RECT 626.850 605.400 628.650 611.250 ;
        RECT 631.350 604.200 633.150 611.250 ;
        RECT 611.550 603.300 615.150 604.200 ;
        RECT 629.550 603.300 633.150 604.200 ;
        RECT 577.950 596.850 580.050 598.950 ;
        RECT 595.950 598.050 598.050 600.150 ;
        RECT 598.950 599.850 601.050 601.950 ;
        RECT 599.100 598.050 600.900 599.850 ;
        RECT 569.100 595.050 570.900 596.850 ;
        RECT 572.100 595.050 573.900 596.850 ;
        RECT 564.450 591.600 567.000 592.650 ;
        RECT 577.950 591.600 579.150 596.850 ;
        RECT 580.950 593.850 583.050 595.950 ;
        RECT 580.950 592.050 582.750 593.850 ;
        RECT 548.550 579.750 550.350 585.600 ;
        RECT 551.550 579.750 553.350 585.600 ;
        RECT 564.450 579.750 566.250 591.600 ;
        RECT 568.650 579.750 570.450 591.600 ;
        RECT 573.300 579.750 575.100 591.600 ;
        RECT 577.500 579.750 579.300 591.600 ;
        RECT 596.400 585.600 597.600 598.050 ;
        RECT 608.100 597.150 609.900 598.950 ;
        RECT 607.950 595.050 610.050 597.150 ;
        RECT 611.550 595.950 612.750 603.300 ;
        RECT 614.100 597.150 615.900 598.950 ;
        RECT 626.100 597.150 627.900 598.950 ;
        RECT 610.950 593.850 613.050 595.950 ;
        RECT 613.950 595.050 616.050 597.150 ;
        RECT 625.950 595.050 628.050 597.150 ;
        RECT 629.550 595.950 630.750 603.300 ;
        RECT 638.700 602.400 640.500 611.250 ;
        RECT 644.100 603.000 645.900 611.250 ;
        RECT 656.550 608.400 658.350 611.250 ;
        RECT 659.550 608.400 661.350 611.250 ;
        RECT 662.550 608.400 664.350 611.250 ;
        RECT 660.450 604.200 661.350 608.400 ;
        RECT 665.550 605.400 667.350 611.250 ;
        RECT 674.550 606.000 676.350 611.250 ;
        RECT 677.550 606.900 679.350 611.250 ;
        RECT 680.550 610.500 688.350 611.250 ;
        RECT 680.550 606.000 682.350 610.500 ;
        RECT 660.450 603.300 663.750 604.200 ;
        RECT 644.100 601.350 648.600 603.000 ;
        RECT 661.950 602.400 663.750 603.300 ;
        RECT 632.100 597.150 633.900 598.950 ;
        RECT 647.400 597.150 648.600 601.350 ;
        RECT 655.950 599.850 658.050 601.950 ;
        RECT 656.100 598.050 657.900 599.850 ;
        RECT 628.950 593.850 631.050 595.950 ;
        RECT 631.950 595.050 634.050 597.150 ;
        RECT 637.950 593.850 640.050 595.950 ;
        RECT 643.950 593.850 646.050 595.950 ;
        RECT 646.950 595.050 649.050 597.150 ;
        RECT 658.950 596.850 661.050 598.950 ;
        RECT 659.100 595.050 660.900 596.850 ;
        RECT 611.550 585.600 612.750 593.850 ;
        RECT 629.550 585.600 630.750 593.850 ;
        RECT 638.100 592.050 639.900 593.850 ;
        RECT 640.950 590.850 643.050 592.950 ;
        RECT 644.250 592.050 646.050 593.850 ;
        RECT 641.100 589.050 642.900 590.850 ;
        RECT 647.700 586.800 648.750 595.050 ;
        RECT 662.700 594.150 663.600 602.400 ;
        RECT 666.000 600.150 667.050 605.400 ;
        RECT 674.550 605.100 682.350 606.000 ;
        RECT 683.550 605.400 685.350 609.600 ;
        RECT 686.550 605.400 688.350 610.500 ;
        RECT 693.750 608.400 695.550 611.250 ;
        RECT 696.750 608.400 698.550 611.250 ;
        RECT 683.850 603.900 684.750 605.400 ;
        RECT 680.400 602.850 684.750 603.900 ;
        RECT 677.100 600.150 678.900 601.950 ;
        RECT 664.950 598.050 667.050 600.150 ;
        RECT 661.950 594.000 663.750 594.150 ;
        RECT 641.700 585.900 648.750 586.800 ;
        RECT 641.700 585.600 643.350 585.900 ;
        RECT 580.800 579.750 582.600 585.600 ;
        RECT 595.650 579.750 597.450 585.600 ;
        RECT 598.650 579.750 600.450 585.600 ;
        RECT 608.550 579.750 610.350 585.600 ;
        RECT 611.550 579.750 613.350 585.600 ;
        RECT 614.550 579.750 616.350 585.600 ;
        RECT 626.550 579.750 628.350 585.600 ;
        RECT 629.550 579.750 631.350 585.600 ;
        RECT 632.550 579.750 634.350 585.600 ;
        RECT 638.550 579.750 640.350 585.600 ;
        RECT 641.550 579.750 643.350 585.600 ;
        RECT 647.550 585.600 648.750 585.900 ;
        RECT 656.550 592.800 663.750 594.000 ;
        RECT 656.550 591.600 657.750 592.800 ;
        RECT 661.950 592.350 663.750 592.800 ;
        RECT 644.550 579.750 646.350 585.000 ;
        RECT 647.550 579.750 649.350 585.600 ;
        RECT 656.550 579.750 658.350 591.600 ;
        RECT 665.100 591.450 666.450 598.050 ;
        RECT 673.950 596.850 676.050 598.950 ;
        RECT 676.950 598.050 679.050 600.150 ;
        RECT 680.400 598.950 681.600 602.850 ;
        RECT 682.500 600.150 684.300 601.950 ;
        RECT 697.050 600.150 698.550 608.400 ;
        RECT 679.950 596.850 682.050 598.950 ;
        RECT 682.950 598.050 685.050 600.150 ;
        RECT 685.950 596.850 688.050 598.950 ;
        RECT 694.950 598.050 698.550 600.150 ;
        RECT 674.100 595.050 675.900 596.850 ;
        RECT 680.550 591.600 681.750 596.850 ;
        RECT 685.950 595.050 687.750 596.850 ;
        RECT 661.050 579.750 662.850 591.450 ;
        RECT 664.050 590.100 666.450 591.450 ;
        RECT 664.050 579.750 665.850 590.100 ;
        RECT 674.550 579.750 676.350 591.600 ;
        RECT 679.050 579.750 682.350 591.600 ;
        RECT 685.050 579.750 686.850 591.600 ;
        RECT 697.050 585.600 698.550 598.050 ;
        RECT 700.650 605.400 702.450 611.250 ;
        RECT 706.050 605.400 707.850 611.250 ;
        RECT 711.600 606.600 713.400 611.250 ;
        RECT 716.250 607.500 718.050 611.250 ;
        RECT 719.250 607.500 721.050 611.250 ;
        RECT 722.250 607.500 724.050 611.250 ;
        RECT 709.200 605.400 713.400 606.600 ;
        RECT 715.950 605.400 718.050 607.500 ;
        RECT 718.950 605.400 721.050 607.500 ;
        RECT 721.950 605.400 724.050 607.500 ;
        RECT 726.000 607.500 727.800 611.250 ;
        RECT 729.000 608.400 730.800 611.250 ;
        RECT 732.000 607.500 733.800 611.250 ;
        RECT 736.500 608.400 738.300 611.250 ;
        RECT 739.500 608.400 741.300 611.250 ;
        RECT 742.500 608.400 744.300 611.250 ;
        RECT 745.500 608.400 747.300 611.250 ;
        RECT 726.000 605.700 728.850 607.500 ;
        RECT 726.750 605.400 728.850 605.700 ;
        RECT 730.950 605.700 733.800 607.500 ;
        RECT 734.700 606.750 736.500 607.200 ;
        RECT 739.950 607.050 741.300 608.400 ;
        RECT 742.950 607.050 744.300 608.400 ;
        RECT 745.950 607.050 747.300 608.400 ;
        RECT 730.950 605.400 733.050 605.700 ;
        RECT 734.700 605.400 738.750 606.750 ;
        RECT 700.650 590.550 701.850 605.400 ;
        RECT 709.200 601.800 710.700 605.400 ;
        RECT 715.350 602.700 722.100 604.500 ;
        RECT 723.000 602.700 729.900 604.500 ;
        RECT 737.850 604.050 738.750 605.400 ;
        RECT 739.950 604.950 742.050 607.050 ;
        RECT 742.950 604.950 745.050 607.050 ;
        RECT 745.950 604.950 748.050 607.050 ;
        RECT 737.850 603.900 742.950 604.050 ;
        RECT 737.850 603.150 745.500 603.900 ;
        RECT 741.150 602.700 745.500 603.150 ;
        RECT 723.000 601.800 724.050 602.700 ;
        RECT 741.150 602.250 742.950 602.700 ;
        RECT 702.900 600.000 710.700 601.800 ;
        RECT 714.150 600.750 724.050 601.800 ;
        RECT 714.150 598.950 715.200 600.750 ;
        RECT 724.950 600.450 732.600 601.800 ;
        RECT 724.950 599.700 725.850 600.450 ;
        RECT 706.950 597.900 715.200 598.950 ;
        RECT 716.250 598.650 725.850 599.700 ;
        RECT 706.950 593.850 709.050 597.900 ;
        RECT 716.250 597.000 717.150 598.650 ;
        RECT 726.750 597.750 730.650 599.550 ;
        RECT 731.550 598.950 732.600 600.450 ;
        RECT 733.950 601.650 736.050 601.950 ;
        RECT 733.950 599.850 737.850 601.650 ;
        RECT 744.450 599.250 745.500 602.700 ;
        RECT 747.000 601.800 748.050 604.950 ;
        RECT 749.700 605.400 751.500 611.250 ;
        RECT 755.100 605.400 756.900 611.250 ;
        RECT 760.500 605.400 762.300 611.250 ;
        RECT 770.550 608.400 772.350 611.250 ;
        RECT 749.700 604.500 751.200 605.400 ;
        RECT 749.700 603.300 758.100 604.500 ;
        RECT 756.300 602.700 758.100 603.300 ;
        RECT 761.100 601.800 762.300 605.400 ;
        RECT 771.150 604.500 772.350 608.400 ;
        RECT 773.850 605.400 775.650 611.250 ;
        RECT 776.850 605.400 778.650 611.250 ;
        RECT 785.550 608.400 787.350 611.250 ;
        RECT 788.550 608.400 790.350 611.250 ;
        RECT 791.550 608.400 793.350 611.250 ;
        RECT 771.150 603.600 776.250 604.500 ;
        RECT 747.000 600.900 762.300 601.800 ;
        RECT 731.550 598.050 743.550 598.950 ;
        RECT 710.100 595.200 717.150 597.000 ;
        RECT 718.500 595.950 720.300 597.750 ;
        RECT 726.750 597.450 728.850 597.750 ;
        RECT 730.950 596.550 733.050 596.850 ;
        RECT 739.800 596.550 741.600 597.150 ;
        RECT 730.950 595.950 741.600 596.550 ;
        RECT 718.500 595.350 741.600 595.950 ;
        RECT 742.500 596.550 743.550 598.050 ;
        RECT 744.450 597.450 746.250 599.250 ;
        RECT 748.050 598.950 759.900 600.000 ;
        RECT 748.050 596.550 749.250 598.950 ;
        RECT 758.100 597.150 759.900 598.950 ;
        RECT 742.500 595.650 749.250 596.550 ;
        RECT 751.950 595.650 754.050 595.950 ;
        RECT 718.500 594.750 733.050 595.350 ;
        RECT 750.150 594.450 754.050 595.650 ;
        RECT 757.950 595.050 760.050 597.150 ;
        RECT 740.100 593.850 754.050 594.450 ;
        RECT 714.000 593.550 753.750 593.850 ;
        RECT 702.750 592.650 704.550 593.250 ;
        RECT 714.000 592.650 742.050 593.550 ;
        RECT 702.750 591.450 715.050 592.650 ;
        RECT 742.950 592.050 745.050 592.350 ;
        RECT 752.700 592.050 754.500 592.650 ;
        RECT 715.950 590.550 718.050 591.750 ;
        RECT 700.650 589.650 718.050 590.550 ;
        RECT 721.950 590.400 742.050 591.750 ;
        RECT 721.950 589.650 724.050 590.400 ;
        RECT 703.500 585.600 704.700 589.650 ;
        RECT 705.600 587.700 707.400 588.300 ;
        RECT 712.350 588.150 714.150 588.300 ;
        RECT 705.600 586.500 711.300 587.700 ;
        RECT 712.350 586.950 721.050 588.150 ;
        RECT 712.350 586.500 714.150 586.950 ;
        RECT 693.750 579.750 695.550 585.600 ;
        RECT 696.750 579.750 698.550 585.600 ;
        RECT 700.500 579.750 702.300 585.600 ;
        RECT 703.500 579.750 705.300 585.600 ;
        RECT 706.500 579.750 708.300 585.600 ;
        RECT 709.500 579.750 711.300 586.500 ;
        RECT 718.950 586.050 721.050 586.950 ;
        RECT 712.500 579.750 714.300 585.600 ;
        RECT 715.800 583.800 717.900 585.900 ;
        RECT 716.400 582.600 717.900 583.800 ;
        RECT 716.250 579.750 718.050 582.600 ;
        RECT 719.250 579.750 721.050 586.050 ;
        RECT 722.550 582.600 723.900 589.650 ;
        RECT 740.100 589.350 742.050 590.400 ;
        RECT 742.950 590.850 754.500 592.050 ;
        RECT 742.950 590.250 745.050 590.850 ;
        RECT 756.000 589.350 757.800 590.100 ;
        RECT 725.100 586.800 729.000 588.600 ;
        RECT 726.000 586.500 729.000 586.800 ;
        RECT 730.950 588.150 733.050 588.600 ;
        RECT 740.100 588.300 757.800 589.350 ;
        RECT 730.950 586.500 733.350 588.150 ;
        RECT 722.250 579.750 724.050 582.600 ;
        RECT 726.000 579.750 727.800 586.500 ;
        RECT 732.000 585.600 733.350 586.500 ;
        RECT 739.950 585.600 742.050 586.050 ;
        RECT 729.000 579.750 730.800 585.600 ;
        RECT 732.000 579.750 733.800 585.600 ;
        RECT 735.750 579.750 737.550 585.600 ;
        RECT 739.500 583.950 742.050 585.600 ;
        RECT 742.950 583.950 745.050 586.050 ;
        RECT 745.950 583.950 748.050 586.050 ;
        RECT 739.500 582.600 740.700 583.950 ;
        RECT 742.950 582.600 743.850 583.950 ;
        RECT 745.950 582.600 747.150 583.950 ;
        RECT 738.750 579.750 740.700 582.600 ;
        RECT 741.750 579.750 743.850 582.600 ;
        RECT 744.750 579.750 747.150 582.600 ;
        RECT 748.500 579.750 750.300 583.050 ;
        RECT 751.500 579.750 753.300 588.300 ;
        RECT 761.100 587.400 762.300 600.900 ;
        RECT 774.000 602.700 776.250 603.600 ;
        RECT 769.950 596.850 772.050 598.950 ;
        RECT 770.100 595.050 771.900 596.850 ;
        RECT 774.000 594.300 775.050 602.700 ;
        RECT 777.150 598.950 778.350 605.400 ;
        RECT 789.450 604.200 790.350 608.400 ;
        RECT 794.550 605.400 796.350 611.250 ;
        RECT 803.550 608.400 805.350 611.250 ;
        RECT 806.550 608.400 808.350 611.250 ;
        RECT 809.550 608.400 811.350 611.250 ;
        RECT 789.450 603.300 792.750 604.200 ;
        RECT 790.950 602.400 792.750 603.300 ;
        RECT 784.950 599.850 787.050 601.950 ;
        RECT 775.950 596.850 778.350 598.950 ;
        RECT 785.100 598.050 786.900 599.850 ;
        RECT 787.950 596.850 790.050 598.950 ;
        RECT 774.000 593.400 776.250 594.300 ;
        RECT 758.250 586.500 762.300 587.400 ;
        RECT 770.550 592.500 776.250 593.400 ;
        RECT 758.250 585.600 759.300 586.500 ;
        RECT 770.550 585.600 771.750 592.500 ;
        RECT 777.150 591.600 778.350 596.850 ;
        RECT 788.100 595.050 789.900 596.850 ;
        RECT 791.700 594.150 792.600 602.400 ;
        RECT 795.000 600.150 796.050 605.400 ;
        RECT 807.000 601.950 808.050 608.400 ;
        RECT 818.550 606.300 820.350 611.250 ;
        RECT 821.550 607.200 823.350 611.250 ;
        RECT 824.550 606.300 826.350 611.250 ;
        RECT 818.550 604.950 826.350 606.300 ;
        RECT 827.550 605.400 829.350 611.250 ;
        RECT 836.550 606.300 838.350 611.250 ;
        RECT 839.550 607.200 841.350 611.250 ;
        RECT 842.550 606.300 844.350 611.250 ;
        RECT 827.550 603.300 828.750 605.400 ;
        RECT 836.550 604.950 844.350 606.300 ;
        RECT 845.550 605.400 847.350 611.250 ;
        RECT 845.550 603.300 846.750 605.400 ;
        RECT 825.000 602.250 828.750 603.300 ;
        RECT 843.000 602.250 846.750 603.300 ;
        RECT 793.950 598.050 796.050 600.150 ;
        RECT 805.950 599.850 808.050 601.950 ;
        RECT 821.100 600.150 822.900 601.950 ;
        RECT 790.950 594.000 792.750 594.150 ;
        RECT 785.550 592.800 792.750 594.000 ;
        RECT 785.550 591.600 786.750 592.800 ;
        RECT 790.950 592.350 792.750 592.800 ;
        RECT 754.500 579.750 756.300 585.600 ;
        RECT 757.500 579.750 759.300 585.600 ;
        RECT 760.500 579.750 762.300 585.600 ;
        RECT 770.550 579.750 772.350 585.600 ;
        RECT 773.850 579.750 775.650 591.600 ;
        RECT 776.850 579.750 778.650 591.600 ;
        RECT 785.550 579.750 787.350 591.600 ;
        RECT 794.100 591.450 795.450 598.050 ;
        RECT 802.950 596.850 805.050 598.950 ;
        RECT 803.100 595.050 804.900 596.850 ;
        RECT 807.000 592.650 808.050 599.850 ;
        RECT 808.950 596.850 811.050 598.950 ;
        RECT 817.950 596.850 820.050 598.950 ;
        RECT 820.950 598.050 823.050 600.150 ;
        RECT 824.850 598.950 826.050 602.250 ;
        RECT 839.100 600.150 840.900 601.950 ;
        RECT 823.950 596.850 826.050 598.950 ;
        RECT 835.950 596.850 838.050 598.950 ;
        RECT 838.950 598.050 841.050 600.150 ;
        RECT 842.850 598.950 844.050 602.250 ;
        RECT 841.950 596.850 844.050 598.950 ;
        RECT 809.100 595.050 810.900 596.850 ;
        RECT 818.100 595.050 819.900 596.850 ;
        RECT 807.000 591.600 809.550 592.650 ;
        RECT 823.950 591.600 825.150 596.850 ;
        RECT 826.950 593.850 829.050 595.950 ;
        RECT 836.100 595.050 837.900 596.850 ;
        RECT 826.950 592.050 828.750 593.850 ;
        RECT 841.950 591.600 843.150 596.850 ;
        RECT 844.950 593.850 847.050 595.950 ;
        RECT 844.950 592.050 846.750 593.850 ;
        RECT 790.050 579.750 791.850 591.450 ;
        RECT 793.050 590.100 795.450 591.450 ;
        RECT 793.050 579.750 794.850 590.100 ;
        RECT 803.550 579.750 805.350 591.600 ;
        RECT 807.750 579.750 809.550 591.600 ;
        RECT 819.300 579.750 821.100 591.600 ;
        RECT 823.500 579.750 825.300 591.600 ;
        RECT 826.800 579.750 828.600 585.600 ;
        RECT 837.300 579.750 839.100 591.600 ;
        RECT 841.500 579.750 843.300 591.600 ;
        RECT 844.800 579.750 846.600 585.600 ;
        RECT 4.650 569.400 6.450 575.250 ;
        RECT 7.650 569.400 9.450 575.250 ;
        RECT 17.550 569.400 19.350 575.250 ;
        RECT 20.550 569.400 22.350 575.250 ;
        RECT 23.550 570.000 25.350 575.250 ;
        RECT 5.400 556.950 6.600 569.400 ;
        RECT 20.700 569.100 22.350 569.400 ;
        RECT 26.550 569.400 28.350 575.250 ;
        RECT 32.550 569.400 34.350 575.250 ;
        RECT 35.550 569.400 37.350 575.250 ;
        RECT 38.550 570.000 40.350 575.250 ;
        RECT 26.550 569.100 27.750 569.400 ;
        RECT 20.700 568.200 27.750 569.100 ;
        RECT 35.700 569.100 37.350 569.400 ;
        RECT 41.550 569.400 43.350 575.250 ;
        RECT 41.550 569.100 42.750 569.400 ;
        RECT 35.700 568.200 42.750 569.100 ;
        RECT 20.100 564.150 21.900 565.950 ;
        RECT 17.100 561.150 18.900 562.950 ;
        RECT 19.950 562.050 22.050 564.150 ;
        RECT 23.250 561.150 25.050 562.950 ;
        RECT 16.950 559.050 19.050 561.150 ;
        RECT 22.950 559.050 25.050 561.150 ;
        RECT 26.700 559.950 27.750 568.200 ;
        RECT 35.100 564.150 36.900 565.950 ;
        RECT 32.100 561.150 33.900 562.950 ;
        RECT 34.950 562.050 37.050 564.150 ;
        RECT 38.250 561.150 40.050 562.950 ;
        RECT 25.950 557.850 28.050 559.950 ;
        RECT 31.950 559.050 34.050 561.150 ;
        RECT 37.950 559.050 40.050 561.150 ;
        RECT 41.700 559.950 42.750 568.200 ;
        RECT 47.550 564.300 49.350 575.250 ;
        RECT 50.550 565.200 52.350 575.250 ;
        RECT 53.550 564.300 55.350 575.250 ;
        RECT 47.550 563.400 55.350 564.300 ;
        RECT 56.550 563.400 58.350 575.250 ;
        RECT 72.150 564.900 73.950 575.250 ;
        RECT 71.550 563.550 73.950 564.900 ;
        RECT 75.150 563.550 76.950 575.250 ;
        RECT 40.950 557.850 43.050 559.950 ;
        RECT 56.700 558.150 57.900 563.400 ;
        RECT 4.950 554.850 7.050 556.950 ;
        RECT 8.100 555.150 9.900 556.950 ;
        RECT 5.400 546.600 6.600 554.850 ;
        RECT 7.950 553.050 10.050 555.150 ;
        RECT 26.400 553.650 27.600 557.850 ;
        RECT 41.400 553.650 42.600 557.850 ;
        RECT 46.950 554.850 49.050 556.950 ;
        RECT 50.100 555.150 51.900 556.950 ;
        RECT 4.650 543.750 6.450 546.600 ;
        RECT 7.650 543.750 9.450 546.600 ;
        RECT 17.700 543.750 19.500 552.600 ;
        RECT 23.100 552.000 27.600 553.650 ;
        RECT 23.100 543.750 24.900 552.000 ;
        RECT 32.700 543.750 34.500 552.600 ;
        RECT 38.100 552.000 42.600 553.650 ;
        RECT 47.100 553.050 48.900 554.850 ;
        RECT 49.950 553.050 52.050 555.150 ;
        RECT 52.950 554.850 55.050 556.950 ;
        RECT 55.950 556.050 58.050 558.150 ;
        RECT 71.550 556.950 72.900 563.550 ;
        RECT 79.650 563.400 81.450 575.250 ;
        RECT 89.550 569.400 91.350 575.250 ;
        RECT 92.550 569.400 94.350 575.250 ;
        RECT 95.550 569.400 97.350 575.250 ;
        RECT 74.250 562.200 76.050 562.650 ;
        RECT 80.250 562.200 81.450 563.400 ;
        RECT 74.250 561.000 81.450 562.200 ;
        RECT 92.550 561.150 93.750 569.400 ;
        RECT 101.550 563.400 103.350 575.250 ;
        RECT 105.750 563.400 107.550 575.250 ;
        RECT 121.050 563.400 122.850 575.250 ;
        RECT 124.050 563.400 125.850 575.250 ;
        RECT 127.650 569.400 129.450 575.250 ;
        RECT 130.650 569.400 132.450 575.250 ;
        RECT 105.000 562.350 107.550 563.400 ;
        RECT 74.250 560.850 76.050 561.000 ;
        RECT 53.100 553.050 54.900 554.850 ;
        RECT 38.100 543.750 39.900 552.000 ;
        RECT 56.700 549.600 57.900 556.050 ;
        RECT 70.950 554.850 73.050 556.950 ;
        RECT 70.950 549.600 72.000 554.850 ;
        RECT 74.400 552.600 75.300 560.850 ;
        RECT 77.100 558.150 78.900 559.950 ;
        RECT 76.950 556.050 79.050 558.150 ;
        RECT 88.950 557.850 91.050 559.950 ;
        RECT 91.950 559.050 94.050 561.150 ;
        RECT 80.100 555.150 81.900 556.950 ;
        RECT 89.100 556.050 90.900 557.850 ;
        RECT 79.950 553.050 82.050 555.150 ;
        RECT 74.250 551.700 76.050 552.600 ;
        RECT 92.550 551.700 93.750 559.050 ;
        RECT 94.950 557.850 97.050 559.950 ;
        RECT 101.100 558.150 102.900 559.950 ;
        RECT 95.100 556.050 96.900 557.850 ;
        RECT 100.950 556.050 103.050 558.150 ;
        RECT 105.000 555.150 106.050 562.350 ;
        RECT 107.100 558.150 108.900 559.950 ;
        RECT 121.650 558.150 122.850 563.400 ;
        RECT 106.950 556.050 109.050 558.150 ;
        RECT 121.650 556.050 124.050 558.150 ;
        RECT 124.950 557.850 127.050 559.950 ;
        RECT 125.100 556.050 126.900 557.850 ;
        RECT 103.950 553.050 106.050 555.150 ;
        RECT 74.250 550.800 77.550 551.700 ;
        RECT 92.550 550.800 96.150 551.700 ;
        RECT 48.000 543.750 49.800 549.600 ;
        RECT 52.200 547.950 57.900 549.600 ;
        RECT 52.200 543.750 54.000 547.950 ;
        RECT 55.500 543.750 57.300 546.600 ;
        RECT 70.650 543.750 72.450 549.600 ;
        RECT 76.650 546.600 77.550 550.800 ;
        RECT 73.650 543.750 75.450 546.600 ;
        RECT 76.650 543.750 78.450 546.600 ;
        RECT 79.650 543.750 81.450 546.600 ;
        RECT 89.850 543.750 91.650 549.600 ;
        RECT 94.350 543.750 96.150 550.800 ;
        RECT 105.000 546.600 106.050 553.050 ;
        RECT 121.650 549.600 122.850 556.050 ;
        RECT 128.100 552.300 129.300 569.400 ;
        RECT 136.650 563.400 138.450 575.250 ;
        RECT 139.650 562.500 141.450 575.250 ;
        RECT 142.650 563.400 144.450 575.250 ;
        RECT 145.650 562.500 147.450 575.250 ;
        RECT 148.650 563.400 150.450 575.250 ;
        RECT 151.650 562.500 153.450 575.250 ;
        RECT 154.650 563.400 156.450 575.250 ;
        RECT 157.650 562.500 159.450 575.250 ;
        RECT 160.650 563.400 162.450 575.250 ;
        RECT 171.450 563.400 173.250 575.250 ;
        RECT 175.650 563.400 177.450 575.250 ;
        RECT 183.450 563.400 185.250 575.250 ;
        RECT 187.650 563.400 189.450 575.250 ;
        RECT 193.650 569.400 195.450 575.250 ;
        RECT 196.650 569.400 198.450 575.250 ;
        RECT 199.650 569.400 201.450 575.250 ;
        RECT 203.550 569.400 205.350 575.250 ;
        RECT 206.550 569.400 208.350 575.250 ;
        RECT 209.550 569.400 211.350 575.250 ;
        RECT 221.550 569.400 223.350 575.250 ;
        RECT 138.750 561.300 141.450 562.500 ;
        RECT 143.700 561.300 147.450 562.500 ;
        RECT 149.700 561.300 153.450 562.500 ;
        RECT 155.550 561.300 159.450 562.500 ;
        RECT 171.450 562.350 174.000 563.400 ;
        RECT 183.450 562.350 186.000 563.400 ;
        RECT 131.100 558.150 132.900 559.950 ;
        RECT 130.950 556.050 133.050 558.150 ;
        RECT 138.750 556.950 139.800 561.300 ;
        RECT 136.950 554.850 139.800 556.950 ;
        RECT 124.950 551.100 132.450 552.300 ;
        RECT 124.950 550.500 126.750 551.100 ;
        RECT 121.650 548.100 124.950 549.600 ;
        RECT 101.550 543.750 103.350 546.600 ;
        RECT 104.550 543.750 106.350 546.600 ;
        RECT 107.550 543.750 109.350 546.600 ;
        RECT 123.150 543.750 124.950 548.100 ;
        RECT 126.150 543.750 127.950 549.600 ;
        RECT 130.650 543.750 132.450 551.100 ;
        RECT 138.750 551.700 139.800 554.850 ;
        RECT 143.700 554.400 144.900 561.300 ;
        RECT 149.700 554.400 150.900 561.300 ;
        RECT 155.550 554.400 156.750 561.300 ;
        RECT 170.100 558.150 171.900 559.950 ;
        RECT 157.950 554.850 160.050 556.950 ;
        RECT 169.950 556.050 172.050 558.150 ;
        RECT 172.950 555.150 174.000 562.350 ;
        RECT 176.100 558.150 177.900 559.950 ;
        RECT 182.100 558.150 183.900 559.950 ;
        RECT 175.950 556.050 178.050 558.150 ;
        RECT 181.950 556.050 184.050 558.150 ;
        RECT 184.950 555.150 186.000 562.350 ;
        RECT 197.250 561.150 198.450 569.400 ;
        RECT 206.550 561.150 207.750 569.400 ;
        RECT 221.550 562.500 222.750 569.400 ;
        RECT 224.850 563.400 226.650 575.250 ;
        RECT 227.850 563.400 229.650 575.250 ;
        RECT 239.550 569.400 241.350 575.250 ;
        RECT 242.550 569.400 244.350 575.250 ;
        RECT 245.550 569.400 247.350 575.250 ;
        RECT 256.650 569.400 258.450 575.250 ;
        RECT 259.650 569.400 261.450 575.250 ;
        RECT 221.550 561.600 227.250 562.500 ;
        RECT 188.100 558.150 189.900 559.950 ;
        RECT 187.950 556.050 190.050 558.150 ;
        RECT 193.950 557.850 196.050 559.950 ;
        RECT 196.950 559.050 199.050 561.150 ;
        RECT 194.100 556.050 195.900 557.850 ;
        RECT 140.700 552.600 144.900 554.400 ;
        RECT 146.700 552.600 150.900 554.400 ;
        RECT 152.700 552.600 156.750 554.400 ;
        RECT 158.100 553.050 159.900 554.850 ;
        RECT 172.950 553.050 175.050 555.150 ;
        RECT 184.950 553.050 187.050 555.150 ;
        RECT 143.700 551.700 144.900 552.600 ;
        RECT 149.700 551.700 150.900 552.600 ;
        RECT 155.550 551.700 156.750 552.600 ;
        RECT 138.750 550.650 141.600 551.700 ;
        RECT 138.900 550.500 141.600 550.650 ;
        RECT 143.700 550.500 147.600 551.700 ;
        RECT 149.700 550.500 153.450 551.700 ;
        RECT 155.550 550.500 159.600 551.700 ;
        RECT 139.800 549.600 141.600 550.500 ;
        RECT 145.800 549.600 147.600 550.500 ;
        RECT 136.650 543.750 138.450 549.600 ;
        RECT 139.650 543.750 141.450 549.600 ;
        RECT 142.650 543.750 144.450 549.600 ;
        RECT 145.650 543.750 147.450 549.600 ;
        RECT 148.650 543.750 150.450 549.600 ;
        RECT 151.650 543.750 153.450 550.500 ;
        RECT 157.800 549.600 159.600 550.500 ;
        RECT 154.650 543.750 156.450 549.600 ;
        RECT 157.650 543.750 159.450 549.600 ;
        RECT 160.650 543.750 162.450 549.600 ;
        RECT 172.950 546.600 174.000 553.050 ;
        RECT 184.950 546.600 186.000 553.050 ;
        RECT 197.250 551.700 198.450 559.050 ;
        RECT 199.950 557.850 202.050 559.950 ;
        RECT 202.950 557.850 205.050 559.950 ;
        RECT 205.950 559.050 208.050 561.150 ;
        RECT 225.000 560.700 227.250 561.600 ;
        RECT 200.100 556.050 201.900 557.850 ;
        RECT 203.100 556.050 204.900 557.850 ;
        RECT 194.850 550.800 198.450 551.700 ;
        RECT 206.550 551.700 207.750 559.050 ;
        RECT 208.950 557.850 211.050 559.950 ;
        RECT 221.100 558.150 222.900 559.950 ;
        RECT 209.100 556.050 210.900 557.850 ;
        RECT 220.950 556.050 223.050 558.150 ;
        RECT 225.000 552.300 226.050 560.700 ;
        RECT 228.150 558.150 229.350 563.400 ;
        RECT 242.550 561.150 243.750 569.400 ;
        RECT 226.950 556.050 229.350 558.150 ;
        RECT 238.950 557.850 241.050 559.950 ;
        RECT 241.950 559.050 244.050 561.150 ;
        RECT 239.100 556.050 240.900 557.850 ;
        RECT 206.550 550.800 210.150 551.700 ;
        RECT 225.000 551.400 227.250 552.300 ;
        RECT 169.650 543.750 171.450 546.600 ;
        RECT 172.650 543.750 174.450 546.600 ;
        RECT 175.650 543.750 177.450 546.600 ;
        RECT 181.650 543.750 183.450 546.600 ;
        RECT 184.650 543.750 186.450 546.600 ;
        RECT 187.650 543.750 189.450 546.600 ;
        RECT 194.850 543.750 196.650 550.800 ;
        RECT 199.350 543.750 201.150 549.600 ;
        RECT 203.850 543.750 205.650 549.600 ;
        RECT 208.350 543.750 210.150 550.800 ;
        RECT 222.150 550.500 227.250 551.400 ;
        RECT 222.150 546.600 223.350 550.500 ;
        RECT 228.150 549.600 229.350 556.050 ;
        RECT 242.550 551.700 243.750 559.050 ;
        RECT 244.950 557.850 247.050 559.950 ;
        RECT 245.100 556.050 246.900 557.850 ;
        RECT 257.400 556.950 258.600 569.400 ;
        RECT 264.300 563.400 266.100 575.250 ;
        RECT 268.500 563.400 270.300 575.250 ;
        RECT 271.800 569.400 273.600 575.250 ;
        RECT 278.550 563.400 280.350 575.250 ;
        RECT 282.750 563.400 284.550 575.250 ;
        RECT 296.550 569.400 298.350 575.250 ;
        RECT 299.550 569.400 301.350 575.250 ;
        RECT 302.550 570.000 304.350 575.250 ;
        RECT 299.700 569.100 301.350 569.400 ;
        RECT 305.550 569.400 307.350 575.250 ;
        RECT 305.550 569.100 306.750 569.400 ;
        RECT 299.700 568.200 306.750 569.100 ;
        RECT 299.100 564.150 300.900 565.950 ;
        RECT 263.100 558.150 264.900 559.950 ;
        RECT 268.950 558.150 270.150 563.400 ;
        RECT 271.950 561.150 273.750 562.950 ;
        RECT 282.000 562.350 284.550 563.400 ;
        RECT 271.950 559.050 274.050 561.150 ;
        RECT 278.100 558.150 279.900 559.950 ;
        RECT 256.950 554.850 259.050 556.950 ;
        RECT 260.100 555.150 261.900 556.950 ;
        RECT 262.950 556.050 265.050 558.150 ;
        RECT 242.550 550.800 246.150 551.700 ;
        RECT 221.550 543.750 223.350 546.600 ;
        RECT 224.850 543.750 226.650 549.600 ;
        RECT 227.850 543.750 229.650 549.600 ;
        RECT 239.850 543.750 241.650 549.600 ;
        RECT 244.350 543.750 246.150 550.800 ;
        RECT 257.400 546.600 258.600 554.850 ;
        RECT 259.950 553.050 262.050 555.150 ;
        RECT 265.950 554.850 268.050 556.950 ;
        RECT 268.950 556.050 271.050 558.150 ;
        RECT 277.950 556.050 280.050 558.150 ;
        RECT 266.100 553.050 267.900 554.850 ;
        RECT 269.850 552.750 271.050 556.050 ;
        RECT 282.000 555.150 283.050 562.350 ;
        RECT 296.100 561.150 297.900 562.950 ;
        RECT 298.950 562.050 301.050 564.150 ;
        RECT 302.250 561.150 304.050 562.950 ;
        RECT 284.100 558.150 285.900 559.950 ;
        RECT 295.950 559.050 298.050 561.150 ;
        RECT 301.950 559.050 304.050 561.150 ;
        RECT 305.700 559.950 306.750 568.200 ;
        RECT 315.450 563.400 317.250 575.250 ;
        RECT 319.650 563.400 321.450 575.250 ;
        RECT 325.650 569.400 327.450 575.250 ;
        RECT 328.650 570.000 330.450 575.250 ;
        RECT 326.250 569.100 327.450 569.400 ;
        RECT 331.650 569.400 333.450 575.250 ;
        RECT 334.650 569.400 336.450 575.250 ;
        RECT 331.650 569.100 333.300 569.400 ;
        RECT 326.250 568.200 333.300 569.100 ;
        RECT 315.450 562.350 318.000 563.400 ;
        RECT 283.950 556.050 286.050 558.150 ;
        RECT 304.950 557.850 307.050 559.950 ;
        RECT 314.100 558.150 315.900 559.950 ;
        RECT 280.950 553.050 283.050 555.150 ;
        RECT 305.400 553.650 306.600 557.850 ;
        RECT 313.950 556.050 316.050 558.150 ;
        RECT 270.000 551.700 273.750 552.750 ;
        RECT 263.550 548.700 271.350 550.050 ;
        RECT 256.650 543.750 258.450 546.600 ;
        RECT 259.650 543.750 261.450 546.600 ;
        RECT 263.550 543.750 265.350 548.700 ;
        RECT 266.550 543.750 268.350 547.800 ;
        RECT 269.550 543.750 271.350 548.700 ;
        RECT 272.550 549.600 273.750 551.700 ;
        RECT 272.550 543.750 274.350 549.600 ;
        RECT 282.000 546.600 283.050 553.050 ;
        RECT 278.550 543.750 280.350 546.600 ;
        RECT 281.550 543.750 283.350 546.600 ;
        RECT 284.550 543.750 286.350 546.600 ;
        RECT 296.700 543.750 298.500 552.600 ;
        RECT 302.100 552.000 306.600 553.650 ;
        RECT 316.950 555.150 318.000 562.350 ;
        RECT 326.250 559.950 327.300 568.200 ;
        RECT 332.100 564.150 333.900 565.950 ;
        RECT 328.950 561.150 330.750 562.950 ;
        RECT 331.950 562.050 334.050 564.150 ;
        RECT 344.550 563.400 346.350 575.250 ;
        RECT 348.750 563.400 350.550 575.250 ;
        RECT 364.650 569.400 366.450 575.250 ;
        RECT 367.650 569.400 369.450 575.250 ;
        RECT 374.550 569.400 376.350 575.250 ;
        RECT 377.550 569.400 379.350 575.250 ;
        RECT 380.550 570.000 382.350 575.250 ;
        RECT 335.100 561.150 336.900 562.950 ;
        RECT 348.000 562.350 350.550 563.400 ;
        RECT 320.100 558.150 321.900 559.950 ;
        RECT 319.950 556.050 322.050 558.150 ;
        RECT 325.950 557.850 328.050 559.950 ;
        RECT 328.950 559.050 331.050 561.150 ;
        RECT 334.950 559.050 337.050 561.150 ;
        RECT 340.950 558.450 343.050 559.050 ;
        RECT 316.950 553.050 319.050 555.150 ;
        RECT 326.400 553.650 327.600 557.850 ;
        RECT 338.550 557.550 343.050 558.450 ;
        RECT 344.100 558.150 345.900 559.950 ;
        RECT 334.950 555.450 337.050 556.050 ;
        RECT 338.550 555.450 339.450 557.550 ;
        RECT 340.950 556.950 343.050 557.550 ;
        RECT 343.950 556.050 346.050 558.150 ;
        RECT 334.950 554.550 339.450 555.450 ;
        RECT 348.000 555.150 349.050 562.350 ;
        RECT 350.100 558.150 351.900 559.950 ;
        RECT 349.950 556.050 352.050 558.150 ;
        RECT 365.400 556.950 366.600 569.400 ;
        RECT 377.700 569.100 379.350 569.400 ;
        RECT 383.550 569.400 385.350 575.250 ;
        RECT 390.750 569.400 392.550 575.250 ;
        RECT 393.750 569.400 395.550 575.250 ;
        RECT 397.500 569.400 399.300 575.250 ;
        RECT 400.500 569.400 402.300 575.250 ;
        RECT 403.500 569.400 405.300 575.250 ;
        RECT 383.550 569.100 384.750 569.400 ;
        RECT 377.700 568.200 384.750 569.100 ;
        RECT 377.100 564.150 378.900 565.950 ;
        RECT 374.100 561.150 375.900 562.950 ;
        RECT 376.950 562.050 379.050 564.150 ;
        RECT 380.250 561.150 382.050 562.950 ;
        RECT 373.950 559.050 376.050 561.150 ;
        RECT 379.950 559.050 382.050 561.150 ;
        RECT 383.700 559.950 384.750 568.200 ;
        RECT 382.950 557.850 385.050 559.950 ;
        RECT 334.950 553.950 337.050 554.550 ;
        RECT 302.100 543.750 303.900 552.000 ;
        RECT 316.950 546.600 318.000 553.050 ;
        RECT 326.400 552.000 330.900 553.650 ;
        RECT 346.950 553.050 349.050 555.150 ;
        RECT 364.950 554.850 367.050 556.950 ;
        RECT 368.100 555.150 369.900 556.950 ;
        RECT 313.650 543.750 315.450 546.600 ;
        RECT 316.650 543.750 318.450 546.600 ;
        RECT 319.650 543.750 321.450 546.600 ;
        RECT 329.100 543.750 330.900 552.000 ;
        RECT 334.500 543.750 336.300 552.600 ;
        RECT 348.000 546.600 349.050 553.050 ;
        RECT 349.950 552.450 352.050 553.050 ;
        RECT 361.950 552.450 364.050 553.050 ;
        RECT 349.950 551.550 364.050 552.450 ;
        RECT 349.950 550.950 352.050 551.550 ;
        RECT 361.950 550.950 364.050 551.550 ;
        RECT 365.400 546.600 366.600 554.850 ;
        RECT 367.950 553.050 370.050 555.150 ;
        RECT 383.400 553.650 384.600 557.850 ;
        RECT 394.050 556.950 395.550 569.400 ;
        RECT 400.500 565.350 401.700 569.400 ;
        RECT 406.500 568.500 408.300 575.250 ;
        RECT 409.500 569.400 411.300 575.250 ;
        RECT 413.250 572.400 415.050 575.250 ;
        RECT 413.400 571.200 414.900 572.400 ;
        RECT 412.800 569.100 414.900 571.200 ;
        RECT 416.250 568.950 418.050 575.250 ;
        RECT 419.250 572.400 421.050 575.250 ;
        RECT 402.600 567.300 408.300 568.500 ;
        RECT 409.350 568.050 411.150 568.500 ;
        RECT 415.950 568.050 418.050 568.950 ;
        RECT 402.600 566.700 404.400 567.300 ;
        RECT 409.350 566.850 418.050 568.050 ;
        RECT 409.350 566.700 411.150 566.850 ;
        RECT 419.550 565.350 420.900 572.400 ;
        RECT 423.000 568.500 424.800 575.250 ;
        RECT 426.000 569.400 427.800 575.250 ;
        RECT 429.000 569.400 430.800 575.250 ;
        RECT 432.750 569.400 434.550 575.250 ;
        RECT 435.750 572.400 437.700 575.250 ;
        RECT 438.750 572.400 440.850 575.250 ;
        RECT 441.750 572.400 444.150 575.250 ;
        RECT 436.500 571.050 437.700 572.400 ;
        RECT 439.950 571.050 440.850 572.400 ;
        RECT 442.950 571.050 444.150 572.400 ;
        RECT 445.500 571.950 447.300 575.250 ;
        RECT 436.500 569.400 439.050 571.050 ;
        RECT 429.000 568.500 430.350 569.400 ;
        RECT 436.950 568.950 439.050 569.400 ;
        RECT 439.950 568.950 442.050 571.050 ;
        RECT 442.950 568.950 445.050 571.050 ;
        RECT 423.000 568.200 426.000 568.500 ;
        RECT 422.100 566.400 426.000 568.200 ;
        RECT 427.950 566.850 430.350 568.500 ;
        RECT 427.950 566.400 430.050 566.850 ;
        RECT 448.500 566.700 450.300 575.250 ;
        RECT 451.500 569.400 453.300 575.250 ;
        RECT 454.500 569.400 456.300 575.250 ;
        RECT 457.500 569.400 459.300 575.250 ;
        RECT 461.550 569.400 463.350 575.250 ;
        RECT 464.550 569.400 466.350 575.250 ;
        RECT 476.550 569.400 478.350 575.250 ;
        RECT 479.550 569.400 481.350 575.250 ;
        RECT 482.550 569.400 484.350 575.250 ;
        RECT 493.650 574.500 501.450 575.250 ;
        RECT 455.250 568.500 456.300 569.400 ;
        RECT 455.250 567.600 459.300 568.500 ;
        RECT 437.100 565.650 454.800 566.700 ;
        RECT 391.950 554.850 395.550 556.950 ;
        RECT 344.550 543.750 346.350 546.600 ;
        RECT 347.550 543.750 349.350 546.600 ;
        RECT 350.550 543.750 352.350 546.600 ;
        RECT 364.650 543.750 366.450 546.600 ;
        RECT 367.650 543.750 369.450 546.600 ;
        RECT 374.700 543.750 376.500 552.600 ;
        RECT 380.100 552.000 384.600 553.650 ;
        RECT 380.100 543.750 381.900 552.000 ;
        RECT 394.050 546.600 395.550 554.850 ;
        RECT 390.750 543.750 392.550 546.600 ;
        RECT 393.750 543.750 395.550 546.600 ;
        RECT 397.650 564.450 415.050 565.350 ;
        RECT 397.650 549.600 398.850 564.450 ;
        RECT 399.750 562.350 412.050 563.550 ;
        RECT 412.950 563.250 415.050 564.450 ;
        RECT 418.950 564.600 421.050 565.350 ;
        RECT 437.100 564.600 439.050 565.650 ;
        RECT 453.000 564.900 454.800 565.650 ;
        RECT 418.950 563.250 439.050 564.600 ;
        RECT 439.950 564.150 442.050 564.750 ;
        RECT 439.950 562.950 451.500 564.150 ;
        RECT 439.950 562.650 442.050 562.950 ;
        RECT 449.700 562.350 451.500 562.950 ;
        RECT 399.750 561.750 401.550 562.350 ;
        RECT 411.000 561.450 439.050 562.350 ;
        RECT 411.000 561.150 450.750 561.450 ;
        RECT 403.950 557.100 406.050 561.150 ;
        RECT 437.100 560.550 451.050 561.150 ;
        RECT 407.100 558.000 414.150 559.800 ;
        RECT 403.950 556.050 412.200 557.100 ;
        RECT 399.900 553.200 407.700 555.000 ;
        RECT 411.150 554.250 412.200 556.050 ;
        RECT 413.250 556.350 414.150 558.000 ;
        RECT 415.500 559.650 430.050 560.250 ;
        RECT 415.500 559.050 438.600 559.650 ;
        RECT 447.150 559.350 451.050 560.550 ;
        RECT 415.500 557.250 417.300 559.050 ;
        RECT 427.950 558.450 438.600 559.050 ;
        RECT 427.950 558.150 430.050 558.450 ;
        RECT 436.800 557.850 438.600 558.450 ;
        RECT 439.500 558.450 446.250 559.350 ;
        RECT 448.950 559.050 451.050 559.350 ;
        RECT 423.750 557.250 425.850 557.550 ;
        RECT 413.250 555.300 422.850 556.350 ;
        RECT 423.750 555.450 427.650 557.250 ;
        RECT 439.500 556.950 440.550 558.450 ;
        RECT 428.550 556.050 440.550 556.950 ;
        RECT 421.950 554.550 422.850 555.300 ;
        RECT 428.550 554.550 429.600 556.050 ;
        RECT 441.450 555.750 443.250 557.550 ;
        RECT 445.050 556.050 446.250 558.450 ;
        RECT 454.950 557.850 457.050 559.950 ;
        RECT 455.100 556.050 456.900 557.850 ;
        RECT 411.150 553.200 421.050 554.250 ;
        RECT 421.950 553.200 429.600 554.550 ;
        RECT 430.950 553.350 434.850 555.150 ;
        RECT 406.200 549.600 407.700 553.200 ;
        RECT 420.000 552.300 421.050 553.200 ;
        RECT 430.950 553.050 433.050 553.350 ;
        RECT 438.150 552.300 439.950 552.750 ;
        RECT 441.450 552.300 442.500 555.750 ;
        RECT 445.050 555.000 456.900 556.050 ;
        RECT 458.100 554.100 459.300 567.600 ;
        RECT 464.400 556.950 465.600 569.400 ;
        RECT 479.550 561.150 480.750 569.400 ;
        RECT 493.650 563.400 495.450 574.500 ;
        RECT 496.650 563.400 498.450 573.600 ;
        RECT 499.650 564.600 501.450 574.500 ;
        RECT 502.650 565.500 504.450 575.250 ;
        RECT 505.650 564.600 507.450 575.250 ;
        RECT 499.650 563.700 507.450 564.600 ;
        RECT 516.300 563.400 518.100 575.250 ;
        RECT 520.500 563.400 522.300 575.250 ;
        RECT 523.800 569.400 525.600 575.250 ;
        RECT 534.450 563.400 536.250 575.250 ;
        RECT 538.650 563.400 540.450 575.250 ;
        RECT 544.650 569.400 546.450 575.250 ;
        RECT 547.650 569.400 549.450 575.250 ;
        RECT 557.550 569.400 559.350 575.250 ;
        RECT 560.550 569.400 562.350 575.250 ;
        RECT 563.550 570.000 565.350 575.250 ;
        RECT 496.800 562.500 498.600 563.400 ;
        RECT 496.800 561.600 500.850 562.500 ;
        RECT 475.950 557.850 478.050 559.950 ;
        RECT 478.950 559.050 481.050 561.150 ;
        RECT 461.100 555.150 462.900 556.950 ;
        RECT 412.350 550.500 419.100 552.300 ;
        RECT 420.000 550.500 426.900 552.300 ;
        RECT 438.150 551.850 442.500 552.300 ;
        RECT 434.850 551.100 442.500 551.850 ;
        RECT 444.000 553.200 459.300 554.100 ;
        RECT 434.850 550.950 439.950 551.100 ;
        RECT 434.850 549.600 435.750 550.950 ;
        RECT 444.000 550.050 445.050 553.200 ;
        RECT 453.300 551.700 455.100 552.300 ;
        RECT 397.650 543.750 399.450 549.600 ;
        RECT 403.050 543.750 404.850 549.600 ;
        RECT 406.200 548.400 410.400 549.600 ;
        RECT 408.600 543.750 410.400 548.400 ;
        RECT 412.950 547.500 415.050 549.600 ;
        RECT 415.950 547.500 418.050 549.600 ;
        RECT 418.950 547.500 421.050 549.600 ;
        RECT 423.750 549.300 425.850 549.600 ;
        RECT 413.250 543.750 415.050 547.500 ;
        RECT 416.250 543.750 418.050 547.500 ;
        RECT 419.250 543.750 421.050 547.500 ;
        RECT 423.000 547.500 425.850 549.300 ;
        RECT 427.950 549.300 430.050 549.600 ;
        RECT 427.950 547.500 430.800 549.300 ;
        RECT 431.700 548.250 435.750 549.600 ;
        RECT 431.700 547.800 433.500 548.250 ;
        RECT 436.950 547.950 439.050 550.050 ;
        RECT 439.950 547.950 442.050 550.050 ;
        RECT 442.950 547.950 445.050 550.050 ;
        RECT 446.700 550.500 455.100 551.700 ;
        RECT 446.700 549.600 448.200 550.500 ;
        RECT 458.100 549.600 459.300 553.200 ;
        RECT 460.950 553.050 463.050 555.150 ;
        RECT 463.950 554.850 466.050 556.950 ;
        RECT 476.100 556.050 477.900 557.850 ;
        RECT 423.000 543.750 424.800 547.500 ;
        RECT 426.000 543.750 427.800 546.600 ;
        RECT 429.000 543.750 430.800 547.500 ;
        RECT 436.950 546.600 438.300 547.950 ;
        RECT 439.950 546.600 441.300 547.950 ;
        RECT 442.950 546.600 444.300 547.950 ;
        RECT 433.500 543.750 435.300 546.600 ;
        RECT 436.500 543.750 438.300 546.600 ;
        RECT 439.500 543.750 441.300 546.600 ;
        RECT 442.500 543.750 444.300 546.600 ;
        RECT 446.700 543.750 448.500 549.600 ;
        RECT 452.100 543.750 453.900 549.600 ;
        RECT 457.500 543.750 459.300 549.600 ;
        RECT 464.400 546.600 465.600 554.850 ;
        RECT 479.550 551.700 480.750 559.050 ;
        RECT 481.950 557.850 484.050 559.950 ;
        RECT 494.100 558.150 495.900 559.950 ;
        RECT 499.950 558.150 500.850 561.600 ;
        RECT 505.950 558.150 507.750 559.950 ;
        RECT 515.100 558.150 516.900 559.950 ;
        RECT 520.950 558.150 522.150 563.400 ;
        RECT 523.950 561.150 525.750 562.950 ;
        RECT 534.450 562.350 537.000 563.400 ;
        RECT 523.950 559.050 526.050 561.150 ;
        RECT 533.100 558.150 534.900 559.950 ;
        RECT 482.100 556.050 483.900 557.850 ;
        RECT 493.950 556.050 496.050 558.150 ;
        RECT 496.950 554.850 499.050 556.950 ;
        RECT 499.950 556.050 502.050 558.150 ;
        RECT 497.250 553.050 499.050 554.850 ;
        RECT 479.550 550.800 483.150 551.700 ;
        RECT 461.550 543.750 463.350 546.600 ;
        RECT 464.550 543.750 466.350 546.600 ;
        RECT 476.850 543.750 478.650 549.600 ;
        RECT 481.350 543.750 483.150 550.800 ;
        RECT 501.000 549.600 502.050 556.050 ;
        RECT 502.950 554.850 505.050 556.950 ;
        RECT 505.950 556.050 508.050 558.150 ;
        RECT 514.950 556.050 517.050 558.150 ;
        RECT 517.950 554.850 520.050 556.950 ;
        RECT 520.950 556.050 523.050 558.150 ;
        RECT 532.950 556.050 535.050 558.150 ;
        RECT 502.950 553.050 504.750 554.850 ;
        RECT 518.100 553.050 519.900 554.850 ;
        RECT 521.850 552.750 523.050 556.050 ;
        RECT 535.950 555.150 537.000 562.350 ;
        RECT 539.100 558.150 540.900 559.950 ;
        RECT 538.950 556.050 541.050 558.150 ;
        RECT 545.400 556.950 546.600 569.400 ;
        RECT 560.700 569.100 562.350 569.400 ;
        RECT 566.550 569.400 568.350 575.250 ;
        RECT 580.650 569.400 582.450 575.250 ;
        RECT 583.650 569.400 585.450 575.250 ;
        RECT 593.400 569.400 595.200 575.250 ;
        RECT 566.550 569.100 567.750 569.400 ;
        RECT 560.700 568.200 567.750 569.100 ;
        RECT 560.100 564.150 561.900 565.950 ;
        RECT 557.100 561.150 558.900 562.950 ;
        RECT 559.950 562.050 562.050 564.150 ;
        RECT 563.250 561.150 565.050 562.950 ;
        RECT 556.950 559.050 559.050 561.150 ;
        RECT 562.950 559.050 565.050 561.150 ;
        RECT 566.700 559.950 567.750 568.200 ;
        RECT 565.950 557.850 568.050 559.950 ;
        RECT 535.950 553.050 538.050 555.150 ;
        RECT 544.950 554.850 547.050 556.950 ;
        RECT 548.100 555.150 549.900 556.950 ;
        RECT 522.000 551.700 525.750 552.750 ;
        RECT 496.800 543.750 498.600 549.600 ;
        RECT 501.000 543.750 502.800 549.600 ;
        RECT 505.200 543.750 507.000 549.600 ;
        RECT 515.550 548.700 523.350 550.050 ;
        RECT 515.550 543.750 517.350 548.700 ;
        RECT 518.550 543.750 520.350 547.800 ;
        RECT 521.550 543.750 523.350 548.700 ;
        RECT 524.550 549.600 525.750 551.700 ;
        RECT 524.550 543.750 526.350 549.600 ;
        RECT 535.950 546.600 537.000 553.050 ;
        RECT 545.400 546.600 546.600 554.850 ;
        RECT 547.950 553.050 550.050 555.150 ;
        RECT 566.400 553.650 567.600 557.850 ;
        RECT 581.400 556.950 582.600 569.400 ;
        RECT 596.700 563.400 598.500 575.250 ;
        RECT 600.900 563.400 602.700 575.250 ;
        RECT 611.550 563.400 613.350 575.250 ;
        RECT 616.050 563.550 617.850 575.250 ;
        RECT 619.050 564.900 620.850 575.250 ;
        RECT 628.650 569.400 630.450 575.250 ;
        RECT 631.650 569.400 633.450 575.250 ;
        RECT 634.650 569.400 636.450 575.250 ;
        RECT 619.050 563.550 621.450 564.900 ;
        RECT 593.250 561.150 595.050 562.950 ;
        RECT 592.950 559.050 595.050 561.150 ;
        RECT 596.850 558.150 598.050 563.400 ;
        RECT 611.550 562.200 612.750 563.400 ;
        RECT 616.950 562.200 618.750 562.650 ;
        RECT 611.550 561.000 618.750 562.200 ;
        RECT 616.950 560.850 618.750 561.000 ;
        RECT 602.100 558.150 603.900 559.950 ;
        RECT 614.100 558.150 615.900 559.950 ;
        RECT 580.950 554.850 583.050 556.950 ;
        RECT 584.100 555.150 585.900 556.950 ;
        RECT 595.950 556.050 598.050 558.150 ;
        RECT 532.650 543.750 534.450 546.600 ;
        RECT 535.650 543.750 537.450 546.600 ;
        RECT 538.650 543.750 540.450 546.600 ;
        RECT 544.650 543.750 546.450 546.600 ;
        RECT 547.650 543.750 549.450 546.600 ;
        RECT 557.700 543.750 559.500 552.600 ;
        RECT 563.100 552.000 567.600 553.650 ;
        RECT 563.100 543.750 564.900 552.000 ;
        RECT 581.400 546.600 582.600 554.850 ;
        RECT 583.950 553.050 586.050 555.150 ;
        RECT 595.950 552.750 597.150 556.050 ;
        RECT 598.950 554.850 601.050 556.950 ;
        RECT 601.950 556.050 604.050 558.150 ;
        RECT 611.100 555.150 612.900 556.950 ;
        RECT 613.950 556.050 616.050 558.150 ;
        RECT 599.100 553.050 600.900 554.850 ;
        RECT 610.950 553.050 613.050 555.150 ;
        RECT 593.250 551.700 597.000 552.750 ;
        RECT 617.700 552.600 618.600 560.850 ;
        RECT 620.100 556.950 621.450 563.550 ;
        RECT 632.250 561.150 633.450 569.400 ;
        RECT 639.300 563.400 641.100 575.250 ;
        RECT 643.500 563.400 645.300 575.250 ;
        RECT 646.800 569.400 648.600 575.250 ;
        RECT 659.400 569.400 661.200 575.250 ;
        RECT 662.700 563.400 664.500 575.250 ;
        RECT 666.900 563.400 668.700 575.250 ;
        RECT 678.150 564.900 679.950 575.250 ;
        RECT 677.550 563.550 679.950 564.900 ;
        RECT 681.150 563.550 682.950 575.250 ;
        RECT 628.950 557.850 631.050 559.950 ;
        RECT 631.950 559.050 634.050 561.150 ;
        RECT 619.950 554.850 622.050 556.950 ;
        RECT 629.100 556.050 630.900 557.850 ;
        RECT 616.950 551.700 618.750 552.600 ;
        RECT 593.250 549.600 594.450 551.700 ;
        RECT 615.450 550.800 618.750 551.700 ;
        RECT 580.650 543.750 582.450 546.600 ;
        RECT 583.650 543.750 585.450 546.600 ;
        RECT 592.650 543.750 594.450 549.600 ;
        RECT 595.650 548.700 603.450 550.050 ;
        RECT 595.650 543.750 597.450 548.700 ;
        RECT 598.650 543.750 600.450 547.800 ;
        RECT 601.650 543.750 603.450 548.700 ;
        RECT 615.450 546.600 616.350 550.800 ;
        RECT 621.000 549.600 622.050 554.850 ;
        RECT 632.250 551.700 633.450 559.050 ;
        RECT 634.950 557.850 637.050 559.950 ;
        RECT 638.100 558.150 639.900 559.950 ;
        RECT 643.950 558.150 645.150 563.400 ;
        RECT 646.950 561.150 648.750 562.950 ;
        RECT 659.250 561.150 661.050 562.950 ;
        RECT 646.950 559.050 649.050 561.150 ;
        RECT 658.950 559.050 661.050 561.150 ;
        RECT 662.850 558.150 664.050 563.400 ;
        RECT 668.100 558.150 669.900 559.950 ;
        RECT 635.100 556.050 636.900 557.850 ;
        RECT 637.950 556.050 640.050 558.150 ;
        RECT 640.950 554.850 643.050 556.950 ;
        RECT 643.950 556.050 646.050 558.150 ;
        RECT 641.100 553.050 642.900 554.850 ;
        RECT 644.850 552.750 646.050 556.050 ;
        RECT 661.950 556.050 664.050 558.150 ;
        RECT 661.950 552.750 663.150 556.050 ;
        RECT 664.950 554.850 667.050 556.950 ;
        RECT 667.950 556.050 670.050 558.150 ;
        RECT 677.550 556.950 678.900 563.550 ;
        RECT 685.650 563.400 687.450 575.250 ;
        RECT 697.650 563.400 699.450 575.250 ;
        RECT 680.250 562.200 682.050 562.650 ;
        RECT 686.250 562.200 687.450 563.400 ;
        RECT 700.650 562.500 702.450 575.250 ;
        RECT 703.650 563.400 705.450 575.250 ;
        RECT 706.650 562.500 708.450 575.250 ;
        RECT 709.650 563.400 711.450 575.250 ;
        RECT 712.650 562.500 714.450 575.250 ;
        RECT 715.650 563.400 717.450 575.250 ;
        RECT 718.650 562.500 720.450 575.250 ;
        RECT 721.650 563.400 723.450 575.250 ;
        RECT 730.650 569.400 732.450 575.250 ;
        RECT 733.650 569.400 735.450 575.250 ;
        RECT 736.650 569.400 738.450 575.250 ;
        RECT 680.250 561.000 687.450 562.200 ;
        RECT 699.750 561.300 702.450 562.500 ;
        RECT 704.700 561.300 708.450 562.500 ;
        RECT 710.700 561.300 714.450 562.500 ;
        RECT 716.550 561.300 720.450 562.500 ;
        RECT 680.250 560.850 682.050 561.000 ;
        RECT 676.950 554.850 679.050 556.950 ;
        RECT 665.100 553.050 666.900 554.850 ;
        RECT 645.000 551.700 648.750 552.750 ;
        RECT 629.850 550.800 633.450 551.700 ;
        RECT 611.550 543.750 613.350 546.600 ;
        RECT 614.550 543.750 616.350 546.600 ;
        RECT 617.550 543.750 619.350 546.600 ;
        RECT 620.550 543.750 622.350 549.600 ;
        RECT 629.850 543.750 631.650 550.800 ;
        RECT 634.350 543.750 636.150 549.600 ;
        RECT 638.550 548.700 646.350 550.050 ;
        RECT 638.550 543.750 640.350 548.700 ;
        RECT 641.550 543.750 643.350 547.800 ;
        RECT 644.550 543.750 646.350 548.700 ;
        RECT 647.550 549.600 648.750 551.700 ;
        RECT 659.250 551.700 663.000 552.750 ;
        RECT 659.250 549.600 660.450 551.700 ;
        RECT 647.550 543.750 649.350 549.600 ;
        RECT 658.650 543.750 660.450 549.600 ;
        RECT 661.650 548.700 669.450 550.050 ;
        RECT 676.950 549.600 678.000 554.850 ;
        RECT 680.400 552.600 681.300 560.850 ;
        RECT 683.100 558.150 684.900 559.950 ;
        RECT 682.950 556.050 685.050 558.150 ;
        RECT 699.750 556.950 700.800 561.300 ;
        RECT 686.100 555.150 687.900 556.950 ;
        RECT 685.950 553.050 688.050 555.150 ;
        RECT 697.950 554.850 700.800 556.950 ;
        RECT 680.250 551.700 682.050 552.600 ;
        RECT 699.750 551.700 700.800 554.850 ;
        RECT 704.700 554.400 705.900 561.300 ;
        RECT 710.700 554.400 711.900 561.300 ;
        RECT 716.550 554.400 717.750 561.300 ;
        RECT 734.250 561.150 735.450 569.400 ;
        RECT 744.300 563.400 746.100 575.250 ;
        RECT 748.500 563.400 750.300 575.250 ;
        RECT 751.800 569.400 753.600 575.250 ;
        RECT 764.400 569.400 766.200 575.250 ;
        RECT 767.700 563.400 769.500 575.250 ;
        RECT 771.900 563.400 773.700 575.250 ;
        RECT 777.750 569.400 779.550 575.250 ;
        RECT 780.750 569.400 782.550 575.250 ;
        RECT 784.500 569.400 786.300 575.250 ;
        RECT 787.500 569.400 789.300 575.250 ;
        RECT 790.500 569.400 792.300 575.250 ;
        RECT 730.950 557.850 733.050 559.950 ;
        RECT 733.950 559.050 736.050 561.150 ;
        RECT 718.950 554.850 721.050 556.950 ;
        RECT 731.100 556.050 732.900 557.850 ;
        RECT 701.700 552.600 705.900 554.400 ;
        RECT 707.700 552.600 711.900 554.400 ;
        RECT 713.700 552.600 717.750 554.400 ;
        RECT 719.100 553.050 720.900 554.850 ;
        RECT 704.700 551.700 705.900 552.600 ;
        RECT 710.700 551.700 711.900 552.600 ;
        RECT 716.550 551.700 717.750 552.600 ;
        RECT 734.250 551.700 735.450 559.050 ;
        RECT 736.950 557.850 739.050 559.950 ;
        RECT 743.100 558.150 744.900 559.950 ;
        RECT 748.950 558.150 750.150 563.400 ;
        RECT 751.950 561.150 753.750 562.950 ;
        RECT 764.250 561.150 766.050 562.950 ;
        RECT 751.950 559.050 754.050 561.150 ;
        RECT 763.950 559.050 766.050 561.150 ;
        RECT 767.850 558.150 769.050 563.400 ;
        RECT 773.100 558.150 774.900 559.950 ;
        RECT 737.100 556.050 738.900 557.850 ;
        RECT 742.950 556.050 745.050 558.150 ;
        RECT 745.950 554.850 748.050 556.950 ;
        RECT 748.950 556.050 751.050 558.150 ;
        RECT 746.100 553.050 747.900 554.850 ;
        RECT 749.850 552.750 751.050 556.050 ;
        RECT 766.950 556.050 769.050 558.150 ;
        RECT 766.950 552.750 768.150 556.050 ;
        RECT 769.950 554.850 772.050 556.950 ;
        RECT 772.950 556.050 775.050 558.150 ;
        RECT 781.050 556.950 782.550 569.400 ;
        RECT 787.500 565.350 788.700 569.400 ;
        RECT 793.500 568.500 795.300 575.250 ;
        RECT 796.500 569.400 798.300 575.250 ;
        RECT 800.250 572.400 802.050 575.250 ;
        RECT 800.400 571.200 801.900 572.400 ;
        RECT 799.800 569.100 801.900 571.200 ;
        RECT 803.250 568.950 805.050 575.250 ;
        RECT 806.250 572.400 808.050 575.250 ;
        RECT 789.600 567.300 795.300 568.500 ;
        RECT 796.350 568.050 798.150 568.500 ;
        RECT 802.950 568.050 805.050 568.950 ;
        RECT 789.600 566.700 791.400 567.300 ;
        RECT 796.350 566.850 805.050 568.050 ;
        RECT 796.350 566.700 798.150 566.850 ;
        RECT 806.550 565.350 807.900 572.400 ;
        RECT 810.000 568.500 811.800 575.250 ;
        RECT 813.000 569.400 814.800 575.250 ;
        RECT 816.000 569.400 817.800 575.250 ;
        RECT 819.750 569.400 821.550 575.250 ;
        RECT 822.750 572.400 824.700 575.250 ;
        RECT 825.750 572.400 827.850 575.250 ;
        RECT 828.750 572.400 831.150 575.250 ;
        RECT 823.500 571.050 824.700 572.400 ;
        RECT 826.950 571.050 827.850 572.400 ;
        RECT 829.950 571.050 831.150 572.400 ;
        RECT 832.500 571.950 834.300 575.250 ;
        RECT 823.500 569.400 826.050 571.050 ;
        RECT 816.000 568.500 817.350 569.400 ;
        RECT 823.950 568.950 826.050 569.400 ;
        RECT 826.950 568.950 829.050 571.050 ;
        RECT 829.950 568.950 832.050 571.050 ;
        RECT 810.000 568.200 813.000 568.500 ;
        RECT 809.100 566.400 813.000 568.200 ;
        RECT 814.950 566.850 817.350 568.500 ;
        RECT 814.950 566.400 817.050 566.850 ;
        RECT 835.500 566.700 837.300 575.250 ;
        RECT 838.500 569.400 840.300 575.250 ;
        RECT 841.500 569.400 843.300 575.250 ;
        RECT 844.500 569.400 846.300 575.250 ;
        RECT 842.250 568.500 843.300 569.400 ;
        RECT 842.250 567.600 846.300 568.500 ;
        RECT 824.100 565.650 841.800 566.700 ;
        RECT 778.950 554.850 782.550 556.950 ;
        RECT 770.100 553.050 771.900 554.850 ;
        RECT 750.000 551.700 753.750 552.750 ;
        RECT 680.250 550.800 683.550 551.700 ;
        RECT 661.650 543.750 663.450 548.700 ;
        RECT 664.650 543.750 666.450 547.800 ;
        RECT 667.650 543.750 669.450 548.700 ;
        RECT 676.650 543.750 678.450 549.600 ;
        RECT 682.650 546.600 683.550 550.800 ;
        RECT 699.750 550.650 702.600 551.700 ;
        RECT 699.900 550.500 702.600 550.650 ;
        RECT 704.700 550.500 708.600 551.700 ;
        RECT 710.700 550.500 714.450 551.700 ;
        RECT 716.550 550.500 720.600 551.700 ;
        RECT 700.800 549.600 702.600 550.500 ;
        RECT 706.800 549.600 708.600 550.500 ;
        RECT 679.650 543.750 681.450 546.600 ;
        RECT 682.650 543.750 684.450 546.600 ;
        RECT 685.650 543.750 687.450 546.600 ;
        RECT 697.650 543.750 699.450 549.600 ;
        RECT 700.650 543.750 702.450 549.600 ;
        RECT 703.650 543.750 705.450 549.600 ;
        RECT 706.650 543.750 708.450 549.600 ;
        RECT 709.650 543.750 711.450 549.600 ;
        RECT 712.650 543.750 714.450 550.500 ;
        RECT 718.800 549.600 720.600 550.500 ;
        RECT 731.850 550.800 735.450 551.700 ;
        RECT 715.650 543.750 717.450 549.600 ;
        RECT 718.650 543.750 720.450 549.600 ;
        RECT 721.650 543.750 723.450 549.600 ;
        RECT 731.850 543.750 733.650 550.800 ;
        RECT 736.350 543.750 738.150 549.600 ;
        RECT 743.550 548.700 751.350 550.050 ;
        RECT 743.550 543.750 745.350 548.700 ;
        RECT 746.550 543.750 748.350 547.800 ;
        RECT 749.550 543.750 751.350 548.700 ;
        RECT 752.550 549.600 753.750 551.700 ;
        RECT 764.250 551.700 768.000 552.750 ;
        RECT 764.250 549.600 765.450 551.700 ;
        RECT 752.550 543.750 754.350 549.600 ;
        RECT 763.650 543.750 765.450 549.600 ;
        RECT 766.650 548.700 774.450 550.050 ;
        RECT 766.650 543.750 768.450 548.700 ;
        RECT 769.650 543.750 771.450 547.800 ;
        RECT 772.650 543.750 774.450 548.700 ;
        RECT 781.050 546.600 782.550 554.850 ;
        RECT 777.750 543.750 779.550 546.600 ;
        RECT 780.750 543.750 782.550 546.600 ;
        RECT 784.650 564.450 802.050 565.350 ;
        RECT 784.650 549.600 785.850 564.450 ;
        RECT 786.750 562.350 799.050 563.550 ;
        RECT 799.950 563.250 802.050 564.450 ;
        RECT 805.950 564.600 808.050 565.350 ;
        RECT 824.100 564.600 826.050 565.650 ;
        RECT 840.000 564.900 841.800 565.650 ;
        RECT 805.950 563.250 826.050 564.600 ;
        RECT 826.950 564.150 829.050 564.750 ;
        RECT 826.950 562.950 838.500 564.150 ;
        RECT 826.950 562.650 829.050 562.950 ;
        RECT 836.700 562.350 838.500 562.950 ;
        RECT 786.750 561.750 788.550 562.350 ;
        RECT 798.000 561.450 826.050 562.350 ;
        RECT 798.000 561.150 837.750 561.450 ;
        RECT 790.950 557.100 793.050 561.150 ;
        RECT 824.100 560.550 838.050 561.150 ;
        RECT 794.100 558.000 801.150 559.800 ;
        RECT 790.950 556.050 799.200 557.100 ;
        RECT 786.900 553.200 794.700 555.000 ;
        RECT 798.150 554.250 799.200 556.050 ;
        RECT 800.250 556.350 801.150 558.000 ;
        RECT 802.500 559.650 817.050 560.250 ;
        RECT 802.500 559.050 825.600 559.650 ;
        RECT 834.150 559.350 838.050 560.550 ;
        RECT 802.500 557.250 804.300 559.050 ;
        RECT 814.950 558.450 825.600 559.050 ;
        RECT 814.950 558.150 817.050 558.450 ;
        RECT 823.800 557.850 825.600 558.450 ;
        RECT 826.500 558.450 833.250 559.350 ;
        RECT 835.950 559.050 838.050 559.350 ;
        RECT 810.750 557.250 812.850 557.550 ;
        RECT 800.250 555.300 809.850 556.350 ;
        RECT 810.750 555.450 814.650 557.250 ;
        RECT 826.500 556.950 827.550 558.450 ;
        RECT 815.550 556.050 827.550 556.950 ;
        RECT 808.950 554.550 809.850 555.300 ;
        RECT 815.550 554.550 816.600 556.050 ;
        RECT 828.450 555.750 830.250 557.550 ;
        RECT 832.050 556.050 833.250 558.450 ;
        RECT 841.950 557.850 844.050 559.950 ;
        RECT 842.100 556.050 843.900 557.850 ;
        RECT 798.150 553.200 808.050 554.250 ;
        RECT 808.950 553.200 816.600 554.550 ;
        RECT 817.950 553.350 821.850 555.150 ;
        RECT 793.200 549.600 794.700 553.200 ;
        RECT 807.000 552.300 808.050 553.200 ;
        RECT 817.950 553.050 820.050 553.350 ;
        RECT 825.150 552.300 826.950 552.750 ;
        RECT 828.450 552.300 829.500 555.750 ;
        RECT 832.050 555.000 843.900 556.050 ;
        RECT 845.100 554.100 846.300 567.600 ;
        RECT 799.350 550.500 806.100 552.300 ;
        RECT 807.000 550.500 813.900 552.300 ;
        RECT 825.150 551.850 829.500 552.300 ;
        RECT 821.850 551.100 829.500 551.850 ;
        RECT 831.000 553.200 846.300 554.100 ;
        RECT 821.850 550.950 826.950 551.100 ;
        RECT 821.850 549.600 822.750 550.950 ;
        RECT 831.000 550.050 832.050 553.200 ;
        RECT 840.300 551.700 842.100 552.300 ;
        RECT 784.650 543.750 786.450 549.600 ;
        RECT 790.050 543.750 791.850 549.600 ;
        RECT 793.200 548.400 797.400 549.600 ;
        RECT 795.600 543.750 797.400 548.400 ;
        RECT 799.950 547.500 802.050 549.600 ;
        RECT 802.950 547.500 805.050 549.600 ;
        RECT 805.950 547.500 808.050 549.600 ;
        RECT 810.750 549.300 812.850 549.600 ;
        RECT 800.250 543.750 802.050 547.500 ;
        RECT 803.250 543.750 805.050 547.500 ;
        RECT 806.250 543.750 808.050 547.500 ;
        RECT 810.000 547.500 812.850 549.300 ;
        RECT 814.950 549.300 817.050 549.600 ;
        RECT 814.950 547.500 817.800 549.300 ;
        RECT 818.700 548.250 822.750 549.600 ;
        RECT 818.700 547.800 820.500 548.250 ;
        RECT 823.950 547.950 826.050 550.050 ;
        RECT 826.950 547.950 829.050 550.050 ;
        RECT 829.950 547.950 832.050 550.050 ;
        RECT 833.700 550.500 842.100 551.700 ;
        RECT 833.700 549.600 835.200 550.500 ;
        RECT 845.100 549.600 846.300 553.200 ;
        RECT 810.000 543.750 811.800 547.500 ;
        RECT 813.000 543.750 814.800 546.600 ;
        RECT 816.000 543.750 817.800 547.500 ;
        RECT 823.950 546.600 825.300 547.950 ;
        RECT 826.950 546.600 828.300 547.950 ;
        RECT 829.950 546.600 831.300 547.950 ;
        RECT 820.500 543.750 822.300 546.600 ;
        RECT 823.500 543.750 825.300 546.600 ;
        RECT 826.500 543.750 828.300 546.600 ;
        RECT 829.500 543.750 831.300 546.600 ;
        RECT 833.700 543.750 835.500 549.600 ;
        RECT 839.100 543.750 840.900 549.600 ;
        RECT 844.500 543.750 846.300 549.600 ;
        RECT 8.850 532.200 10.650 539.250 ;
        RECT 13.350 533.400 15.150 539.250 ;
        RECT 8.850 531.300 12.450 532.200 ;
        RECT 8.100 525.150 9.900 526.950 ;
        RECT 7.950 523.050 10.050 525.150 ;
        RECT 11.250 523.950 12.450 531.300 ;
        RECT 23.100 531.000 24.900 539.250 ;
        RECT 20.400 529.350 24.900 531.000 ;
        RECT 28.500 530.400 30.300 539.250 ;
        RECT 41.850 532.200 43.650 539.250 ;
        RECT 46.350 533.400 48.150 539.250 ;
        RECT 41.850 531.300 45.450 532.200 ;
        RECT 14.100 525.150 15.900 526.950 ;
        RECT 20.400 525.150 21.600 529.350 ;
        RECT 41.100 525.150 42.900 526.950 ;
        RECT 10.950 521.850 13.050 523.950 ;
        RECT 13.950 523.050 16.050 525.150 ;
        RECT 19.950 523.050 22.050 525.150 ;
        RECT 11.250 513.600 12.450 521.850 ;
        RECT 20.250 514.800 21.300 523.050 ;
        RECT 22.950 521.850 25.050 523.950 ;
        RECT 28.950 521.850 31.050 523.950 ;
        RECT 40.950 523.050 43.050 525.150 ;
        RECT 44.250 523.950 45.450 531.300 ;
        RECT 62.100 531.000 63.900 539.250 ;
        RECT 59.400 529.350 63.900 531.000 ;
        RECT 67.500 530.400 69.300 539.250 ;
        RECT 74.850 533.400 76.650 539.250 ;
        RECT 79.350 532.200 81.150 539.250 ;
        RECT 77.550 531.300 81.150 532.200 ;
        RECT 47.100 525.150 48.900 526.950 ;
        RECT 59.400 525.150 60.600 529.350 ;
        RECT 74.100 525.150 75.900 526.950 ;
        RECT 43.950 521.850 46.050 523.950 ;
        RECT 46.950 523.050 49.050 525.150 ;
        RECT 58.950 523.050 61.050 525.150 ;
        RECT 22.950 520.050 24.750 521.850 ;
        RECT 25.950 518.850 28.050 520.950 ;
        RECT 29.100 520.050 30.900 521.850 ;
        RECT 26.100 517.050 27.900 518.850 ;
        RECT 20.250 513.900 27.300 514.800 ;
        RECT 20.250 513.600 21.450 513.900 ;
        RECT 7.650 507.750 9.450 513.600 ;
        RECT 10.650 507.750 12.450 513.600 ;
        RECT 13.650 507.750 15.450 513.600 ;
        RECT 19.650 507.750 21.450 513.600 ;
        RECT 25.650 513.600 27.300 513.900 ;
        RECT 44.250 513.600 45.450 521.850 ;
        RECT 59.250 514.800 60.300 523.050 ;
        RECT 61.950 521.850 64.050 523.950 ;
        RECT 67.950 521.850 70.050 523.950 ;
        RECT 73.950 523.050 76.050 525.150 ;
        RECT 77.550 523.950 78.750 531.300 ;
        RECT 89.700 530.400 91.500 539.250 ;
        RECT 95.100 531.000 96.900 539.250 ;
        RECT 95.100 529.350 99.600 531.000 ;
        RECT 104.700 530.400 106.500 539.250 ;
        RECT 110.100 531.000 111.900 539.250 ;
        RECT 110.100 529.350 114.600 531.000 ;
        RECT 125.700 530.400 127.500 539.250 ;
        RECT 131.100 531.000 132.900 539.250 ;
        RECT 141.000 533.400 142.800 539.250 ;
        RECT 145.200 535.050 147.000 539.250 ;
        RECT 148.500 536.400 150.300 539.250 ;
        RECT 164.250 536.400 166.350 539.250 ;
        RECT 167.550 536.400 169.350 539.250 ;
        RECT 170.550 536.400 172.350 539.250 ;
        RECT 173.550 536.400 175.350 539.250 ;
        RECT 168.300 535.500 169.350 536.400 ;
        RECT 174.300 535.500 175.350 536.400 ;
        RECT 145.200 533.400 150.900 535.050 ;
        RECT 168.300 534.600 179.100 535.500 ;
        RECT 131.100 529.350 135.600 531.000 ;
        RECT 80.100 525.150 81.900 526.950 ;
        RECT 98.400 525.150 99.600 529.350 ;
        RECT 113.400 525.150 114.600 529.350 ;
        RECT 134.400 525.150 135.600 529.350 ;
        RECT 140.100 528.150 141.900 529.950 ;
        RECT 139.950 526.050 142.050 528.150 ;
        RECT 142.950 527.850 145.050 529.950 ;
        RECT 146.100 528.150 147.900 529.950 ;
        RECT 143.100 526.050 144.900 527.850 ;
        RECT 145.950 526.050 148.050 528.150 ;
        RECT 149.700 526.950 150.900 533.400 ;
        RECT 170.100 528.150 171.900 529.950 ;
        RECT 177.900 528.150 179.100 534.600 ;
        RECT 191.550 531.900 193.350 539.250 ;
        RECT 196.050 533.400 197.850 539.250 ;
        RECT 199.050 534.900 200.850 539.250 ;
        RECT 199.050 533.400 202.350 534.900 ;
        RECT 197.250 531.900 199.050 532.500 ;
        RECT 191.550 530.700 199.050 531.900 ;
        RECT 76.950 521.850 79.050 523.950 ;
        RECT 79.950 523.050 82.050 525.150 ;
        RECT 88.950 521.850 91.050 523.950 ;
        RECT 94.950 521.850 97.050 523.950 ;
        RECT 97.950 523.050 100.050 525.150 ;
        RECT 61.950 520.050 63.750 521.850 ;
        RECT 64.950 518.850 67.050 520.950 ;
        RECT 68.100 520.050 69.900 521.850 ;
        RECT 65.100 517.050 66.900 518.850 ;
        RECT 59.250 513.900 66.300 514.800 ;
        RECT 59.250 513.600 60.450 513.900 ;
        RECT 22.650 507.750 24.450 513.000 ;
        RECT 25.650 507.750 27.450 513.600 ;
        RECT 28.650 507.750 30.450 513.600 ;
        RECT 40.650 507.750 42.450 513.600 ;
        RECT 43.650 507.750 45.450 513.600 ;
        RECT 46.650 507.750 48.450 513.600 ;
        RECT 58.650 507.750 60.450 513.600 ;
        RECT 64.650 513.600 66.300 513.900 ;
        RECT 77.550 513.600 78.750 521.850 ;
        RECT 89.100 520.050 90.900 521.850 ;
        RECT 91.950 518.850 94.050 520.950 ;
        RECT 95.250 520.050 97.050 521.850 ;
        RECT 92.100 517.050 93.900 518.850 ;
        RECT 98.700 514.800 99.750 523.050 ;
        RECT 103.950 521.850 106.050 523.950 ;
        RECT 109.950 521.850 112.050 523.950 ;
        RECT 112.950 523.050 115.050 525.150 ;
        RECT 104.100 520.050 105.900 521.850 ;
        RECT 106.950 518.850 109.050 520.950 ;
        RECT 110.250 520.050 112.050 521.850 ;
        RECT 107.100 517.050 108.900 518.850 ;
        RECT 113.700 514.800 114.750 523.050 ;
        RECT 124.950 521.850 127.050 523.950 ;
        RECT 130.950 521.850 133.050 523.950 ;
        RECT 133.950 523.050 136.050 525.150 ;
        RECT 148.950 524.850 151.050 526.950 ;
        RECT 163.950 524.850 166.050 526.950 ;
        RECT 169.950 526.050 172.050 528.150 ;
        RECT 172.950 524.850 175.050 526.950 ;
        RECT 177.900 526.050 181.050 528.150 ;
        RECT 125.100 520.050 126.900 521.850 ;
        RECT 127.950 518.850 130.050 520.950 ;
        RECT 131.250 520.050 133.050 521.850 ;
        RECT 128.100 517.050 129.900 518.850 ;
        RECT 134.700 514.800 135.750 523.050 ;
        RECT 149.700 519.600 150.900 524.850 ;
        RECT 164.100 523.050 165.900 524.850 ;
        RECT 173.100 523.050 174.900 524.850 ;
        RECT 177.900 520.800 179.100 526.050 ;
        RECT 190.950 524.850 193.050 526.950 ;
        RECT 191.100 523.050 192.900 524.850 ;
        RECT 177.900 519.600 181.350 520.800 ;
        RECT 92.700 513.900 99.750 514.800 ;
        RECT 92.700 513.600 94.350 513.900 ;
        RECT 61.650 507.750 63.450 513.000 ;
        RECT 64.650 507.750 66.450 513.600 ;
        RECT 67.650 507.750 69.450 513.600 ;
        RECT 74.550 507.750 76.350 513.600 ;
        RECT 77.550 507.750 79.350 513.600 ;
        RECT 80.550 507.750 82.350 513.600 ;
        RECT 89.550 507.750 91.350 513.600 ;
        RECT 92.550 507.750 94.350 513.600 ;
        RECT 98.550 513.600 99.750 513.900 ;
        RECT 107.700 513.900 114.750 514.800 ;
        RECT 107.700 513.600 109.350 513.900 ;
        RECT 95.550 507.750 97.350 513.000 ;
        RECT 98.550 507.750 100.350 513.600 ;
        RECT 104.550 507.750 106.350 513.600 ;
        RECT 107.550 507.750 109.350 513.600 ;
        RECT 113.550 513.600 114.750 513.900 ;
        RECT 128.700 513.900 135.750 514.800 ;
        RECT 128.700 513.600 130.350 513.900 ;
        RECT 110.550 507.750 112.350 513.000 ;
        RECT 113.550 507.750 115.350 513.600 ;
        RECT 125.550 507.750 127.350 513.600 ;
        RECT 128.550 507.750 130.350 513.600 ;
        RECT 134.550 513.600 135.750 513.900 ;
        RECT 140.550 518.700 148.350 519.600 ;
        RECT 131.550 507.750 133.350 513.000 ;
        RECT 134.550 507.750 136.350 513.600 ;
        RECT 140.550 507.750 142.350 518.700 ;
        RECT 143.550 507.750 145.350 517.800 ;
        RECT 146.550 507.750 148.350 518.700 ;
        RECT 149.550 507.750 151.350 519.600 ;
        RECT 161.550 517.500 169.350 518.400 ;
        RECT 161.550 507.750 163.350 517.500 ;
        RECT 164.550 507.750 166.350 516.600 ;
        RECT 167.550 508.500 169.350 517.500 ;
        RECT 170.550 517.200 178.950 518.100 ;
        RECT 170.550 509.400 172.350 517.200 ;
        RECT 173.550 508.500 175.350 516.300 ;
        RECT 167.550 507.750 175.350 508.500 ;
        RECT 177.150 508.500 178.950 517.200 ;
        RECT 180.150 517.200 181.350 519.600 ;
        RECT 180.150 509.400 181.950 517.200 ;
        RECT 183.150 508.500 184.950 517.800 ;
        RECT 194.700 513.600 195.900 530.700 ;
        RECT 201.150 526.950 202.350 533.400 ;
        RECT 212.850 532.200 214.650 539.250 ;
        RECT 217.350 533.400 219.150 539.250 ;
        RECT 226.650 536.400 228.450 539.250 ;
        RECT 229.650 536.400 231.450 539.250 ;
        RECT 232.650 536.400 234.450 539.250 ;
        RECT 212.850 531.300 216.450 532.200 ;
        RECT 197.100 525.150 198.900 526.950 ;
        RECT 196.950 523.050 199.050 525.150 ;
        RECT 199.950 524.850 202.350 526.950 ;
        RECT 212.100 525.150 213.900 526.950 ;
        RECT 201.150 519.600 202.350 524.850 ;
        RECT 211.950 523.050 214.050 525.150 ;
        RECT 215.250 523.950 216.450 531.300 ;
        RECT 229.950 529.950 231.000 536.400 ;
        RECT 242.100 531.000 243.900 539.250 ;
        RECT 229.950 527.850 232.050 529.950 ;
        RECT 239.400 529.350 243.900 531.000 ;
        RECT 247.500 530.400 249.300 539.250 ;
        RECT 257.550 536.400 259.350 539.250 ;
        RECT 260.550 536.400 262.350 539.250 ;
        RECT 263.550 536.400 265.350 539.250 ;
        RECT 261.000 529.950 262.050 536.400 ;
        RECT 272.550 531.900 274.350 539.250 ;
        RECT 277.050 533.400 278.850 539.250 ;
        RECT 280.050 534.900 281.850 539.250 ;
        RECT 280.050 533.400 283.350 534.900 ;
        RECT 278.250 531.900 280.050 532.500 ;
        RECT 272.550 530.700 280.050 531.900 ;
        RECT 218.100 525.150 219.900 526.950 ;
        RECT 214.950 521.850 217.050 523.950 ;
        RECT 217.950 523.050 220.050 525.150 ;
        RECT 226.950 524.850 229.050 526.950 ;
        RECT 227.100 523.050 228.900 524.850 ;
        RECT 177.150 507.750 184.950 508.500 ;
        RECT 191.550 507.750 193.350 513.600 ;
        RECT 194.550 507.750 196.350 513.600 ;
        RECT 198.150 507.750 199.950 519.600 ;
        RECT 201.150 507.750 202.950 519.600 ;
        RECT 215.250 513.600 216.450 521.850 ;
        RECT 229.950 520.650 231.000 527.850 ;
        RECT 232.950 524.850 235.050 526.950 ;
        RECT 239.400 525.150 240.600 529.350 ;
        RECT 259.950 527.850 262.050 529.950 ;
        RECT 233.100 523.050 234.900 524.850 ;
        RECT 238.950 523.050 241.050 525.150 ;
        RECT 256.950 524.850 259.050 526.950 ;
        RECT 228.450 519.600 231.000 520.650 ;
        RECT 211.650 507.750 213.450 513.600 ;
        RECT 214.650 507.750 216.450 513.600 ;
        RECT 217.650 507.750 219.450 513.600 ;
        RECT 228.450 507.750 230.250 519.600 ;
        RECT 232.650 507.750 234.450 519.600 ;
        RECT 239.250 514.800 240.300 523.050 ;
        RECT 241.950 521.850 244.050 523.950 ;
        RECT 247.950 521.850 250.050 523.950 ;
        RECT 257.100 523.050 258.900 524.850 ;
        RECT 241.950 520.050 243.750 521.850 ;
        RECT 244.950 518.850 247.050 520.950 ;
        RECT 248.100 520.050 249.900 521.850 ;
        RECT 261.000 520.650 262.050 527.850 ;
        RECT 262.950 524.850 265.050 526.950 ;
        RECT 271.950 524.850 274.050 526.950 ;
        RECT 263.100 523.050 264.900 524.850 ;
        RECT 272.100 523.050 273.900 524.850 ;
        RECT 261.000 519.600 263.550 520.650 ;
        RECT 245.100 517.050 246.900 518.850 ;
        RECT 239.250 513.900 246.300 514.800 ;
        RECT 239.250 513.600 240.450 513.900 ;
        RECT 238.650 507.750 240.450 513.600 ;
        RECT 244.650 513.600 246.300 513.900 ;
        RECT 241.650 507.750 243.450 513.000 ;
        RECT 244.650 507.750 246.450 513.600 ;
        RECT 247.650 507.750 249.450 513.600 ;
        RECT 257.550 507.750 259.350 519.600 ;
        RECT 261.750 507.750 263.550 519.600 ;
        RECT 275.700 513.600 276.900 530.700 ;
        RECT 282.150 526.950 283.350 533.400 ;
        RECT 287.700 530.400 289.500 539.250 ;
        RECT 293.100 531.000 294.900 539.250 ;
        RECT 308.550 531.900 310.350 539.250 ;
        RECT 313.050 533.400 314.850 539.250 ;
        RECT 316.050 534.900 317.850 539.250 ;
        RECT 316.050 533.400 319.350 534.900 ;
        RECT 314.250 531.900 316.050 532.500 ;
        RECT 293.100 529.350 297.600 531.000 ;
        RECT 308.550 530.700 316.050 531.900 ;
        RECT 278.100 525.150 279.900 526.950 ;
        RECT 277.950 523.050 280.050 525.150 ;
        RECT 280.950 524.850 283.350 526.950 ;
        RECT 296.400 525.150 297.600 529.350 ;
        RECT 282.150 519.600 283.350 524.850 ;
        RECT 286.950 521.850 289.050 523.950 ;
        RECT 292.950 521.850 295.050 523.950 ;
        RECT 295.950 523.050 298.050 525.150 ;
        RECT 307.950 524.850 310.050 526.950 ;
        RECT 308.100 523.050 309.900 524.850 ;
        RECT 287.100 520.050 288.900 521.850 ;
        RECT 272.550 507.750 274.350 513.600 ;
        RECT 275.550 507.750 277.350 513.600 ;
        RECT 279.150 507.750 280.950 519.600 ;
        RECT 282.150 507.750 283.950 519.600 ;
        RECT 289.950 518.850 292.050 520.950 ;
        RECT 293.250 520.050 295.050 521.850 ;
        RECT 290.100 517.050 291.900 518.850 ;
        RECT 296.700 514.800 297.750 523.050 ;
        RECT 290.700 513.900 297.750 514.800 ;
        RECT 290.700 513.600 292.350 513.900 ;
        RECT 287.550 507.750 289.350 513.600 ;
        RECT 290.550 507.750 292.350 513.600 ;
        RECT 296.550 513.600 297.750 513.900 ;
        RECT 311.700 513.600 312.900 530.700 ;
        RECT 318.150 526.950 319.350 533.400 ;
        RECT 326.700 530.400 328.500 539.250 ;
        RECT 332.100 531.000 333.900 539.250 ;
        RECT 350.850 532.200 352.650 539.250 ;
        RECT 355.350 533.400 357.150 539.250 ;
        RECT 359.550 536.400 361.350 539.250 ;
        RECT 362.550 536.400 364.350 539.250 ;
        RECT 365.550 536.400 367.350 539.250 ;
        RECT 363.450 532.200 364.350 536.400 ;
        RECT 368.550 533.400 370.350 539.250 ;
        RECT 383.700 536.400 385.500 539.250 ;
        RECT 387.000 535.050 388.800 539.250 ;
        RECT 383.100 533.400 388.800 535.050 ;
        RECT 391.200 533.400 393.000 539.250 ;
        RECT 398.550 534.300 400.350 539.250 ;
        RECT 401.550 535.200 403.350 539.250 ;
        RECT 404.550 534.300 406.350 539.250 ;
        RECT 350.850 531.300 354.450 532.200 ;
        RECT 363.450 531.300 366.750 532.200 ;
        RECT 332.100 529.350 336.600 531.000 ;
        RECT 314.100 525.150 315.900 526.950 ;
        RECT 313.950 523.050 316.050 525.150 ;
        RECT 316.950 524.850 319.350 526.950 ;
        RECT 335.400 525.150 336.600 529.350 ;
        RECT 350.100 525.150 351.900 526.950 ;
        RECT 318.150 519.600 319.350 524.850 ;
        RECT 325.950 521.850 328.050 523.950 ;
        RECT 331.950 521.850 334.050 523.950 ;
        RECT 334.950 523.050 337.050 525.150 ;
        RECT 349.950 523.050 352.050 525.150 ;
        RECT 353.250 523.950 354.450 531.300 ;
        RECT 364.950 530.400 366.750 531.300 ;
        RECT 358.950 527.850 361.050 529.950 ;
        RECT 356.100 525.150 357.900 526.950 ;
        RECT 359.100 526.050 360.900 527.850 ;
        RECT 326.100 520.050 327.900 521.850 ;
        RECT 293.550 507.750 295.350 513.000 ;
        RECT 296.550 507.750 298.350 513.600 ;
        RECT 308.550 507.750 310.350 513.600 ;
        RECT 311.550 507.750 313.350 513.600 ;
        RECT 315.150 507.750 316.950 519.600 ;
        RECT 318.150 507.750 319.950 519.600 ;
        RECT 328.950 518.850 331.050 520.950 ;
        RECT 332.250 520.050 334.050 521.850 ;
        RECT 329.100 517.050 330.900 518.850 ;
        RECT 335.700 514.800 336.750 523.050 ;
        RECT 352.950 521.850 355.050 523.950 ;
        RECT 355.950 523.050 358.050 525.150 ;
        RECT 361.950 524.850 364.050 526.950 ;
        RECT 362.100 523.050 363.900 524.850 ;
        RECT 365.700 522.150 366.600 530.400 ;
        RECT 369.000 528.150 370.050 533.400 ;
        RECT 367.950 526.050 370.050 528.150 ;
        RECT 383.100 526.950 384.300 533.400 ;
        RECT 398.550 532.950 406.350 534.300 ;
        RECT 407.550 533.400 409.350 539.250 ;
        RECT 416.550 534.300 418.350 539.250 ;
        RECT 419.550 535.200 421.350 539.250 ;
        RECT 422.550 534.300 424.350 539.250 ;
        RECT 407.550 531.300 408.750 533.400 ;
        RECT 416.550 532.950 424.350 534.300 ;
        RECT 425.550 533.400 427.350 539.250 ;
        RECT 432.750 536.400 434.550 539.250 ;
        RECT 435.750 536.400 437.550 539.250 ;
        RECT 425.550 531.300 426.750 533.400 ;
        RECT 405.000 530.250 408.750 531.300 ;
        RECT 423.000 530.250 426.750 531.300 ;
        RECT 386.100 528.150 387.900 529.950 ;
        RECT 364.950 522.000 366.750 522.150 ;
        RECT 329.700 513.900 336.750 514.800 ;
        RECT 329.700 513.600 331.350 513.900 ;
        RECT 326.550 507.750 328.350 513.600 ;
        RECT 329.550 507.750 331.350 513.600 ;
        RECT 335.550 513.600 336.750 513.900 ;
        RECT 353.250 513.600 354.450 521.850 ;
        RECT 359.550 520.800 366.750 522.000 ;
        RECT 359.550 519.600 360.750 520.800 ;
        RECT 364.950 520.350 366.750 520.800 ;
        RECT 332.550 507.750 334.350 513.000 ;
        RECT 335.550 507.750 337.350 513.600 ;
        RECT 349.650 507.750 351.450 513.600 ;
        RECT 352.650 507.750 354.450 513.600 ;
        RECT 355.650 507.750 357.450 513.600 ;
        RECT 359.550 507.750 361.350 519.600 ;
        RECT 368.100 519.450 369.450 526.050 ;
        RECT 382.950 524.850 385.050 526.950 ;
        RECT 385.950 526.050 388.050 528.150 ;
        RECT 388.950 527.850 391.050 529.950 ;
        RECT 392.100 528.150 393.900 529.950 ;
        RECT 401.100 528.150 402.900 529.950 ;
        RECT 389.100 526.050 390.900 527.850 ;
        RECT 391.950 526.050 394.050 528.150 ;
        RECT 397.950 524.850 400.050 526.950 ;
        RECT 400.950 526.050 403.050 528.150 ;
        RECT 404.850 526.950 406.050 530.250 ;
        RECT 419.100 528.150 420.900 529.950 ;
        RECT 403.950 524.850 406.050 526.950 ;
        RECT 415.950 524.850 418.050 526.950 ;
        RECT 418.950 526.050 421.050 528.150 ;
        RECT 422.850 526.950 424.050 530.250 ;
        RECT 436.050 528.150 437.550 536.400 ;
        RECT 421.950 524.850 424.050 526.950 ;
        RECT 433.950 526.050 437.550 528.150 ;
        RECT 383.100 519.600 384.300 524.850 ;
        RECT 398.100 523.050 399.900 524.850 ;
        RECT 403.950 519.600 405.150 524.850 ;
        RECT 406.950 521.850 409.050 523.950 ;
        RECT 416.100 523.050 417.900 524.850 ;
        RECT 406.950 520.050 408.750 521.850 ;
        RECT 421.950 519.600 423.150 524.850 ;
        RECT 424.950 521.850 427.050 523.950 ;
        RECT 424.950 520.050 426.750 521.850 ;
        RECT 364.050 507.750 365.850 519.450 ;
        RECT 367.050 518.100 369.450 519.450 ;
        RECT 367.050 507.750 368.850 518.100 ;
        RECT 382.650 507.750 384.450 519.600 ;
        RECT 385.650 518.700 393.450 519.600 ;
        RECT 385.650 507.750 387.450 518.700 ;
        RECT 388.650 507.750 390.450 517.800 ;
        RECT 391.650 507.750 393.450 518.700 ;
        RECT 399.300 507.750 401.100 519.600 ;
        RECT 403.500 507.750 405.300 519.600 ;
        RECT 406.800 507.750 408.600 513.600 ;
        RECT 417.300 507.750 419.100 519.600 ;
        RECT 421.500 507.750 423.300 519.600 ;
        RECT 436.050 513.600 437.550 526.050 ;
        RECT 439.650 533.400 441.450 539.250 ;
        RECT 445.050 533.400 446.850 539.250 ;
        RECT 450.600 534.600 452.400 539.250 ;
        RECT 455.250 535.500 457.050 539.250 ;
        RECT 458.250 535.500 460.050 539.250 ;
        RECT 461.250 535.500 463.050 539.250 ;
        RECT 448.200 533.400 452.400 534.600 ;
        RECT 454.950 533.400 457.050 535.500 ;
        RECT 457.950 533.400 460.050 535.500 ;
        RECT 460.950 533.400 463.050 535.500 ;
        RECT 465.000 535.500 466.800 539.250 ;
        RECT 468.000 536.400 469.800 539.250 ;
        RECT 471.000 535.500 472.800 539.250 ;
        RECT 475.500 536.400 477.300 539.250 ;
        RECT 478.500 536.400 480.300 539.250 ;
        RECT 481.500 536.400 483.300 539.250 ;
        RECT 484.500 536.400 486.300 539.250 ;
        RECT 465.000 533.700 467.850 535.500 ;
        RECT 465.750 533.400 467.850 533.700 ;
        RECT 469.950 533.700 472.800 535.500 ;
        RECT 473.700 534.750 475.500 535.200 ;
        RECT 478.950 535.050 480.300 536.400 ;
        RECT 481.950 535.050 483.300 536.400 ;
        RECT 484.950 535.050 486.300 536.400 ;
        RECT 469.950 533.400 472.050 533.700 ;
        RECT 473.700 533.400 477.750 534.750 ;
        RECT 439.650 518.550 440.850 533.400 ;
        RECT 448.200 529.800 449.700 533.400 ;
        RECT 454.350 530.700 461.100 532.500 ;
        RECT 462.000 530.700 468.900 532.500 ;
        RECT 476.850 532.050 477.750 533.400 ;
        RECT 478.950 532.950 481.050 535.050 ;
        RECT 481.950 532.950 484.050 535.050 ;
        RECT 484.950 532.950 487.050 535.050 ;
        RECT 476.850 531.900 481.950 532.050 ;
        RECT 476.850 531.150 484.500 531.900 ;
        RECT 480.150 530.700 484.500 531.150 ;
        RECT 462.000 529.800 463.050 530.700 ;
        RECT 480.150 530.250 481.950 530.700 ;
        RECT 441.900 528.000 449.700 529.800 ;
        RECT 453.150 528.750 463.050 529.800 ;
        RECT 453.150 526.950 454.200 528.750 ;
        RECT 463.950 528.450 471.600 529.800 ;
        RECT 463.950 527.700 464.850 528.450 ;
        RECT 445.950 525.900 454.200 526.950 ;
        RECT 455.250 526.650 464.850 527.700 ;
        RECT 445.950 521.850 448.050 525.900 ;
        RECT 455.250 525.000 456.150 526.650 ;
        RECT 465.750 525.750 469.650 527.550 ;
        RECT 470.550 526.950 471.600 528.450 ;
        RECT 472.950 529.650 475.050 529.950 ;
        RECT 472.950 527.850 476.850 529.650 ;
        RECT 483.450 527.250 484.500 530.700 ;
        RECT 486.000 529.800 487.050 532.950 ;
        RECT 488.700 533.400 490.500 539.250 ;
        RECT 494.100 533.400 495.900 539.250 ;
        RECT 499.500 533.400 501.300 539.250 ;
        RECT 504.000 533.400 505.800 539.250 ;
        RECT 508.200 533.400 510.000 539.250 ;
        RECT 512.400 533.400 514.200 539.250 ;
        RECT 488.700 532.500 490.200 533.400 ;
        RECT 488.700 531.300 497.100 532.500 ;
        RECT 495.300 530.700 497.100 531.300 ;
        RECT 500.100 529.800 501.300 533.400 ;
        RECT 486.000 528.900 501.300 529.800 ;
        RECT 470.550 526.050 482.550 526.950 ;
        RECT 449.100 523.200 456.150 525.000 ;
        RECT 457.500 523.950 459.300 525.750 ;
        RECT 465.750 525.450 467.850 525.750 ;
        RECT 469.950 524.550 472.050 524.850 ;
        RECT 478.800 524.550 480.600 525.150 ;
        RECT 469.950 523.950 480.600 524.550 ;
        RECT 457.500 523.350 480.600 523.950 ;
        RECT 481.500 524.550 482.550 526.050 ;
        RECT 483.450 525.450 485.250 527.250 ;
        RECT 487.050 526.950 498.900 528.000 ;
        RECT 487.050 524.550 488.250 526.950 ;
        RECT 497.100 525.150 498.900 526.950 ;
        RECT 481.500 523.650 488.250 524.550 ;
        RECT 490.950 523.650 493.050 523.950 ;
        RECT 457.500 522.750 472.050 523.350 ;
        RECT 489.150 522.450 493.050 523.650 ;
        RECT 496.950 523.050 499.050 525.150 ;
        RECT 479.100 521.850 493.050 522.450 ;
        RECT 453.000 521.550 492.750 521.850 ;
        RECT 441.750 520.650 443.550 521.250 ;
        RECT 453.000 520.650 481.050 521.550 ;
        RECT 441.750 519.450 454.050 520.650 ;
        RECT 481.950 520.050 484.050 520.350 ;
        RECT 491.700 520.050 493.500 520.650 ;
        RECT 454.950 518.550 457.050 519.750 ;
        RECT 439.650 517.650 457.050 518.550 ;
        RECT 460.950 518.400 481.050 519.750 ;
        RECT 460.950 517.650 463.050 518.400 ;
        RECT 442.500 513.600 443.700 517.650 ;
        RECT 444.600 515.700 446.400 516.300 ;
        RECT 451.350 516.150 453.150 516.300 ;
        RECT 444.600 514.500 450.300 515.700 ;
        RECT 451.350 514.950 460.050 516.150 ;
        RECT 451.350 514.500 453.150 514.950 ;
        RECT 424.800 507.750 426.600 513.600 ;
        RECT 432.750 507.750 434.550 513.600 ;
        RECT 435.750 507.750 437.550 513.600 ;
        RECT 439.500 507.750 441.300 513.600 ;
        RECT 442.500 507.750 444.300 513.600 ;
        RECT 445.500 507.750 447.300 513.600 ;
        RECT 448.500 507.750 450.300 514.500 ;
        RECT 457.950 514.050 460.050 514.950 ;
        RECT 451.500 507.750 453.300 513.600 ;
        RECT 454.800 511.800 456.900 513.900 ;
        RECT 455.400 510.600 456.900 511.800 ;
        RECT 455.250 507.750 457.050 510.600 ;
        RECT 458.250 507.750 460.050 514.050 ;
        RECT 461.550 510.600 462.900 517.650 ;
        RECT 479.100 517.350 481.050 518.400 ;
        RECT 481.950 518.850 493.500 520.050 ;
        RECT 481.950 518.250 484.050 518.850 ;
        RECT 495.000 517.350 496.800 518.100 ;
        RECT 464.100 514.800 468.000 516.600 ;
        RECT 465.000 514.500 468.000 514.800 ;
        RECT 469.950 516.150 472.050 516.600 ;
        RECT 479.100 516.300 496.800 517.350 ;
        RECT 469.950 514.500 472.350 516.150 ;
        RECT 461.250 507.750 463.050 510.600 ;
        RECT 465.000 507.750 466.800 514.500 ;
        RECT 471.000 513.600 472.350 514.500 ;
        RECT 478.950 513.600 481.050 514.050 ;
        RECT 468.000 507.750 469.800 513.600 ;
        RECT 471.000 507.750 472.800 513.600 ;
        RECT 474.750 507.750 476.550 513.600 ;
        RECT 478.500 511.950 481.050 513.600 ;
        RECT 481.950 511.950 484.050 514.050 ;
        RECT 484.950 511.950 487.050 514.050 ;
        RECT 478.500 510.600 479.700 511.950 ;
        RECT 481.950 510.600 482.850 511.950 ;
        RECT 484.950 510.600 486.150 511.950 ;
        RECT 477.750 507.750 479.700 510.600 ;
        RECT 480.750 507.750 482.850 510.600 ;
        RECT 483.750 507.750 486.150 510.600 ;
        RECT 487.500 507.750 489.300 511.050 ;
        RECT 490.500 507.750 492.300 516.300 ;
        RECT 500.100 515.400 501.300 528.900 ;
        RECT 506.250 528.150 508.050 529.950 ;
        RECT 502.950 524.850 505.050 526.950 ;
        RECT 505.950 526.050 508.050 528.150 ;
        RECT 508.950 526.950 510.000 533.400 ;
        RECT 527.700 530.400 529.500 539.250 ;
        RECT 533.100 531.000 534.900 539.250 ;
        RECT 549.000 533.400 550.800 539.250 ;
        RECT 553.200 533.400 555.000 539.250 ;
        RECT 557.400 533.400 559.200 539.250 ;
        RECT 572.550 536.400 574.350 539.250 ;
        RECT 575.550 536.400 577.350 539.250 ;
        RECT 511.950 528.150 513.750 529.950 ;
        RECT 533.100 529.350 537.600 531.000 ;
        RECT 508.950 524.850 511.050 526.950 ;
        RECT 511.950 526.050 514.050 528.150 ;
        RECT 514.950 524.850 517.050 526.950 ;
        RECT 536.400 525.150 537.600 529.350 ;
        RECT 551.250 528.150 553.050 529.950 ;
        RECT 503.250 523.050 505.050 524.850 ;
        RECT 510.150 521.400 511.050 524.850 ;
        RECT 515.100 523.050 516.900 524.850 ;
        RECT 526.950 521.850 529.050 523.950 ;
        RECT 532.950 521.850 535.050 523.950 ;
        RECT 535.950 523.050 538.050 525.150 ;
        RECT 547.950 524.850 550.050 526.950 ;
        RECT 550.950 526.050 553.050 528.150 ;
        RECT 553.950 526.950 555.000 533.400 ;
        RECT 556.950 528.150 558.750 529.950 ;
        RECT 553.950 524.850 556.050 526.950 ;
        RECT 556.950 526.050 559.050 528.150 ;
        RECT 571.950 527.850 574.050 529.950 ;
        RECT 575.400 528.150 576.600 536.400 ;
        RECT 587.850 532.200 589.650 539.250 ;
        RECT 592.350 533.400 594.150 539.250 ;
        RECT 599.550 536.400 601.350 539.250 ;
        RECT 602.550 536.400 604.350 539.250 ;
        RECT 605.550 536.400 607.350 539.250 ;
        RECT 614.550 536.400 616.350 539.250 ;
        RECT 617.550 536.400 619.350 539.250 ;
        RECT 620.550 536.400 622.350 539.250 ;
        RECT 626.550 536.400 628.350 539.250 ;
        RECT 629.550 536.400 631.350 539.250 ;
        RECT 587.850 531.300 591.450 532.200 ;
        RECT 559.950 524.850 562.050 526.950 ;
        RECT 572.100 526.050 573.900 527.850 ;
        RECT 574.950 526.050 577.050 528.150 ;
        RECT 548.250 523.050 550.050 524.850 ;
        RECT 510.150 520.500 514.200 521.400 ;
        RECT 512.400 519.600 514.200 520.500 ;
        RECT 527.100 520.050 528.900 521.850 ;
        RECT 497.250 514.500 501.300 515.400 ;
        RECT 503.550 518.400 511.350 519.300 ;
        RECT 497.250 513.600 498.300 514.500 ;
        RECT 493.500 507.750 495.300 513.600 ;
        RECT 496.500 507.750 498.300 513.600 ;
        RECT 499.500 507.750 501.300 513.600 ;
        RECT 503.550 507.750 505.350 518.400 ;
        RECT 506.550 507.750 508.350 517.500 ;
        RECT 509.550 508.500 511.350 518.400 ;
        RECT 512.550 509.400 514.350 519.600 ;
        RECT 515.550 508.500 517.350 519.600 ;
        RECT 529.950 518.850 532.050 520.950 ;
        RECT 533.250 520.050 535.050 521.850 ;
        RECT 530.100 517.050 531.900 518.850 ;
        RECT 536.700 514.800 537.750 523.050 ;
        RECT 555.150 521.400 556.050 524.850 ;
        RECT 560.100 523.050 561.900 524.850 ;
        RECT 555.150 520.500 559.200 521.400 ;
        RECT 557.400 519.600 559.200 520.500 ;
        RECT 530.700 513.900 537.750 514.800 ;
        RECT 530.700 513.600 532.350 513.900 ;
        RECT 509.550 507.750 517.350 508.500 ;
        RECT 527.550 507.750 529.350 513.600 ;
        RECT 530.550 507.750 532.350 513.600 ;
        RECT 536.550 513.600 537.750 513.900 ;
        RECT 548.550 518.400 556.350 519.300 ;
        RECT 533.550 507.750 535.350 513.000 ;
        RECT 536.550 507.750 538.350 513.600 ;
        RECT 548.550 507.750 550.350 518.400 ;
        RECT 551.550 507.750 553.350 517.500 ;
        RECT 554.550 508.500 556.350 518.400 ;
        RECT 557.550 509.400 559.350 519.600 ;
        RECT 560.550 508.500 562.350 519.600 ;
        RECT 575.400 513.600 576.600 526.050 ;
        RECT 587.100 525.150 588.900 526.950 ;
        RECT 586.950 523.050 589.050 525.150 ;
        RECT 590.250 523.950 591.450 531.300 ;
        RECT 603.000 529.950 604.050 536.400 ;
        RECT 604.950 531.450 607.050 532.050 ;
        RECT 604.950 530.550 609.450 531.450 ;
        RECT 604.950 529.950 607.050 530.550 ;
        RECT 601.950 527.850 604.050 529.950 ;
        RECT 608.550 529.050 609.450 530.550 ;
        RECT 618.000 529.950 619.050 536.400 ;
        RECT 593.100 525.150 594.900 526.950 ;
        RECT 589.950 521.850 592.050 523.950 ;
        RECT 592.950 523.050 595.050 525.150 ;
        RECT 598.950 524.850 601.050 526.950 ;
        RECT 599.100 523.050 600.900 524.850 ;
        RECT 590.250 513.600 591.450 521.850 ;
        RECT 603.000 520.650 604.050 527.850 ;
        RECT 607.950 526.950 610.050 529.050 ;
        RECT 616.950 527.850 619.050 529.950 ;
        RECT 625.950 527.850 628.050 529.950 ;
        RECT 629.400 528.150 630.600 536.400 ;
        RECT 641.550 534.300 643.350 539.250 ;
        RECT 644.550 535.200 646.350 539.250 ;
        RECT 647.550 534.300 649.350 539.250 ;
        RECT 641.550 532.950 649.350 534.300 ;
        RECT 650.550 533.400 652.350 539.250 ;
        RECT 656.550 536.400 658.350 539.250 ;
        RECT 659.550 536.400 661.350 539.250 ;
        RECT 662.550 536.400 664.350 539.250 ;
        RECT 650.550 531.300 651.750 533.400 ;
        RECT 648.000 530.250 651.750 531.300 ;
        RECT 644.100 528.150 645.900 529.950 ;
        RECT 604.950 524.850 607.050 526.950 ;
        RECT 613.950 524.850 616.050 526.950 ;
        RECT 605.100 523.050 606.900 524.850 ;
        RECT 614.100 523.050 615.900 524.850 ;
        RECT 618.000 520.650 619.050 527.850 ;
        RECT 619.950 524.850 622.050 526.950 ;
        RECT 626.100 526.050 627.900 527.850 ;
        RECT 628.950 526.050 631.050 528.150 ;
        RECT 620.100 523.050 621.900 524.850 ;
        RECT 603.000 519.600 605.550 520.650 ;
        RECT 618.000 519.600 620.550 520.650 ;
        RECT 554.550 507.750 562.350 508.500 ;
        RECT 572.550 507.750 574.350 513.600 ;
        RECT 575.550 507.750 577.350 513.600 ;
        RECT 586.650 507.750 588.450 513.600 ;
        RECT 589.650 507.750 591.450 513.600 ;
        RECT 592.650 507.750 594.450 513.600 ;
        RECT 599.550 507.750 601.350 519.600 ;
        RECT 603.750 507.750 605.550 519.600 ;
        RECT 614.550 507.750 616.350 519.600 ;
        RECT 618.750 507.750 620.550 519.600 ;
        RECT 629.400 513.600 630.600 526.050 ;
        RECT 640.950 524.850 643.050 526.950 ;
        RECT 643.950 526.050 646.050 528.150 ;
        RECT 647.850 526.950 649.050 530.250 ;
        RECT 660.000 529.950 661.050 536.400 ;
        RECT 674.850 532.200 676.650 539.250 ;
        RECT 679.350 533.400 681.150 539.250 ;
        RECT 684.750 536.400 686.550 539.250 ;
        RECT 687.750 536.400 689.550 539.250 ;
        RECT 674.850 531.300 678.450 532.200 ;
        RECT 658.950 527.850 661.050 529.950 ;
        RECT 646.950 524.850 649.050 526.950 ;
        RECT 655.950 524.850 658.050 526.950 ;
        RECT 641.100 523.050 642.900 524.850 ;
        RECT 646.950 519.600 648.150 524.850 ;
        RECT 649.950 521.850 652.050 523.950 ;
        RECT 656.100 523.050 657.900 524.850 ;
        RECT 649.950 520.050 651.750 521.850 ;
        RECT 660.000 520.650 661.050 527.850 ;
        RECT 661.950 524.850 664.050 526.950 ;
        RECT 674.100 525.150 675.900 526.950 ;
        RECT 662.100 523.050 663.900 524.850 ;
        RECT 673.950 523.050 676.050 525.150 ;
        RECT 677.250 523.950 678.450 531.300 ;
        RECT 688.050 528.150 689.550 536.400 ;
        RECT 680.100 525.150 681.900 526.950 ;
        RECT 685.950 526.050 689.550 528.150 ;
        RECT 676.950 521.850 679.050 523.950 ;
        RECT 679.950 523.050 682.050 525.150 ;
        RECT 660.000 519.600 662.550 520.650 ;
        RECT 626.550 507.750 628.350 513.600 ;
        RECT 629.550 507.750 631.350 513.600 ;
        RECT 642.300 507.750 644.100 519.600 ;
        RECT 646.500 507.750 648.300 519.600 ;
        RECT 649.800 507.750 651.600 513.600 ;
        RECT 656.550 507.750 658.350 519.600 ;
        RECT 660.750 507.750 662.550 519.600 ;
        RECT 677.250 513.600 678.450 521.850 ;
        RECT 688.050 513.600 689.550 526.050 ;
        RECT 691.650 533.400 693.450 539.250 ;
        RECT 697.050 533.400 698.850 539.250 ;
        RECT 702.600 534.600 704.400 539.250 ;
        RECT 707.250 535.500 709.050 539.250 ;
        RECT 710.250 535.500 712.050 539.250 ;
        RECT 713.250 535.500 715.050 539.250 ;
        RECT 700.200 533.400 704.400 534.600 ;
        RECT 706.950 533.400 709.050 535.500 ;
        RECT 709.950 533.400 712.050 535.500 ;
        RECT 712.950 533.400 715.050 535.500 ;
        RECT 717.000 535.500 718.800 539.250 ;
        RECT 720.000 536.400 721.800 539.250 ;
        RECT 723.000 535.500 724.800 539.250 ;
        RECT 727.500 536.400 729.300 539.250 ;
        RECT 730.500 536.400 732.300 539.250 ;
        RECT 733.500 536.400 735.300 539.250 ;
        RECT 736.500 536.400 738.300 539.250 ;
        RECT 717.000 533.700 719.850 535.500 ;
        RECT 717.750 533.400 719.850 533.700 ;
        RECT 721.950 533.700 724.800 535.500 ;
        RECT 725.700 534.750 727.500 535.200 ;
        RECT 730.950 535.050 732.300 536.400 ;
        RECT 733.950 535.050 735.300 536.400 ;
        RECT 736.950 535.050 738.300 536.400 ;
        RECT 721.950 533.400 724.050 533.700 ;
        RECT 725.700 533.400 729.750 534.750 ;
        RECT 691.650 518.550 692.850 533.400 ;
        RECT 700.200 529.800 701.700 533.400 ;
        RECT 706.350 530.700 713.100 532.500 ;
        RECT 714.000 530.700 720.900 532.500 ;
        RECT 728.850 532.050 729.750 533.400 ;
        RECT 730.950 532.950 733.050 535.050 ;
        RECT 733.950 532.950 736.050 535.050 ;
        RECT 736.950 532.950 739.050 535.050 ;
        RECT 728.850 531.900 733.950 532.050 ;
        RECT 728.850 531.150 736.500 531.900 ;
        RECT 732.150 530.700 736.500 531.150 ;
        RECT 714.000 529.800 715.050 530.700 ;
        RECT 732.150 530.250 733.950 530.700 ;
        RECT 693.900 528.000 701.700 529.800 ;
        RECT 705.150 528.750 715.050 529.800 ;
        RECT 705.150 526.950 706.200 528.750 ;
        RECT 715.950 528.450 723.600 529.800 ;
        RECT 715.950 527.700 716.850 528.450 ;
        RECT 697.950 525.900 706.200 526.950 ;
        RECT 707.250 526.650 716.850 527.700 ;
        RECT 697.950 521.850 700.050 525.900 ;
        RECT 707.250 525.000 708.150 526.650 ;
        RECT 717.750 525.750 721.650 527.550 ;
        RECT 722.550 526.950 723.600 528.450 ;
        RECT 724.950 529.650 727.050 529.950 ;
        RECT 724.950 527.850 728.850 529.650 ;
        RECT 735.450 527.250 736.500 530.700 ;
        RECT 738.000 529.800 739.050 532.950 ;
        RECT 740.700 533.400 742.500 539.250 ;
        RECT 746.100 533.400 747.900 539.250 ;
        RECT 751.500 533.400 753.300 539.250 ;
        RECT 740.700 532.500 742.200 533.400 ;
        RECT 740.700 531.300 749.100 532.500 ;
        RECT 747.300 530.700 749.100 531.300 ;
        RECT 752.100 529.800 753.300 533.400 ;
        RECT 758.550 534.300 760.350 539.250 ;
        RECT 761.550 535.200 763.350 539.250 ;
        RECT 764.550 534.300 766.350 539.250 ;
        RECT 758.550 532.950 766.350 534.300 ;
        RECT 767.550 533.400 769.350 539.250 ;
        RECT 776.850 533.400 778.650 539.250 ;
        RECT 757.950 531.450 760.050 532.050 ;
        RECT 738.000 528.900 753.300 529.800 ;
        RECT 722.550 526.050 734.550 526.950 ;
        RECT 701.100 523.200 708.150 525.000 ;
        RECT 709.500 523.950 711.300 525.750 ;
        RECT 717.750 525.450 719.850 525.750 ;
        RECT 721.950 524.550 724.050 524.850 ;
        RECT 730.800 524.550 732.600 525.150 ;
        RECT 721.950 523.950 732.600 524.550 ;
        RECT 709.500 523.350 732.600 523.950 ;
        RECT 733.500 524.550 734.550 526.050 ;
        RECT 735.450 525.450 737.250 527.250 ;
        RECT 739.050 526.950 750.900 528.000 ;
        RECT 739.050 524.550 740.250 526.950 ;
        RECT 749.100 525.150 750.900 526.950 ;
        RECT 733.500 523.650 740.250 524.550 ;
        RECT 742.950 523.650 745.050 523.950 ;
        RECT 709.500 522.750 724.050 523.350 ;
        RECT 741.150 522.450 745.050 523.650 ;
        RECT 748.950 523.050 751.050 525.150 ;
        RECT 731.100 521.850 745.050 522.450 ;
        RECT 705.000 521.550 744.750 521.850 ;
        RECT 693.750 520.650 695.550 521.250 ;
        RECT 705.000 520.650 733.050 521.550 ;
        RECT 693.750 519.450 706.050 520.650 ;
        RECT 733.950 520.050 736.050 520.350 ;
        RECT 743.700 520.050 745.500 520.650 ;
        RECT 706.950 518.550 709.050 519.750 ;
        RECT 691.650 517.650 709.050 518.550 ;
        RECT 712.950 518.400 733.050 519.750 ;
        RECT 712.950 517.650 715.050 518.400 ;
        RECT 694.500 513.600 695.700 517.650 ;
        RECT 696.600 515.700 698.400 516.300 ;
        RECT 703.350 516.150 705.150 516.300 ;
        RECT 696.600 514.500 702.300 515.700 ;
        RECT 703.350 514.950 712.050 516.150 ;
        RECT 703.350 514.500 705.150 514.950 ;
        RECT 673.650 507.750 675.450 513.600 ;
        RECT 676.650 507.750 678.450 513.600 ;
        RECT 679.650 507.750 681.450 513.600 ;
        RECT 684.750 507.750 686.550 513.600 ;
        RECT 687.750 507.750 689.550 513.600 ;
        RECT 691.500 507.750 693.300 513.600 ;
        RECT 694.500 507.750 696.300 513.600 ;
        RECT 697.500 507.750 699.300 513.600 ;
        RECT 700.500 507.750 702.300 514.500 ;
        RECT 709.950 514.050 712.050 514.950 ;
        RECT 703.500 507.750 705.300 513.600 ;
        RECT 706.800 511.800 708.900 513.900 ;
        RECT 707.400 510.600 708.900 511.800 ;
        RECT 707.250 507.750 709.050 510.600 ;
        RECT 710.250 507.750 712.050 514.050 ;
        RECT 713.550 510.600 714.900 517.650 ;
        RECT 731.100 517.350 733.050 518.400 ;
        RECT 733.950 518.850 745.500 520.050 ;
        RECT 733.950 518.250 736.050 518.850 ;
        RECT 747.000 517.350 748.800 518.100 ;
        RECT 716.100 514.800 720.000 516.600 ;
        RECT 717.000 514.500 720.000 514.800 ;
        RECT 721.950 516.150 724.050 516.600 ;
        RECT 731.100 516.300 748.800 517.350 ;
        RECT 721.950 514.500 724.350 516.150 ;
        RECT 713.250 507.750 715.050 510.600 ;
        RECT 717.000 507.750 718.800 514.500 ;
        RECT 723.000 513.600 724.350 514.500 ;
        RECT 730.950 513.600 733.050 514.050 ;
        RECT 720.000 507.750 721.800 513.600 ;
        RECT 723.000 507.750 724.800 513.600 ;
        RECT 726.750 507.750 728.550 513.600 ;
        RECT 730.500 511.950 733.050 513.600 ;
        RECT 733.950 511.950 736.050 514.050 ;
        RECT 736.950 511.950 739.050 514.050 ;
        RECT 730.500 510.600 731.700 511.950 ;
        RECT 733.950 510.600 734.850 511.950 ;
        RECT 736.950 510.600 738.150 511.950 ;
        RECT 729.750 507.750 731.700 510.600 ;
        RECT 732.750 507.750 734.850 510.600 ;
        RECT 735.750 507.750 738.150 510.600 ;
        RECT 739.500 507.750 741.300 511.050 ;
        RECT 742.500 507.750 744.300 516.300 ;
        RECT 752.100 515.400 753.300 528.900 ;
        RECT 755.550 530.550 760.050 531.450 ;
        RECT 767.550 531.300 768.750 533.400 ;
        RECT 781.350 532.200 783.150 539.250 ;
        RECT 789.750 536.400 791.550 539.250 ;
        RECT 792.750 536.400 794.550 539.250 ;
        RECT 755.550 520.050 756.450 530.550 ;
        RECT 757.950 529.950 760.050 530.550 ;
        RECT 765.000 530.250 768.750 531.300 ;
        RECT 779.550 531.300 783.150 532.200 ;
        RECT 761.100 528.150 762.900 529.950 ;
        RECT 757.950 524.850 760.050 526.950 ;
        RECT 760.950 526.050 763.050 528.150 ;
        RECT 764.850 526.950 766.050 530.250 ;
        RECT 763.950 524.850 766.050 526.950 ;
        RECT 776.100 525.150 777.900 526.950 ;
        RECT 758.100 523.050 759.900 524.850 ;
        RECT 754.950 517.950 757.050 520.050 ;
        RECT 763.950 519.600 765.150 524.850 ;
        RECT 766.950 521.850 769.050 523.950 ;
        RECT 775.950 523.050 778.050 525.150 ;
        RECT 779.550 523.950 780.750 531.300 ;
        RECT 793.050 528.150 794.550 536.400 ;
        RECT 782.100 525.150 783.900 526.950 ;
        RECT 790.950 526.050 794.550 528.150 ;
        RECT 778.950 521.850 781.050 523.950 ;
        RECT 781.950 523.050 784.050 525.150 ;
        RECT 766.950 520.050 768.750 521.850 ;
        RECT 749.250 514.500 753.300 515.400 ;
        RECT 749.250 513.600 750.300 514.500 ;
        RECT 745.500 507.750 747.300 513.600 ;
        RECT 748.500 507.750 750.300 513.600 ;
        RECT 751.500 507.750 753.300 513.600 ;
        RECT 759.300 507.750 761.100 519.600 ;
        RECT 763.500 507.750 765.300 519.600 ;
        RECT 779.550 513.600 780.750 521.850 ;
        RECT 793.050 513.600 794.550 526.050 ;
        RECT 796.650 533.400 798.450 539.250 ;
        RECT 802.050 533.400 803.850 539.250 ;
        RECT 807.600 534.600 809.400 539.250 ;
        RECT 812.250 535.500 814.050 539.250 ;
        RECT 815.250 535.500 817.050 539.250 ;
        RECT 818.250 535.500 820.050 539.250 ;
        RECT 805.200 533.400 809.400 534.600 ;
        RECT 811.950 533.400 814.050 535.500 ;
        RECT 814.950 533.400 817.050 535.500 ;
        RECT 817.950 533.400 820.050 535.500 ;
        RECT 822.000 535.500 823.800 539.250 ;
        RECT 825.000 536.400 826.800 539.250 ;
        RECT 828.000 535.500 829.800 539.250 ;
        RECT 832.500 536.400 834.300 539.250 ;
        RECT 835.500 536.400 837.300 539.250 ;
        RECT 838.500 536.400 840.300 539.250 ;
        RECT 841.500 536.400 843.300 539.250 ;
        RECT 822.000 533.700 824.850 535.500 ;
        RECT 822.750 533.400 824.850 533.700 ;
        RECT 826.950 533.700 829.800 535.500 ;
        RECT 830.700 534.750 832.500 535.200 ;
        RECT 835.950 535.050 837.300 536.400 ;
        RECT 838.950 535.050 840.300 536.400 ;
        RECT 841.950 535.050 843.300 536.400 ;
        RECT 826.950 533.400 829.050 533.700 ;
        RECT 830.700 533.400 834.750 534.750 ;
        RECT 796.650 518.550 797.850 533.400 ;
        RECT 805.200 529.800 806.700 533.400 ;
        RECT 811.350 530.700 818.100 532.500 ;
        RECT 819.000 530.700 825.900 532.500 ;
        RECT 833.850 532.050 834.750 533.400 ;
        RECT 835.950 532.950 838.050 535.050 ;
        RECT 838.950 532.950 841.050 535.050 ;
        RECT 841.950 532.950 844.050 535.050 ;
        RECT 833.850 531.900 838.950 532.050 ;
        RECT 833.850 531.150 841.500 531.900 ;
        RECT 837.150 530.700 841.500 531.150 ;
        RECT 819.000 529.800 820.050 530.700 ;
        RECT 837.150 530.250 838.950 530.700 ;
        RECT 798.900 528.000 806.700 529.800 ;
        RECT 810.150 528.750 820.050 529.800 ;
        RECT 810.150 526.950 811.200 528.750 ;
        RECT 820.950 528.450 828.600 529.800 ;
        RECT 820.950 527.700 821.850 528.450 ;
        RECT 802.950 525.900 811.200 526.950 ;
        RECT 812.250 526.650 821.850 527.700 ;
        RECT 802.950 521.850 805.050 525.900 ;
        RECT 812.250 525.000 813.150 526.650 ;
        RECT 822.750 525.750 826.650 527.550 ;
        RECT 827.550 526.950 828.600 528.450 ;
        RECT 829.950 529.650 832.050 529.950 ;
        RECT 829.950 527.850 833.850 529.650 ;
        RECT 840.450 527.250 841.500 530.700 ;
        RECT 843.000 529.800 844.050 532.950 ;
        RECT 845.700 533.400 847.500 539.250 ;
        RECT 851.100 533.400 852.900 539.250 ;
        RECT 856.500 533.400 858.300 539.250 ;
        RECT 845.700 532.500 847.200 533.400 ;
        RECT 845.700 531.300 854.100 532.500 ;
        RECT 852.300 530.700 854.100 531.300 ;
        RECT 857.100 529.800 858.300 533.400 ;
        RECT 843.000 528.900 858.300 529.800 ;
        RECT 827.550 526.050 839.550 526.950 ;
        RECT 806.100 523.200 813.150 525.000 ;
        RECT 814.500 523.950 816.300 525.750 ;
        RECT 822.750 525.450 824.850 525.750 ;
        RECT 826.950 524.550 829.050 524.850 ;
        RECT 835.800 524.550 837.600 525.150 ;
        RECT 826.950 523.950 837.600 524.550 ;
        RECT 814.500 523.350 837.600 523.950 ;
        RECT 838.500 524.550 839.550 526.050 ;
        RECT 840.450 525.450 842.250 527.250 ;
        RECT 844.050 526.950 855.900 528.000 ;
        RECT 844.050 524.550 845.250 526.950 ;
        RECT 854.100 525.150 855.900 526.950 ;
        RECT 838.500 523.650 845.250 524.550 ;
        RECT 847.950 523.650 850.050 523.950 ;
        RECT 814.500 522.750 829.050 523.350 ;
        RECT 846.150 522.450 850.050 523.650 ;
        RECT 853.950 523.050 856.050 525.150 ;
        RECT 836.100 521.850 850.050 522.450 ;
        RECT 810.000 521.550 849.750 521.850 ;
        RECT 798.750 520.650 800.550 521.250 ;
        RECT 810.000 520.650 838.050 521.550 ;
        RECT 798.750 519.450 811.050 520.650 ;
        RECT 838.950 520.050 841.050 520.350 ;
        RECT 848.700 520.050 850.500 520.650 ;
        RECT 811.950 518.550 814.050 519.750 ;
        RECT 796.650 517.650 814.050 518.550 ;
        RECT 817.950 518.400 838.050 519.750 ;
        RECT 817.950 517.650 820.050 518.400 ;
        RECT 799.500 513.600 800.700 517.650 ;
        RECT 801.600 515.700 803.400 516.300 ;
        RECT 808.350 516.150 810.150 516.300 ;
        RECT 801.600 514.500 807.300 515.700 ;
        RECT 808.350 514.950 817.050 516.150 ;
        RECT 808.350 514.500 810.150 514.950 ;
        RECT 766.800 507.750 768.600 513.600 ;
        RECT 776.550 507.750 778.350 513.600 ;
        RECT 779.550 507.750 781.350 513.600 ;
        RECT 782.550 507.750 784.350 513.600 ;
        RECT 789.750 507.750 791.550 513.600 ;
        RECT 792.750 507.750 794.550 513.600 ;
        RECT 796.500 507.750 798.300 513.600 ;
        RECT 799.500 507.750 801.300 513.600 ;
        RECT 802.500 507.750 804.300 513.600 ;
        RECT 805.500 507.750 807.300 514.500 ;
        RECT 814.950 514.050 817.050 514.950 ;
        RECT 808.500 507.750 810.300 513.600 ;
        RECT 811.800 511.800 813.900 513.900 ;
        RECT 812.400 510.600 813.900 511.800 ;
        RECT 812.250 507.750 814.050 510.600 ;
        RECT 815.250 507.750 817.050 514.050 ;
        RECT 818.550 510.600 819.900 517.650 ;
        RECT 836.100 517.350 838.050 518.400 ;
        RECT 838.950 518.850 850.500 520.050 ;
        RECT 838.950 518.250 841.050 518.850 ;
        RECT 852.000 517.350 853.800 518.100 ;
        RECT 821.100 514.800 825.000 516.600 ;
        RECT 822.000 514.500 825.000 514.800 ;
        RECT 826.950 516.150 829.050 516.600 ;
        RECT 836.100 516.300 853.800 517.350 ;
        RECT 826.950 514.500 829.350 516.150 ;
        RECT 818.250 507.750 820.050 510.600 ;
        RECT 822.000 507.750 823.800 514.500 ;
        RECT 828.000 513.600 829.350 514.500 ;
        RECT 835.950 513.600 838.050 514.050 ;
        RECT 825.000 507.750 826.800 513.600 ;
        RECT 828.000 507.750 829.800 513.600 ;
        RECT 831.750 507.750 833.550 513.600 ;
        RECT 835.500 511.950 838.050 513.600 ;
        RECT 838.950 511.950 841.050 514.050 ;
        RECT 841.950 511.950 844.050 514.050 ;
        RECT 835.500 510.600 836.700 511.950 ;
        RECT 838.950 510.600 839.850 511.950 ;
        RECT 841.950 510.600 843.150 511.950 ;
        RECT 834.750 507.750 836.700 510.600 ;
        RECT 837.750 507.750 839.850 510.600 ;
        RECT 840.750 507.750 843.150 510.600 ;
        RECT 844.500 507.750 846.300 511.050 ;
        RECT 847.500 507.750 849.300 516.300 ;
        RECT 857.100 515.400 858.300 528.900 ;
        RECT 854.250 514.500 858.300 515.400 ;
        RECT 854.250 513.600 855.300 514.500 ;
        RECT 850.500 507.750 852.300 513.600 ;
        RECT 853.500 507.750 855.300 513.600 ;
        RECT 856.500 507.750 858.300 513.600 ;
        RECT 7.650 497.400 9.450 503.250 ;
        RECT 10.650 497.400 12.450 503.250 ;
        RECT 8.400 484.950 9.600 497.400 ;
        RECT 17.550 491.400 19.350 503.250 ;
        RECT 22.050 491.550 23.850 503.250 ;
        RECT 25.050 492.900 26.850 503.250 ;
        RECT 38.400 497.400 40.200 503.250 ;
        RECT 25.050 491.550 27.450 492.900 ;
        RECT 17.550 490.200 18.750 491.400 ;
        RECT 22.950 490.200 24.750 490.650 ;
        RECT 17.550 489.000 24.750 490.200 ;
        RECT 22.950 488.850 24.750 489.000 ;
        RECT 20.100 486.150 21.900 487.950 ;
        RECT 7.950 482.850 10.050 484.950 ;
        RECT 11.100 483.150 12.900 484.950 ;
        RECT 17.100 483.150 18.900 484.950 ;
        RECT 19.950 484.050 22.050 486.150 ;
        RECT 8.400 474.600 9.600 482.850 ;
        RECT 10.950 481.050 13.050 483.150 ;
        RECT 16.950 481.050 19.050 483.150 ;
        RECT 23.700 480.600 24.600 488.850 ;
        RECT 26.100 484.950 27.450 491.550 ;
        RECT 41.700 491.400 43.500 503.250 ;
        RECT 45.900 491.400 47.700 503.250 ;
        RECT 54.300 491.400 56.100 503.250 ;
        RECT 58.500 491.400 60.300 503.250 ;
        RECT 61.800 497.400 63.600 503.250 ;
        RECT 71.550 491.400 73.350 503.250 ;
        RECT 76.050 491.550 77.850 503.250 ;
        RECT 79.050 492.900 80.850 503.250 ;
        RECT 89.550 497.400 91.350 503.250 ;
        RECT 92.550 497.400 94.350 503.250 ;
        RECT 95.550 498.000 97.350 503.250 ;
        RECT 92.700 497.100 94.350 497.400 ;
        RECT 98.550 497.400 100.350 503.250 ;
        RECT 98.550 497.100 99.750 497.400 ;
        RECT 92.700 496.200 99.750 497.100 ;
        RECT 79.050 491.550 81.450 492.900 ;
        RECT 92.100 492.150 93.900 493.950 ;
        RECT 38.250 489.150 40.050 490.950 ;
        RECT 37.950 487.050 40.050 489.150 ;
        RECT 41.850 486.150 43.050 491.400 ;
        RECT 47.100 486.150 48.900 487.950 ;
        RECT 53.100 486.150 54.900 487.950 ;
        RECT 58.950 486.150 60.150 491.400 ;
        RECT 61.950 489.150 63.750 490.950 ;
        RECT 71.550 490.200 72.750 491.400 ;
        RECT 76.950 490.200 78.750 490.650 ;
        RECT 61.950 487.050 64.050 489.150 ;
        RECT 71.550 489.000 78.750 490.200 ;
        RECT 76.950 488.850 78.750 489.000 ;
        RECT 74.100 486.150 75.900 487.950 ;
        RECT 25.950 482.850 28.050 484.950 ;
        RECT 22.950 479.700 24.750 480.600 ;
        RECT 21.450 478.800 24.750 479.700 ;
        RECT 21.450 474.600 22.350 478.800 ;
        RECT 27.000 477.600 28.050 482.850 ;
        RECT 40.950 484.050 43.050 486.150 ;
        RECT 40.950 480.750 42.150 484.050 ;
        RECT 43.950 482.850 46.050 484.950 ;
        RECT 46.950 484.050 49.050 486.150 ;
        RECT 52.950 484.050 55.050 486.150 ;
        RECT 55.950 482.850 58.050 484.950 ;
        RECT 58.950 484.050 61.050 486.150 ;
        RECT 44.100 481.050 45.900 482.850 ;
        RECT 56.100 481.050 57.900 482.850 ;
        RECT 59.850 480.750 61.050 484.050 ;
        RECT 71.100 483.150 72.900 484.950 ;
        RECT 73.950 484.050 76.050 486.150 ;
        RECT 70.950 481.050 73.050 483.150 ;
        RECT 38.250 479.700 42.000 480.750 ;
        RECT 60.000 479.700 63.750 480.750 ;
        RECT 77.700 480.600 78.600 488.850 ;
        RECT 80.100 484.950 81.450 491.550 ;
        RECT 89.100 489.150 90.900 490.950 ;
        RECT 91.950 490.050 94.050 492.150 ;
        RECT 95.250 489.150 97.050 490.950 ;
        RECT 88.950 487.050 91.050 489.150 ;
        RECT 94.950 487.050 97.050 489.150 ;
        RECT 98.700 487.950 99.750 496.200 ;
        RECT 108.300 491.400 110.100 503.250 ;
        RECT 112.500 491.400 114.300 503.250 ;
        RECT 115.800 497.400 117.600 503.250 ;
        RECT 122.700 497.400 124.500 503.250 ;
        RECT 125.700 497.400 127.500 503.250 ;
        RECT 128.700 497.400 130.500 503.250 ;
        RECT 125.700 496.500 126.750 497.400 ;
        RECT 122.700 495.600 126.750 496.500 ;
        RECT 97.950 485.850 100.050 487.950 ;
        RECT 107.100 486.150 108.900 487.950 ;
        RECT 112.950 486.150 114.150 491.400 ;
        RECT 115.950 489.150 117.750 490.950 ;
        RECT 115.950 487.050 118.050 489.150 ;
        RECT 79.950 482.850 82.050 484.950 ;
        RECT 76.950 479.700 78.750 480.600 ;
        RECT 38.250 477.600 39.450 479.700 ;
        RECT 7.650 471.750 9.450 474.600 ;
        RECT 10.650 471.750 12.450 474.600 ;
        RECT 17.550 471.750 19.350 474.600 ;
        RECT 20.550 471.750 22.350 474.600 ;
        RECT 23.550 471.750 25.350 474.600 ;
        RECT 26.550 471.750 28.350 477.600 ;
        RECT 37.650 471.750 39.450 477.600 ;
        RECT 40.650 476.700 48.450 478.050 ;
        RECT 40.650 471.750 42.450 476.700 ;
        RECT 43.650 471.750 45.450 475.800 ;
        RECT 46.650 471.750 48.450 476.700 ;
        RECT 53.550 476.700 61.350 478.050 ;
        RECT 53.550 471.750 55.350 476.700 ;
        RECT 56.550 471.750 58.350 475.800 ;
        RECT 59.550 471.750 61.350 476.700 ;
        RECT 62.550 477.600 63.750 479.700 ;
        RECT 75.450 478.800 78.750 479.700 ;
        RECT 62.550 471.750 64.350 477.600 ;
        RECT 75.450 474.600 76.350 478.800 ;
        RECT 81.000 477.600 82.050 482.850 ;
        RECT 82.950 483.450 85.050 484.050 ;
        RECT 88.950 483.450 91.050 484.050 ;
        RECT 82.950 482.550 91.050 483.450 ;
        RECT 82.950 481.950 85.050 482.550 ;
        RECT 88.950 481.950 91.050 482.550 ;
        RECT 98.400 481.650 99.600 485.850 ;
        RECT 106.950 484.050 109.050 486.150 ;
        RECT 109.950 482.850 112.050 484.950 ;
        RECT 112.950 484.050 115.050 486.150 ;
        RECT 71.550 471.750 73.350 474.600 ;
        RECT 74.550 471.750 76.350 474.600 ;
        RECT 77.550 471.750 79.350 474.600 ;
        RECT 80.550 471.750 82.350 477.600 ;
        RECT 89.700 471.750 91.500 480.600 ;
        RECT 95.100 480.000 99.600 481.650 ;
        RECT 110.100 481.050 111.900 482.850 ;
        RECT 113.850 480.750 115.050 484.050 ;
        RECT 122.700 482.100 123.900 495.600 ;
        RECT 131.700 494.700 133.500 503.250 ;
        RECT 134.700 499.950 136.500 503.250 ;
        RECT 137.850 500.400 140.250 503.250 ;
        RECT 141.150 500.400 143.250 503.250 ;
        RECT 144.300 500.400 146.250 503.250 ;
        RECT 137.850 499.050 139.050 500.400 ;
        RECT 141.150 499.050 142.050 500.400 ;
        RECT 144.300 499.050 145.500 500.400 ;
        RECT 136.950 496.950 139.050 499.050 ;
        RECT 139.950 496.950 142.050 499.050 ;
        RECT 142.950 497.400 145.500 499.050 ;
        RECT 147.450 497.400 149.250 503.250 ;
        RECT 151.200 497.400 153.000 503.250 ;
        RECT 154.200 497.400 156.000 503.250 ;
        RECT 142.950 496.950 145.050 497.400 ;
        RECT 151.650 496.500 153.000 497.400 ;
        RECT 157.200 496.500 159.000 503.250 ;
        RECT 160.950 500.400 162.750 503.250 ;
        RECT 151.650 494.850 154.050 496.500 ;
        RECT 127.200 493.650 144.900 494.700 ;
        RECT 151.950 494.400 154.050 494.850 ;
        RECT 156.000 496.200 159.000 496.500 ;
        RECT 156.000 494.400 159.900 496.200 ;
        RECT 127.200 492.900 129.000 493.650 ;
        RECT 139.950 492.150 142.050 492.750 ;
        RECT 130.500 490.950 142.050 492.150 ;
        RECT 142.950 492.600 144.900 493.650 ;
        RECT 161.100 493.350 162.450 500.400 ;
        RECT 163.950 496.950 165.750 503.250 ;
        RECT 166.950 500.400 168.750 503.250 ;
        RECT 167.100 499.200 168.600 500.400 ;
        RECT 167.100 497.100 169.200 499.200 ;
        RECT 170.700 497.400 172.500 503.250 ;
        RECT 163.950 496.050 166.050 496.950 ;
        RECT 173.700 496.500 175.500 503.250 ;
        RECT 176.700 497.400 178.500 503.250 ;
        RECT 179.700 497.400 181.500 503.250 ;
        RECT 182.700 497.400 184.500 503.250 ;
        RECT 186.450 497.400 188.250 503.250 ;
        RECT 189.450 497.400 191.250 503.250 ;
        RECT 197.550 497.400 199.350 503.250 ;
        RECT 200.550 497.400 202.350 503.250 ;
        RECT 203.550 498.000 205.350 503.250 ;
        RECT 170.850 496.050 172.650 496.500 ;
        RECT 163.950 494.850 172.650 496.050 ;
        RECT 173.700 495.300 179.400 496.500 ;
        RECT 170.850 494.700 172.650 494.850 ;
        RECT 177.600 494.700 179.400 495.300 ;
        RECT 180.300 493.350 181.500 497.400 ;
        RECT 160.950 492.600 163.050 493.350 ;
        RECT 142.950 491.250 163.050 492.600 ;
        RECT 166.950 492.450 184.350 493.350 ;
        RECT 166.950 491.250 169.050 492.450 ;
        RECT 130.500 490.350 132.300 490.950 ;
        RECT 139.950 490.650 142.050 490.950 ;
        RECT 169.950 490.350 182.250 491.550 ;
        RECT 142.950 489.450 171.000 490.350 ;
        RECT 180.450 489.750 182.250 490.350 ;
        RECT 131.250 489.150 171.000 489.450 ;
        RECT 130.950 488.550 144.900 489.150 ;
        RECT 124.950 485.850 127.050 487.950 ;
        RECT 130.950 487.350 134.850 488.550 ;
        RECT 151.950 487.650 166.500 488.250 ;
        RECT 130.950 487.050 133.050 487.350 ;
        RECT 135.750 486.450 142.500 487.350 ;
        RECT 125.100 484.050 126.900 485.850 ;
        RECT 135.750 484.050 136.950 486.450 ;
        RECT 125.100 483.000 136.950 484.050 ;
        RECT 138.750 483.750 140.550 485.550 ;
        RECT 141.450 484.950 142.500 486.450 ;
        RECT 143.400 487.050 166.500 487.650 ;
        RECT 143.400 486.450 154.050 487.050 ;
        RECT 143.400 485.850 145.200 486.450 ;
        RECT 151.950 486.150 154.050 486.450 ;
        RECT 156.150 485.250 158.250 485.550 ;
        RECT 164.700 485.250 166.500 487.050 ;
        RECT 167.850 486.000 174.900 487.800 ;
        RECT 141.450 484.050 153.450 484.950 ;
        RECT 122.700 481.200 138.000 482.100 ;
        RECT 95.100 471.750 96.900 480.000 ;
        RECT 114.000 479.700 117.750 480.750 ;
        RECT 107.550 476.700 115.350 478.050 ;
        RECT 107.550 471.750 109.350 476.700 ;
        RECT 110.550 471.750 112.350 475.800 ;
        RECT 113.550 471.750 115.350 476.700 ;
        RECT 116.550 477.600 117.750 479.700 ;
        RECT 122.700 477.600 123.900 481.200 ;
        RECT 126.900 479.700 128.700 480.300 ;
        RECT 126.900 478.500 135.300 479.700 ;
        RECT 133.800 477.600 135.300 478.500 ;
        RECT 116.550 471.750 118.350 477.600 ;
        RECT 122.700 471.750 124.500 477.600 ;
        RECT 128.100 471.750 129.900 477.600 ;
        RECT 133.500 471.750 135.300 477.600 ;
        RECT 136.950 478.050 138.000 481.200 ;
        RECT 139.500 480.300 140.550 483.750 ;
        RECT 147.150 481.350 151.050 483.150 ;
        RECT 148.950 481.050 151.050 481.350 ;
        RECT 152.400 482.550 153.450 484.050 ;
        RECT 154.350 483.450 158.250 485.250 ;
        RECT 167.850 484.350 168.750 486.000 ;
        RECT 175.950 485.100 178.050 489.150 ;
        RECT 159.150 483.300 168.750 484.350 ;
        RECT 169.800 484.050 178.050 485.100 ;
        RECT 159.150 482.550 160.050 483.300 ;
        RECT 152.400 481.200 160.050 482.550 ;
        RECT 169.800 482.250 170.850 484.050 ;
        RECT 160.950 481.200 170.850 482.250 ;
        RECT 174.300 481.200 182.100 483.000 ;
        RECT 142.050 480.300 143.850 480.750 ;
        RECT 160.950 480.300 162.000 481.200 ;
        RECT 139.500 479.850 143.850 480.300 ;
        RECT 139.500 479.100 147.150 479.850 ;
        RECT 142.050 478.950 147.150 479.100 ;
        RECT 136.950 475.950 139.050 478.050 ;
        RECT 139.950 475.950 142.050 478.050 ;
        RECT 142.950 475.950 145.050 478.050 ;
        RECT 146.250 477.600 147.150 478.950 ;
        RECT 155.100 478.500 162.000 480.300 ;
        RECT 162.900 478.500 169.650 480.300 ;
        RECT 174.300 477.600 175.800 481.200 ;
        RECT 183.150 477.600 184.350 492.450 ;
        RECT 146.250 476.250 150.300 477.600 ;
        RECT 151.950 477.300 154.050 477.600 ;
        RECT 137.700 474.600 139.050 475.950 ;
        RECT 140.700 474.600 142.050 475.950 ;
        RECT 143.700 474.600 145.050 475.950 ;
        RECT 148.500 475.800 150.300 476.250 ;
        RECT 151.200 475.500 154.050 477.300 ;
        RECT 156.150 477.300 158.250 477.600 ;
        RECT 156.150 475.500 159.000 477.300 ;
        RECT 137.700 471.750 139.500 474.600 ;
        RECT 140.700 471.750 142.500 474.600 ;
        RECT 143.700 471.750 145.500 474.600 ;
        RECT 146.700 471.750 148.500 474.600 ;
        RECT 151.200 471.750 153.000 475.500 ;
        RECT 154.200 471.750 156.000 474.600 ;
        RECT 157.200 471.750 159.000 475.500 ;
        RECT 160.950 475.500 163.050 477.600 ;
        RECT 163.950 475.500 166.050 477.600 ;
        RECT 166.950 475.500 169.050 477.600 ;
        RECT 171.600 476.400 175.800 477.600 ;
        RECT 160.950 471.750 162.750 475.500 ;
        RECT 163.950 471.750 165.750 475.500 ;
        RECT 166.950 471.750 168.750 475.500 ;
        RECT 171.600 471.750 173.400 476.400 ;
        RECT 177.150 471.750 178.950 477.600 ;
        RECT 182.550 471.750 184.350 477.600 ;
        RECT 186.450 484.950 187.950 497.400 ;
        RECT 200.700 497.100 202.350 497.400 ;
        RECT 206.550 497.400 208.350 503.250 ;
        RECT 206.550 497.100 207.750 497.400 ;
        RECT 200.700 496.200 207.750 497.100 ;
        RECT 200.100 492.150 201.900 493.950 ;
        RECT 197.100 489.150 198.900 490.950 ;
        RECT 199.950 490.050 202.050 492.150 ;
        RECT 203.250 489.150 205.050 490.950 ;
        RECT 196.950 487.050 199.050 489.150 ;
        RECT 202.950 487.050 205.050 489.150 ;
        RECT 206.700 487.950 207.750 496.200 ;
        RECT 215.550 491.400 217.350 503.250 ;
        RECT 219.750 491.400 221.550 503.250 ;
        RECT 233.400 497.400 235.200 503.250 ;
        RECT 236.700 491.400 238.500 503.250 ;
        RECT 240.900 491.400 242.700 503.250 ;
        RECT 249.300 491.400 251.100 503.250 ;
        RECT 253.500 491.400 255.300 503.250 ;
        RECT 256.800 497.400 258.600 503.250 ;
        RECT 270.450 491.400 272.250 503.250 ;
        RECT 274.650 491.400 276.450 503.250 ;
        RECT 288.450 491.400 290.250 503.250 ;
        RECT 292.650 491.400 294.450 503.250 ;
        RECT 299.550 497.400 301.350 503.250 ;
        RECT 302.550 497.400 304.350 503.250 ;
        RECT 219.000 490.350 221.550 491.400 ;
        RECT 205.950 485.850 208.050 487.950 ;
        RECT 215.100 486.150 216.900 487.950 ;
        RECT 186.450 482.850 190.050 484.950 ;
        RECT 186.450 474.600 187.950 482.850 ;
        RECT 206.400 481.650 207.600 485.850 ;
        RECT 214.950 484.050 217.050 486.150 ;
        RECT 219.000 483.150 220.050 490.350 ;
        RECT 233.250 489.150 235.050 490.950 ;
        RECT 221.100 486.150 222.900 487.950 ;
        RECT 232.950 487.050 235.050 489.150 ;
        RECT 236.850 486.150 238.050 491.400 ;
        RECT 242.100 486.150 243.900 487.950 ;
        RECT 248.100 486.150 249.900 487.950 ;
        RECT 253.950 486.150 255.150 491.400 ;
        RECT 256.950 489.150 258.750 490.950 ;
        RECT 270.450 490.350 273.000 491.400 ;
        RECT 288.450 490.350 291.000 491.400 ;
        RECT 256.950 487.050 259.050 489.150 ;
        RECT 269.100 486.150 270.900 487.950 ;
        RECT 220.950 484.050 223.050 486.150 ;
        RECT 235.950 484.050 238.050 486.150 ;
        RECT 186.450 471.750 188.250 474.600 ;
        RECT 189.450 471.750 191.250 474.600 ;
        RECT 197.700 471.750 199.500 480.600 ;
        RECT 203.100 480.000 207.600 481.650 ;
        RECT 217.950 481.050 220.050 483.150 ;
        RECT 203.100 471.750 204.900 480.000 ;
        RECT 219.000 474.600 220.050 481.050 ;
        RECT 235.950 480.750 237.150 484.050 ;
        RECT 238.950 482.850 241.050 484.950 ;
        RECT 241.950 484.050 244.050 486.150 ;
        RECT 247.950 484.050 250.050 486.150 ;
        RECT 250.950 482.850 253.050 484.950 ;
        RECT 253.950 484.050 256.050 486.150 ;
        RECT 268.950 484.050 271.050 486.150 ;
        RECT 239.100 481.050 240.900 482.850 ;
        RECT 251.100 481.050 252.900 482.850 ;
        RECT 254.850 480.750 256.050 484.050 ;
        RECT 271.950 483.150 273.000 490.350 ;
        RECT 275.100 486.150 276.900 487.950 ;
        RECT 287.100 486.150 288.900 487.950 ;
        RECT 274.950 484.050 277.050 486.150 ;
        RECT 286.950 484.050 289.050 486.150 ;
        RECT 289.950 483.150 291.000 490.350 ;
        RECT 293.100 486.150 294.900 487.950 ;
        RECT 299.100 486.150 300.900 487.950 ;
        RECT 292.950 484.050 295.050 486.150 ;
        RECT 298.950 484.050 301.050 486.150 ;
        RECT 271.950 481.050 274.050 483.150 ;
        RECT 289.950 481.050 292.050 483.150 ;
        RECT 233.250 479.700 237.000 480.750 ;
        RECT 255.000 479.700 258.750 480.750 ;
        RECT 233.250 477.600 234.450 479.700 ;
        RECT 215.550 471.750 217.350 474.600 ;
        RECT 218.550 471.750 220.350 474.600 ;
        RECT 221.550 471.750 223.350 474.600 ;
        RECT 232.650 471.750 234.450 477.600 ;
        RECT 235.650 476.700 243.450 478.050 ;
        RECT 235.650 471.750 237.450 476.700 ;
        RECT 238.650 471.750 240.450 475.800 ;
        RECT 241.650 471.750 243.450 476.700 ;
        RECT 248.550 476.700 256.350 478.050 ;
        RECT 248.550 471.750 250.350 476.700 ;
        RECT 251.550 471.750 253.350 475.800 ;
        RECT 254.550 471.750 256.350 476.700 ;
        RECT 257.550 477.600 258.750 479.700 ;
        RECT 257.550 471.750 259.350 477.600 ;
        RECT 271.950 474.600 273.000 481.050 ;
        RECT 289.950 474.600 291.000 481.050 ;
        RECT 302.700 480.300 303.900 497.400 ;
        RECT 306.150 491.400 307.950 503.250 ;
        RECT 309.150 491.400 310.950 503.250 ;
        RECT 319.650 497.400 321.450 503.250 ;
        RECT 322.650 498.000 324.450 503.250 ;
        RECT 320.250 497.100 321.450 497.400 ;
        RECT 325.650 497.400 327.450 503.250 ;
        RECT 328.650 497.400 330.450 503.250 ;
        RECT 335.550 497.400 337.350 503.250 ;
        RECT 338.550 497.400 340.350 503.250 ;
        RECT 325.650 497.100 327.300 497.400 ;
        RECT 320.250 496.200 327.300 497.100 ;
        RECT 304.950 485.850 307.050 487.950 ;
        RECT 309.150 486.150 310.350 491.400 ;
        RECT 320.250 487.950 321.300 496.200 ;
        RECT 326.100 492.150 327.900 493.950 ;
        RECT 322.950 489.150 324.750 490.950 ;
        RECT 325.950 490.050 328.050 492.150 ;
        RECT 329.100 489.150 330.900 490.950 ;
        RECT 305.100 484.050 306.900 485.850 ;
        RECT 307.950 484.050 310.350 486.150 ;
        RECT 319.950 485.850 322.050 487.950 ;
        RECT 322.950 487.050 325.050 489.150 ;
        RECT 328.950 487.050 331.050 489.150 ;
        RECT 299.550 479.100 307.050 480.300 ;
        RECT 268.650 471.750 270.450 474.600 ;
        RECT 271.650 471.750 273.450 474.600 ;
        RECT 274.650 471.750 276.450 474.600 ;
        RECT 286.650 471.750 288.450 474.600 ;
        RECT 289.650 471.750 291.450 474.600 ;
        RECT 292.650 471.750 294.450 474.600 ;
        RECT 299.550 471.750 301.350 479.100 ;
        RECT 305.250 478.500 307.050 479.100 ;
        RECT 309.150 477.600 310.350 484.050 ;
        RECT 320.400 481.650 321.600 485.850 ;
        RECT 338.400 484.950 339.600 497.400 ;
        RECT 348.300 491.400 350.100 503.250 ;
        RECT 352.500 491.400 354.300 503.250 ;
        RECT 355.800 497.400 357.600 503.250 ;
        RECT 368.550 497.400 370.350 503.250 ;
        RECT 371.550 497.400 373.350 503.250 ;
        RECT 380.550 497.400 382.350 503.250 ;
        RECT 383.550 497.400 385.350 503.250 ;
        RECT 386.550 498.000 388.350 503.250 ;
        RECT 347.100 486.150 348.900 487.950 ;
        RECT 352.950 486.150 354.150 491.400 ;
        RECT 355.950 489.150 357.750 490.950 ;
        RECT 355.950 487.050 358.050 489.150 ;
        RECT 335.100 483.150 336.900 484.950 ;
        RECT 320.400 480.000 324.900 481.650 ;
        RECT 334.950 481.050 337.050 483.150 ;
        RECT 337.950 482.850 340.050 484.950 ;
        RECT 346.950 484.050 349.050 486.150 ;
        RECT 349.950 482.850 352.050 484.950 ;
        RECT 352.950 484.050 355.050 486.150 ;
        RECT 371.400 484.950 372.600 497.400 ;
        RECT 383.700 497.100 385.350 497.400 ;
        RECT 389.550 497.400 391.350 503.250 ;
        RECT 401.400 497.400 403.200 503.250 ;
        RECT 389.550 497.100 390.750 497.400 ;
        RECT 383.700 496.200 390.750 497.100 ;
        RECT 383.100 492.150 384.900 493.950 ;
        RECT 380.100 489.150 381.900 490.950 ;
        RECT 382.950 490.050 385.050 492.150 ;
        RECT 386.250 489.150 388.050 490.950 ;
        RECT 379.950 487.050 382.050 489.150 ;
        RECT 385.950 487.050 388.050 489.150 ;
        RECT 389.700 487.950 390.750 496.200 ;
        RECT 404.700 491.400 406.500 503.250 ;
        RECT 408.900 491.400 410.700 503.250 ;
        RECT 419.400 497.400 421.200 503.250 ;
        RECT 422.700 491.400 424.500 503.250 ;
        RECT 426.900 491.400 428.700 503.250 ;
        RECT 434.550 497.400 436.350 503.250 ;
        RECT 437.550 497.400 439.350 503.250 ;
        RECT 440.550 497.400 442.350 503.250 ;
        RECT 433.950 492.450 436.050 493.050 ;
        RECT 431.550 491.550 436.050 492.450 ;
        RECT 401.250 489.150 403.050 490.950 ;
        RECT 388.950 485.850 391.050 487.950 ;
        RECT 400.950 487.050 403.050 489.150 ;
        RECT 404.850 486.150 406.050 491.400 ;
        RECT 419.250 489.150 421.050 490.950 ;
        RECT 410.100 486.150 411.900 487.950 ;
        RECT 418.950 487.050 421.050 489.150 ;
        RECT 422.850 486.150 424.050 491.400 ;
        RECT 428.100 486.150 429.900 487.950 ;
        RECT 304.050 471.750 305.850 477.600 ;
        RECT 307.050 476.100 310.350 477.600 ;
        RECT 307.050 471.750 308.850 476.100 ;
        RECT 323.100 471.750 324.900 480.000 ;
        RECT 328.500 471.750 330.300 480.600 ;
        RECT 338.400 474.600 339.600 482.850 ;
        RECT 350.100 481.050 351.900 482.850 ;
        RECT 353.850 480.750 355.050 484.050 ;
        RECT 368.100 483.150 369.900 484.950 ;
        RECT 367.950 481.050 370.050 483.150 ;
        RECT 370.950 482.850 373.050 484.950 ;
        RECT 354.000 479.700 357.750 480.750 ;
        RECT 347.550 476.700 355.350 478.050 ;
        RECT 335.550 471.750 337.350 474.600 ;
        RECT 338.550 471.750 340.350 474.600 ;
        RECT 347.550 471.750 349.350 476.700 ;
        RECT 350.550 471.750 352.350 475.800 ;
        RECT 353.550 471.750 355.350 476.700 ;
        RECT 356.550 477.600 357.750 479.700 ;
        RECT 356.550 471.750 358.350 477.600 ;
        RECT 371.400 474.600 372.600 482.850 ;
        RECT 389.400 481.650 390.600 485.850 ;
        RECT 368.550 471.750 370.350 474.600 ;
        RECT 371.550 471.750 373.350 474.600 ;
        RECT 380.700 471.750 382.500 480.600 ;
        RECT 386.100 480.000 390.600 481.650 ;
        RECT 403.950 484.050 406.050 486.150 ;
        RECT 403.950 480.750 405.150 484.050 ;
        RECT 406.950 482.850 409.050 484.950 ;
        RECT 409.950 484.050 412.050 486.150 ;
        RECT 421.950 484.050 424.050 486.150 ;
        RECT 407.100 481.050 408.900 482.850 ;
        RECT 421.950 480.750 423.150 484.050 ;
        RECT 424.950 482.850 427.050 484.950 ;
        RECT 427.950 484.050 430.050 486.150 ;
        RECT 425.100 481.050 426.900 482.850 ;
        RECT 386.100 471.750 387.900 480.000 ;
        RECT 401.250 479.700 405.000 480.750 ;
        RECT 419.250 479.700 423.000 480.750 ;
        RECT 431.550 480.450 432.450 491.550 ;
        RECT 433.950 490.950 436.050 491.550 ;
        RECT 437.550 489.150 438.750 497.400 ;
        RECT 447.300 491.400 449.100 503.250 ;
        RECT 451.500 491.400 453.300 503.250 ;
        RECT 454.800 497.400 456.600 503.250 ;
        RECT 464.400 497.400 466.200 503.250 ;
        RECT 467.700 491.400 469.500 503.250 ;
        RECT 471.900 491.400 473.700 503.250 ;
        RECT 476.700 497.400 478.500 503.250 ;
        RECT 479.700 497.400 481.500 503.250 ;
        RECT 482.700 497.400 484.500 503.250 ;
        RECT 479.700 496.500 480.750 497.400 ;
        RECT 476.700 495.600 480.750 496.500 ;
        RECT 433.950 485.850 436.050 487.950 ;
        RECT 436.950 487.050 439.050 489.150 ;
        RECT 434.100 484.050 435.900 485.850 ;
        RECT 433.950 480.450 436.050 481.050 ;
        RECT 401.250 477.600 402.450 479.700 ;
        RECT 400.650 471.750 402.450 477.600 ;
        RECT 403.650 476.700 411.450 478.050 ;
        RECT 419.250 477.600 420.450 479.700 ;
        RECT 431.550 479.550 436.050 480.450 ;
        RECT 433.950 478.950 436.050 479.550 ;
        RECT 437.550 479.700 438.750 487.050 ;
        RECT 439.950 485.850 442.050 487.950 ;
        RECT 446.100 486.150 447.900 487.950 ;
        RECT 451.950 486.150 453.150 491.400 ;
        RECT 454.950 489.150 456.750 490.950 ;
        RECT 464.250 489.150 466.050 490.950 ;
        RECT 454.950 487.050 457.050 489.150 ;
        RECT 463.950 487.050 466.050 489.150 ;
        RECT 467.850 486.150 469.050 491.400 ;
        RECT 473.100 486.150 474.900 487.950 ;
        RECT 440.100 484.050 441.900 485.850 ;
        RECT 445.950 484.050 448.050 486.150 ;
        RECT 448.950 482.850 451.050 484.950 ;
        RECT 451.950 484.050 454.050 486.150 ;
        RECT 449.100 481.050 450.900 482.850 ;
        RECT 452.850 480.750 454.050 484.050 ;
        RECT 466.950 484.050 469.050 486.150 ;
        RECT 466.950 480.750 468.150 484.050 ;
        RECT 469.950 482.850 472.050 484.950 ;
        RECT 472.950 484.050 475.050 486.150 ;
        RECT 470.100 481.050 471.900 482.850 ;
        RECT 476.700 482.100 477.900 495.600 ;
        RECT 485.700 494.700 487.500 503.250 ;
        RECT 488.700 499.950 490.500 503.250 ;
        RECT 491.850 500.400 494.250 503.250 ;
        RECT 495.150 500.400 497.250 503.250 ;
        RECT 498.300 500.400 500.250 503.250 ;
        RECT 491.850 499.050 493.050 500.400 ;
        RECT 495.150 499.050 496.050 500.400 ;
        RECT 498.300 499.050 499.500 500.400 ;
        RECT 490.950 496.950 493.050 499.050 ;
        RECT 493.950 496.950 496.050 499.050 ;
        RECT 496.950 497.400 499.500 499.050 ;
        RECT 501.450 497.400 503.250 503.250 ;
        RECT 505.200 497.400 507.000 503.250 ;
        RECT 508.200 497.400 510.000 503.250 ;
        RECT 496.950 496.950 499.050 497.400 ;
        RECT 505.650 496.500 507.000 497.400 ;
        RECT 511.200 496.500 513.000 503.250 ;
        RECT 514.950 500.400 516.750 503.250 ;
        RECT 505.650 494.850 508.050 496.500 ;
        RECT 481.200 493.650 498.900 494.700 ;
        RECT 505.950 494.400 508.050 494.850 ;
        RECT 510.000 496.200 513.000 496.500 ;
        RECT 510.000 494.400 513.900 496.200 ;
        RECT 481.200 492.900 483.000 493.650 ;
        RECT 493.950 492.150 496.050 492.750 ;
        RECT 484.500 490.950 496.050 492.150 ;
        RECT 496.950 492.600 498.900 493.650 ;
        RECT 515.100 493.350 516.450 500.400 ;
        RECT 517.950 496.950 519.750 503.250 ;
        RECT 520.950 500.400 522.750 503.250 ;
        RECT 521.100 499.200 522.600 500.400 ;
        RECT 521.100 497.100 523.200 499.200 ;
        RECT 524.700 497.400 526.500 503.250 ;
        RECT 517.950 496.050 520.050 496.950 ;
        RECT 527.700 496.500 529.500 503.250 ;
        RECT 530.700 497.400 532.500 503.250 ;
        RECT 533.700 497.400 535.500 503.250 ;
        RECT 536.700 497.400 538.500 503.250 ;
        RECT 540.450 497.400 542.250 503.250 ;
        RECT 543.450 497.400 545.250 503.250 ;
        RECT 548.550 497.400 550.350 503.250 ;
        RECT 551.550 497.400 553.350 503.250 ;
        RECT 554.550 498.000 556.350 503.250 ;
        RECT 524.850 496.050 526.650 496.500 ;
        RECT 517.950 494.850 526.650 496.050 ;
        RECT 527.700 495.300 533.400 496.500 ;
        RECT 524.850 494.700 526.650 494.850 ;
        RECT 531.600 494.700 533.400 495.300 ;
        RECT 534.300 493.350 535.500 497.400 ;
        RECT 514.950 492.600 517.050 493.350 ;
        RECT 496.950 491.250 517.050 492.600 ;
        RECT 520.950 492.450 538.350 493.350 ;
        RECT 520.950 491.250 523.050 492.450 ;
        RECT 484.500 490.350 486.300 490.950 ;
        RECT 493.950 490.650 496.050 490.950 ;
        RECT 523.950 490.350 536.250 491.550 ;
        RECT 496.950 489.450 525.000 490.350 ;
        RECT 534.450 489.750 536.250 490.350 ;
        RECT 485.250 489.150 525.000 489.450 ;
        RECT 484.950 488.550 498.900 489.150 ;
        RECT 478.950 485.850 481.050 487.950 ;
        RECT 484.950 487.350 488.850 488.550 ;
        RECT 505.950 487.650 520.500 488.250 ;
        RECT 484.950 487.050 487.050 487.350 ;
        RECT 489.750 486.450 496.500 487.350 ;
        RECT 479.100 484.050 480.900 485.850 ;
        RECT 489.750 484.050 490.950 486.450 ;
        RECT 479.100 483.000 490.950 484.050 ;
        RECT 492.750 483.750 494.550 485.550 ;
        RECT 495.450 484.950 496.500 486.450 ;
        RECT 497.400 487.050 520.500 487.650 ;
        RECT 497.400 486.450 508.050 487.050 ;
        RECT 497.400 485.850 499.200 486.450 ;
        RECT 505.950 486.150 508.050 486.450 ;
        RECT 510.150 485.250 512.250 485.550 ;
        RECT 518.700 485.250 520.500 487.050 ;
        RECT 521.850 486.000 528.900 487.800 ;
        RECT 495.450 484.050 507.450 484.950 ;
        RECT 476.700 481.200 492.000 482.100 ;
        RECT 453.000 479.700 456.750 480.750 ;
        RECT 437.550 478.800 441.150 479.700 ;
        RECT 403.650 471.750 405.450 476.700 ;
        RECT 406.650 471.750 408.450 475.800 ;
        RECT 409.650 471.750 411.450 476.700 ;
        RECT 418.650 471.750 420.450 477.600 ;
        RECT 421.650 476.700 429.450 478.050 ;
        RECT 421.650 471.750 423.450 476.700 ;
        RECT 424.650 471.750 426.450 475.800 ;
        RECT 427.650 471.750 429.450 476.700 ;
        RECT 434.850 471.750 436.650 477.600 ;
        RECT 439.350 471.750 441.150 478.800 ;
        RECT 446.550 476.700 454.350 478.050 ;
        RECT 446.550 471.750 448.350 476.700 ;
        RECT 449.550 471.750 451.350 475.800 ;
        RECT 452.550 471.750 454.350 476.700 ;
        RECT 455.550 477.600 456.750 479.700 ;
        RECT 464.250 479.700 468.000 480.750 ;
        RECT 464.250 477.600 465.450 479.700 ;
        RECT 455.550 471.750 457.350 477.600 ;
        RECT 463.650 471.750 465.450 477.600 ;
        RECT 466.650 476.700 474.450 478.050 ;
        RECT 466.650 471.750 468.450 476.700 ;
        RECT 469.650 471.750 471.450 475.800 ;
        RECT 472.650 471.750 474.450 476.700 ;
        RECT 476.700 477.600 477.900 481.200 ;
        RECT 480.900 479.700 482.700 480.300 ;
        RECT 480.900 478.500 489.300 479.700 ;
        RECT 487.800 477.600 489.300 478.500 ;
        RECT 476.700 471.750 478.500 477.600 ;
        RECT 482.100 471.750 483.900 477.600 ;
        RECT 487.500 471.750 489.300 477.600 ;
        RECT 490.950 478.050 492.000 481.200 ;
        RECT 493.500 480.300 494.550 483.750 ;
        RECT 501.150 481.350 505.050 483.150 ;
        RECT 502.950 481.050 505.050 481.350 ;
        RECT 506.400 482.550 507.450 484.050 ;
        RECT 508.350 483.450 512.250 485.250 ;
        RECT 521.850 484.350 522.750 486.000 ;
        RECT 529.950 485.100 532.050 489.150 ;
        RECT 513.150 483.300 522.750 484.350 ;
        RECT 523.800 484.050 532.050 485.100 ;
        RECT 513.150 482.550 514.050 483.300 ;
        RECT 506.400 481.200 514.050 482.550 ;
        RECT 523.800 482.250 524.850 484.050 ;
        RECT 514.950 481.200 524.850 482.250 ;
        RECT 528.300 481.200 536.100 483.000 ;
        RECT 496.050 480.300 497.850 480.750 ;
        RECT 514.950 480.300 516.000 481.200 ;
        RECT 493.500 479.850 497.850 480.300 ;
        RECT 493.500 479.100 501.150 479.850 ;
        RECT 496.050 478.950 501.150 479.100 ;
        RECT 490.950 475.950 493.050 478.050 ;
        RECT 493.950 475.950 496.050 478.050 ;
        RECT 496.950 475.950 499.050 478.050 ;
        RECT 500.250 477.600 501.150 478.950 ;
        RECT 509.100 478.500 516.000 480.300 ;
        RECT 516.900 478.500 523.650 480.300 ;
        RECT 528.300 477.600 529.800 481.200 ;
        RECT 537.150 477.600 538.350 492.450 ;
        RECT 500.250 476.250 504.300 477.600 ;
        RECT 505.950 477.300 508.050 477.600 ;
        RECT 491.700 474.600 493.050 475.950 ;
        RECT 494.700 474.600 496.050 475.950 ;
        RECT 497.700 474.600 499.050 475.950 ;
        RECT 502.500 475.800 504.300 476.250 ;
        RECT 505.200 475.500 508.050 477.300 ;
        RECT 510.150 477.300 512.250 477.600 ;
        RECT 510.150 475.500 513.000 477.300 ;
        RECT 491.700 471.750 493.500 474.600 ;
        RECT 494.700 471.750 496.500 474.600 ;
        RECT 497.700 471.750 499.500 474.600 ;
        RECT 500.700 471.750 502.500 474.600 ;
        RECT 505.200 471.750 507.000 475.500 ;
        RECT 508.200 471.750 510.000 474.600 ;
        RECT 511.200 471.750 513.000 475.500 ;
        RECT 514.950 475.500 517.050 477.600 ;
        RECT 517.950 475.500 520.050 477.600 ;
        RECT 520.950 475.500 523.050 477.600 ;
        RECT 525.600 476.400 529.800 477.600 ;
        RECT 514.950 471.750 516.750 475.500 ;
        RECT 517.950 471.750 519.750 475.500 ;
        RECT 520.950 471.750 522.750 475.500 ;
        RECT 525.600 471.750 527.400 476.400 ;
        RECT 531.150 471.750 532.950 477.600 ;
        RECT 536.550 471.750 538.350 477.600 ;
        RECT 540.450 484.950 541.950 497.400 ;
        RECT 551.700 497.100 553.350 497.400 ;
        RECT 557.550 497.400 559.350 503.250 ;
        RECT 564.750 497.400 566.550 503.250 ;
        RECT 567.750 497.400 569.550 503.250 ;
        RECT 571.500 497.400 573.300 503.250 ;
        RECT 574.500 497.400 576.300 503.250 ;
        RECT 577.500 497.400 579.300 503.250 ;
        RECT 557.550 497.100 558.750 497.400 ;
        RECT 551.700 496.200 558.750 497.100 ;
        RECT 551.100 492.150 552.900 493.950 ;
        RECT 548.100 489.150 549.900 490.950 ;
        RECT 550.950 490.050 553.050 492.150 ;
        RECT 554.250 489.150 556.050 490.950 ;
        RECT 547.950 487.050 550.050 489.150 ;
        RECT 553.950 487.050 556.050 489.150 ;
        RECT 557.700 487.950 558.750 496.200 ;
        RECT 556.950 485.850 559.050 487.950 ;
        RECT 540.450 482.850 544.050 484.950 ;
        RECT 540.450 474.600 541.950 482.850 ;
        RECT 557.400 481.650 558.600 485.850 ;
        RECT 568.050 484.950 569.550 497.400 ;
        RECT 574.500 493.350 575.700 497.400 ;
        RECT 580.500 496.500 582.300 503.250 ;
        RECT 583.500 497.400 585.300 503.250 ;
        RECT 587.250 500.400 589.050 503.250 ;
        RECT 587.400 499.200 588.900 500.400 ;
        RECT 586.800 497.100 588.900 499.200 ;
        RECT 590.250 496.950 592.050 503.250 ;
        RECT 593.250 500.400 595.050 503.250 ;
        RECT 576.600 495.300 582.300 496.500 ;
        RECT 583.350 496.050 585.150 496.500 ;
        RECT 589.950 496.050 592.050 496.950 ;
        RECT 576.600 494.700 578.400 495.300 ;
        RECT 583.350 494.850 592.050 496.050 ;
        RECT 583.350 494.700 585.150 494.850 ;
        RECT 593.550 493.350 594.900 500.400 ;
        RECT 597.000 496.500 598.800 503.250 ;
        RECT 600.000 497.400 601.800 503.250 ;
        RECT 603.000 497.400 604.800 503.250 ;
        RECT 606.750 497.400 608.550 503.250 ;
        RECT 609.750 500.400 611.700 503.250 ;
        RECT 612.750 500.400 614.850 503.250 ;
        RECT 615.750 500.400 618.150 503.250 ;
        RECT 610.500 499.050 611.700 500.400 ;
        RECT 613.950 499.050 614.850 500.400 ;
        RECT 616.950 499.050 618.150 500.400 ;
        RECT 619.500 499.950 621.300 503.250 ;
        RECT 610.500 497.400 613.050 499.050 ;
        RECT 603.000 496.500 604.350 497.400 ;
        RECT 610.950 496.950 613.050 497.400 ;
        RECT 613.950 496.950 616.050 499.050 ;
        RECT 616.950 496.950 619.050 499.050 ;
        RECT 597.000 496.200 600.000 496.500 ;
        RECT 596.100 494.400 600.000 496.200 ;
        RECT 601.950 494.850 604.350 496.500 ;
        RECT 601.950 494.400 604.050 494.850 ;
        RECT 622.500 494.700 624.300 503.250 ;
        RECT 625.500 497.400 627.300 503.250 ;
        RECT 628.500 497.400 630.300 503.250 ;
        RECT 631.500 497.400 633.300 503.250 ;
        RECT 643.650 497.400 645.450 503.250 ;
        RECT 646.650 497.400 648.450 503.250 ;
        RECT 651.750 497.400 653.550 503.250 ;
        RECT 654.750 497.400 656.550 503.250 ;
        RECT 658.500 497.400 660.300 503.250 ;
        RECT 661.500 497.400 663.300 503.250 ;
        RECT 664.500 497.400 666.300 503.250 ;
        RECT 629.250 496.500 630.300 497.400 ;
        RECT 629.250 495.600 633.300 496.500 ;
        RECT 611.100 493.650 628.800 494.700 ;
        RECT 565.950 482.850 569.550 484.950 ;
        RECT 540.450 471.750 542.250 474.600 ;
        RECT 543.450 471.750 545.250 474.600 ;
        RECT 548.700 471.750 550.500 480.600 ;
        RECT 554.100 480.000 558.600 481.650 ;
        RECT 554.100 471.750 555.900 480.000 ;
        RECT 568.050 474.600 569.550 482.850 ;
        RECT 564.750 471.750 566.550 474.600 ;
        RECT 567.750 471.750 569.550 474.600 ;
        RECT 571.650 492.450 589.050 493.350 ;
        RECT 571.650 477.600 572.850 492.450 ;
        RECT 573.750 490.350 586.050 491.550 ;
        RECT 586.950 491.250 589.050 492.450 ;
        RECT 592.950 492.600 595.050 493.350 ;
        RECT 611.100 492.600 613.050 493.650 ;
        RECT 627.000 492.900 628.800 493.650 ;
        RECT 592.950 491.250 613.050 492.600 ;
        RECT 613.950 492.150 616.050 492.750 ;
        RECT 613.950 490.950 625.500 492.150 ;
        RECT 613.950 490.650 616.050 490.950 ;
        RECT 623.700 490.350 625.500 490.950 ;
        RECT 573.750 489.750 575.550 490.350 ;
        RECT 585.000 489.450 613.050 490.350 ;
        RECT 585.000 489.150 624.750 489.450 ;
        RECT 577.950 485.100 580.050 489.150 ;
        RECT 611.100 488.550 625.050 489.150 ;
        RECT 581.100 486.000 588.150 487.800 ;
        RECT 577.950 484.050 586.200 485.100 ;
        RECT 573.900 481.200 581.700 483.000 ;
        RECT 585.150 482.250 586.200 484.050 ;
        RECT 587.250 484.350 588.150 486.000 ;
        RECT 589.500 487.650 604.050 488.250 ;
        RECT 589.500 487.050 612.600 487.650 ;
        RECT 621.150 487.350 625.050 488.550 ;
        RECT 589.500 485.250 591.300 487.050 ;
        RECT 601.950 486.450 612.600 487.050 ;
        RECT 601.950 486.150 604.050 486.450 ;
        RECT 610.800 485.850 612.600 486.450 ;
        RECT 613.500 486.450 620.250 487.350 ;
        RECT 622.950 487.050 625.050 487.350 ;
        RECT 597.750 485.250 599.850 485.550 ;
        RECT 587.250 483.300 596.850 484.350 ;
        RECT 597.750 483.450 601.650 485.250 ;
        RECT 613.500 484.950 614.550 486.450 ;
        RECT 602.550 484.050 614.550 484.950 ;
        RECT 595.950 482.550 596.850 483.300 ;
        RECT 602.550 482.550 603.600 484.050 ;
        RECT 615.450 483.750 617.250 485.550 ;
        RECT 619.050 484.050 620.250 486.450 ;
        RECT 628.950 485.850 631.050 487.950 ;
        RECT 629.100 484.050 630.900 485.850 ;
        RECT 585.150 481.200 595.050 482.250 ;
        RECT 595.950 481.200 603.600 482.550 ;
        RECT 604.950 481.350 608.850 483.150 ;
        RECT 580.200 477.600 581.700 481.200 ;
        RECT 594.000 480.300 595.050 481.200 ;
        RECT 604.950 481.050 607.050 481.350 ;
        RECT 612.150 480.300 613.950 480.750 ;
        RECT 615.450 480.300 616.500 483.750 ;
        RECT 619.050 483.000 630.900 484.050 ;
        RECT 632.100 482.100 633.300 495.600 ;
        RECT 644.400 484.950 645.600 497.400 ;
        RECT 655.050 484.950 656.550 497.400 ;
        RECT 661.500 493.350 662.700 497.400 ;
        RECT 667.500 496.500 669.300 503.250 ;
        RECT 670.500 497.400 672.300 503.250 ;
        RECT 674.250 500.400 676.050 503.250 ;
        RECT 674.400 499.200 675.900 500.400 ;
        RECT 673.800 497.100 675.900 499.200 ;
        RECT 677.250 496.950 679.050 503.250 ;
        RECT 680.250 500.400 682.050 503.250 ;
        RECT 663.600 495.300 669.300 496.500 ;
        RECT 670.350 496.050 672.150 496.500 ;
        RECT 676.950 496.050 679.050 496.950 ;
        RECT 663.600 494.700 665.400 495.300 ;
        RECT 670.350 494.850 679.050 496.050 ;
        RECT 670.350 494.700 672.150 494.850 ;
        RECT 680.550 493.350 681.900 500.400 ;
        RECT 684.000 496.500 685.800 503.250 ;
        RECT 687.000 497.400 688.800 503.250 ;
        RECT 690.000 497.400 691.800 503.250 ;
        RECT 693.750 497.400 695.550 503.250 ;
        RECT 696.750 500.400 698.700 503.250 ;
        RECT 699.750 500.400 701.850 503.250 ;
        RECT 702.750 500.400 705.150 503.250 ;
        RECT 697.500 499.050 698.700 500.400 ;
        RECT 700.950 499.050 701.850 500.400 ;
        RECT 703.950 499.050 705.150 500.400 ;
        RECT 706.500 499.950 708.300 503.250 ;
        RECT 697.500 497.400 700.050 499.050 ;
        RECT 690.000 496.500 691.350 497.400 ;
        RECT 697.950 496.950 700.050 497.400 ;
        RECT 700.950 496.950 703.050 499.050 ;
        RECT 703.950 496.950 706.050 499.050 ;
        RECT 684.000 496.200 687.000 496.500 ;
        RECT 683.100 494.400 687.000 496.200 ;
        RECT 688.950 494.850 691.350 496.500 ;
        RECT 688.950 494.400 691.050 494.850 ;
        RECT 709.500 494.700 711.300 503.250 ;
        RECT 712.500 497.400 714.300 503.250 ;
        RECT 715.500 497.400 717.300 503.250 ;
        RECT 718.500 497.400 720.300 503.250 ;
        RECT 716.250 496.500 717.300 497.400 ;
        RECT 716.250 495.600 720.300 496.500 ;
        RECT 698.100 493.650 715.800 494.700 ;
        RECT 643.950 482.850 646.050 484.950 ;
        RECT 647.100 483.150 648.900 484.950 ;
        RECT 586.350 478.500 593.100 480.300 ;
        RECT 594.000 478.500 600.900 480.300 ;
        RECT 612.150 479.850 616.500 480.300 ;
        RECT 608.850 479.100 616.500 479.850 ;
        RECT 618.000 481.200 633.300 482.100 ;
        RECT 608.850 478.950 613.950 479.100 ;
        RECT 608.850 477.600 609.750 478.950 ;
        RECT 618.000 478.050 619.050 481.200 ;
        RECT 627.300 479.700 629.100 480.300 ;
        RECT 571.650 471.750 573.450 477.600 ;
        RECT 577.050 471.750 578.850 477.600 ;
        RECT 580.200 476.400 584.400 477.600 ;
        RECT 582.600 471.750 584.400 476.400 ;
        RECT 586.950 475.500 589.050 477.600 ;
        RECT 589.950 475.500 592.050 477.600 ;
        RECT 592.950 475.500 595.050 477.600 ;
        RECT 597.750 477.300 599.850 477.600 ;
        RECT 587.250 471.750 589.050 475.500 ;
        RECT 590.250 471.750 592.050 475.500 ;
        RECT 593.250 471.750 595.050 475.500 ;
        RECT 597.000 475.500 599.850 477.300 ;
        RECT 601.950 477.300 604.050 477.600 ;
        RECT 601.950 475.500 604.800 477.300 ;
        RECT 605.700 476.250 609.750 477.600 ;
        RECT 605.700 475.800 607.500 476.250 ;
        RECT 610.950 475.950 613.050 478.050 ;
        RECT 613.950 475.950 616.050 478.050 ;
        RECT 616.950 475.950 619.050 478.050 ;
        RECT 620.700 478.500 629.100 479.700 ;
        RECT 620.700 477.600 622.200 478.500 ;
        RECT 632.100 477.600 633.300 481.200 ;
        RECT 597.000 471.750 598.800 475.500 ;
        RECT 600.000 471.750 601.800 474.600 ;
        RECT 603.000 471.750 604.800 475.500 ;
        RECT 610.950 474.600 612.300 475.950 ;
        RECT 613.950 474.600 615.300 475.950 ;
        RECT 616.950 474.600 618.300 475.950 ;
        RECT 607.500 471.750 609.300 474.600 ;
        RECT 610.500 471.750 612.300 474.600 ;
        RECT 613.500 471.750 615.300 474.600 ;
        RECT 616.500 471.750 618.300 474.600 ;
        RECT 620.700 471.750 622.500 477.600 ;
        RECT 626.100 471.750 627.900 477.600 ;
        RECT 631.500 471.750 633.300 477.600 ;
        RECT 644.400 474.600 645.600 482.850 ;
        RECT 646.950 481.050 649.050 483.150 ;
        RECT 652.950 482.850 656.550 484.950 ;
        RECT 655.050 474.600 656.550 482.850 ;
        RECT 643.650 471.750 645.450 474.600 ;
        RECT 646.650 471.750 648.450 474.600 ;
        RECT 651.750 471.750 653.550 474.600 ;
        RECT 654.750 471.750 656.550 474.600 ;
        RECT 658.650 492.450 676.050 493.350 ;
        RECT 658.650 477.600 659.850 492.450 ;
        RECT 660.750 490.350 673.050 491.550 ;
        RECT 673.950 491.250 676.050 492.450 ;
        RECT 679.950 492.600 682.050 493.350 ;
        RECT 698.100 492.600 700.050 493.650 ;
        RECT 714.000 492.900 715.800 493.650 ;
        RECT 679.950 491.250 700.050 492.600 ;
        RECT 700.950 492.150 703.050 492.750 ;
        RECT 700.950 490.950 712.500 492.150 ;
        RECT 700.950 490.650 703.050 490.950 ;
        RECT 710.700 490.350 712.500 490.950 ;
        RECT 660.750 489.750 662.550 490.350 ;
        RECT 672.000 489.450 700.050 490.350 ;
        RECT 672.000 489.150 711.750 489.450 ;
        RECT 664.950 485.100 667.050 489.150 ;
        RECT 698.100 488.550 712.050 489.150 ;
        RECT 668.100 486.000 675.150 487.800 ;
        RECT 664.950 484.050 673.200 485.100 ;
        RECT 660.900 481.200 668.700 483.000 ;
        RECT 672.150 482.250 673.200 484.050 ;
        RECT 674.250 484.350 675.150 486.000 ;
        RECT 676.500 487.650 691.050 488.250 ;
        RECT 676.500 487.050 699.600 487.650 ;
        RECT 708.150 487.350 712.050 488.550 ;
        RECT 676.500 485.250 678.300 487.050 ;
        RECT 688.950 486.450 699.600 487.050 ;
        RECT 688.950 486.150 691.050 486.450 ;
        RECT 697.800 485.850 699.600 486.450 ;
        RECT 700.500 486.450 707.250 487.350 ;
        RECT 709.950 487.050 712.050 487.350 ;
        RECT 684.750 485.250 686.850 485.550 ;
        RECT 674.250 483.300 683.850 484.350 ;
        RECT 684.750 483.450 688.650 485.250 ;
        RECT 700.500 484.950 701.550 486.450 ;
        RECT 689.550 484.050 701.550 484.950 ;
        RECT 682.950 482.550 683.850 483.300 ;
        RECT 689.550 482.550 690.600 484.050 ;
        RECT 702.450 483.750 704.250 485.550 ;
        RECT 706.050 484.050 707.250 486.450 ;
        RECT 715.950 485.850 718.050 487.950 ;
        RECT 716.100 484.050 717.900 485.850 ;
        RECT 672.150 481.200 682.050 482.250 ;
        RECT 682.950 481.200 690.600 482.550 ;
        RECT 691.950 481.350 695.850 483.150 ;
        RECT 667.200 477.600 668.700 481.200 ;
        RECT 681.000 480.300 682.050 481.200 ;
        RECT 691.950 481.050 694.050 481.350 ;
        RECT 699.150 480.300 700.950 480.750 ;
        RECT 702.450 480.300 703.500 483.750 ;
        RECT 706.050 483.000 717.900 484.050 ;
        RECT 719.100 482.100 720.300 495.600 ;
        RECT 727.650 491.400 729.450 503.250 ;
        RECT 730.650 491.400 732.450 503.250 ;
        RECT 734.550 497.400 736.350 503.250 ;
        RECT 728.400 486.150 729.600 491.400 ;
        RECT 734.550 490.500 735.750 497.400 ;
        RECT 737.850 491.400 739.650 503.250 ;
        RECT 740.850 491.400 742.650 503.250 ;
        RECT 749.550 491.400 751.350 503.250 ;
        RECT 753.750 491.400 755.550 503.250 ;
        RECT 764.550 497.400 766.350 503.250 ;
        RECT 767.550 497.400 769.350 503.250 ;
        RECT 770.550 498.000 772.350 503.250 ;
        RECT 767.700 497.100 769.350 497.400 ;
        RECT 773.550 497.400 775.350 503.250 ;
        RECT 780.750 497.400 782.550 503.250 ;
        RECT 783.750 497.400 785.550 503.250 ;
        RECT 787.500 497.400 789.300 503.250 ;
        RECT 790.500 497.400 792.300 503.250 ;
        RECT 793.500 497.400 795.300 503.250 ;
        RECT 773.550 497.100 774.750 497.400 ;
        RECT 767.700 496.200 774.750 497.100 ;
        RECT 767.100 492.150 768.900 493.950 ;
        RECT 734.550 489.600 740.250 490.500 ;
        RECT 738.000 488.700 740.250 489.600 ;
        RECT 734.100 486.150 735.900 487.950 ;
        RECT 727.950 484.050 730.050 486.150 ;
        RECT 673.350 478.500 680.100 480.300 ;
        RECT 681.000 478.500 687.900 480.300 ;
        RECT 699.150 479.850 703.500 480.300 ;
        RECT 695.850 479.100 703.500 479.850 ;
        RECT 705.000 481.200 720.300 482.100 ;
        RECT 695.850 478.950 700.950 479.100 ;
        RECT 695.850 477.600 696.750 478.950 ;
        RECT 705.000 478.050 706.050 481.200 ;
        RECT 714.300 479.700 716.100 480.300 ;
        RECT 658.650 471.750 660.450 477.600 ;
        RECT 664.050 471.750 665.850 477.600 ;
        RECT 667.200 476.400 671.400 477.600 ;
        RECT 669.600 471.750 671.400 476.400 ;
        RECT 673.950 475.500 676.050 477.600 ;
        RECT 676.950 475.500 679.050 477.600 ;
        RECT 679.950 475.500 682.050 477.600 ;
        RECT 684.750 477.300 686.850 477.600 ;
        RECT 674.250 471.750 676.050 475.500 ;
        RECT 677.250 471.750 679.050 475.500 ;
        RECT 680.250 471.750 682.050 475.500 ;
        RECT 684.000 475.500 686.850 477.300 ;
        RECT 688.950 477.300 691.050 477.600 ;
        RECT 688.950 475.500 691.800 477.300 ;
        RECT 692.700 476.250 696.750 477.600 ;
        RECT 692.700 475.800 694.500 476.250 ;
        RECT 697.950 475.950 700.050 478.050 ;
        RECT 700.950 475.950 703.050 478.050 ;
        RECT 703.950 475.950 706.050 478.050 ;
        RECT 707.700 478.500 716.100 479.700 ;
        RECT 707.700 477.600 709.200 478.500 ;
        RECT 719.100 477.600 720.300 481.200 ;
        RECT 728.400 477.600 729.600 484.050 ;
        RECT 730.950 482.850 733.050 484.950 ;
        RECT 733.950 484.050 736.050 486.150 ;
        RECT 731.100 481.050 732.900 482.850 ;
        RECT 738.000 480.300 739.050 488.700 ;
        RECT 741.150 486.150 742.350 491.400 ;
        RECT 753.000 490.350 755.550 491.400 ;
        RECT 749.100 486.150 750.900 487.950 ;
        RECT 739.950 484.050 742.350 486.150 ;
        RECT 748.950 484.050 751.050 486.150 ;
        RECT 738.000 479.400 740.250 480.300 ;
        RECT 735.150 478.500 740.250 479.400 ;
        RECT 684.000 471.750 685.800 475.500 ;
        RECT 687.000 471.750 688.800 474.600 ;
        RECT 690.000 471.750 691.800 475.500 ;
        RECT 697.950 474.600 699.300 475.950 ;
        RECT 700.950 474.600 702.300 475.950 ;
        RECT 703.950 474.600 705.300 475.950 ;
        RECT 694.500 471.750 696.300 474.600 ;
        RECT 697.500 471.750 699.300 474.600 ;
        RECT 700.500 471.750 702.300 474.600 ;
        RECT 703.500 471.750 705.300 474.600 ;
        RECT 707.700 471.750 709.500 477.600 ;
        RECT 713.100 471.750 714.900 477.600 ;
        RECT 718.500 471.750 720.300 477.600 ;
        RECT 727.650 471.750 729.450 477.600 ;
        RECT 730.650 471.750 732.450 477.600 ;
        RECT 735.150 474.600 736.350 478.500 ;
        RECT 741.150 477.600 742.350 484.050 ;
        RECT 753.000 483.150 754.050 490.350 ;
        RECT 764.100 489.150 765.900 490.950 ;
        RECT 766.950 490.050 769.050 492.150 ;
        RECT 770.250 489.150 772.050 490.950 ;
        RECT 755.100 486.150 756.900 487.950 ;
        RECT 763.950 487.050 766.050 489.150 ;
        RECT 769.950 487.050 772.050 489.150 ;
        RECT 773.700 487.950 774.750 496.200 ;
        RECT 754.950 484.050 757.050 486.150 ;
        RECT 772.950 485.850 775.050 487.950 ;
        RECT 751.950 481.050 754.050 483.150 ;
        RECT 773.400 481.650 774.600 485.850 ;
        RECT 784.050 484.950 785.550 497.400 ;
        RECT 790.500 493.350 791.700 497.400 ;
        RECT 796.500 496.500 798.300 503.250 ;
        RECT 799.500 497.400 801.300 503.250 ;
        RECT 803.250 500.400 805.050 503.250 ;
        RECT 803.400 499.200 804.900 500.400 ;
        RECT 802.800 497.100 804.900 499.200 ;
        RECT 806.250 496.950 808.050 503.250 ;
        RECT 809.250 500.400 811.050 503.250 ;
        RECT 792.600 495.300 798.300 496.500 ;
        RECT 799.350 496.050 801.150 496.500 ;
        RECT 805.950 496.050 808.050 496.950 ;
        RECT 792.600 494.700 794.400 495.300 ;
        RECT 799.350 494.850 808.050 496.050 ;
        RECT 799.350 494.700 801.150 494.850 ;
        RECT 809.550 493.350 810.900 500.400 ;
        RECT 813.000 496.500 814.800 503.250 ;
        RECT 816.000 497.400 817.800 503.250 ;
        RECT 819.000 497.400 820.800 503.250 ;
        RECT 822.750 497.400 824.550 503.250 ;
        RECT 825.750 500.400 827.700 503.250 ;
        RECT 828.750 500.400 830.850 503.250 ;
        RECT 831.750 500.400 834.150 503.250 ;
        RECT 826.500 499.050 827.700 500.400 ;
        RECT 829.950 499.050 830.850 500.400 ;
        RECT 832.950 499.050 834.150 500.400 ;
        RECT 835.500 499.950 837.300 503.250 ;
        RECT 826.500 497.400 829.050 499.050 ;
        RECT 819.000 496.500 820.350 497.400 ;
        RECT 826.950 496.950 829.050 497.400 ;
        RECT 829.950 496.950 832.050 499.050 ;
        RECT 832.950 496.950 835.050 499.050 ;
        RECT 813.000 496.200 816.000 496.500 ;
        RECT 812.100 494.400 816.000 496.200 ;
        RECT 817.950 494.850 820.350 496.500 ;
        RECT 817.950 494.400 820.050 494.850 ;
        RECT 838.500 494.700 840.300 503.250 ;
        RECT 841.500 497.400 843.300 503.250 ;
        RECT 844.500 497.400 846.300 503.250 ;
        RECT 847.500 497.400 849.300 503.250 ;
        RECT 845.250 496.500 846.300 497.400 ;
        RECT 845.250 495.600 849.300 496.500 ;
        RECT 827.100 493.650 844.800 494.700 ;
        RECT 781.950 482.850 785.550 484.950 ;
        RECT 734.550 471.750 736.350 474.600 ;
        RECT 737.850 471.750 739.650 477.600 ;
        RECT 740.850 471.750 742.650 477.600 ;
        RECT 753.000 474.600 754.050 481.050 ;
        RECT 749.550 471.750 751.350 474.600 ;
        RECT 752.550 471.750 754.350 474.600 ;
        RECT 755.550 471.750 757.350 474.600 ;
        RECT 764.700 471.750 766.500 480.600 ;
        RECT 770.100 480.000 774.600 481.650 ;
        RECT 770.100 471.750 771.900 480.000 ;
        RECT 784.050 474.600 785.550 482.850 ;
        RECT 780.750 471.750 782.550 474.600 ;
        RECT 783.750 471.750 785.550 474.600 ;
        RECT 787.650 492.450 805.050 493.350 ;
        RECT 787.650 477.600 788.850 492.450 ;
        RECT 789.750 490.350 802.050 491.550 ;
        RECT 802.950 491.250 805.050 492.450 ;
        RECT 808.950 492.600 811.050 493.350 ;
        RECT 827.100 492.600 829.050 493.650 ;
        RECT 843.000 492.900 844.800 493.650 ;
        RECT 808.950 491.250 829.050 492.600 ;
        RECT 829.950 492.150 832.050 492.750 ;
        RECT 829.950 490.950 841.500 492.150 ;
        RECT 829.950 490.650 832.050 490.950 ;
        RECT 839.700 490.350 841.500 490.950 ;
        RECT 789.750 489.750 791.550 490.350 ;
        RECT 801.000 489.450 829.050 490.350 ;
        RECT 801.000 489.150 840.750 489.450 ;
        RECT 793.950 485.100 796.050 489.150 ;
        RECT 827.100 488.550 841.050 489.150 ;
        RECT 797.100 486.000 804.150 487.800 ;
        RECT 793.950 484.050 802.200 485.100 ;
        RECT 789.900 481.200 797.700 483.000 ;
        RECT 801.150 482.250 802.200 484.050 ;
        RECT 803.250 484.350 804.150 486.000 ;
        RECT 805.500 487.650 820.050 488.250 ;
        RECT 805.500 487.050 828.600 487.650 ;
        RECT 837.150 487.350 841.050 488.550 ;
        RECT 805.500 485.250 807.300 487.050 ;
        RECT 817.950 486.450 828.600 487.050 ;
        RECT 817.950 486.150 820.050 486.450 ;
        RECT 826.800 485.850 828.600 486.450 ;
        RECT 829.500 486.450 836.250 487.350 ;
        RECT 838.950 487.050 841.050 487.350 ;
        RECT 813.750 485.250 815.850 485.550 ;
        RECT 803.250 483.300 812.850 484.350 ;
        RECT 813.750 483.450 817.650 485.250 ;
        RECT 829.500 484.950 830.550 486.450 ;
        RECT 818.550 484.050 830.550 484.950 ;
        RECT 811.950 482.550 812.850 483.300 ;
        RECT 818.550 482.550 819.600 484.050 ;
        RECT 831.450 483.750 833.250 485.550 ;
        RECT 835.050 484.050 836.250 486.450 ;
        RECT 844.950 485.850 847.050 487.950 ;
        RECT 845.100 484.050 846.900 485.850 ;
        RECT 801.150 481.200 811.050 482.250 ;
        RECT 811.950 481.200 819.600 482.550 ;
        RECT 820.950 481.350 824.850 483.150 ;
        RECT 796.200 477.600 797.700 481.200 ;
        RECT 810.000 480.300 811.050 481.200 ;
        RECT 820.950 481.050 823.050 481.350 ;
        RECT 828.150 480.300 829.950 480.750 ;
        RECT 831.450 480.300 832.500 483.750 ;
        RECT 835.050 483.000 846.900 484.050 ;
        RECT 848.100 482.100 849.300 495.600 ;
        RECT 802.350 478.500 809.100 480.300 ;
        RECT 810.000 478.500 816.900 480.300 ;
        RECT 828.150 479.850 832.500 480.300 ;
        RECT 824.850 479.100 832.500 479.850 ;
        RECT 834.000 481.200 849.300 482.100 ;
        RECT 824.850 478.950 829.950 479.100 ;
        RECT 824.850 477.600 825.750 478.950 ;
        RECT 834.000 478.050 835.050 481.200 ;
        RECT 843.300 479.700 845.100 480.300 ;
        RECT 787.650 471.750 789.450 477.600 ;
        RECT 793.050 471.750 794.850 477.600 ;
        RECT 796.200 476.400 800.400 477.600 ;
        RECT 798.600 471.750 800.400 476.400 ;
        RECT 802.950 475.500 805.050 477.600 ;
        RECT 805.950 475.500 808.050 477.600 ;
        RECT 808.950 475.500 811.050 477.600 ;
        RECT 813.750 477.300 815.850 477.600 ;
        RECT 803.250 471.750 805.050 475.500 ;
        RECT 806.250 471.750 808.050 475.500 ;
        RECT 809.250 471.750 811.050 475.500 ;
        RECT 813.000 475.500 815.850 477.300 ;
        RECT 817.950 477.300 820.050 477.600 ;
        RECT 817.950 475.500 820.800 477.300 ;
        RECT 821.700 476.250 825.750 477.600 ;
        RECT 821.700 475.800 823.500 476.250 ;
        RECT 826.950 475.950 829.050 478.050 ;
        RECT 829.950 475.950 832.050 478.050 ;
        RECT 832.950 475.950 835.050 478.050 ;
        RECT 836.700 478.500 845.100 479.700 ;
        RECT 836.700 477.600 838.200 478.500 ;
        RECT 848.100 477.600 849.300 481.200 ;
        RECT 813.000 471.750 814.800 475.500 ;
        RECT 816.000 471.750 817.800 474.600 ;
        RECT 819.000 471.750 820.800 475.500 ;
        RECT 826.950 474.600 828.300 475.950 ;
        RECT 829.950 474.600 831.300 475.950 ;
        RECT 832.950 474.600 834.300 475.950 ;
        RECT 823.500 471.750 825.300 474.600 ;
        RECT 826.500 471.750 828.300 474.600 ;
        RECT 829.500 471.750 831.300 474.600 ;
        RECT 832.500 471.750 834.300 474.600 ;
        RECT 836.700 471.750 838.500 477.600 ;
        RECT 842.100 471.750 843.900 477.600 ;
        RECT 847.500 471.750 849.300 477.600 ;
        RECT 8.850 460.200 10.650 467.250 ;
        RECT 13.350 461.400 15.150 467.250 ;
        RECT 22.650 464.400 24.450 467.250 ;
        RECT 25.650 464.400 27.450 467.250 ;
        RECT 28.650 464.400 30.450 467.250 ;
        RECT 8.850 459.300 12.450 460.200 ;
        RECT 8.100 453.150 9.900 454.950 ;
        RECT 7.950 451.050 10.050 453.150 ;
        RECT 11.250 451.950 12.450 459.300 ;
        RECT 25.950 457.950 27.000 464.400 ;
        RECT 35.550 459.900 37.350 467.250 ;
        RECT 40.050 461.400 41.850 467.250 ;
        RECT 43.050 462.900 44.850 467.250 ;
        RECT 43.050 461.400 46.350 462.900 ;
        RECT 55.650 461.400 57.450 467.250 ;
        RECT 41.250 459.900 43.050 460.500 ;
        RECT 35.550 458.700 43.050 459.900 ;
        RECT 25.950 455.850 28.050 457.950 ;
        RECT 14.100 453.150 15.900 454.950 ;
        RECT 10.950 449.850 13.050 451.950 ;
        RECT 13.950 451.050 16.050 453.150 ;
        RECT 22.950 452.850 25.050 454.950 ;
        RECT 23.100 451.050 24.900 452.850 ;
        RECT 11.250 441.600 12.450 449.850 ;
        RECT 25.950 448.650 27.000 455.850 ;
        RECT 28.950 452.850 31.050 454.950 ;
        RECT 34.950 452.850 37.050 454.950 ;
        RECT 29.100 451.050 30.900 452.850 ;
        RECT 35.100 451.050 36.900 452.850 ;
        RECT 24.450 447.600 27.000 448.650 ;
        RECT 7.650 435.750 9.450 441.600 ;
        RECT 10.650 435.750 12.450 441.600 ;
        RECT 13.650 435.750 15.450 441.600 ;
        RECT 24.450 435.750 26.250 447.600 ;
        RECT 28.650 435.750 30.450 447.600 ;
        RECT 38.700 441.600 39.900 458.700 ;
        RECT 45.150 454.950 46.350 461.400 ;
        RECT 56.250 459.300 57.450 461.400 ;
        RECT 58.650 462.300 60.450 467.250 ;
        RECT 61.650 463.200 63.450 467.250 ;
        RECT 64.650 462.300 66.450 467.250 ;
        RECT 71.550 464.400 73.350 467.250 ;
        RECT 74.550 464.400 76.350 467.250 ;
        RECT 77.550 464.400 79.350 467.250 ;
        RECT 88.650 464.400 90.450 467.250 ;
        RECT 91.650 464.400 93.450 467.250 ;
        RECT 94.650 464.400 96.450 467.250 ;
        RECT 58.650 460.950 66.450 462.300 ;
        RECT 56.250 458.250 60.000 459.300 ;
        RECT 41.100 453.150 42.900 454.950 ;
        RECT 40.950 451.050 43.050 453.150 ;
        RECT 43.950 452.850 46.350 454.950 ;
        RECT 58.950 454.950 60.150 458.250 ;
        RECT 75.000 457.950 76.050 464.400 ;
        RECT 62.100 456.150 63.900 457.950 ;
        RECT 58.950 452.850 61.050 454.950 ;
        RECT 61.950 454.050 64.050 456.150 ;
        RECT 73.950 455.850 76.050 457.950 ;
        RECT 64.950 452.850 67.050 454.950 ;
        RECT 70.950 452.850 73.050 454.950 ;
        RECT 45.150 447.600 46.350 452.850 ;
        RECT 55.950 449.850 58.050 451.950 ;
        RECT 56.250 448.050 58.050 449.850 ;
        RECT 59.850 447.600 61.050 452.850 ;
        RECT 65.100 451.050 66.900 452.850 ;
        RECT 71.100 451.050 72.900 452.850 ;
        RECT 75.000 448.650 76.050 455.850 ;
        RECT 91.950 457.950 93.000 464.400 ;
        RECT 94.950 459.450 97.050 460.050 ;
        RECT 100.950 459.450 103.050 460.050 ;
        RECT 94.950 458.550 103.050 459.450 ;
        RECT 94.950 457.950 97.050 458.550 ;
        RECT 100.950 457.950 103.050 458.550 ;
        RECT 104.700 458.400 106.500 467.250 ;
        RECT 110.100 459.000 111.900 467.250 ;
        RECT 122.550 464.400 124.350 467.250 ;
        RECT 125.550 464.400 127.350 467.250 ;
        RECT 134.550 464.400 136.350 467.250 ;
        RECT 137.550 464.400 139.350 467.250 ;
        RECT 91.950 455.850 94.050 457.950 ;
        RECT 110.100 457.350 114.600 459.000 ;
        RECT 76.950 452.850 79.050 454.950 ;
        RECT 88.950 452.850 91.050 454.950 ;
        RECT 77.100 451.050 78.900 452.850 ;
        RECT 89.100 451.050 90.900 452.850 ;
        RECT 91.950 448.650 93.000 455.850 ;
        RECT 94.950 452.850 97.050 454.950 ;
        RECT 113.400 453.150 114.600 457.350 ;
        RECT 121.950 455.850 124.050 457.950 ;
        RECT 125.400 456.150 126.600 464.400 ;
        RECT 122.100 454.050 123.900 455.850 ;
        RECT 124.950 454.050 127.050 456.150 ;
        RECT 133.950 455.850 136.050 457.950 ;
        RECT 137.400 456.150 138.600 464.400 ;
        RECT 143.700 461.400 145.500 467.250 ;
        RECT 149.100 461.400 150.900 467.250 ;
        RECT 154.500 461.400 156.300 467.250 ;
        RECT 158.700 464.400 160.500 467.250 ;
        RECT 161.700 464.400 163.500 467.250 ;
        RECT 164.700 464.400 166.500 467.250 ;
        RECT 167.700 464.400 169.500 467.250 ;
        RECT 158.700 463.050 160.050 464.400 ;
        RECT 161.700 463.050 163.050 464.400 ;
        RECT 164.700 463.050 166.050 464.400 ;
        RECT 172.200 463.500 174.000 467.250 ;
        RECT 175.200 464.400 177.000 467.250 ;
        RECT 178.200 463.500 180.000 467.250 ;
        RECT 143.700 457.800 144.900 461.400 ;
        RECT 154.800 460.500 156.300 461.400 ;
        RECT 147.900 459.300 156.300 460.500 ;
        RECT 157.950 460.950 160.050 463.050 ;
        RECT 160.950 460.950 163.050 463.050 ;
        RECT 163.950 460.950 166.050 463.050 ;
        RECT 169.500 462.750 171.300 463.200 ;
        RECT 167.250 461.400 171.300 462.750 ;
        RECT 172.200 461.700 175.050 463.500 ;
        RECT 172.950 461.400 175.050 461.700 ;
        RECT 177.150 461.700 180.000 463.500 ;
        RECT 181.950 463.500 183.750 467.250 ;
        RECT 184.950 463.500 186.750 467.250 ;
        RECT 187.950 463.500 189.750 467.250 ;
        RECT 177.150 461.400 179.250 461.700 ;
        RECT 181.950 461.400 184.050 463.500 ;
        RECT 184.950 461.400 187.050 463.500 ;
        RECT 187.950 461.400 190.050 463.500 ;
        RECT 192.600 462.600 194.400 467.250 ;
        RECT 192.600 461.400 196.800 462.600 ;
        RECT 198.150 461.400 199.950 467.250 ;
        RECT 203.550 461.400 205.350 467.250 ;
        RECT 147.900 458.700 149.700 459.300 ;
        RECT 157.950 457.800 159.000 460.950 ;
        RECT 167.250 460.050 168.150 461.400 ;
        RECT 163.050 459.900 168.150 460.050 ;
        RECT 143.700 456.900 159.000 457.800 ;
        RECT 160.500 459.150 168.150 459.900 ;
        RECT 160.500 458.700 164.850 459.150 ;
        RECT 176.100 458.700 183.000 460.500 ;
        RECT 183.900 458.700 190.650 460.500 ;
        RECT 134.100 454.050 135.900 455.850 ;
        RECT 136.950 454.050 139.050 456.150 ;
        RECT 95.100 451.050 96.900 452.850 ;
        RECT 103.950 449.850 106.050 451.950 ;
        RECT 109.950 449.850 112.050 451.950 ;
        RECT 112.950 451.050 115.050 453.150 ;
        RECT 75.000 447.600 77.550 448.650 ;
        RECT 35.550 435.750 37.350 441.600 ;
        RECT 38.550 435.750 40.350 441.600 ;
        RECT 42.150 435.750 43.950 447.600 ;
        RECT 45.150 435.750 46.950 447.600 ;
        RECT 56.400 435.750 58.200 441.600 ;
        RECT 59.700 435.750 61.500 447.600 ;
        RECT 63.900 435.750 65.700 447.600 ;
        RECT 71.550 435.750 73.350 447.600 ;
        RECT 75.750 435.750 77.550 447.600 ;
        RECT 90.450 447.600 93.000 448.650 ;
        RECT 104.100 448.050 105.900 449.850 ;
        RECT 90.450 435.750 92.250 447.600 ;
        RECT 94.650 435.750 96.450 447.600 ;
        RECT 106.950 446.850 109.050 448.950 ;
        RECT 110.250 448.050 112.050 449.850 ;
        RECT 107.100 445.050 108.900 446.850 ;
        RECT 113.700 442.800 114.750 451.050 ;
        RECT 107.700 441.900 114.750 442.800 ;
        RECT 107.700 441.600 109.350 441.900 ;
        RECT 104.550 435.750 106.350 441.600 ;
        RECT 107.550 435.750 109.350 441.600 ;
        RECT 113.550 441.600 114.750 441.900 ;
        RECT 125.400 441.600 126.600 454.050 ;
        RECT 137.400 441.600 138.600 454.050 ;
        RECT 143.700 443.400 144.900 456.900 ;
        RECT 146.100 454.950 157.950 456.000 ;
        RECT 160.500 455.250 161.550 458.700 ;
        RECT 163.050 458.250 164.850 458.700 ;
        RECT 169.950 457.650 172.050 457.950 ;
        RECT 181.950 457.800 183.000 458.700 ;
        RECT 195.300 457.800 196.800 461.400 ;
        RECT 168.150 455.850 172.050 457.650 ;
        RECT 173.400 456.450 181.050 457.800 ;
        RECT 181.950 456.750 191.850 457.800 ;
        RECT 146.100 453.150 147.900 454.950 ;
        RECT 145.950 451.050 148.050 453.150 ;
        RECT 156.750 452.550 157.950 454.950 ;
        RECT 159.750 453.450 161.550 455.250 ;
        RECT 173.400 454.950 174.450 456.450 ;
        RECT 180.150 455.700 181.050 456.450 ;
        RECT 162.450 454.050 174.450 454.950 ;
        RECT 162.450 452.550 163.500 454.050 ;
        RECT 175.350 453.750 179.250 455.550 ;
        RECT 180.150 454.650 189.750 455.700 ;
        RECT 177.150 453.450 179.250 453.750 ;
        RECT 151.950 451.650 154.050 451.950 ;
        RECT 156.750 451.650 163.500 452.550 ;
        RECT 164.400 452.550 166.200 453.150 ;
        RECT 172.950 452.550 175.050 452.850 ;
        RECT 164.400 451.950 175.050 452.550 ;
        RECT 185.700 451.950 187.500 453.750 ;
        RECT 151.950 450.450 155.850 451.650 ;
        RECT 164.400 451.350 187.500 451.950 ;
        RECT 172.950 450.750 187.500 451.350 ;
        RECT 188.850 453.000 189.750 454.650 ;
        RECT 190.800 454.950 191.850 456.750 ;
        RECT 195.300 456.000 203.100 457.800 ;
        RECT 190.800 453.900 199.050 454.950 ;
        RECT 188.850 451.200 195.900 453.000 ;
        RECT 151.950 449.850 165.900 450.450 ;
        RECT 196.950 449.850 199.050 453.900 ;
        RECT 152.250 449.550 192.000 449.850 ;
        RECT 163.950 448.650 192.000 449.550 ;
        RECT 201.450 448.650 203.250 449.250 ;
        RECT 151.500 448.050 153.300 448.650 ;
        RECT 160.950 448.050 163.050 448.350 ;
        RECT 151.500 446.850 163.050 448.050 ;
        RECT 160.950 446.250 163.050 446.850 ;
        RECT 163.950 446.400 184.050 447.750 ;
        RECT 148.200 445.350 150.000 446.100 ;
        RECT 163.950 445.350 165.900 446.400 ;
        RECT 181.950 445.650 184.050 446.400 ;
        RECT 187.950 446.550 190.050 447.750 ;
        RECT 190.950 447.450 203.250 448.650 ;
        RECT 204.150 446.550 205.350 461.400 ;
        RECT 187.950 445.650 205.350 446.550 ;
        RECT 207.450 464.400 209.250 467.250 ;
        RECT 210.450 464.400 212.250 467.250 ;
        RECT 207.450 456.150 208.950 464.400 ;
        RECT 223.650 461.400 225.450 467.250 ;
        RECT 224.250 459.300 225.450 461.400 ;
        RECT 226.650 462.300 228.450 467.250 ;
        RECT 229.650 463.200 231.450 467.250 ;
        RECT 232.650 462.300 234.450 467.250 ;
        RECT 226.650 460.950 234.450 462.300 ;
        RECT 241.650 461.400 243.450 467.250 ;
        RECT 242.250 459.300 243.450 461.400 ;
        RECT 244.650 462.300 246.450 467.250 ;
        RECT 247.650 463.200 249.450 467.250 ;
        RECT 250.650 462.300 252.450 467.250 ;
        RECT 259.650 464.400 261.450 467.250 ;
        RECT 262.650 464.400 264.450 467.250 ;
        RECT 265.650 464.400 267.450 467.250 ;
        RECT 244.650 460.950 252.450 462.300 ;
        RECT 224.250 458.250 228.000 459.300 ;
        RECT 242.250 458.250 246.000 459.300 ;
        RECT 207.450 454.050 211.050 456.150 ;
        RECT 226.950 454.950 228.150 458.250 ;
        RECT 230.100 456.150 231.900 457.950 ;
        RECT 148.200 444.300 165.900 445.350 ;
        RECT 143.700 442.500 147.750 443.400 ;
        RECT 146.700 441.600 147.750 442.500 ;
        RECT 110.550 435.750 112.350 441.000 ;
        RECT 113.550 435.750 115.350 441.600 ;
        RECT 122.550 435.750 124.350 441.600 ;
        RECT 125.550 435.750 127.350 441.600 ;
        RECT 134.550 435.750 136.350 441.600 ;
        RECT 137.550 435.750 139.350 441.600 ;
        RECT 143.700 435.750 145.500 441.600 ;
        RECT 146.700 435.750 148.500 441.600 ;
        RECT 149.700 435.750 151.500 441.600 ;
        RECT 152.700 435.750 154.500 444.300 ;
        RECT 172.950 444.150 175.050 444.600 ;
        RECT 172.650 442.500 175.050 444.150 ;
        RECT 177.000 442.800 180.900 444.600 ;
        RECT 177.000 442.500 180.000 442.800 ;
        RECT 157.950 439.950 160.050 442.050 ;
        RECT 160.950 439.950 163.050 442.050 ;
        RECT 163.950 441.600 166.050 442.050 ;
        RECT 172.650 441.600 174.000 442.500 ;
        RECT 163.950 439.950 166.500 441.600 ;
        RECT 155.700 435.750 157.500 439.050 ;
        RECT 158.850 438.600 160.050 439.950 ;
        RECT 162.150 438.600 163.050 439.950 ;
        RECT 165.300 438.600 166.500 439.950 ;
        RECT 158.850 435.750 161.250 438.600 ;
        RECT 162.150 435.750 164.250 438.600 ;
        RECT 165.300 435.750 167.250 438.600 ;
        RECT 168.450 435.750 170.250 441.600 ;
        RECT 172.200 435.750 174.000 441.600 ;
        RECT 175.200 435.750 177.000 441.600 ;
        RECT 178.200 435.750 180.000 442.500 ;
        RECT 182.100 438.600 183.450 445.650 ;
        RECT 191.850 444.150 193.650 444.300 ;
        RECT 184.950 442.950 193.650 444.150 ;
        RECT 198.600 443.700 200.400 444.300 ;
        RECT 184.950 442.050 187.050 442.950 ;
        RECT 191.850 442.500 193.650 442.950 ;
        RECT 194.700 442.500 200.400 443.700 ;
        RECT 181.950 435.750 183.750 438.600 ;
        RECT 184.950 435.750 186.750 442.050 ;
        RECT 188.100 439.800 190.200 441.900 ;
        RECT 188.100 438.600 189.600 439.800 ;
        RECT 187.950 435.750 189.750 438.600 ;
        RECT 191.700 435.750 193.500 441.600 ;
        RECT 194.700 435.750 196.500 442.500 ;
        RECT 201.300 441.600 202.500 445.650 ;
        RECT 207.450 441.600 208.950 454.050 ;
        RECT 226.950 452.850 229.050 454.950 ;
        RECT 229.950 454.050 232.050 456.150 ;
        RECT 244.950 454.950 246.150 458.250 ;
        RECT 262.950 457.950 264.000 464.400 ;
        RECT 272.550 459.900 274.350 467.250 ;
        RECT 277.050 461.400 278.850 467.250 ;
        RECT 280.050 462.900 281.850 467.250 ;
        RECT 280.050 461.400 283.350 462.900 ;
        RECT 278.250 459.900 280.050 460.500 ;
        RECT 272.550 458.700 280.050 459.900 ;
        RECT 248.100 456.150 249.900 457.950 ;
        RECT 232.950 452.850 235.050 454.950 ;
        RECT 244.950 452.850 247.050 454.950 ;
        RECT 247.950 454.050 250.050 456.150 ;
        RECT 262.950 455.850 265.050 457.950 ;
        RECT 250.950 452.850 253.050 454.950 ;
        RECT 259.950 452.850 262.050 454.950 ;
        RECT 223.950 449.850 226.050 451.950 ;
        RECT 224.250 448.050 226.050 449.850 ;
        RECT 227.850 447.600 229.050 452.850 ;
        RECT 233.100 451.050 234.900 452.850 ;
        RECT 241.950 449.850 244.050 451.950 ;
        RECT 242.250 448.050 244.050 449.850 ;
        RECT 245.850 447.600 247.050 452.850 ;
        RECT 251.100 451.050 252.900 452.850 ;
        RECT 260.100 451.050 261.900 452.850 ;
        RECT 262.950 448.650 264.000 455.850 ;
        RECT 265.950 452.850 268.050 454.950 ;
        RECT 271.950 452.850 274.050 454.950 ;
        RECT 266.100 451.050 267.900 452.850 ;
        RECT 272.100 451.050 273.900 452.850 ;
        RECT 261.450 447.600 264.000 448.650 ;
        RECT 197.700 435.750 199.500 441.600 ;
        RECT 200.700 435.750 202.500 441.600 ;
        RECT 203.700 435.750 205.500 441.600 ;
        RECT 207.450 435.750 209.250 441.600 ;
        RECT 210.450 435.750 212.250 441.600 ;
        RECT 224.400 435.750 226.200 441.600 ;
        RECT 227.700 435.750 229.500 447.600 ;
        RECT 231.900 435.750 233.700 447.600 ;
        RECT 242.400 435.750 244.200 441.600 ;
        RECT 245.700 435.750 247.500 447.600 ;
        RECT 249.900 435.750 251.700 447.600 ;
        RECT 261.450 435.750 263.250 447.600 ;
        RECT 265.650 435.750 267.450 447.600 ;
        RECT 275.700 441.600 276.900 458.700 ;
        RECT 282.150 454.950 283.350 461.400 ;
        RECT 290.700 458.400 292.500 467.250 ;
        RECT 296.100 459.000 297.900 467.250 ;
        RECT 296.100 457.350 300.600 459.000 ;
        RECT 311.700 458.400 313.500 467.250 ;
        RECT 317.100 459.000 318.900 467.250 ;
        RECT 332.850 460.200 334.650 467.250 ;
        RECT 337.350 461.400 339.150 467.250 ;
        RECT 317.100 457.350 321.600 459.000 ;
        RECT 328.950 457.950 331.050 460.050 ;
        RECT 332.850 459.300 336.450 460.200 ;
        RECT 278.100 453.150 279.900 454.950 ;
        RECT 277.950 451.050 280.050 453.150 ;
        RECT 280.950 452.850 283.350 454.950 ;
        RECT 299.400 453.150 300.600 457.350 ;
        RECT 313.950 456.450 316.050 457.050 ;
        RECT 308.550 455.550 316.050 456.450 ;
        RECT 282.150 447.600 283.350 452.850 ;
        RECT 289.950 449.850 292.050 451.950 ;
        RECT 295.950 449.850 298.050 451.950 ;
        RECT 298.950 451.050 301.050 453.150 ;
        RECT 290.100 448.050 291.900 449.850 ;
        RECT 272.550 435.750 274.350 441.600 ;
        RECT 275.550 435.750 277.350 441.600 ;
        RECT 279.150 435.750 280.950 447.600 ;
        RECT 282.150 435.750 283.950 447.600 ;
        RECT 292.950 446.850 295.050 448.950 ;
        RECT 296.250 448.050 298.050 449.850 ;
        RECT 293.100 445.050 294.900 446.850 ;
        RECT 299.700 442.800 300.750 451.050 ;
        RECT 308.550 448.050 309.450 455.550 ;
        RECT 313.950 454.950 316.050 455.550 ;
        RECT 320.400 453.150 321.600 457.350 ;
        RECT 310.950 449.850 313.050 451.950 ;
        RECT 316.950 449.850 319.050 451.950 ;
        RECT 319.950 451.050 322.050 453.150 ;
        RECT 311.100 448.050 312.900 449.850 ;
        RECT 307.950 445.950 310.050 448.050 ;
        RECT 313.950 446.850 316.050 448.950 ;
        RECT 317.250 448.050 319.050 449.850 ;
        RECT 314.100 445.050 315.900 446.850 ;
        RECT 320.700 442.800 321.750 451.050 ;
        RECT 329.550 447.450 330.450 457.950 ;
        RECT 332.100 453.150 333.900 454.950 ;
        RECT 331.950 451.050 334.050 453.150 ;
        RECT 335.250 451.950 336.450 459.300 ;
        RECT 347.100 459.000 348.900 467.250 ;
        RECT 344.400 457.350 348.900 459.000 ;
        RECT 352.500 458.400 354.300 467.250 ;
        RECT 362.550 462.300 364.350 467.250 ;
        RECT 365.550 463.200 367.350 467.250 ;
        RECT 368.550 462.300 370.350 467.250 ;
        RECT 362.550 460.950 370.350 462.300 ;
        RECT 371.550 461.400 373.350 467.250 ;
        RECT 379.650 464.400 381.450 467.250 ;
        RECT 382.650 464.400 384.450 467.250 ;
        RECT 394.650 464.400 396.450 467.250 ;
        RECT 397.650 464.400 399.450 467.250 ;
        RECT 400.650 464.400 402.450 467.250 ;
        RECT 407.250 464.400 409.350 467.250 ;
        RECT 410.550 464.400 412.350 467.250 ;
        RECT 413.550 464.400 415.350 467.250 ;
        RECT 416.550 464.400 418.350 467.250 ;
        RECT 431.550 464.400 433.350 467.250 ;
        RECT 434.550 464.400 436.350 467.250 ;
        RECT 371.550 459.300 372.750 461.400 ;
        RECT 369.000 458.250 372.750 459.300 ;
        RECT 338.100 453.150 339.900 454.950 ;
        RECT 344.400 453.150 345.600 457.350 ;
        RECT 365.100 456.150 366.900 457.950 ;
        RECT 334.950 449.850 337.050 451.950 ;
        RECT 337.950 451.050 340.050 453.150 ;
        RECT 343.950 451.050 346.050 453.150 ;
        RECT 361.950 452.850 364.050 454.950 ;
        RECT 364.950 454.050 367.050 456.150 ;
        RECT 368.850 454.950 370.050 458.250 ;
        RECT 380.400 456.150 381.600 464.400 ;
        RECT 394.950 459.450 397.050 460.050 ;
        RECT 392.550 458.550 397.050 459.450 ;
        RECT 367.950 452.850 370.050 454.950 ;
        RECT 379.950 454.050 382.050 456.150 ;
        RECT 382.950 455.850 385.050 457.950 ;
        RECT 383.100 454.050 384.900 455.850 ;
        RECT 331.950 447.450 334.050 448.050 ;
        RECT 329.550 446.550 334.050 447.450 ;
        RECT 331.950 445.950 334.050 446.550 ;
        RECT 293.700 441.900 300.750 442.800 ;
        RECT 293.700 441.600 295.350 441.900 ;
        RECT 290.550 435.750 292.350 441.600 ;
        RECT 293.550 435.750 295.350 441.600 ;
        RECT 299.550 441.600 300.750 441.900 ;
        RECT 314.700 441.900 321.750 442.800 ;
        RECT 314.700 441.600 316.350 441.900 ;
        RECT 296.550 435.750 298.350 441.000 ;
        RECT 299.550 435.750 301.350 441.600 ;
        RECT 311.550 435.750 313.350 441.600 ;
        RECT 314.550 435.750 316.350 441.600 ;
        RECT 320.550 441.600 321.750 441.900 ;
        RECT 335.250 441.600 336.450 449.850 ;
        RECT 344.250 442.800 345.300 451.050 ;
        RECT 346.950 449.850 349.050 451.950 ;
        RECT 352.950 449.850 355.050 451.950 ;
        RECT 362.100 451.050 363.900 452.850 ;
        RECT 346.950 448.050 348.750 449.850 ;
        RECT 349.950 446.850 352.050 448.950 ;
        RECT 353.100 448.050 354.900 449.850 ;
        RECT 367.950 447.600 369.150 452.850 ;
        RECT 370.950 449.850 373.050 451.950 ;
        RECT 370.950 448.050 372.750 449.850 ;
        RECT 350.100 445.050 351.900 446.850 ;
        RECT 344.250 441.900 351.300 442.800 ;
        RECT 344.250 441.600 345.450 441.900 ;
        RECT 317.550 435.750 319.350 441.000 ;
        RECT 320.550 435.750 322.350 441.600 ;
        RECT 331.650 435.750 333.450 441.600 ;
        RECT 334.650 435.750 336.450 441.600 ;
        RECT 337.650 435.750 339.450 441.600 ;
        RECT 343.650 435.750 345.450 441.600 ;
        RECT 349.650 441.600 351.300 441.900 ;
        RECT 346.650 435.750 348.450 441.000 ;
        RECT 349.650 435.750 351.450 441.600 ;
        RECT 352.650 435.750 354.450 441.600 ;
        RECT 363.300 435.750 365.100 447.600 ;
        RECT 367.500 435.750 369.300 447.600 ;
        RECT 380.400 441.600 381.600 454.050 ;
        RECT 385.950 453.450 388.050 454.050 ;
        RECT 392.550 453.450 393.450 458.550 ;
        RECT 394.950 457.950 397.050 458.550 ;
        RECT 397.950 457.950 399.000 464.400 ;
        RECT 411.300 463.500 412.350 464.400 ;
        RECT 417.300 463.500 418.350 464.400 ;
        RECT 411.300 462.600 422.100 463.500 ;
        RECT 397.950 455.850 400.050 457.950 ;
        RECT 413.100 456.150 414.900 457.950 ;
        RECT 420.900 456.150 422.100 462.600 ;
        RECT 385.950 452.550 393.450 453.450 ;
        RECT 394.950 452.850 397.050 454.950 ;
        RECT 385.950 451.950 388.050 452.550 ;
        RECT 395.100 451.050 396.900 452.850 ;
        RECT 397.950 448.650 399.000 455.850 ;
        RECT 400.950 452.850 403.050 454.950 ;
        RECT 406.950 452.850 409.050 454.950 ;
        RECT 412.950 454.050 415.050 456.150 ;
        RECT 415.950 452.850 418.050 454.950 ;
        RECT 420.900 454.050 424.050 456.150 ;
        RECT 430.950 455.850 433.050 457.950 ;
        RECT 434.400 456.150 435.600 464.400 ;
        RECT 442.650 461.400 444.450 467.250 ;
        RECT 443.250 459.300 444.450 461.400 ;
        RECT 445.650 462.300 447.450 467.250 ;
        RECT 448.650 463.200 450.450 467.250 ;
        RECT 451.650 462.300 453.450 467.250 ;
        RECT 445.650 460.950 453.450 462.300 ;
        RECT 455.550 462.300 457.350 467.250 ;
        RECT 458.550 463.200 460.350 467.250 ;
        RECT 461.550 462.300 463.350 467.250 ;
        RECT 455.550 460.950 463.350 462.300 ;
        RECT 464.550 461.400 466.350 467.250 ;
        RECT 476.550 464.400 478.350 467.250 ;
        RECT 479.550 464.400 481.350 467.250 ;
        RECT 475.950 462.450 478.050 463.050 ;
        RECT 473.550 461.550 478.050 462.450 ;
        RECT 464.550 459.300 465.750 461.400 ;
        RECT 443.250 458.250 447.000 459.300 ;
        RECT 462.000 458.250 465.750 459.300 ;
        RECT 431.100 454.050 432.900 455.850 ;
        RECT 433.950 454.050 436.050 456.150 ;
        RECT 445.950 454.950 447.150 458.250 ;
        RECT 449.100 456.150 450.900 457.950 ;
        RECT 458.100 456.150 459.900 457.950 ;
        RECT 401.100 451.050 402.900 452.850 ;
        RECT 407.100 451.050 408.900 452.850 ;
        RECT 416.100 451.050 417.900 452.850 ;
        RECT 396.450 447.600 399.000 448.650 ;
        RECT 420.900 448.800 422.100 454.050 ;
        RECT 420.900 447.600 424.350 448.800 ;
        RECT 370.800 435.750 372.600 441.600 ;
        RECT 379.650 435.750 381.450 441.600 ;
        RECT 382.650 435.750 384.450 441.600 ;
        RECT 396.450 435.750 398.250 447.600 ;
        RECT 400.650 435.750 402.450 447.600 ;
        RECT 404.550 445.500 412.350 446.400 ;
        RECT 404.550 435.750 406.350 445.500 ;
        RECT 407.550 435.750 409.350 444.600 ;
        RECT 410.550 436.500 412.350 445.500 ;
        RECT 413.550 445.200 421.950 446.100 ;
        RECT 413.550 437.400 415.350 445.200 ;
        RECT 416.550 436.500 418.350 444.300 ;
        RECT 410.550 435.750 418.350 436.500 ;
        RECT 420.150 436.500 421.950 445.200 ;
        RECT 423.150 445.200 424.350 447.600 ;
        RECT 423.150 437.400 424.950 445.200 ;
        RECT 426.150 436.500 427.950 445.800 ;
        RECT 434.400 441.600 435.600 454.050 ;
        RECT 445.950 452.850 448.050 454.950 ;
        RECT 448.950 454.050 451.050 456.150 ;
        RECT 451.950 452.850 454.050 454.950 ;
        RECT 454.950 452.850 457.050 454.950 ;
        RECT 457.950 454.050 460.050 456.150 ;
        RECT 461.850 454.950 463.050 458.250 ;
        RECT 460.950 452.850 463.050 454.950 ;
        RECT 442.950 449.850 445.050 451.950 ;
        RECT 443.250 448.050 445.050 449.850 ;
        RECT 446.850 447.600 448.050 452.850 ;
        RECT 452.100 451.050 453.900 452.850 ;
        RECT 455.100 451.050 456.900 452.850 ;
        RECT 460.950 447.600 462.150 452.850 ;
        RECT 463.950 449.850 466.050 451.950 ;
        RECT 473.550 450.450 474.450 461.550 ;
        RECT 475.950 460.950 478.050 461.550 ;
        RECT 475.950 455.850 478.050 457.950 ;
        RECT 479.400 456.150 480.600 464.400 ;
        RECT 485.700 458.400 487.500 467.250 ;
        RECT 491.100 459.000 492.900 467.250 ;
        RECT 491.100 457.350 495.600 459.000 ;
        RECT 496.950 457.950 499.050 460.050 ;
        RECT 506.700 458.400 508.500 467.250 ;
        RECT 512.100 459.000 513.900 467.250 ;
        RECT 487.950 456.450 490.050 457.050 ;
        RECT 476.100 454.050 477.900 455.850 ;
        RECT 478.950 454.050 481.050 456.150 ;
        RECT 482.550 455.550 490.050 456.450 ;
        RECT 475.950 450.450 478.050 451.050 ;
        RECT 463.950 448.050 465.750 449.850 ;
        RECT 473.550 449.550 478.050 450.450 ;
        RECT 475.950 448.950 478.050 449.550 ;
        RECT 420.150 435.750 427.950 436.500 ;
        RECT 431.550 435.750 433.350 441.600 ;
        RECT 434.550 435.750 436.350 441.600 ;
        RECT 443.400 435.750 445.200 441.600 ;
        RECT 446.700 435.750 448.500 447.600 ;
        RECT 450.900 435.750 452.700 447.600 ;
        RECT 456.300 435.750 458.100 447.600 ;
        RECT 460.500 435.750 462.300 447.600 ;
        RECT 479.400 441.600 480.600 454.050 ;
        RECT 482.550 444.450 483.450 455.550 ;
        RECT 487.950 454.950 490.050 455.550 ;
        RECT 494.400 453.150 495.600 457.350 ;
        RECT 484.950 449.850 487.050 451.950 ;
        RECT 490.950 449.850 493.050 451.950 ;
        RECT 493.950 451.050 496.050 453.150 ;
        RECT 485.100 448.050 486.900 449.850 ;
        RECT 487.950 446.850 490.050 448.950 ;
        RECT 491.250 448.050 493.050 449.850 ;
        RECT 488.100 445.050 489.900 446.850 ;
        RECT 484.950 444.450 487.050 445.050 ;
        RECT 482.550 443.550 487.050 444.450 ;
        RECT 484.950 442.950 487.050 443.550 ;
        RECT 494.700 442.800 495.750 451.050 ;
        RECT 497.550 447.450 498.450 457.950 ;
        RECT 512.100 457.350 516.600 459.000 ;
        RECT 527.700 458.400 529.500 467.250 ;
        RECT 533.100 459.000 534.900 467.250 ;
        RECT 550.650 464.400 552.450 467.250 ;
        RECT 553.650 464.400 555.450 467.250 ;
        RECT 558.750 464.400 560.550 467.250 ;
        RECT 561.750 464.400 563.550 467.250 ;
        RECT 533.100 457.350 537.600 459.000 ;
        RECT 502.950 454.950 505.050 457.050 ;
        RECT 499.950 453.450 502.050 454.050 ;
        RECT 503.550 453.450 504.450 454.950 ;
        RECT 499.950 452.550 504.450 453.450 ;
        RECT 515.400 453.150 516.600 457.350 ;
        RECT 523.950 456.450 526.050 457.050 ;
        RECT 529.950 456.450 532.050 457.050 ;
        RECT 523.950 455.550 532.050 456.450 ;
        RECT 523.950 454.950 526.050 455.550 ;
        RECT 529.950 454.950 532.050 455.550 ;
        RECT 536.400 453.150 537.600 457.350 ;
        RECT 551.400 456.150 552.600 464.400 ;
        RECT 550.950 454.050 553.050 456.150 ;
        RECT 553.950 455.850 556.050 457.950 ;
        RECT 562.050 456.150 563.550 464.400 ;
        RECT 554.100 454.050 555.900 455.850 ;
        RECT 559.950 454.050 563.550 456.150 ;
        RECT 499.950 451.950 502.050 452.550 ;
        RECT 505.950 449.850 508.050 451.950 ;
        RECT 511.950 449.850 514.050 451.950 ;
        RECT 514.950 451.050 517.050 453.150 ;
        RECT 506.100 448.050 507.900 449.850 ;
        RECT 502.950 447.450 505.050 448.050 ;
        RECT 497.550 446.550 505.050 447.450 ;
        RECT 508.950 446.850 511.050 448.950 ;
        RECT 512.250 448.050 514.050 449.850 ;
        RECT 502.950 445.950 505.050 446.550 ;
        RECT 509.100 445.050 510.900 446.850 ;
        RECT 515.700 442.800 516.750 451.050 ;
        RECT 526.950 449.850 529.050 451.950 ;
        RECT 532.950 449.850 535.050 451.950 ;
        RECT 535.950 451.050 538.050 453.150 ;
        RECT 527.100 448.050 528.900 449.850 ;
        RECT 529.950 446.850 532.050 448.950 ;
        RECT 533.250 448.050 535.050 449.850 ;
        RECT 530.100 445.050 531.900 446.850 ;
        RECT 536.700 442.800 537.750 451.050 ;
        RECT 488.700 441.900 495.750 442.800 ;
        RECT 488.700 441.600 490.350 441.900 ;
        RECT 463.800 435.750 465.600 441.600 ;
        RECT 476.550 435.750 478.350 441.600 ;
        RECT 479.550 435.750 481.350 441.600 ;
        RECT 485.550 435.750 487.350 441.600 ;
        RECT 488.550 435.750 490.350 441.600 ;
        RECT 494.550 441.600 495.750 441.900 ;
        RECT 509.700 441.900 516.750 442.800 ;
        RECT 509.700 441.600 511.350 441.900 ;
        RECT 491.550 435.750 493.350 441.000 ;
        RECT 494.550 435.750 496.350 441.600 ;
        RECT 506.550 435.750 508.350 441.600 ;
        RECT 509.550 435.750 511.350 441.600 ;
        RECT 515.550 441.600 516.750 441.900 ;
        RECT 530.700 441.900 537.750 442.800 ;
        RECT 530.700 441.600 532.350 441.900 ;
        RECT 512.550 435.750 514.350 441.000 ;
        RECT 515.550 435.750 517.350 441.600 ;
        RECT 527.550 435.750 529.350 441.600 ;
        RECT 530.550 435.750 532.350 441.600 ;
        RECT 536.550 441.600 537.750 441.900 ;
        RECT 551.400 441.600 552.600 454.050 ;
        RECT 562.050 441.600 563.550 454.050 ;
        RECT 565.650 461.400 567.450 467.250 ;
        RECT 571.050 461.400 572.850 467.250 ;
        RECT 576.600 462.600 578.400 467.250 ;
        RECT 581.250 463.500 583.050 467.250 ;
        RECT 584.250 463.500 586.050 467.250 ;
        RECT 587.250 463.500 589.050 467.250 ;
        RECT 574.200 461.400 578.400 462.600 ;
        RECT 580.950 461.400 583.050 463.500 ;
        RECT 583.950 461.400 586.050 463.500 ;
        RECT 586.950 461.400 589.050 463.500 ;
        RECT 591.000 463.500 592.800 467.250 ;
        RECT 594.000 464.400 595.800 467.250 ;
        RECT 597.000 463.500 598.800 467.250 ;
        RECT 601.500 464.400 603.300 467.250 ;
        RECT 604.500 464.400 606.300 467.250 ;
        RECT 607.500 464.400 609.300 467.250 ;
        RECT 610.500 464.400 612.300 467.250 ;
        RECT 591.000 461.700 593.850 463.500 ;
        RECT 591.750 461.400 593.850 461.700 ;
        RECT 595.950 461.700 598.800 463.500 ;
        RECT 599.700 462.750 601.500 463.200 ;
        RECT 604.950 463.050 606.300 464.400 ;
        RECT 607.950 463.050 609.300 464.400 ;
        RECT 610.950 463.050 612.300 464.400 ;
        RECT 595.950 461.400 598.050 461.700 ;
        RECT 599.700 461.400 603.750 462.750 ;
        RECT 565.650 446.550 566.850 461.400 ;
        RECT 574.200 457.800 575.700 461.400 ;
        RECT 580.350 458.700 587.100 460.500 ;
        RECT 588.000 458.700 594.900 460.500 ;
        RECT 602.850 460.050 603.750 461.400 ;
        RECT 604.950 460.950 607.050 463.050 ;
        RECT 607.950 460.950 610.050 463.050 ;
        RECT 610.950 460.950 613.050 463.050 ;
        RECT 602.850 459.900 607.950 460.050 ;
        RECT 602.850 459.150 610.500 459.900 ;
        RECT 606.150 458.700 610.500 459.150 ;
        RECT 588.000 457.800 589.050 458.700 ;
        RECT 606.150 458.250 607.950 458.700 ;
        RECT 567.900 456.000 575.700 457.800 ;
        RECT 579.150 456.750 589.050 457.800 ;
        RECT 579.150 454.950 580.200 456.750 ;
        RECT 589.950 456.450 597.600 457.800 ;
        RECT 589.950 455.700 590.850 456.450 ;
        RECT 571.950 453.900 580.200 454.950 ;
        RECT 581.250 454.650 590.850 455.700 ;
        RECT 571.950 449.850 574.050 453.900 ;
        RECT 581.250 453.000 582.150 454.650 ;
        RECT 591.750 453.750 595.650 455.550 ;
        RECT 596.550 454.950 597.600 456.450 ;
        RECT 598.950 457.650 601.050 457.950 ;
        RECT 598.950 455.850 602.850 457.650 ;
        RECT 609.450 455.250 610.500 458.700 ;
        RECT 612.000 457.800 613.050 460.950 ;
        RECT 614.700 461.400 616.500 467.250 ;
        RECT 620.100 461.400 621.900 467.250 ;
        RECT 625.500 461.400 627.300 467.250 ;
        RECT 632.550 464.400 634.350 467.250 ;
        RECT 635.550 464.400 637.350 467.250 ;
        RECT 614.700 460.500 616.200 461.400 ;
        RECT 614.700 459.300 623.100 460.500 ;
        RECT 621.300 458.700 623.100 459.300 ;
        RECT 626.100 457.800 627.300 461.400 ;
        RECT 612.000 456.900 627.300 457.800 ;
        RECT 596.550 454.050 608.550 454.950 ;
        RECT 575.100 451.200 582.150 453.000 ;
        RECT 583.500 451.950 585.300 453.750 ;
        RECT 591.750 453.450 593.850 453.750 ;
        RECT 595.950 452.550 598.050 452.850 ;
        RECT 604.800 452.550 606.600 453.150 ;
        RECT 595.950 451.950 606.600 452.550 ;
        RECT 583.500 451.350 606.600 451.950 ;
        RECT 607.500 452.550 608.550 454.050 ;
        RECT 609.450 453.450 611.250 455.250 ;
        RECT 613.050 454.950 624.900 456.000 ;
        RECT 613.050 452.550 614.250 454.950 ;
        RECT 623.100 453.150 624.900 454.950 ;
        RECT 607.500 451.650 614.250 452.550 ;
        RECT 616.950 451.650 619.050 451.950 ;
        RECT 583.500 450.750 598.050 451.350 ;
        RECT 615.150 450.450 619.050 451.650 ;
        RECT 622.950 451.050 625.050 453.150 ;
        RECT 605.100 449.850 619.050 450.450 ;
        RECT 579.000 449.550 618.750 449.850 ;
        RECT 567.750 448.650 569.550 449.250 ;
        RECT 579.000 448.650 607.050 449.550 ;
        RECT 567.750 447.450 580.050 448.650 ;
        RECT 607.950 448.050 610.050 448.350 ;
        RECT 617.700 448.050 619.500 448.650 ;
        RECT 580.950 446.550 583.050 447.750 ;
        RECT 565.650 445.650 583.050 446.550 ;
        RECT 586.950 446.400 607.050 447.750 ;
        RECT 586.950 445.650 589.050 446.400 ;
        RECT 568.500 441.600 569.700 445.650 ;
        RECT 570.600 443.700 572.400 444.300 ;
        RECT 577.350 444.150 579.150 444.300 ;
        RECT 570.600 442.500 576.300 443.700 ;
        RECT 577.350 442.950 586.050 444.150 ;
        RECT 577.350 442.500 579.150 442.950 ;
        RECT 533.550 435.750 535.350 441.000 ;
        RECT 536.550 435.750 538.350 441.600 ;
        RECT 550.650 435.750 552.450 441.600 ;
        RECT 553.650 435.750 555.450 441.600 ;
        RECT 558.750 435.750 560.550 441.600 ;
        RECT 561.750 435.750 563.550 441.600 ;
        RECT 565.500 435.750 567.300 441.600 ;
        RECT 568.500 435.750 570.300 441.600 ;
        RECT 571.500 435.750 573.300 441.600 ;
        RECT 574.500 435.750 576.300 442.500 ;
        RECT 583.950 442.050 586.050 442.950 ;
        RECT 577.500 435.750 579.300 441.600 ;
        RECT 580.800 439.800 582.900 441.900 ;
        RECT 581.400 438.600 582.900 439.800 ;
        RECT 581.250 435.750 583.050 438.600 ;
        RECT 584.250 435.750 586.050 442.050 ;
        RECT 587.550 438.600 588.900 445.650 ;
        RECT 605.100 445.350 607.050 446.400 ;
        RECT 607.950 446.850 619.500 448.050 ;
        RECT 607.950 446.250 610.050 446.850 ;
        RECT 621.000 445.350 622.800 446.100 ;
        RECT 590.100 442.800 594.000 444.600 ;
        RECT 591.000 442.500 594.000 442.800 ;
        RECT 595.950 444.150 598.050 444.600 ;
        RECT 605.100 444.300 622.800 445.350 ;
        RECT 595.950 442.500 598.350 444.150 ;
        RECT 587.250 435.750 589.050 438.600 ;
        RECT 591.000 435.750 592.800 442.500 ;
        RECT 597.000 441.600 598.350 442.500 ;
        RECT 604.950 441.600 607.050 442.050 ;
        RECT 594.000 435.750 595.800 441.600 ;
        RECT 597.000 435.750 598.800 441.600 ;
        RECT 600.750 435.750 602.550 441.600 ;
        RECT 604.500 439.950 607.050 441.600 ;
        RECT 607.950 439.950 610.050 442.050 ;
        RECT 610.950 439.950 613.050 442.050 ;
        RECT 604.500 438.600 605.700 439.950 ;
        RECT 607.950 438.600 608.850 439.950 ;
        RECT 610.950 438.600 612.150 439.950 ;
        RECT 603.750 435.750 605.700 438.600 ;
        RECT 606.750 435.750 608.850 438.600 ;
        RECT 609.750 435.750 612.150 438.600 ;
        RECT 613.500 435.750 615.300 439.050 ;
        RECT 616.500 435.750 618.300 444.300 ;
        RECT 626.100 443.400 627.300 456.900 ;
        RECT 631.950 455.850 634.050 457.950 ;
        RECT 635.400 456.150 636.600 464.400 ;
        RECT 647.550 462.300 649.350 467.250 ;
        RECT 650.550 463.200 652.350 467.250 ;
        RECT 653.550 462.300 655.350 467.250 ;
        RECT 647.550 460.950 655.350 462.300 ;
        RECT 656.550 461.400 658.350 467.250 ;
        RECT 668.550 462.300 670.350 467.250 ;
        RECT 671.550 463.200 673.350 467.250 ;
        RECT 674.550 462.300 676.350 467.250 ;
        RECT 656.550 459.300 657.750 461.400 ;
        RECT 668.550 460.950 676.350 462.300 ;
        RECT 677.550 461.400 679.350 467.250 ;
        RECT 686.550 462.300 688.350 467.250 ;
        RECT 689.550 463.200 691.350 467.250 ;
        RECT 692.550 462.300 694.350 467.250 ;
        RECT 677.550 459.300 678.750 461.400 ;
        RECT 686.550 460.950 694.350 462.300 ;
        RECT 695.550 461.400 697.350 467.250 ;
        RECT 695.550 459.300 696.750 461.400 ;
        RECT 654.000 458.250 657.750 459.300 ;
        RECT 675.000 458.250 678.750 459.300 ;
        RECT 693.000 458.250 696.750 459.300 ;
        RECT 710.100 459.000 711.900 467.250 ;
        RECT 650.100 456.150 651.900 457.950 ;
        RECT 632.100 454.050 633.900 455.850 ;
        RECT 634.950 454.050 637.050 456.150 ;
        RECT 623.250 442.500 627.300 443.400 ;
        RECT 623.250 441.600 624.300 442.500 ;
        RECT 635.400 441.600 636.600 454.050 ;
        RECT 646.950 452.850 649.050 454.950 ;
        RECT 649.950 454.050 652.050 456.150 ;
        RECT 653.850 454.950 655.050 458.250 ;
        RECT 671.100 456.150 672.900 457.950 ;
        RECT 652.950 452.850 655.050 454.950 ;
        RECT 667.950 452.850 670.050 454.950 ;
        RECT 670.950 454.050 673.050 456.150 ;
        RECT 674.850 454.950 676.050 458.250 ;
        RECT 689.100 456.150 690.900 457.950 ;
        RECT 673.950 452.850 676.050 454.950 ;
        RECT 685.950 452.850 688.050 454.950 ;
        RECT 688.950 454.050 691.050 456.150 ;
        RECT 692.850 454.950 694.050 458.250 ;
        RECT 707.400 457.350 711.900 459.000 ;
        RECT 715.500 458.400 717.300 467.250 ;
        RECT 724.650 461.400 726.450 467.250 ;
        RECT 727.650 464.400 729.450 467.250 ;
        RECT 730.650 464.400 732.450 467.250 ;
        RECT 733.650 464.400 735.450 467.250 ;
        RECT 694.950 456.450 697.050 457.050 ;
        RECT 703.950 456.450 706.050 457.050 ;
        RECT 694.950 455.550 706.050 456.450 ;
        RECT 694.950 454.950 697.050 455.550 ;
        RECT 703.950 454.950 706.050 455.550 ;
        RECT 691.950 452.850 694.050 454.950 ;
        RECT 707.400 453.150 708.600 457.350 ;
        RECT 724.950 456.150 726.000 461.400 ;
        RECT 730.650 460.200 731.550 464.400 ;
        RECT 728.250 459.300 731.550 460.200 ;
        RECT 743.850 460.200 745.650 467.250 ;
        RECT 748.350 461.400 750.150 467.250 ;
        RECT 758.850 460.200 760.650 467.250 ;
        RECT 763.350 461.400 765.150 467.250 ;
        RECT 769.650 464.400 771.450 467.250 ;
        RECT 772.650 464.400 774.450 467.250 ;
        RECT 777.750 464.400 779.550 467.250 ;
        RECT 780.750 464.400 782.550 467.250 ;
        RECT 743.850 459.300 747.450 460.200 ;
        RECT 758.850 459.300 762.450 460.200 ;
        RECT 728.250 458.400 730.050 459.300 ;
        RECT 724.950 454.050 727.050 456.150 ;
        RECT 647.100 451.050 648.900 452.850 ;
        RECT 652.950 447.600 654.150 452.850 ;
        RECT 655.950 449.850 658.050 451.950 ;
        RECT 668.100 451.050 669.900 452.850 ;
        RECT 655.950 448.050 657.750 449.850 ;
        RECT 673.950 447.600 675.150 452.850 ;
        RECT 676.950 449.850 679.050 451.950 ;
        RECT 686.100 451.050 687.900 452.850 ;
        RECT 676.950 448.050 678.750 449.850 ;
        RECT 691.950 447.600 693.150 452.850 ;
        RECT 694.950 449.850 697.050 451.950 ;
        RECT 706.950 451.050 709.050 453.150 ;
        RECT 694.950 448.050 696.750 449.850 ;
        RECT 619.500 435.750 621.300 441.600 ;
        RECT 622.500 435.750 624.300 441.600 ;
        RECT 625.500 435.750 627.300 441.600 ;
        RECT 632.550 435.750 634.350 441.600 ;
        RECT 635.550 435.750 637.350 441.600 ;
        RECT 648.300 435.750 650.100 447.600 ;
        RECT 652.500 435.750 654.300 447.600 ;
        RECT 655.800 435.750 657.600 441.600 ;
        RECT 669.300 435.750 671.100 447.600 ;
        RECT 673.500 435.750 675.300 447.600 ;
        RECT 676.800 435.750 678.600 441.600 ;
        RECT 687.300 435.750 689.100 447.600 ;
        RECT 691.500 435.750 693.300 447.600 ;
        RECT 707.250 442.800 708.300 451.050 ;
        RECT 709.950 449.850 712.050 451.950 ;
        RECT 715.950 449.850 718.050 451.950 ;
        RECT 709.950 448.050 711.750 449.850 ;
        RECT 712.950 446.850 715.050 448.950 ;
        RECT 716.100 448.050 717.900 449.850 ;
        RECT 725.550 447.450 726.900 454.050 ;
        RECT 728.400 450.150 729.300 458.400 ;
        RECT 733.950 455.850 736.050 457.950 ;
        RECT 730.950 452.850 733.050 454.950 ;
        RECT 734.100 454.050 735.900 455.850 ;
        RECT 743.100 453.150 744.900 454.950 ;
        RECT 731.100 451.050 732.900 452.850 ;
        RECT 742.950 451.050 745.050 453.150 ;
        RECT 746.250 451.950 747.450 459.300 ;
        RECT 749.100 453.150 750.900 454.950 ;
        RECT 758.100 453.150 759.900 454.950 ;
        RECT 728.250 450.000 730.050 450.150 ;
        RECT 728.250 448.800 735.450 450.000 ;
        RECT 745.950 449.850 748.050 451.950 ;
        RECT 748.950 451.050 751.050 453.150 ;
        RECT 757.950 451.050 760.050 453.150 ;
        RECT 761.250 451.950 762.450 459.300 ;
        RECT 770.400 456.150 771.600 464.400 ;
        RECT 764.100 453.150 765.900 454.950 ;
        RECT 769.950 454.050 772.050 456.150 ;
        RECT 772.950 455.850 775.050 457.950 ;
        RECT 781.050 456.150 782.550 464.400 ;
        RECT 773.100 454.050 774.900 455.850 ;
        RECT 778.950 454.050 782.550 456.150 ;
        RECT 760.950 449.850 763.050 451.950 ;
        RECT 763.950 451.050 766.050 453.150 ;
        RECT 728.250 448.350 730.050 448.800 ;
        RECT 734.250 447.600 735.450 448.800 ;
        RECT 713.100 445.050 714.900 446.850 ;
        RECT 725.550 446.100 727.950 447.450 ;
        RECT 707.250 441.900 714.300 442.800 ;
        RECT 707.250 441.600 708.450 441.900 ;
        RECT 694.800 435.750 696.600 441.600 ;
        RECT 706.650 435.750 708.450 441.600 ;
        RECT 712.650 441.600 714.300 441.900 ;
        RECT 709.650 435.750 711.450 441.000 ;
        RECT 712.650 435.750 714.450 441.600 ;
        RECT 715.650 435.750 717.450 441.600 ;
        RECT 726.150 435.750 727.950 446.100 ;
        RECT 729.150 435.750 730.950 447.450 ;
        RECT 733.650 435.750 735.450 447.600 ;
        RECT 746.250 441.600 747.450 449.850 ;
        RECT 761.250 441.600 762.450 449.850 ;
        RECT 770.400 441.600 771.600 454.050 ;
        RECT 781.050 441.600 782.550 454.050 ;
        RECT 784.650 461.400 786.450 467.250 ;
        RECT 790.050 461.400 791.850 467.250 ;
        RECT 795.600 462.600 797.400 467.250 ;
        RECT 800.250 463.500 802.050 467.250 ;
        RECT 803.250 463.500 805.050 467.250 ;
        RECT 806.250 463.500 808.050 467.250 ;
        RECT 793.200 461.400 797.400 462.600 ;
        RECT 799.950 461.400 802.050 463.500 ;
        RECT 802.950 461.400 805.050 463.500 ;
        RECT 805.950 461.400 808.050 463.500 ;
        RECT 810.000 463.500 811.800 467.250 ;
        RECT 813.000 464.400 814.800 467.250 ;
        RECT 816.000 463.500 817.800 467.250 ;
        RECT 820.500 464.400 822.300 467.250 ;
        RECT 823.500 464.400 825.300 467.250 ;
        RECT 826.500 464.400 828.300 467.250 ;
        RECT 829.500 464.400 831.300 467.250 ;
        RECT 810.000 461.700 812.850 463.500 ;
        RECT 810.750 461.400 812.850 461.700 ;
        RECT 814.950 461.700 817.800 463.500 ;
        RECT 818.700 462.750 820.500 463.200 ;
        RECT 823.950 463.050 825.300 464.400 ;
        RECT 826.950 463.050 828.300 464.400 ;
        RECT 829.950 463.050 831.300 464.400 ;
        RECT 814.950 461.400 817.050 461.700 ;
        RECT 818.700 461.400 822.750 462.750 ;
        RECT 784.650 446.550 785.850 461.400 ;
        RECT 793.200 457.800 794.700 461.400 ;
        RECT 799.350 458.700 806.100 460.500 ;
        RECT 807.000 458.700 813.900 460.500 ;
        RECT 821.850 460.050 822.750 461.400 ;
        RECT 823.950 460.950 826.050 463.050 ;
        RECT 826.950 460.950 829.050 463.050 ;
        RECT 829.950 460.950 832.050 463.050 ;
        RECT 821.850 459.900 826.950 460.050 ;
        RECT 821.850 459.150 829.500 459.900 ;
        RECT 825.150 458.700 829.500 459.150 ;
        RECT 807.000 457.800 808.050 458.700 ;
        RECT 825.150 458.250 826.950 458.700 ;
        RECT 786.900 456.000 794.700 457.800 ;
        RECT 798.150 456.750 808.050 457.800 ;
        RECT 798.150 454.950 799.200 456.750 ;
        RECT 808.950 456.450 816.600 457.800 ;
        RECT 808.950 455.700 809.850 456.450 ;
        RECT 790.950 453.900 799.200 454.950 ;
        RECT 800.250 454.650 809.850 455.700 ;
        RECT 790.950 449.850 793.050 453.900 ;
        RECT 800.250 453.000 801.150 454.650 ;
        RECT 810.750 453.750 814.650 455.550 ;
        RECT 815.550 454.950 816.600 456.450 ;
        RECT 817.950 457.650 820.050 457.950 ;
        RECT 817.950 455.850 821.850 457.650 ;
        RECT 828.450 455.250 829.500 458.700 ;
        RECT 831.000 457.800 832.050 460.950 ;
        RECT 833.700 461.400 835.500 467.250 ;
        RECT 839.100 461.400 840.900 467.250 ;
        RECT 844.500 461.400 846.300 467.250 ;
        RECT 833.700 460.500 835.200 461.400 ;
        RECT 833.700 459.300 842.100 460.500 ;
        RECT 840.300 458.700 842.100 459.300 ;
        RECT 845.100 457.800 846.300 461.400 ;
        RECT 831.000 456.900 846.300 457.800 ;
        RECT 815.550 454.050 827.550 454.950 ;
        RECT 794.100 451.200 801.150 453.000 ;
        RECT 802.500 451.950 804.300 453.750 ;
        RECT 810.750 453.450 812.850 453.750 ;
        RECT 814.950 452.550 817.050 452.850 ;
        RECT 823.800 452.550 825.600 453.150 ;
        RECT 814.950 451.950 825.600 452.550 ;
        RECT 802.500 451.350 825.600 451.950 ;
        RECT 826.500 452.550 827.550 454.050 ;
        RECT 828.450 453.450 830.250 455.250 ;
        RECT 832.050 454.950 843.900 456.000 ;
        RECT 832.050 452.550 833.250 454.950 ;
        RECT 842.100 453.150 843.900 454.950 ;
        RECT 826.500 451.650 833.250 452.550 ;
        RECT 835.950 451.650 838.050 451.950 ;
        RECT 802.500 450.750 817.050 451.350 ;
        RECT 834.150 450.450 838.050 451.650 ;
        RECT 841.950 451.050 844.050 453.150 ;
        RECT 824.100 449.850 838.050 450.450 ;
        RECT 798.000 449.550 837.750 449.850 ;
        RECT 786.750 448.650 788.550 449.250 ;
        RECT 798.000 448.650 826.050 449.550 ;
        RECT 786.750 447.450 799.050 448.650 ;
        RECT 826.950 448.050 829.050 448.350 ;
        RECT 836.700 448.050 838.500 448.650 ;
        RECT 799.950 446.550 802.050 447.750 ;
        RECT 784.650 445.650 802.050 446.550 ;
        RECT 805.950 446.400 826.050 447.750 ;
        RECT 805.950 445.650 808.050 446.400 ;
        RECT 787.500 441.600 788.700 445.650 ;
        RECT 789.600 443.700 791.400 444.300 ;
        RECT 796.350 444.150 798.150 444.300 ;
        RECT 789.600 442.500 795.300 443.700 ;
        RECT 796.350 442.950 805.050 444.150 ;
        RECT 796.350 442.500 798.150 442.950 ;
        RECT 742.650 435.750 744.450 441.600 ;
        RECT 745.650 435.750 747.450 441.600 ;
        RECT 748.650 435.750 750.450 441.600 ;
        RECT 757.650 435.750 759.450 441.600 ;
        RECT 760.650 435.750 762.450 441.600 ;
        RECT 763.650 435.750 765.450 441.600 ;
        RECT 769.650 435.750 771.450 441.600 ;
        RECT 772.650 435.750 774.450 441.600 ;
        RECT 777.750 435.750 779.550 441.600 ;
        RECT 780.750 435.750 782.550 441.600 ;
        RECT 784.500 435.750 786.300 441.600 ;
        RECT 787.500 435.750 789.300 441.600 ;
        RECT 790.500 435.750 792.300 441.600 ;
        RECT 793.500 435.750 795.300 442.500 ;
        RECT 802.950 442.050 805.050 442.950 ;
        RECT 796.500 435.750 798.300 441.600 ;
        RECT 799.800 439.800 801.900 441.900 ;
        RECT 800.400 438.600 801.900 439.800 ;
        RECT 800.250 435.750 802.050 438.600 ;
        RECT 803.250 435.750 805.050 442.050 ;
        RECT 806.550 438.600 807.900 445.650 ;
        RECT 824.100 445.350 826.050 446.400 ;
        RECT 826.950 446.850 838.500 448.050 ;
        RECT 826.950 446.250 829.050 446.850 ;
        RECT 840.000 445.350 841.800 446.100 ;
        RECT 809.100 442.800 813.000 444.600 ;
        RECT 810.000 442.500 813.000 442.800 ;
        RECT 814.950 444.150 817.050 444.600 ;
        RECT 824.100 444.300 841.800 445.350 ;
        RECT 814.950 442.500 817.350 444.150 ;
        RECT 806.250 435.750 808.050 438.600 ;
        RECT 810.000 435.750 811.800 442.500 ;
        RECT 816.000 441.600 817.350 442.500 ;
        RECT 823.950 441.600 826.050 442.050 ;
        RECT 813.000 435.750 814.800 441.600 ;
        RECT 816.000 435.750 817.800 441.600 ;
        RECT 819.750 435.750 821.550 441.600 ;
        RECT 823.500 439.950 826.050 441.600 ;
        RECT 826.950 439.950 829.050 442.050 ;
        RECT 829.950 439.950 832.050 442.050 ;
        RECT 823.500 438.600 824.700 439.950 ;
        RECT 826.950 438.600 827.850 439.950 ;
        RECT 829.950 438.600 831.150 439.950 ;
        RECT 822.750 435.750 824.700 438.600 ;
        RECT 825.750 435.750 827.850 438.600 ;
        RECT 828.750 435.750 831.150 438.600 ;
        RECT 832.500 435.750 834.300 439.050 ;
        RECT 835.500 435.750 837.300 444.300 ;
        RECT 845.100 443.400 846.300 456.900 ;
        RECT 842.250 442.500 846.300 443.400 ;
        RECT 842.250 441.600 843.300 442.500 ;
        RECT 838.500 435.750 840.300 441.600 ;
        RECT 841.500 435.750 843.300 441.600 ;
        RECT 844.500 435.750 846.300 441.600 ;
        RECT 7.650 425.400 9.450 431.250 ;
        RECT 10.650 425.400 12.450 431.250 ;
        RECT 8.400 412.950 9.600 425.400 ;
        RECT 21.300 419.400 23.100 431.250 ;
        RECT 25.500 419.400 27.300 431.250 ;
        RECT 28.800 425.400 30.600 431.250 ;
        RECT 40.650 425.400 42.450 431.250 ;
        RECT 43.650 425.400 45.450 431.250 ;
        RECT 46.650 425.400 48.450 431.250 ;
        RECT 53.400 425.400 55.200 431.250 ;
        RECT 20.100 414.150 21.900 415.950 ;
        RECT 25.950 414.150 27.150 419.400 ;
        RECT 28.950 417.150 30.750 418.950 ;
        RECT 44.250 417.150 45.450 425.400 ;
        RECT 56.700 419.400 58.500 431.250 ;
        RECT 60.900 419.400 62.700 431.250 ;
        RECT 72.300 419.400 74.100 431.250 ;
        RECT 76.500 419.400 78.300 431.250 ;
        RECT 79.800 425.400 81.600 431.250 ;
        RECT 88.650 425.400 90.450 431.250 ;
        RECT 91.650 425.400 93.450 431.250 ;
        RECT 94.650 425.400 96.450 431.250 ;
        RECT 53.250 417.150 55.050 418.950 ;
        RECT 28.950 415.050 31.050 417.150 ;
        RECT 7.950 410.850 10.050 412.950 ;
        RECT 11.100 411.150 12.900 412.950 ;
        RECT 19.950 412.050 22.050 414.150 ;
        RECT 8.400 402.600 9.600 410.850 ;
        RECT 10.950 409.050 13.050 411.150 ;
        RECT 22.950 410.850 25.050 412.950 ;
        RECT 25.950 412.050 28.050 414.150 ;
        RECT 40.950 413.850 43.050 415.950 ;
        RECT 43.950 415.050 46.050 417.150 ;
        RECT 41.100 412.050 42.900 413.850 ;
        RECT 23.100 409.050 24.900 410.850 ;
        RECT 26.850 408.750 28.050 412.050 ;
        RECT 27.000 407.700 30.750 408.750 ;
        RECT 44.250 407.700 45.450 415.050 ;
        RECT 46.950 413.850 49.050 415.950 ;
        RECT 52.950 415.050 55.050 417.150 ;
        RECT 56.850 414.150 58.050 419.400 ;
        RECT 62.100 414.150 63.900 415.950 ;
        RECT 71.100 414.150 72.900 415.950 ;
        RECT 76.950 414.150 78.150 419.400 ;
        RECT 79.950 417.150 81.750 418.950 ;
        RECT 92.250 417.150 93.450 425.400 ;
        RECT 94.950 420.450 97.050 421.050 ;
        RECT 94.950 419.550 99.450 420.450 ;
        RECT 94.950 418.950 97.050 419.550 ;
        RECT 79.950 415.050 82.050 417.150 ;
        RECT 47.100 412.050 48.900 413.850 ;
        RECT 55.950 412.050 58.050 414.150 ;
        RECT 55.950 408.750 57.150 412.050 ;
        RECT 58.950 410.850 61.050 412.950 ;
        RECT 61.950 412.050 64.050 414.150 ;
        RECT 70.950 412.050 73.050 414.150 ;
        RECT 73.950 410.850 76.050 412.950 ;
        RECT 76.950 412.050 79.050 414.150 ;
        RECT 88.950 413.850 91.050 415.950 ;
        RECT 91.950 415.050 94.050 417.150 ;
        RECT 89.100 412.050 90.900 413.850 ;
        RECT 59.100 409.050 60.900 410.850 ;
        RECT 74.100 409.050 75.900 410.850 ;
        RECT 77.850 408.750 79.050 412.050 ;
        RECT 20.550 404.700 28.350 406.050 ;
        RECT 7.650 399.750 9.450 402.600 ;
        RECT 10.650 399.750 12.450 402.600 ;
        RECT 20.550 399.750 22.350 404.700 ;
        RECT 23.550 399.750 25.350 403.800 ;
        RECT 26.550 399.750 28.350 404.700 ;
        RECT 29.550 405.600 30.750 407.700 ;
        RECT 41.850 406.800 45.450 407.700 ;
        RECT 53.250 407.700 57.000 408.750 ;
        RECT 78.000 407.700 81.750 408.750 ;
        RECT 92.250 407.700 93.450 415.050 ;
        RECT 94.950 413.850 97.050 415.950 ;
        RECT 95.100 412.050 96.900 413.850 ;
        RECT 98.550 409.050 99.450 419.550 ;
        RECT 102.300 419.400 104.100 431.250 ;
        RECT 106.500 419.400 108.300 431.250 ;
        RECT 109.800 425.400 111.600 431.250 ;
        RECT 122.400 425.400 124.200 431.250 ;
        RECT 125.700 419.400 127.500 431.250 ;
        RECT 129.900 419.400 131.700 431.250 ;
        RECT 141.450 419.400 143.250 431.250 ;
        RECT 145.650 419.400 147.450 431.250 ;
        RECT 152.550 419.400 154.350 431.250 ;
        RECT 155.550 419.400 157.350 431.250 ;
        RECT 164.550 425.400 166.350 431.250 ;
        RECT 167.550 425.400 169.350 431.250 ;
        RECT 170.550 426.000 172.350 431.250 ;
        RECT 167.700 425.100 169.350 425.400 ;
        RECT 173.550 425.400 175.350 431.250 ;
        RECT 180.750 425.400 182.550 431.250 ;
        RECT 183.750 425.400 185.550 431.250 ;
        RECT 187.500 425.400 189.300 431.250 ;
        RECT 190.500 425.400 192.300 431.250 ;
        RECT 193.500 425.400 195.300 431.250 ;
        RECT 173.550 425.100 174.750 425.400 ;
        RECT 167.700 424.200 174.750 425.100 ;
        RECT 167.100 420.150 168.900 421.950 ;
        RECT 101.100 414.150 102.900 415.950 ;
        RECT 106.950 414.150 108.150 419.400 ;
        RECT 109.950 417.150 111.750 418.950 ;
        RECT 122.250 417.150 124.050 418.950 ;
        RECT 109.950 415.050 112.050 417.150 ;
        RECT 121.950 415.050 124.050 417.150 ;
        RECT 125.850 414.150 127.050 419.400 ;
        RECT 141.450 418.350 144.000 419.400 ;
        RECT 131.100 414.150 132.900 415.950 ;
        RECT 140.100 414.150 141.900 415.950 ;
        RECT 100.950 412.050 103.050 414.150 ;
        RECT 103.950 410.850 106.050 412.950 ;
        RECT 106.950 412.050 109.050 414.150 ;
        RECT 104.100 409.050 105.900 410.850 ;
        RECT 29.550 399.750 31.350 405.600 ;
        RECT 41.850 399.750 43.650 406.800 ;
        RECT 53.250 405.600 54.450 407.700 ;
        RECT 46.350 399.750 48.150 405.600 ;
        RECT 52.650 399.750 54.450 405.600 ;
        RECT 55.650 404.700 63.450 406.050 ;
        RECT 55.650 399.750 57.450 404.700 ;
        RECT 58.650 399.750 60.450 403.800 ;
        RECT 61.650 399.750 63.450 404.700 ;
        RECT 71.550 404.700 79.350 406.050 ;
        RECT 71.550 399.750 73.350 404.700 ;
        RECT 74.550 399.750 76.350 403.800 ;
        RECT 77.550 399.750 79.350 404.700 ;
        RECT 80.550 405.600 81.750 407.700 ;
        RECT 89.850 406.800 93.450 407.700 ;
        RECT 97.950 406.950 100.050 409.050 ;
        RECT 107.850 408.750 109.050 412.050 ;
        RECT 124.950 412.050 127.050 414.150 ;
        RECT 124.950 408.750 126.150 412.050 ;
        RECT 127.950 410.850 130.050 412.950 ;
        RECT 130.950 412.050 133.050 414.150 ;
        RECT 139.950 412.050 142.050 414.150 ;
        RECT 142.950 411.150 144.000 418.350 ;
        RECT 146.100 414.150 147.900 415.950 ;
        RECT 155.400 414.150 156.600 419.400 ;
        RECT 164.100 417.150 165.900 418.950 ;
        RECT 166.950 418.050 169.050 420.150 ;
        RECT 170.250 417.150 172.050 418.950 ;
        RECT 163.950 415.050 166.050 417.150 ;
        RECT 169.950 415.050 172.050 417.150 ;
        RECT 173.700 415.950 174.750 424.200 ;
        RECT 145.950 412.050 148.050 414.150 ;
        RECT 128.100 409.050 129.900 410.850 ;
        RECT 142.950 409.050 145.050 411.150 ;
        RECT 151.950 410.850 154.050 412.950 ;
        RECT 154.950 412.050 157.050 414.150 ;
        RECT 172.950 413.850 175.050 415.950 ;
        RECT 152.100 409.050 153.900 410.850 ;
        RECT 108.000 407.700 111.750 408.750 ;
        RECT 80.550 399.750 82.350 405.600 ;
        RECT 89.850 399.750 91.650 406.800 ;
        RECT 94.350 399.750 96.150 405.600 ;
        RECT 101.550 404.700 109.350 406.050 ;
        RECT 101.550 399.750 103.350 404.700 ;
        RECT 104.550 399.750 106.350 403.800 ;
        RECT 107.550 399.750 109.350 404.700 ;
        RECT 110.550 405.600 111.750 407.700 ;
        RECT 122.250 407.700 126.000 408.750 ;
        RECT 122.250 405.600 123.450 407.700 ;
        RECT 110.550 399.750 112.350 405.600 ;
        RECT 121.650 399.750 123.450 405.600 ;
        RECT 124.650 404.700 132.450 406.050 ;
        RECT 124.650 399.750 126.450 404.700 ;
        RECT 127.650 399.750 129.450 403.800 ;
        RECT 130.650 399.750 132.450 404.700 ;
        RECT 142.950 402.600 144.000 409.050 ;
        RECT 155.400 405.600 156.600 412.050 ;
        RECT 173.400 409.650 174.600 413.850 ;
        RECT 184.050 412.950 185.550 425.400 ;
        RECT 190.500 421.350 191.700 425.400 ;
        RECT 196.500 424.500 198.300 431.250 ;
        RECT 199.500 425.400 201.300 431.250 ;
        RECT 203.250 428.400 205.050 431.250 ;
        RECT 203.400 427.200 204.900 428.400 ;
        RECT 202.800 425.100 204.900 427.200 ;
        RECT 206.250 424.950 208.050 431.250 ;
        RECT 209.250 428.400 211.050 431.250 ;
        RECT 192.600 423.300 198.300 424.500 ;
        RECT 199.350 424.050 201.150 424.500 ;
        RECT 205.950 424.050 208.050 424.950 ;
        RECT 192.600 422.700 194.400 423.300 ;
        RECT 199.350 422.850 208.050 424.050 ;
        RECT 199.350 422.700 201.150 422.850 ;
        RECT 209.550 421.350 210.900 428.400 ;
        RECT 213.000 424.500 214.800 431.250 ;
        RECT 216.000 425.400 217.800 431.250 ;
        RECT 219.000 425.400 220.800 431.250 ;
        RECT 222.750 425.400 224.550 431.250 ;
        RECT 225.750 428.400 227.700 431.250 ;
        RECT 228.750 428.400 230.850 431.250 ;
        RECT 231.750 428.400 234.150 431.250 ;
        RECT 226.500 427.050 227.700 428.400 ;
        RECT 229.950 427.050 230.850 428.400 ;
        RECT 232.950 427.050 234.150 428.400 ;
        RECT 235.500 427.950 237.300 431.250 ;
        RECT 226.500 425.400 229.050 427.050 ;
        RECT 219.000 424.500 220.350 425.400 ;
        RECT 226.950 424.950 229.050 425.400 ;
        RECT 229.950 424.950 232.050 427.050 ;
        RECT 232.950 424.950 235.050 427.050 ;
        RECT 213.000 424.200 216.000 424.500 ;
        RECT 212.100 422.400 216.000 424.200 ;
        RECT 217.950 422.850 220.350 424.500 ;
        RECT 217.950 422.400 220.050 422.850 ;
        RECT 238.500 422.700 240.300 431.250 ;
        RECT 241.500 425.400 243.300 431.250 ;
        RECT 244.500 425.400 246.300 431.250 ;
        RECT 247.500 425.400 249.300 431.250 ;
        RECT 245.250 424.500 246.300 425.400 ;
        RECT 245.250 423.600 249.300 424.500 ;
        RECT 227.100 421.650 244.800 422.700 ;
        RECT 181.950 410.850 185.550 412.950 ;
        RECT 139.650 399.750 141.450 402.600 ;
        RECT 142.650 399.750 144.450 402.600 ;
        RECT 145.650 399.750 147.450 402.600 ;
        RECT 152.550 399.750 154.350 405.600 ;
        RECT 155.550 399.750 157.350 405.600 ;
        RECT 164.700 399.750 166.500 408.600 ;
        RECT 170.100 408.000 174.600 409.650 ;
        RECT 170.100 399.750 171.900 408.000 ;
        RECT 184.050 402.600 185.550 410.850 ;
        RECT 180.750 399.750 182.550 402.600 ;
        RECT 183.750 399.750 185.550 402.600 ;
        RECT 187.650 420.450 205.050 421.350 ;
        RECT 187.650 405.600 188.850 420.450 ;
        RECT 189.750 418.350 202.050 419.550 ;
        RECT 202.950 419.250 205.050 420.450 ;
        RECT 208.950 420.600 211.050 421.350 ;
        RECT 227.100 420.600 229.050 421.650 ;
        RECT 243.000 420.900 244.800 421.650 ;
        RECT 208.950 419.250 229.050 420.600 ;
        RECT 229.950 420.150 232.050 420.750 ;
        RECT 229.950 418.950 241.500 420.150 ;
        RECT 229.950 418.650 232.050 418.950 ;
        RECT 239.700 418.350 241.500 418.950 ;
        RECT 189.750 417.750 191.550 418.350 ;
        RECT 201.000 417.450 229.050 418.350 ;
        RECT 201.000 417.150 240.750 417.450 ;
        RECT 193.950 413.100 196.050 417.150 ;
        RECT 227.100 416.550 241.050 417.150 ;
        RECT 197.100 414.000 204.150 415.800 ;
        RECT 193.950 412.050 202.200 413.100 ;
        RECT 189.900 409.200 197.700 411.000 ;
        RECT 201.150 410.250 202.200 412.050 ;
        RECT 203.250 412.350 204.150 414.000 ;
        RECT 205.500 415.650 220.050 416.250 ;
        RECT 205.500 415.050 228.600 415.650 ;
        RECT 237.150 415.350 241.050 416.550 ;
        RECT 205.500 413.250 207.300 415.050 ;
        RECT 217.950 414.450 228.600 415.050 ;
        RECT 217.950 414.150 220.050 414.450 ;
        RECT 226.800 413.850 228.600 414.450 ;
        RECT 229.500 414.450 236.250 415.350 ;
        RECT 238.950 415.050 241.050 415.350 ;
        RECT 213.750 413.250 215.850 413.550 ;
        RECT 203.250 411.300 212.850 412.350 ;
        RECT 213.750 411.450 217.650 413.250 ;
        RECT 229.500 412.950 230.550 414.450 ;
        RECT 218.550 412.050 230.550 412.950 ;
        RECT 211.950 410.550 212.850 411.300 ;
        RECT 218.550 410.550 219.600 412.050 ;
        RECT 231.450 411.750 233.250 413.550 ;
        RECT 235.050 412.050 236.250 414.450 ;
        RECT 244.950 413.850 247.050 415.950 ;
        RECT 245.100 412.050 246.900 413.850 ;
        RECT 201.150 409.200 211.050 410.250 ;
        RECT 211.950 409.200 219.600 410.550 ;
        RECT 220.950 409.350 224.850 411.150 ;
        RECT 196.200 405.600 197.700 409.200 ;
        RECT 210.000 408.300 211.050 409.200 ;
        RECT 220.950 409.050 223.050 409.350 ;
        RECT 228.150 408.300 229.950 408.750 ;
        RECT 231.450 408.300 232.500 411.750 ;
        RECT 235.050 411.000 246.900 412.050 ;
        RECT 248.100 410.100 249.300 423.600 ;
        RECT 255.300 419.400 257.100 431.250 ;
        RECT 259.500 419.400 261.300 431.250 ;
        RECT 262.800 425.400 264.600 431.250 ;
        RECT 275.400 425.400 277.200 431.250 ;
        RECT 278.700 419.400 280.500 431.250 ;
        RECT 282.900 419.400 284.700 431.250 ;
        RECT 287.550 425.400 289.350 431.250 ;
        RECT 290.550 425.400 292.350 431.250 ;
        RECT 301.650 425.400 303.450 431.250 ;
        RECT 304.650 426.000 306.450 431.250 ;
        RECT 254.100 414.150 255.900 415.950 ;
        RECT 259.950 414.150 261.150 419.400 ;
        RECT 262.950 417.150 264.750 418.950 ;
        RECT 275.250 417.150 277.050 418.950 ;
        RECT 262.950 415.050 265.050 417.150 ;
        RECT 274.950 415.050 277.050 417.150 ;
        RECT 278.850 414.150 280.050 419.400 ;
        RECT 284.100 414.150 285.900 415.950 ;
        RECT 253.950 412.050 256.050 414.150 ;
        RECT 256.950 410.850 259.050 412.950 ;
        RECT 259.950 412.050 262.050 414.150 ;
        RECT 202.350 406.500 209.100 408.300 ;
        RECT 210.000 406.500 216.900 408.300 ;
        RECT 228.150 407.850 232.500 408.300 ;
        RECT 224.850 407.100 232.500 407.850 ;
        RECT 234.000 409.200 249.300 410.100 ;
        RECT 224.850 406.950 229.950 407.100 ;
        RECT 224.850 405.600 225.750 406.950 ;
        RECT 234.000 406.050 235.050 409.200 ;
        RECT 243.300 407.700 245.100 408.300 ;
        RECT 187.650 399.750 189.450 405.600 ;
        RECT 193.050 399.750 194.850 405.600 ;
        RECT 196.200 404.400 200.400 405.600 ;
        RECT 198.600 399.750 200.400 404.400 ;
        RECT 202.950 403.500 205.050 405.600 ;
        RECT 205.950 403.500 208.050 405.600 ;
        RECT 208.950 403.500 211.050 405.600 ;
        RECT 213.750 405.300 215.850 405.600 ;
        RECT 203.250 399.750 205.050 403.500 ;
        RECT 206.250 399.750 208.050 403.500 ;
        RECT 209.250 399.750 211.050 403.500 ;
        RECT 213.000 403.500 215.850 405.300 ;
        RECT 217.950 405.300 220.050 405.600 ;
        RECT 217.950 403.500 220.800 405.300 ;
        RECT 221.700 404.250 225.750 405.600 ;
        RECT 221.700 403.800 223.500 404.250 ;
        RECT 226.950 403.950 229.050 406.050 ;
        RECT 229.950 403.950 232.050 406.050 ;
        RECT 232.950 403.950 235.050 406.050 ;
        RECT 236.700 406.500 245.100 407.700 ;
        RECT 236.700 405.600 238.200 406.500 ;
        RECT 248.100 405.600 249.300 409.200 ;
        RECT 257.100 409.050 258.900 410.850 ;
        RECT 260.850 408.750 262.050 412.050 ;
        RECT 277.950 412.050 280.050 414.150 ;
        RECT 277.950 408.750 279.150 412.050 ;
        RECT 280.950 410.850 283.050 412.950 ;
        RECT 283.950 412.050 286.050 414.150 ;
        RECT 290.400 412.950 291.600 425.400 ;
        RECT 302.250 425.100 303.450 425.400 ;
        RECT 307.650 425.400 309.450 431.250 ;
        RECT 310.650 425.400 312.450 431.250 ;
        RECT 320.400 425.400 322.200 431.250 ;
        RECT 307.650 425.100 309.300 425.400 ;
        RECT 302.250 424.200 309.300 425.100 ;
        RECT 302.250 415.950 303.300 424.200 ;
        RECT 308.100 420.150 309.900 421.950 ;
        RECT 304.950 417.150 306.750 418.950 ;
        RECT 307.950 418.050 310.050 420.150 ;
        RECT 323.700 419.400 325.500 431.250 ;
        RECT 327.900 419.400 329.700 431.250 ;
        RECT 335.550 425.400 337.350 431.250 ;
        RECT 338.550 425.400 340.350 431.250 ;
        RECT 341.550 425.400 343.350 431.250 ;
        RECT 347.550 425.400 349.350 431.250 ;
        RECT 350.550 425.400 352.350 431.250 ;
        RECT 353.550 426.000 355.350 431.250 ;
        RECT 311.100 417.150 312.900 418.950 ;
        RECT 320.250 417.150 322.050 418.950 ;
        RECT 301.950 413.850 304.050 415.950 ;
        RECT 304.950 415.050 307.050 417.150 ;
        RECT 310.950 415.050 313.050 417.150 ;
        RECT 319.950 415.050 322.050 417.150 ;
        RECT 323.850 414.150 325.050 419.400 ;
        RECT 338.550 417.150 339.750 425.400 ;
        RECT 350.700 425.100 352.350 425.400 ;
        RECT 356.550 425.400 358.350 431.250 ;
        RECT 368.550 425.400 370.350 431.250 ;
        RECT 371.550 425.400 373.350 431.250 ;
        RECT 374.550 426.000 376.350 431.250 ;
        RECT 356.550 425.100 357.750 425.400 ;
        RECT 350.700 424.200 357.750 425.100 ;
        RECT 371.700 425.100 373.350 425.400 ;
        RECT 377.550 425.400 379.350 431.250 ;
        RECT 377.550 425.100 378.750 425.400 ;
        RECT 371.700 424.200 378.750 425.100 ;
        RECT 350.100 420.150 351.900 421.950 ;
        RECT 347.100 417.150 348.900 418.950 ;
        RECT 349.950 418.050 352.050 420.150 ;
        RECT 353.250 417.150 355.050 418.950 ;
        RECT 329.100 414.150 330.900 415.950 ;
        RECT 287.100 411.150 288.900 412.950 ;
        RECT 281.100 409.050 282.900 410.850 ;
        RECT 286.950 409.050 289.050 411.150 ;
        RECT 289.950 410.850 292.050 412.950 ;
        RECT 261.000 407.700 264.750 408.750 ;
        RECT 213.000 399.750 214.800 403.500 ;
        RECT 216.000 399.750 217.800 402.600 ;
        RECT 219.000 399.750 220.800 403.500 ;
        RECT 226.950 402.600 228.300 403.950 ;
        RECT 229.950 402.600 231.300 403.950 ;
        RECT 232.950 402.600 234.300 403.950 ;
        RECT 223.500 399.750 225.300 402.600 ;
        RECT 226.500 399.750 228.300 402.600 ;
        RECT 229.500 399.750 231.300 402.600 ;
        RECT 232.500 399.750 234.300 402.600 ;
        RECT 236.700 399.750 238.500 405.600 ;
        RECT 242.100 399.750 243.900 405.600 ;
        RECT 247.500 399.750 249.300 405.600 ;
        RECT 254.550 404.700 262.350 406.050 ;
        RECT 254.550 399.750 256.350 404.700 ;
        RECT 257.550 399.750 259.350 403.800 ;
        RECT 260.550 399.750 262.350 404.700 ;
        RECT 263.550 405.600 264.750 407.700 ;
        RECT 275.250 407.700 279.000 408.750 ;
        RECT 275.250 405.600 276.450 407.700 ;
        RECT 263.550 399.750 265.350 405.600 ;
        RECT 274.650 399.750 276.450 405.600 ;
        RECT 277.650 404.700 285.450 406.050 ;
        RECT 277.650 399.750 279.450 404.700 ;
        RECT 280.650 399.750 282.450 403.800 ;
        RECT 283.650 399.750 285.450 404.700 ;
        RECT 290.400 402.600 291.600 410.850 ;
        RECT 302.400 409.650 303.600 413.850 ;
        RECT 322.950 412.050 325.050 414.150 ;
        RECT 302.400 408.000 306.900 409.650 ;
        RECT 322.950 408.750 324.150 412.050 ;
        RECT 325.950 410.850 328.050 412.950 ;
        RECT 328.950 412.050 331.050 414.150 ;
        RECT 334.950 413.850 337.050 415.950 ;
        RECT 337.950 415.050 340.050 417.150 ;
        RECT 335.100 412.050 336.900 413.850 ;
        RECT 326.100 409.050 327.900 410.850 ;
        RECT 287.550 399.750 289.350 402.600 ;
        RECT 290.550 399.750 292.350 402.600 ;
        RECT 305.100 399.750 306.900 408.000 ;
        RECT 310.500 399.750 312.300 408.600 ;
        RECT 320.250 407.700 324.000 408.750 ;
        RECT 338.550 407.700 339.750 415.050 ;
        RECT 340.950 413.850 343.050 415.950 ;
        RECT 346.950 415.050 349.050 417.150 ;
        RECT 352.950 415.050 355.050 417.150 ;
        RECT 356.700 415.950 357.750 424.200 ;
        RECT 371.100 420.150 372.900 421.950 ;
        RECT 368.100 417.150 369.900 418.950 ;
        RECT 370.950 418.050 373.050 420.150 ;
        RECT 374.250 417.150 376.050 418.950 ;
        RECT 355.950 413.850 358.050 415.950 ;
        RECT 367.950 415.050 370.050 417.150 ;
        RECT 373.950 415.050 376.050 417.150 ;
        RECT 377.700 415.950 378.750 424.200 ;
        RECT 384.300 419.400 386.100 431.250 ;
        RECT 388.500 419.400 390.300 431.250 ;
        RECT 391.800 425.400 393.600 431.250 ;
        RECT 400.650 425.400 402.450 431.250 ;
        RECT 403.650 425.400 405.450 431.250 ;
        RECT 406.650 425.400 408.450 431.250 ;
        RECT 412.650 425.400 414.450 431.250 ;
        RECT 415.650 425.400 417.450 431.250 ;
        RECT 425.550 425.400 427.350 431.250 ;
        RECT 428.550 425.400 430.350 431.250 ;
        RECT 431.550 426.000 433.350 431.250 ;
        RECT 376.950 413.850 379.050 415.950 ;
        RECT 383.100 414.150 384.900 415.950 ;
        RECT 388.950 414.150 390.150 419.400 ;
        RECT 391.950 417.150 393.750 418.950 ;
        RECT 404.250 417.150 405.450 425.400 ;
        RECT 391.950 415.050 394.050 417.150 ;
        RECT 341.100 412.050 342.900 413.850 ;
        RECT 356.400 409.650 357.600 413.850 ;
        RECT 377.400 409.650 378.600 413.850 ;
        RECT 382.950 412.050 385.050 414.150 ;
        RECT 385.950 410.850 388.050 412.950 ;
        RECT 388.950 412.050 391.050 414.150 ;
        RECT 400.950 413.850 403.050 415.950 ;
        RECT 403.950 415.050 406.050 417.150 ;
        RECT 401.100 412.050 402.900 413.850 ;
        RECT 320.250 405.600 321.450 407.700 ;
        RECT 338.550 406.800 342.150 407.700 ;
        RECT 319.650 399.750 321.450 405.600 ;
        RECT 322.650 404.700 330.450 406.050 ;
        RECT 322.650 399.750 324.450 404.700 ;
        RECT 325.650 399.750 327.450 403.800 ;
        RECT 328.650 399.750 330.450 404.700 ;
        RECT 335.850 399.750 337.650 405.600 ;
        RECT 340.350 399.750 342.150 406.800 ;
        RECT 347.700 399.750 349.500 408.600 ;
        RECT 353.100 408.000 357.600 409.650 ;
        RECT 353.100 399.750 354.900 408.000 ;
        RECT 368.700 399.750 370.500 408.600 ;
        RECT 374.100 408.000 378.600 409.650 ;
        RECT 386.100 409.050 387.900 410.850 ;
        RECT 389.850 408.750 391.050 412.050 ;
        RECT 374.100 399.750 375.900 408.000 ;
        RECT 390.000 407.700 393.750 408.750 ;
        RECT 404.250 407.700 405.450 415.050 ;
        RECT 406.950 413.850 409.050 415.950 ;
        RECT 407.100 412.050 408.900 413.850 ;
        RECT 413.400 412.950 414.600 425.400 ;
        RECT 428.700 425.100 430.350 425.400 ;
        RECT 434.550 425.400 436.350 431.250 ;
        RECT 446.550 425.400 448.350 431.250 ;
        RECT 449.550 425.400 451.350 431.250 ;
        RECT 452.550 426.000 454.350 431.250 ;
        RECT 434.550 425.100 435.750 425.400 ;
        RECT 428.700 424.200 435.750 425.100 ;
        RECT 449.700 425.100 451.350 425.400 ;
        RECT 455.550 425.400 457.350 431.250 ;
        RECT 455.550 425.100 456.750 425.400 ;
        RECT 449.700 424.200 456.750 425.100 ;
        RECT 428.100 420.150 429.900 421.950 ;
        RECT 425.100 417.150 426.900 418.950 ;
        RECT 427.950 418.050 430.050 420.150 ;
        RECT 431.250 417.150 433.050 418.950 ;
        RECT 424.950 415.050 427.050 417.150 ;
        RECT 430.950 415.050 433.050 417.150 ;
        RECT 434.700 415.950 435.750 424.200 ;
        RECT 449.100 420.150 450.900 421.950 ;
        RECT 446.100 417.150 447.900 418.950 ;
        RECT 448.950 418.050 451.050 420.150 ;
        RECT 452.250 417.150 454.050 418.950 ;
        RECT 433.950 413.850 436.050 415.950 ;
        RECT 445.950 415.050 448.050 417.150 ;
        RECT 451.950 415.050 454.050 417.150 ;
        RECT 455.700 415.950 456.750 424.200 ;
        RECT 465.300 419.400 467.100 431.250 ;
        RECT 469.500 419.400 471.300 431.250 ;
        RECT 472.800 425.400 474.600 431.250 ;
        RECT 486.300 419.400 488.100 431.250 ;
        RECT 490.500 419.400 492.300 431.250 ;
        RECT 493.800 425.400 495.600 431.250 ;
        RECT 500.550 419.400 502.350 431.250 ;
        RECT 505.050 419.550 506.850 431.250 ;
        RECT 508.050 420.900 509.850 431.250 ;
        RECT 508.050 419.550 510.450 420.900 ;
        RECT 454.950 413.850 457.050 415.950 ;
        RECT 464.100 414.150 465.900 415.950 ;
        RECT 469.950 414.150 471.150 419.400 ;
        RECT 472.950 417.150 474.750 418.950 ;
        RECT 472.950 415.050 475.050 417.150 ;
        RECT 485.100 414.150 486.900 415.950 ;
        RECT 490.950 414.150 492.150 419.400 ;
        RECT 493.950 417.150 495.750 418.950 ;
        RECT 500.550 418.200 501.750 419.400 ;
        RECT 505.950 418.200 507.750 418.650 ;
        RECT 493.950 415.050 496.050 417.150 ;
        RECT 500.550 417.000 507.750 418.200 ;
        RECT 505.950 416.850 507.750 417.000 ;
        RECT 503.100 414.150 504.900 415.950 ;
        RECT 412.950 410.850 415.050 412.950 ;
        RECT 416.100 411.150 417.900 412.950 ;
        RECT 383.550 404.700 391.350 406.050 ;
        RECT 383.550 399.750 385.350 404.700 ;
        RECT 386.550 399.750 388.350 403.800 ;
        RECT 389.550 399.750 391.350 404.700 ;
        RECT 392.550 405.600 393.750 407.700 ;
        RECT 401.850 406.800 405.450 407.700 ;
        RECT 392.550 399.750 394.350 405.600 ;
        RECT 401.850 399.750 403.650 406.800 ;
        RECT 406.350 399.750 408.150 405.600 ;
        RECT 413.400 402.600 414.600 410.850 ;
        RECT 415.950 409.050 418.050 411.150 ;
        RECT 434.400 409.650 435.600 413.850 ;
        RECT 455.400 409.650 456.600 413.850 ;
        RECT 463.950 412.050 466.050 414.150 ;
        RECT 466.950 410.850 469.050 412.950 ;
        RECT 469.950 412.050 472.050 414.150 ;
        RECT 484.950 412.050 487.050 414.150 ;
        RECT 412.650 399.750 414.450 402.600 ;
        RECT 415.650 399.750 417.450 402.600 ;
        RECT 425.700 399.750 427.500 408.600 ;
        RECT 431.100 408.000 435.600 409.650 ;
        RECT 431.100 399.750 432.900 408.000 ;
        RECT 446.700 399.750 448.500 408.600 ;
        RECT 452.100 408.000 456.600 409.650 ;
        RECT 467.100 409.050 468.900 410.850 ;
        RECT 470.850 408.750 472.050 412.050 ;
        RECT 487.950 410.850 490.050 412.950 ;
        RECT 490.950 412.050 493.050 414.150 ;
        RECT 488.100 409.050 489.900 410.850 ;
        RECT 491.850 408.750 493.050 412.050 ;
        RECT 500.100 411.150 501.900 412.950 ;
        RECT 502.950 412.050 505.050 414.150 ;
        RECT 499.950 409.050 502.050 411.150 ;
        RECT 452.100 399.750 453.900 408.000 ;
        RECT 471.000 407.700 474.750 408.750 ;
        RECT 492.000 407.700 495.750 408.750 ;
        RECT 506.700 408.600 507.600 416.850 ;
        RECT 509.100 412.950 510.450 419.550 ;
        RECT 521.550 419.400 523.350 431.250 ;
        RECT 525.750 419.400 527.550 431.250 ;
        RECT 533.550 420.300 535.350 431.250 ;
        RECT 536.550 421.200 538.350 431.250 ;
        RECT 539.550 420.300 541.350 431.250 ;
        RECT 533.550 419.400 541.350 420.300 ;
        RECT 542.550 419.400 544.350 431.250 ;
        RECT 548.550 425.400 550.350 431.250 ;
        RECT 551.550 425.400 553.350 431.250 ;
        RECT 557.550 425.400 559.350 431.250 ;
        RECT 560.550 425.400 562.350 431.250 ;
        RECT 572.550 425.400 574.350 431.250 ;
        RECT 525.000 418.350 527.550 419.400 ;
        RECT 521.100 414.150 522.900 415.950 ;
        RECT 508.950 410.850 511.050 412.950 ;
        RECT 520.950 412.050 523.050 414.150 ;
        RECT 525.000 411.150 526.050 418.350 ;
        RECT 527.100 414.150 528.900 415.950 ;
        RECT 542.700 414.150 543.900 419.400 ;
        RECT 526.950 412.050 529.050 414.150 ;
        RECT 505.950 407.700 507.750 408.600 ;
        RECT 464.550 404.700 472.350 406.050 ;
        RECT 464.550 399.750 466.350 404.700 ;
        RECT 467.550 399.750 469.350 403.800 ;
        RECT 470.550 399.750 472.350 404.700 ;
        RECT 473.550 405.600 474.750 407.700 ;
        RECT 473.550 399.750 475.350 405.600 ;
        RECT 485.550 404.700 493.350 406.050 ;
        RECT 485.550 399.750 487.350 404.700 ;
        RECT 488.550 399.750 490.350 403.800 ;
        RECT 491.550 399.750 493.350 404.700 ;
        RECT 494.550 405.600 495.750 407.700 ;
        RECT 504.450 406.800 507.750 407.700 ;
        RECT 494.550 399.750 496.350 405.600 ;
        RECT 504.450 402.600 505.350 406.800 ;
        RECT 510.000 405.600 511.050 410.850 ;
        RECT 523.950 409.050 526.050 411.150 ;
        RECT 532.950 410.850 535.050 412.950 ;
        RECT 536.100 411.150 537.900 412.950 ;
        RECT 533.100 409.050 534.900 410.850 ;
        RECT 535.950 409.050 538.050 411.150 ;
        RECT 538.950 410.850 541.050 412.950 ;
        RECT 541.950 412.050 544.050 414.150 ;
        RECT 551.400 412.950 552.600 425.400 ;
        RECT 560.400 412.950 561.600 425.400 ;
        RECT 572.550 418.500 573.750 425.400 ;
        RECT 575.850 419.400 577.650 431.250 ;
        RECT 578.850 419.400 580.650 431.250 ;
        RECT 586.650 419.400 588.450 431.250 ;
        RECT 572.550 417.600 578.250 418.500 ;
        RECT 576.000 416.700 578.250 417.600 ;
        RECT 572.100 414.150 573.900 415.950 ;
        RECT 539.100 409.050 540.900 410.850 ;
        RECT 500.550 399.750 502.350 402.600 ;
        RECT 503.550 399.750 505.350 402.600 ;
        RECT 506.550 399.750 508.350 402.600 ;
        RECT 509.550 399.750 511.350 405.600 ;
        RECT 525.000 402.600 526.050 409.050 ;
        RECT 542.700 405.600 543.900 412.050 ;
        RECT 548.100 411.150 549.900 412.950 ;
        RECT 547.950 409.050 550.050 411.150 ;
        RECT 550.950 410.850 553.050 412.950 ;
        RECT 557.100 411.150 558.900 412.950 ;
        RECT 521.550 399.750 523.350 402.600 ;
        RECT 524.550 399.750 526.350 402.600 ;
        RECT 527.550 399.750 529.350 402.600 ;
        RECT 534.000 399.750 535.800 405.600 ;
        RECT 538.200 403.950 543.900 405.600 ;
        RECT 538.200 399.750 540.000 403.950 ;
        RECT 551.400 402.600 552.600 410.850 ;
        RECT 556.950 409.050 559.050 411.150 ;
        RECT 559.950 410.850 562.050 412.950 ;
        RECT 571.950 412.050 574.050 414.150 ;
        RECT 560.400 402.600 561.600 410.850 ;
        RECT 576.000 408.300 577.050 416.700 ;
        RECT 579.150 414.150 580.350 419.400 ;
        RECT 589.650 418.500 591.450 431.250 ;
        RECT 592.650 419.400 594.450 431.250 ;
        RECT 595.650 418.500 597.450 431.250 ;
        RECT 598.650 419.400 600.450 431.250 ;
        RECT 601.650 418.500 603.450 431.250 ;
        RECT 604.650 419.400 606.450 431.250 ;
        RECT 607.650 418.500 609.450 431.250 ;
        RECT 610.650 419.400 612.450 431.250 ;
        RECT 620.400 425.400 622.200 431.250 ;
        RECT 616.950 421.950 619.050 424.050 ;
        RECT 577.950 412.050 580.350 414.150 ;
        RECT 588.750 417.300 591.450 418.500 ;
        RECT 593.700 417.300 597.450 418.500 ;
        RECT 599.700 417.300 603.450 418.500 ;
        RECT 605.550 417.300 609.450 418.500 ;
        RECT 588.750 412.950 589.800 417.300 ;
        RECT 576.000 407.400 578.250 408.300 ;
        RECT 573.150 406.500 578.250 407.400 ;
        RECT 573.150 402.600 574.350 406.500 ;
        RECT 579.150 405.600 580.350 412.050 ;
        RECT 586.950 410.850 589.800 412.950 ;
        RECT 588.750 407.700 589.800 410.850 ;
        RECT 593.700 410.400 594.900 417.300 ;
        RECT 599.700 410.400 600.900 417.300 ;
        RECT 605.550 410.400 606.750 417.300 ;
        RECT 607.950 410.850 610.050 412.950 ;
        RECT 617.550 411.450 618.450 421.950 ;
        RECT 623.700 419.400 625.500 431.250 ;
        RECT 627.900 419.400 629.700 431.250 ;
        RECT 633.750 425.400 635.550 431.250 ;
        RECT 636.750 425.400 638.550 431.250 ;
        RECT 640.500 425.400 642.300 431.250 ;
        RECT 643.500 425.400 645.300 431.250 ;
        RECT 646.500 425.400 648.300 431.250 ;
        RECT 620.250 417.150 622.050 418.950 ;
        RECT 619.950 415.050 622.050 417.150 ;
        RECT 623.850 414.150 625.050 419.400 ;
        RECT 629.100 414.150 630.900 415.950 ;
        RECT 622.950 412.050 625.050 414.150 ;
        RECT 619.950 411.450 622.050 412.050 ;
        RECT 590.700 408.600 594.900 410.400 ;
        RECT 596.700 408.600 600.900 410.400 ;
        RECT 602.700 408.600 606.750 410.400 ;
        RECT 608.100 409.050 609.900 410.850 ;
        RECT 617.550 410.550 622.050 411.450 ;
        RECT 619.950 409.950 622.050 410.550 ;
        RECT 622.950 408.750 624.150 412.050 ;
        RECT 625.950 410.850 628.050 412.950 ;
        RECT 628.950 412.050 631.050 414.150 ;
        RECT 637.050 412.950 638.550 425.400 ;
        RECT 643.500 421.350 644.700 425.400 ;
        RECT 649.500 424.500 651.300 431.250 ;
        RECT 652.500 425.400 654.300 431.250 ;
        RECT 656.250 428.400 658.050 431.250 ;
        RECT 656.400 427.200 657.900 428.400 ;
        RECT 655.800 425.100 657.900 427.200 ;
        RECT 659.250 424.950 661.050 431.250 ;
        RECT 662.250 428.400 664.050 431.250 ;
        RECT 645.600 423.300 651.300 424.500 ;
        RECT 652.350 424.050 654.150 424.500 ;
        RECT 658.950 424.050 661.050 424.950 ;
        RECT 645.600 422.700 647.400 423.300 ;
        RECT 652.350 422.850 661.050 424.050 ;
        RECT 652.350 422.700 654.150 422.850 ;
        RECT 662.550 421.350 663.900 428.400 ;
        RECT 666.000 424.500 667.800 431.250 ;
        RECT 669.000 425.400 670.800 431.250 ;
        RECT 672.000 425.400 673.800 431.250 ;
        RECT 675.750 425.400 677.550 431.250 ;
        RECT 678.750 428.400 680.700 431.250 ;
        RECT 681.750 428.400 683.850 431.250 ;
        RECT 684.750 428.400 687.150 431.250 ;
        RECT 679.500 427.050 680.700 428.400 ;
        RECT 682.950 427.050 683.850 428.400 ;
        RECT 685.950 427.050 687.150 428.400 ;
        RECT 688.500 427.950 690.300 431.250 ;
        RECT 679.500 425.400 682.050 427.050 ;
        RECT 672.000 424.500 673.350 425.400 ;
        RECT 679.950 424.950 682.050 425.400 ;
        RECT 682.950 424.950 685.050 427.050 ;
        RECT 685.950 424.950 688.050 427.050 ;
        RECT 666.000 424.200 669.000 424.500 ;
        RECT 665.100 422.400 669.000 424.200 ;
        RECT 670.950 422.850 673.350 424.500 ;
        RECT 670.950 422.400 673.050 422.850 ;
        RECT 691.500 422.700 693.300 431.250 ;
        RECT 694.500 425.400 696.300 431.250 ;
        RECT 697.500 425.400 699.300 431.250 ;
        RECT 700.500 425.400 702.300 431.250 ;
        RECT 707.550 425.400 709.350 431.250 ;
        RECT 710.550 425.400 712.350 431.250 ;
        RECT 713.550 425.400 715.350 431.250 ;
        RECT 722.550 425.400 724.350 431.250 ;
        RECT 725.550 425.400 727.350 431.250 ;
        RECT 728.550 425.400 730.350 431.250 ;
        RECT 739.650 425.400 741.450 431.250 ;
        RECT 742.650 425.400 744.450 431.250 ;
        RECT 745.650 425.400 747.450 431.250 ;
        RECT 698.250 424.500 699.300 425.400 ;
        RECT 698.250 423.600 702.300 424.500 ;
        RECT 680.100 421.650 697.800 422.700 ;
        RECT 634.950 410.850 638.550 412.950 ;
        RECT 626.100 409.050 627.900 410.850 ;
        RECT 593.700 407.700 594.900 408.600 ;
        RECT 599.700 407.700 600.900 408.600 ;
        RECT 605.550 407.700 606.750 408.600 ;
        RECT 620.250 407.700 624.000 408.750 ;
        RECT 588.750 406.650 591.600 407.700 ;
        RECT 588.900 406.500 591.600 406.650 ;
        RECT 593.700 406.500 597.600 407.700 ;
        RECT 599.700 406.500 603.450 407.700 ;
        RECT 605.550 406.500 609.600 407.700 ;
        RECT 589.800 405.600 591.600 406.500 ;
        RECT 595.800 405.600 597.600 406.500 ;
        RECT 541.500 399.750 543.300 402.600 ;
        RECT 548.550 399.750 550.350 402.600 ;
        RECT 551.550 399.750 553.350 402.600 ;
        RECT 557.550 399.750 559.350 402.600 ;
        RECT 560.550 399.750 562.350 402.600 ;
        RECT 572.550 399.750 574.350 402.600 ;
        RECT 575.850 399.750 577.650 405.600 ;
        RECT 578.850 399.750 580.650 405.600 ;
        RECT 586.650 399.750 588.450 405.600 ;
        RECT 589.650 399.750 591.450 405.600 ;
        RECT 592.650 399.750 594.450 405.600 ;
        RECT 595.650 399.750 597.450 405.600 ;
        RECT 598.650 399.750 600.450 405.600 ;
        RECT 601.650 399.750 603.450 406.500 ;
        RECT 607.800 405.600 609.600 406.500 ;
        RECT 620.250 405.600 621.450 407.700 ;
        RECT 604.650 399.750 606.450 405.600 ;
        RECT 607.650 399.750 609.450 405.600 ;
        RECT 610.650 399.750 612.450 405.600 ;
        RECT 619.650 399.750 621.450 405.600 ;
        RECT 622.650 404.700 630.450 406.050 ;
        RECT 622.650 399.750 624.450 404.700 ;
        RECT 625.650 399.750 627.450 403.800 ;
        RECT 628.650 399.750 630.450 404.700 ;
        RECT 637.050 402.600 638.550 410.850 ;
        RECT 633.750 399.750 635.550 402.600 ;
        RECT 636.750 399.750 638.550 402.600 ;
        RECT 640.650 420.450 658.050 421.350 ;
        RECT 640.650 405.600 641.850 420.450 ;
        RECT 642.750 418.350 655.050 419.550 ;
        RECT 655.950 419.250 658.050 420.450 ;
        RECT 661.950 420.600 664.050 421.350 ;
        RECT 680.100 420.600 682.050 421.650 ;
        RECT 696.000 420.900 697.800 421.650 ;
        RECT 661.950 419.250 682.050 420.600 ;
        RECT 682.950 420.150 685.050 420.750 ;
        RECT 682.950 418.950 694.500 420.150 ;
        RECT 682.950 418.650 685.050 418.950 ;
        RECT 692.700 418.350 694.500 418.950 ;
        RECT 642.750 417.750 644.550 418.350 ;
        RECT 654.000 417.450 682.050 418.350 ;
        RECT 654.000 417.150 693.750 417.450 ;
        RECT 646.950 413.100 649.050 417.150 ;
        RECT 680.100 416.550 694.050 417.150 ;
        RECT 650.100 414.000 657.150 415.800 ;
        RECT 646.950 412.050 655.200 413.100 ;
        RECT 642.900 409.200 650.700 411.000 ;
        RECT 654.150 410.250 655.200 412.050 ;
        RECT 656.250 412.350 657.150 414.000 ;
        RECT 658.500 415.650 673.050 416.250 ;
        RECT 658.500 415.050 681.600 415.650 ;
        RECT 690.150 415.350 694.050 416.550 ;
        RECT 658.500 413.250 660.300 415.050 ;
        RECT 670.950 414.450 681.600 415.050 ;
        RECT 670.950 414.150 673.050 414.450 ;
        RECT 679.800 413.850 681.600 414.450 ;
        RECT 682.500 414.450 689.250 415.350 ;
        RECT 691.950 415.050 694.050 415.350 ;
        RECT 666.750 413.250 668.850 413.550 ;
        RECT 656.250 411.300 665.850 412.350 ;
        RECT 666.750 411.450 670.650 413.250 ;
        RECT 682.500 412.950 683.550 414.450 ;
        RECT 671.550 412.050 683.550 412.950 ;
        RECT 664.950 410.550 665.850 411.300 ;
        RECT 671.550 410.550 672.600 412.050 ;
        RECT 684.450 411.750 686.250 413.550 ;
        RECT 688.050 412.050 689.250 414.450 ;
        RECT 697.950 413.850 700.050 415.950 ;
        RECT 698.100 412.050 699.900 413.850 ;
        RECT 654.150 409.200 664.050 410.250 ;
        RECT 664.950 409.200 672.600 410.550 ;
        RECT 673.950 409.350 677.850 411.150 ;
        RECT 649.200 405.600 650.700 409.200 ;
        RECT 663.000 408.300 664.050 409.200 ;
        RECT 673.950 409.050 676.050 409.350 ;
        RECT 681.150 408.300 682.950 408.750 ;
        RECT 684.450 408.300 685.500 411.750 ;
        RECT 688.050 411.000 699.900 412.050 ;
        RECT 701.100 410.100 702.300 423.600 ;
        RECT 710.550 417.150 711.750 425.400 ;
        RECT 721.950 420.450 724.050 421.050 ;
        RECT 719.550 419.550 724.050 420.450 ;
        RECT 706.950 413.850 709.050 415.950 ;
        RECT 709.950 415.050 712.050 417.150 ;
        RECT 707.100 412.050 708.900 413.850 ;
        RECT 655.350 406.500 662.100 408.300 ;
        RECT 663.000 406.500 669.900 408.300 ;
        RECT 681.150 407.850 685.500 408.300 ;
        RECT 677.850 407.100 685.500 407.850 ;
        RECT 687.000 409.200 702.300 410.100 ;
        RECT 677.850 406.950 682.950 407.100 ;
        RECT 677.850 405.600 678.750 406.950 ;
        RECT 687.000 406.050 688.050 409.200 ;
        RECT 696.300 407.700 698.100 408.300 ;
        RECT 640.650 399.750 642.450 405.600 ;
        RECT 646.050 399.750 647.850 405.600 ;
        RECT 649.200 404.400 653.400 405.600 ;
        RECT 651.600 399.750 653.400 404.400 ;
        RECT 655.950 403.500 658.050 405.600 ;
        RECT 658.950 403.500 661.050 405.600 ;
        RECT 661.950 403.500 664.050 405.600 ;
        RECT 666.750 405.300 668.850 405.600 ;
        RECT 656.250 399.750 658.050 403.500 ;
        RECT 659.250 399.750 661.050 403.500 ;
        RECT 662.250 399.750 664.050 403.500 ;
        RECT 666.000 403.500 668.850 405.300 ;
        RECT 670.950 405.300 673.050 405.600 ;
        RECT 670.950 403.500 673.800 405.300 ;
        RECT 674.700 404.250 678.750 405.600 ;
        RECT 674.700 403.800 676.500 404.250 ;
        RECT 679.950 403.950 682.050 406.050 ;
        RECT 682.950 403.950 685.050 406.050 ;
        RECT 685.950 403.950 688.050 406.050 ;
        RECT 689.700 406.500 698.100 407.700 ;
        RECT 689.700 405.600 691.200 406.500 ;
        RECT 701.100 405.600 702.300 409.200 ;
        RECT 710.550 407.700 711.750 415.050 ;
        RECT 712.950 413.850 715.050 415.950 ;
        RECT 713.100 412.050 714.900 413.850 ;
        RECT 719.550 408.450 720.450 419.550 ;
        RECT 721.950 418.950 724.050 419.550 ;
        RECT 725.550 417.150 726.750 425.400 ;
        RECT 743.250 417.150 744.450 425.400 ;
        RECT 753.300 419.400 755.100 431.250 ;
        RECT 757.500 419.400 759.300 431.250 ;
        RECT 760.800 425.400 762.600 431.250 ;
        RECT 772.650 425.400 774.450 431.250 ;
        RECT 775.650 425.400 777.450 431.250 ;
        RECT 780.750 425.400 782.550 431.250 ;
        RECT 783.750 425.400 785.550 431.250 ;
        RECT 787.500 425.400 789.300 431.250 ;
        RECT 790.500 425.400 792.300 431.250 ;
        RECT 793.500 425.400 795.300 431.250 ;
        RECT 721.950 413.850 724.050 415.950 ;
        RECT 724.950 415.050 727.050 417.150 ;
        RECT 722.100 412.050 723.900 413.850 ;
        RECT 721.950 408.450 724.050 409.050 ;
        RECT 710.550 406.800 714.150 407.700 ;
        RECT 719.550 407.550 724.050 408.450 ;
        RECT 721.950 406.950 724.050 407.550 ;
        RECT 725.550 407.700 726.750 415.050 ;
        RECT 727.950 413.850 730.050 415.950 ;
        RECT 739.950 413.850 742.050 415.950 ;
        RECT 742.950 415.050 745.050 417.150 ;
        RECT 728.100 412.050 729.900 413.850 ;
        RECT 740.100 412.050 741.900 413.850 ;
        RECT 743.250 407.700 744.450 415.050 ;
        RECT 745.950 413.850 748.050 415.950 ;
        RECT 752.100 414.150 753.900 415.950 ;
        RECT 757.950 414.150 759.150 419.400 ;
        RECT 760.950 417.150 762.750 418.950 ;
        RECT 760.950 415.050 763.050 417.150 ;
        RECT 746.100 412.050 747.900 413.850 ;
        RECT 751.950 412.050 754.050 414.150 ;
        RECT 754.950 410.850 757.050 412.950 ;
        RECT 757.950 412.050 760.050 414.150 ;
        RECT 773.400 412.950 774.600 425.400 ;
        RECT 784.050 412.950 785.550 425.400 ;
        RECT 790.500 421.350 791.700 425.400 ;
        RECT 796.500 424.500 798.300 431.250 ;
        RECT 799.500 425.400 801.300 431.250 ;
        RECT 803.250 428.400 805.050 431.250 ;
        RECT 803.400 427.200 804.900 428.400 ;
        RECT 802.800 425.100 804.900 427.200 ;
        RECT 806.250 424.950 808.050 431.250 ;
        RECT 809.250 428.400 811.050 431.250 ;
        RECT 792.600 423.300 798.300 424.500 ;
        RECT 799.350 424.050 801.150 424.500 ;
        RECT 805.950 424.050 808.050 424.950 ;
        RECT 792.600 422.700 794.400 423.300 ;
        RECT 799.350 422.850 808.050 424.050 ;
        RECT 799.350 422.700 801.150 422.850 ;
        RECT 809.550 421.350 810.900 428.400 ;
        RECT 813.000 424.500 814.800 431.250 ;
        RECT 816.000 425.400 817.800 431.250 ;
        RECT 819.000 425.400 820.800 431.250 ;
        RECT 822.750 425.400 824.550 431.250 ;
        RECT 825.750 428.400 827.700 431.250 ;
        RECT 828.750 428.400 830.850 431.250 ;
        RECT 831.750 428.400 834.150 431.250 ;
        RECT 826.500 427.050 827.700 428.400 ;
        RECT 829.950 427.050 830.850 428.400 ;
        RECT 832.950 427.050 834.150 428.400 ;
        RECT 835.500 427.950 837.300 431.250 ;
        RECT 826.500 425.400 829.050 427.050 ;
        RECT 819.000 424.500 820.350 425.400 ;
        RECT 826.950 424.950 829.050 425.400 ;
        RECT 829.950 424.950 832.050 427.050 ;
        RECT 832.950 424.950 835.050 427.050 ;
        RECT 813.000 424.200 816.000 424.500 ;
        RECT 812.100 422.400 816.000 424.200 ;
        RECT 817.950 422.850 820.350 424.500 ;
        RECT 817.950 422.400 820.050 422.850 ;
        RECT 838.500 422.700 840.300 431.250 ;
        RECT 841.500 425.400 843.300 431.250 ;
        RECT 844.500 425.400 846.300 431.250 ;
        RECT 847.500 425.400 849.300 431.250 ;
        RECT 845.250 424.500 846.300 425.400 ;
        RECT 845.250 423.600 849.300 424.500 ;
        RECT 827.100 421.650 844.800 422.700 ;
        RECT 755.100 409.050 756.900 410.850 ;
        RECT 758.850 408.750 760.050 412.050 ;
        RECT 772.950 410.850 775.050 412.950 ;
        RECT 776.100 411.150 777.900 412.950 ;
        RECT 759.000 407.700 762.750 408.750 ;
        RECT 725.550 406.800 729.150 407.700 ;
        RECT 666.000 399.750 667.800 403.500 ;
        RECT 669.000 399.750 670.800 402.600 ;
        RECT 672.000 399.750 673.800 403.500 ;
        RECT 679.950 402.600 681.300 403.950 ;
        RECT 682.950 402.600 684.300 403.950 ;
        RECT 685.950 402.600 687.300 403.950 ;
        RECT 676.500 399.750 678.300 402.600 ;
        RECT 679.500 399.750 681.300 402.600 ;
        RECT 682.500 399.750 684.300 402.600 ;
        RECT 685.500 399.750 687.300 402.600 ;
        RECT 689.700 399.750 691.500 405.600 ;
        RECT 695.100 399.750 696.900 405.600 ;
        RECT 700.500 399.750 702.300 405.600 ;
        RECT 707.850 399.750 709.650 405.600 ;
        RECT 712.350 399.750 714.150 406.800 ;
        RECT 722.850 399.750 724.650 405.600 ;
        RECT 727.350 399.750 729.150 406.800 ;
        RECT 740.850 406.800 744.450 407.700 ;
        RECT 740.850 399.750 742.650 406.800 ;
        RECT 745.350 399.750 747.150 405.600 ;
        RECT 752.550 404.700 760.350 406.050 ;
        RECT 752.550 399.750 754.350 404.700 ;
        RECT 755.550 399.750 757.350 403.800 ;
        RECT 758.550 399.750 760.350 404.700 ;
        RECT 761.550 405.600 762.750 407.700 ;
        RECT 761.550 399.750 763.350 405.600 ;
        RECT 773.400 402.600 774.600 410.850 ;
        RECT 775.950 409.050 778.050 411.150 ;
        RECT 781.950 410.850 785.550 412.950 ;
        RECT 784.050 402.600 785.550 410.850 ;
        RECT 772.650 399.750 774.450 402.600 ;
        RECT 775.650 399.750 777.450 402.600 ;
        RECT 780.750 399.750 782.550 402.600 ;
        RECT 783.750 399.750 785.550 402.600 ;
        RECT 787.650 420.450 805.050 421.350 ;
        RECT 787.650 405.600 788.850 420.450 ;
        RECT 789.750 418.350 802.050 419.550 ;
        RECT 802.950 419.250 805.050 420.450 ;
        RECT 808.950 420.600 811.050 421.350 ;
        RECT 827.100 420.600 829.050 421.650 ;
        RECT 843.000 420.900 844.800 421.650 ;
        RECT 808.950 419.250 829.050 420.600 ;
        RECT 829.950 420.150 832.050 420.750 ;
        RECT 829.950 418.950 841.500 420.150 ;
        RECT 829.950 418.650 832.050 418.950 ;
        RECT 839.700 418.350 841.500 418.950 ;
        RECT 789.750 417.750 791.550 418.350 ;
        RECT 801.000 417.450 829.050 418.350 ;
        RECT 801.000 417.150 840.750 417.450 ;
        RECT 793.950 413.100 796.050 417.150 ;
        RECT 827.100 416.550 841.050 417.150 ;
        RECT 797.100 414.000 804.150 415.800 ;
        RECT 793.950 412.050 802.200 413.100 ;
        RECT 789.900 409.200 797.700 411.000 ;
        RECT 801.150 410.250 802.200 412.050 ;
        RECT 803.250 412.350 804.150 414.000 ;
        RECT 805.500 415.650 820.050 416.250 ;
        RECT 805.500 415.050 828.600 415.650 ;
        RECT 837.150 415.350 841.050 416.550 ;
        RECT 805.500 413.250 807.300 415.050 ;
        RECT 817.950 414.450 828.600 415.050 ;
        RECT 817.950 414.150 820.050 414.450 ;
        RECT 826.800 413.850 828.600 414.450 ;
        RECT 829.500 414.450 836.250 415.350 ;
        RECT 838.950 415.050 841.050 415.350 ;
        RECT 813.750 413.250 815.850 413.550 ;
        RECT 803.250 411.300 812.850 412.350 ;
        RECT 813.750 411.450 817.650 413.250 ;
        RECT 829.500 412.950 830.550 414.450 ;
        RECT 818.550 412.050 830.550 412.950 ;
        RECT 811.950 410.550 812.850 411.300 ;
        RECT 818.550 410.550 819.600 412.050 ;
        RECT 831.450 411.750 833.250 413.550 ;
        RECT 835.050 412.050 836.250 414.450 ;
        RECT 844.950 413.850 847.050 415.950 ;
        RECT 845.100 412.050 846.900 413.850 ;
        RECT 801.150 409.200 811.050 410.250 ;
        RECT 811.950 409.200 819.600 410.550 ;
        RECT 820.950 409.350 824.850 411.150 ;
        RECT 796.200 405.600 797.700 409.200 ;
        RECT 810.000 408.300 811.050 409.200 ;
        RECT 820.950 409.050 823.050 409.350 ;
        RECT 828.150 408.300 829.950 408.750 ;
        RECT 831.450 408.300 832.500 411.750 ;
        RECT 835.050 411.000 846.900 412.050 ;
        RECT 848.100 410.100 849.300 423.600 ;
        RECT 802.350 406.500 809.100 408.300 ;
        RECT 810.000 406.500 816.900 408.300 ;
        RECT 828.150 407.850 832.500 408.300 ;
        RECT 824.850 407.100 832.500 407.850 ;
        RECT 834.000 409.200 849.300 410.100 ;
        RECT 824.850 406.950 829.950 407.100 ;
        RECT 824.850 405.600 825.750 406.950 ;
        RECT 834.000 406.050 835.050 409.200 ;
        RECT 843.300 407.700 845.100 408.300 ;
        RECT 787.650 399.750 789.450 405.600 ;
        RECT 793.050 399.750 794.850 405.600 ;
        RECT 796.200 404.400 800.400 405.600 ;
        RECT 798.600 399.750 800.400 404.400 ;
        RECT 802.950 403.500 805.050 405.600 ;
        RECT 805.950 403.500 808.050 405.600 ;
        RECT 808.950 403.500 811.050 405.600 ;
        RECT 813.750 405.300 815.850 405.600 ;
        RECT 803.250 399.750 805.050 403.500 ;
        RECT 806.250 399.750 808.050 403.500 ;
        RECT 809.250 399.750 811.050 403.500 ;
        RECT 813.000 403.500 815.850 405.300 ;
        RECT 817.950 405.300 820.050 405.600 ;
        RECT 817.950 403.500 820.800 405.300 ;
        RECT 821.700 404.250 825.750 405.600 ;
        RECT 821.700 403.800 823.500 404.250 ;
        RECT 826.950 403.950 829.050 406.050 ;
        RECT 829.950 403.950 832.050 406.050 ;
        RECT 832.950 403.950 835.050 406.050 ;
        RECT 836.700 406.500 845.100 407.700 ;
        RECT 836.700 405.600 838.200 406.500 ;
        RECT 848.100 405.600 849.300 409.200 ;
        RECT 813.000 399.750 814.800 403.500 ;
        RECT 816.000 399.750 817.800 402.600 ;
        RECT 819.000 399.750 820.800 403.500 ;
        RECT 826.950 402.600 828.300 403.950 ;
        RECT 829.950 402.600 831.300 403.950 ;
        RECT 832.950 402.600 834.300 403.950 ;
        RECT 823.500 399.750 825.300 402.600 ;
        RECT 826.500 399.750 828.300 402.600 ;
        RECT 829.500 399.750 831.300 402.600 ;
        RECT 832.500 399.750 834.300 402.600 ;
        RECT 836.700 399.750 838.500 405.600 ;
        RECT 842.100 399.750 843.900 405.600 ;
        RECT 847.500 399.750 849.300 405.600 ;
        RECT 8.850 388.200 10.650 395.250 ;
        RECT 13.350 389.400 15.150 395.250 ;
        RECT 20.550 392.400 22.350 395.250 ;
        RECT 23.550 392.400 25.350 395.250 ;
        RECT 8.850 387.300 12.450 388.200 ;
        RECT 8.100 381.150 9.900 382.950 ;
        RECT 7.950 379.050 10.050 381.150 ;
        RECT 11.250 379.950 12.450 387.300 ;
        RECT 19.950 383.850 22.050 385.950 ;
        RECT 23.400 384.150 24.600 392.400 ;
        RECT 35.850 388.200 37.650 395.250 ;
        RECT 40.350 389.400 42.150 395.250 ;
        RECT 50.850 388.200 52.650 395.250 ;
        RECT 55.350 389.400 57.150 395.250 ;
        RECT 62.850 389.400 64.650 395.250 ;
        RECT 67.350 388.200 69.150 395.250 ;
        RECT 76.650 392.400 78.450 395.250 ;
        RECT 79.650 392.400 81.450 395.250 ;
        RECT 82.650 392.400 84.450 395.250 ;
        RECT 92.550 392.400 94.350 395.250 ;
        RECT 95.550 392.400 97.350 395.250 ;
        RECT 98.550 392.400 100.350 395.250 ;
        RECT 110.550 392.400 112.350 395.250 ;
        RECT 113.550 392.400 115.350 395.250 ;
        RECT 116.550 392.400 118.350 395.250 ;
        RECT 124.650 392.400 126.450 395.250 ;
        RECT 127.650 392.400 129.450 395.250 ;
        RECT 130.650 392.400 132.450 395.250 ;
        RECT 35.850 387.300 39.450 388.200 ;
        RECT 50.850 387.300 54.450 388.200 ;
        RECT 14.100 381.150 15.900 382.950 ;
        RECT 20.100 382.050 21.900 383.850 ;
        RECT 22.950 382.050 25.050 384.150 ;
        RECT 10.950 377.850 13.050 379.950 ;
        RECT 13.950 379.050 16.050 381.150 ;
        RECT 11.250 369.600 12.450 377.850 ;
        RECT 23.400 369.600 24.600 382.050 ;
        RECT 35.100 381.150 36.900 382.950 ;
        RECT 34.950 379.050 37.050 381.150 ;
        RECT 38.250 379.950 39.450 387.300 ;
        RECT 41.100 381.150 42.900 382.950 ;
        RECT 50.100 381.150 51.900 382.950 ;
        RECT 37.950 377.850 40.050 379.950 ;
        RECT 40.950 379.050 43.050 381.150 ;
        RECT 49.950 379.050 52.050 381.150 ;
        RECT 53.250 379.950 54.450 387.300 ;
        RECT 65.550 387.300 69.150 388.200 ;
        RECT 56.100 381.150 57.900 382.950 ;
        RECT 62.100 381.150 63.900 382.950 ;
        RECT 52.950 377.850 55.050 379.950 ;
        RECT 55.950 379.050 58.050 381.150 ;
        RECT 61.950 379.050 64.050 381.150 ;
        RECT 65.550 379.950 66.750 387.300 ;
        RECT 79.950 385.950 81.000 392.400 ;
        RECT 96.000 385.950 97.050 392.400 ;
        RECT 114.000 385.950 115.050 392.400 ;
        RECT 79.950 383.850 82.050 385.950 ;
        RECT 94.950 383.850 97.050 385.950 ;
        RECT 112.950 383.850 115.050 385.950 ;
        RECT 68.100 381.150 69.900 382.950 ;
        RECT 64.950 377.850 67.050 379.950 ;
        RECT 67.950 379.050 70.050 381.150 ;
        RECT 76.950 380.850 79.050 382.950 ;
        RECT 77.100 379.050 78.900 380.850 ;
        RECT 38.250 369.600 39.450 377.850 ;
        RECT 53.250 369.600 54.450 377.850 ;
        RECT 65.550 369.600 66.750 377.850 ;
        RECT 79.950 376.650 81.000 383.850 ;
        RECT 82.950 380.850 85.050 382.950 ;
        RECT 91.950 380.850 94.050 382.950 ;
        RECT 83.100 379.050 84.900 380.850 ;
        RECT 92.100 379.050 93.900 380.850 ;
        RECT 78.450 375.600 81.000 376.650 ;
        RECT 96.000 376.650 97.050 383.850 ;
        RECT 97.950 380.850 100.050 382.950 ;
        RECT 109.950 380.850 112.050 382.950 ;
        RECT 98.100 379.050 99.900 380.850 ;
        RECT 110.100 379.050 111.900 380.850 ;
        RECT 114.000 376.650 115.050 383.850 ;
        RECT 127.950 385.950 129.000 392.400 ;
        RECT 140.850 389.400 142.650 395.250 ;
        RECT 145.350 388.200 147.150 395.250 ;
        RECT 160.650 392.400 162.450 395.250 ;
        RECT 163.650 392.400 165.450 395.250 ;
        RECT 143.550 387.300 147.150 388.200 ;
        RECT 127.950 383.850 130.050 385.950 ;
        RECT 115.950 380.850 118.050 382.950 ;
        RECT 124.950 380.850 127.050 382.950 ;
        RECT 116.100 379.050 117.900 380.850 ;
        RECT 125.100 379.050 126.900 380.850 ;
        RECT 127.950 376.650 129.000 383.850 ;
        RECT 130.950 380.850 133.050 382.950 ;
        RECT 140.100 381.150 141.900 382.950 ;
        RECT 131.100 379.050 132.900 380.850 ;
        RECT 139.950 379.050 142.050 381.150 ;
        RECT 143.550 379.950 144.750 387.300 ;
        RECT 161.400 384.150 162.600 392.400 ;
        RECT 170.850 389.400 172.650 395.250 ;
        RECT 175.350 388.200 177.150 395.250 ;
        RECT 185.850 389.400 187.650 395.250 ;
        RECT 190.350 388.200 192.150 395.250 ;
        RECT 173.550 387.300 177.150 388.200 ;
        RECT 188.550 387.300 192.150 388.200 ;
        RECT 203.550 387.900 205.350 395.250 ;
        RECT 208.050 389.400 209.850 395.250 ;
        RECT 211.050 390.900 212.850 395.250 ;
        RECT 211.050 389.400 214.350 390.900 ;
        RECT 218.850 389.400 220.650 395.250 ;
        RECT 209.250 387.900 211.050 388.500 ;
        RECT 146.100 381.150 147.900 382.950 ;
        RECT 160.950 382.050 163.050 384.150 ;
        RECT 163.950 383.850 166.050 385.950 ;
        RECT 164.100 382.050 165.900 383.850 ;
        RECT 142.950 377.850 145.050 379.950 ;
        RECT 145.950 379.050 148.050 381.150 ;
        RECT 96.000 375.600 98.550 376.650 ;
        RECT 114.000 375.600 116.550 376.650 ;
        RECT 7.650 363.750 9.450 369.600 ;
        RECT 10.650 363.750 12.450 369.600 ;
        RECT 13.650 363.750 15.450 369.600 ;
        RECT 20.550 363.750 22.350 369.600 ;
        RECT 23.550 363.750 25.350 369.600 ;
        RECT 34.650 363.750 36.450 369.600 ;
        RECT 37.650 363.750 39.450 369.600 ;
        RECT 40.650 363.750 42.450 369.600 ;
        RECT 49.650 363.750 51.450 369.600 ;
        RECT 52.650 363.750 54.450 369.600 ;
        RECT 55.650 363.750 57.450 369.600 ;
        RECT 62.550 363.750 64.350 369.600 ;
        RECT 65.550 363.750 67.350 369.600 ;
        RECT 68.550 363.750 70.350 369.600 ;
        RECT 78.450 363.750 80.250 375.600 ;
        RECT 82.650 363.750 84.450 375.600 ;
        RECT 92.550 363.750 94.350 375.600 ;
        RECT 96.750 363.750 98.550 375.600 ;
        RECT 110.550 363.750 112.350 375.600 ;
        RECT 114.750 363.750 116.550 375.600 ;
        RECT 126.450 375.600 129.000 376.650 ;
        RECT 126.450 363.750 128.250 375.600 ;
        RECT 130.650 363.750 132.450 375.600 ;
        RECT 143.550 369.600 144.750 377.850 ;
        RECT 145.950 375.450 148.050 376.050 ;
        RECT 157.950 375.450 160.050 376.050 ;
        RECT 145.950 374.550 160.050 375.450 ;
        RECT 145.950 373.950 148.050 374.550 ;
        RECT 157.950 373.950 160.050 374.550 ;
        RECT 161.400 369.600 162.600 382.050 ;
        RECT 170.100 381.150 171.900 382.950 ;
        RECT 169.950 379.050 172.050 381.150 ;
        RECT 173.550 379.950 174.750 387.300 ;
        RECT 176.100 381.150 177.900 382.950 ;
        RECT 185.100 381.150 186.900 382.950 ;
        RECT 172.950 377.850 175.050 379.950 ;
        RECT 175.950 379.050 178.050 381.150 ;
        RECT 184.950 379.050 187.050 381.150 ;
        RECT 188.550 379.950 189.750 387.300 ;
        RECT 203.550 386.700 211.050 387.900 ;
        RECT 191.100 381.150 192.900 382.950 ;
        RECT 187.950 377.850 190.050 379.950 ;
        RECT 190.950 379.050 193.050 381.150 ;
        RECT 202.950 380.850 205.050 382.950 ;
        RECT 203.100 379.050 204.900 380.850 ;
        RECT 163.950 375.450 166.050 376.050 ;
        RECT 169.950 375.450 172.050 376.050 ;
        RECT 163.950 374.550 172.050 375.450 ;
        RECT 163.950 373.950 166.050 374.550 ;
        RECT 169.950 373.950 172.050 374.550 ;
        RECT 173.550 369.600 174.750 377.850 ;
        RECT 188.550 369.600 189.750 377.850 ;
        RECT 206.700 369.600 207.900 386.700 ;
        RECT 213.150 382.950 214.350 389.400 ;
        RECT 223.350 388.200 225.150 395.250 ;
        RECT 231.000 389.400 232.800 395.250 ;
        RECT 235.200 391.050 237.000 395.250 ;
        RECT 238.500 392.400 240.300 395.250 ;
        RECT 235.200 389.400 240.900 391.050 ;
        RECT 247.650 389.400 249.450 395.250 ;
        RECT 221.550 387.300 225.150 388.200 ;
        RECT 209.100 381.150 210.900 382.950 ;
        RECT 208.950 379.050 211.050 381.150 ;
        RECT 211.950 380.850 214.350 382.950 ;
        RECT 218.100 381.150 219.900 382.950 ;
        RECT 213.150 375.600 214.350 380.850 ;
        RECT 217.950 379.050 220.050 381.150 ;
        RECT 221.550 379.950 222.750 387.300 ;
        RECT 230.100 384.150 231.900 385.950 ;
        RECT 224.100 381.150 225.900 382.950 ;
        RECT 229.950 382.050 232.050 384.150 ;
        RECT 232.950 383.850 235.050 385.950 ;
        RECT 236.100 384.150 237.900 385.950 ;
        RECT 233.100 382.050 234.900 383.850 ;
        RECT 235.950 382.050 238.050 384.150 ;
        RECT 239.700 382.950 240.900 389.400 ;
        RECT 248.250 387.300 249.450 389.400 ;
        RECT 250.650 390.300 252.450 395.250 ;
        RECT 253.650 391.200 255.450 395.250 ;
        RECT 256.650 390.300 258.450 395.250 ;
        RECT 250.650 388.950 258.450 390.300 ;
        RECT 268.650 394.500 276.450 395.250 ;
        RECT 268.650 389.400 270.450 394.500 ;
        RECT 271.650 389.400 273.450 393.600 ;
        RECT 274.650 390.000 276.450 394.500 ;
        RECT 277.650 390.900 279.450 395.250 ;
        RECT 280.650 390.000 282.450 395.250 ;
        RECT 272.250 387.900 273.150 389.400 ;
        RECT 274.650 389.100 282.450 390.000 ;
        RECT 292.650 389.400 294.450 395.250 ;
        RECT 248.250 386.250 252.000 387.300 ;
        RECT 272.250 386.850 276.600 387.900 ;
        RECT 250.950 382.950 252.150 386.250 ;
        RECT 254.100 384.150 255.900 385.950 ;
        RECT 272.700 384.150 274.500 385.950 ;
        RECT 220.950 377.850 223.050 379.950 ;
        RECT 223.950 379.050 226.050 381.150 ;
        RECT 238.950 380.850 241.050 382.950 ;
        RECT 250.950 380.850 253.050 382.950 ;
        RECT 253.950 382.050 256.050 384.150 ;
        RECT 256.950 380.850 259.050 382.950 ;
        RECT 268.950 380.850 271.050 382.950 ;
        RECT 271.950 382.050 274.050 384.150 ;
        RECT 275.400 382.950 276.600 386.850 ;
        RECT 293.250 387.300 294.450 389.400 ;
        RECT 295.650 390.300 297.450 395.250 ;
        RECT 298.650 391.200 300.450 395.250 ;
        RECT 301.650 390.300 303.450 395.250 ;
        RECT 311.550 392.400 313.350 395.250 ;
        RECT 314.550 392.400 316.350 395.250 ;
        RECT 295.650 388.950 303.450 390.300 ;
        RECT 293.250 386.250 297.000 387.300 ;
        RECT 278.100 384.150 279.900 385.950 ;
        RECT 274.950 380.850 277.050 382.950 ;
        RECT 277.950 382.050 280.050 384.150 ;
        RECT 295.950 382.950 297.150 386.250 ;
        RECT 299.100 384.150 300.900 385.950 ;
        RECT 280.950 380.850 283.050 382.950 ;
        RECT 295.950 380.850 298.050 382.950 ;
        RECT 298.950 382.050 301.050 384.150 ;
        RECT 310.950 383.850 313.050 385.950 ;
        RECT 314.400 384.150 315.600 392.400 ;
        RECT 323.550 389.400 325.350 395.250 ;
        RECT 326.550 389.400 328.350 395.250 ;
        RECT 334.650 392.400 336.450 395.250 ;
        RECT 337.650 392.400 339.450 395.250 ;
        RECT 340.650 392.400 342.450 395.250 ;
        RECT 352.650 392.400 354.450 395.250 ;
        RECT 355.650 392.400 357.450 395.250 ;
        RECT 358.650 392.400 360.450 395.250 ;
        RECT 371.700 392.400 373.500 395.250 ;
        RECT 323.100 384.150 324.900 385.950 ;
        RECT 301.950 380.850 304.050 382.950 ;
        RECT 311.100 382.050 312.900 383.850 ;
        RECT 313.950 382.050 316.050 384.150 ;
        RECT 322.950 382.050 325.050 384.150 ;
        RECT 326.400 382.950 327.600 389.400 ;
        RECT 337.950 385.950 339.000 392.400 ;
        RECT 355.950 385.950 357.000 392.400 ;
        RECT 375.000 391.050 376.800 395.250 ;
        RECT 371.100 389.400 376.800 391.050 ;
        RECT 379.200 389.400 381.000 395.250 ;
        RECT 389.550 392.400 391.350 395.250 ;
        RECT 392.550 392.400 394.350 395.250 ;
        RECT 395.550 392.400 397.350 395.250 ;
        RECT 402.750 392.400 404.550 395.250 ;
        RECT 405.750 392.400 407.550 395.250 ;
        RECT 337.950 383.850 340.050 385.950 ;
        RECT 355.950 383.850 358.050 385.950 ;
        RECT 140.550 363.750 142.350 369.600 ;
        RECT 143.550 363.750 145.350 369.600 ;
        RECT 146.550 363.750 148.350 369.600 ;
        RECT 160.650 363.750 162.450 369.600 ;
        RECT 163.650 363.750 165.450 369.600 ;
        RECT 170.550 363.750 172.350 369.600 ;
        RECT 173.550 363.750 175.350 369.600 ;
        RECT 176.550 363.750 178.350 369.600 ;
        RECT 185.550 363.750 187.350 369.600 ;
        RECT 188.550 363.750 190.350 369.600 ;
        RECT 191.550 363.750 193.350 369.600 ;
        RECT 203.550 363.750 205.350 369.600 ;
        RECT 206.550 363.750 208.350 369.600 ;
        RECT 210.150 363.750 211.950 375.600 ;
        RECT 213.150 363.750 214.950 375.600 ;
        RECT 221.550 369.600 222.750 377.850 ;
        RECT 239.700 375.600 240.900 380.850 ;
        RECT 247.950 377.850 250.050 379.950 ;
        RECT 248.250 376.050 250.050 377.850 ;
        RECT 251.850 375.600 253.050 380.850 ;
        RECT 257.100 379.050 258.900 380.850 ;
        RECT 269.250 379.050 271.050 380.850 ;
        RECT 275.250 375.600 276.450 380.850 ;
        RECT 281.100 379.050 282.900 380.850 ;
        RECT 292.950 377.850 295.050 379.950 ;
        RECT 293.250 376.050 295.050 377.850 ;
        RECT 296.850 375.600 298.050 380.850 ;
        RECT 302.100 379.050 303.900 380.850 ;
        RECT 230.550 374.700 238.350 375.600 ;
        RECT 218.550 363.750 220.350 369.600 ;
        RECT 221.550 363.750 223.350 369.600 ;
        RECT 224.550 363.750 226.350 369.600 ;
        RECT 230.550 363.750 232.350 374.700 ;
        RECT 233.550 363.750 235.350 373.800 ;
        RECT 236.550 363.750 238.350 374.700 ;
        RECT 239.550 363.750 241.350 375.600 ;
        RECT 248.400 363.750 250.200 369.600 ;
        RECT 251.700 363.750 253.500 375.600 ;
        RECT 255.900 363.750 257.700 375.600 ;
        RECT 270.150 363.750 271.950 375.600 ;
        RECT 274.650 363.750 277.950 375.600 ;
        RECT 280.650 363.750 282.450 375.600 ;
        RECT 293.400 363.750 295.200 369.600 ;
        RECT 296.700 363.750 298.500 375.600 ;
        RECT 300.900 363.750 302.700 375.600 ;
        RECT 314.400 369.600 315.600 382.050 ;
        RECT 325.950 380.850 328.050 382.950 ;
        RECT 334.950 380.850 337.050 382.950 ;
        RECT 326.400 375.600 327.600 380.850 ;
        RECT 335.100 379.050 336.900 380.850 ;
        RECT 337.950 376.650 339.000 383.850 ;
        RECT 340.950 380.850 343.050 382.950 ;
        RECT 352.950 380.850 355.050 382.950 ;
        RECT 341.100 379.050 342.900 380.850 ;
        RECT 353.100 379.050 354.900 380.850 ;
        RECT 355.950 376.650 357.000 383.850 ;
        RECT 371.100 382.950 372.300 389.400 ;
        RECT 393.000 385.950 394.050 392.400 ;
        RECT 374.100 384.150 375.900 385.950 ;
        RECT 358.950 380.850 361.050 382.950 ;
        RECT 370.950 380.850 373.050 382.950 ;
        RECT 373.950 382.050 376.050 384.150 ;
        RECT 376.950 383.850 379.050 385.950 ;
        RECT 380.100 384.150 381.900 385.950 ;
        RECT 377.100 382.050 378.900 383.850 ;
        RECT 379.950 382.050 382.050 384.150 ;
        RECT 391.950 383.850 394.050 385.950 ;
        RECT 406.050 384.150 407.550 392.400 ;
        RECT 388.950 380.850 391.050 382.950 ;
        RECT 359.100 379.050 360.900 380.850 ;
        RECT 336.450 375.600 339.000 376.650 ;
        RECT 354.450 375.600 357.000 376.650 ;
        RECT 371.100 375.600 372.300 380.850 ;
        RECT 389.100 379.050 390.900 380.850 ;
        RECT 393.000 376.650 394.050 383.850 ;
        RECT 394.950 380.850 397.050 382.950 ;
        RECT 403.950 382.050 407.550 384.150 ;
        RECT 395.100 379.050 396.900 380.850 ;
        RECT 393.000 375.600 395.550 376.650 ;
        RECT 311.550 363.750 313.350 369.600 ;
        RECT 314.550 363.750 316.350 369.600 ;
        RECT 323.550 363.750 325.350 375.600 ;
        RECT 326.550 363.750 328.350 375.600 ;
        RECT 336.450 363.750 338.250 375.600 ;
        RECT 340.650 363.750 342.450 375.600 ;
        RECT 354.450 363.750 356.250 375.600 ;
        RECT 358.650 363.750 360.450 375.600 ;
        RECT 370.650 363.750 372.450 375.600 ;
        RECT 373.650 374.700 381.450 375.600 ;
        RECT 373.650 363.750 375.450 374.700 ;
        RECT 376.650 363.750 378.450 373.800 ;
        RECT 379.650 363.750 381.450 374.700 ;
        RECT 389.550 363.750 391.350 375.600 ;
        RECT 393.750 363.750 395.550 375.600 ;
        RECT 406.050 369.600 407.550 382.050 ;
        RECT 409.650 389.400 411.450 395.250 ;
        RECT 415.050 389.400 416.850 395.250 ;
        RECT 420.600 390.600 422.400 395.250 ;
        RECT 425.250 391.500 427.050 395.250 ;
        RECT 428.250 391.500 430.050 395.250 ;
        RECT 431.250 391.500 433.050 395.250 ;
        RECT 418.200 389.400 422.400 390.600 ;
        RECT 424.950 389.400 427.050 391.500 ;
        RECT 427.950 389.400 430.050 391.500 ;
        RECT 430.950 389.400 433.050 391.500 ;
        RECT 435.000 391.500 436.800 395.250 ;
        RECT 438.000 392.400 439.800 395.250 ;
        RECT 441.000 391.500 442.800 395.250 ;
        RECT 445.500 392.400 447.300 395.250 ;
        RECT 448.500 392.400 450.300 395.250 ;
        RECT 451.500 392.400 453.300 395.250 ;
        RECT 454.500 392.400 456.300 395.250 ;
        RECT 435.000 389.700 437.850 391.500 ;
        RECT 435.750 389.400 437.850 389.700 ;
        RECT 439.950 389.700 442.800 391.500 ;
        RECT 443.700 390.750 445.500 391.200 ;
        RECT 448.950 391.050 450.300 392.400 ;
        RECT 451.950 391.050 453.300 392.400 ;
        RECT 454.950 391.050 456.300 392.400 ;
        RECT 439.950 389.400 442.050 389.700 ;
        RECT 443.700 389.400 447.750 390.750 ;
        RECT 409.650 374.550 410.850 389.400 ;
        RECT 418.200 385.800 419.700 389.400 ;
        RECT 424.350 386.700 431.100 388.500 ;
        RECT 432.000 386.700 438.900 388.500 ;
        RECT 446.850 388.050 447.750 389.400 ;
        RECT 448.950 388.950 451.050 391.050 ;
        RECT 451.950 388.950 454.050 391.050 ;
        RECT 454.950 388.950 457.050 391.050 ;
        RECT 446.850 387.900 451.950 388.050 ;
        RECT 446.850 387.150 454.500 387.900 ;
        RECT 450.150 386.700 454.500 387.150 ;
        RECT 432.000 385.800 433.050 386.700 ;
        RECT 450.150 386.250 451.950 386.700 ;
        RECT 411.900 384.000 419.700 385.800 ;
        RECT 423.150 384.750 433.050 385.800 ;
        RECT 423.150 382.950 424.200 384.750 ;
        RECT 433.950 384.450 441.600 385.800 ;
        RECT 433.950 383.700 434.850 384.450 ;
        RECT 415.950 381.900 424.200 382.950 ;
        RECT 425.250 382.650 434.850 383.700 ;
        RECT 415.950 377.850 418.050 381.900 ;
        RECT 425.250 381.000 426.150 382.650 ;
        RECT 435.750 381.750 439.650 383.550 ;
        RECT 440.550 382.950 441.600 384.450 ;
        RECT 442.950 385.650 445.050 385.950 ;
        RECT 442.950 383.850 446.850 385.650 ;
        RECT 453.450 383.250 454.500 386.700 ;
        RECT 456.000 385.800 457.050 388.950 ;
        RECT 458.700 389.400 460.500 395.250 ;
        RECT 464.100 389.400 465.900 395.250 ;
        RECT 469.500 389.400 471.300 395.250 ;
        RECT 479.550 392.400 481.350 395.250 ;
        RECT 482.550 392.400 484.350 395.250 ;
        RECT 485.550 392.400 487.350 395.250 ;
        RECT 458.700 388.500 460.200 389.400 ;
        RECT 458.700 387.300 467.100 388.500 ;
        RECT 465.300 386.700 467.100 387.300 ;
        RECT 470.100 385.800 471.300 389.400 ;
        RECT 483.000 385.950 484.050 392.400 ;
        RECT 491.550 387.900 493.350 395.250 ;
        RECT 496.050 389.400 497.850 395.250 ;
        RECT 499.050 390.900 500.850 395.250 ;
        RECT 512.550 392.400 514.350 395.250 ;
        RECT 499.050 389.400 502.350 390.900 ;
        RECT 497.250 387.900 499.050 388.500 ;
        RECT 491.550 386.700 499.050 387.900 ;
        RECT 456.000 384.900 471.300 385.800 ;
        RECT 440.550 382.050 452.550 382.950 ;
        RECT 419.100 379.200 426.150 381.000 ;
        RECT 427.500 379.950 429.300 381.750 ;
        RECT 435.750 381.450 437.850 381.750 ;
        RECT 439.950 380.550 442.050 380.850 ;
        RECT 448.800 380.550 450.600 381.150 ;
        RECT 439.950 379.950 450.600 380.550 ;
        RECT 427.500 379.350 450.600 379.950 ;
        RECT 451.500 380.550 452.550 382.050 ;
        RECT 453.450 381.450 455.250 383.250 ;
        RECT 457.050 382.950 468.900 384.000 ;
        RECT 457.050 380.550 458.250 382.950 ;
        RECT 467.100 381.150 468.900 382.950 ;
        RECT 451.500 379.650 458.250 380.550 ;
        RECT 460.950 379.650 463.050 379.950 ;
        RECT 427.500 378.750 442.050 379.350 ;
        RECT 459.150 378.450 463.050 379.650 ;
        RECT 466.950 379.050 469.050 381.150 ;
        RECT 449.100 377.850 463.050 378.450 ;
        RECT 423.000 377.550 462.750 377.850 ;
        RECT 411.750 376.650 413.550 377.250 ;
        RECT 423.000 376.650 451.050 377.550 ;
        RECT 411.750 375.450 424.050 376.650 ;
        RECT 451.950 376.050 454.050 376.350 ;
        RECT 461.700 376.050 463.500 376.650 ;
        RECT 424.950 374.550 427.050 375.750 ;
        RECT 409.650 373.650 427.050 374.550 ;
        RECT 430.950 374.400 451.050 375.750 ;
        RECT 430.950 373.650 433.050 374.400 ;
        RECT 412.500 369.600 413.700 373.650 ;
        RECT 414.600 371.700 416.400 372.300 ;
        RECT 421.350 372.150 423.150 372.300 ;
        RECT 414.600 370.500 420.300 371.700 ;
        RECT 421.350 370.950 430.050 372.150 ;
        RECT 421.350 370.500 423.150 370.950 ;
        RECT 402.750 363.750 404.550 369.600 ;
        RECT 405.750 363.750 407.550 369.600 ;
        RECT 409.500 363.750 411.300 369.600 ;
        RECT 412.500 363.750 414.300 369.600 ;
        RECT 415.500 363.750 417.300 369.600 ;
        RECT 418.500 363.750 420.300 370.500 ;
        RECT 427.950 370.050 430.050 370.950 ;
        RECT 421.500 363.750 423.300 369.600 ;
        RECT 424.800 367.800 426.900 369.900 ;
        RECT 425.400 366.600 426.900 367.800 ;
        RECT 425.250 363.750 427.050 366.600 ;
        RECT 428.250 363.750 430.050 370.050 ;
        RECT 431.550 366.600 432.900 373.650 ;
        RECT 449.100 373.350 451.050 374.400 ;
        RECT 451.950 374.850 463.500 376.050 ;
        RECT 451.950 374.250 454.050 374.850 ;
        RECT 465.000 373.350 466.800 374.100 ;
        RECT 434.100 370.800 438.000 372.600 ;
        RECT 435.000 370.500 438.000 370.800 ;
        RECT 439.950 372.150 442.050 372.600 ;
        RECT 449.100 372.300 466.800 373.350 ;
        RECT 439.950 370.500 442.350 372.150 ;
        RECT 431.250 363.750 433.050 366.600 ;
        RECT 435.000 363.750 436.800 370.500 ;
        RECT 441.000 369.600 442.350 370.500 ;
        RECT 448.950 369.600 451.050 370.050 ;
        RECT 438.000 363.750 439.800 369.600 ;
        RECT 441.000 363.750 442.800 369.600 ;
        RECT 444.750 363.750 446.550 369.600 ;
        RECT 448.500 367.950 451.050 369.600 ;
        RECT 451.950 367.950 454.050 370.050 ;
        RECT 454.950 367.950 457.050 370.050 ;
        RECT 448.500 366.600 449.700 367.950 ;
        RECT 451.950 366.600 452.850 367.950 ;
        RECT 454.950 366.600 456.150 367.950 ;
        RECT 447.750 363.750 449.700 366.600 ;
        RECT 450.750 363.750 452.850 366.600 ;
        RECT 453.750 363.750 456.150 366.600 ;
        RECT 457.500 363.750 459.300 367.050 ;
        RECT 460.500 363.750 462.300 372.300 ;
        RECT 470.100 371.400 471.300 384.900 ;
        RECT 481.950 383.850 484.050 385.950 ;
        RECT 478.950 380.850 481.050 382.950 ;
        RECT 479.100 379.050 480.900 380.850 ;
        RECT 483.000 376.650 484.050 383.850 ;
        RECT 484.950 380.850 487.050 382.950 ;
        RECT 490.950 380.850 493.050 382.950 ;
        RECT 485.100 379.050 486.900 380.850 ;
        RECT 491.100 379.050 492.900 380.850 ;
        RECT 483.000 375.600 485.550 376.650 ;
        RECT 467.250 370.500 471.300 371.400 ;
        RECT 467.250 369.600 468.300 370.500 ;
        RECT 463.500 363.750 465.300 369.600 ;
        RECT 466.500 363.750 468.300 369.600 ;
        RECT 469.500 363.750 471.300 369.600 ;
        RECT 479.550 363.750 481.350 375.600 ;
        RECT 483.750 363.750 485.550 375.600 ;
        RECT 494.700 369.600 495.900 386.700 ;
        RECT 501.150 382.950 502.350 389.400 ;
        RECT 513.150 388.500 514.350 392.400 ;
        RECT 515.850 389.400 517.650 395.250 ;
        RECT 518.850 389.400 520.650 395.250 ;
        RECT 513.150 387.600 518.250 388.500 ;
        RECT 516.000 386.700 518.250 387.600 ;
        RECT 497.100 381.150 498.900 382.950 ;
        RECT 496.950 379.050 499.050 381.150 ;
        RECT 499.950 380.850 502.350 382.950 ;
        RECT 511.950 380.850 514.050 382.950 ;
        RECT 501.150 375.600 502.350 380.850 ;
        RECT 512.100 379.050 513.900 380.850 ;
        RECT 516.000 378.300 517.050 386.700 ;
        RECT 519.150 382.950 520.350 389.400 ;
        RECT 530.700 386.400 532.500 395.250 ;
        RECT 536.100 387.000 537.900 395.250 ;
        RECT 546.750 392.400 548.550 395.250 ;
        RECT 549.750 392.400 551.550 395.250 ;
        RECT 536.100 385.350 540.600 387.000 ;
        RECT 517.950 380.850 520.350 382.950 ;
        RECT 539.400 381.150 540.600 385.350 ;
        RECT 550.050 384.150 551.550 392.400 ;
        RECT 547.950 382.050 551.550 384.150 ;
        RECT 516.000 377.400 518.250 378.300 ;
        RECT 512.550 376.500 518.250 377.400 ;
        RECT 491.550 363.750 493.350 369.600 ;
        RECT 494.550 363.750 496.350 369.600 ;
        RECT 498.150 363.750 499.950 375.600 ;
        RECT 501.150 363.750 502.950 375.600 ;
        RECT 512.550 369.600 513.750 376.500 ;
        RECT 519.150 375.600 520.350 380.850 ;
        RECT 529.950 377.850 532.050 379.950 ;
        RECT 535.950 377.850 538.050 379.950 ;
        RECT 538.950 379.050 541.050 381.150 ;
        RECT 530.100 376.050 531.900 377.850 ;
        RECT 512.550 363.750 514.350 369.600 ;
        RECT 515.850 363.750 517.650 375.600 ;
        RECT 518.850 363.750 520.650 375.600 ;
        RECT 532.950 374.850 535.050 376.950 ;
        RECT 536.250 376.050 538.050 377.850 ;
        RECT 533.100 373.050 534.900 374.850 ;
        RECT 539.700 370.800 540.750 379.050 ;
        RECT 533.700 369.900 540.750 370.800 ;
        RECT 533.700 369.600 535.350 369.900 ;
        RECT 530.550 363.750 532.350 369.600 ;
        RECT 533.550 363.750 535.350 369.600 ;
        RECT 539.550 369.600 540.750 369.900 ;
        RECT 550.050 369.600 551.550 382.050 ;
        RECT 553.650 389.400 555.450 395.250 ;
        RECT 559.050 389.400 560.850 395.250 ;
        RECT 564.600 390.600 566.400 395.250 ;
        RECT 569.250 391.500 571.050 395.250 ;
        RECT 572.250 391.500 574.050 395.250 ;
        RECT 575.250 391.500 577.050 395.250 ;
        RECT 562.200 389.400 566.400 390.600 ;
        RECT 568.950 389.400 571.050 391.500 ;
        RECT 571.950 389.400 574.050 391.500 ;
        RECT 574.950 389.400 577.050 391.500 ;
        RECT 579.000 391.500 580.800 395.250 ;
        RECT 582.000 392.400 583.800 395.250 ;
        RECT 585.000 391.500 586.800 395.250 ;
        RECT 589.500 392.400 591.300 395.250 ;
        RECT 592.500 392.400 594.300 395.250 ;
        RECT 595.500 392.400 597.300 395.250 ;
        RECT 598.500 392.400 600.300 395.250 ;
        RECT 579.000 389.700 581.850 391.500 ;
        RECT 579.750 389.400 581.850 389.700 ;
        RECT 583.950 389.700 586.800 391.500 ;
        RECT 587.700 390.750 589.500 391.200 ;
        RECT 592.950 391.050 594.300 392.400 ;
        RECT 595.950 391.050 597.300 392.400 ;
        RECT 598.950 391.050 600.300 392.400 ;
        RECT 583.950 389.400 586.050 389.700 ;
        RECT 587.700 389.400 591.750 390.750 ;
        RECT 553.650 374.550 554.850 389.400 ;
        RECT 562.200 385.800 563.700 389.400 ;
        RECT 568.350 386.700 575.100 388.500 ;
        RECT 576.000 386.700 582.900 388.500 ;
        RECT 590.850 388.050 591.750 389.400 ;
        RECT 592.950 388.950 595.050 391.050 ;
        RECT 595.950 388.950 598.050 391.050 ;
        RECT 598.950 388.950 601.050 391.050 ;
        RECT 590.850 387.900 595.950 388.050 ;
        RECT 590.850 387.150 598.500 387.900 ;
        RECT 594.150 386.700 598.500 387.150 ;
        RECT 576.000 385.800 577.050 386.700 ;
        RECT 594.150 386.250 595.950 386.700 ;
        RECT 555.900 384.000 563.700 385.800 ;
        RECT 567.150 384.750 577.050 385.800 ;
        RECT 567.150 382.950 568.200 384.750 ;
        RECT 577.950 384.450 585.600 385.800 ;
        RECT 577.950 383.700 578.850 384.450 ;
        RECT 559.950 381.900 568.200 382.950 ;
        RECT 569.250 382.650 578.850 383.700 ;
        RECT 559.950 377.850 562.050 381.900 ;
        RECT 569.250 381.000 570.150 382.650 ;
        RECT 579.750 381.750 583.650 383.550 ;
        RECT 584.550 382.950 585.600 384.450 ;
        RECT 586.950 385.650 589.050 385.950 ;
        RECT 586.950 383.850 590.850 385.650 ;
        RECT 597.450 383.250 598.500 386.700 ;
        RECT 600.000 385.800 601.050 388.950 ;
        RECT 602.700 389.400 604.500 395.250 ;
        RECT 608.100 389.400 609.900 395.250 ;
        RECT 613.500 389.400 615.300 395.250 ;
        RECT 620.550 392.400 622.350 395.250 ;
        RECT 623.550 392.400 625.350 395.250 ;
        RECT 635.700 392.400 637.500 395.250 ;
        RECT 602.700 388.500 604.200 389.400 ;
        RECT 602.700 387.300 611.100 388.500 ;
        RECT 609.300 386.700 611.100 387.300 ;
        RECT 614.100 385.800 615.300 389.400 ;
        RECT 600.000 384.900 615.300 385.800 ;
        RECT 584.550 382.050 596.550 382.950 ;
        RECT 563.100 379.200 570.150 381.000 ;
        RECT 571.500 379.950 573.300 381.750 ;
        RECT 579.750 381.450 581.850 381.750 ;
        RECT 583.950 380.550 586.050 380.850 ;
        RECT 592.800 380.550 594.600 381.150 ;
        RECT 583.950 379.950 594.600 380.550 ;
        RECT 571.500 379.350 594.600 379.950 ;
        RECT 595.500 380.550 596.550 382.050 ;
        RECT 597.450 381.450 599.250 383.250 ;
        RECT 601.050 382.950 612.900 384.000 ;
        RECT 601.050 380.550 602.250 382.950 ;
        RECT 611.100 381.150 612.900 382.950 ;
        RECT 595.500 379.650 602.250 380.550 ;
        RECT 604.950 379.650 607.050 379.950 ;
        RECT 571.500 378.750 586.050 379.350 ;
        RECT 603.150 378.450 607.050 379.650 ;
        RECT 610.950 379.050 613.050 381.150 ;
        RECT 593.100 377.850 607.050 378.450 ;
        RECT 567.000 377.550 606.750 377.850 ;
        RECT 555.750 376.650 557.550 377.250 ;
        RECT 567.000 376.650 595.050 377.550 ;
        RECT 555.750 375.450 568.050 376.650 ;
        RECT 595.950 376.050 598.050 376.350 ;
        RECT 605.700 376.050 607.500 376.650 ;
        RECT 568.950 374.550 571.050 375.750 ;
        RECT 553.650 373.650 571.050 374.550 ;
        RECT 574.950 374.400 595.050 375.750 ;
        RECT 574.950 373.650 577.050 374.400 ;
        RECT 556.500 369.600 557.700 373.650 ;
        RECT 558.600 371.700 560.400 372.300 ;
        RECT 565.350 372.150 567.150 372.300 ;
        RECT 558.600 370.500 564.300 371.700 ;
        RECT 565.350 370.950 574.050 372.150 ;
        RECT 565.350 370.500 567.150 370.950 ;
        RECT 536.550 363.750 538.350 369.000 ;
        RECT 539.550 363.750 541.350 369.600 ;
        RECT 546.750 363.750 548.550 369.600 ;
        RECT 549.750 363.750 551.550 369.600 ;
        RECT 553.500 363.750 555.300 369.600 ;
        RECT 556.500 363.750 558.300 369.600 ;
        RECT 559.500 363.750 561.300 369.600 ;
        RECT 562.500 363.750 564.300 370.500 ;
        RECT 571.950 370.050 574.050 370.950 ;
        RECT 565.500 363.750 567.300 369.600 ;
        RECT 568.800 367.800 570.900 369.900 ;
        RECT 569.400 366.600 570.900 367.800 ;
        RECT 569.250 363.750 571.050 366.600 ;
        RECT 572.250 363.750 574.050 370.050 ;
        RECT 575.550 366.600 576.900 373.650 ;
        RECT 593.100 373.350 595.050 374.400 ;
        RECT 595.950 374.850 607.500 376.050 ;
        RECT 595.950 374.250 598.050 374.850 ;
        RECT 609.000 373.350 610.800 374.100 ;
        RECT 578.100 370.800 582.000 372.600 ;
        RECT 579.000 370.500 582.000 370.800 ;
        RECT 583.950 372.150 586.050 372.600 ;
        RECT 593.100 372.300 610.800 373.350 ;
        RECT 583.950 370.500 586.350 372.150 ;
        RECT 575.250 363.750 577.050 366.600 ;
        RECT 579.000 363.750 580.800 370.500 ;
        RECT 585.000 369.600 586.350 370.500 ;
        RECT 592.950 369.600 595.050 370.050 ;
        RECT 582.000 363.750 583.800 369.600 ;
        RECT 585.000 363.750 586.800 369.600 ;
        RECT 588.750 363.750 590.550 369.600 ;
        RECT 592.500 367.950 595.050 369.600 ;
        RECT 595.950 367.950 598.050 370.050 ;
        RECT 598.950 367.950 601.050 370.050 ;
        RECT 592.500 366.600 593.700 367.950 ;
        RECT 595.950 366.600 596.850 367.950 ;
        RECT 598.950 366.600 600.150 367.950 ;
        RECT 591.750 363.750 593.700 366.600 ;
        RECT 594.750 363.750 596.850 366.600 ;
        RECT 597.750 363.750 600.150 366.600 ;
        RECT 601.500 363.750 603.300 367.050 ;
        RECT 604.500 363.750 606.300 372.300 ;
        RECT 614.100 371.400 615.300 384.900 ;
        RECT 619.950 383.850 622.050 385.950 ;
        RECT 623.400 384.150 624.600 392.400 ;
        RECT 639.000 391.050 640.800 395.250 ;
        RECT 635.100 389.400 640.800 391.050 ;
        RECT 643.200 389.400 645.000 395.250 ;
        RECT 620.100 382.050 621.900 383.850 ;
        RECT 622.950 382.050 625.050 384.150 ;
        RECT 635.100 382.950 636.300 389.400 ;
        RECT 653.100 387.000 654.900 395.250 ;
        RECT 638.100 384.150 639.900 385.950 ;
        RECT 611.250 370.500 615.300 371.400 ;
        RECT 611.250 369.600 612.300 370.500 ;
        RECT 623.400 369.600 624.600 382.050 ;
        RECT 634.950 380.850 637.050 382.950 ;
        RECT 637.950 382.050 640.050 384.150 ;
        RECT 640.950 383.850 643.050 385.950 ;
        RECT 644.100 384.150 645.900 385.950 ;
        RECT 650.400 385.350 654.900 387.000 ;
        RECT 658.500 386.400 660.300 395.250 ;
        RECT 667.650 392.400 669.450 395.250 ;
        RECT 670.650 392.400 672.450 395.250 ;
        RECT 641.100 382.050 642.900 383.850 ;
        RECT 643.950 382.050 646.050 384.150 ;
        RECT 650.400 381.150 651.600 385.350 ;
        RECT 668.400 384.150 669.600 392.400 ;
        RECT 676.350 389.400 678.150 395.250 ;
        RECT 679.350 389.400 681.150 395.250 ;
        RECT 682.650 392.400 684.450 395.250 ;
        RECT 667.950 382.050 670.050 384.150 ;
        RECT 670.950 383.850 673.050 385.950 ;
        RECT 671.100 382.050 672.900 383.850 ;
        RECT 676.650 382.950 677.850 389.400 ;
        RECT 682.650 388.500 683.850 392.400 ;
        RECT 691.650 389.400 693.450 395.250 ;
        RECT 678.750 387.600 683.850 388.500 ;
        RECT 678.750 386.700 681.000 387.600 ;
        RECT 635.100 375.600 636.300 380.850 ;
        RECT 649.950 379.050 652.050 381.150 ;
        RECT 607.500 363.750 609.300 369.600 ;
        RECT 610.500 363.750 612.300 369.600 ;
        RECT 613.500 363.750 615.300 369.600 ;
        RECT 620.550 363.750 622.350 369.600 ;
        RECT 623.550 363.750 625.350 369.600 ;
        RECT 634.650 363.750 636.450 375.600 ;
        RECT 637.650 374.700 645.450 375.600 ;
        RECT 637.650 363.750 639.450 374.700 ;
        RECT 640.650 363.750 642.450 373.800 ;
        RECT 643.650 363.750 645.450 374.700 ;
        RECT 650.250 370.800 651.300 379.050 ;
        RECT 652.950 377.850 655.050 379.950 ;
        RECT 658.950 377.850 661.050 379.950 ;
        RECT 652.950 376.050 654.750 377.850 ;
        RECT 655.950 374.850 658.050 376.950 ;
        RECT 659.100 376.050 660.900 377.850 ;
        RECT 656.100 373.050 657.900 374.850 ;
        RECT 650.250 369.900 657.300 370.800 ;
        RECT 650.250 369.600 651.450 369.900 ;
        RECT 649.650 363.750 651.450 369.600 ;
        RECT 655.650 369.600 657.300 369.900 ;
        RECT 668.400 369.600 669.600 382.050 ;
        RECT 676.650 380.850 679.050 382.950 ;
        RECT 676.650 375.600 677.850 380.850 ;
        RECT 679.950 378.300 681.000 386.700 ;
        RECT 692.250 387.300 693.450 389.400 ;
        RECT 694.650 390.300 696.450 395.250 ;
        RECT 697.650 391.200 699.450 395.250 ;
        RECT 700.650 390.300 702.450 395.250 ;
        RECT 694.650 388.950 702.450 390.300 ;
        RECT 704.700 389.400 706.500 395.250 ;
        RECT 710.100 389.400 711.900 395.250 ;
        RECT 715.500 389.400 717.300 395.250 ;
        RECT 719.700 392.400 721.500 395.250 ;
        RECT 722.700 392.400 724.500 395.250 ;
        RECT 725.700 392.400 727.500 395.250 ;
        RECT 728.700 392.400 730.500 395.250 ;
        RECT 719.700 391.050 721.050 392.400 ;
        RECT 722.700 391.050 724.050 392.400 ;
        RECT 725.700 391.050 727.050 392.400 ;
        RECT 733.200 391.500 735.000 395.250 ;
        RECT 736.200 392.400 738.000 395.250 ;
        RECT 739.200 391.500 741.000 395.250 ;
        RECT 692.250 386.250 696.000 387.300 ;
        RECT 685.950 384.450 688.050 385.050 ;
        RECT 691.950 384.450 694.050 385.050 ;
        RECT 685.950 383.550 694.050 384.450 ;
        RECT 685.950 382.950 688.050 383.550 ;
        RECT 691.950 382.950 694.050 383.550 ;
        RECT 694.950 382.950 696.150 386.250 ;
        RECT 698.100 384.150 699.900 385.950 ;
        RECT 704.700 385.800 705.900 389.400 ;
        RECT 715.800 388.500 717.300 389.400 ;
        RECT 708.900 387.300 717.300 388.500 ;
        RECT 718.950 388.950 721.050 391.050 ;
        RECT 721.950 388.950 724.050 391.050 ;
        RECT 724.950 388.950 727.050 391.050 ;
        RECT 730.500 390.750 732.300 391.200 ;
        RECT 728.250 389.400 732.300 390.750 ;
        RECT 733.200 389.700 736.050 391.500 ;
        RECT 733.950 389.400 736.050 389.700 ;
        RECT 738.150 389.700 741.000 391.500 ;
        RECT 742.950 391.500 744.750 395.250 ;
        RECT 745.950 391.500 747.750 395.250 ;
        RECT 748.950 391.500 750.750 395.250 ;
        RECT 738.150 389.400 740.250 389.700 ;
        RECT 742.950 389.400 745.050 391.500 ;
        RECT 745.950 389.400 748.050 391.500 ;
        RECT 748.950 389.400 751.050 391.500 ;
        RECT 753.600 390.600 755.400 395.250 ;
        RECT 753.600 389.400 757.800 390.600 ;
        RECT 759.150 389.400 760.950 395.250 ;
        RECT 764.550 389.400 766.350 395.250 ;
        RECT 708.900 386.700 710.700 387.300 ;
        RECT 718.950 385.800 720.000 388.950 ;
        RECT 728.250 388.050 729.150 389.400 ;
        RECT 724.050 387.900 729.150 388.050 ;
        RECT 704.700 384.900 720.000 385.800 ;
        RECT 721.500 387.150 729.150 387.900 ;
        RECT 721.500 386.700 725.850 387.150 ;
        RECT 737.100 386.700 744.000 388.500 ;
        RECT 744.900 386.700 751.650 388.500 ;
        RECT 682.950 380.850 685.050 382.950 ;
        RECT 694.950 380.850 697.050 382.950 ;
        RECT 697.950 382.050 700.050 384.150 ;
        RECT 700.950 380.850 703.050 382.950 ;
        RECT 683.100 379.050 684.900 380.850 ;
        RECT 678.750 377.400 681.000 378.300 ;
        RECT 691.950 377.850 694.050 379.950 ;
        RECT 678.750 376.500 684.450 377.400 ;
        RECT 652.650 363.750 654.450 369.000 ;
        RECT 655.650 363.750 657.450 369.600 ;
        RECT 658.650 363.750 660.450 369.600 ;
        RECT 667.650 363.750 669.450 369.600 ;
        RECT 670.650 363.750 672.450 369.600 ;
        RECT 676.350 363.750 678.150 375.600 ;
        RECT 679.350 363.750 681.150 375.600 ;
        RECT 683.250 369.600 684.450 376.500 ;
        RECT 692.250 376.050 694.050 377.850 ;
        RECT 695.850 375.600 697.050 380.850 ;
        RECT 701.100 379.050 702.900 380.850 ;
        RECT 682.650 363.750 684.450 369.600 ;
        RECT 692.400 363.750 694.200 369.600 ;
        RECT 695.700 363.750 697.500 375.600 ;
        RECT 699.900 363.750 701.700 375.600 ;
        RECT 704.700 371.400 705.900 384.900 ;
        RECT 707.100 382.950 718.950 384.000 ;
        RECT 721.500 383.250 722.550 386.700 ;
        RECT 724.050 386.250 725.850 386.700 ;
        RECT 730.950 385.650 733.050 385.950 ;
        RECT 742.950 385.800 744.000 386.700 ;
        RECT 756.300 385.800 757.800 389.400 ;
        RECT 729.150 383.850 733.050 385.650 ;
        RECT 734.400 384.450 742.050 385.800 ;
        RECT 742.950 384.750 752.850 385.800 ;
        RECT 707.100 381.150 708.900 382.950 ;
        RECT 706.950 379.050 709.050 381.150 ;
        RECT 717.750 380.550 718.950 382.950 ;
        RECT 720.750 381.450 722.550 383.250 ;
        RECT 734.400 382.950 735.450 384.450 ;
        RECT 741.150 383.700 742.050 384.450 ;
        RECT 723.450 382.050 735.450 382.950 ;
        RECT 723.450 380.550 724.500 382.050 ;
        RECT 736.350 381.750 740.250 383.550 ;
        RECT 741.150 382.650 750.750 383.700 ;
        RECT 738.150 381.450 740.250 381.750 ;
        RECT 712.950 379.650 715.050 379.950 ;
        RECT 717.750 379.650 724.500 380.550 ;
        RECT 725.400 380.550 727.200 381.150 ;
        RECT 733.950 380.550 736.050 380.850 ;
        RECT 725.400 379.950 736.050 380.550 ;
        RECT 746.700 379.950 748.500 381.750 ;
        RECT 712.950 378.450 716.850 379.650 ;
        RECT 725.400 379.350 748.500 379.950 ;
        RECT 733.950 378.750 748.500 379.350 ;
        RECT 749.850 381.000 750.750 382.650 ;
        RECT 751.800 382.950 752.850 384.750 ;
        RECT 756.300 384.000 764.100 385.800 ;
        RECT 751.800 381.900 760.050 382.950 ;
        RECT 749.850 379.200 756.900 381.000 ;
        RECT 712.950 377.850 726.900 378.450 ;
        RECT 757.950 377.850 760.050 381.900 ;
        RECT 713.250 377.550 753.000 377.850 ;
        RECT 724.950 376.650 753.000 377.550 ;
        RECT 762.450 376.650 764.250 377.250 ;
        RECT 712.500 376.050 714.300 376.650 ;
        RECT 721.950 376.050 724.050 376.350 ;
        RECT 712.500 374.850 724.050 376.050 ;
        RECT 721.950 374.250 724.050 374.850 ;
        RECT 724.950 374.400 745.050 375.750 ;
        RECT 709.200 373.350 711.000 374.100 ;
        RECT 724.950 373.350 726.900 374.400 ;
        RECT 742.950 373.650 745.050 374.400 ;
        RECT 748.950 374.550 751.050 375.750 ;
        RECT 751.950 375.450 764.250 376.650 ;
        RECT 765.150 374.550 766.350 389.400 ;
        RECT 748.950 373.650 766.350 374.550 ;
        RECT 768.450 392.400 770.250 395.250 ;
        RECT 771.450 392.400 773.250 395.250 ;
        RECT 768.450 384.150 769.950 392.400 ;
        RECT 782.550 390.300 784.350 395.250 ;
        RECT 785.550 391.200 787.350 395.250 ;
        RECT 788.550 390.300 790.350 395.250 ;
        RECT 782.550 388.950 790.350 390.300 ;
        RECT 791.550 389.400 793.350 395.250 ;
        RECT 791.550 387.300 792.750 389.400 ;
        RECT 789.000 386.250 792.750 387.300 ;
        RECT 803.100 387.000 804.900 395.250 ;
        RECT 785.100 384.150 786.900 385.950 ;
        RECT 768.450 382.050 772.050 384.150 ;
        RECT 709.200 372.300 726.900 373.350 ;
        RECT 704.700 370.500 708.750 371.400 ;
        RECT 707.700 369.600 708.750 370.500 ;
        RECT 704.700 363.750 706.500 369.600 ;
        RECT 707.700 363.750 709.500 369.600 ;
        RECT 710.700 363.750 712.500 369.600 ;
        RECT 713.700 363.750 715.500 372.300 ;
        RECT 733.950 372.150 736.050 372.600 ;
        RECT 733.650 370.500 736.050 372.150 ;
        RECT 738.000 370.800 741.900 372.600 ;
        RECT 738.000 370.500 741.000 370.800 ;
        RECT 718.950 367.950 721.050 370.050 ;
        RECT 721.950 367.950 724.050 370.050 ;
        RECT 724.950 369.600 727.050 370.050 ;
        RECT 733.650 369.600 735.000 370.500 ;
        RECT 724.950 367.950 727.500 369.600 ;
        RECT 716.700 363.750 718.500 367.050 ;
        RECT 719.850 366.600 721.050 367.950 ;
        RECT 723.150 366.600 724.050 367.950 ;
        RECT 726.300 366.600 727.500 367.950 ;
        RECT 719.850 363.750 722.250 366.600 ;
        RECT 723.150 363.750 725.250 366.600 ;
        RECT 726.300 363.750 728.250 366.600 ;
        RECT 729.450 363.750 731.250 369.600 ;
        RECT 733.200 363.750 735.000 369.600 ;
        RECT 736.200 363.750 738.000 369.600 ;
        RECT 739.200 363.750 741.000 370.500 ;
        RECT 743.100 366.600 744.450 373.650 ;
        RECT 752.850 372.150 754.650 372.300 ;
        RECT 745.950 370.950 754.650 372.150 ;
        RECT 759.600 371.700 761.400 372.300 ;
        RECT 745.950 370.050 748.050 370.950 ;
        RECT 752.850 370.500 754.650 370.950 ;
        RECT 755.700 370.500 761.400 371.700 ;
        RECT 742.950 363.750 744.750 366.600 ;
        RECT 745.950 363.750 747.750 370.050 ;
        RECT 749.100 367.800 751.200 369.900 ;
        RECT 749.100 366.600 750.600 367.800 ;
        RECT 748.950 363.750 750.750 366.600 ;
        RECT 752.700 363.750 754.500 369.600 ;
        RECT 755.700 363.750 757.500 370.500 ;
        RECT 762.300 369.600 763.500 373.650 ;
        RECT 768.450 369.600 769.950 382.050 ;
        RECT 781.950 380.850 784.050 382.950 ;
        RECT 784.950 382.050 787.050 384.150 ;
        RECT 788.850 382.950 790.050 386.250 ;
        RECT 800.400 385.350 804.900 387.000 ;
        RECT 808.500 386.400 810.300 395.250 ;
        RECT 815.550 392.400 817.350 395.250 ;
        RECT 818.550 392.400 820.350 395.250 ;
        RECT 790.950 384.450 793.050 385.050 ;
        RECT 796.950 384.450 799.050 385.050 ;
        RECT 790.950 383.550 799.050 384.450 ;
        RECT 790.950 382.950 793.050 383.550 ;
        RECT 796.950 382.950 799.050 383.550 ;
        RECT 787.950 380.850 790.050 382.950 ;
        RECT 800.400 381.150 801.600 385.350 ;
        RECT 814.950 383.850 817.050 385.950 ;
        RECT 818.400 384.150 819.600 392.400 ;
        RECT 827.850 389.400 829.650 395.250 ;
        RECT 832.350 388.200 834.150 395.250 ;
        RECT 847.650 389.400 849.450 395.250 ;
        RECT 850.650 392.400 852.450 395.250 ;
        RECT 853.650 392.400 855.450 395.250 ;
        RECT 856.650 392.400 858.450 395.250 ;
        RECT 830.550 387.300 834.150 388.200 ;
        RECT 815.100 382.050 816.900 383.850 ;
        RECT 817.950 382.050 820.050 384.150 ;
        RECT 782.100 379.050 783.900 380.850 ;
        RECT 787.950 375.600 789.150 380.850 ;
        RECT 790.950 377.850 793.050 379.950 ;
        RECT 799.950 379.050 802.050 381.150 ;
        RECT 790.950 376.050 792.750 377.850 ;
        RECT 758.700 363.750 760.500 369.600 ;
        RECT 761.700 363.750 763.500 369.600 ;
        RECT 764.700 363.750 766.500 369.600 ;
        RECT 768.450 363.750 770.250 369.600 ;
        RECT 771.450 363.750 773.250 369.600 ;
        RECT 783.300 363.750 785.100 375.600 ;
        RECT 787.500 363.750 789.300 375.600 ;
        RECT 800.250 370.800 801.300 379.050 ;
        RECT 802.950 377.850 805.050 379.950 ;
        RECT 808.950 377.850 811.050 379.950 ;
        RECT 802.950 376.050 804.750 377.850 ;
        RECT 805.950 374.850 808.050 376.950 ;
        RECT 809.100 376.050 810.900 377.850 ;
        RECT 806.100 373.050 807.900 374.850 ;
        RECT 800.250 369.900 807.300 370.800 ;
        RECT 800.250 369.600 801.450 369.900 ;
        RECT 790.800 363.750 792.600 369.600 ;
        RECT 799.650 363.750 801.450 369.600 ;
        RECT 805.650 369.600 807.300 369.900 ;
        RECT 818.400 369.600 819.600 382.050 ;
        RECT 827.100 381.150 828.900 382.950 ;
        RECT 826.950 379.050 829.050 381.150 ;
        RECT 830.550 379.950 831.750 387.300 ;
        RECT 847.950 384.150 849.000 389.400 ;
        RECT 853.650 388.200 854.550 392.400 ;
        RECT 851.250 387.300 854.550 388.200 ;
        RECT 851.250 386.400 853.050 387.300 ;
        RECT 833.100 381.150 834.900 382.950 ;
        RECT 847.950 382.050 850.050 384.150 ;
        RECT 829.950 377.850 832.050 379.950 ;
        RECT 832.950 379.050 835.050 381.150 ;
        RECT 830.550 369.600 831.750 377.850 ;
        RECT 848.550 375.450 849.900 382.050 ;
        RECT 851.400 378.150 852.300 386.400 ;
        RECT 856.950 383.850 859.050 385.950 ;
        RECT 853.950 380.850 856.050 382.950 ;
        RECT 857.100 382.050 858.900 383.850 ;
        RECT 854.100 379.050 855.900 380.850 ;
        RECT 851.250 378.000 853.050 378.150 ;
        RECT 851.250 376.800 858.450 378.000 ;
        RECT 851.250 376.350 853.050 376.800 ;
        RECT 857.250 375.600 858.450 376.800 ;
        RECT 848.550 374.100 850.950 375.450 ;
        RECT 802.650 363.750 804.450 369.000 ;
        RECT 805.650 363.750 807.450 369.600 ;
        RECT 808.650 363.750 810.450 369.600 ;
        RECT 815.550 363.750 817.350 369.600 ;
        RECT 818.550 363.750 820.350 369.600 ;
        RECT 827.550 363.750 829.350 369.600 ;
        RECT 830.550 363.750 832.350 369.600 ;
        RECT 833.550 363.750 835.350 369.600 ;
        RECT 849.150 363.750 850.950 374.100 ;
        RECT 852.150 363.750 853.950 375.450 ;
        RECT 856.650 363.750 858.450 375.600 ;
        RECT 9.150 348.900 10.950 359.250 ;
        RECT 8.550 347.550 10.950 348.900 ;
        RECT 12.150 347.550 13.950 359.250 ;
        RECT 8.550 340.950 9.900 347.550 ;
        RECT 16.650 347.400 18.450 359.250 ;
        RECT 25.650 353.400 27.450 359.250 ;
        RECT 28.650 353.400 30.450 359.250 ;
        RECT 31.650 353.400 33.450 359.250 ;
        RECT 11.250 346.200 13.050 346.650 ;
        RECT 17.250 346.200 18.450 347.400 ;
        RECT 11.250 345.000 18.450 346.200 ;
        RECT 29.250 345.150 30.450 353.400 ;
        RECT 42.450 347.400 44.250 359.250 ;
        RECT 46.650 347.400 48.450 359.250 ;
        RECT 53.550 348.300 55.350 359.250 ;
        RECT 56.550 349.200 58.350 359.250 ;
        RECT 59.550 348.300 61.350 359.250 ;
        RECT 53.550 347.400 61.350 348.300 ;
        RECT 62.550 347.400 64.350 359.250 ;
        RECT 78.450 347.400 80.250 359.250 ;
        RECT 82.650 347.400 84.450 359.250 ;
        RECT 86.550 347.400 88.350 359.250 ;
        RECT 90.750 347.400 92.550 359.250 ;
        RECT 98.550 353.400 100.350 359.250 ;
        RECT 101.550 353.400 103.350 359.250 ;
        RECT 113.550 353.400 115.350 359.250 ;
        RECT 116.550 353.400 118.350 359.250 ;
        RECT 119.550 354.000 121.350 359.250 ;
        RECT 42.450 346.350 45.000 347.400 ;
        RECT 11.250 344.850 13.050 345.000 ;
        RECT 7.950 338.850 10.050 340.950 ;
        RECT 7.950 333.600 9.000 338.850 ;
        RECT 11.400 336.600 12.300 344.850 ;
        RECT 14.100 342.150 15.900 343.950 ;
        RECT 13.950 340.050 16.050 342.150 ;
        RECT 25.950 341.850 28.050 343.950 ;
        RECT 28.950 343.050 31.050 345.150 ;
        RECT 17.100 339.150 18.900 340.950 ;
        RECT 26.100 340.050 27.900 341.850 ;
        RECT 16.950 337.050 19.050 339.150 ;
        RECT 11.250 335.700 13.050 336.600 ;
        RECT 29.250 335.700 30.450 343.050 ;
        RECT 31.950 341.850 34.050 343.950 ;
        RECT 41.100 342.150 42.900 343.950 ;
        RECT 32.100 340.050 33.900 341.850 ;
        RECT 40.950 340.050 43.050 342.150 ;
        RECT 11.250 334.800 14.550 335.700 ;
        RECT 7.650 327.750 9.450 333.600 ;
        RECT 13.650 330.600 14.550 334.800 ;
        RECT 26.850 334.800 30.450 335.700 ;
        RECT 43.950 339.150 45.000 346.350 ;
        RECT 47.100 342.150 48.900 343.950 ;
        RECT 62.700 342.150 63.900 347.400 ;
        RECT 78.450 346.350 81.000 347.400 ;
        RECT 77.100 342.150 78.900 343.950 ;
        RECT 46.950 340.050 49.050 342.150 ;
        RECT 43.950 337.050 46.050 339.150 ;
        RECT 52.950 338.850 55.050 340.950 ;
        RECT 56.100 339.150 57.900 340.950 ;
        RECT 53.100 337.050 54.900 338.850 ;
        RECT 55.950 337.050 58.050 339.150 ;
        RECT 58.950 338.850 61.050 340.950 ;
        RECT 61.950 340.050 64.050 342.150 ;
        RECT 76.950 340.050 79.050 342.150 ;
        RECT 59.100 337.050 60.900 338.850 ;
        RECT 10.650 327.750 12.450 330.600 ;
        RECT 13.650 327.750 15.450 330.600 ;
        RECT 16.650 327.750 18.450 330.600 ;
        RECT 26.850 327.750 28.650 334.800 ;
        RECT 31.350 327.750 33.150 333.600 ;
        RECT 43.950 330.600 45.000 337.050 ;
        RECT 62.700 333.600 63.900 340.050 ;
        RECT 40.650 327.750 42.450 330.600 ;
        RECT 43.650 327.750 45.450 330.600 ;
        RECT 46.650 327.750 48.450 330.600 ;
        RECT 54.000 327.750 55.800 333.600 ;
        RECT 58.200 331.950 63.900 333.600 ;
        RECT 79.950 339.150 81.000 346.350 ;
        RECT 90.000 346.350 92.550 347.400 ;
        RECT 83.100 342.150 84.900 343.950 ;
        RECT 86.100 342.150 87.900 343.950 ;
        RECT 82.950 340.050 85.050 342.150 ;
        RECT 85.950 340.050 88.050 342.150 ;
        RECT 90.000 339.150 91.050 346.350 ;
        RECT 92.100 342.150 93.900 343.950 ;
        RECT 91.950 340.050 94.050 342.150 ;
        RECT 101.400 340.950 102.600 353.400 ;
        RECT 116.700 353.100 118.350 353.400 ;
        RECT 122.550 353.400 124.350 359.250 ;
        RECT 133.650 353.400 135.450 359.250 ;
        RECT 136.650 353.400 138.450 359.250 ;
        RECT 139.650 353.400 141.450 359.250 ;
        RECT 148.650 353.400 150.450 359.250 ;
        RECT 151.650 353.400 153.450 359.250 ;
        RECT 154.650 353.400 156.450 359.250 ;
        RECT 161.550 353.400 163.350 359.250 ;
        RECT 164.550 353.400 166.350 359.250 ;
        RECT 167.550 353.400 169.350 359.250 ;
        RECT 122.550 353.100 123.750 353.400 ;
        RECT 116.700 352.200 123.750 353.100 ;
        RECT 116.100 348.150 117.900 349.950 ;
        RECT 113.100 345.150 114.900 346.950 ;
        RECT 115.950 346.050 118.050 348.150 ;
        RECT 119.250 345.150 121.050 346.950 ;
        RECT 112.950 343.050 115.050 345.150 ;
        RECT 118.950 343.050 121.050 345.150 ;
        RECT 122.700 343.950 123.750 352.200 ;
        RECT 124.950 348.450 127.050 349.050 ;
        RECT 133.950 348.450 136.050 349.050 ;
        RECT 124.950 347.550 136.050 348.450 ;
        RECT 124.950 346.950 127.050 347.550 ;
        RECT 133.950 346.950 136.050 347.550 ;
        RECT 137.250 345.150 138.450 353.400 ;
        RECT 139.950 348.450 142.050 349.050 ;
        RECT 145.950 348.450 148.050 349.050 ;
        RECT 139.950 347.550 148.050 348.450 ;
        RECT 139.950 346.950 142.050 347.550 ;
        RECT 145.950 346.950 148.050 347.550 ;
        RECT 152.250 345.150 153.450 353.400 ;
        RECT 164.550 345.150 165.750 353.400 ;
        RECT 175.650 347.400 177.450 359.250 ;
        RECT 178.650 348.300 180.450 359.250 ;
        RECT 181.650 349.200 183.450 359.250 ;
        RECT 184.650 348.300 186.450 359.250 ;
        RECT 178.650 347.400 186.450 348.300 ;
        RECT 195.300 347.400 197.100 359.250 ;
        RECT 199.500 347.400 201.300 359.250 ;
        RECT 202.800 353.400 204.600 359.250 ;
        RECT 213.450 347.400 215.250 359.250 ;
        RECT 217.650 347.400 219.450 359.250 ;
        RECT 228.300 347.400 230.100 359.250 ;
        RECT 232.500 347.400 234.300 359.250 ;
        RECT 235.800 353.400 237.600 359.250 ;
        RECT 245.550 348.300 247.350 359.250 ;
        RECT 248.550 349.200 250.350 359.250 ;
        RECT 251.550 348.300 253.350 359.250 ;
        RECT 245.550 347.400 253.350 348.300 ;
        RECT 254.550 347.400 256.350 359.250 ;
        RECT 268.350 347.400 270.150 359.250 ;
        RECT 271.350 347.400 273.150 359.250 ;
        RECT 274.650 353.400 276.450 359.250 ;
        RECT 280.650 353.400 282.450 359.250 ;
        RECT 283.650 353.400 285.450 359.250 ;
        RECT 286.650 353.400 288.450 359.250 ;
        RECT 121.950 341.850 124.050 343.950 ;
        RECT 133.950 341.850 136.050 343.950 ;
        RECT 136.950 343.050 139.050 345.150 ;
        RECT 98.100 339.150 99.900 340.950 ;
        RECT 79.950 337.050 82.050 339.150 ;
        RECT 88.950 337.050 91.050 339.150 ;
        RECT 97.950 337.050 100.050 339.150 ;
        RECT 100.950 338.850 103.050 340.950 ;
        RECT 58.200 327.750 60.000 331.950 ;
        RECT 79.950 330.600 81.000 337.050 ;
        RECT 90.000 330.600 91.050 337.050 ;
        RECT 101.400 330.600 102.600 338.850 ;
        RECT 122.400 337.650 123.600 341.850 ;
        RECT 134.100 340.050 135.900 341.850 ;
        RECT 61.500 327.750 63.300 330.600 ;
        RECT 76.650 327.750 78.450 330.600 ;
        RECT 79.650 327.750 81.450 330.600 ;
        RECT 82.650 327.750 84.450 330.600 ;
        RECT 86.550 327.750 88.350 330.600 ;
        RECT 89.550 327.750 91.350 330.600 ;
        RECT 92.550 327.750 94.350 330.600 ;
        RECT 98.550 327.750 100.350 330.600 ;
        RECT 101.550 327.750 103.350 330.600 ;
        RECT 113.700 327.750 115.500 336.600 ;
        RECT 119.100 336.000 123.600 337.650 ;
        RECT 119.100 327.750 120.900 336.000 ;
        RECT 137.250 335.700 138.450 343.050 ;
        RECT 139.950 341.850 142.050 343.950 ;
        RECT 148.950 341.850 151.050 343.950 ;
        RECT 151.950 343.050 154.050 345.150 ;
        RECT 140.100 340.050 141.900 341.850 ;
        RECT 149.100 340.050 150.900 341.850 ;
        RECT 152.250 335.700 153.450 343.050 ;
        RECT 154.950 341.850 157.050 343.950 ;
        RECT 160.950 341.850 163.050 343.950 ;
        RECT 163.950 343.050 166.050 345.150 ;
        RECT 155.100 340.050 156.900 341.850 ;
        RECT 161.100 340.050 162.900 341.850 ;
        RECT 134.850 334.800 138.450 335.700 ;
        RECT 149.850 334.800 153.450 335.700 ;
        RECT 164.550 335.700 165.750 343.050 ;
        RECT 166.950 341.850 169.050 343.950 ;
        RECT 176.100 342.150 177.300 347.400 ;
        RECT 178.950 345.450 181.050 346.050 ;
        RECT 178.950 344.550 192.450 345.450 ;
        RECT 178.950 343.950 181.050 344.550 ;
        RECT 167.100 340.050 168.900 341.850 ;
        RECT 175.950 340.050 178.050 342.150 ;
        RECT 164.550 334.800 168.150 335.700 ;
        RECT 134.850 327.750 136.650 334.800 ;
        RECT 139.350 327.750 141.150 333.600 ;
        RECT 149.850 327.750 151.650 334.800 ;
        RECT 154.350 327.750 156.150 333.600 ;
        RECT 161.850 327.750 163.650 333.600 ;
        RECT 166.350 327.750 168.150 334.800 ;
        RECT 176.100 333.600 177.300 340.050 ;
        RECT 178.950 338.850 181.050 340.950 ;
        RECT 182.100 339.150 183.900 340.950 ;
        RECT 179.100 337.050 180.900 338.850 ;
        RECT 181.950 337.050 184.050 339.150 ;
        RECT 184.950 338.850 187.050 340.950 ;
        RECT 185.100 337.050 186.900 338.850 ;
        RECT 191.550 336.450 192.450 344.550 ;
        RECT 194.100 342.150 195.900 343.950 ;
        RECT 199.950 342.150 201.150 347.400 ;
        RECT 202.950 345.150 204.750 346.950 ;
        RECT 213.450 346.350 216.000 347.400 ;
        RECT 202.950 343.050 205.050 345.150 ;
        RECT 212.100 342.150 213.900 343.950 ;
        RECT 193.950 340.050 196.050 342.150 ;
        RECT 196.950 338.850 199.050 340.950 ;
        RECT 199.950 340.050 202.050 342.150 ;
        RECT 211.950 340.050 214.050 342.150 ;
        RECT 197.100 337.050 198.900 338.850 ;
        RECT 193.950 336.450 196.050 337.050 ;
        RECT 200.850 336.750 202.050 340.050 ;
        RECT 214.950 339.150 216.000 346.350 ;
        RECT 218.100 342.150 219.900 343.950 ;
        RECT 227.100 342.150 228.900 343.950 ;
        RECT 232.950 342.150 234.150 347.400 ;
        RECT 235.950 345.150 237.750 346.950 ;
        RECT 235.950 343.050 238.050 345.150 ;
        RECT 254.700 342.150 255.900 347.400 ;
        RECT 268.650 342.150 269.850 347.400 ;
        RECT 275.250 346.500 276.450 353.400 ;
        RECT 270.750 345.600 276.450 346.500 ;
        RECT 270.750 344.700 273.000 345.600 ;
        RECT 284.250 345.150 285.450 353.400 ;
        RECT 295.050 347.400 296.850 359.250 ;
        RECT 298.050 347.400 299.850 359.250 ;
        RECT 301.650 353.400 303.450 359.250 ;
        RECT 304.650 353.400 306.450 359.250 ;
        RECT 217.950 340.050 220.050 342.150 ;
        RECT 226.950 340.050 229.050 342.150 ;
        RECT 214.950 337.050 217.050 339.150 ;
        RECT 229.950 338.850 232.050 340.950 ;
        RECT 232.950 340.050 235.050 342.150 ;
        RECT 230.100 337.050 231.900 338.850 ;
        RECT 191.550 335.550 196.050 336.450 ;
        RECT 201.000 335.700 204.750 336.750 ;
        RECT 193.950 334.950 196.050 335.550 ;
        RECT 176.100 331.950 181.800 333.600 ;
        RECT 176.700 327.750 178.500 330.600 ;
        RECT 180.000 327.750 181.800 331.950 ;
        RECT 184.200 327.750 186.000 333.600 ;
        RECT 194.550 332.700 202.350 334.050 ;
        RECT 194.550 327.750 196.350 332.700 ;
        RECT 197.550 327.750 199.350 331.800 ;
        RECT 200.550 327.750 202.350 332.700 ;
        RECT 203.550 333.600 204.750 335.700 ;
        RECT 203.550 327.750 205.350 333.600 ;
        RECT 214.950 330.600 216.000 337.050 ;
        RECT 233.850 336.750 235.050 340.050 ;
        RECT 244.950 338.850 247.050 340.950 ;
        RECT 248.100 339.150 249.900 340.950 ;
        RECT 245.100 337.050 246.900 338.850 ;
        RECT 247.950 337.050 250.050 339.150 ;
        RECT 250.950 338.850 253.050 340.950 ;
        RECT 253.950 340.050 256.050 342.150 ;
        RECT 268.650 340.050 271.050 342.150 ;
        RECT 251.100 337.050 252.900 338.850 ;
        RECT 234.000 335.700 237.750 336.750 ;
        RECT 227.550 332.700 235.350 334.050 ;
        RECT 211.650 327.750 213.450 330.600 ;
        RECT 214.650 327.750 216.450 330.600 ;
        RECT 217.650 327.750 219.450 330.600 ;
        RECT 227.550 327.750 229.350 332.700 ;
        RECT 230.550 327.750 232.350 331.800 ;
        RECT 233.550 327.750 235.350 332.700 ;
        RECT 236.550 333.600 237.750 335.700 ;
        RECT 254.700 333.600 255.900 340.050 ;
        RECT 268.650 333.600 269.850 340.050 ;
        RECT 271.950 336.300 273.000 344.700 ;
        RECT 275.100 342.150 276.900 343.950 ;
        RECT 274.950 340.050 277.050 342.150 ;
        RECT 280.950 341.850 283.050 343.950 ;
        RECT 283.950 343.050 286.050 345.150 ;
        RECT 281.100 340.050 282.900 341.850 ;
        RECT 270.750 335.400 273.000 336.300 ;
        RECT 284.250 335.700 285.450 343.050 ;
        RECT 286.950 341.850 289.050 343.950 ;
        RECT 295.650 342.150 296.850 347.400 ;
        RECT 287.100 340.050 288.900 341.850 ;
        RECT 295.650 340.050 298.050 342.150 ;
        RECT 298.950 341.850 301.050 343.950 ;
        RECT 299.100 340.050 300.900 341.850 ;
        RECT 270.750 334.500 275.850 335.400 ;
        RECT 236.550 327.750 238.350 333.600 ;
        RECT 246.000 327.750 247.800 333.600 ;
        RECT 250.200 331.950 255.900 333.600 ;
        RECT 250.200 327.750 252.000 331.950 ;
        RECT 253.500 327.750 255.300 330.600 ;
        RECT 268.350 327.750 270.150 333.600 ;
        RECT 271.350 327.750 273.150 333.600 ;
        RECT 274.650 330.600 275.850 334.500 ;
        RECT 281.850 334.800 285.450 335.700 ;
        RECT 274.650 327.750 276.450 330.600 ;
        RECT 281.850 327.750 283.650 334.800 ;
        RECT 295.650 333.600 296.850 340.050 ;
        RECT 302.100 336.300 303.300 353.400 ;
        RECT 312.300 347.400 314.100 359.250 ;
        RECT 316.500 347.400 318.300 359.250 ;
        RECT 319.800 353.400 321.600 359.250 ;
        RECT 331.650 347.400 333.450 359.250 ;
        RECT 334.650 347.400 336.450 359.250 ;
        RECT 343.650 347.400 345.450 359.250 ;
        RECT 346.650 348.300 348.450 359.250 ;
        RECT 349.650 349.200 351.450 359.250 ;
        RECT 352.650 348.300 354.450 359.250 ;
        RECT 346.650 347.400 354.450 348.300 ;
        RECT 360.300 347.400 362.100 359.250 ;
        RECT 364.500 347.400 366.300 359.250 ;
        RECT 367.800 353.400 369.600 359.250 ;
        RECT 379.050 347.400 380.850 359.250 ;
        RECT 382.050 347.400 383.850 359.250 ;
        RECT 385.650 353.400 387.450 359.250 ;
        RECT 388.650 353.400 390.450 359.250 ;
        RECT 305.100 342.150 306.900 343.950 ;
        RECT 311.100 342.150 312.900 343.950 ;
        RECT 316.950 342.150 318.150 347.400 ;
        RECT 319.950 345.150 321.750 346.950 ;
        RECT 319.950 343.050 322.050 345.150 ;
        RECT 332.400 342.150 333.600 347.400 ;
        RECT 344.100 342.150 345.300 347.400 ;
        RECT 359.100 342.150 360.900 343.950 ;
        RECT 364.950 342.150 366.150 347.400 ;
        RECT 367.950 345.150 369.750 346.950 ;
        RECT 367.950 343.050 370.050 345.150 ;
        RECT 379.650 342.150 380.850 347.400 ;
        RECT 304.950 340.050 307.050 342.150 ;
        RECT 310.950 340.050 313.050 342.150 ;
        RECT 313.950 338.850 316.050 340.950 ;
        RECT 316.950 340.050 319.050 342.150 ;
        RECT 331.950 340.050 334.050 342.150 ;
        RECT 314.100 337.050 315.900 338.850 ;
        RECT 317.850 336.750 319.050 340.050 ;
        RECT 298.950 335.100 306.450 336.300 ;
        RECT 318.000 335.700 321.750 336.750 ;
        RECT 298.950 334.500 300.750 335.100 ;
        RECT 286.350 327.750 288.150 333.600 ;
        RECT 295.650 332.100 298.950 333.600 ;
        RECT 297.150 327.750 298.950 332.100 ;
        RECT 300.150 327.750 301.950 333.600 ;
        RECT 304.650 327.750 306.450 335.100 ;
        RECT 311.550 332.700 319.350 334.050 ;
        RECT 311.550 327.750 313.350 332.700 ;
        RECT 314.550 327.750 316.350 331.800 ;
        RECT 317.550 327.750 319.350 332.700 ;
        RECT 320.550 333.600 321.750 335.700 ;
        RECT 332.400 333.600 333.600 340.050 ;
        RECT 334.950 338.850 337.050 340.950 ;
        RECT 343.950 340.050 346.050 342.150 ;
        RECT 335.100 337.050 336.900 338.850 ;
        RECT 344.100 333.600 345.300 340.050 ;
        RECT 346.950 338.850 349.050 340.950 ;
        RECT 350.100 339.150 351.900 340.950 ;
        RECT 347.100 337.050 348.900 338.850 ;
        RECT 349.950 337.050 352.050 339.150 ;
        RECT 352.950 338.850 355.050 340.950 ;
        RECT 358.950 340.050 361.050 342.150 ;
        RECT 361.950 338.850 364.050 340.950 ;
        RECT 364.950 340.050 367.050 342.150 ;
        RECT 353.100 337.050 354.900 338.850 ;
        RECT 362.100 337.050 363.900 338.850 ;
        RECT 365.850 336.750 367.050 340.050 ;
        RECT 379.650 340.050 382.050 342.150 ;
        RECT 382.950 341.850 385.050 343.950 ;
        RECT 383.100 340.050 384.900 341.850 ;
        RECT 366.000 335.700 369.750 336.750 ;
        RECT 320.550 327.750 322.350 333.600 ;
        RECT 331.650 327.750 333.450 333.600 ;
        RECT 334.650 327.750 336.450 333.600 ;
        RECT 344.100 331.950 349.800 333.600 ;
        RECT 344.700 327.750 346.500 330.600 ;
        RECT 348.000 327.750 349.800 331.950 ;
        RECT 352.200 327.750 354.000 333.600 ;
        RECT 359.550 332.700 367.350 334.050 ;
        RECT 359.550 327.750 361.350 332.700 ;
        RECT 362.550 327.750 364.350 331.800 ;
        RECT 365.550 327.750 367.350 332.700 ;
        RECT 368.550 333.600 369.750 335.700 ;
        RECT 379.650 333.600 380.850 340.050 ;
        RECT 386.100 336.300 387.300 353.400 ;
        RECT 399.450 347.400 401.250 359.250 ;
        RECT 403.650 347.400 405.450 359.250 ;
        RECT 410.550 347.400 412.350 359.250 ;
        RECT 414.750 347.400 416.550 359.250 ;
        RECT 425.550 347.400 427.350 359.250 ;
        RECT 429.750 347.400 431.550 359.250 ;
        RECT 399.450 346.350 402.000 347.400 ;
        RECT 389.100 342.150 390.900 343.950 ;
        RECT 398.100 342.150 399.900 343.950 ;
        RECT 388.950 340.050 391.050 342.150 ;
        RECT 397.950 340.050 400.050 342.150 ;
        RECT 400.950 339.150 402.000 346.350 ;
        RECT 414.000 346.350 416.550 347.400 ;
        RECT 429.000 346.350 431.550 347.400 ;
        RECT 444.450 347.400 446.250 359.250 ;
        RECT 448.650 347.400 450.450 359.250 ;
        RECT 455.550 347.400 457.350 359.250 ;
        RECT 459.750 347.400 461.550 359.250 ;
        RECT 472.650 347.400 474.450 359.250 ;
        RECT 475.650 347.400 477.450 359.250 ;
        RECT 485.550 348.600 487.350 359.250 ;
        RECT 488.550 349.500 490.350 359.250 ;
        RECT 491.550 358.500 499.350 359.250 ;
        RECT 491.550 348.600 493.350 358.500 ;
        RECT 485.550 347.700 493.350 348.600 ;
        RECT 494.550 347.400 496.350 357.600 ;
        RECT 497.550 347.400 499.350 358.500 ;
        RECT 505.650 353.400 507.450 359.250 ;
        RECT 508.650 353.400 510.450 359.250 ;
        RECT 444.450 346.350 447.000 347.400 ;
        RECT 404.100 342.150 405.900 343.950 ;
        RECT 410.100 342.150 411.900 343.950 ;
        RECT 403.950 340.050 406.050 342.150 ;
        RECT 409.950 340.050 412.050 342.150 ;
        RECT 414.000 339.150 415.050 346.350 ;
        RECT 416.100 342.150 417.900 343.950 ;
        RECT 425.100 342.150 426.900 343.950 ;
        RECT 415.950 340.050 418.050 342.150 ;
        RECT 424.950 340.050 427.050 342.150 ;
        RECT 429.000 339.150 430.050 346.350 ;
        RECT 431.100 342.150 432.900 343.950 ;
        RECT 443.100 342.150 444.900 343.950 ;
        RECT 430.950 340.050 433.050 342.150 ;
        RECT 442.950 340.050 445.050 342.150 ;
        RECT 400.950 337.050 403.050 339.150 ;
        RECT 412.950 337.050 415.050 339.150 ;
        RECT 427.950 337.050 430.050 339.150 ;
        RECT 382.950 335.100 390.450 336.300 ;
        RECT 382.950 334.500 384.750 335.100 ;
        RECT 368.550 327.750 370.350 333.600 ;
        RECT 379.650 332.100 382.950 333.600 ;
        RECT 381.150 327.750 382.950 332.100 ;
        RECT 384.150 327.750 385.950 333.600 ;
        RECT 388.650 327.750 390.450 335.100 ;
        RECT 400.950 330.600 402.000 337.050 ;
        RECT 414.000 330.600 415.050 337.050 ;
        RECT 429.000 330.600 430.050 337.050 ;
        RECT 445.950 339.150 447.000 346.350 ;
        RECT 459.000 346.350 461.550 347.400 ;
        RECT 451.950 343.950 454.050 346.050 ;
        RECT 449.100 342.150 450.900 343.950 ;
        RECT 448.950 340.050 451.050 342.150 ;
        RECT 445.950 337.050 448.050 339.150 ;
        RECT 445.950 330.600 447.000 337.050 ;
        RECT 448.950 336.450 451.050 337.050 ;
        RECT 452.550 336.450 453.450 343.950 ;
        RECT 455.100 342.150 456.900 343.950 ;
        RECT 454.950 340.050 457.050 342.150 ;
        RECT 459.000 339.150 460.050 346.350 ;
        RECT 461.100 342.150 462.900 343.950 ;
        RECT 473.400 342.150 474.600 347.400 ;
        RECT 494.400 346.500 496.200 347.400 ;
        RECT 492.150 345.600 496.200 346.500 ;
        RECT 485.250 342.150 487.050 343.950 ;
        RECT 492.150 342.150 493.050 345.600 ;
        RECT 497.100 342.150 498.900 343.950 ;
        RECT 460.950 340.050 463.050 342.150 ;
        RECT 472.950 340.050 475.050 342.150 ;
        RECT 457.950 337.050 460.050 339.150 ;
        RECT 448.950 335.550 453.450 336.450 ;
        RECT 448.950 334.950 451.050 335.550 ;
        RECT 459.000 330.600 460.050 337.050 ;
        RECT 473.400 333.600 474.600 340.050 ;
        RECT 475.950 338.850 478.050 340.950 ;
        RECT 484.950 340.050 487.050 342.150 ;
        RECT 487.950 338.850 490.050 340.950 ;
        RECT 476.100 337.050 477.900 338.850 ;
        RECT 488.250 337.050 490.050 338.850 ;
        RECT 490.950 340.050 493.050 342.150 ;
        RECT 490.950 333.600 492.000 340.050 ;
        RECT 493.950 338.850 496.050 340.950 ;
        RECT 496.950 340.050 499.050 342.150 ;
        RECT 506.400 340.950 507.600 353.400 ;
        RECT 522.450 347.400 524.250 359.250 ;
        RECT 526.650 347.400 528.450 359.250 ;
        RECT 530.550 353.400 532.350 359.250 ;
        RECT 522.450 346.350 525.000 347.400 ;
        RECT 521.100 342.150 522.900 343.950 ;
        RECT 505.950 338.850 508.050 340.950 ;
        RECT 509.100 339.150 510.900 340.950 ;
        RECT 520.950 340.050 523.050 342.150 ;
        RECT 523.950 339.150 525.000 346.350 ;
        RECT 530.550 346.500 531.750 353.400 ;
        RECT 533.850 347.400 535.650 359.250 ;
        RECT 536.850 347.400 538.650 359.250 ;
        RECT 542.550 353.400 544.350 359.250 ;
        RECT 530.550 345.600 536.250 346.500 ;
        RECT 534.000 344.700 536.250 345.600 ;
        RECT 527.100 342.150 528.900 343.950 ;
        RECT 530.100 342.150 531.900 343.950 ;
        RECT 526.950 340.050 529.050 342.150 ;
        RECT 529.950 340.050 532.050 342.150 ;
        RECT 493.950 337.050 495.750 338.850 ;
        RECT 397.650 327.750 399.450 330.600 ;
        RECT 400.650 327.750 402.450 330.600 ;
        RECT 403.650 327.750 405.450 330.600 ;
        RECT 410.550 327.750 412.350 330.600 ;
        RECT 413.550 327.750 415.350 330.600 ;
        RECT 416.550 327.750 418.350 330.600 ;
        RECT 425.550 327.750 427.350 330.600 ;
        RECT 428.550 327.750 430.350 330.600 ;
        RECT 431.550 327.750 433.350 330.600 ;
        RECT 442.650 327.750 444.450 330.600 ;
        RECT 445.650 327.750 447.450 330.600 ;
        RECT 448.650 327.750 450.450 330.600 ;
        RECT 455.550 327.750 457.350 330.600 ;
        RECT 458.550 327.750 460.350 330.600 ;
        RECT 461.550 327.750 463.350 330.600 ;
        RECT 472.650 327.750 474.450 333.600 ;
        RECT 475.650 327.750 477.450 333.600 ;
        RECT 486.000 327.750 487.800 333.600 ;
        RECT 490.200 327.750 492.000 333.600 ;
        RECT 494.400 327.750 496.200 333.600 ;
        RECT 506.400 330.600 507.600 338.850 ;
        RECT 508.950 337.050 511.050 339.150 ;
        RECT 523.950 337.050 526.050 339.150 ;
        RECT 523.950 330.600 525.000 337.050 ;
        RECT 534.000 336.300 535.050 344.700 ;
        RECT 537.150 342.150 538.350 347.400 ;
        RECT 542.550 346.500 543.750 353.400 ;
        RECT 545.850 347.400 547.650 359.250 ;
        RECT 548.850 347.400 550.650 359.250 ;
        RECT 562.650 353.400 564.450 359.250 ;
        RECT 565.650 353.400 567.450 359.250 ;
        RECT 568.650 353.400 570.450 359.250 ;
        RECT 581.400 353.400 583.200 359.250 ;
        RECT 542.550 345.600 548.250 346.500 ;
        RECT 546.000 344.700 548.250 345.600 ;
        RECT 542.100 342.150 543.900 343.950 ;
        RECT 535.950 340.050 538.350 342.150 ;
        RECT 541.950 340.050 544.050 342.150 ;
        RECT 534.000 335.400 536.250 336.300 ;
        RECT 531.150 334.500 536.250 335.400 ;
        RECT 531.150 330.600 532.350 334.500 ;
        RECT 537.150 333.600 538.350 340.050 ;
        RECT 546.000 336.300 547.050 344.700 ;
        RECT 549.150 342.150 550.350 347.400 ;
        RECT 566.250 345.150 567.450 353.400 ;
        RECT 584.700 347.400 586.500 359.250 ;
        RECT 588.900 347.400 590.700 359.250 ;
        RECT 598.650 347.400 600.450 359.250 ;
        RECT 601.650 347.400 603.450 359.250 ;
        RECT 606.750 353.400 608.550 359.250 ;
        RECT 609.750 353.400 611.550 359.250 ;
        RECT 613.500 353.400 615.300 359.250 ;
        RECT 616.500 353.400 618.300 359.250 ;
        RECT 619.500 353.400 621.300 359.250 ;
        RECT 581.250 345.150 583.050 346.950 ;
        RECT 547.950 340.050 550.350 342.150 ;
        RECT 562.950 341.850 565.050 343.950 ;
        RECT 565.950 343.050 568.050 345.150 ;
        RECT 563.100 340.050 564.900 341.850 ;
        RECT 546.000 335.400 548.250 336.300 ;
        RECT 543.150 334.500 548.250 335.400 ;
        RECT 505.650 327.750 507.450 330.600 ;
        RECT 508.650 327.750 510.450 330.600 ;
        RECT 520.650 327.750 522.450 330.600 ;
        RECT 523.650 327.750 525.450 330.600 ;
        RECT 526.650 327.750 528.450 330.600 ;
        RECT 530.550 327.750 532.350 330.600 ;
        RECT 533.850 327.750 535.650 333.600 ;
        RECT 536.850 327.750 538.650 333.600 ;
        RECT 543.150 330.600 544.350 334.500 ;
        RECT 549.150 333.600 550.350 340.050 ;
        RECT 566.250 335.700 567.450 343.050 ;
        RECT 568.950 341.850 571.050 343.950 ;
        RECT 580.950 343.050 583.050 345.150 ;
        RECT 584.850 342.150 586.050 347.400 ;
        RECT 590.100 342.150 591.900 343.950 ;
        RECT 599.400 342.150 600.600 347.400 ;
        RECT 569.100 340.050 570.900 341.850 ;
        RECT 583.950 340.050 586.050 342.150 ;
        RECT 583.950 336.750 585.150 340.050 ;
        RECT 586.950 338.850 589.050 340.950 ;
        RECT 589.950 340.050 592.050 342.150 ;
        RECT 598.950 340.050 601.050 342.150 ;
        RECT 610.050 340.950 611.550 353.400 ;
        RECT 616.500 349.350 617.700 353.400 ;
        RECT 622.500 352.500 624.300 359.250 ;
        RECT 625.500 353.400 627.300 359.250 ;
        RECT 629.250 356.400 631.050 359.250 ;
        RECT 629.400 355.200 630.900 356.400 ;
        RECT 628.800 353.100 630.900 355.200 ;
        RECT 632.250 352.950 634.050 359.250 ;
        RECT 635.250 356.400 637.050 359.250 ;
        RECT 618.600 351.300 624.300 352.500 ;
        RECT 625.350 352.050 627.150 352.500 ;
        RECT 631.950 352.050 634.050 352.950 ;
        RECT 618.600 350.700 620.400 351.300 ;
        RECT 625.350 350.850 634.050 352.050 ;
        RECT 625.350 350.700 627.150 350.850 ;
        RECT 635.550 349.350 636.900 356.400 ;
        RECT 639.000 352.500 640.800 359.250 ;
        RECT 642.000 353.400 643.800 359.250 ;
        RECT 645.000 353.400 646.800 359.250 ;
        RECT 648.750 353.400 650.550 359.250 ;
        RECT 651.750 356.400 653.700 359.250 ;
        RECT 654.750 356.400 656.850 359.250 ;
        RECT 657.750 356.400 660.150 359.250 ;
        RECT 652.500 355.050 653.700 356.400 ;
        RECT 655.950 355.050 656.850 356.400 ;
        RECT 658.950 355.050 660.150 356.400 ;
        RECT 661.500 355.950 663.300 359.250 ;
        RECT 652.500 353.400 655.050 355.050 ;
        RECT 645.000 352.500 646.350 353.400 ;
        RECT 652.950 352.950 655.050 353.400 ;
        RECT 655.950 352.950 658.050 355.050 ;
        RECT 658.950 352.950 661.050 355.050 ;
        RECT 639.000 352.200 642.000 352.500 ;
        RECT 638.100 350.400 642.000 352.200 ;
        RECT 643.950 350.850 646.350 352.500 ;
        RECT 643.950 350.400 646.050 350.850 ;
        RECT 664.500 350.700 666.300 359.250 ;
        RECT 667.500 353.400 669.300 359.250 ;
        RECT 670.500 353.400 672.300 359.250 ;
        RECT 673.500 353.400 675.300 359.250 ;
        RECT 677.700 353.400 679.500 359.250 ;
        RECT 680.700 353.400 682.500 359.250 ;
        RECT 683.700 353.400 685.500 359.250 ;
        RECT 671.250 352.500 672.300 353.400 ;
        RECT 680.700 352.500 681.750 353.400 ;
        RECT 671.250 351.600 675.300 352.500 ;
        RECT 653.100 349.650 670.800 350.700 ;
        RECT 587.100 337.050 588.900 338.850 ;
        RECT 563.850 334.800 567.450 335.700 ;
        RECT 581.250 335.700 585.000 336.750 ;
        RECT 542.550 327.750 544.350 330.600 ;
        RECT 545.850 327.750 547.650 333.600 ;
        RECT 548.850 327.750 550.650 333.600 ;
        RECT 563.850 327.750 565.650 334.800 ;
        RECT 581.250 333.600 582.450 335.700 ;
        RECT 568.350 327.750 570.150 333.600 ;
        RECT 580.650 327.750 582.450 333.600 ;
        RECT 583.650 332.700 591.450 334.050 ;
        RECT 599.400 333.600 600.600 340.050 ;
        RECT 601.950 338.850 604.050 340.950 ;
        RECT 607.950 338.850 611.550 340.950 ;
        RECT 602.100 337.050 603.900 338.850 ;
        RECT 583.650 327.750 585.450 332.700 ;
        RECT 586.650 327.750 588.450 331.800 ;
        RECT 589.650 327.750 591.450 332.700 ;
        RECT 598.650 327.750 600.450 333.600 ;
        RECT 601.650 327.750 603.450 333.600 ;
        RECT 610.050 330.600 611.550 338.850 ;
        RECT 606.750 327.750 608.550 330.600 ;
        RECT 609.750 327.750 611.550 330.600 ;
        RECT 613.650 348.450 631.050 349.350 ;
        RECT 613.650 333.600 614.850 348.450 ;
        RECT 615.750 346.350 628.050 347.550 ;
        RECT 628.950 347.250 631.050 348.450 ;
        RECT 634.950 348.600 637.050 349.350 ;
        RECT 653.100 348.600 655.050 349.650 ;
        RECT 669.000 348.900 670.800 349.650 ;
        RECT 634.950 347.250 655.050 348.600 ;
        RECT 655.950 348.150 658.050 348.750 ;
        RECT 655.950 346.950 667.500 348.150 ;
        RECT 655.950 346.650 658.050 346.950 ;
        RECT 665.700 346.350 667.500 346.950 ;
        RECT 615.750 345.750 617.550 346.350 ;
        RECT 627.000 345.450 655.050 346.350 ;
        RECT 627.000 345.150 666.750 345.450 ;
        RECT 619.950 341.100 622.050 345.150 ;
        RECT 653.100 344.550 667.050 345.150 ;
        RECT 623.100 342.000 630.150 343.800 ;
        RECT 619.950 340.050 628.200 341.100 ;
        RECT 615.900 337.200 623.700 339.000 ;
        RECT 627.150 338.250 628.200 340.050 ;
        RECT 629.250 340.350 630.150 342.000 ;
        RECT 631.500 343.650 646.050 344.250 ;
        RECT 631.500 343.050 654.600 343.650 ;
        RECT 663.150 343.350 667.050 344.550 ;
        RECT 631.500 341.250 633.300 343.050 ;
        RECT 643.950 342.450 654.600 343.050 ;
        RECT 643.950 342.150 646.050 342.450 ;
        RECT 652.800 341.850 654.600 342.450 ;
        RECT 655.500 342.450 662.250 343.350 ;
        RECT 664.950 343.050 667.050 343.350 ;
        RECT 639.750 341.250 641.850 341.550 ;
        RECT 629.250 339.300 638.850 340.350 ;
        RECT 639.750 339.450 643.650 341.250 ;
        RECT 655.500 340.950 656.550 342.450 ;
        RECT 644.550 340.050 656.550 340.950 ;
        RECT 637.950 338.550 638.850 339.300 ;
        RECT 644.550 338.550 645.600 340.050 ;
        RECT 657.450 339.750 659.250 341.550 ;
        RECT 661.050 340.050 662.250 342.450 ;
        RECT 670.950 341.850 673.050 343.950 ;
        RECT 671.100 340.050 672.900 341.850 ;
        RECT 627.150 337.200 637.050 338.250 ;
        RECT 637.950 337.200 645.600 338.550 ;
        RECT 646.950 337.350 650.850 339.150 ;
        RECT 622.200 333.600 623.700 337.200 ;
        RECT 636.000 336.300 637.050 337.200 ;
        RECT 646.950 337.050 649.050 337.350 ;
        RECT 654.150 336.300 655.950 336.750 ;
        RECT 657.450 336.300 658.500 339.750 ;
        RECT 661.050 339.000 672.900 340.050 ;
        RECT 674.100 338.100 675.300 351.600 ;
        RECT 628.350 334.500 635.100 336.300 ;
        RECT 636.000 334.500 642.900 336.300 ;
        RECT 654.150 335.850 658.500 336.300 ;
        RECT 650.850 335.100 658.500 335.850 ;
        RECT 660.000 337.200 675.300 338.100 ;
        RECT 650.850 334.950 655.950 335.100 ;
        RECT 650.850 333.600 651.750 334.950 ;
        RECT 660.000 334.050 661.050 337.200 ;
        RECT 669.300 335.700 671.100 336.300 ;
        RECT 613.650 327.750 615.450 333.600 ;
        RECT 619.050 327.750 620.850 333.600 ;
        RECT 622.200 332.400 626.400 333.600 ;
        RECT 624.600 327.750 626.400 332.400 ;
        RECT 628.950 331.500 631.050 333.600 ;
        RECT 631.950 331.500 634.050 333.600 ;
        RECT 634.950 331.500 637.050 333.600 ;
        RECT 639.750 333.300 641.850 333.600 ;
        RECT 629.250 327.750 631.050 331.500 ;
        RECT 632.250 327.750 634.050 331.500 ;
        RECT 635.250 327.750 637.050 331.500 ;
        RECT 639.000 331.500 641.850 333.300 ;
        RECT 643.950 333.300 646.050 333.600 ;
        RECT 643.950 331.500 646.800 333.300 ;
        RECT 647.700 332.250 651.750 333.600 ;
        RECT 647.700 331.800 649.500 332.250 ;
        RECT 652.950 331.950 655.050 334.050 ;
        RECT 655.950 331.950 658.050 334.050 ;
        RECT 658.950 331.950 661.050 334.050 ;
        RECT 662.700 334.500 671.100 335.700 ;
        RECT 662.700 333.600 664.200 334.500 ;
        RECT 674.100 333.600 675.300 337.200 ;
        RECT 639.000 327.750 640.800 331.500 ;
        RECT 642.000 327.750 643.800 330.600 ;
        RECT 645.000 327.750 646.800 331.500 ;
        RECT 652.950 330.600 654.300 331.950 ;
        RECT 655.950 330.600 657.300 331.950 ;
        RECT 658.950 330.600 660.300 331.950 ;
        RECT 649.500 327.750 651.300 330.600 ;
        RECT 652.500 327.750 654.300 330.600 ;
        RECT 655.500 327.750 657.300 330.600 ;
        RECT 658.500 327.750 660.300 330.600 ;
        RECT 662.700 327.750 664.500 333.600 ;
        RECT 668.100 327.750 669.900 333.600 ;
        RECT 673.500 327.750 675.300 333.600 ;
        RECT 677.700 351.600 681.750 352.500 ;
        RECT 677.700 338.100 678.900 351.600 ;
        RECT 686.700 350.700 688.500 359.250 ;
        RECT 689.700 355.950 691.500 359.250 ;
        RECT 692.850 356.400 695.250 359.250 ;
        RECT 696.150 356.400 698.250 359.250 ;
        RECT 699.300 356.400 701.250 359.250 ;
        RECT 692.850 355.050 694.050 356.400 ;
        RECT 696.150 355.050 697.050 356.400 ;
        RECT 699.300 355.050 700.500 356.400 ;
        RECT 691.950 352.950 694.050 355.050 ;
        RECT 694.950 352.950 697.050 355.050 ;
        RECT 697.950 353.400 700.500 355.050 ;
        RECT 702.450 353.400 704.250 359.250 ;
        RECT 706.200 353.400 708.000 359.250 ;
        RECT 709.200 353.400 711.000 359.250 ;
        RECT 697.950 352.950 700.050 353.400 ;
        RECT 706.650 352.500 708.000 353.400 ;
        RECT 712.200 352.500 714.000 359.250 ;
        RECT 715.950 356.400 717.750 359.250 ;
        RECT 706.650 350.850 709.050 352.500 ;
        RECT 682.200 349.650 699.900 350.700 ;
        RECT 706.950 350.400 709.050 350.850 ;
        RECT 711.000 352.200 714.000 352.500 ;
        RECT 711.000 350.400 714.900 352.200 ;
        RECT 682.200 348.900 684.000 349.650 ;
        RECT 694.950 348.150 697.050 348.750 ;
        RECT 685.500 346.950 697.050 348.150 ;
        RECT 697.950 348.600 699.900 349.650 ;
        RECT 716.100 349.350 717.450 356.400 ;
        RECT 718.950 352.950 720.750 359.250 ;
        RECT 721.950 356.400 723.750 359.250 ;
        RECT 722.100 355.200 723.600 356.400 ;
        RECT 722.100 353.100 724.200 355.200 ;
        RECT 725.700 353.400 727.500 359.250 ;
        RECT 718.950 352.050 721.050 352.950 ;
        RECT 728.700 352.500 730.500 359.250 ;
        RECT 731.700 353.400 733.500 359.250 ;
        RECT 734.700 353.400 736.500 359.250 ;
        RECT 737.700 353.400 739.500 359.250 ;
        RECT 741.450 353.400 743.250 359.250 ;
        RECT 744.450 353.400 746.250 359.250 ;
        RECT 725.850 352.050 727.650 352.500 ;
        RECT 718.950 350.850 727.650 352.050 ;
        RECT 728.700 351.300 734.400 352.500 ;
        RECT 725.850 350.700 727.650 350.850 ;
        RECT 732.600 350.700 734.400 351.300 ;
        RECT 735.300 349.350 736.500 353.400 ;
        RECT 715.950 348.600 718.050 349.350 ;
        RECT 697.950 347.250 718.050 348.600 ;
        RECT 721.950 348.450 739.350 349.350 ;
        RECT 721.950 347.250 724.050 348.450 ;
        RECT 685.500 346.350 687.300 346.950 ;
        RECT 694.950 346.650 697.050 346.950 ;
        RECT 724.950 346.350 737.250 347.550 ;
        RECT 697.950 345.450 726.000 346.350 ;
        RECT 735.450 345.750 737.250 346.350 ;
        RECT 686.250 345.150 726.000 345.450 ;
        RECT 685.950 344.550 699.900 345.150 ;
        RECT 679.950 341.850 682.050 343.950 ;
        RECT 685.950 343.350 689.850 344.550 ;
        RECT 706.950 343.650 721.500 344.250 ;
        RECT 685.950 343.050 688.050 343.350 ;
        RECT 690.750 342.450 697.500 343.350 ;
        RECT 680.100 340.050 681.900 341.850 ;
        RECT 690.750 340.050 691.950 342.450 ;
        RECT 680.100 339.000 691.950 340.050 ;
        RECT 693.750 339.750 695.550 341.550 ;
        RECT 696.450 340.950 697.500 342.450 ;
        RECT 698.400 343.050 721.500 343.650 ;
        RECT 698.400 342.450 709.050 343.050 ;
        RECT 698.400 341.850 700.200 342.450 ;
        RECT 706.950 342.150 709.050 342.450 ;
        RECT 711.150 341.250 713.250 341.550 ;
        RECT 719.700 341.250 721.500 343.050 ;
        RECT 722.850 342.000 729.900 343.800 ;
        RECT 696.450 340.050 708.450 340.950 ;
        RECT 677.700 337.200 693.000 338.100 ;
        RECT 677.700 333.600 678.900 337.200 ;
        RECT 681.900 335.700 683.700 336.300 ;
        RECT 681.900 334.500 690.300 335.700 ;
        RECT 688.800 333.600 690.300 334.500 ;
        RECT 677.700 327.750 679.500 333.600 ;
        RECT 683.100 327.750 684.900 333.600 ;
        RECT 688.500 327.750 690.300 333.600 ;
        RECT 691.950 334.050 693.000 337.200 ;
        RECT 694.500 336.300 695.550 339.750 ;
        RECT 702.150 337.350 706.050 339.150 ;
        RECT 703.950 337.050 706.050 337.350 ;
        RECT 707.400 338.550 708.450 340.050 ;
        RECT 709.350 339.450 713.250 341.250 ;
        RECT 722.850 340.350 723.750 342.000 ;
        RECT 730.950 341.100 733.050 345.150 ;
        RECT 714.150 339.300 723.750 340.350 ;
        RECT 724.800 340.050 733.050 341.100 ;
        RECT 714.150 338.550 715.050 339.300 ;
        RECT 707.400 337.200 715.050 338.550 ;
        RECT 724.800 338.250 725.850 340.050 ;
        RECT 715.950 337.200 725.850 338.250 ;
        RECT 729.300 337.200 737.100 339.000 ;
        RECT 697.050 336.300 698.850 336.750 ;
        RECT 715.950 336.300 717.000 337.200 ;
        RECT 694.500 335.850 698.850 336.300 ;
        RECT 694.500 335.100 702.150 335.850 ;
        RECT 697.050 334.950 702.150 335.100 ;
        RECT 691.950 331.950 694.050 334.050 ;
        RECT 694.950 331.950 697.050 334.050 ;
        RECT 697.950 331.950 700.050 334.050 ;
        RECT 701.250 333.600 702.150 334.950 ;
        RECT 710.100 334.500 717.000 336.300 ;
        RECT 717.900 334.500 724.650 336.300 ;
        RECT 729.300 333.600 730.800 337.200 ;
        RECT 738.150 333.600 739.350 348.450 ;
        RECT 701.250 332.250 705.300 333.600 ;
        RECT 706.950 333.300 709.050 333.600 ;
        RECT 692.700 330.600 694.050 331.950 ;
        RECT 695.700 330.600 697.050 331.950 ;
        RECT 698.700 330.600 700.050 331.950 ;
        RECT 703.500 331.800 705.300 332.250 ;
        RECT 706.200 331.500 709.050 333.300 ;
        RECT 711.150 333.300 713.250 333.600 ;
        RECT 711.150 331.500 714.000 333.300 ;
        RECT 692.700 327.750 694.500 330.600 ;
        RECT 695.700 327.750 697.500 330.600 ;
        RECT 698.700 327.750 700.500 330.600 ;
        RECT 701.700 327.750 703.500 330.600 ;
        RECT 706.200 327.750 708.000 331.500 ;
        RECT 709.200 327.750 711.000 330.600 ;
        RECT 712.200 327.750 714.000 331.500 ;
        RECT 715.950 331.500 718.050 333.600 ;
        RECT 718.950 331.500 721.050 333.600 ;
        RECT 721.950 331.500 724.050 333.600 ;
        RECT 726.600 332.400 730.800 333.600 ;
        RECT 715.950 327.750 717.750 331.500 ;
        RECT 718.950 327.750 720.750 331.500 ;
        RECT 721.950 327.750 723.750 331.500 ;
        RECT 726.600 327.750 728.400 332.400 ;
        RECT 732.150 327.750 733.950 333.600 ;
        RECT 737.550 327.750 739.350 333.600 ;
        RECT 741.450 340.950 742.950 353.400 ;
        RECT 759.450 347.400 761.250 359.250 ;
        RECT 763.650 347.400 765.450 359.250 ;
        RECT 773.550 347.400 775.350 359.250 ;
        RECT 777.750 347.400 779.550 359.250 ;
        RECT 791.550 353.400 793.350 359.250 ;
        RECT 794.550 353.400 796.350 359.250 ;
        RECT 797.550 354.000 799.350 359.250 ;
        RECT 794.700 353.100 796.350 353.400 ;
        RECT 800.550 353.400 802.350 359.250 ;
        RECT 809.400 353.400 811.200 359.250 ;
        RECT 800.550 353.100 801.750 353.400 ;
        RECT 794.700 352.200 801.750 353.100 ;
        RECT 794.100 348.150 795.900 349.950 ;
        RECT 759.450 346.350 762.000 347.400 ;
        RECT 758.100 342.150 759.900 343.950 ;
        RECT 741.450 338.850 745.050 340.950 ;
        RECT 757.950 340.050 760.050 342.150 ;
        RECT 760.950 339.150 762.000 346.350 ;
        RECT 777.000 346.350 779.550 347.400 ;
        RECT 764.100 342.150 765.900 343.950 ;
        RECT 773.100 342.150 774.900 343.950 ;
        RECT 763.950 340.050 766.050 342.150 ;
        RECT 772.950 340.050 775.050 342.150 ;
        RECT 777.000 339.150 778.050 346.350 ;
        RECT 791.100 345.150 792.900 346.950 ;
        RECT 793.950 346.050 796.050 348.150 ;
        RECT 797.250 345.150 799.050 346.950 ;
        RECT 779.100 342.150 780.900 343.950 ;
        RECT 790.950 343.050 793.050 345.150 ;
        RECT 796.950 343.050 799.050 345.150 ;
        RECT 800.700 343.950 801.750 352.200 ;
        RECT 812.700 347.400 814.500 359.250 ;
        RECT 816.900 347.400 818.700 359.250 ;
        RECT 828.450 347.400 830.250 359.250 ;
        RECT 832.650 347.400 834.450 359.250 ;
        RECT 839.550 347.400 841.350 359.250 ;
        RECT 843.750 347.400 845.550 359.250 ;
        RECT 809.250 345.150 811.050 346.950 ;
        RECT 778.950 340.050 781.050 342.150 ;
        RECT 799.950 341.850 802.050 343.950 ;
        RECT 808.950 343.050 811.050 345.150 ;
        RECT 812.850 342.150 814.050 347.400 ;
        RECT 828.450 346.350 831.000 347.400 ;
        RECT 818.100 342.150 819.900 343.950 ;
        RECT 827.100 342.150 828.900 343.950 ;
        RECT 741.450 330.600 742.950 338.850 ;
        RECT 760.950 337.050 763.050 339.150 ;
        RECT 775.950 337.050 778.050 339.150 ;
        RECT 784.950 339.450 787.050 340.050 ;
        RECT 790.950 339.450 793.050 340.050 ;
        RECT 784.950 338.550 793.050 339.450 ;
        RECT 784.950 337.950 787.050 338.550 ;
        RECT 790.950 337.950 793.050 338.550 ;
        RECT 800.400 337.650 801.600 341.850 ;
        RECT 760.950 330.600 762.000 337.050 ;
        RECT 777.000 330.600 778.050 337.050 ;
        RECT 741.450 327.750 743.250 330.600 ;
        RECT 744.450 327.750 746.250 330.600 ;
        RECT 757.650 327.750 759.450 330.600 ;
        RECT 760.650 327.750 762.450 330.600 ;
        RECT 763.650 327.750 765.450 330.600 ;
        RECT 773.550 327.750 775.350 330.600 ;
        RECT 776.550 327.750 778.350 330.600 ;
        RECT 779.550 327.750 781.350 330.600 ;
        RECT 791.700 327.750 793.500 336.600 ;
        RECT 797.100 336.000 801.600 337.650 ;
        RECT 811.950 340.050 814.050 342.150 ;
        RECT 811.950 336.750 813.150 340.050 ;
        RECT 814.950 338.850 817.050 340.950 ;
        RECT 817.950 340.050 820.050 342.150 ;
        RECT 826.950 340.050 829.050 342.150 ;
        RECT 829.950 339.150 831.000 346.350 ;
        RECT 843.000 346.350 845.550 347.400 ;
        RECT 833.100 342.150 834.900 343.950 ;
        RECT 839.100 342.150 840.900 343.950 ;
        RECT 832.950 340.050 835.050 342.150 ;
        RECT 838.950 340.050 841.050 342.150 ;
        RECT 843.000 339.150 844.050 346.350 ;
        RECT 845.100 342.150 846.900 343.950 ;
        RECT 844.950 340.050 847.050 342.150 ;
        RECT 815.100 337.050 816.900 338.850 ;
        RECT 829.950 337.050 832.050 339.150 ;
        RECT 841.950 337.050 844.050 339.150 ;
        RECT 797.100 327.750 798.900 336.000 ;
        RECT 809.250 335.700 813.000 336.750 ;
        RECT 809.250 333.600 810.450 335.700 ;
        RECT 808.650 327.750 810.450 333.600 ;
        RECT 811.650 332.700 819.450 334.050 ;
        RECT 811.650 327.750 813.450 332.700 ;
        RECT 814.650 327.750 816.450 331.800 ;
        RECT 817.650 327.750 819.450 332.700 ;
        RECT 829.950 330.600 831.000 337.050 ;
        RECT 843.000 330.600 844.050 337.050 ;
        RECT 826.650 327.750 828.450 330.600 ;
        RECT 829.650 327.750 831.450 330.600 ;
        RECT 832.650 327.750 834.450 330.600 ;
        RECT 839.550 327.750 841.350 330.600 ;
        RECT 842.550 327.750 844.350 330.600 ;
        RECT 845.550 327.750 847.350 330.600 ;
        RECT 10.800 317.400 12.600 323.250 ;
        RECT 15.000 317.400 16.800 323.250 ;
        RECT 19.200 317.400 21.000 323.250 ;
        RECT 26.550 317.400 28.350 323.250 ;
        RECT 29.550 317.400 31.350 323.250 ;
        RECT 41.850 317.400 43.650 323.250 ;
        RECT 11.250 312.150 13.050 313.950 ;
        RECT 7.950 308.850 10.050 310.950 ;
        RECT 10.950 310.050 13.050 312.150 ;
        RECT 15.000 310.950 16.050 317.400 ;
        RECT 13.950 308.850 16.050 310.950 ;
        RECT 16.950 312.150 18.750 313.950 ;
        RECT 26.100 312.150 27.900 313.950 ;
        RECT 16.950 310.050 19.050 312.150 ;
        RECT 19.950 308.850 22.050 310.950 ;
        RECT 25.950 310.050 28.050 312.150 ;
        RECT 29.400 310.950 30.600 317.400 ;
        RECT 46.350 316.200 48.150 323.250 ;
        RECT 54.000 317.400 55.800 323.250 ;
        RECT 58.200 319.050 60.000 323.250 ;
        RECT 61.500 320.400 63.300 323.250 ;
        RECT 58.200 317.400 63.900 319.050 ;
        RECT 44.550 315.300 48.150 316.200 ;
        RECT 28.950 308.850 31.050 310.950 ;
        RECT 41.100 309.150 42.900 310.950 ;
        RECT 8.100 307.050 9.900 308.850 ;
        RECT 13.950 305.400 14.850 308.850 ;
        RECT 19.950 307.050 21.750 308.850 ;
        RECT 10.800 304.500 14.850 305.400 ;
        RECT 10.800 303.600 12.600 304.500 ;
        RECT 29.400 303.600 30.600 308.850 ;
        RECT 40.950 307.050 43.050 309.150 ;
        RECT 44.550 307.950 45.750 315.300 ;
        RECT 53.100 312.150 54.900 313.950 ;
        RECT 47.100 309.150 48.900 310.950 ;
        RECT 52.950 310.050 55.050 312.150 ;
        RECT 55.950 311.850 58.050 313.950 ;
        RECT 59.100 312.150 60.900 313.950 ;
        RECT 56.100 310.050 57.900 311.850 ;
        RECT 58.950 310.050 61.050 312.150 ;
        RECT 62.700 310.950 63.900 317.400 ;
        RECT 68.550 318.300 70.350 323.250 ;
        RECT 71.550 319.200 73.350 323.250 ;
        RECT 74.550 318.300 76.350 323.250 ;
        RECT 68.550 316.950 76.350 318.300 ;
        RECT 77.550 317.400 79.350 323.250 ;
        RECT 85.650 320.400 87.450 323.250 ;
        RECT 88.650 320.400 90.450 323.250 ;
        RECT 91.650 320.400 93.450 323.250 ;
        RECT 104.700 320.400 106.500 323.250 ;
        RECT 77.550 315.300 78.750 317.400 ;
        RECT 75.000 314.250 78.750 315.300 ;
        RECT 71.100 312.150 72.900 313.950 ;
        RECT 43.950 305.850 46.050 307.950 ;
        RECT 46.950 307.050 49.050 309.150 ;
        RECT 61.950 308.850 64.050 310.950 ;
        RECT 67.950 308.850 70.050 310.950 ;
        RECT 70.950 310.050 73.050 312.150 ;
        RECT 74.850 310.950 76.050 314.250 ;
        RECT 88.950 313.950 90.000 320.400 ;
        RECT 108.000 319.050 109.800 323.250 ;
        RECT 104.100 317.400 109.800 319.050 ;
        RECT 112.200 317.400 114.000 323.250 ;
        RECT 116.550 320.400 118.350 323.250 ;
        RECT 119.550 320.400 121.350 323.250 ;
        RECT 122.550 320.400 124.350 323.250 ;
        RECT 88.950 311.850 91.050 313.950 ;
        RECT 73.950 308.850 76.050 310.950 ;
        RECT 85.950 308.850 88.050 310.950 ;
        RECT 7.650 292.500 9.450 303.600 ;
        RECT 10.650 293.400 12.450 303.600 ;
        RECT 13.650 302.400 21.450 303.300 ;
        RECT 13.650 292.500 15.450 302.400 ;
        RECT 7.650 291.750 15.450 292.500 ;
        RECT 16.650 291.750 18.450 301.500 ;
        RECT 19.650 291.750 21.450 302.400 ;
        RECT 26.550 291.750 28.350 303.600 ;
        RECT 29.550 291.750 31.350 303.600 ;
        RECT 44.550 297.600 45.750 305.850 ;
        RECT 62.700 303.600 63.900 308.850 ;
        RECT 68.100 307.050 69.900 308.850 ;
        RECT 73.950 303.600 75.150 308.850 ;
        RECT 76.950 305.850 79.050 307.950 ;
        RECT 86.100 307.050 87.900 308.850 ;
        RECT 76.950 304.050 78.750 305.850 ;
        RECT 88.950 304.650 90.000 311.850 ;
        RECT 104.100 310.950 105.300 317.400 ;
        RECT 120.000 313.950 121.050 320.400 ;
        RECT 134.850 316.200 136.650 323.250 ;
        RECT 139.350 317.400 141.150 323.250 ;
        RECT 134.850 315.300 138.450 316.200 ;
        RECT 107.100 312.150 108.900 313.950 ;
        RECT 91.950 308.850 94.050 310.950 ;
        RECT 103.950 308.850 106.050 310.950 ;
        RECT 106.950 310.050 109.050 312.150 ;
        RECT 109.950 311.850 112.050 313.950 ;
        RECT 113.100 312.150 114.900 313.950 ;
        RECT 110.100 310.050 111.900 311.850 ;
        RECT 112.950 310.050 115.050 312.150 ;
        RECT 118.950 311.850 121.050 313.950 ;
        RECT 115.950 308.850 118.050 310.950 ;
        RECT 92.100 307.050 93.900 308.850 ;
        RECT 87.450 303.600 90.000 304.650 ;
        RECT 104.100 303.600 105.300 308.850 ;
        RECT 116.100 307.050 117.900 308.850 ;
        RECT 120.000 304.650 121.050 311.850 ;
        RECT 121.950 308.850 124.050 310.950 ;
        RECT 134.100 309.150 135.900 310.950 ;
        RECT 122.100 307.050 123.900 308.850 ;
        RECT 133.950 307.050 136.050 309.150 ;
        RECT 137.250 307.950 138.450 315.300 ;
        RECT 152.100 315.000 153.900 323.250 ;
        RECT 149.400 313.350 153.900 315.000 ;
        RECT 157.500 314.400 159.300 323.250 ;
        RECT 169.650 317.400 171.450 323.250 ;
        RECT 170.250 315.300 171.450 317.400 ;
        RECT 172.650 318.300 174.450 323.250 ;
        RECT 175.650 319.200 177.450 323.250 ;
        RECT 178.650 318.300 180.450 323.250 ;
        RECT 185.550 320.400 187.350 323.250 ;
        RECT 188.550 320.400 190.350 323.250 ;
        RECT 172.650 316.950 180.450 318.300 ;
        RECT 170.250 314.250 174.000 315.300 ;
        RECT 140.100 309.150 141.900 310.950 ;
        RECT 149.400 309.150 150.600 313.350 ;
        RECT 154.950 312.450 157.050 313.050 ;
        RECT 163.950 312.450 166.050 313.050 ;
        RECT 169.950 312.450 172.050 313.050 ;
        RECT 154.950 311.550 162.450 312.450 ;
        RECT 154.950 310.950 157.050 311.550 ;
        RECT 136.950 305.850 139.050 307.950 ;
        RECT 139.950 307.050 142.050 309.150 ;
        RECT 148.950 307.050 151.050 309.150 ;
        RECT 120.000 303.600 122.550 304.650 ;
        RECT 53.550 302.700 61.350 303.600 ;
        RECT 41.550 291.750 43.350 297.600 ;
        RECT 44.550 291.750 46.350 297.600 ;
        RECT 47.550 291.750 49.350 297.600 ;
        RECT 53.550 291.750 55.350 302.700 ;
        RECT 56.550 291.750 58.350 301.800 ;
        RECT 59.550 291.750 61.350 302.700 ;
        RECT 62.550 291.750 64.350 303.600 ;
        RECT 69.300 291.750 71.100 303.600 ;
        RECT 73.500 291.750 75.300 303.600 ;
        RECT 76.800 291.750 78.600 297.600 ;
        RECT 87.450 291.750 89.250 303.600 ;
        RECT 91.650 291.750 93.450 303.600 ;
        RECT 103.650 291.750 105.450 303.600 ;
        RECT 106.650 302.700 114.450 303.600 ;
        RECT 106.650 291.750 108.450 302.700 ;
        RECT 109.650 291.750 111.450 301.800 ;
        RECT 112.650 291.750 114.450 302.700 ;
        RECT 116.550 291.750 118.350 303.600 ;
        RECT 120.750 291.750 122.550 303.600 ;
        RECT 137.250 297.600 138.450 305.850 ;
        RECT 149.250 298.800 150.300 307.050 ;
        RECT 151.950 305.850 154.050 307.950 ;
        RECT 157.950 305.850 160.050 307.950 ;
        RECT 161.550 307.050 162.450 311.550 ;
        RECT 163.950 311.550 172.050 312.450 ;
        RECT 163.950 310.950 166.050 311.550 ;
        RECT 169.950 310.950 172.050 311.550 ;
        RECT 172.950 310.950 174.150 314.250 ;
        RECT 176.100 312.150 177.900 313.950 ;
        RECT 172.950 308.850 175.050 310.950 ;
        RECT 175.950 310.050 178.050 312.150 ;
        RECT 184.950 311.850 187.050 313.950 ;
        RECT 188.400 312.150 189.600 320.400 ;
        RECT 201.000 317.400 202.800 323.250 ;
        RECT 205.200 317.400 207.000 323.250 ;
        RECT 209.400 317.400 211.200 323.250 ;
        RECT 222.000 317.400 223.800 323.250 ;
        RECT 226.200 317.400 228.000 323.250 ;
        RECT 230.400 317.400 232.200 323.250 ;
        RECT 235.950 319.950 238.050 322.050 ;
        RECT 203.250 312.150 205.050 313.950 ;
        RECT 178.950 308.850 181.050 310.950 ;
        RECT 185.100 310.050 186.900 311.850 ;
        RECT 187.950 310.050 190.050 312.150 ;
        RECT 151.950 304.050 153.750 305.850 ;
        RECT 154.950 302.850 157.050 304.950 ;
        RECT 158.100 304.050 159.900 305.850 ;
        RECT 160.950 304.950 163.050 307.050 ;
        RECT 169.950 305.850 172.050 307.950 ;
        RECT 170.250 304.050 172.050 305.850 ;
        RECT 173.850 303.600 175.050 308.850 ;
        RECT 179.100 307.050 180.900 308.850 ;
        RECT 155.100 301.050 156.900 302.850 ;
        RECT 149.250 297.900 156.300 298.800 ;
        RECT 149.250 297.600 150.450 297.900 ;
        RECT 133.650 291.750 135.450 297.600 ;
        RECT 136.650 291.750 138.450 297.600 ;
        RECT 139.650 291.750 141.450 297.600 ;
        RECT 148.650 291.750 150.450 297.600 ;
        RECT 154.650 297.600 156.300 297.900 ;
        RECT 151.650 291.750 153.450 297.000 ;
        RECT 154.650 291.750 156.450 297.600 ;
        RECT 157.650 291.750 159.450 297.600 ;
        RECT 170.400 291.750 172.200 297.600 ;
        RECT 173.700 291.750 175.500 303.600 ;
        RECT 177.900 291.750 179.700 303.600 ;
        RECT 188.400 297.600 189.600 310.050 ;
        RECT 199.950 308.850 202.050 310.950 ;
        RECT 202.950 310.050 205.050 312.150 ;
        RECT 205.950 310.950 207.000 317.400 ;
        RECT 208.950 312.150 210.750 313.950 ;
        RECT 224.250 312.150 226.050 313.950 ;
        RECT 205.950 308.850 208.050 310.950 ;
        RECT 208.950 310.050 211.050 312.150 ;
        RECT 211.950 308.850 214.050 310.950 ;
        RECT 220.950 308.850 223.050 310.950 ;
        RECT 223.950 310.050 226.050 312.150 ;
        RECT 226.950 310.950 228.000 317.400 ;
        RECT 229.950 312.150 231.750 313.950 ;
        RECT 226.950 308.850 229.050 310.950 ;
        RECT 229.950 310.050 232.050 312.150 ;
        RECT 232.950 308.850 235.050 310.950 ;
        RECT 200.250 307.050 202.050 308.850 ;
        RECT 207.150 305.400 208.050 308.850 ;
        RECT 212.100 307.050 213.900 308.850 ;
        RECT 221.250 307.050 223.050 308.850 ;
        RECT 228.150 305.400 229.050 308.850 ;
        RECT 233.100 307.050 234.900 308.850 ;
        RECT 236.550 306.450 237.450 319.950 ;
        RECT 243.000 317.400 244.800 323.250 ;
        RECT 247.200 319.050 249.000 323.250 ;
        RECT 250.500 320.400 252.300 323.250 ;
        RECT 247.200 317.400 252.900 319.050 ;
        RECT 242.100 312.150 243.900 313.950 ;
        RECT 241.950 310.050 244.050 312.150 ;
        RECT 244.950 311.850 247.050 313.950 ;
        RECT 248.100 312.150 249.900 313.950 ;
        RECT 245.100 310.050 246.900 311.850 ;
        RECT 247.950 310.050 250.050 312.150 ;
        RECT 251.700 310.950 252.900 317.400 ;
        RECT 260.550 318.000 262.350 323.250 ;
        RECT 263.550 318.900 265.350 323.250 ;
        RECT 266.550 322.500 274.350 323.250 ;
        RECT 266.550 318.000 268.350 322.500 ;
        RECT 260.550 317.100 268.350 318.000 ;
        RECT 269.550 317.400 271.350 321.600 ;
        RECT 272.550 317.400 274.350 322.500 ;
        RECT 283.650 320.400 285.450 323.250 ;
        RECT 286.650 320.400 288.450 323.250 ;
        RECT 289.650 320.400 291.450 323.250 ;
        RECT 296.550 320.400 298.350 323.250 ;
        RECT 299.550 320.400 301.350 323.250 ;
        RECT 302.550 320.400 304.350 323.250 ;
        RECT 314.700 320.400 316.500 323.250 ;
        RECT 269.850 315.900 270.750 317.400 ;
        RECT 266.400 314.850 270.750 315.900 ;
        RECT 263.100 312.150 264.900 313.950 ;
        RECT 250.950 308.850 253.050 310.950 ;
        RECT 259.950 308.850 262.050 310.950 ;
        RECT 262.950 310.050 265.050 312.150 ;
        RECT 266.400 310.950 267.600 314.850 ;
        RECT 286.950 313.950 288.000 320.400 ;
        RECT 300.000 313.950 301.050 320.400 ;
        RECT 318.000 319.050 319.800 323.250 ;
        RECT 268.500 312.150 270.300 313.950 ;
        RECT 265.950 308.850 268.050 310.950 ;
        RECT 268.950 310.050 271.050 312.150 ;
        RECT 286.950 311.850 289.050 313.950 ;
        RECT 298.950 311.850 301.050 313.950 ;
        RECT 271.950 308.850 274.050 310.950 ;
        RECT 283.950 308.850 286.050 310.950 ;
        RECT 238.950 306.450 241.050 307.050 ;
        RECT 236.550 305.550 241.050 306.450 ;
        RECT 207.150 304.500 211.200 305.400 ;
        RECT 228.150 304.500 232.200 305.400 ;
        RECT 238.950 304.950 241.050 305.550 ;
        RECT 209.400 303.600 211.200 304.500 ;
        RECT 230.400 303.600 232.200 304.500 ;
        RECT 251.700 303.600 252.900 308.850 ;
        RECT 260.100 307.050 261.900 308.850 ;
        RECT 266.550 303.600 267.750 308.850 ;
        RECT 271.950 307.050 273.750 308.850 ;
        RECT 284.100 307.050 285.900 308.850 ;
        RECT 286.950 304.650 288.000 311.850 ;
        RECT 289.950 308.850 292.050 310.950 ;
        RECT 295.950 308.850 298.050 310.950 ;
        RECT 290.100 307.050 291.900 308.850 ;
        RECT 296.100 307.050 297.900 308.850 ;
        RECT 285.450 303.600 288.000 304.650 ;
        RECT 300.000 304.650 301.050 311.850 ;
        RECT 314.100 317.400 319.800 319.050 ;
        RECT 322.200 317.400 324.000 323.250 ;
        RECT 314.100 310.950 315.300 317.400 ;
        RECT 332.850 316.200 334.650 323.250 ;
        RECT 337.350 317.400 339.150 323.250 ;
        RECT 347.850 316.200 349.650 323.250 ;
        RECT 352.350 317.400 354.150 323.250 ;
        RECT 361.650 317.400 363.450 323.250 ;
        RECT 332.850 315.300 336.450 316.200 ;
        RECT 347.850 315.300 351.450 316.200 ;
        RECT 317.100 312.150 318.900 313.950 ;
        RECT 301.950 308.850 304.050 310.950 ;
        RECT 313.950 308.850 316.050 310.950 ;
        RECT 316.950 310.050 319.050 312.150 ;
        RECT 319.950 311.850 322.050 313.950 ;
        RECT 323.100 312.150 324.900 313.950 ;
        RECT 320.100 310.050 321.900 311.850 ;
        RECT 322.950 310.050 325.050 312.150 ;
        RECT 332.100 309.150 333.900 310.950 ;
        RECT 302.100 307.050 303.900 308.850 ;
        RECT 300.000 303.600 302.550 304.650 ;
        RECT 314.100 303.600 315.300 308.850 ;
        RECT 331.950 307.050 334.050 309.150 ;
        RECT 335.250 307.950 336.450 315.300 ;
        RECT 338.100 309.150 339.900 310.950 ;
        RECT 347.100 309.150 348.900 310.950 ;
        RECT 334.950 305.850 337.050 307.950 ;
        RECT 337.950 307.050 340.050 309.150 ;
        RECT 346.950 307.050 349.050 309.150 ;
        RECT 350.250 307.950 351.450 315.300 ;
        RECT 362.250 315.300 363.450 317.400 ;
        RECT 364.650 318.300 366.450 323.250 ;
        RECT 367.650 319.200 369.450 323.250 ;
        RECT 370.650 318.300 372.450 323.250 ;
        RECT 364.650 316.950 372.450 318.300 ;
        RECT 380.850 316.200 382.650 323.250 ;
        RECT 385.350 317.400 387.150 323.250 ;
        RECT 394.650 317.400 396.450 323.250 ;
        RECT 380.850 315.300 384.450 316.200 ;
        RECT 362.250 314.250 366.000 315.300 ;
        RECT 364.950 310.950 366.150 314.250 ;
        RECT 368.100 312.150 369.900 313.950 ;
        RECT 353.100 309.150 354.900 310.950 ;
        RECT 349.950 305.850 352.050 307.950 ;
        RECT 352.950 307.050 355.050 309.150 ;
        RECT 364.950 308.850 367.050 310.950 ;
        RECT 367.950 310.050 370.050 312.150 ;
        RECT 370.950 308.850 373.050 310.950 ;
        RECT 380.100 309.150 381.900 310.950 ;
        RECT 361.950 305.850 364.050 307.950 ;
        RECT 200.550 302.400 208.350 303.300 ;
        RECT 185.550 291.750 187.350 297.600 ;
        RECT 188.550 291.750 190.350 297.600 ;
        RECT 200.550 291.750 202.350 302.400 ;
        RECT 203.550 291.750 205.350 301.500 ;
        RECT 206.550 292.500 208.350 302.400 ;
        RECT 209.550 293.400 211.350 303.600 ;
        RECT 212.550 292.500 214.350 303.600 ;
        RECT 206.550 291.750 214.350 292.500 ;
        RECT 221.550 302.400 229.350 303.300 ;
        RECT 221.550 291.750 223.350 302.400 ;
        RECT 224.550 291.750 226.350 301.500 ;
        RECT 227.550 292.500 229.350 302.400 ;
        RECT 230.550 293.400 232.350 303.600 ;
        RECT 233.550 292.500 235.350 303.600 ;
        RECT 227.550 291.750 235.350 292.500 ;
        RECT 242.550 302.700 250.350 303.600 ;
        RECT 242.550 291.750 244.350 302.700 ;
        RECT 245.550 291.750 247.350 301.800 ;
        RECT 248.550 291.750 250.350 302.700 ;
        RECT 251.550 291.750 253.350 303.600 ;
        RECT 260.550 291.750 262.350 303.600 ;
        RECT 265.050 291.750 268.350 303.600 ;
        RECT 271.050 291.750 272.850 303.600 ;
        RECT 285.450 291.750 287.250 303.600 ;
        RECT 289.650 291.750 291.450 303.600 ;
        RECT 296.550 291.750 298.350 303.600 ;
        RECT 300.750 291.750 302.550 303.600 ;
        RECT 313.650 291.750 315.450 303.600 ;
        RECT 316.650 302.700 324.450 303.600 ;
        RECT 316.650 291.750 318.450 302.700 ;
        RECT 319.650 291.750 321.450 301.800 ;
        RECT 322.650 291.750 324.450 302.700 ;
        RECT 335.250 297.600 336.450 305.850 ;
        RECT 350.250 297.600 351.450 305.850 ;
        RECT 362.250 304.050 364.050 305.850 ;
        RECT 365.850 303.600 367.050 308.850 ;
        RECT 371.100 307.050 372.900 308.850 ;
        RECT 379.950 307.050 382.050 309.150 ;
        RECT 383.250 307.950 384.450 315.300 ;
        RECT 395.250 315.300 396.450 317.400 ;
        RECT 397.650 318.300 399.450 323.250 ;
        RECT 400.650 319.200 402.450 323.250 ;
        RECT 403.650 318.300 405.450 323.250 ;
        RECT 397.650 316.950 405.450 318.300 ;
        RECT 415.800 317.400 417.600 323.250 ;
        RECT 420.000 317.400 421.800 323.250 ;
        RECT 424.200 317.400 426.000 323.250 ;
        RECT 431.550 318.000 433.350 323.250 ;
        RECT 434.550 318.900 436.350 323.250 ;
        RECT 437.550 322.500 445.350 323.250 ;
        RECT 437.550 318.000 439.350 322.500 ;
        RECT 395.250 314.250 399.000 315.300 ;
        RECT 397.950 310.950 399.150 314.250 ;
        RECT 401.100 312.150 402.900 313.950 ;
        RECT 416.250 312.150 418.050 313.950 ;
        RECT 386.100 309.150 387.900 310.950 ;
        RECT 382.950 305.850 385.050 307.950 ;
        RECT 385.950 307.050 388.050 309.150 ;
        RECT 397.950 308.850 400.050 310.950 ;
        RECT 400.950 310.050 403.050 312.150 ;
        RECT 403.950 308.850 406.050 310.950 ;
        RECT 412.950 308.850 415.050 310.950 ;
        RECT 415.950 310.050 418.050 312.150 ;
        RECT 420.000 310.950 421.050 317.400 ;
        RECT 431.550 317.100 439.350 318.000 ;
        RECT 440.550 317.400 442.350 321.600 ;
        RECT 443.550 317.400 445.350 322.500 ;
        RECT 454.650 320.400 456.450 323.250 ;
        RECT 457.650 320.400 459.450 323.250 ;
        RECT 440.850 315.900 441.750 317.400 ;
        RECT 437.400 314.850 441.750 315.900 ;
        RECT 418.950 308.850 421.050 310.950 ;
        RECT 421.950 312.150 423.750 313.950 ;
        RECT 434.100 312.150 435.900 313.950 ;
        RECT 421.950 310.050 424.050 312.150 ;
        RECT 424.950 308.850 427.050 310.950 ;
        RECT 430.950 308.850 433.050 310.950 ;
        RECT 433.950 310.050 436.050 312.150 ;
        RECT 437.400 310.950 438.600 314.850 ;
        RECT 439.500 312.150 441.300 313.950 ;
        RECT 455.400 312.150 456.600 320.400 ;
        RECT 467.550 318.300 469.350 323.250 ;
        RECT 470.550 319.200 472.350 323.250 ;
        RECT 473.550 318.300 475.350 323.250 ;
        RECT 467.550 316.950 475.350 318.300 ;
        RECT 476.550 317.400 478.350 323.250 ;
        RECT 476.550 315.300 477.750 317.400 ;
        RECT 485.850 316.200 487.650 323.250 ;
        RECT 490.350 317.400 492.150 323.250 ;
        RECT 485.850 315.300 489.450 316.200 ;
        RECT 474.000 314.250 477.750 315.300 ;
        RECT 436.950 308.850 439.050 310.950 ;
        RECT 439.950 310.050 442.050 312.150 ;
        RECT 442.950 308.850 445.050 310.950 ;
        RECT 454.950 310.050 457.050 312.150 ;
        RECT 457.950 311.850 460.050 313.950 ;
        RECT 470.100 312.150 471.900 313.950 ;
        RECT 458.100 310.050 459.900 311.850 ;
        RECT 394.950 305.850 397.050 307.950 ;
        RECT 331.650 291.750 333.450 297.600 ;
        RECT 334.650 291.750 336.450 297.600 ;
        RECT 337.650 291.750 339.450 297.600 ;
        RECT 346.650 291.750 348.450 297.600 ;
        RECT 349.650 291.750 351.450 297.600 ;
        RECT 352.650 291.750 354.450 297.600 ;
        RECT 362.400 291.750 364.200 297.600 ;
        RECT 365.700 291.750 367.500 303.600 ;
        RECT 369.900 291.750 371.700 303.600 ;
        RECT 383.250 297.600 384.450 305.850 ;
        RECT 395.250 304.050 397.050 305.850 ;
        RECT 398.850 303.600 400.050 308.850 ;
        RECT 404.100 307.050 405.900 308.850 ;
        RECT 413.100 307.050 414.900 308.850 ;
        RECT 418.950 305.400 419.850 308.850 ;
        RECT 424.950 307.050 426.750 308.850 ;
        RECT 431.100 307.050 432.900 308.850 ;
        RECT 415.800 304.500 419.850 305.400 ;
        RECT 415.800 303.600 417.600 304.500 ;
        RECT 437.550 303.600 438.750 308.850 ;
        RECT 442.950 307.050 444.750 308.850 ;
        RECT 379.650 291.750 381.450 297.600 ;
        RECT 382.650 291.750 384.450 297.600 ;
        RECT 385.650 291.750 387.450 297.600 ;
        RECT 395.400 291.750 397.200 297.600 ;
        RECT 398.700 291.750 400.500 303.600 ;
        RECT 402.900 291.750 404.700 303.600 ;
        RECT 412.650 292.500 414.450 303.600 ;
        RECT 415.650 293.400 417.450 303.600 ;
        RECT 418.650 302.400 426.450 303.300 ;
        RECT 418.650 292.500 420.450 302.400 ;
        RECT 412.650 291.750 420.450 292.500 ;
        RECT 421.650 291.750 423.450 301.500 ;
        RECT 424.650 291.750 426.450 302.400 ;
        RECT 431.550 291.750 433.350 303.600 ;
        RECT 436.050 291.750 439.350 303.600 ;
        RECT 442.050 291.750 443.850 303.600 ;
        RECT 455.400 297.600 456.600 310.050 ;
        RECT 466.950 308.850 469.050 310.950 ;
        RECT 469.950 310.050 472.050 312.150 ;
        RECT 473.850 310.950 475.050 314.250 ;
        RECT 472.950 308.850 475.050 310.950 ;
        RECT 485.100 309.150 486.900 310.950 ;
        RECT 467.100 307.050 468.900 308.850 ;
        RECT 472.950 303.600 474.150 308.850 ;
        RECT 475.950 305.850 478.050 307.950 ;
        RECT 484.950 307.050 487.050 309.150 ;
        RECT 488.250 307.950 489.450 315.300 ;
        RECT 503.100 315.000 504.900 323.250 ;
        RECT 500.400 313.350 504.900 315.000 ;
        RECT 508.500 314.400 510.300 323.250 ;
        RECT 515.550 320.400 517.350 323.250 ;
        RECT 518.550 320.400 520.350 323.250 ;
        RECT 533.250 320.400 535.350 323.250 ;
        RECT 536.550 320.400 538.350 323.250 ;
        RECT 539.550 320.400 541.350 323.250 ;
        RECT 542.550 320.400 544.350 323.250 ;
        RECT 491.100 309.150 492.900 310.950 ;
        RECT 500.400 309.150 501.600 313.350 ;
        RECT 514.950 311.850 517.050 313.950 ;
        RECT 518.400 312.150 519.600 320.400 ;
        RECT 537.300 319.500 538.350 320.400 ;
        RECT 543.300 319.500 544.350 320.400 ;
        RECT 537.300 318.600 548.100 319.500 ;
        RECT 520.950 315.450 523.050 316.050 ;
        RECT 532.950 315.450 535.050 316.050 ;
        RECT 520.950 314.550 535.050 315.450 ;
        RECT 520.950 313.950 523.050 314.550 ;
        RECT 532.950 313.950 535.050 314.550 ;
        RECT 539.100 312.150 540.900 313.950 ;
        RECT 546.900 312.150 548.100 318.600 ;
        RECT 562.650 317.400 564.450 323.250 ;
        RECT 565.650 320.400 567.450 323.250 ;
        RECT 568.650 320.400 570.450 323.250 ;
        RECT 571.650 320.400 573.450 323.250 ;
        RECT 562.950 312.150 564.000 317.400 ;
        RECT 568.650 316.200 569.550 320.400 ;
        RECT 566.250 315.300 569.550 316.200 ;
        RECT 584.850 316.200 586.650 323.250 ;
        RECT 589.350 317.400 591.150 323.250 ;
        RECT 601.650 317.400 603.450 323.250 ;
        RECT 604.650 320.400 606.450 323.250 ;
        RECT 607.650 320.400 609.450 323.250 ;
        RECT 610.650 320.400 612.450 323.250 ;
        RECT 584.850 315.300 588.450 316.200 ;
        RECT 595.950 315.450 598.050 316.050 ;
        RECT 566.250 314.400 568.050 315.300 ;
        RECT 515.100 310.050 516.900 311.850 ;
        RECT 517.950 310.050 520.050 312.150 ;
        RECT 487.950 305.850 490.050 307.950 ;
        RECT 490.950 307.050 493.050 309.150 ;
        RECT 499.950 307.050 502.050 309.150 ;
        RECT 475.950 304.050 477.750 305.850 ;
        RECT 454.650 291.750 456.450 297.600 ;
        RECT 457.650 291.750 459.450 297.600 ;
        RECT 468.300 291.750 470.100 303.600 ;
        RECT 472.500 291.750 474.300 303.600 ;
        RECT 488.250 297.600 489.450 305.850 ;
        RECT 500.250 298.800 501.300 307.050 ;
        RECT 502.950 305.850 505.050 307.950 ;
        RECT 508.950 305.850 511.050 307.950 ;
        RECT 502.950 304.050 504.750 305.850 ;
        RECT 505.950 302.850 508.050 304.950 ;
        RECT 509.100 304.050 510.900 305.850 ;
        RECT 506.100 301.050 507.900 302.850 ;
        RECT 500.250 297.900 507.300 298.800 ;
        RECT 500.250 297.600 501.450 297.900 ;
        RECT 475.800 291.750 477.600 297.600 ;
        RECT 484.650 291.750 486.450 297.600 ;
        RECT 487.650 291.750 489.450 297.600 ;
        RECT 490.650 291.750 492.450 297.600 ;
        RECT 499.650 291.750 501.450 297.600 ;
        RECT 505.650 297.600 507.300 297.900 ;
        RECT 518.400 297.600 519.600 310.050 ;
        RECT 532.950 308.850 535.050 310.950 ;
        RECT 538.950 310.050 541.050 312.150 ;
        RECT 541.950 308.850 544.050 310.950 ;
        RECT 546.900 310.050 550.050 312.150 ;
        RECT 562.950 310.050 565.050 312.150 ;
        RECT 533.100 307.050 534.900 308.850 ;
        RECT 542.100 307.050 543.900 308.850 ;
        RECT 546.900 304.800 548.100 310.050 ;
        RECT 546.900 303.600 550.350 304.800 ;
        RECT 530.550 301.500 538.350 302.400 ;
        RECT 502.650 291.750 504.450 297.000 ;
        RECT 505.650 291.750 507.450 297.600 ;
        RECT 508.650 291.750 510.450 297.600 ;
        RECT 515.550 291.750 517.350 297.600 ;
        RECT 518.550 291.750 520.350 297.600 ;
        RECT 530.550 291.750 532.350 301.500 ;
        RECT 533.550 291.750 535.350 300.600 ;
        RECT 536.550 292.500 538.350 301.500 ;
        RECT 539.550 301.200 547.950 302.100 ;
        RECT 539.550 293.400 541.350 301.200 ;
        RECT 542.550 292.500 544.350 300.300 ;
        RECT 536.550 291.750 544.350 292.500 ;
        RECT 546.150 292.500 547.950 301.200 ;
        RECT 549.150 301.200 550.350 303.600 ;
        RECT 563.550 303.450 564.900 310.050 ;
        RECT 566.400 306.150 567.300 314.400 ;
        RECT 571.950 311.850 574.050 313.950 ;
        RECT 568.950 308.850 571.050 310.950 ;
        RECT 572.100 310.050 573.900 311.850 ;
        RECT 584.100 309.150 585.900 310.950 ;
        RECT 569.100 307.050 570.900 308.850 ;
        RECT 583.950 307.050 586.050 309.150 ;
        RECT 587.250 307.950 588.450 315.300 ;
        RECT 593.550 314.550 598.050 315.450 ;
        RECT 590.100 309.150 591.900 310.950 ;
        RECT 566.250 306.000 568.050 306.150 ;
        RECT 566.250 304.800 573.450 306.000 ;
        RECT 586.950 305.850 589.050 307.950 ;
        RECT 589.950 307.050 592.050 309.150 ;
        RECT 566.250 304.350 568.050 304.800 ;
        RECT 572.250 303.600 573.450 304.800 ;
        RECT 563.550 302.100 565.950 303.450 ;
        RECT 549.150 293.400 550.950 301.200 ;
        RECT 552.150 292.500 553.950 301.800 ;
        RECT 546.150 291.750 553.950 292.500 ;
        RECT 564.150 291.750 565.950 302.100 ;
        RECT 567.150 291.750 568.950 303.450 ;
        RECT 571.650 291.750 573.450 303.600 ;
        RECT 587.250 297.600 588.450 305.850 ;
        RECT 589.950 303.450 592.050 304.050 ;
        RECT 593.550 303.450 594.450 314.550 ;
        RECT 595.950 313.950 598.050 314.550 ;
        RECT 601.950 312.150 603.000 317.400 ;
        RECT 607.650 316.200 608.550 320.400 ;
        RECT 614.850 317.400 616.650 323.250 ;
        RECT 619.350 316.200 621.150 323.250 ;
        RECT 632.700 320.400 634.500 323.250 ;
        RECT 636.000 319.050 637.800 323.250 ;
        RECT 605.250 315.300 608.550 316.200 ;
        RECT 617.550 315.300 621.150 316.200 ;
        RECT 632.100 317.400 637.800 319.050 ;
        RECT 640.200 317.400 642.000 323.250 ;
        RECT 647.550 318.300 649.350 323.250 ;
        RECT 650.550 319.200 652.350 323.250 ;
        RECT 653.550 318.300 655.350 323.250 ;
        RECT 605.250 314.400 607.050 315.300 ;
        RECT 601.950 310.050 604.050 312.150 ;
        RECT 589.950 302.550 594.450 303.450 ;
        RECT 602.550 303.450 603.900 310.050 ;
        RECT 605.400 306.150 606.300 314.400 ;
        RECT 610.950 311.850 613.050 313.950 ;
        RECT 607.950 308.850 610.050 310.950 ;
        RECT 611.100 310.050 612.900 311.850 ;
        RECT 614.100 309.150 615.900 310.950 ;
        RECT 608.100 307.050 609.900 308.850 ;
        RECT 613.950 307.050 616.050 309.150 ;
        RECT 617.550 307.950 618.750 315.300 ;
        RECT 632.100 310.950 633.300 317.400 ;
        RECT 647.550 316.950 655.350 318.300 ;
        RECT 656.550 317.400 658.350 323.250 ;
        RECT 670.650 320.400 672.450 323.250 ;
        RECT 673.650 320.400 675.450 323.250 ;
        RECT 676.650 320.400 678.450 323.250 ;
        RECT 656.550 315.300 657.750 317.400 ;
        RECT 654.000 314.250 657.750 315.300 ;
        RECT 635.100 312.150 636.900 313.950 ;
        RECT 620.100 309.150 621.900 310.950 ;
        RECT 605.250 306.000 607.050 306.150 ;
        RECT 605.250 304.800 612.450 306.000 ;
        RECT 616.950 305.850 619.050 307.950 ;
        RECT 619.950 307.050 622.050 309.150 ;
        RECT 631.950 308.850 634.050 310.950 ;
        RECT 634.950 310.050 637.050 312.150 ;
        RECT 637.950 311.850 640.050 313.950 ;
        RECT 641.100 312.150 642.900 313.950 ;
        RECT 650.100 312.150 651.900 313.950 ;
        RECT 638.100 310.050 639.900 311.850 ;
        RECT 640.950 310.050 643.050 312.150 ;
        RECT 646.950 308.850 649.050 310.950 ;
        RECT 649.950 310.050 652.050 312.150 ;
        RECT 653.850 310.950 655.050 314.250 ;
        RECT 673.950 313.950 675.000 320.400 ;
        RECT 683.850 316.200 685.650 323.250 ;
        RECT 688.350 317.400 690.150 323.250 ;
        RECT 700.650 317.400 702.450 323.250 ;
        RECT 676.950 315.450 679.050 316.050 ;
        RECT 676.950 314.550 681.450 315.450 ;
        RECT 683.850 315.300 687.450 316.200 ;
        RECT 676.950 313.950 679.050 314.550 ;
        RECT 673.950 311.850 676.050 313.950 ;
        RECT 652.950 308.850 655.050 310.950 ;
        RECT 670.950 308.850 673.050 310.950 ;
        RECT 605.250 304.350 607.050 304.800 ;
        RECT 611.250 303.600 612.450 304.800 ;
        RECT 589.950 301.950 592.050 302.550 ;
        RECT 602.550 302.100 604.950 303.450 ;
        RECT 583.650 291.750 585.450 297.600 ;
        RECT 586.650 291.750 588.450 297.600 ;
        RECT 589.650 291.750 591.450 297.600 ;
        RECT 603.150 291.750 604.950 302.100 ;
        RECT 606.150 291.750 607.950 303.450 ;
        RECT 610.650 291.750 612.450 303.600 ;
        RECT 617.550 297.600 618.750 305.850 ;
        RECT 632.100 303.600 633.300 308.850 ;
        RECT 647.100 307.050 648.900 308.850 ;
        RECT 652.950 303.600 654.150 308.850 ;
        RECT 655.950 305.850 658.050 307.950 ;
        RECT 671.100 307.050 672.900 308.850 ;
        RECT 655.950 304.050 657.750 305.850 ;
        RECT 673.950 304.650 675.000 311.850 ;
        RECT 676.950 308.850 679.050 310.950 ;
        RECT 677.100 307.050 678.900 308.850 ;
        RECT 672.450 303.600 675.000 304.650 ;
        RECT 680.550 304.050 681.450 314.550 ;
        RECT 683.100 309.150 684.900 310.950 ;
        RECT 682.950 307.050 685.050 309.150 ;
        RECT 686.250 307.950 687.450 315.300 ;
        RECT 701.250 315.300 702.450 317.400 ;
        RECT 703.650 318.300 705.450 323.250 ;
        RECT 706.650 319.200 708.450 323.250 ;
        RECT 709.650 318.300 711.450 323.250 ;
        RECT 719.550 320.400 721.350 323.250 ;
        RECT 703.650 316.950 711.450 318.300 ;
        RECT 720.150 316.500 721.350 320.400 ;
        RECT 722.850 317.400 724.650 323.250 ;
        RECT 725.850 317.400 727.650 323.250 ;
        RECT 739.650 320.400 741.450 323.250 ;
        RECT 742.650 320.400 744.450 323.250 ;
        RECT 720.150 315.600 725.250 316.500 ;
        RECT 701.250 314.250 705.000 315.300 ;
        RECT 723.000 314.700 725.250 315.600 ;
        RECT 703.950 310.950 705.150 314.250 ;
        RECT 707.100 312.150 708.900 313.950 ;
        RECT 689.100 309.150 690.900 310.950 ;
        RECT 685.950 305.850 688.050 307.950 ;
        RECT 688.950 307.050 691.050 309.150 ;
        RECT 703.950 308.850 706.050 310.950 ;
        RECT 706.950 310.050 709.050 312.150 ;
        RECT 709.950 308.850 712.050 310.950 ;
        RECT 718.950 308.850 721.050 310.950 ;
        RECT 700.950 305.850 703.050 307.950 ;
        RECT 614.550 291.750 616.350 297.600 ;
        RECT 617.550 291.750 619.350 297.600 ;
        RECT 620.550 291.750 622.350 297.600 ;
        RECT 631.650 291.750 633.450 303.600 ;
        RECT 634.650 302.700 642.450 303.600 ;
        RECT 634.650 291.750 636.450 302.700 ;
        RECT 637.650 291.750 639.450 301.800 ;
        RECT 640.650 291.750 642.450 302.700 ;
        RECT 648.300 291.750 650.100 303.600 ;
        RECT 652.500 291.750 654.300 303.600 ;
        RECT 655.800 291.750 657.600 297.600 ;
        RECT 672.450 291.750 674.250 303.600 ;
        RECT 676.650 291.750 678.450 303.600 ;
        RECT 679.950 301.950 682.050 304.050 ;
        RECT 686.250 297.600 687.450 305.850 ;
        RECT 701.250 304.050 703.050 305.850 ;
        RECT 704.850 303.600 706.050 308.850 ;
        RECT 710.100 307.050 711.900 308.850 ;
        RECT 719.100 307.050 720.900 308.850 ;
        RECT 723.000 306.300 724.050 314.700 ;
        RECT 726.150 310.950 727.350 317.400 ;
        RECT 740.400 312.150 741.600 320.400 ;
        RECT 755.100 315.000 756.900 323.250 ;
        RECT 724.950 308.850 727.350 310.950 ;
        RECT 739.950 310.050 742.050 312.150 ;
        RECT 742.950 311.850 745.050 313.950 ;
        RECT 752.400 313.350 756.900 315.000 ;
        RECT 760.500 314.400 762.300 323.250 ;
        RECT 766.650 320.400 768.450 323.250 ;
        RECT 769.650 320.400 771.450 323.250 ;
        RECT 772.650 320.400 774.450 323.250 ;
        RECT 769.950 313.950 771.000 320.400 ;
        RECT 782.550 318.300 784.350 323.250 ;
        RECT 785.550 319.200 787.350 323.250 ;
        RECT 788.550 318.300 790.350 323.250 ;
        RECT 782.550 316.950 790.350 318.300 ;
        RECT 791.550 317.400 793.350 323.250 ;
        RECT 791.550 315.300 792.750 317.400 ;
        RECT 789.000 314.250 792.750 315.300 ;
        RECT 803.100 315.000 804.900 323.250 ;
        RECT 743.100 310.050 744.900 311.850 ;
        RECT 723.000 305.400 725.250 306.300 ;
        RECT 719.550 304.500 725.250 305.400 ;
        RECT 682.650 291.750 684.450 297.600 ;
        RECT 685.650 291.750 687.450 297.600 ;
        RECT 688.650 291.750 690.450 297.600 ;
        RECT 701.400 291.750 703.200 297.600 ;
        RECT 704.700 291.750 706.500 303.600 ;
        RECT 708.900 291.750 710.700 303.600 ;
        RECT 719.550 297.600 720.750 304.500 ;
        RECT 726.150 303.600 727.350 308.850 ;
        RECT 719.550 291.750 721.350 297.600 ;
        RECT 722.850 291.750 724.650 303.600 ;
        RECT 725.850 291.750 727.650 303.600 ;
        RECT 740.400 297.600 741.600 310.050 ;
        RECT 752.400 309.150 753.600 313.350 ;
        RECT 769.950 311.850 772.050 313.950 ;
        RECT 785.100 312.150 786.900 313.950 ;
        RECT 751.950 307.050 754.050 309.150 ;
        RECT 766.950 308.850 769.050 310.950 ;
        RECT 752.250 298.800 753.300 307.050 ;
        RECT 754.950 305.850 757.050 307.950 ;
        RECT 760.950 305.850 763.050 307.950 ;
        RECT 767.100 307.050 768.900 308.850 ;
        RECT 754.950 304.050 756.750 305.850 ;
        RECT 757.950 302.850 760.050 304.950 ;
        RECT 761.100 304.050 762.900 305.850 ;
        RECT 769.950 304.650 771.000 311.850 ;
        RECT 772.950 308.850 775.050 310.950 ;
        RECT 781.950 308.850 784.050 310.950 ;
        RECT 784.950 310.050 787.050 312.150 ;
        RECT 788.850 310.950 790.050 314.250 ;
        RECT 787.950 308.850 790.050 310.950 ;
        RECT 800.400 313.350 804.900 315.000 ;
        RECT 808.500 314.400 810.300 323.250 ;
        RECT 814.650 317.400 816.450 323.250 ;
        RECT 817.650 320.400 819.450 323.250 ;
        RECT 820.650 320.400 822.450 323.250 ;
        RECT 823.650 320.400 825.450 323.250 ;
        RECT 800.400 309.150 801.600 313.350 ;
        RECT 814.950 312.150 816.000 317.400 ;
        RECT 820.650 316.200 821.550 320.400 ;
        RECT 833.850 317.400 835.650 323.250 ;
        RECT 838.350 316.200 840.150 323.250 ;
        RECT 848.550 320.400 850.350 323.250 ;
        RECT 851.550 320.400 853.350 323.250 ;
        RECT 854.550 320.400 856.350 323.250 ;
        RECT 818.250 315.300 821.550 316.200 ;
        RECT 836.550 315.300 840.150 316.200 ;
        RECT 818.250 314.400 820.050 315.300 ;
        RECT 814.950 310.050 817.050 312.150 ;
        RECT 773.100 307.050 774.900 308.850 ;
        RECT 782.100 307.050 783.900 308.850 ;
        RECT 768.450 303.600 771.000 304.650 ;
        RECT 787.950 303.600 789.150 308.850 ;
        RECT 790.950 305.850 793.050 307.950 ;
        RECT 799.950 307.050 802.050 309.150 ;
        RECT 790.950 304.050 792.750 305.850 ;
        RECT 758.100 301.050 759.900 302.850 ;
        RECT 752.250 297.900 759.300 298.800 ;
        RECT 752.250 297.600 753.450 297.900 ;
        RECT 739.650 291.750 741.450 297.600 ;
        RECT 742.650 291.750 744.450 297.600 ;
        RECT 751.650 291.750 753.450 297.600 ;
        RECT 757.650 297.600 759.300 297.900 ;
        RECT 754.650 291.750 756.450 297.000 ;
        RECT 757.650 291.750 759.450 297.600 ;
        RECT 760.650 291.750 762.450 297.600 ;
        RECT 768.450 291.750 770.250 303.600 ;
        RECT 772.650 291.750 774.450 303.600 ;
        RECT 783.300 291.750 785.100 303.600 ;
        RECT 787.500 291.750 789.300 303.600 ;
        RECT 800.250 298.800 801.300 307.050 ;
        RECT 802.950 305.850 805.050 307.950 ;
        RECT 808.950 305.850 811.050 307.950 ;
        RECT 802.950 304.050 804.750 305.850 ;
        RECT 805.950 302.850 808.050 304.950 ;
        RECT 809.100 304.050 810.900 305.850 ;
        RECT 815.550 303.450 816.900 310.050 ;
        RECT 818.400 306.150 819.300 314.400 ;
        RECT 823.950 311.850 826.050 313.950 ;
        RECT 820.950 308.850 823.050 310.950 ;
        RECT 824.100 310.050 825.900 311.850 ;
        RECT 833.100 309.150 834.900 310.950 ;
        RECT 821.100 307.050 822.900 308.850 ;
        RECT 832.950 307.050 835.050 309.150 ;
        RECT 836.550 307.950 837.750 315.300 ;
        RECT 852.000 313.950 853.050 320.400 ;
        RECT 850.950 311.850 853.050 313.950 ;
        RECT 839.100 309.150 840.900 310.950 ;
        RECT 818.250 306.000 820.050 306.150 ;
        RECT 818.250 304.800 825.450 306.000 ;
        RECT 835.950 305.850 838.050 307.950 ;
        RECT 838.950 307.050 841.050 309.150 ;
        RECT 847.950 308.850 850.050 310.950 ;
        RECT 848.100 307.050 849.900 308.850 ;
        RECT 818.250 304.350 820.050 304.800 ;
        RECT 824.250 303.600 825.450 304.800 ;
        RECT 806.100 301.050 807.900 302.850 ;
        RECT 815.550 302.100 817.950 303.450 ;
        RECT 800.250 297.900 807.300 298.800 ;
        RECT 800.250 297.600 801.450 297.900 ;
        RECT 790.800 291.750 792.600 297.600 ;
        RECT 799.650 291.750 801.450 297.600 ;
        RECT 805.650 297.600 807.300 297.900 ;
        RECT 802.650 291.750 804.450 297.000 ;
        RECT 805.650 291.750 807.450 297.600 ;
        RECT 808.650 291.750 810.450 297.600 ;
        RECT 816.150 291.750 817.950 302.100 ;
        RECT 819.150 291.750 820.950 303.450 ;
        RECT 823.650 291.750 825.450 303.600 ;
        RECT 836.550 297.600 837.750 305.850 ;
        RECT 852.000 304.650 853.050 311.850 ;
        RECT 853.950 308.850 856.050 310.950 ;
        RECT 854.100 307.050 855.900 308.850 ;
        RECT 852.000 303.600 854.550 304.650 ;
        RECT 833.550 291.750 835.350 297.600 ;
        RECT 836.550 291.750 838.350 297.600 ;
        RECT 839.550 291.750 841.350 297.600 ;
        RECT 848.550 291.750 850.350 303.600 ;
        RECT 852.750 291.750 854.550 303.600 ;
        RECT 2.700 281.400 4.500 287.250 ;
        RECT 5.700 281.400 7.500 287.250 ;
        RECT 8.700 281.400 10.500 287.250 ;
        RECT 5.700 280.500 6.750 281.400 ;
        RECT 2.700 279.600 6.750 280.500 ;
        RECT 2.700 266.100 3.900 279.600 ;
        RECT 11.700 278.700 13.500 287.250 ;
        RECT 14.700 283.950 16.500 287.250 ;
        RECT 17.850 284.400 20.250 287.250 ;
        RECT 21.150 284.400 23.250 287.250 ;
        RECT 24.300 284.400 26.250 287.250 ;
        RECT 17.850 283.050 19.050 284.400 ;
        RECT 21.150 283.050 22.050 284.400 ;
        RECT 24.300 283.050 25.500 284.400 ;
        RECT 16.950 280.950 19.050 283.050 ;
        RECT 19.950 280.950 22.050 283.050 ;
        RECT 22.950 281.400 25.500 283.050 ;
        RECT 27.450 281.400 29.250 287.250 ;
        RECT 31.200 281.400 33.000 287.250 ;
        RECT 34.200 281.400 36.000 287.250 ;
        RECT 22.950 280.950 25.050 281.400 ;
        RECT 31.650 280.500 33.000 281.400 ;
        RECT 37.200 280.500 39.000 287.250 ;
        RECT 40.950 284.400 42.750 287.250 ;
        RECT 31.650 278.850 34.050 280.500 ;
        RECT 7.200 277.650 24.900 278.700 ;
        RECT 31.950 278.400 34.050 278.850 ;
        RECT 36.000 280.200 39.000 280.500 ;
        RECT 36.000 278.400 39.900 280.200 ;
        RECT 7.200 276.900 9.000 277.650 ;
        RECT 19.950 276.150 22.050 276.750 ;
        RECT 10.500 274.950 22.050 276.150 ;
        RECT 22.950 276.600 24.900 277.650 ;
        RECT 41.100 277.350 42.450 284.400 ;
        RECT 43.950 280.950 45.750 287.250 ;
        RECT 46.950 284.400 48.750 287.250 ;
        RECT 47.100 283.200 48.600 284.400 ;
        RECT 47.100 281.100 49.200 283.200 ;
        RECT 50.700 281.400 52.500 287.250 ;
        RECT 43.950 280.050 46.050 280.950 ;
        RECT 53.700 280.500 55.500 287.250 ;
        RECT 56.700 281.400 58.500 287.250 ;
        RECT 59.700 281.400 61.500 287.250 ;
        RECT 62.700 281.400 64.500 287.250 ;
        RECT 66.450 281.400 68.250 287.250 ;
        RECT 69.450 281.400 71.250 287.250 ;
        RECT 76.650 281.400 78.450 287.250 ;
        RECT 79.650 282.000 81.450 287.250 ;
        RECT 50.850 280.050 52.650 280.500 ;
        RECT 43.950 278.850 52.650 280.050 ;
        RECT 53.700 279.300 59.400 280.500 ;
        RECT 50.850 278.700 52.650 278.850 ;
        RECT 57.600 278.700 59.400 279.300 ;
        RECT 60.300 277.350 61.500 281.400 ;
        RECT 40.950 276.600 43.050 277.350 ;
        RECT 22.950 275.250 43.050 276.600 ;
        RECT 46.950 276.450 64.350 277.350 ;
        RECT 46.950 275.250 49.050 276.450 ;
        RECT 10.500 274.350 12.300 274.950 ;
        RECT 19.950 274.650 22.050 274.950 ;
        RECT 49.950 274.350 62.250 275.550 ;
        RECT 22.950 273.450 51.000 274.350 ;
        RECT 60.450 273.750 62.250 274.350 ;
        RECT 11.250 273.150 51.000 273.450 ;
        RECT 10.950 272.550 24.900 273.150 ;
        RECT 4.950 269.850 7.050 271.950 ;
        RECT 10.950 271.350 14.850 272.550 ;
        RECT 31.950 271.650 46.500 272.250 ;
        RECT 10.950 271.050 13.050 271.350 ;
        RECT 15.750 270.450 22.500 271.350 ;
        RECT 5.100 268.050 6.900 269.850 ;
        RECT 15.750 268.050 16.950 270.450 ;
        RECT 5.100 267.000 16.950 268.050 ;
        RECT 18.750 267.750 20.550 269.550 ;
        RECT 21.450 268.950 22.500 270.450 ;
        RECT 23.400 271.050 46.500 271.650 ;
        RECT 23.400 270.450 34.050 271.050 ;
        RECT 23.400 269.850 25.200 270.450 ;
        RECT 31.950 270.150 34.050 270.450 ;
        RECT 36.150 269.250 38.250 269.550 ;
        RECT 44.700 269.250 46.500 271.050 ;
        RECT 47.850 270.000 54.900 271.800 ;
        RECT 21.450 268.050 33.450 268.950 ;
        RECT 2.700 265.200 18.000 266.100 ;
        RECT 2.700 261.600 3.900 265.200 ;
        RECT 6.900 263.700 8.700 264.300 ;
        RECT 6.900 262.500 15.300 263.700 ;
        RECT 13.800 261.600 15.300 262.500 ;
        RECT 2.700 255.750 4.500 261.600 ;
        RECT 8.100 255.750 9.900 261.600 ;
        RECT 13.500 255.750 15.300 261.600 ;
        RECT 16.950 262.050 18.000 265.200 ;
        RECT 19.500 264.300 20.550 267.750 ;
        RECT 27.150 265.350 31.050 267.150 ;
        RECT 28.950 265.050 31.050 265.350 ;
        RECT 32.400 266.550 33.450 268.050 ;
        RECT 34.350 267.450 38.250 269.250 ;
        RECT 47.850 268.350 48.750 270.000 ;
        RECT 55.950 269.100 58.050 273.150 ;
        RECT 39.150 267.300 48.750 268.350 ;
        RECT 49.800 268.050 58.050 269.100 ;
        RECT 39.150 266.550 40.050 267.300 ;
        RECT 32.400 265.200 40.050 266.550 ;
        RECT 49.800 266.250 50.850 268.050 ;
        RECT 40.950 265.200 50.850 266.250 ;
        RECT 54.300 265.200 62.100 267.000 ;
        RECT 22.050 264.300 23.850 264.750 ;
        RECT 40.950 264.300 42.000 265.200 ;
        RECT 19.500 263.850 23.850 264.300 ;
        RECT 19.500 263.100 27.150 263.850 ;
        RECT 22.050 262.950 27.150 263.100 ;
        RECT 16.950 259.950 19.050 262.050 ;
        RECT 19.950 259.950 22.050 262.050 ;
        RECT 22.950 259.950 25.050 262.050 ;
        RECT 26.250 261.600 27.150 262.950 ;
        RECT 35.100 262.500 42.000 264.300 ;
        RECT 42.900 262.500 49.650 264.300 ;
        RECT 54.300 261.600 55.800 265.200 ;
        RECT 63.150 261.600 64.350 276.450 ;
        RECT 26.250 260.250 30.300 261.600 ;
        RECT 31.950 261.300 34.050 261.600 ;
        RECT 17.700 258.600 19.050 259.950 ;
        RECT 20.700 258.600 22.050 259.950 ;
        RECT 23.700 258.600 25.050 259.950 ;
        RECT 28.500 259.800 30.300 260.250 ;
        RECT 31.200 259.500 34.050 261.300 ;
        RECT 36.150 261.300 38.250 261.600 ;
        RECT 36.150 259.500 39.000 261.300 ;
        RECT 17.700 255.750 19.500 258.600 ;
        RECT 20.700 255.750 22.500 258.600 ;
        RECT 23.700 255.750 25.500 258.600 ;
        RECT 26.700 255.750 28.500 258.600 ;
        RECT 31.200 255.750 33.000 259.500 ;
        RECT 34.200 255.750 36.000 258.600 ;
        RECT 37.200 255.750 39.000 259.500 ;
        RECT 40.950 259.500 43.050 261.600 ;
        RECT 43.950 259.500 46.050 261.600 ;
        RECT 46.950 259.500 49.050 261.600 ;
        RECT 51.600 260.400 55.800 261.600 ;
        RECT 40.950 255.750 42.750 259.500 ;
        RECT 43.950 255.750 45.750 259.500 ;
        RECT 46.950 255.750 48.750 259.500 ;
        RECT 51.600 255.750 53.400 260.400 ;
        RECT 57.150 255.750 58.950 261.600 ;
        RECT 62.550 255.750 64.350 261.600 ;
        RECT 66.450 268.950 67.950 281.400 ;
        RECT 77.250 281.100 78.450 281.400 ;
        RECT 82.650 281.400 84.450 287.250 ;
        RECT 85.650 281.400 87.450 287.250 ;
        RECT 82.650 281.100 84.300 281.400 ;
        RECT 77.250 280.200 84.300 281.100 ;
        RECT 77.250 271.950 78.300 280.200 ;
        RECT 83.100 276.150 84.900 277.950 ;
        RECT 79.950 273.150 81.750 274.950 ;
        RECT 82.950 274.050 85.050 276.150 ;
        RECT 92.550 275.400 94.350 287.250 ;
        RECT 95.550 275.400 97.350 287.250 ;
        RECT 111.450 275.400 113.250 287.250 ;
        RECT 115.650 275.400 117.450 287.250 ;
        RECT 119.550 275.400 121.350 287.250 ;
        RECT 123.750 275.400 125.550 287.250 ;
        RECT 139.650 281.400 141.450 287.250 ;
        RECT 142.650 282.000 144.450 287.250 ;
        RECT 86.100 273.150 87.900 274.950 ;
        RECT 76.950 269.850 79.050 271.950 ;
        RECT 79.950 271.050 82.050 273.150 ;
        RECT 85.950 271.050 88.050 273.150 ;
        RECT 95.400 270.150 96.600 275.400 ;
        RECT 111.450 274.350 114.000 275.400 ;
        RECT 110.100 270.150 111.900 271.950 ;
        RECT 66.450 266.850 70.050 268.950 ;
        RECT 66.450 258.600 67.950 266.850 ;
        RECT 77.400 265.650 78.600 269.850 ;
        RECT 91.950 266.850 94.050 268.950 ;
        RECT 94.950 268.050 97.050 270.150 ;
        RECT 109.950 268.050 112.050 270.150 ;
        RECT 77.400 264.000 81.900 265.650 ;
        RECT 92.100 265.050 93.900 266.850 ;
        RECT 66.450 255.750 68.250 258.600 ;
        RECT 69.450 255.750 71.250 258.600 ;
        RECT 80.100 255.750 81.900 264.000 ;
        RECT 85.500 255.750 87.300 264.600 ;
        RECT 95.400 261.600 96.600 268.050 ;
        RECT 112.950 267.150 114.000 274.350 ;
        RECT 123.000 274.350 125.550 275.400 ;
        RECT 140.250 281.100 141.450 281.400 ;
        RECT 145.650 281.400 147.450 287.250 ;
        RECT 148.650 281.400 150.450 287.250 ;
        RECT 152.550 281.400 154.350 287.250 ;
        RECT 155.550 281.400 157.350 287.250 ;
        RECT 158.550 282.000 160.350 287.250 ;
        RECT 145.650 281.100 147.300 281.400 ;
        RECT 140.250 280.200 147.300 281.100 ;
        RECT 155.700 281.100 157.350 281.400 ;
        RECT 161.550 281.400 163.350 287.250 ;
        RECT 161.550 281.100 162.750 281.400 ;
        RECT 155.700 280.200 162.750 281.100 ;
        RECT 116.100 270.150 117.900 271.950 ;
        RECT 119.100 270.150 120.900 271.950 ;
        RECT 115.950 268.050 118.050 270.150 ;
        RECT 118.950 268.050 121.050 270.150 ;
        RECT 123.000 267.150 124.050 274.350 ;
        RECT 140.250 271.950 141.300 280.200 ;
        RECT 146.100 276.150 147.900 277.950 ;
        RECT 155.100 276.150 156.900 277.950 ;
        RECT 142.950 273.150 144.750 274.950 ;
        RECT 145.950 274.050 148.050 276.150 ;
        RECT 149.100 273.150 150.900 274.950 ;
        RECT 152.100 273.150 153.900 274.950 ;
        RECT 154.950 274.050 157.050 276.150 ;
        RECT 158.250 273.150 160.050 274.950 ;
        RECT 125.100 270.150 126.900 271.950 ;
        RECT 124.950 268.050 127.050 270.150 ;
        RECT 139.950 269.850 142.050 271.950 ;
        RECT 142.950 271.050 145.050 273.150 ;
        RECT 148.950 271.050 151.050 273.150 ;
        RECT 151.950 271.050 154.050 273.150 ;
        RECT 157.950 271.050 160.050 273.150 ;
        RECT 161.700 271.950 162.750 280.200 ;
        RECT 175.050 275.400 176.850 287.250 ;
        RECT 178.050 275.400 179.850 287.250 ;
        RECT 181.650 281.400 183.450 287.250 ;
        RECT 184.650 281.400 186.450 287.250 ;
        RECT 193.650 281.400 195.450 287.250 ;
        RECT 196.650 281.400 198.450 287.250 ;
        RECT 199.650 281.400 201.450 287.250 ;
        RECT 160.950 269.850 163.050 271.950 ;
        RECT 175.650 270.150 176.850 275.400 ;
        RECT 112.950 265.050 115.050 267.150 ;
        RECT 121.950 265.050 124.050 267.150 ;
        RECT 92.550 255.750 94.350 261.600 ;
        RECT 95.550 255.750 97.350 261.600 ;
        RECT 112.950 258.600 114.000 265.050 ;
        RECT 123.000 258.600 124.050 265.050 ;
        RECT 140.400 265.650 141.600 269.850 ;
        RECT 161.400 265.650 162.600 269.850 ;
        RECT 140.400 264.000 144.900 265.650 ;
        RECT 109.650 255.750 111.450 258.600 ;
        RECT 112.650 255.750 114.450 258.600 ;
        RECT 115.650 255.750 117.450 258.600 ;
        RECT 119.550 255.750 121.350 258.600 ;
        RECT 122.550 255.750 124.350 258.600 ;
        RECT 125.550 255.750 127.350 258.600 ;
        RECT 143.100 255.750 144.900 264.000 ;
        RECT 148.500 255.750 150.300 264.600 ;
        RECT 152.700 255.750 154.500 264.600 ;
        RECT 158.100 264.000 162.600 265.650 ;
        RECT 175.650 268.050 178.050 270.150 ;
        RECT 178.950 269.850 181.050 271.950 ;
        RECT 179.100 268.050 180.900 269.850 ;
        RECT 158.100 255.750 159.900 264.000 ;
        RECT 175.650 261.600 176.850 268.050 ;
        RECT 182.100 264.300 183.300 281.400 ;
        RECT 197.250 273.150 198.450 281.400 ;
        RECT 208.650 275.400 210.450 287.250 ;
        RECT 211.650 276.300 213.450 287.250 ;
        RECT 214.650 277.200 216.450 287.250 ;
        RECT 217.650 276.300 219.450 287.250 ;
        RECT 211.650 275.400 219.450 276.300 ;
        RECT 225.300 275.400 227.100 287.250 ;
        RECT 229.500 275.400 231.300 287.250 ;
        RECT 232.800 281.400 234.600 287.250 ;
        RECT 242.550 281.400 244.350 287.250 ;
        RECT 245.550 281.400 247.350 287.250 ;
        RECT 248.550 281.400 250.350 287.250 ;
        RECT 259.650 281.400 261.450 287.250 ;
        RECT 262.650 281.400 264.450 287.250 ;
        RECT 265.650 281.400 267.450 287.250 ;
        RECT 272.550 281.400 274.350 287.250 ;
        RECT 275.550 281.400 277.350 287.250 ;
        RECT 278.550 281.400 280.350 287.250 ;
        RECT 287.550 281.400 289.350 287.250 ;
        RECT 290.550 281.400 292.350 287.250 ;
        RECT 293.550 281.400 295.350 287.250 ;
        RECT 185.100 270.150 186.900 271.950 ;
        RECT 184.950 268.050 187.050 270.150 ;
        RECT 193.950 269.850 196.050 271.950 ;
        RECT 196.950 271.050 199.050 273.150 ;
        RECT 194.100 268.050 195.900 269.850 ;
        RECT 178.950 263.100 186.450 264.300 ;
        RECT 197.250 263.700 198.450 271.050 ;
        RECT 199.950 269.850 202.050 271.950 ;
        RECT 209.100 270.150 210.300 275.400 ;
        RECT 224.100 270.150 225.900 271.950 ;
        RECT 229.950 270.150 231.150 275.400 ;
        RECT 232.950 273.150 234.750 274.950 ;
        RECT 245.550 273.150 246.750 281.400 ;
        RECT 263.250 273.150 264.450 281.400 ;
        RECT 275.550 273.150 276.750 281.400 ;
        RECT 290.550 273.150 291.750 281.400 ;
        RECT 299.550 276.300 301.350 287.250 ;
        RECT 302.550 277.200 304.350 287.250 ;
        RECT 305.550 276.300 307.350 287.250 ;
        RECT 299.550 275.400 307.350 276.300 ;
        RECT 308.550 275.400 310.350 287.250 ;
        RECT 318.300 275.400 320.100 287.250 ;
        RECT 322.500 275.400 324.300 287.250 ;
        RECT 325.800 281.400 327.600 287.250 ;
        RECT 336.300 275.400 338.100 287.250 ;
        RECT 340.500 275.400 342.300 287.250 ;
        RECT 343.800 281.400 345.600 287.250 ;
        RECT 353.550 281.400 355.350 287.250 ;
        RECT 356.550 281.400 358.350 287.250 ;
        RECT 359.550 281.400 361.350 287.250 ;
        RECT 352.950 276.450 355.050 277.050 ;
        RECT 350.550 275.550 355.050 276.450 ;
        RECT 232.950 271.050 235.050 273.150 ;
        RECT 200.100 268.050 201.900 269.850 ;
        RECT 208.950 268.050 211.050 270.150 ;
        RECT 178.950 262.500 180.750 263.100 ;
        RECT 175.650 260.100 178.950 261.600 ;
        RECT 177.150 255.750 178.950 260.100 ;
        RECT 180.150 255.750 181.950 261.600 ;
        RECT 184.650 255.750 186.450 263.100 ;
        RECT 194.850 262.800 198.450 263.700 ;
        RECT 194.850 255.750 196.650 262.800 ;
        RECT 209.100 261.600 210.300 268.050 ;
        RECT 211.950 266.850 214.050 268.950 ;
        RECT 215.100 267.150 216.900 268.950 ;
        RECT 212.100 265.050 213.900 266.850 ;
        RECT 214.950 265.050 217.050 267.150 ;
        RECT 217.950 266.850 220.050 268.950 ;
        RECT 223.950 268.050 226.050 270.150 ;
        RECT 226.950 266.850 229.050 268.950 ;
        RECT 229.950 268.050 232.050 270.150 ;
        RECT 241.950 269.850 244.050 271.950 ;
        RECT 244.950 271.050 247.050 273.150 ;
        RECT 242.100 268.050 243.900 269.850 ;
        RECT 218.100 265.050 219.900 266.850 ;
        RECT 227.100 265.050 228.900 266.850 ;
        RECT 230.850 264.750 232.050 268.050 ;
        RECT 231.000 263.700 234.750 264.750 ;
        RECT 199.350 255.750 201.150 261.600 ;
        RECT 209.100 259.950 214.800 261.600 ;
        RECT 209.700 255.750 211.500 258.600 ;
        RECT 213.000 255.750 214.800 259.950 ;
        RECT 217.200 255.750 219.000 261.600 ;
        RECT 224.550 260.700 232.350 262.050 ;
        RECT 224.550 255.750 226.350 260.700 ;
        RECT 227.550 255.750 229.350 259.800 ;
        RECT 230.550 255.750 232.350 260.700 ;
        RECT 233.550 261.600 234.750 263.700 ;
        RECT 245.550 263.700 246.750 271.050 ;
        RECT 247.950 269.850 250.050 271.950 ;
        RECT 259.950 269.850 262.050 271.950 ;
        RECT 262.950 271.050 265.050 273.150 ;
        RECT 248.100 268.050 249.900 269.850 ;
        RECT 260.100 268.050 261.900 269.850 ;
        RECT 263.250 263.700 264.450 271.050 ;
        RECT 265.950 269.850 268.050 271.950 ;
        RECT 271.950 269.850 274.050 271.950 ;
        RECT 274.950 271.050 277.050 273.150 ;
        RECT 266.100 268.050 267.900 269.850 ;
        RECT 272.100 268.050 273.900 269.850 ;
        RECT 245.550 262.800 249.150 263.700 ;
        RECT 233.550 255.750 235.350 261.600 ;
        RECT 242.850 255.750 244.650 261.600 ;
        RECT 247.350 255.750 249.150 262.800 ;
        RECT 260.850 262.800 264.450 263.700 ;
        RECT 275.550 263.700 276.750 271.050 ;
        RECT 277.950 269.850 280.050 271.950 ;
        RECT 286.950 269.850 289.050 271.950 ;
        RECT 289.950 271.050 292.050 273.150 ;
        RECT 278.100 268.050 279.900 269.850 ;
        RECT 287.100 268.050 288.900 269.850 ;
        RECT 290.550 263.700 291.750 271.050 ;
        RECT 292.950 269.850 295.050 271.950 ;
        RECT 308.700 270.150 309.900 275.400 ;
        RECT 317.100 270.150 318.900 271.950 ;
        RECT 322.950 270.150 324.150 275.400 ;
        RECT 325.950 273.150 327.750 274.950 ;
        RECT 325.950 271.050 328.050 273.150 ;
        RECT 335.100 270.150 336.900 271.950 ;
        RECT 340.950 270.150 342.150 275.400 ;
        RECT 343.950 273.150 345.750 274.950 ;
        RECT 343.950 271.050 346.050 273.150 ;
        RECT 293.100 268.050 294.900 269.850 ;
        RECT 298.950 266.850 301.050 268.950 ;
        RECT 302.100 267.150 303.900 268.950 ;
        RECT 299.100 265.050 300.900 266.850 ;
        RECT 301.950 265.050 304.050 267.150 ;
        RECT 304.950 266.850 307.050 268.950 ;
        RECT 307.950 268.050 310.050 270.150 ;
        RECT 316.950 268.050 319.050 270.150 ;
        RECT 305.100 265.050 306.900 266.850 ;
        RECT 275.550 262.800 279.150 263.700 ;
        RECT 290.550 262.800 294.150 263.700 ;
        RECT 260.850 255.750 262.650 262.800 ;
        RECT 265.350 255.750 267.150 261.600 ;
        RECT 272.850 255.750 274.650 261.600 ;
        RECT 277.350 255.750 279.150 262.800 ;
        RECT 287.850 255.750 289.650 261.600 ;
        RECT 292.350 255.750 294.150 262.800 ;
        RECT 308.700 261.600 309.900 268.050 ;
        RECT 319.950 266.850 322.050 268.950 ;
        RECT 322.950 268.050 325.050 270.150 ;
        RECT 334.950 268.050 337.050 270.150 ;
        RECT 320.100 265.050 321.900 266.850 ;
        RECT 323.850 264.750 325.050 268.050 ;
        RECT 337.950 266.850 340.050 268.950 ;
        RECT 340.950 268.050 343.050 270.150 ;
        RECT 338.100 265.050 339.900 266.850 ;
        RECT 341.850 264.750 343.050 268.050 ;
        RECT 343.950 267.450 346.050 268.050 ;
        RECT 350.550 267.450 351.450 275.550 ;
        RECT 352.950 274.950 355.050 275.550 ;
        RECT 356.550 273.150 357.750 281.400 ;
        RECT 364.950 274.950 367.050 277.050 ;
        RECT 370.650 275.400 372.450 287.250 ;
        RECT 373.650 275.400 375.450 287.250 ;
        RECT 382.650 275.400 384.450 287.250 ;
        RECT 385.650 276.300 387.450 287.250 ;
        RECT 388.650 277.200 390.450 287.250 ;
        RECT 391.650 276.300 393.450 287.250 ;
        RECT 385.650 275.400 393.450 276.300 ;
        RECT 399.300 275.400 401.100 287.250 ;
        RECT 403.500 275.400 405.300 287.250 ;
        RECT 406.800 281.400 408.600 287.250 ;
        RECT 420.300 275.400 422.100 287.250 ;
        RECT 424.500 275.400 426.300 287.250 ;
        RECT 427.800 281.400 429.600 287.250 ;
        RECT 436.650 281.400 438.450 287.250 ;
        RECT 439.650 282.000 441.450 287.250 ;
        RECT 437.250 281.100 438.450 281.400 ;
        RECT 442.650 281.400 444.450 287.250 ;
        RECT 445.650 281.400 447.450 287.250 ;
        RECT 454.650 281.400 456.450 287.250 ;
        RECT 457.650 281.400 459.450 287.250 ;
        RECT 460.650 281.400 462.450 287.250 ;
        RECT 467.550 281.400 469.350 287.250 ;
        RECT 470.550 281.400 472.350 287.250 ;
        RECT 473.550 281.400 475.350 287.250 ;
        RECT 482.550 281.400 484.350 287.250 ;
        RECT 485.550 281.400 487.350 287.250 ;
        RECT 488.550 281.400 490.350 287.250 ;
        RECT 442.650 281.100 444.300 281.400 ;
        RECT 437.250 280.200 444.300 281.100 ;
        RECT 352.950 269.850 355.050 271.950 ;
        RECT 355.950 271.050 358.050 273.150 ;
        RECT 353.100 268.050 354.900 269.850 ;
        RECT 343.950 266.550 351.450 267.450 ;
        RECT 343.950 265.950 346.050 266.550 ;
        RECT 324.000 263.700 327.750 264.750 ;
        RECT 342.000 263.700 345.750 264.750 ;
        RECT 300.000 255.750 301.800 261.600 ;
        RECT 304.200 259.950 309.900 261.600 ;
        RECT 317.550 260.700 325.350 262.050 ;
        RECT 304.200 255.750 306.000 259.950 ;
        RECT 307.500 255.750 309.300 258.600 ;
        RECT 317.550 255.750 319.350 260.700 ;
        RECT 320.550 255.750 322.350 259.800 ;
        RECT 323.550 255.750 325.350 260.700 ;
        RECT 326.550 261.600 327.750 263.700 ;
        RECT 326.550 255.750 328.350 261.600 ;
        RECT 335.550 260.700 343.350 262.050 ;
        RECT 335.550 255.750 337.350 260.700 ;
        RECT 338.550 255.750 340.350 259.800 ;
        RECT 341.550 255.750 343.350 260.700 ;
        RECT 344.550 261.600 345.750 263.700 ;
        RECT 356.550 263.700 357.750 271.050 ;
        RECT 358.950 269.850 361.050 271.950 ;
        RECT 359.100 268.050 360.900 269.850 ;
        RECT 365.550 267.450 366.450 274.950 ;
        RECT 371.400 270.150 372.600 275.400 ;
        RECT 376.950 273.450 379.050 274.050 ;
        RECT 376.950 272.550 381.450 273.450 ;
        RECT 376.950 271.950 379.050 272.550 ;
        RECT 370.950 268.050 373.050 270.150 ;
        RECT 367.950 267.450 370.050 268.050 ;
        RECT 365.550 266.550 370.050 267.450 ;
        RECT 367.950 265.950 370.050 266.550 ;
        RECT 356.550 262.800 360.150 263.700 ;
        RECT 344.550 255.750 346.350 261.600 ;
        RECT 353.850 255.750 355.650 261.600 ;
        RECT 358.350 255.750 360.150 262.800 ;
        RECT 371.400 261.600 372.600 268.050 ;
        RECT 373.950 266.850 376.050 268.950 ;
        RECT 374.100 265.050 375.900 266.850 ;
        RECT 380.550 265.050 381.450 272.550 ;
        RECT 383.100 270.150 384.300 275.400 ;
        RECT 394.950 271.950 397.050 274.050 ;
        RECT 382.950 268.050 385.050 270.150 ;
        RECT 379.950 262.950 382.050 265.050 ;
        RECT 383.100 261.600 384.300 268.050 ;
        RECT 385.950 266.850 388.050 268.950 ;
        RECT 389.100 267.150 390.900 268.950 ;
        RECT 386.100 265.050 387.900 266.850 ;
        RECT 388.950 265.050 391.050 267.150 ;
        RECT 391.950 266.850 394.050 268.950 ;
        RECT 392.100 265.050 393.900 266.850 ;
        RECT 395.550 264.450 396.450 271.950 ;
        RECT 398.100 270.150 399.900 271.950 ;
        RECT 403.950 270.150 405.150 275.400 ;
        RECT 406.950 273.150 408.750 274.950 ;
        RECT 406.950 271.050 409.050 273.150 ;
        RECT 419.100 270.150 420.900 271.950 ;
        RECT 424.950 270.150 426.150 275.400 ;
        RECT 430.950 274.950 433.050 277.050 ;
        RECT 427.950 273.150 429.750 274.950 ;
        RECT 427.950 271.050 430.050 273.150 ;
        RECT 397.950 268.050 400.050 270.150 ;
        RECT 400.950 266.850 403.050 268.950 ;
        RECT 403.950 268.050 406.050 270.150 ;
        RECT 418.950 268.050 421.050 270.150 ;
        RECT 401.100 265.050 402.900 266.850 ;
        RECT 397.950 264.450 400.050 265.050 ;
        RECT 404.850 264.750 406.050 268.050 ;
        RECT 421.950 266.850 424.050 268.950 ;
        RECT 424.950 268.050 427.050 270.150 ;
        RECT 422.100 265.050 423.900 266.850 ;
        RECT 425.850 264.750 427.050 268.050 ;
        RECT 427.950 267.450 430.050 268.050 ;
        RECT 431.550 267.450 432.450 274.950 ;
        RECT 437.250 271.950 438.300 280.200 ;
        RECT 443.100 276.150 444.900 277.950 ;
        RECT 439.950 273.150 441.750 274.950 ;
        RECT 442.950 274.050 445.050 276.150 ;
        RECT 446.100 273.150 447.900 274.950 ;
        RECT 458.250 273.150 459.450 281.400 ;
        RECT 466.950 276.450 469.050 277.050 ;
        RECT 464.550 275.550 469.050 276.450 ;
        RECT 436.950 269.850 439.050 271.950 ;
        RECT 439.950 271.050 442.050 273.150 ;
        RECT 445.950 271.050 448.050 273.150 ;
        RECT 454.950 269.850 457.050 271.950 ;
        RECT 457.950 271.050 460.050 273.150 ;
        RECT 427.950 266.550 432.450 267.450 ;
        RECT 427.950 265.950 430.050 266.550 ;
        RECT 437.400 265.650 438.600 269.850 ;
        RECT 455.100 268.050 456.900 269.850 ;
        RECT 395.550 263.550 400.050 264.450 ;
        RECT 405.000 263.700 408.750 264.750 ;
        RECT 426.000 263.700 429.750 264.750 ;
        RECT 437.400 264.000 441.900 265.650 ;
        RECT 397.950 262.950 400.050 263.550 ;
        RECT 370.650 255.750 372.450 261.600 ;
        RECT 373.650 255.750 375.450 261.600 ;
        RECT 383.100 259.950 388.800 261.600 ;
        RECT 383.700 255.750 385.500 258.600 ;
        RECT 387.000 255.750 388.800 259.950 ;
        RECT 391.200 255.750 393.000 261.600 ;
        RECT 398.550 260.700 406.350 262.050 ;
        RECT 398.550 255.750 400.350 260.700 ;
        RECT 401.550 255.750 403.350 259.800 ;
        RECT 404.550 255.750 406.350 260.700 ;
        RECT 407.550 261.600 408.750 263.700 ;
        RECT 407.550 255.750 409.350 261.600 ;
        RECT 419.550 260.700 427.350 262.050 ;
        RECT 419.550 255.750 421.350 260.700 ;
        RECT 422.550 255.750 424.350 259.800 ;
        RECT 425.550 255.750 427.350 260.700 ;
        RECT 428.550 261.600 429.750 263.700 ;
        RECT 428.550 255.750 430.350 261.600 ;
        RECT 440.100 255.750 441.900 264.000 ;
        RECT 445.500 255.750 447.300 264.600 ;
        RECT 458.250 263.700 459.450 271.050 ;
        RECT 460.950 269.850 463.050 271.950 ;
        RECT 461.100 268.050 462.900 269.850 ;
        RECT 464.550 265.050 465.450 275.550 ;
        RECT 466.950 274.950 469.050 275.550 ;
        RECT 470.550 273.150 471.750 281.400 ;
        RECT 485.550 273.150 486.750 281.400 ;
        RECT 490.950 274.950 493.050 277.050 ;
        RECT 494.550 276.600 496.350 287.250 ;
        RECT 497.550 277.500 499.350 287.250 ;
        RECT 500.550 286.500 508.350 287.250 ;
        RECT 500.550 276.600 502.350 286.500 ;
        RECT 494.550 275.700 502.350 276.600 ;
        RECT 503.550 275.400 505.350 285.600 ;
        RECT 506.550 275.400 508.350 286.500 ;
        RECT 518.550 276.600 520.350 287.250 ;
        RECT 521.550 277.500 523.350 287.250 ;
        RECT 524.550 286.500 532.350 287.250 ;
        RECT 524.550 276.600 526.350 286.500 ;
        RECT 518.550 275.700 526.350 276.600 ;
        RECT 527.550 275.400 529.350 285.600 ;
        RECT 530.550 275.400 532.350 286.500 ;
        RECT 538.650 281.400 540.450 287.250 ;
        RECT 541.650 281.400 543.450 287.250 ;
        RECT 550.650 286.500 558.450 287.250 ;
        RECT 466.950 269.850 469.050 271.950 ;
        RECT 469.950 271.050 472.050 273.150 ;
        RECT 467.100 268.050 468.900 269.850 ;
        RECT 455.850 262.800 459.450 263.700 ;
        RECT 463.950 262.950 466.050 265.050 ;
        RECT 470.550 263.700 471.750 271.050 ;
        RECT 472.950 269.850 475.050 271.950 ;
        RECT 481.950 269.850 484.050 271.950 ;
        RECT 484.950 271.050 487.050 273.150 ;
        RECT 473.100 268.050 474.900 269.850 ;
        RECT 482.100 268.050 483.900 269.850 ;
        RECT 485.550 263.700 486.750 271.050 ;
        RECT 487.950 269.850 490.050 271.950 ;
        RECT 488.100 268.050 489.900 269.850 ;
        RECT 491.550 265.050 492.450 274.950 ;
        RECT 503.400 274.500 505.200 275.400 ;
        RECT 527.400 274.500 529.200 275.400 ;
        RECT 501.150 273.600 505.200 274.500 ;
        RECT 525.150 273.600 529.200 274.500 ;
        RECT 494.250 270.150 496.050 271.950 ;
        RECT 501.150 270.150 502.050 273.600 ;
        RECT 506.100 270.150 507.900 271.950 ;
        RECT 518.250 270.150 520.050 271.950 ;
        RECT 525.150 270.150 526.050 273.600 ;
        RECT 530.100 270.150 531.900 271.950 ;
        RECT 493.950 268.050 496.050 270.150 ;
        RECT 496.950 266.850 499.050 268.950 ;
        RECT 497.250 265.050 499.050 266.850 ;
        RECT 499.950 268.050 502.050 270.150 ;
        RECT 470.550 262.800 474.150 263.700 ;
        RECT 485.550 262.800 489.150 263.700 ;
        RECT 490.950 262.950 493.050 265.050 ;
        RECT 455.850 255.750 457.650 262.800 ;
        RECT 460.350 255.750 462.150 261.600 ;
        RECT 467.850 255.750 469.650 261.600 ;
        RECT 472.350 255.750 474.150 262.800 ;
        RECT 482.850 255.750 484.650 261.600 ;
        RECT 487.350 255.750 489.150 262.800 ;
        RECT 499.950 261.600 501.000 268.050 ;
        RECT 502.950 266.850 505.050 268.950 ;
        RECT 505.950 268.050 508.050 270.150 ;
        RECT 517.950 268.050 520.050 270.150 ;
        RECT 520.950 266.850 523.050 268.950 ;
        RECT 502.950 265.050 504.750 266.850 ;
        RECT 521.250 265.050 523.050 266.850 ;
        RECT 523.950 268.050 526.050 270.150 ;
        RECT 517.950 264.450 520.050 265.050 ;
        RECT 515.550 263.550 520.050 264.450 ;
        RECT 495.000 255.750 496.800 261.600 ;
        RECT 499.200 255.750 501.000 261.600 ;
        RECT 503.400 255.750 505.200 261.600 ;
        RECT 508.950 261.450 511.050 262.050 ;
        RECT 515.550 261.450 516.450 263.550 ;
        RECT 517.950 262.950 520.050 263.550 ;
        RECT 523.950 261.600 525.000 268.050 ;
        RECT 526.950 266.850 529.050 268.950 ;
        RECT 529.950 268.050 532.050 270.150 ;
        RECT 539.400 268.950 540.600 281.400 ;
        RECT 550.650 275.400 552.450 286.500 ;
        RECT 553.650 275.400 555.450 285.600 ;
        RECT 556.650 276.600 558.450 286.500 ;
        RECT 559.650 277.500 561.450 287.250 ;
        RECT 562.650 276.600 564.450 287.250 ;
        RECT 556.650 275.700 564.450 276.600 ;
        RECT 569.550 276.300 571.350 287.250 ;
        RECT 572.550 277.200 574.350 287.250 ;
        RECT 575.550 276.300 577.350 287.250 ;
        RECT 569.550 275.400 577.350 276.300 ;
        RECT 578.550 275.400 580.350 287.250 ;
        RECT 586.650 281.400 588.450 287.250 ;
        RECT 589.650 281.400 591.450 287.250 ;
        RECT 553.800 274.500 555.600 275.400 ;
        RECT 553.800 273.600 557.850 274.500 ;
        RECT 551.100 270.150 552.900 271.950 ;
        RECT 556.950 270.150 557.850 273.600 ;
        RECT 562.950 270.150 564.750 271.950 ;
        RECT 578.700 270.150 579.900 275.400 ;
        RECT 538.950 266.850 541.050 268.950 ;
        RECT 542.100 267.150 543.900 268.950 ;
        RECT 550.950 268.050 553.050 270.150 ;
        RECT 526.950 265.050 528.750 266.850 ;
        RECT 508.950 260.550 516.450 261.450 ;
        RECT 508.950 259.950 511.050 260.550 ;
        RECT 519.000 255.750 520.800 261.600 ;
        RECT 523.200 255.750 525.000 261.600 ;
        RECT 527.400 255.750 529.200 261.600 ;
        RECT 539.400 258.600 540.600 266.850 ;
        RECT 541.950 265.050 544.050 267.150 ;
        RECT 553.950 266.850 556.050 268.950 ;
        RECT 556.950 268.050 559.050 270.150 ;
        RECT 554.250 265.050 556.050 266.850 ;
        RECT 550.950 264.450 553.050 265.050 ;
        RECT 548.550 263.550 553.050 264.450 ;
        RECT 541.950 261.450 544.050 262.050 ;
        RECT 548.550 261.450 549.450 263.550 ;
        RECT 550.950 262.950 553.050 263.550 ;
        RECT 558.000 261.600 559.050 268.050 ;
        RECT 559.950 266.850 562.050 268.950 ;
        RECT 562.950 268.050 565.050 270.150 ;
        RECT 559.950 265.050 561.750 266.850 ;
        RECT 565.950 265.950 568.050 268.050 ;
        RECT 568.950 266.850 571.050 268.950 ;
        RECT 572.100 267.150 573.900 268.950 ;
        RECT 562.950 264.450 565.050 265.050 ;
        RECT 566.550 264.450 567.450 265.950 ;
        RECT 569.100 265.050 570.900 266.850 ;
        RECT 571.950 265.050 574.050 267.150 ;
        RECT 574.950 266.850 577.050 268.950 ;
        RECT 577.950 268.050 580.050 270.150 ;
        RECT 587.400 268.950 588.600 281.400 ;
        RECT 594.300 275.400 596.100 287.250 ;
        RECT 598.500 275.400 600.300 287.250 ;
        RECT 601.800 281.400 603.600 287.250 ;
        RECT 608.550 281.400 610.350 287.250 ;
        RECT 611.550 281.400 613.350 287.250 ;
        RECT 617.550 281.400 619.350 287.250 ;
        RECT 620.550 281.400 622.350 287.250 ;
        RECT 623.550 281.400 625.350 287.250 ;
        RECT 629.550 281.400 631.350 287.250 ;
        RECT 632.550 281.400 634.350 287.250 ;
        RECT 635.550 281.400 637.350 287.250 ;
        RECT 593.100 270.150 594.900 271.950 ;
        RECT 598.950 270.150 600.150 275.400 ;
        RECT 601.950 273.150 603.750 274.950 ;
        RECT 607.950 273.450 610.050 274.050 ;
        RECT 601.950 271.050 604.050 273.150 ;
        RECT 605.550 272.550 610.050 273.450 ;
        RECT 575.100 265.050 576.900 266.850 ;
        RECT 562.950 263.550 567.450 264.450 ;
        RECT 562.950 262.950 565.050 263.550 ;
        RECT 578.700 261.600 579.900 268.050 ;
        RECT 586.950 266.850 589.050 268.950 ;
        RECT 590.100 267.150 591.900 268.950 ;
        RECT 592.950 268.050 595.050 270.150 ;
        RECT 541.950 260.550 549.450 261.450 ;
        RECT 541.950 259.950 544.050 260.550 ;
        RECT 538.650 255.750 540.450 258.600 ;
        RECT 541.650 255.750 543.450 258.600 ;
        RECT 553.800 255.750 555.600 261.600 ;
        RECT 558.000 255.750 559.800 261.600 ;
        RECT 562.200 255.750 564.000 261.600 ;
        RECT 570.000 255.750 571.800 261.600 ;
        RECT 574.200 259.950 579.900 261.600 ;
        RECT 574.200 255.750 576.000 259.950 ;
        RECT 587.400 258.600 588.600 266.850 ;
        RECT 589.950 265.050 592.050 267.150 ;
        RECT 595.950 266.850 598.050 268.950 ;
        RECT 598.950 268.050 601.050 270.150 ;
        RECT 596.100 265.050 597.900 266.850 ;
        RECT 599.850 264.750 601.050 268.050 ;
        RECT 601.950 267.450 604.050 268.050 ;
        RECT 605.550 267.450 606.450 272.550 ;
        RECT 607.950 271.950 610.050 272.550 ;
        RECT 611.400 268.950 612.600 281.400 ;
        RECT 620.550 273.150 621.750 281.400 ;
        RECT 632.550 273.150 633.750 281.400 ;
        RECT 637.950 277.950 640.050 280.050 ;
        RECT 616.950 269.850 619.050 271.950 ;
        RECT 619.950 271.050 622.050 273.150 ;
        RECT 601.950 266.550 606.450 267.450 ;
        RECT 608.100 267.150 609.900 268.950 ;
        RECT 601.950 265.950 604.050 266.550 ;
        RECT 607.950 265.050 610.050 267.150 ;
        RECT 610.950 266.850 613.050 268.950 ;
        RECT 617.100 268.050 618.900 269.850 ;
        RECT 600.000 263.700 603.750 264.750 ;
        RECT 593.550 260.700 601.350 262.050 ;
        RECT 577.500 255.750 579.300 258.600 ;
        RECT 586.650 255.750 588.450 258.600 ;
        RECT 589.650 255.750 591.450 258.600 ;
        RECT 593.550 255.750 595.350 260.700 ;
        RECT 596.550 255.750 598.350 259.800 ;
        RECT 599.550 255.750 601.350 260.700 ;
        RECT 602.550 261.600 603.750 263.700 ;
        RECT 602.550 255.750 604.350 261.600 ;
        RECT 611.400 258.600 612.600 266.850 ;
        RECT 620.550 263.700 621.750 271.050 ;
        RECT 622.950 269.850 625.050 271.950 ;
        RECT 628.950 269.850 631.050 271.950 ;
        RECT 631.950 271.050 634.050 273.150 ;
        RECT 623.100 268.050 624.900 269.850 ;
        RECT 629.100 268.050 630.900 269.850 ;
        RECT 632.550 263.700 633.750 271.050 ;
        RECT 634.950 269.850 637.050 271.950 ;
        RECT 635.100 268.050 636.900 269.850 ;
        RECT 620.550 262.800 624.150 263.700 ;
        RECT 632.550 262.800 636.150 263.700 ;
        RECT 608.550 255.750 610.350 258.600 ;
        RECT 611.550 255.750 613.350 258.600 ;
        RECT 617.850 255.750 619.650 261.600 ;
        RECT 622.350 255.750 624.150 262.800 ;
        RECT 629.850 255.750 631.650 261.600 ;
        RECT 634.350 255.750 636.150 262.800 ;
        RECT 638.550 261.450 639.450 277.950 ;
        RECT 649.650 275.400 651.450 287.250 ;
        RECT 652.650 276.300 654.450 287.250 ;
        RECT 655.650 277.200 657.450 287.250 ;
        RECT 658.650 276.300 660.450 287.250 ;
        RECT 652.650 275.400 660.450 276.300 ;
        RECT 667.050 275.400 668.850 287.250 ;
        RECT 670.050 275.400 671.850 287.250 ;
        RECT 673.650 281.400 675.450 287.250 ;
        RECT 676.650 281.400 678.450 287.250 ;
        RECT 686.550 281.400 688.350 287.250 ;
        RECT 689.550 281.400 691.350 287.250 ;
        RECT 692.550 282.000 694.350 287.250 ;
        RECT 650.100 270.150 651.300 275.400 ;
        RECT 667.650 270.150 668.850 275.400 ;
        RECT 649.950 268.050 652.050 270.150 ;
        RECT 646.950 261.450 649.050 262.050 ;
        RECT 638.550 260.550 649.050 261.450 ;
        RECT 646.950 259.950 649.050 260.550 ;
        RECT 650.100 261.600 651.300 268.050 ;
        RECT 652.950 266.850 655.050 268.950 ;
        RECT 656.100 267.150 657.900 268.950 ;
        RECT 653.100 265.050 654.900 266.850 ;
        RECT 655.950 265.050 658.050 267.150 ;
        RECT 658.950 266.850 661.050 268.950 ;
        RECT 667.650 268.050 670.050 270.150 ;
        RECT 670.950 269.850 673.050 271.950 ;
        RECT 671.100 268.050 672.900 269.850 ;
        RECT 659.100 265.050 660.900 266.850 ;
        RECT 667.650 261.600 668.850 268.050 ;
        RECT 674.100 264.300 675.300 281.400 ;
        RECT 689.700 281.100 691.350 281.400 ;
        RECT 695.550 281.400 697.350 287.250 ;
        RECT 701.550 281.400 703.350 287.250 ;
        RECT 704.550 281.400 706.350 287.250 ;
        RECT 716.550 281.400 718.350 287.250 ;
        RECT 719.550 281.400 721.350 287.250 ;
        RECT 722.550 282.000 724.350 287.250 ;
        RECT 695.550 281.100 696.750 281.400 ;
        RECT 689.700 280.200 696.750 281.100 ;
        RECT 689.100 276.150 690.900 277.950 ;
        RECT 682.950 271.950 685.050 274.050 ;
        RECT 686.100 273.150 687.900 274.950 ;
        RECT 688.950 274.050 691.050 276.150 ;
        RECT 692.250 273.150 694.050 274.950 ;
        RECT 677.100 270.150 678.900 271.950 ;
        RECT 676.950 268.050 679.050 270.150 ;
        RECT 683.550 267.450 684.450 271.950 ;
        RECT 685.950 271.050 688.050 273.150 ;
        RECT 691.950 271.050 694.050 273.150 ;
        RECT 695.700 271.950 696.750 280.200 ;
        RECT 694.950 269.850 697.050 271.950 ;
        RECT 685.950 267.450 688.050 268.050 ;
        RECT 683.550 266.550 688.050 267.450 ;
        RECT 685.950 265.950 688.050 266.550 ;
        RECT 695.400 265.650 696.600 269.850 ;
        RECT 704.400 268.950 705.600 281.400 ;
        RECT 719.700 281.100 721.350 281.400 ;
        RECT 725.550 281.400 727.350 287.250 ;
        RECT 736.650 281.400 738.450 287.250 ;
        RECT 739.650 281.400 741.450 287.250 ;
        RECT 742.650 281.400 744.450 287.250 ;
        RECT 725.550 281.100 726.750 281.400 ;
        RECT 719.700 280.200 726.750 281.100 ;
        RECT 719.100 276.150 720.900 277.950 ;
        RECT 716.100 273.150 717.900 274.950 ;
        RECT 718.950 274.050 721.050 276.150 ;
        RECT 722.250 273.150 724.050 274.950 ;
        RECT 715.950 271.050 718.050 273.150 ;
        RECT 721.950 271.050 724.050 273.150 ;
        RECT 725.700 271.950 726.750 280.200 ;
        RECT 736.950 276.450 739.050 277.050 ;
        RECT 734.550 275.550 739.050 276.450 ;
        RECT 724.950 269.850 727.050 271.950 ;
        RECT 701.100 267.150 702.900 268.950 ;
        RECT 670.950 263.100 678.450 264.300 ;
        RECT 670.950 262.500 672.750 263.100 ;
        RECT 650.100 259.950 655.800 261.600 ;
        RECT 650.700 255.750 652.500 258.600 ;
        RECT 654.000 255.750 655.800 259.950 ;
        RECT 658.200 255.750 660.000 261.600 ;
        RECT 667.650 260.100 670.950 261.600 ;
        RECT 669.150 255.750 670.950 260.100 ;
        RECT 672.150 255.750 673.950 261.600 ;
        RECT 676.650 255.750 678.450 263.100 ;
        RECT 686.700 255.750 688.500 264.600 ;
        RECT 692.100 264.000 696.600 265.650 ;
        RECT 700.950 265.050 703.050 267.150 ;
        RECT 703.950 266.850 706.050 268.950 ;
        RECT 692.100 255.750 693.900 264.000 ;
        RECT 704.400 258.600 705.600 266.850 ;
        RECT 725.400 265.650 726.600 269.850 ;
        RECT 701.550 255.750 703.350 258.600 ;
        RECT 704.550 255.750 706.350 258.600 ;
        RECT 716.700 255.750 718.500 264.600 ;
        RECT 722.100 264.000 726.600 265.650 ;
        RECT 727.950 264.450 730.050 265.050 ;
        RECT 734.550 264.450 735.450 275.550 ;
        RECT 736.950 274.950 739.050 275.550 ;
        RECT 740.250 273.150 741.450 281.400 ;
        RECT 751.650 275.400 753.450 287.250 ;
        RECT 754.650 276.300 756.450 287.250 ;
        RECT 757.650 277.200 759.450 287.250 ;
        RECT 760.650 276.300 762.450 287.250 ;
        RECT 770.400 281.400 772.200 287.250 ;
        RECT 754.650 275.400 762.450 276.300 ;
        RECT 773.700 275.400 775.500 287.250 ;
        RECT 777.900 275.400 779.700 287.250 ;
        RECT 782.700 281.400 784.500 287.250 ;
        RECT 785.700 281.400 787.500 287.250 ;
        RECT 788.700 281.400 790.500 287.250 ;
        RECT 785.700 280.500 786.750 281.400 ;
        RECT 782.700 279.600 786.750 280.500 ;
        RECT 736.950 269.850 739.050 271.950 ;
        RECT 739.950 271.050 742.050 273.150 ;
        RECT 737.100 268.050 738.900 269.850 ;
        RECT 722.100 255.750 723.900 264.000 ;
        RECT 727.950 263.550 735.450 264.450 ;
        RECT 740.250 263.700 741.450 271.050 ;
        RECT 742.950 269.850 745.050 271.950 ;
        RECT 752.100 270.150 753.300 275.400 ;
        RECT 770.250 273.150 772.050 274.950 ;
        RECT 769.950 271.050 772.050 273.150 ;
        RECT 773.850 270.150 775.050 275.400 ;
        RECT 779.100 270.150 780.900 271.950 ;
        RECT 743.100 268.050 744.900 269.850 ;
        RECT 751.950 268.050 754.050 270.150 ;
        RECT 727.950 262.950 730.050 263.550 ;
        RECT 737.850 262.800 741.450 263.700 ;
        RECT 737.850 255.750 739.650 262.800 ;
        RECT 752.100 261.600 753.300 268.050 ;
        RECT 754.950 266.850 757.050 268.950 ;
        RECT 758.100 267.150 759.900 268.950 ;
        RECT 755.100 265.050 756.900 266.850 ;
        RECT 757.950 265.050 760.050 267.150 ;
        RECT 760.950 266.850 763.050 268.950 ;
        RECT 772.950 268.050 775.050 270.150 ;
        RECT 761.100 265.050 762.900 266.850 ;
        RECT 772.950 264.750 774.150 268.050 ;
        RECT 775.950 266.850 778.050 268.950 ;
        RECT 778.950 268.050 781.050 270.150 ;
        RECT 776.100 265.050 777.900 266.850 ;
        RECT 782.700 266.100 783.900 279.600 ;
        RECT 791.700 278.700 793.500 287.250 ;
        RECT 794.700 283.950 796.500 287.250 ;
        RECT 797.850 284.400 800.250 287.250 ;
        RECT 801.150 284.400 803.250 287.250 ;
        RECT 804.300 284.400 806.250 287.250 ;
        RECT 797.850 283.050 799.050 284.400 ;
        RECT 801.150 283.050 802.050 284.400 ;
        RECT 804.300 283.050 805.500 284.400 ;
        RECT 796.950 280.950 799.050 283.050 ;
        RECT 799.950 280.950 802.050 283.050 ;
        RECT 802.950 281.400 805.500 283.050 ;
        RECT 807.450 281.400 809.250 287.250 ;
        RECT 811.200 281.400 813.000 287.250 ;
        RECT 814.200 281.400 816.000 287.250 ;
        RECT 802.950 280.950 805.050 281.400 ;
        RECT 811.650 280.500 813.000 281.400 ;
        RECT 817.200 280.500 819.000 287.250 ;
        RECT 820.950 284.400 822.750 287.250 ;
        RECT 811.650 278.850 814.050 280.500 ;
        RECT 787.200 277.650 804.900 278.700 ;
        RECT 811.950 278.400 814.050 278.850 ;
        RECT 816.000 280.200 819.000 280.500 ;
        RECT 816.000 278.400 819.900 280.200 ;
        RECT 787.200 276.900 789.000 277.650 ;
        RECT 799.950 276.150 802.050 276.750 ;
        RECT 790.500 274.950 802.050 276.150 ;
        RECT 802.950 276.600 804.900 277.650 ;
        RECT 821.100 277.350 822.450 284.400 ;
        RECT 823.950 280.950 825.750 287.250 ;
        RECT 826.950 284.400 828.750 287.250 ;
        RECT 827.100 283.200 828.600 284.400 ;
        RECT 827.100 281.100 829.200 283.200 ;
        RECT 830.700 281.400 832.500 287.250 ;
        RECT 823.950 280.050 826.050 280.950 ;
        RECT 833.700 280.500 835.500 287.250 ;
        RECT 836.700 281.400 838.500 287.250 ;
        RECT 839.700 281.400 841.500 287.250 ;
        RECT 842.700 281.400 844.500 287.250 ;
        RECT 846.450 281.400 848.250 287.250 ;
        RECT 849.450 281.400 851.250 287.250 ;
        RECT 830.850 280.050 832.650 280.500 ;
        RECT 823.950 278.850 832.650 280.050 ;
        RECT 833.700 279.300 839.400 280.500 ;
        RECT 830.850 278.700 832.650 278.850 ;
        RECT 837.600 278.700 839.400 279.300 ;
        RECT 840.300 277.350 841.500 281.400 ;
        RECT 820.950 276.600 823.050 277.350 ;
        RECT 802.950 275.250 823.050 276.600 ;
        RECT 826.950 276.450 844.350 277.350 ;
        RECT 826.950 275.250 829.050 276.450 ;
        RECT 790.500 274.350 792.300 274.950 ;
        RECT 799.950 274.650 802.050 274.950 ;
        RECT 829.950 274.350 842.250 275.550 ;
        RECT 802.950 273.450 831.000 274.350 ;
        RECT 840.450 273.750 842.250 274.350 ;
        RECT 791.250 273.150 831.000 273.450 ;
        RECT 790.950 272.550 804.900 273.150 ;
        RECT 784.950 269.850 787.050 271.950 ;
        RECT 790.950 271.350 794.850 272.550 ;
        RECT 811.950 271.650 826.500 272.250 ;
        RECT 790.950 271.050 793.050 271.350 ;
        RECT 795.750 270.450 802.500 271.350 ;
        RECT 785.100 268.050 786.900 269.850 ;
        RECT 795.750 268.050 796.950 270.450 ;
        RECT 785.100 267.000 796.950 268.050 ;
        RECT 798.750 267.750 800.550 269.550 ;
        RECT 801.450 268.950 802.500 270.450 ;
        RECT 803.400 271.050 826.500 271.650 ;
        RECT 803.400 270.450 814.050 271.050 ;
        RECT 803.400 269.850 805.200 270.450 ;
        RECT 811.950 270.150 814.050 270.450 ;
        RECT 816.150 269.250 818.250 269.550 ;
        RECT 824.700 269.250 826.500 271.050 ;
        RECT 827.850 270.000 834.900 271.800 ;
        RECT 801.450 268.050 813.450 268.950 ;
        RECT 782.700 265.200 798.000 266.100 ;
        RECT 770.250 263.700 774.000 264.750 ;
        RECT 770.250 261.600 771.450 263.700 ;
        RECT 742.350 255.750 744.150 261.600 ;
        RECT 752.100 259.950 757.800 261.600 ;
        RECT 752.700 255.750 754.500 258.600 ;
        RECT 756.000 255.750 757.800 259.950 ;
        RECT 760.200 255.750 762.000 261.600 ;
        RECT 769.650 255.750 771.450 261.600 ;
        RECT 772.650 260.700 780.450 262.050 ;
        RECT 772.650 255.750 774.450 260.700 ;
        RECT 775.650 255.750 777.450 259.800 ;
        RECT 778.650 255.750 780.450 260.700 ;
        RECT 782.700 261.600 783.900 265.200 ;
        RECT 786.900 263.700 788.700 264.300 ;
        RECT 786.900 262.500 795.300 263.700 ;
        RECT 793.800 261.600 795.300 262.500 ;
        RECT 782.700 255.750 784.500 261.600 ;
        RECT 788.100 255.750 789.900 261.600 ;
        RECT 793.500 255.750 795.300 261.600 ;
        RECT 796.950 262.050 798.000 265.200 ;
        RECT 799.500 264.300 800.550 267.750 ;
        RECT 807.150 265.350 811.050 267.150 ;
        RECT 808.950 265.050 811.050 265.350 ;
        RECT 812.400 266.550 813.450 268.050 ;
        RECT 814.350 267.450 818.250 269.250 ;
        RECT 827.850 268.350 828.750 270.000 ;
        RECT 835.950 269.100 838.050 273.150 ;
        RECT 819.150 267.300 828.750 268.350 ;
        RECT 829.800 268.050 838.050 269.100 ;
        RECT 819.150 266.550 820.050 267.300 ;
        RECT 812.400 265.200 820.050 266.550 ;
        RECT 829.800 266.250 830.850 268.050 ;
        RECT 820.950 265.200 830.850 266.250 ;
        RECT 834.300 265.200 842.100 267.000 ;
        RECT 802.050 264.300 803.850 264.750 ;
        RECT 820.950 264.300 822.000 265.200 ;
        RECT 799.500 263.850 803.850 264.300 ;
        RECT 799.500 263.100 807.150 263.850 ;
        RECT 802.050 262.950 807.150 263.100 ;
        RECT 796.950 259.950 799.050 262.050 ;
        RECT 799.950 259.950 802.050 262.050 ;
        RECT 802.950 259.950 805.050 262.050 ;
        RECT 806.250 261.600 807.150 262.950 ;
        RECT 815.100 262.500 822.000 264.300 ;
        RECT 822.900 262.500 829.650 264.300 ;
        RECT 834.300 261.600 835.800 265.200 ;
        RECT 843.150 261.600 844.350 276.450 ;
        RECT 806.250 260.250 810.300 261.600 ;
        RECT 811.950 261.300 814.050 261.600 ;
        RECT 797.700 258.600 799.050 259.950 ;
        RECT 800.700 258.600 802.050 259.950 ;
        RECT 803.700 258.600 805.050 259.950 ;
        RECT 808.500 259.800 810.300 260.250 ;
        RECT 811.200 259.500 814.050 261.300 ;
        RECT 816.150 261.300 818.250 261.600 ;
        RECT 816.150 259.500 819.000 261.300 ;
        RECT 797.700 255.750 799.500 258.600 ;
        RECT 800.700 255.750 802.500 258.600 ;
        RECT 803.700 255.750 805.500 258.600 ;
        RECT 806.700 255.750 808.500 258.600 ;
        RECT 811.200 255.750 813.000 259.500 ;
        RECT 814.200 255.750 816.000 258.600 ;
        RECT 817.200 255.750 819.000 259.500 ;
        RECT 820.950 259.500 823.050 261.600 ;
        RECT 823.950 259.500 826.050 261.600 ;
        RECT 826.950 259.500 829.050 261.600 ;
        RECT 831.600 260.400 835.800 261.600 ;
        RECT 820.950 255.750 822.750 259.500 ;
        RECT 823.950 255.750 825.750 259.500 ;
        RECT 826.950 255.750 828.750 259.500 ;
        RECT 831.600 255.750 833.400 260.400 ;
        RECT 837.150 255.750 838.950 261.600 ;
        RECT 842.550 255.750 844.350 261.600 ;
        RECT 846.450 268.950 847.950 281.400 ;
        RECT 846.450 266.850 850.050 268.950 ;
        RECT 846.450 258.600 847.950 266.850 ;
        RECT 846.450 255.750 848.250 258.600 ;
        RECT 849.450 255.750 851.250 258.600 ;
        RECT 7.650 245.400 9.450 251.250 ;
        RECT 10.650 245.400 12.450 251.250 ;
        RECT 20.550 246.300 22.350 251.250 ;
        RECT 23.550 247.200 25.350 251.250 ;
        RECT 26.550 246.300 28.350 251.250 ;
        RECT 8.400 238.950 9.600 245.400 ;
        RECT 20.550 244.950 28.350 246.300 ;
        RECT 29.550 245.400 31.350 251.250 ;
        RECT 38.550 246.300 40.350 251.250 ;
        RECT 41.550 247.200 43.350 251.250 ;
        RECT 44.550 246.300 46.350 251.250 ;
        RECT 29.550 243.300 30.750 245.400 ;
        RECT 38.550 244.950 46.350 246.300 ;
        RECT 47.550 245.400 49.350 251.250 ;
        RECT 55.650 245.400 57.450 251.250 ;
        RECT 47.550 243.300 48.750 245.400 ;
        RECT 27.000 242.250 30.750 243.300 ;
        RECT 45.000 242.250 48.750 243.300 ;
        RECT 56.250 243.300 57.450 245.400 ;
        RECT 58.650 246.300 60.450 251.250 ;
        RECT 61.650 247.200 63.450 251.250 ;
        RECT 64.650 246.300 66.450 251.250 ;
        RECT 58.650 244.950 66.450 246.300 ;
        RECT 56.250 242.250 60.000 243.300 ;
        RECT 11.100 240.150 12.900 241.950 ;
        RECT 23.100 240.150 24.900 241.950 ;
        RECT 7.950 236.850 10.050 238.950 ;
        RECT 10.950 238.050 13.050 240.150 ;
        RECT 19.950 236.850 22.050 238.950 ;
        RECT 22.950 238.050 25.050 240.150 ;
        RECT 26.850 238.950 28.050 242.250 ;
        RECT 41.100 240.150 42.900 241.950 ;
        RECT 25.950 236.850 28.050 238.950 ;
        RECT 37.950 236.850 40.050 238.950 ;
        RECT 40.950 238.050 43.050 240.150 ;
        RECT 44.850 238.950 46.050 242.250 ;
        RECT 43.950 236.850 46.050 238.950 ;
        RECT 58.950 238.950 60.150 242.250 ;
        RECT 70.950 241.950 73.050 244.050 ;
        RECT 74.700 242.400 76.500 251.250 ;
        RECT 80.100 243.000 81.900 251.250 ;
        RECT 93.000 245.400 94.800 251.250 ;
        RECT 97.200 247.050 99.000 251.250 ;
        RECT 100.500 248.400 102.300 251.250 ;
        RECT 106.950 247.950 109.050 250.050 ;
        RECT 110.550 248.400 112.350 251.250 ;
        RECT 113.550 248.400 115.350 251.250 ;
        RECT 116.550 248.400 118.350 251.250 ;
        RECT 97.200 245.400 102.900 247.050 ;
        RECT 62.100 240.150 63.900 241.950 ;
        RECT 58.950 236.850 61.050 238.950 ;
        RECT 61.950 238.050 64.050 240.150 ;
        RECT 64.950 236.850 67.050 238.950 ;
        RECT 8.400 231.600 9.600 236.850 ;
        RECT 20.100 235.050 21.900 236.850 ;
        RECT 25.950 231.600 27.150 236.850 ;
        RECT 28.950 233.850 31.050 235.950 ;
        RECT 38.100 235.050 39.900 236.850 ;
        RECT 28.950 232.050 30.750 233.850 ;
        RECT 43.950 231.600 45.150 236.850 ;
        RECT 46.950 233.850 49.050 235.950 ;
        RECT 55.950 233.850 58.050 235.950 ;
        RECT 46.950 232.050 48.750 233.850 ;
        RECT 56.250 232.050 58.050 233.850 ;
        RECT 59.850 231.600 61.050 236.850 ;
        RECT 65.100 235.050 66.900 236.850 ;
        RECT 71.550 235.050 72.450 241.950 ;
        RECT 80.100 241.350 84.600 243.000 ;
        RECT 83.400 237.150 84.600 241.350 ;
        RECT 92.100 240.150 93.900 241.950 ;
        RECT 91.950 238.050 94.050 240.150 ;
        RECT 94.950 239.850 97.050 241.950 ;
        RECT 98.100 240.150 99.900 241.950 ;
        RECT 95.100 238.050 96.900 239.850 ;
        RECT 97.950 238.050 100.050 240.150 ;
        RECT 101.700 238.950 102.900 245.400 ;
        RECT 70.950 232.950 73.050 235.050 ;
        RECT 73.950 233.850 76.050 235.950 ;
        RECT 79.950 233.850 82.050 235.950 ;
        RECT 82.950 235.050 85.050 237.150 ;
        RECT 100.950 236.850 103.050 238.950 ;
        RECT 107.550 238.050 108.450 247.950 ;
        RECT 114.000 241.950 115.050 248.400 ;
        RECT 128.550 246.300 130.350 251.250 ;
        RECT 131.550 247.200 133.350 251.250 ;
        RECT 134.550 246.300 136.350 251.250 ;
        RECT 128.550 244.950 136.350 246.300 ;
        RECT 137.550 245.400 139.350 251.250 ;
        RECT 146.550 248.400 148.350 251.250 ;
        RECT 149.550 248.400 151.350 251.250 ;
        RECT 152.550 248.400 154.350 251.250 ;
        RECT 163.650 248.400 165.450 251.250 ;
        RECT 166.650 248.400 168.450 251.250 ;
        RECT 169.650 248.400 171.450 251.250 ;
        RECT 176.550 248.400 178.350 251.250 ;
        RECT 179.550 248.400 181.350 251.250 ;
        RECT 137.550 243.300 138.750 245.400 ;
        RECT 135.000 242.250 138.750 243.300 ;
        RECT 112.950 239.850 115.050 241.950 ;
        RECT 131.100 240.150 132.900 241.950 ;
        RECT 74.100 232.050 75.900 233.850 ;
        RECT 7.650 219.750 9.450 231.600 ;
        RECT 10.650 219.750 12.450 231.600 ;
        RECT 21.300 219.750 23.100 231.600 ;
        RECT 25.500 219.750 27.300 231.600 ;
        RECT 28.800 219.750 30.600 225.600 ;
        RECT 39.300 219.750 41.100 231.600 ;
        RECT 43.500 219.750 45.300 231.600 ;
        RECT 46.800 219.750 48.600 225.600 ;
        RECT 56.400 219.750 58.200 225.600 ;
        RECT 59.700 219.750 61.500 231.600 ;
        RECT 63.900 219.750 65.700 231.600 ;
        RECT 76.950 230.850 79.050 232.950 ;
        RECT 80.250 232.050 82.050 233.850 ;
        RECT 77.100 229.050 78.900 230.850 ;
        RECT 83.700 226.800 84.750 235.050 ;
        RECT 101.700 231.600 102.900 236.850 ;
        RECT 106.950 235.950 109.050 238.050 ;
        RECT 109.950 236.850 112.050 238.950 ;
        RECT 110.100 235.050 111.900 236.850 ;
        RECT 114.000 232.650 115.050 239.850 ;
        RECT 115.950 236.850 118.050 238.950 ;
        RECT 127.950 236.850 130.050 238.950 ;
        RECT 130.950 238.050 133.050 240.150 ;
        RECT 134.850 238.950 136.050 242.250 ;
        RECT 139.950 241.950 142.050 244.050 ;
        RECT 150.000 241.950 151.050 248.400 ;
        RECT 133.950 236.850 136.050 238.950 ;
        RECT 116.100 235.050 117.900 236.850 ;
        RECT 128.100 235.050 129.900 236.850 ;
        RECT 114.000 231.600 116.550 232.650 ;
        RECT 133.950 231.600 135.150 236.850 ;
        RECT 136.950 233.850 139.050 235.950 ;
        RECT 136.950 232.050 138.750 233.850 ;
        RECT 77.700 225.900 84.750 226.800 ;
        RECT 77.700 225.600 79.350 225.900 ;
        RECT 74.550 219.750 76.350 225.600 ;
        RECT 77.550 219.750 79.350 225.600 ;
        RECT 83.550 225.600 84.750 225.900 ;
        RECT 92.550 230.700 100.350 231.600 ;
        RECT 80.550 219.750 82.350 225.000 ;
        RECT 83.550 219.750 85.350 225.600 ;
        RECT 92.550 219.750 94.350 230.700 ;
        RECT 95.550 219.750 97.350 229.800 ;
        RECT 98.550 219.750 100.350 230.700 ;
        RECT 101.550 219.750 103.350 231.600 ;
        RECT 110.550 219.750 112.350 231.600 ;
        RECT 114.750 219.750 116.550 231.600 ;
        RECT 129.300 219.750 131.100 231.600 ;
        RECT 133.500 219.750 135.300 231.600 ;
        RECT 136.950 228.450 139.050 229.050 ;
        RECT 140.550 228.450 141.450 241.950 ;
        RECT 148.950 239.850 151.050 241.950 ;
        RECT 145.950 236.850 148.050 238.950 ;
        RECT 146.100 235.050 147.900 236.850 ;
        RECT 150.000 232.650 151.050 239.850 ;
        RECT 166.950 241.950 168.000 248.400 ;
        RECT 166.950 239.850 169.050 241.950 ;
        RECT 175.950 239.850 178.050 241.950 ;
        RECT 179.400 240.150 180.600 248.400 ;
        RECT 188.550 246.300 190.350 251.250 ;
        RECT 191.550 247.200 193.350 251.250 ;
        RECT 194.550 246.300 196.350 251.250 ;
        RECT 188.550 244.950 196.350 246.300 ;
        RECT 197.550 245.400 199.350 251.250 ;
        RECT 197.550 243.300 198.750 245.400 ;
        RECT 195.000 242.250 198.750 243.300 ;
        RECT 206.550 243.900 208.350 251.250 ;
        RECT 211.050 245.400 212.850 251.250 ;
        RECT 214.050 246.900 215.850 251.250 ;
        RECT 214.050 245.400 217.350 246.900 ;
        RECT 224.850 245.400 226.650 251.250 ;
        RECT 212.250 243.900 214.050 244.500 ;
        RECT 206.550 242.700 214.050 243.900 ;
        RECT 191.100 240.150 192.900 241.950 ;
        RECT 151.950 236.850 154.050 238.950 ;
        RECT 163.950 236.850 166.050 238.950 ;
        RECT 152.100 235.050 153.900 236.850 ;
        RECT 164.100 235.050 165.900 236.850 ;
        RECT 166.950 232.650 168.000 239.850 ;
        RECT 169.950 236.850 172.050 238.950 ;
        RECT 176.100 238.050 177.900 239.850 ;
        RECT 178.950 238.050 181.050 240.150 ;
        RECT 170.100 235.050 171.900 236.850 ;
        RECT 150.000 231.600 152.550 232.650 ;
        RECT 136.950 227.550 141.450 228.450 ;
        RECT 136.950 226.950 139.050 227.550 ;
        RECT 136.800 219.750 138.600 225.600 ;
        RECT 146.550 219.750 148.350 231.600 ;
        RECT 150.750 219.750 152.550 231.600 ;
        RECT 165.450 231.600 168.000 232.650 ;
        RECT 165.450 219.750 167.250 231.600 ;
        RECT 169.650 219.750 171.450 231.600 ;
        RECT 179.400 225.600 180.600 238.050 ;
        RECT 187.950 236.850 190.050 238.950 ;
        RECT 190.950 238.050 193.050 240.150 ;
        RECT 194.850 238.950 196.050 242.250 ;
        RECT 193.950 236.850 196.050 238.950 ;
        RECT 205.950 236.850 208.050 238.950 ;
        RECT 188.100 235.050 189.900 236.850 ;
        RECT 193.950 231.600 195.150 236.850 ;
        RECT 196.950 233.850 199.050 235.950 ;
        RECT 206.100 235.050 207.900 236.850 ;
        RECT 196.950 232.050 198.750 233.850 ;
        RECT 176.550 219.750 178.350 225.600 ;
        RECT 179.550 219.750 181.350 225.600 ;
        RECT 189.300 219.750 191.100 231.600 ;
        RECT 193.500 219.750 195.300 231.600 ;
        RECT 209.700 225.600 210.900 242.700 ;
        RECT 216.150 238.950 217.350 245.400 ;
        RECT 229.350 244.200 231.150 251.250 ;
        RECT 239.850 245.400 241.650 251.250 ;
        RECT 244.350 244.200 246.150 251.250 ;
        RECT 256.650 245.400 258.450 251.250 ;
        RECT 227.550 243.300 231.150 244.200 ;
        RECT 242.550 243.300 246.150 244.200 ;
        RECT 257.250 243.300 258.450 245.400 ;
        RECT 259.650 246.300 261.450 251.250 ;
        RECT 262.650 247.200 264.450 251.250 ;
        RECT 265.650 246.300 267.450 251.250 ;
        RECT 272.550 248.400 274.350 251.250 ;
        RECT 275.550 248.400 277.350 251.250 ;
        RECT 259.650 244.950 267.450 246.300 ;
        RECT 212.100 237.150 213.900 238.950 ;
        RECT 211.950 235.050 214.050 237.150 ;
        RECT 214.950 236.850 217.350 238.950 ;
        RECT 224.100 237.150 225.900 238.950 ;
        RECT 216.150 231.600 217.350 236.850 ;
        RECT 223.950 235.050 226.050 237.150 ;
        RECT 227.550 235.950 228.750 243.300 ;
        RECT 230.100 237.150 231.900 238.950 ;
        RECT 239.100 237.150 240.900 238.950 ;
        RECT 226.950 233.850 229.050 235.950 ;
        RECT 229.950 235.050 232.050 237.150 ;
        RECT 238.950 235.050 241.050 237.150 ;
        RECT 242.550 235.950 243.750 243.300 ;
        RECT 257.250 242.250 261.000 243.300 ;
        RECT 259.950 238.950 261.150 242.250 ;
        RECT 263.100 240.150 264.900 241.950 ;
        RECT 245.100 237.150 246.900 238.950 ;
        RECT 241.950 233.850 244.050 235.950 ;
        RECT 244.950 235.050 247.050 237.150 ;
        RECT 259.950 236.850 262.050 238.950 ;
        RECT 262.950 238.050 265.050 240.150 ;
        RECT 271.950 239.850 274.050 241.950 ;
        RECT 275.400 240.150 276.600 248.400 ;
        RECT 287.850 244.200 289.650 251.250 ;
        RECT 292.350 245.400 294.150 251.250 ;
        RECT 299.850 245.400 301.650 251.250 ;
        RECT 304.350 244.200 306.150 251.250 ;
        RECT 287.850 243.300 291.450 244.200 ;
        RECT 265.950 236.850 268.050 238.950 ;
        RECT 272.100 238.050 273.900 239.850 ;
        RECT 274.950 238.050 277.050 240.150 ;
        RECT 256.950 233.850 259.050 235.950 ;
        RECT 196.800 219.750 198.600 225.600 ;
        RECT 206.550 219.750 208.350 225.600 ;
        RECT 209.550 219.750 211.350 225.600 ;
        RECT 213.150 219.750 214.950 231.600 ;
        RECT 216.150 219.750 217.950 231.600 ;
        RECT 227.550 225.600 228.750 233.850 ;
        RECT 242.550 225.600 243.750 233.850 ;
        RECT 257.250 232.050 259.050 233.850 ;
        RECT 260.850 231.600 262.050 236.850 ;
        RECT 266.100 235.050 267.900 236.850 ;
        RECT 224.550 219.750 226.350 225.600 ;
        RECT 227.550 219.750 229.350 225.600 ;
        RECT 230.550 219.750 232.350 225.600 ;
        RECT 239.550 219.750 241.350 225.600 ;
        RECT 242.550 219.750 244.350 225.600 ;
        RECT 245.550 219.750 247.350 225.600 ;
        RECT 257.400 219.750 259.200 225.600 ;
        RECT 260.700 219.750 262.500 231.600 ;
        RECT 264.900 219.750 266.700 231.600 ;
        RECT 275.400 225.600 276.600 238.050 ;
        RECT 287.100 237.150 288.900 238.950 ;
        RECT 286.950 235.050 289.050 237.150 ;
        RECT 290.250 235.950 291.450 243.300 ;
        RECT 302.550 243.300 306.150 244.200 ;
        RECT 311.700 245.400 313.500 251.250 ;
        RECT 317.100 245.400 318.900 251.250 ;
        RECT 322.500 245.400 324.300 251.250 ;
        RECT 326.700 248.400 328.500 251.250 ;
        RECT 329.700 248.400 331.500 251.250 ;
        RECT 332.700 248.400 334.500 251.250 ;
        RECT 335.700 248.400 337.500 251.250 ;
        RECT 326.700 247.050 328.050 248.400 ;
        RECT 329.700 247.050 331.050 248.400 ;
        RECT 332.700 247.050 334.050 248.400 ;
        RECT 340.200 247.500 342.000 251.250 ;
        RECT 343.200 248.400 345.000 251.250 ;
        RECT 346.200 247.500 348.000 251.250 ;
        RECT 293.100 237.150 294.900 238.950 ;
        RECT 299.100 237.150 300.900 238.950 ;
        RECT 289.950 233.850 292.050 235.950 ;
        RECT 292.950 235.050 295.050 237.150 ;
        RECT 298.950 235.050 301.050 237.150 ;
        RECT 302.550 235.950 303.750 243.300 ;
        RECT 311.700 241.800 312.900 245.400 ;
        RECT 322.800 244.500 324.300 245.400 ;
        RECT 315.900 243.300 324.300 244.500 ;
        RECT 325.950 244.950 328.050 247.050 ;
        RECT 328.950 244.950 331.050 247.050 ;
        RECT 331.950 244.950 334.050 247.050 ;
        RECT 337.500 246.750 339.300 247.200 ;
        RECT 335.250 245.400 339.300 246.750 ;
        RECT 340.200 245.700 343.050 247.500 ;
        RECT 340.950 245.400 343.050 245.700 ;
        RECT 345.150 245.700 348.000 247.500 ;
        RECT 349.950 247.500 351.750 251.250 ;
        RECT 352.950 247.500 354.750 251.250 ;
        RECT 355.950 247.500 357.750 251.250 ;
        RECT 345.150 245.400 347.250 245.700 ;
        RECT 349.950 245.400 352.050 247.500 ;
        RECT 352.950 245.400 355.050 247.500 ;
        RECT 355.950 245.400 358.050 247.500 ;
        RECT 360.600 246.600 362.400 251.250 ;
        RECT 360.600 245.400 364.800 246.600 ;
        RECT 366.150 245.400 367.950 251.250 ;
        RECT 371.550 245.400 373.350 251.250 ;
        RECT 315.900 242.700 317.700 243.300 ;
        RECT 325.950 241.800 327.000 244.950 ;
        RECT 335.250 244.050 336.150 245.400 ;
        RECT 331.050 243.900 336.150 244.050 ;
        RECT 311.700 240.900 327.000 241.800 ;
        RECT 328.500 243.150 336.150 243.900 ;
        RECT 328.500 242.700 332.850 243.150 ;
        RECT 344.100 242.700 351.000 244.500 ;
        RECT 351.900 242.700 358.650 244.500 ;
        RECT 305.100 237.150 306.900 238.950 ;
        RECT 301.950 233.850 304.050 235.950 ;
        RECT 304.950 235.050 307.050 237.150 ;
        RECT 290.250 225.600 291.450 233.850 ;
        RECT 302.550 225.600 303.750 233.850 ;
        RECT 311.700 227.400 312.900 240.900 ;
        RECT 314.100 238.950 325.950 240.000 ;
        RECT 328.500 239.250 329.550 242.700 ;
        RECT 331.050 242.250 332.850 242.700 ;
        RECT 337.950 241.650 340.050 241.950 ;
        RECT 349.950 241.800 351.000 242.700 ;
        RECT 363.300 241.800 364.800 245.400 ;
        RECT 336.150 239.850 340.050 241.650 ;
        RECT 341.400 240.450 349.050 241.800 ;
        RECT 349.950 240.750 359.850 241.800 ;
        RECT 314.100 237.150 315.900 238.950 ;
        RECT 313.950 235.050 316.050 237.150 ;
        RECT 324.750 236.550 325.950 238.950 ;
        RECT 327.750 237.450 329.550 239.250 ;
        RECT 341.400 238.950 342.450 240.450 ;
        RECT 348.150 239.700 349.050 240.450 ;
        RECT 330.450 238.050 342.450 238.950 ;
        RECT 330.450 236.550 331.500 238.050 ;
        RECT 343.350 237.750 347.250 239.550 ;
        RECT 348.150 238.650 357.750 239.700 ;
        RECT 345.150 237.450 347.250 237.750 ;
        RECT 319.950 235.650 322.050 235.950 ;
        RECT 324.750 235.650 331.500 236.550 ;
        RECT 332.400 236.550 334.200 237.150 ;
        RECT 340.950 236.550 343.050 236.850 ;
        RECT 332.400 235.950 343.050 236.550 ;
        RECT 353.700 235.950 355.500 237.750 ;
        RECT 319.950 234.450 323.850 235.650 ;
        RECT 332.400 235.350 355.500 235.950 ;
        RECT 340.950 234.750 355.500 235.350 ;
        RECT 356.850 237.000 357.750 238.650 ;
        RECT 358.800 238.950 359.850 240.750 ;
        RECT 363.300 240.000 371.100 241.800 ;
        RECT 358.800 237.900 367.050 238.950 ;
        RECT 356.850 235.200 363.900 237.000 ;
        RECT 319.950 233.850 333.900 234.450 ;
        RECT 364.950 233.850 367.050 237.900 ;
        RECT 320.250 233.550 360.000 233.850 ;
        RECT 331.950 232.650 360.000 233.550 ;
        RECT 369.450 232.650 371.250 233.250 ;
        RECT 319.500 232.050 321.300 232.650 ;
        RECT 328.950 232.050 331.050 232.350 ;
        RECT 319.500 230.850 331.050 232.050 ;
        RECT 328.950 230.250 331.050 230.850 ;
        RECT 331.950 230.400 352.050 231.750 ;
        RECT 316.200 229.350 318.000 230.100 ;
        RECT 331.950 229.350 333.900 230.400 ;
        RECT 349.950 229.650 352.050 230.400 ;
        RECT 355.950 230.550 358.050 231.750 ;
        RECT 358.950 231.450 371.250 232.650 ;
        RECT 372.150 230.550 373.350 245.400 ;
        RECT 355.950 229.650 373.350 230.550 ;
        RECT 375.450 248.400 377.250 251.250 ;
        RECT 378.450 248.400 380.250 251.250 ;
        RECT 391.650 250.500 399.450 251.250 ;
        RECT 375.450 240.150 376.950 248.400 ;
        RECT 391.650 245.400 393.450 250.500 ;
        RECT 394.650 245.400 396.450 249.600 ;
        RECT 397.650 246.000 399.450 250.500 ;
        RECT 400.650 246.900 402.450 251.250 ;
        RECT 403.650 246.000 405.450 251.250 ;
        RECT 395.250 243.900 396.150 245.400 ;
        RECT 397.650 245.100 405.450 246.000 ;
        RECT 410.850 245.400 412.650 251.250 ;
        RECT 415.350 244.200 417.150 251.250 ;
        RECT 395.250 242.850 399.600 243.900 ;
        RECT 395.700 240.150 397.500 241.950 ;
        RECT 375.450 238.050 379.050 240.150 ;
        RECT 316.200 228.300 333.900 229.350 ;
        RECT 311.700 226.500 315.750 227.400 ;
        RECT 314.700 225.600 315.750 226.500 ;
        RECT 272.550 219.750 274.350 225.600 ;
        RECT 275.550 219.750 277.350 225.600 ;
        RECT 286.650 219.750 288.450 225.600 ;
        RECT 289.650 219.750 291.450 225.600 ;
        RECT 292.650 219.750 294.450 225.600 ;
        RECT 299.550 219.750 301.350 225.600 ;
        RECT 302.550 219.750 304.350 225.600 ;
        RECT 305.550 219.750 307.350 225.600 ;
        RECT 311.700 219.750 313.500 225.600 ;
        RECT 314.700 219.750 316.500 225.600 ;
        RECT 317.700 219.750 319.500 225.600 ;
        RECT 320.700 219.750 322.500 228.300 ;
        RECT 340.950 228.150 343.050 228.600 ;
        RECT 340.650 226.500 343.050 228.150 ;
        RECT 345.000 226.800 348.900 228.600 ;
        RECT 345.000 226.500 348.000 226.800 ;
        RECT 325.950 223.950 328.050 226.050 ;
        RECT 328.950 223.950 331.050 226.050 ;
        RECT 331.950 225.600 334.050 226.050 ;
        RECT 340.650 225.600 342.000 226.500 ;
        RECT 331.950 223.950 334.500 225.600 ;
        RECT 323.700 219.750 325.500 223.050 ;
        RECT 326.850 222.600 328.050 223.950 ;
        RECT 330.150 222.600 331.050 223.950 ;
        RECT 333.300 222.600 334.500 223.950 ;
        RECT 326.850 219.750 329.250 222.600 ;
        RECT 330.150 219.750 332.250 222.600 ;
        RECT 333.300 219.750 335.250 222.600 ;
        RECT 336.450 219.750 338.250 225.600 ;
        RECT 340.200 219.750 342.000 225.600 ;
        RECT 343.200 219.750 345.000 225.600 ;
        RECT 346.200 219.750 348.000 226.500 ;
        RECT 350.100 222.600 351.450 229.650 ;
        RECT 359.850 228.150 361.650 228.300 ;
        RECT 352.950 226.950 361.650 228.150 ;
        RECT 366.600 227.700 368.400 228.300 ;
        RECT 352.950 226.050 355.050 226.950 ;
        RECT 359.850 226.500 361.650 226.950 ;
        RECT 362.700 226.500 368.400 227.700 ;
        RECT 349.950 219.750 351.750 222.600 ;
        RECT 352.950 219.750 354.750 226.050 ;
        RECT 356.100 223.800 358.200 225.900 ;
        RECT 356.100 222.600 357.600 223.800 ;
        RECT 355.950 219.750 357.750 222.600 ;
        RECT 359.700 219.750 361.500 225.600 ;
        RECT 362.700 219.750 364.500 226.500 ;
        RECT 369.300 225.600 370.500 229.650 ;
        RECT 375.450 225.600 376.950 238.050 ;
        RECT 391.950 236.850 394.050 238.950 ;
        RECT 394.950 238.050 397.050 240.150 ;
        RECT 398.400 238.950 399.600 242.850 ;
        RECT 413.550 243.300 417.150 244.200 ;
        RECT 401.100 240.150 402.900 241.950 ;
        RECT 397.950 236.850 400.050 238.950 ;
        RECT 400.950 238.050 403.050 240.150 ;
        RECT 403.950 236.850 406.050 238.950 ;
        RECT 410.100 237.150 411.900 238.950 ;
        RECT 392.250 235.050 394.050 236.850 ;
        RECT 398.250 231.600 399.450 236.850 ;
        RECT 404.100 235.050 405.900 236.850 ;
        RECT 409.950 235.050 412.050 237.150 ;
        RECT 413.550 235.950 414.750 243.300 ;
        RECT 425.700 242.400 427.500 251.250 ;
        RECT 431.100 243.000 432.900 251.250 ;
        RECT 447.000 245.400 448.800 251.250 ;
        RECT 451.200 247.050 453.000 251.250 ;
        RECT 454.500 248.400 456.300 251.250 ;
        RECT 451.200 245.400 456.900 247.050 ;
        RECT 431.100 241.350 435.600 243.000 ;
        RECT 442.950 241.950 445.050 244.050 ;
        RECT 416.100 237.150 417.900 238.950 ;
        RECT 434.400 237.150 435.600 241.350 ;
        RECT 412.950 233.850 415.050 235.950 ;
        RECT 415.950 235.050 418.050 237.150 ;
        RECT 424.950 233.850 427.050 235.950 ;
        RECT 430.950 233.850 433.050 235.950 ;
        RECT 433.950 235.050 436.050 237.150 ;
        RECT 365.700 219.750 367.500 225.600 ;
        RECT 368.700 219.750 370.500 225.600 ;
        RECT 371.700 219.750 373.500 225.600 ;
        RECT 375.450 219.750 377.250 225.600 ;
        RECT 378.450 219.750 380.250 225.600 ;
        RECT 393.150 219.750 394.950 231.600 ;
        RECT 397.650 219.750 400.950 231.600 ;
        RECT 403.650 219.750 405.450 231.600 ;
        RECT 413.550 225.600 414.750 233.850 ;
        RECT 425.100 232.050 426.900 233.850 ;
        RECT 427.950 230.850 430.050 232.950 ;
        RECT 431.250 232.050 433.050 233.850 ;
        RECT 428.100 229.050 429.900 230.850 ;
        RECT 434.700 226.800 435.750 235.050 ;
        RECT 428.700 225.900 435.750 226.800 ;
        RECT 428.700 225.600 430.350 225.900 ;
        RECT 410.550 219.750 412.350 225.600 ;
        RECT 413.550 219.750 415.350 225.600 ;
        RECT 416.550 219.750 418.350 225.600 ;
        RECT 425.550 219.750 427.350 225.600 ;
        RECT 428.550 219.750 430.350 225.600 ;
        RECT 434.550 225.600 435.750 225.900 ;
        RECT 431.550 219.750 433.350 225.000 ;
        RECT 434.550 219.750 436.350 225.600 ;
        RECT 439.950 222.450 442.050 223.050 ;
        RECT 443.550 222.450 444.450 241.950 ;
        RECT 446.100 240.150 447.900 241.950 ;
        RECT 445.950 238.050 448.050 240.150 ;
        RECT 448.950 239.850 451.050 241.950 ;
        RECT 452.100 240.150 453.900 241.950 ;
        RECT 449.100 238.050 450.900 239.850 ;
        RECT 451.950 238.050 454.050 240.150 ;
        RECT 455.700 238.950 456.900 245.400 ;
        RECT 461.550 246.000 463.350 251.250 ;
        RECT 464.550 246.900 466.350 251.250 ;
        RECT 467.550 250.500 475.350 251.250 ;
        RECT 467.550 246.000 469.350 250.500 ;
        RECT 461.550 245.100 469.350 246.000 ;
        RECT 470.550 245.400 472.350 249.600 ;
        RECT 473.550 245.400 475.350 250.500 ;
        RECT 470.850 243.900 471.750 245.400 ;
        RECT 467.400 242.850 471.750 243.900 ;
        RECT 488.100 243.000 489.900 251.250 ;
        RECT 464.100 240.150 465.900 241.950 ;
        RECT 454.950 236.850 457.050 238.950 ;
        RECT 460.950 236.850 463.050 238.950 ;
        RECT 463.950 238.050 466.050 240.150 ;
        RECT 467.400 238.950 468.600 242.850 ;
        RECT 469.500 240.150 471.300 241.950 ;
        RECT 485.400 241.350 489.900 243.000 ;
        RECT 493.500 242.400 495.300 251.250 ;
        RECT 502.650 248.400 504.450 251.250 ;
        RECT 505.650 248.400 507.450 251.250 ;
        RECT 466.950 236.850 469.050 238.950 ;
        RECT 469.950 238.050 472.050 240.150 ;
        RECT 472.950 236.850 475.050 238.950 ;
        RECT 485.400 237.150 486.600 241.350 ;
        RECT 503.400 240.150 504.600 248.400 ;
        RECT 512.850 245.400 514.650 251.250 ;
        RECT 517.350 244.200 519.150 251.250 ;
        RECT 528.000 245.400 529.800 251.250 ;
        RECT 532.200 247.050 534.000 251.250 ;
        RECT 535.500 248.400 537.300 251.250 ;
        RECT 532.200 245.400 537.900 247.050 ;
        RECT 511.950 243.450 514.050 244.050 ;
        RECT 509.550 242.550 514.050 243.450 ;
        RECT 502.950 238.050 505.050 240.150 ;
        RECT 505.950 239.850 508.050 241.950 ;
        RECT 506.100 238.050 507.900 239.850 ;
        RECT 455.700 231.600 456.900 236.850 ;
        RECT 461.100 235.050 462.900 236.850 ;
        RECT 467.550 231.600 468.750 236.850 ;
        RECT 472.950 235.050 474.750 236.850 ;
        RECT 484.950 235.050 487.050 237.150 ;
        RECT 439.950 221.550 444.450 222.450 ;
        RECT 446.550 230.700 454.350 231.600 ;
        RECT 439.950 220.950 442.050 221.550 ;
        RECT 446.550 219.750 448.350 230.700 ;
        RECT 449.550 219.750 451.350 229.800 ;
        RECT 452.550 219.750 454.350 230.700 ;
        RECT 455.550 219.750 457.350 231.600 ;
        RECT 461.550 219.750 463.350 231.600 ;
        RECT 466.050 219.750 469.350 231.600 ;
        RECT 472.050 219.750 473.850 231.600 ;
        RECT 485.250 226.800 486.300 235.050 ;
        RECT 487.950 233.850 490.050 235.950 ;
        RECT 493.950 233.850 496.050 235.950 ;
        RECT 487.950 232.050 489.750 233.850 ;
        RECT 490.950 230.850 493.050 232.950 ;
        RECT 494.100 232.050 495.900 233.850 ;
        RECT 491.100 229.050 492.900 230.850 ;
        RECT 485.250 225.900 492.300 226.800 ;
        RECT 485.250 225.600 486.450 225.900 ;
        RECT 484.650 219.750 486.450 225.600 ;
        RECT 490.650 225.600 492.300 225.900 ;
        RECT 503.400 225.600 504.600 238.050 ;
        RECT 505.950 234.450 508.050 235.050 ;
        RECT 509.550 234.450 510.450 242.550 ;
        RECT 511.950 241.950 514.050 242.550 ;
        RECT 515.550 243.300 519.150 244.200 ;
        RECT 512.100 237.150 513.900 238.950 ;
        RECT 511.950 235.050 514.050 237.150 ;
        RECT 515.550 235.950 516.750 243.300 ;
        RECT 527.100 240.150 528.900 241.950 ;
        RECT 518.100 237.150 519.900 238.950 ;
        RECT 526.950 238.050 529.050 240.150 ;
        RECT 529.950 239.850 532.050 241.950 ;
        RECT 533.100 240.150 534.900 241.950 ;
        RECT 530.100 238.050 531.900 239.850 ;
        RECT 532.950 238.050 535.050 240.150 ;
        RECT 536.700 238.950 537.900 245.400 ;
        RECT 548.850 244.200 550.650 251.250 ;
        RECT 553.350 245.400 555.150 251.250 ;
        RECT 548.850 243.300 552.450 244.200 ;
        RECT 505.950 233.550 510.450 234.450 ;
        RECT 514.950 233.850 517.050 235.950 ;
        RECT 517.950 235.050 520.050 237.150 ;
        RECT 535.950 236.850 538.050 238.950 ;
        RECT 548.100 237.150 549.900 238.950 ;
        RECT 505.950 232.950 508.050 233.550 ;
        RECT 515.550 225.600 516.750 233.850 ;
        RECT 536.700 231.600 537.900 236.850 ;
        RECT 547.950 235.050 550.050 237.150 ;
        RECT 551.250 235.950 552.450 243.300 ;
        RECT 566.100 243.000 567.900 251.250 ;
        RECT 563.400 241.350 567.900 243.000 ;
        RECT 571.500 242.400 573.300 251.250 ;
        RECT 577.650 248.400 579.450 251.250 ;
        RECT 580.650 248.400 582.450 251.250 ;
        RECT 583.650 248.400 585.450 251.250 ;
        RECT 580.950 241.950 582.000 248.400 ;
        RECT 594.000 245.400 595.800 251.250 ;
        RECT 598.200 247.050 600.000 251.250 ;
        RECT 601.500 248.400 603.300 251.250 ;
        RECT 598.200 245.400 603.900 247.050 ;
        RECT 583.950 243.450 586.050 244.050 ;
        RECT 583.950 242.550 591.450 243.450 ;
        RECT 583.950 241.950 586.050 242.550 ;
        RECT 554.100 237.150 555.900 238.950 ;
        RECT 563.400 237.150 564.600 241.350 ;
        RECT 580.950 239.850 583.050 241.950 ;
        RECT 550.950 233.850 553.050 235.950 ;
        RECT 553.950 235.050 556.050 237.150 ;
        RECT 562.950 235.050 565.050 237.150 ;
        RECT 577.950 236.850 580.050 238.950 ;
        RECT 527.550 230.700 535.350 231.600 ;
        RECT 487.650 219.750 489.450 225.000 ;
        RECT 490.650 219.750 492.450 225.600 ;
        RECT 493.650 219.750 495.450 225.600 ;
        RECT 502.650 219.750 504.450 225.600 ;
        RECT 505.650 219.750 507.450 225.600 ;
        RECT 512.550 219.750 514.350 225.600 ;
        RECT 515.550 219.750 517.350 225.600 ;
        RECT 518.550 219.750 520.350 225.600 ;
        RECT 527.550 219.750 529.350 230.700 ;
        RECT 530.550 219.750 532.350 229.800 ;
        RECT 533.550 219.750 535.350 230.700 ;
        RECT 536.550 219.750 538.350 231.600 ;
        RECT 551.250 225.600 552.450 233.850 ;
        RECT 563.250 226.800 564.300 235.050 ;
        RECT 565.950 233.850 568.050 235.950 ;
        RECT 571.950 233.850 574.050 235.950 ;
        RECT 578.100 235.050 579.900 236.850 ;
        RECT 565.950 232.050 567.750 233.850 ;
        RECT 568.950 230.850 571.050 232.950 ;
        RECT 572.100 232.050 573.900 233.850 ;
        RECT 580.950 232.650 582.000 239.850 ;
        RECT 583.950 236.850 586.050 238.950 ;
        RECT 584.100 235.050 585.900 236.850 ;
        RECT 590.550 234.450 591.450 242.550 ;
        RECT 593.100 240.150 594.900 241.950 ;
        RECT 592.950 238.050 595.050 240.150 ;
        RECT 595.950 239.850 598.050 241.950 ;
        RECT 599.100 240.150 600.900 241.950 ;
        RECT 596.100 238.050 597.900 239.850 ;
        RECT 598.950 238.050 601.050 240.150 ;
        RECT 602.700 238.950 603.900 245.400 ;
        RECT 608.700 242.400 610.500 251.250 ;
        RECT 614.100 243.000 615.900 251.250 ;
        RECT 624.000 245.400 625.800 251.250 ;
        RECT 628.200 247.050 630.000 251.250 ;
        RECT 631.500 248.400 633.300 251.250 ;
        RECT 628.200 245.400 633.900 247.050 ;
        RECT 643.650 245.400 645.450 251.250 ;
        RECT 614.100 241.350 618.600 243.000 ;
        RECT 601.950 236.850 604.050 238.950 ;
        RECT 617.400 237.150 618.600 241.350 ;
        RECT 623.100 240.150 624.900 241.950 ;
        RECT 622.950 238.050 625.050 240.150 ;
        RECT 625.950 239.850 628.050 241.950 ;
        RECT 629.100 240.150 630.900 241.950 ;
        RECT 626.100 238.050 627.900 239.850 ;
        RECT 628.950 238.050 631.050 240.150 ;
        RECT 632.700 238.950 633.900 245.400 ;
        RECT 644.250 243.300 645.450 245.400 ;
        RECT 646.650 246.300 648.450 251.250 ;
        RECT 649.650 247.200 651.450 251.250 ;
        RECT 652.650 246.300 654.450 251.250 ;
        RECT 664.650 248.400 666.450 251.250 ;
        RECT 667.650 248.400 669.450 251.250 ;
        RECT 646.650 244.950 654.450 246.300 ;
        RECT 644.250 242.250 648.000 243.300 ;
        RECT 646.950 238.950 648.150 242.250 ;
        RECT 650.100 240.150 651.900 241.950 ;
        RECT 665.400 240.150 666.600 248.400 ;
        RECT 671.550 246.300 673.350 251.250 ;
        RECT 674.550 247.200 676.350 251.250 ;
        RECT 677.550 246.300 679.350 251.250 ;
        RECT 671.550 244.950 679.350 246.300 ;
        RECT 680.550 245.400 682.350 251.250 ;
        RECT 692.550 248.400 694.350 251.250 ;
        RECT 695.550 248.400 697.350 251.250 ;
        RECT 698.550 248.400 700.350 251.250 ;
        RECT 680.550 243.300 681.750 245.400 ;
        RECT 678.000 242.250 681.750 243.300 ;
        RECT 592.950 234.450 595.050 235.050 ;
        RECT 590.550 233.550 595.050 234.450 ;
        RECT 592.950 232.950 595.050 233.550 ;
        RECT 579.450 231.600 582.000 232.650 ;
        RECT 602.700 231.600 603.900 236.850 ;
        RECT 607.950 233.850 610.050 235.950 ;
        RECT 613.950 233.850 616.050 235.950 ;
        RECT 616.950 235.050 619.050 237.150 ;
        RECT 631.950 236.850 634.050 238.950 ;
        RECT 646.950 236.850 649.050 238.950 ;
        RECT 649.950 238.050 652.050 240.150 ;
        RECT 652.950 236.850 655.050 238.950 ;
        RECT 664.950 238.050 667.050 240.150 ;
        RECT 667.950 239.850 670.050 241.950 ;
        RECT 674.100 240.150 675.900 241.950 ;
        RECT 668.100 238.050 669.900 239.850 ;
        RECT 608.100 232.050 609.900 233.850 ;
        RECT 569.100 229.050 570.900 230.850 ;
        RECT 563.250 225.900 570.300 226.800 ;
        RECT 563.250 225.600 564.450 225.900 ;
        RECT 547.650 219.750 549.450 225.600 ;
        RECT 550.650 219.750 552.450 225.600 ;
        RECT 553.650 219.750 555.450 225.600 ;
        RECT 562.650 219.750 564.450 225.600 ;
        RECT 568.650 225.600 570.300 225.900 ;
        RECT 565.650 219.750 567.450 225.000 ;
        RECT 568.650 219.750 570.450 225.600 ;
        RECT 571.650 219.750 573.450 225.600 ;
        RECT 579.450 219.750 581.250 231.600 ;
        RECT 583.650 219.750 585.450 231.600 ;
        RECT 593.550 230.700 601.350 231.600 ;
        RECT 593.550 219.750 595.350 230.700 ;
        RECT 596.550 219.750 598.350 229.800 ;
        RECT 599.550 219.750 601.350 230.700 ;
        RECT 602.550 219.750 604.350 231.600 ;
        RECT 610.950 230.850 613.050 232.950 ;
        RECT 614.250 232.050 616.050 233.850 ;
        RECT 611.100 229.050 612.900 230.850 ;
        RECT 617.700 226.800 618.750 235.050 ;
        RECT 619.950 234.450 622.050 235.050 ;
        RECT 628.950 234.450 631.050 235.050 ;
        RECT 619.950 233.550 631.050 234.450 ;
        RECT 619.950 232.950 622.050 233.550 ;
        RECT 628.950 232.950 631.050 233.550 ;
        RECT 632.700 231.600 633.900 236.850 ;
        RECT 643.950 233.850 646.050 235.950 ;
        RECT 644.250 232.050 646.050 233.850 ;
        RECT 647.850 231.600 649.050 236.850 ;
        RECT 653.100 235.050 654.900 236.850 ;
        RECT 611.700 225.900 618.750 226.800 ;
        RECT 611.700 225.600 613.350 225.900 ;
        RECT 608.550 219.750 610.350 225.600 ;
        RECT 611.550 219.750 613.350 225.600 ;
        RECT 617.550 225.600 618.750 225.900 ;
        RECT 623.550 230.700 631.350 231.600 ;
        RECT 614.550 219.750 616.350 225.000 ;
        RECT 617.550 219.750 619.350 225.600 ;
        RECT 623.550 219.750 625.350 230.700 ;
        RECT 626.550 219.750 628.350 229.800 ;
        RECT 629.550 219.750 631.350 230.700 ;
        RECT 632.550 219.750 634.350 231.600 ;
        RECT 644.400 219.750 646.200 225.600 ;
        RECT 647.700 219.750 649.500 231.600 ;
        RECT 651.900 219.750 653.700 231.600 ;
        RECT 665.400 225.600 666.600 238.050 ;
        RECT 670.950 236.850 673.050 238.950 ;
        RECT 673.950 238.050 676.050 240.150 ;
        RECT 677.850 238.950 679.050 242.250 ;
        RECT 696.000 241.950 697.050 248.400 ;
        RECT 710.850 244.200 712.650 251.250 ;
        RECT 715.350 245.400 717.150 251.250 ;
        RECT 722.550 248.400 724.350 251.250 ;
        RECT 725.550 248.400 727.350 251.250 ;
        RECT 728.550 248.400 730.350 251.250 ;
        RECT 739.650 248.400 741.450 251.250 ;
        RECT 742.650 248.400 744.450 251.250 ;
        RECT 745.650 248.400 747.450 251.250 ;
        RECT 752.550 248.400 754.350 251.250 ;
        RECT 755.550 248.400 757.350 251.250 ;
        RECT 758.550 248.400 760.350 251.250 ;
        RECT 710.850 243.300 714.450 244.200 ;
        RECT 694.950 239.850 697.050 241.950 ;
        RECT 676.950 236.850 679.050 238.950 ;
        RECT 691.950 236.850 694.050 238.950 ;
        RECT 671.100 235.050 672.900 236.850 ;
        RECT 676.950 231.600 678.150 236.850 ;
        RECT 679.950 233.850 682.050 235.950 ;
        RECT 692.100 235.050 693.900 236.850 ;
        RECT 679.950 232.050 681.750 233.850 ;
        RECT 696.000 232.650 697.050 239.850 ;
        RECT 697.950 236.850 700.050 238.950 ;
        RECT 710.100 237.150 711.900 238.950 ;
        RECT 698.100 235.050 699.900 236.850 ;
        RECT 709.950 235.050 712.050 237.150 ;
        RECT 713.250 235.950 714.450 243.300 ;
        RECT 726.000 241.950 727.050 248.400 ;
        RECT 724.950 239.850 727.050 241.950 ;
        RECT 716.100 237.150 717.900 238.950 ;
        RECT 712.950 233.850 715.050 235.950 ;
        RECT 715.950 235.050 718.050 237.150 ;
        RECT 721.950 236.850 724.050 238.950 ;
        RECT 722.100 235.050 723.900 236.850 ;
        RECT 696.000 231.600 698.550 232.650 ;
        RECT 664.650 219.750 666.450 225.600 ;
        RECT 667.650 219.750 669.450 225.600 ;
        RECT 672.300 219.750 674.100 231.600 ;
        RECT 676.500 219.750 678.300 231.600 ;
        RECT 679.800 219.750 681.600 225.600 ;
        RECT 692.550 219.750 694.350 231.600 ;
        RECT 696.750 219.750 698.550 231.600 ;
        RECT 713.250 225.600 714.450 233.850 ;
        RECT 726.000 232.650 727.050 239.850 ;
        RECT 742.950 241.950 744.000 248.400 ;
        RECT 756.000 241.950 757.050 248.400 ;
        RECT 767.550 246.300 769.350 251.250 ;
        RECT 770.550 247.200 772.350 251.250 ;
        RECT 773.550 246.300 775.350 251.250 ;
        RECT 767.550 244.950 775.350 246.300 ;
        RECT 776.550 245.400 778.350 251.250 ;
        RECT 787.650 245.400 789.450 251.250 ;
        RECT 757.950 243.450 760.050 244.050 ;
        RECT 763.950 243.450 766.050 244.050 ;
        RECT 757.950 242.550 766.050 243.450 ;
        RECT 776.550 243.300 777.750 245.400 ;
        RECT 757.950 241.950 760.050 242.550 ;
        RECT 763.950 241.950 766.050 242.550 ;
        RECT 774.000 242.250 777.750 243.300 ;
        RECT 788.250 243.300 789.450 245.400 ;
        RECT 790.650 246.300 792.450 251.250 ;
        RECT 793.650 247.200 795.450 251.250 ;
        RECT 796.650 246.300 798.450 251.250 ;
        RECT 803.550 248.400 805.350 251.250 ;
        RECT 806.550 248.400 808.350 251.250 ;
        RECT 809.550 248.400 811.350 251.250 ;
        RECT 790.650 244.950 798.450 246.300 ;
        RECT 788.250 242.250 792.000 243.300 ;
        RECT 742.950 239.850 745.050 241.950 ;
        RECT 754.950 239.850 757.050 241.950 ;
        RECT 770.100 240.150 771.900 241.950 ;
        RECT 727.950 236.850 730.050 238.950 ;
        RECT 739.950 236.850 742.050 238.950 ;
        RECT 728.100 235.050 729.900 236.850 ;
        RECT 740.100 235.050 741.900 236.850 ;
        RECT 742.950 232.650 744.000 239.850 ;
        RECT 745.950 236.850 748.050 238.950 ;
        RECT 751.950 236.850 754.050 238.950 ;
        RECT 746.100 235.050 747.900 236.850 ;
        RECT 752.100 235.050 753.900 236.850 ;
        RECT 726.000 231.600 728.550 232.650 ;
        RECT 709.650 219.750 711.450 225.600 ;
        RECT 712.650 219.750 714.450 225.600 ;
        RECT 715.650 219.750 717.450 225.600 ;
        RECT 722.550 219.750 724.350 231.600 ;
        RECT 726.750 219.750 728.550 231.600 ;
        RECT 741.450 231.600 744.000 232.650 ;
        RECT 756.000 232.650 757.050 239.850 ;
        RECT 757.950 236.850 760.050 238.950 ;
        RECT 766.950 236.850 769.050 238.950 ;
        RECT 769.950 238.050 772.050 240.150 ;
        RECT 773.850 238.950 775.050 242.250 ;
        RECT 775.950 240.450 778.050 241.050 ;
        RECT 787.950 240.450 790.050 241.050 ;
        RECT 775.950 239.550 790.050 240.450 ;
        RECT 775.950 238.950 778.050 239.550 ;
        RECT 787.950 238.950 790.050 239.550 ;
        RECT 790.950 238.950 792.150 242.250 ;
        RECT 807.000 241.950 808.050 248.400 ;
        RECT 823.650 245.400 825.450 251.250 ;
        RECT 826.650 245.400 828.450 251.250 ;
        RECT 833.550 245.400 835.350 251.250 ;
        RECT 836.550 245.400 838.350 251.250 ;
        RECT 794.100 240.150 795.900 241.950 ;
        RECT 772.950 236.850 775.050 238.950 ;
        RECT 790.950 236.850 793.050 238.950 ;
        RECT 793.950 238.050 796.050 240.150 ;
        RECT 805.950 239.850 808.050 241.950 ;
        RECT 796.950 236.850 799.050 238.950 ;
        RECT 802.950 236.850 805.050 238.950 ;
        RECT 758.100 235.050 759.900 236.850 ;
        RECT 767.100 235.050 768.900 236.850 ;
        RECT 756.000 231.600 758.550 232.650 ;
        RECT 772.950 231.600 774.150 236.850 ;
        RECT 775.950 233.850 778.050 235.950 ;
        RECT 787.950 233.850 790.050 235.950 ;
        RECT 775.950 232.050 777.750 233.850 ;
        RECT 788.250 232.050 790.050 233.850 ;
        RECT 791.850 231.600 793.050 236.850 ;
        RECT 797.100 235.050 798.900 236.850 ;
        RECT 803.100 235.050 804.900 236.850 ;
        RECT 807.000 232.650 808.050 239.850 ;
        RECT 824.400 238.950 825.600 245.400 ;
        RECT 827.100 240.150 828.900 241.950 ;
        RECT 833.100 240.150 834.900 241.950 ;
        RECT 808.950 236.850 811.050 238.950 ;
        RECT 823.950 236.850 826.050 238.950 ;
        RECT 826.950 238.050 829.050 240.150 ;
        RECT 832.950 238.050 835.050 240.150 ;
        RECT 836.400 238.950 837.600 245.400 ;
        RECT 845.850 244.200 847.650 251.250 ;
        RECT 850.350 245.400 852.150 251.250 ;
        RECT 845.850 243.300 849.450 244.200 ;
        RECT 835.950 236.850 838.050 238.950 ;
        RECT 845.100 237.150 846.900 238.950 ;
        RECT 809.100 235.050 810.900 236.850 ;
        RECT 807.000 231.600 809.550 232.650 ;
        RECT 824.400 231.600 825.600 236.850 ;
        RECT 836.400 231.600 837.600 236.850 ;
        RECT 844.950 235.050 847.050 237.150 ;
        RECT 848.250 235.950 849.450 243.300 ;
        RECT 851.100 237.150 852.900 238.950 ;
        RECT 847.950 233.850 850.050 235.950 ;
        RECT 850.950 235.050 853.050 237.150 ;
        RECT 741.450 219.750 743.250 231.600 ;
        RECT 745.650 219.750 747.450 231.600 ;
        RECT 752.550 219.750 754.350 231.600 ;
        RECT 756.750 219.750 758.550 231.600 ;
        RECT 768.300 219.750 770.100 231.600 ;
        RECT 772.500 219.750 774.300 231.600 ;
        RECT 775.800 219.750 777.600 225.600 ;
        RECT 788.400 219.750 790.200 225.600 ;
        RECT 791.700 219.750 793.500 231.600 ;
        RECT 795.900 219.750 797.700 231.600 ;
        RECT 803.550 219.750 805.350 231.600 ;
        RECT 807.750 219.750 809.550 231.600 ;
        RECT 823.650 219.750 825.450 231.600 ;
        RECT 826.650 219.750 828.450 231.600 ;
        RECT 833.550 219.750 835.350 231.600 ;
        RECT 836.550 219.750 838.350 231.600 ;
        RECT 848.250 225.600 849.450 233.850 ;
        RECT 844.650 219.750 846.450 225.600 ;
        RECT 847.650 219.750 849.450 225.600 ;
        RECT 850.650 219.750 852.450 225.600 ;
        RECT 7.650 203.400 9.450 215.250 ;
        RECT 10.650 203.400 12.450 215.250 ;
        RECT 24.450 203.400 26.250 215.250 ;
        RECT 28.650 203.400 30.450 215.250 ;
        RECT 34.650 209.400 36.450 215.250 ;
        RECT 37.650 209.400 39.450 215.250 ;
        RECT 40.650 209.400 42.450 215.250 ;
        RECT 46.650 209.400 48.450 215.250 ;
        RECT 49.650 210.000 51.450 215.250 ;
        RECT 8.400 198.150 9.600 203.400 ;
        RECT 24.450 202.350 27.000 203.400 ;
        RECT 23.100 198.150 24.900 199.950 ;
        RECT 7.950 196.050 10.050 198.150 ;
        RECT 8.400 189.600 9.600 196.050 ;
        RECT 10.950 194.850 13.050 196.950 ;
        RECT 22.950 196.050 25.050 198.150 ;
        RECT 25.950 195.150 27.000 202.350 ;
        RECT 38.250 201.150 39.450 209.400 ;
        RECT 47.250 209.100 48.450 209.400 ;
        RECT 52.650 209.400 54.450 215.250 ;
        RECT 55.650 209.400 57.450 215.250 ;
        RECT 64.650 209.400 66.450 215.250 ;
        RECT 67.650 209.400 69.450 215.250 ;
        RECT 70.650 209.400 72.450 215.250 ;
        RECT 82.650 209.400 84.450 215.250 ;
        RECT 85.650 209.400 87.450 215.250 ;
        RECT 88.650 209.400 90.450 215.250 ;
        RECT 92.550 209.400 94.350 215.250 ;
        RECT 95.550 209.400 97.350 215.250 ;
        RECT 52.650 209.100 54.300 209.400 ;
        RECT 47.250 208.200 54.300 209.100 ;
        RECT 29.100 198.150 30.900 199.950 ;
        RECT 28.950 196.050 31.050 198.150 ;
        RECT 34.950 197.850 37.050 199.950 ;
        RECT 37.950 199.050 40.050 201.150 ;
        RECT 47.250 199.950 48.300 208.200 ;
        RECT 53.100 204.150 54.900 205.950 ;
        RECT 64.950 204.450 67.050 205.050 ;
        RECT 49.950 201.150 51.750 202.950 ;
        RECT 52.950 202.050 55.050 204.150 ;
        RECT 62.550 203.550 67.050 204.450 ;
        RECT 56.100 201.150 57.900 202.950 ;
        RECT 35.100 196.050 36.900 197.850 ;
        RECT 11.100 193.050 12.900 194.850 ;
        RECT 25.950 193.050 28.050 195.150 ;
        RECT 7.650 183.750 9.450 189.600 ;
        RECT 10.650 183.750 12.450 189.600 ;
        RECT 25.950 186.600 27.000 193.050 ;
        RECT 38.250 191.700 39.450 199.050 ;
        RECT 40.950 197.850 43.050 199.950 ;
        RECT 46.950 197.850 49.050 199.950 ;
        RECT 49.950 199.050 52.050 201.150 ;
        RECT 55.950 199.050 58.050 201.150 ;
        RECT 41.100 196.050 42.900 197.850 ;
        RECT 47.400 193.650 48.600 197.850 ;
        RECT 52.950 195.450 55.050 196.050 ;
        RECT 62.550 195.450 63.450 203.550 ;
        RECT 64.950 202.950 67.050 203.550 ;
        RECT 68.250 201.150 69.450 209.400 ;
        RECT 86.250 201.150 87.450 209.400 ;
        RECT 64.950 197.850 67.050 199.950 ;
        RECT 67.950 199.050 70.050 201.150 ;
        RECT 65.100 196.050 66.900 197.850 ;
        RECT 52.950 194.550 63.450 195.450 ;
        RECT 52.950 193.950 55.050 194.550 ;
        RECT 47.400 192.000 51.900 193.650 ;
        RECT 35.850 190.800 39.450 191.700 ;
        RECT 22.650 183.750 24.450 186.600 ;
        RECT 25.650 183.750 27.450 186.600 ;
        RECT 28.650 183.750 30.450 186.600 ;
        RECT 35.850 183.750 37.650 190.800 ;
        RECT 40.350 183.750 42.150 189.600 ;
        RECT 50.100 183.750 51.900 192.000 ;
        RECT 55.500 183.750 57.300 192.600 ;
        RECT 68.250 191.700 69.450 199.050 ;
        RECT 70.950 197.850 73.050 199.950 ;
        RECT 82.950 197.850 85.050 199.950 ;
        RECT 85.950 199.050 88.050 201.150 ;
        RECT 71.100 196.050 72.900 197.850 ;
        RECT 83.100 196.050 84.900 197.850 ;
        RECT 86.250 191.700 87.450 199.050 ;
        RECT 88.950 197.850 91.050 199.950 ;
        RECT 92.100 198.150 93.900 199.950 ;
        RECT 89.100 196.050 90.900 197.850 ;
        RECT 91.950 196.050 94.050 198.150 ;
        RECT 95.700 192.300 96.900 209.400 ;
        RECT 99.150 203.400 100.950 215.250 ;
        RECT 102.150 203.400 103.950 215.250 ;
        RECT 110.550 209.400 112.350 215.250 ;
        RECT 113.550 209.400 115.350 215.250 ;
        RECT 116.550 210.000 118.350 215.250 ;
        RECT 113.700 209.100 115.350 209.400 ;
        RECT 119.550 209.400 121.350 215.250 ;
        RECT 127.650 209.400 129.450 215.250 ;
        RECT 130.650 209.400 132.450 215.250 ;
        RECT 133.650 209.400 135.450 215.250 ;
        RECT 146.400 209.400 148.200 215.250 ;
        RECT 119.550 209.100 120.750 209.400 ;
        RECT 113.700 208.200 120.750 209.100 ;
        RECT 113.100 204.150 114.900 205.950 ;
        RECT 97.950 197.850 100.050 199.950 ;
        RECT 102.150 198.150 103.350 203.400 ;
        RECT 110.100 201.150 111.900 202.950 ;
        RECT 112.950 202.050 115.050 204.150 ;
        RECT 116.250 201.150 118.050 202.950 ;
        RECT 109.950 199.050 112.050 201.150 ;
        RECT 115.950 199.050 118.050 201.150 ;
        RECT 119.700 199.950 120.750 208.200 ;
        RECT 131.250 201.150 132.450 209.400 ;
        RECT 149.700 203.400 151.500 215.250 ;
        RECT 153.900 203.400 155.700 215.250 ;
        RECT 164.550 209.400 166.350 215.250 ;
        RECT 167.550 209.400 169.350 215.250 ;
        RECT 170.550 210.000 172.350 215.250 ;
        RECT 167.700 209.100 169.350 209.400 ;
        RECT 173.550 209.400 175.350 215.250 ;
        RECT 182.400 209.400 184.200 215.250 ;
        RECT 173.550 209.100 174.750 209.400 ;
        RECT 167.700 208.200 174.750 209.100 ;
        RECT 167.100 204.150 168.900 205.950 ;
        RECT 146.250 201.150 148.050 202.950 ;
        RECT 98.100 196.050 99.900 197.850 ;
        RECT 100.950 196.050 103.350 198.150 ;
        RECT 118.950 197.850 121.050 199.950 ;
        RECT 127.950 197.850 130.050 199.950 ;
        RECT 130.950 199.050 133.050 201.150 ;
        RECT 65.850 190.800 69.450 191.700 ;
        RECT 83.850 190.800 87.450 191.700 ;
        RECT 92.550 191.100 100.050 192.300 ;
        RECT 65.850 183.750 67.650 190.800 ;
        RECT 70.350 183.750 72.150 189.600 ;
        RECT 83.850 183.750 85.650 190.800 ;
        RECT 88.350 183.750 90.150 189.600 ;
        RECT 92.550 183.750 94.350 191.100 ;
        RECT 98.250 190.500 100.050 191.100 ;
        RECT 102.150 189.600 103.350 196.050 ;
        RECT 119.400 193.650 120.600 197.850 ;
        RECT 128.100 196.050 129.900 197.850 ;
        RECT 97.050 183.750 98.850 189.600 ;
        RECT 100.050 188.100 103.350 189.600 ;
        RECT 100.050 183.750 101.850 188.100 ;
        RECT 110.700 183.750 112.500 192.600 ;
        RECT 116.100 192.000 120.600 193.650 ;
        RECT 116.100 183.750 117.900 192.000 ;
        RECT 131.250 191.700 132.450 199.050 ;
        RECT 133.950 197.850 136.050 199.950 ;
        RECT 145.950 199.050 148.050 201.150 ;
        RECT 149.850 198.150 151.050 203.400 ;
        RECT 164.100 201.150 165.900 202.950 ;
        RECT 166.950 202.050 169.050 204.150 ;
        RECT 170.250 201.150 172.050 202.950 ;
        RECT 155.100 198.150 156.900 199.950 ;
        RECT 163.950 199.050 166.050 201.150 ;
        RECT 169.950 199.050 172.050 201.150 ;
        RECT 173.700 199.950 174.750 208.200 ;
        RECT 185.700 203.400 187.500 215.250 ;
        RECT 189.900 203.400 191.700 215.250 ;
        RECT 197.550 209.400 199.350 215.250 ;
        RECT 200.550 209.400 202.350 215.250 ;
        RECT 182.250 201.150 184.050 202.950 ;
        RECT 134.100 196.050 135.900 197.850 ;
        RECT 148.950 196.050 151.050 198.150 ;
        RECT 139.950 195.450 142.050 196.050 ;
        RECT 145.950 195.450 148.050 196.050 ;
        RECT 139.950 194.550 148.050 195.450 ;
        RECT 139.950 193.950 142.050 194.550 ;
        RECT 145.950 193.950 148.050 194.550 ;
        RECT 148.950 192.750 150.150 196.050 ;
        RECT 151.950 194.850 154.050 196.950 ;
        RECT 154.950 196.050 157.050 198.150 ;
        RECT 172.950 197.850 175.050 199.950 ;
        RECT 181.950 199.050 184.050 201.150 ;
        RECT 185.850 198.150 187.050 203.400 ;
        RECT 191.100 198.150 192.900 199.950 ;
        RECT 152.100 193.050 153.900 194.850 ;
        RECT 173.400 193.650 174.600 197.850 ;
        RECT 128.850 190.800 132.450 191.700 ;
        RECT 146.250 191.700 150.000 192.750 ;
        RECT 128.850 183.750 130.650 190.800 ;
        RECT 146.250 189.600 147.450 191.700 ;
        RECT 133.350 183.750 135.150 189.600 ;
        RECT 145.650 183.750 147.450 189.600 ;
        RECT 148.650 188.700 156.450 190.050 ;
        RECT 148.650 183.750 150.450 188.700 ;
        RECT 151.650 183.750 153.450 187.800 ;
        RECT 154.650 183.750 156.450 188.700 ;
        RECT 164.700 183.750 166.500 192.600 ;
        RECT 170.100 192.000 174.600 193.650 ;
        RECT 184.950 196.050 187.050 198.150 ;
        RECT 184.950 192.750 186.150 196.050 ;
        RECT 187.950 194.850 190.050 196.950 ;
        RECT 190.950 196.050 193.050 198.150 ;
        RECT 200.400 196.950 201.600 209.400 ;
        RECT 213.150 203.400 214.950 215.250 ;
        RECT 217.650 203.400 220.950 215.250 ;
        RECT 223.650 203.400 225.450 215.250 ;
        RECT 232.650 209.400 234.450 215.250 ;
        RECT 235.650 209.400 237.450 215.250 ;
        RECT 242.550 209.400 244.350 215.250 ;
        RECT 245.550 209.400 247.350 215.250 ;
        RECT 248.550 210.000 250.350 215.250 ;
        RECT 212.250 198.150 214.050 199.950 ;
        RECT 218.250 198.150 219.450 203.400 ;
        RECT 224.100 198.150 225.900 199.950 ;
        RECT 197.100 195.150 198.900 196.950 ;
        RECT 188.100 193.050 189.900 194.850 ;
        RECT 196.950 193.050 199.050 195.150 ;
        RECT 199.950 194.850 202.050 196.950 ;
        RECT 211.950 196.050 214.050 198.150 ;
        RECT 214.950 194.850 217.050 196.950 ;
        RECT 217.950 196.050 220.050 198.150 ;
        RECT 170.100 183.750 171.900 192.000 ;
        RECT 182.250 191.700 186.000 192.750 ;
        RECT 182.250 189.600 183.450 191.700 ;
        RECT 181.650 183.750 183.450 189.600 ;
        RECT 184.650 188.700 192.450 190.050 ;
        RECT 184.650 183.750 186.450 188.700 ;
        RECT 187.650 183.750 189.450 187.800 ;
        RECT 190.650 183.750 192.450 188.700 ;
        RECT 200.400 186.600 201.600 194.850 ;
        RECT 215.700 193.050 217.500 194.850 ;
        RECT 218.400 192.150 219.600 196.050 ;
        RECT 220.950 194.850 223.050 196.950 ;
        RECT 223.950 196.050 226.050 198.150 ;
        RECT 233.400 196.950 234.600 209.400 ;
        RECT 245.700 209.100 247.350 209.400 ;
        RECT 251.550 209.400 253.350 215.250 ;
        RECT 251.550 209.100 252.750 209.400 ;
        RECT 245.700 208.200 252.750 209.100 ;
        RECT 245.100 204.150 246.900 205.950 ;
        RECT 238.950 199.950 241.050 202.050 ;
        RECT 242.100 201.150 243.900 202.950 ;
        RECT 244.950 202.050 247.050 204.150 ;
        RECT 248.250 201.150 250.050 202.950 ;
        RECT 232.950 194.850 235.050 196.950 ;
        RECT 236.100 195.150 237.900 196.950 ;
        RECT 239.550 195.450 240.450 199.950 ;
        RECT 241.950 199.050 244.050 201.150 ;
        RECT 247.950 199.050 250.050 201.150 ;
        RECT 251.700 199.950 252.750 208.200 ;
        RECT 264.450 203.400 266.250 215.250 ;
        RECT 268.650 203.400 270.450 215.250 ;
        RECT 277.650 209.400 279.450 215.250 ;
        RECT 280.650 209.400 282.450 215.250 ;
        RECT 289.650 209.400 291.450 215.250 ;
        RECT 292.650 209.400 294.450 215.250 ;
        RECT 295.650 209.400 297.450 215.250 ;
        RECT 301.650 209.400 303.450 215.250 ;
        RECT 304.650 210.000 306.450 215.250 ;
        RECT 264.450 202.350 267.000 203.400 ;
        RECT 250.950 197.850 253.050 199.950 ;
        RECT 263.100 198.150 264.900 199.950 ;
        RECT 244.950 195.450 247.050 196.050 ;
        RECT 221.100 193.050 222.900 194.850 ;
        RECT 215.250 191.100 219.600 192.150 ;
        RECT 215.250 189.600 216.150 191.100 ;
        RECT 197.550 183.750 199.350 186.600 ;
        RECT 200.550 183.750 202.350 186.600 ;
        RECT 211.650 184.500 213.450 189.600 ;
        RECT 214.650 185.400 216.450 189.600 ;
        RECT 217.650 189.000 225.450 189.900 ;
        RECT 217.650 184.500 219.450 189.000 ;
        RECT 211.650 183.750 219.450 184.500 ;
        RECT 220.650 183.750 222.450 188.100 ;
        RECT 223.650 183.750 225.450 189.000 ;
        RECT 233.400 186.600 234.600 194.850 ;
        RECT 235.950 193.050 238.050 195.150 ;
        RECT 239.550 194.550 247.050 195.450 ;
        RECT 244.950 193.950 247.050 194.550 ;
        RECT 251.400 193.650 252.600 197.850 ;
        RECT 262.950 196.050 265.050 198.150 ;
        RECT 232.650 183.750 234.450 186.600 ;
        RECT 235.650 183.750 237.450 186.600 ;
        RECT 242.700 183.750 244.500 192.600 ;
        RECT 248.100 192.000 252.600 193.650 ;
        RECT 265.950 195.150 267.000 202.350 ;
        RECT 269.100 198.150 270.900 199.950 ;
        RECT 268.950 196.050 271.050 198.150 ;
        RECT 278.400 196.950 279.600 209.400 ;
        RECT 293.250 201.150 294.450 209.400 ;
        RECT 302.250 209.100 303.450 209.400 ;
        RECT 307.650 209.400 309.450 215.250 ;
        RECT 310.650 209.400 312.450 215.250 ;
        RECT 307.650 209.100 309.300 209.400 ;
        RECT 302.250 208.200 309.300 209.100 ;
        RECT 289.950 197.850 292.050 199.950 ;
        RECT 292.950 199.050 295.050 201.150 ;
        RECT 302.250 199.950 303.300 208.200 ;
        RECT 308.100 204.150 309.900 205.950 ;
        RECT 304.950 201.150 306.750 202.950 ;
        RECT 307.950 202.050 310.050 204.150 ;
        RECT 319.050 203.400 320.850 215.250 ;
        RECT 322.050 203.400 323.850 215.250 ;
        RECT 325.650 209.400 327.450 215.250 ;
        RECT 328.650 209.400 330.450 215.250 ;
        RECT 338.550 209.400 340.350 215.250 ;
        RECT 341.550 209.400 343.350 215.250 ;
        RECT 344.550 210.000 346.350 215.250 ;
        RECT 311.100 201.150 312.900 202.950 ;
        RECT 265.950 193.050 268.050 195.150 ;
        RECT 277.950 194.850 280.050 196.950 ;
        RECT 281.100 195.150 282.900 196.950 ;
        RECT 290.100 196.050 291.900 197.850 ;
        RECT 248.100 183.750 249.900 192.000 ;
        RECT 265.950 186.600 267.000 193.050 ;
        RECT 278.400 186.600 279.600 194.850 ;
        RECT 280.950 193.050 283.050 195.150 ;
        RECT 293.250 191.700 294.450 199.050 ;
        RECT 295.950 197.850 298.050 199.950 ;
        RECT 301.950 197.850 304.050 199.950 ;
        RECT 304.950 199.050 307.050 201.150 ;
        RECT 310.950 199.050 313.050 201.150 ;
        RECT 313.950 199.950 316.050 202.050 ;
        RECT 296.100 196.050 297.900 197.850 ;
        RECT 302.400 193.650 303.600 197.850 ;
        RECT 310.950 195.450 313.050 196.050 ;
        RECT 314.550 195.450 315.450 199.950 ;
        RECT 310.950 194.550 315.450 195.450 ;
        RECT 319.650 198.150 320.850 203.400 ;
        RECT 319.650 196.050 322.050 198.150 ;
        RECT 322.950 197.850 325.050 199.950 ;
        RECT 323.100 196.050 324.900 197.850 ;
        RECT 310.950 193.950 313.050 194.550 ;
        RECT 302.400 192.000 306.900 193.650 ;
        RECT 290.850 190.800 294.450 191.700 ;
        RECT 262.650 183.750 264.450 186.600 ;
        RECT 265.650 183.750 267.450 186.600 ;
        RECT 268.650 183.750 270.450 186.600 ;
        RECT 277.650 183.750 279.450 186.600 ;
        RECT 280.650 183.750 282.450 186.600 ;
        RECT 290.850 183.750 292.650 190.800 ;
        RECT 295.350 183.750 297.150 189.600 ;
        RECT 305.100 183.750 306.900 192.000 ;
        RECT 310.500 183.750 312.300 192.600 ;
        RECT 319.650 189.600 320.850 196.050 ;
        RECT 326.100 192.300 327.300 209.400 ;
        RECT 341.700 209.100 343.350 209.400 ;
        RECT 347.550 209.400 349.350 215.250 ;
        RECT 347.550 209.100 348.750 209.400 ;
        RECT 341.700 208.200 348.750 209.100 ;
        RECT 341.100 204.150 342.900 205.950 ;
        RECT 338.100 201.150 339.900 202.950 ;
        RECT 340.950 202.050 343.050 204.150 ;
        RECT 344.250 201.150 346.050 202.950 ;
        RECT 329.100 198.150 330.900 199.950 ;
        RECT 337.950 199.050 340.050 201.150 ;
        RECT 343.950 199.050 346.050 201.150 ;
        RECT 347.700 199.950 348.750 208.200 ;
        RECT 353.550 204.300 355.350 215.250 ;
        RECT 356.550 205.200 358.350 215.250 ;
        RECT 359.550 204.300 361.350 215.250 ;
        RECT 353.550 203.400 361.350 204.300 ;
        RECT 362.550 203.400 364.350 215.250 ;
        RECT 376.650 214.500 384.450 215.250 ;
        RECT 376.650 203.400 378.450 214.500 ;
        RECT 379.650 203.400 381.450 213.600 ;
        RECT 382.650 204.600 384.450 214.500 ;
        RECT 385.650 205.500 387.450 215.250 ;
        RECT 388.650 204.600 390.450 215.250 ;
        RECT 382.650 203.700 390.450 204.600 ;
        RECT 402.450 203.400 404.250 215.250 ;
        RECT 406.650 203.400 408.450 215.250 ;
        RECT 414.150 204.900 415.950 215.250 ;
        RECT 413.550 203.550 415.950 204.900 ;
        RECT 417.150 203.550 418.950 215.250 ;
        RECT 328.950 196.050 331.050 198.150 ;
        RECT 346.950 197.850 349.050 199.950 ;
        RECT 362.700 198.150 363.900 203.400 ;
        RECT 379.800 202.500 381.600 203.400 ;
        RECT 379.800 201.600 383.850 202.500 ;
        RECT 402.450 202.350 405.000 203.400 ;
        RECT 377.100 198.150 378.900 199.950 ;
        RECT 382.950 198.150 383.850 201.600 ;
        RECT 388.950 198.150 390.750 199.950 ;
        RECT 401.100 198.150 402.900 199.950 ;
        RECT 347.400 193.650 348.600 197.850 ;
        RECT 352.950 194.850 355.050 196.950 ;
        RECT 356.100 195.150 357.900 196.950 ;
        RECT 322.950 191.100 330.450 192.300 ;
        RECT 322.950 190.500 324.750 191.100 ;
        RECT 319.650 188.100 322.950 189.600 ;
        RECT 321.150 183.750 322.950 188.100 ;
        RECT 324.150 183.750 325.950 189.600 ;
        RECT 328.650 183.750 330.450 191.100 ;
        RECT 338.700 183.750 340.500 192.600 ;
        RECT 344.100 192.000 348.600 193.650 ;
        RECT 353.100 193.050 354.900 194.850 ;
        RECT 355.950 193.050 358.050 195.150 ;
        RECT 358.950 194.850 361.050 196.950 ;
        RECT 361.950 196.050 364.050 198.150 ;
        RECT 376.950 196.050 379.050 198.150 ;
        RECT 359.100 193.050 360.900 194.850 ;
        RECT 344.100 183.750 345.900 192.000 ;
        RECT 362.700 189.600 363.900 196.050 ;
        RECT 379.950 194.850 382.050 196.950 ;
        RECT 382.950 196.050 385.050 198.150 ;
        RECT 380.250 193.050 382.050 194.850 ;
        RECT 384.000 189.600 385.050 196.050 ;
        RECT 385.950 194.850 388.050 196.950 ;
        RECT 388.950 196.050 391.050 198.150 ;
        RECT 400.950 196.050 403.050 198.150 ;
        RECT 403.950 195.150 405.000 202.350 ;
        RECT 407.100 198.150 408.900 199.950 ;
        RECT 406.950 196.050 409.050 198.150 ;
        RECT 413.550 196.950 414.900 203.550 ;
        RECT 421.650 203.400 423.450 215.250 ;
        RECT 425.550 203.400 427.350 215.250 ;
        RECT 429.750 203.400 431.550 215.250 ;
        RECT 440.550 209.400 442.350 215.250 ;
        RECT 443.550 209.400 445.350 215.250 ;
        RECT 454.650 214.500 462.450 215.250 ;
        RECT 416.250 202.200 418.050 202.650 ;
        RECT 422.250 202.200 423.450 203.400 ;
        RECT 416.250 201.000 423.450 202.200 ;
        RECT 429.000 202.350 431.550 203.400 ;
        RECT 416.250 200.850 418.050 201.000 ;
        RECT 385.950 193.050 387.750 194.850 ;
        RECT 403.950 193.050 406.050 195.150 ;
        RECT 412.950 194.850 415.050 196.950 ;
        RECT 354.000 183.750 355.800 189.600 ;
        RECT 358.200 187.950 363.900 189.600 ;
        RECT 358.200 183.750 360.000 187.950 ;
        RECT 361.500 183.750 363.300 186.600 ;
        RECT 379.800 183.750 381.600 189.600 ;
        RECT 384.000 183.750 385.800 189.600 ;
        RECT 388.200 183.750 390.000 189.600 ;
        RECT 403.950 186.600 405.000 193.050 ;
        RECT 412.950 189.600 414.000 194.850 ;
        RECT 416.400 192.600 417.300 200.850 ;
        RECT 419.100 198.150 420.900 199.950 ;
        RECT 425.100 198.150 426.900 199.950 ;
        RECT 418.950 196.050 421.050 198.150 ;
        RECT 422.100 195.150 423.900 196.950 ;
        RECT 424.950 196.050 427.050 198.150 ;
        RECT 429.000 195.150 430.050 202.350 ;
        RECT 431.100 198.150 432.900 199.950 ;
        RECT 430.950 196.050 433.050 198.150 ;
        RECT 443.400 196.950 444.600 209.400 ;
        RECT 454.650 203.400 456.450 214.500 ;
        RECT 457.650 203.400 459.450 213.600 ;
        RECT 460.650 204.600 462.450 214.500 ;
        RECT 463.650 205.500 465.450 215.250 ;
        RECT 466.650 204.600 468.450 215.250 ;
        RECT 460.650 203.700 468.450 204.600 ;
        RECT 473.550 204.300 475.350 215.250 ;
        RECT 476.550 205.200 478.350 215.250 ;
        RECT 479.550 204.300 481.350 215.250 ;
        RECT 473.550 203.400 481.350 204.300 ;
        RECT 482.550 203.400 484.350 215.250 ;
        RECT 492.300 203.400 494.100 215.250 ;
        RECT 496.500 203.400 498.300 215.250 ;
        RECT 499.800 209.400 501.600 215.250 ;
        RECT 509.550 209.400 511.350 215.250 ;
        RECT 512.550 209.400 514.350 215.250 ;
        RECT 515.550 210.000 517.350 215.250 ;
        RECT 512.700 209.100 514.350 209.400 ;
        RECT 518.550 209.400 520.350 215.250 ;
        RECT 518.550 209.100 519.750 209.400 ;
        RECT 512.700 208.200 519.750 209.100 ;
        RECT 499.950 207.450 502.050 208.050 ;
        RECT 508.950 207.450 511.050 208.050 ;
        RECT 499.950 206.550 511.050 207.450 ;
        RECT 499.950 205.950 502.050 206.550 ;
        RECT 508.950 205.950 511.050 206.550 ;
        RECT 512.100 204.150 513.900 205.950 ;
        RECT 457.800 202.500 459.600 203.400 ;
        RECT 457.800 201.600 461.850 202.500 ;
        RECT 455.100 198.150 456.900 199.950 ;
        RECT 460.950 198.150 461.850 201.600 ;
        RECT 466.950 198.150 468.750 199.950 ;
        RECT 482.700 198.150 483.900 203.400 ;
        RECT 491.100 198.150 492.900 199.950 ;
        RECT 496.950 198.150 498.150 203.400 ;
        RECT 499.950 201.150 501.750 202.950 ;
        RECT 509.100 201.150 510.900 202.950 ;
        RECT 511.950 202.050 514.050 204.150 ;
        RECT 515.250 201.150 517.050 202.950 ;
        RECT 499.950 199.050 502.050 201.150 ;
        RECT 508.950 199.050 511.050 201.150 ;
        RECT 514.950 199.050 517.050 201.150 ;
        RECT 518.700 199.950 519.750 208.200 ;
        RECT 527.550 205.500 529.350 215.250 ;
        RECT 530.550 206.400 532.350 215.250 ;
        RECT 533.550 214.500 541.350 215.250 ;
        RECT 533.550 205.500 535.350 214.500 ;
        RECT 527.550 204.600 535.350 205.500 ;
        RECT 536.550 205.800 538.350 213.600 ;
        RECT 539.550 206.700 541.350 214.500 ;
        RECT 543.150 214.500 550.950 215.250 ;
        RECT 543.150 205.800 544.950 214.500 ;
        RECT 536.550 204.900 544.950 205.800 ;
        RECT 546.150 205.800 547.950 213.600 ;
        RECT 546.150 203.400 547.350 205.800 ;
        RECT 549.150 205.200 550.950 214.500 ;
        RECT 559.650 209.400 561.450 215.250 ;
        RECT 562.650 210.000 564.450 215.250 ;
        RECT 560.250 209.100 561.450 209.400 ;
        RECT 565.650 209.400 567.450 215.250 ;
        RECT 568.650 209.400 570.450 215.250 ;
        RECT 580.650 209.400 582.450 215.250 ;
        RECT 583.650 209.400 585.450 215.250 ;
        RECT 592.650 209.400 594.450 215.250 ;
        RECT 595.650 209.400 597.450 215.250 ;
        RECT 608.400 209.400 610.200 215.250 ;
        RECT 565.650 209.100 567.300 209.400 ;
        RECT 560.250 208.200 567.300 209.100 ;
        RECT 543.900 202.200 547.350 203.400 ;
        RECT 440.100 195.150 441.900 196.950 ;
        RECT 421.950 193.050 424.050 195.150 ;
        RECT 427.950 193.050 430.050 195.150 ;
        RECT 439.950 193.050 442.050 195.150 ;
        RECT 442.950 194.850 445.050 196.950 ;
        RECT 454.950 196.050 457.050 198.150 ;
        RECT 457.950 194.850 460.050 196.950 ;
        RECT 460.950 196.050 463.050 198.150 ;
        RECT 416.250 191.700 418.050 192.600 ;
        RECT 416.250 190.800 419.550 191.700 ;
        RECT 400.650 183.750 402.450 186.600 ;
        RECT 403.650 183.750 405.450 186.600 ;
        RECT 406.650 183.750 408.450 186.600 ;
        RECT 412.650 183.750 414.450 189.600 ;
        RECT 418.650 186.600 419.550 190.800 ;
        RECT 429.000 186.600 430.050 193.050 ;
        RECT 443.400 186.600 444.600 194.850 ;
        RECT 458.250 193.050 460.050 194.850 ;
        RECT 462.000 189.600 463.050 196.050 ;
        RECT 463.950 194.850 466.050 196.950 ;
        RECT 466.950 196.050 469.050 198.150 ;
        RECT 472.950 194.850 475.050 196.950 ;
        RECT 476.100 195.150 477.900 196.950 ;
        RECT 463.950 193.050 465.750 194.850 ;
        RECT 473.100 193.050 474.900 194.850 ;
        RECT 475.950 193.050 478.050 195.150 ;
        RECT 478.950 194.850 481.050 196.950 ;
        RECT 481.950 196.050 484.050 198.150 ;
        RECT 490.950 196.050 493.050 198.150 ;
        RECT 479.100 193.050 480.900 194.850 ;
        RECT 482.700 189.600 483.900 196.050 ;
        RECT 493.950 194.850 496.050 196.950 ;
        RECT 496.950 196.050 499.050 198.150 ;
        RECT 517.950 197.850 520.050 199.950 ;
        RECT 530.100 198.150 531.900 199.950 ;
        RECT 539.100 198.150 540.900 199.950 ;
        RECT 494.100 193.050 495.900 194.850 ;
        RECT 497.850 192.750 499.050 196.050 ;
        RECT 511.950 195.450 514.050 196.050 ;
        RECT 506.550 194.550 514.050 195.450 ;
        RECT 506.550 193.050 507.450 194.550 ;
        RECT 511.950 193.950 514.050 194.550 ;
        RECT 518.400 193.650 519.600 197.850 ;
        RECT 529.950 196.050 532.050 198.150 ;
        RECT 535.950 194.850 538.050 196.950 ;
        RECT 538.950 196.050 541.050 198.150 ;
        RECT 543.900 196.950 545.100 202.200 ;
        RECT 560.250 199.950 561.300 208.200 ;
        RECT 566.100 204.150 567.900 205.950 ;
        RECT 562.950 201.150 564.750 202.950 ;
        RECT 565.950 202.050 568.050 204.150 ;
        RECT 569.100 201.150 570.900 202.950 ;
        RECT 559.950 197.850 562.050 199.950 ;
        RECT 562.950 199.050 565.050 201.150 ;
        RECT 568.950 199.050 571.050 201.150 ;
        RECT 543.900 194.850 547.050 196.950 ;
        RECT 498.000 191.700 501.750 192.750 ;
        RECT 415.650 183.750 417.450 186.600 ;
        RECT 418.650 183.750 420.450 186.600 ;
        RECT 421.650 183.750 423.450 186.600 ;
        RECT 425.550 183.750 427.350 186.600 ;
        RECT 428.550 183.750 430.350 186.600 ;
        RECT 431.550 183.750 433.350 186.600 ;
        RECT 440.550 183.750 442.350 186.600 ;
        RECT 443.550 183.750 445.350 186.600 ;
        RECT 457.800 183.750 459.600 189.600 ;
        RECT 462.000 183.750 463.800 189.600 ;
        RECT 466.200 183.750 468.000 189.600 ;
        RECT 474.000 183.750 475.800 189.600 ;
        RECT 478.200 187.950 483.900 189.600 ;
        RECT 491.550 188.700 499.350 190.050 ;
        RECT 478.200 183.750 480.000 187.950 ;
        RECT 481.500 183.750 483.300 186.600 ;
        RECT 491.550 183.750 493.350 188.700 ;
        RECT 494.550 183.750 496.350 187.800 ;
        RECT 497.550 183.750 499.350 188.700 ;
        RECT 500.550 189.600 501.750 191.700 ;
        RECT 505.950 190.950 508.050 193.050 ;
        RECT 500.550 183.750 502.350 189.600 ;
        RECT 509.700 183.750 511.500 192.600 ;
        RECT 515.100 192.000 519.600 193.650 ;
        RECT 536.100 193.050 537.900 194.850 ;
        RECT 515.100 183.750 516.900 192.000 ;
        RECT 543.900 188.400 545.100 194.850 ;
        RECT 560.400 193.650 561.600 197.850 ;
        RECT 581.400 196.950 582.600 209.400 ;
        RECT 593.400 196.950 594.600 209.400 ;
        RECT 611.700 203.400 613.500 215.250 ;
        RECT 615.900 203.400 617.700 215.250 ;
        RECT 620.550 209.400 622.350 215.250 ;
        RECT 623.550 209.400 625.350 215.250 ;
        RECT 626.550 210.000 628.350 215.250 ;
        RECT 623.700 209.100 625.350 209.400 ;
        RECT 629.550 209.400 631.350 215.250 ;
        RECT 629.550 209.100 630.750 209.400 ;
        RECT 623.700 208.200 630.750 209.100 ;
        RECT 623.100 204.150 624.900 205.950 ;
        RECT 595.950 201.450 598.050 202.050 ;
        RECT 595.950 200.550 600.450 201.450 ;
        RECT 608.250 201.150 610.050 202.950 ;
        RECT 595.950 199.950 598.050 200.550 ;
        RECT 580.950 194.850 583.050 196.950 ;
        RECT 584.100 195.150 585.900 196.950 ;
        RECT 560.400 192.000 564.900 193.650 ;
        RECT 534.300 187.500 545.100 188.400 ;
        RECT 547.950 189.450 550.050 190.050 ;
        RECT 559.950 189.450 562.050 190.050 ;
        RECT 547.950 188.550 562.050 189.450 ;
        RECT 547.950 187.950 550.050 188.550 ;
        RECT 559.950 187.950 562.050 188.550 ;
        RECT 534.300 186.600 535.350 187.500 ;
        RECT 540.300 186.600 541.350 187.500 ;
        RECT 530.250 183.750 532.350 186.600 ;
        RECT 533.550 183.750 535.350 186.600 ;
        RECT 536.550 183.750 538.350 186.600 ;
        RECT 539.550 183.750 541.350 186.600 ;
        RECT 563.100 183.750 564.900 192.000 ;
        RECT 568.500 183.750 570.300 192.600 ;
        RECT 581.400 186.600 582.600 194.850 ;
        RECT 583.950 193.050 586.050 195.150 ;
        RECT 592.950 194.850 595.050 196.950 ;
        RECT 596.100 195.150 597.900 196.950 ;
        RECT 599.550 196.050 600.450 200.550 ;
        RECT 607.950 199.050 610.050 201.150 ;
        RECT 611.850 198.150 613.050 203.400 ;
        RECT 620.100 201.150 621.900 202.950 ;
        RECT 622.950 202.050 625.050 204.150 ;
        RECT 626.250 201.150 628.050 202.950 ;
        RECT 617.100 198.150 618.900 199.950 ;
        RECT 619.950 199.050 622.050 201.150 ;
        RECT 625.950 199.050 628.050 201.150 ;
        RECT 629.700 199.950 630.750 208.200 ;
        RECT 639.300 203.400 641.100 215.250 ;
        RECT 643.500 203.400 645.300 215.250 ;
        RECT 646.800 209.400 648.600 215.250 ;
        RECT 663.450 203.400 665.250 215.250 ;
        RECT 667.650 203.400 669.450 215.250 ;
        RECT 674.550 203.400 676.350 215.250 ;
        RECT 677.550 203.400 679.350 215.250 ;
        RECT 680.550 203.400 682.350 215.250 ;
        RECT 693.450 203.400 695.250 215.250 ;
        RECT 697.650 203.400 699.450 215.250 ;
        RECT 704.550 209.400 706.350 215.250 ;
        RECT 707.550 209.400 709.350 215.250 ;
        RECT 610.950 196.050 613.050 198.150 ;
        RECT 593.400 186.600 594.600 194.850 ;
        RECT 595.950 193.050 598.050 195.150 ;
        RECT 598.950 193.950 601.050 196.050 ;
        RECT 610.950 192.750 612.150 196.050 ;
        RECT 613.950 194.850 616.050 196.950 ;
        RECT 616.950 196.050 619.050 198.150 ;
        RECT 628.950 197.850 631.050 199.950 ;
        RECT 638.100 198.150 639.900 199.950 ;
        RECT 643.950 198.150 645.150 203.400 ;
        RECT 646.950 201.150 648.750 202.950 ;
        RECT 663.450 202.350 666.000 203.400 ;
        RECT 646.950 199.050 649.050 201.150 ;
        RECT 662.100 198.150 663.900 199.950 ;
        RECT 614.100 193.050 615.900 194.850 ;
        RECT 629.400 193.650 630.600 197.850 ;
        RECT 637.950 196.050 640.050 198.150 ;
        RECT 640.950 194.850 643.050 196.950 ;
        RECT 643.950 196.050 646.050 198.150 ;
        RECT 661.950 196.050 664.050 198.150 ;
        RECT 608.250 191.700 612.000 192.750 ;
        RECT 608.250 189.600 609.450 191.700 ;
        RECT 580.650 183.750 582.450 186.600 ;
        RECT 583.650 183.750 585.450 186.600 ;
        RECT 592.650 183.750 594.450 186.600 ;
        RECT 595.650 183.750 597.450 186.600 ;
        RECT 607.650 183.750 609.450 189.600 ;
        RECT 610.650 188.700 618.450 190.050 ;
        RECT 610.650 183.750 612.450 188.700 ;
        RECT 613.650 183.750 615.450 187.800 ;
        RECT 616.650 183.750 618.450 188.700 ;
        RECT 620.700 183.750 622.500 192.600 ;
        RECT 626.100 192.000 630.600 193.650 ;
        RECT 641.100 193.050 642.900 194.850 ;
        RECT 644.850 192.750 646.050 196.050 ;
        RECT 664.950 195.150 666.000 202.350 ;
        RECT 668.100 198.150 669.900 199.950 ;
        RECT 667.950 196.050 670.050 198.150 ;
        RECT 677.850 196.950 679.200 203.400 ;
        RECT 693.450 202.350 696.000 203.400 ;
        RECT 692.100 198.150 693.900 199.950 ;
        RECT 664.950 193.050 667.050 195.150 ;
        RECT 673.950 194.850 676.050 196.950 ;
        RECT 677.850 194.850 682.050 196.950 ;
        RECT 691.950 196.050 694.050 198.150 ;
        RECT 694.950 195.150 696.000 202.350 ;
        RECT 698.100 198.150 699.900 199.950 ;
        RECT 697.950 196.050 700.050 198.150 ;
        RECT 707.400 196.950 708.600 209.400 ;
        RECT 717.300 203.400 719.100 215.250 ;
        RECT 721.500 203.400 723.300 215.250 ;
        RECT 724.800 209.400 726.600 215.250 ;
        RECT 736.650 209.400 738.450 215.250 ;
        RECT 739.650 210.000 741.450 215.250 ;
        RECT 737.250 209.100 738.450 209.400 ;
        RECT 742.650 209.400 744.450 215.250 ;
        RECT 745.650 209.400 747.450 215.250 ;
        RECT 755.400 209.400 757.200 215.250 ;
        RECT 742.650 209.100 744.300 209.400 ;
        RECT 737.250 208.200 744.300 209.100 ;
        RECT 716.100 198.150 717.900 199.950 ;
        RECT 721.950 198.150 723.150 203.400 ;
        RECT 724.950 201.150 726.750 202.950 ;
        RECT 724.950 199.050 727.050 201.150 ;
        RECT 737.250 199.950 738.300 208.200 ;
        RECT 743.100 204.150 744.900 205.950 ;
        RECT 739.950 201.150 741.750 202.950 ;
        RECT 742.950 202.050 745.050 204.150 ;
        RECT 758.700 203.400 760.500 215.250 ;
        RECT 762.900 203.400 764.700 215.250 ;
        RECT 770.550 203.400 772.350 215.250 ;
        RECT 774.750 203.400 776.550 215.250 ;
        RECT 789.150 204.900 790.950 215.250 ;
        RECT 746.100 201.150 747.900 202.950 ;
        RECT 755.250 201.150 757.050 202.950 ;
        RECT 704.100 195.150 705.900 196.950 ;
        RECT 674.100 193.050 675.900 194.850 ;
        RECT 626.100 183.750 627.900 192.000 ;
        RECT 645.000 191.700 648.750 192.750 ;
        RECT 638.550 188.700 646.350 190.050 ;
        RECT 638.550 183.750 640.350 188.700 ;
        RECT 641.550 183.750 643.350 187.800 ;
        RECT 644.550 183.750 646.350 188.700 ;
        RECT 647.550 189.600 648.750 191.700 ;
        RECT 647.550 183.750 649.350 189.600 ;
        RECT 664.950 186.600 666.000 193.050 ;
        RECT 677.850 189.600 679.200 194.850 ;
        RECT 694.950 193.050 697.050 195.150 ;
        RECT 703.950 193.050 706.050 195.150 ;
        RECT 706.950 194.850 709.050 196.950 ;
        RECT 715.950 196.050 718.050 198.150 ;
        RECT 718.950 194.850 721.050 196.950 ;
        RECT 721.950 196.050 724.050 198.150 ;
        RECT 736.950 197.850 739.050 199.950 ;
        RECT 739.950 199.050 742.050 201.150 ;
        RECT 745.950 199.050 748.050 201.150 ;
        RECT 754.950 199.050 757.050 201.150 ;
        RECT 758.850 198.150 760.050 203.400 ;
        RECT 774.000 202.350 776.550 203.400 ;
        RECT 788.550 203.550 790.950 204.900 ;
        RECT 792.150 203.550 793.950 215.250 ;
        RECT 764.100 198.150 765.900 199.950 ;
        RECT 770.100 198.150 771.900 199.950 ;
        RECT 661.650 183.750 663.450 186.600 ;
        RECT 664.650 183.750 666.450 186.600 ;
        RECT 667.650 183.750 669.450 186.600 ;
        RECT 674.550 183.750 676.350 189.600 ;
        RECT 677.550 183.750 679.350 189.600 ;
        RECT 680.550 183.750 682.350 189.600 ;
        RECT 694.950 186.600 696.000 193.050 ;
        RECT 707.400 186.600 708.600 194.850 ;
        RECT 719.100 193.050 720.900 194.850 ;
        RECT 722.850 192.750 724.050 196.050 ;
        RECT 737.400 193.650 738.600 197.850 ;
        RECT 757.950 196.050 760.050 198.150 ;
        RECT 723.000 191.700 726.750 192.750 ;
        RECT 737.400 192.000 741.900 193.650 ;
        RECT 757.950 192.750 759.150 196.050 ;
        RECT 760.950 194.850 763.050 196.950 ;
        RECT 763.950 196.050 766.050 198.150 ;
        RECT 769.950 196.050 772.050 198.150 ;
        RECT 774.000 195.150 775.050 202.350 ;
        RECT 776.100 198.150 777.900 199.950 ;
        RECT 775.950 196.050 778.050 198.150 ;
        RECT 788.550 196.950 789.900 203.550 ;
        RECT 796.650 203.400 798.450 215.250 ;
        RECT 807.150 204.900 808.950 215.250 ;
        RECT 791.250 202.200 793.050 202.650 ;
        RECT 797.250 202.200 798.450 203.400 ;
        RECT 791.250 201.000 798.450 202.200 ;
        RECT 806.550 203.550 808.950 204.900 ;
        RECT 810.150 203.550 811.950 215.250 ;
        RECT 791.250 200.850 793.050 201.000 ;
        RECT 761.100 193.050 762.900 194.850 ;
        RECT 772.950 193.050 775.050 195.150 ;
        RECT 716.550 188.700 724.350 190.050 ;
        RECT 691.650 183.750 693.450 186.600 ;
        RECT 694.650 183.750 696.450 186.600 ;
        RECT 697.650 183.750 699.450 186.600 ;
        RECT 704.550 183.750 706.350 186.600 ;
        RECT 707.550 183.750 709.350 186.600 ;
        RECT 716.550 183.750 718.350 188.700 ;
        RECT 719.550 183.750 721.350 187.800 ;
        RECT 722.550 183.750 724.350 188.700 ;
        RECT 725.550 189.600 726.750 191.700 ;
        RECT 725.550 183.750 727.350 189.600 ;
        RECT 740.100 183.750 741.900 192.000 ;
        RECT 745.500 183.750 747.300 192.600 ;
        RECT 755.250 191.700 759.000 192.750 ;
        RECT 755.250 189.600 756.450 191.700 ;
        RECT 754.650 183.750 756.450 189.600 ;
        RECT 757.650 188.700 765.450 190.050 ;
        RECT 757.650 183.750 759.450 188.700 ;
        RECT 760.650 183.750 762.450 187.800 ;
        RECT 763.650 183.750 765.450 188.700 ;
        RECT 774.000 186.600 775.050 193.050 ;
        RECT 787.950 194.850 790.050 196.950 ;
        RECT 787.950 189.600 789.000 194.850 ;
        RECT 791.400 192.600 792.300 200.850 ;
        RECT 794.100 198.150 795.900 199.950 ;
        RECT 793.950 196.050 796.050 198.150 ;
        RECT 806.550 196.950 807.900 203.550 ;
        RECT 814.650 203.400 816.450 215.250 ;
        RECT 823.650 209.400 825.450 215.250 ;
        RECT 826.650 210.000 828.450 215.250 ;
        RECT 809.250 202.200 811.050 202.650 ;
        RECT 815.250 202.200 816.450 203.400 ;
        RECT 809.250 201.000 816.450 202.200 ;
        RECT 824.250 209.100 825.450 209.400 ;
        RECT 829.650 209.400 831.450 215.250 ;
        RECT 832.650 209.400 834.450 215.250 ;
        RECT 829.650 209.100 831.300 209.400 ;
        RECT 824.250 208.200 831.300 209.100 ;
        RECT 809.250 200.850 811.050 201.000 ;
        RECT 797.100 195.150 798.900 196.950 ;
        RECT 796.950 193.050 799.050 195.150 ;
        RECT 805.950 194.850 808.050 196.950 ;
        RECT 791.250 191.700 793.050 192.600 ;
        RECT 791.250 190.800 794.550 191.700 ;
        RECT 770.550 183.750 772.350 186.600 ;
        RECT 773.550 183.750 775.350 186.600 ;
        RECT 776.550 183.750 778.350 186.600 ;
        RECT 787.650 183.750 789.450 189.600 ;
        RECT 793.650 186.600 794.550 190.800 ;
        RECT 805.950 189.600 807.000 194.850 ;
        RECT 809.400 192.600 810.300 200.850 ;
        RECT 824.250 199.950 825.300 208.200 ;
        RECT 830.100 204.150 831.900 205.950 ;
        RECT 839.550 204.600 841.350 215.250 ;
        RECT 842.550 205.500 844.350 215.250 ;
        RECT 845.550 214.500 853.350 215.250 ;
        RECT 845.550 204.600 847.350 214.500 ;
        RECT 826.950 201.150 828.750 202.950 ;
        RECT 829.950 202.050 832.050 204.150 ;
        RECT 839.550 203.700 847.350 204.600 ;
        RECT 848.550 203.400 850.350 213.600 ;
        RECT 851.550 203.400 853.350 214.500 ;
        RECT 833.100 201.150 834.900 202.950 ;
        RECT 848.400 202.500 850.200 203.400 ;
        RECT 846.150 201.600 850.200 202.500 ;
        RECT 812.100 198.150 813.900 199.950 ;
        RECT 811.950 196.050 814.050 198.150 ;
        RECT 823.950 197.850 826.050 199.950 ;
        RECT 826.950 199.050 829.050 201.150 ;
        RECT 832.950 199.050 835.050 201.150 ;
        RECT 839.250 198.150 841.050 199.950 ;
        RECT 846.150 198.150 847.050 201.600 ;
        RECT 851.100 198.150 852.900 199.950 ;
        RECT 815.100 195.150 816.900 196.950 ;
        RECT 814.950 193.050 817.050 195.150 ;
        RECT 824.400 193.650 825.600 197.850 ;
        RECT 838.950 196.050 841.050 198.150 ;
        RECT 841.950 194.850 844.050 196.950 ;
        RECT 809.250 191.700 811.050 192.600 ;
        RECT 824.400 192.000 828.900 193.650 ;
        RECT 842.250 193.050 844.050 194.850 ;
        RECT 844.950 196.050 847.050 198.150 ;
        RECT 809.250 190.800 812.550 191.700 ;
        RECT 790.650 183.750 792.450 186.600 ;
        RECT 793.650 183.750 795.450 186.600 ;
        RECT 796.650 183.750 798.450 186.600 ;
        RECT 805.650 183.750 807.450 189.600 ;
        RECT 811.650 186.600 812.550 190.800 ;
        RECT 808.650 183.750 810.450 186.600 ;
        RECT 811.650 183.750 813.450 186.600 ;
        RECT 814.650 183.750 816.450 186.600 ;
        RECT 827.100 183.750 828.900 192.000 ;
        RECT 832.500 183.750 834.300 192.600 ;
        RECT 844.950 189.600 846.000 196.050 ;
        RECT 847.950 194.850 850.050 196.950 ;
        RECT 850.950 196.050 853.050 198.150 ;
        RECT 847.950 193.050 849.750 194.850 ;
        RECT 840.000 183.750 841.800 189.600 ;
        RECT 844.200 183.750 846.000 189.600 ;
        RECT 848.400 183.750 850.200 189.600 ;
        RECT 8.850 172.200 10.650 179.250 ;
        RECT 13.350 173.400 15.150 179.250 ;
        RECT 25.650 176.400 27.450 179.250 ;
        RECT 28.650 176.400 30.450 179.250 ;
        RECT 8.850 171.300 12.450 172.200 ;
        RECT 8.100 165.150 9.900 166.950 ;
        RECT 7.950 163.050 10.050 165.150 ;
        RECT 11.250 163.950 12.450 171.300 ;
        RECT 26.400 168.150 27.600 176.400 ;
        RECT 39.000 173.400 40.800 179.250 ;
        RECT 43.200 175.050 45.000 179.250 ;
        RECT 46.500 176.400 48.300 179.250 ;
        RECT 43.200 173.400 48.900 175.050 ;
        RECT 14.100 165.150 15.900 166.950 ;
        RECT 25.950 166.050 28.050 168.150 ;
        RECT 28.950 167.850 31.050 169.950 ;
        RECT 38.100 168.150 39.900 169.950 ;
        RECT 29.100 166.050 30.900 167.850 ;
        RECT 37.950 166.050 40.050 168.150 ;
        RECT 40.950 167.850 43.050 169.950 ;
        RECT 44.100 168.150 45.900 169.950 ;
        RECT 41.100 166.050 42.900 167.850 ;
        RECT 43.950 166.050 46.050 168.150 ;
        RECT 47.700 166.950 48.900 173.400 ;
        RECT 62.100 171.000 63.900 179.250 ;
        RECT 59.400 169.350 63.900 171.000 ;
        RECT 67.500 170.400 69.300 179.250 ;
        RECT 74.700 176.400 76.500 179.250 ;
        RECT 78.000 175.050 79.800 179.250 ;
        RECT 74.100 173.400 79.800 175.050 ;
        RECT 82.200 173.400 84.000 179.250 ;
        RECT 10.950 161.850 13.050 163.950 ;
        RECT 13.950 163.050 16.050 165.150 ;
        RECT 11.250 153.600 12.450 161.850 ;
        RECT 26.400 153.600 27.600 166.050 ;
        RECT 46.950 164.850 49.050 166.950 ;
        RECT 59.400 165.150 60.600 169.350 ;
        RECT 67.950 168.450 70.050 169.050 ;
        RECT 65.550 167.550 70.050 168.450 ;
        RECT 65.550 166.050 66.450 167.550 ;
        RECT 67.950 166.950 70.050 167.550 ;
        RECT 74.100 166.950 75.300 173.400 ;
        RECT 98.100 171.000 99.900 179.250 ;
        RECT 77.100 168.150 78.900 169.950 ;
        RECT 47.700 159.600 48.900 164.850 ;
        RECT 58.950 163.050 61.050 165.150 ;
        RECT 64.950 163.950 67.050 166.050 ;
        RECT 73.950 164.850 76.050 166.950 ;
        RECT 76.950 166.050 79.050 168.150 ;
        RECT 79.950 167.850 82.050 169.950 ;
        RECT 83.100 168.150 84.900 169.950 ;
        RECT 95.400 169.350 99.900 171.000 ;
        RECT 103.500 170.400 105.300 179.250 ;
        RECT 107.700 170.400 109.500 179.250 ;
        RECT 113.100 171.000 114.900 179.250 ;
        RECT 125.850 173.400 127.650 179.250 ;
        RECT 130.350 172.200 132.150 179.250 ;
        RECT 128.550 171.300 132.150 172.200 ;
        RECT 113.100 169.350 117.600 171.000 ;
        RECT 80.100 166.050 81.900 167.850 ;
        RECT 82.950 166.050 85.050 168.150 ;
        RECT 95.400 165.150 96.600 169.350 ;
        RECT 116.400 165.150 117.600 169.350 ;
        RECT 125.100 165.150 126.900 166.950 ;
        RECT 38.550 158.700 46.350 159.600 ;
        RECT 7.650 147.750 9.450 153.600 ;
        RECT 10.650 147.750 12.450 153.600 ;
        RECT 13.650 147.750 15.450 153.600 ;
        RECT 25.650 147.750 27.450 153.600 ;
        RECT 28.650 147.750 30.450 153.600 ;
        RECT 38.550 147.750 40.350 158.700 ;
        RECT 41.550 147.750 43.350 157.800 ;
        RECT 44.550 147.750 46.350 158.700 ;
        RECT 47.550 147.750 49.350 159.600 ;
        RECT 59.250 154.800 60.300 163.050 ;
        RECT 61.950 161.850 64.050 163.950 ;
        RECT 67.950 161.850 70.050 163.950 ;
        RECT 61.950 160.050 63.750 161.850 ;
        RECT 64.950 158.850 67.050 160.950 ;
        RECT 68.100 160.050 69.900 161.850 ;
        RECT 74.100 159.600 75.300 164.850 ;
        RECT 94.950 163.050 97.050 165.150 ;
        RECT 65.100 157.050 66.900 158.850 ;
        RECT 59.250 153.900 66.300 154.800 ;
        RECT 59.250 153.600 60.450 153.900 ;
        RECT 58.650 147.750 60.450 153.600 ;
        RECT 64.650 153.600 66.300 153.900 ;
        RECT 61.650 147.750 63.450 153.000 ;
        RECT 64.650 147.750 66.450 153.600 ;
        RECT 67.650 147.750 69.450 153.600 ;
        RECT 73.650 147.750 75.450 159.600 ;
        RECT 76.650 158.700 84.450 159.600 ;
        RECT 76.650 147.750 78.450 158.700 ;
        RECT 79.650 147.750 81.450 157.800 ;
        RECT 82.650 147.750 84.450 158.700 ;
        RECT 95.250 154.800 96.300 163.050 ;
        RECT 97.950 161.850 100.050 163.950 ;
        RECT 103.950 161.850 106.050 163.950 ;
        RECT 106.950 161.850 109.050 163.950 ;
        RECT 112.950 161.850 115.050 163.950 ;
        RECT 115.950 163.050 118.050 165.150 ;
        RECT 124.950 163.050 127.050 165.150 ;
        RECT 128.550 163.950 129.750 171.300 ;
        RECT 137.700 170.400 139.500 179.250 ;
        RECT 143.100 171.000 144.900 179.250 ;
        RECT 145.950 174.450 148.050 175.050 ;
        RECT 145.950 173.550 150.450 174.450 ;
        RECT 145.950 172.950 148.050 173.550 ;
        RECT 143.100 169.350 147.600 171.000 ;
        RECT 131.100 165.150 132.900 166.950 ;
        RECT 146.400 165.150 147.600 169.350 ;
        RECT 97.950 160.050 99.750 161.850 ;
        RECT 100.950 158.850 103.050 160.950 ;
        RECT 104.100 160.050 105.900 161.850 ;
        RECT 107.100 160.050 108.900 161.850 ;
        RECT 109.950 158.850 112.050 160.950 ;
        RECT 113.250 160.050 115.050 161.850 ;
        RECT 101.100 157.050 102.900 158.850 ;
        RECT 110.100 157.050 111.900 158.850 ;
        RECT 116.700 154.800 117.750 163.050 ;
        RECT 127.950 161.850 130.050 163.950 ;
        RECT 130.950 163.050 133.050 165.150 ;
        RECT 136.950 161.850 139.050 163.950 ;
        RECT 142.950 161.850 145.050 163.950 ;
        RECT 145.950 163.050 148.050 165.150 ;
        RECT 95.250 153.900 102.300 154.800 ;
        RECT 95.250 153.600 96.450 153.900 ;
        RECT 94.650 147.750 96.450 153.600 ;
        RECT 100.650 153.600 102.300 153.900 ;
        RECT 110.700 153.900 117.750 154.800 ;
        RECT 110.700 153.600 112.350 153.900 ;
        RECT 97.650 147.750 99.450 153.000 ;
        RECT 100.650 147.750 102.450 153.600 ;
        RECT 103.650 147.750 105.450 153.600 ;
        RECT 107.550 147.750 109.350 153.600 ;
        RECT 110.550 147.750 112.350 153.600 ;
        RECT 116.550 153.600 117.750 153.900 ;
        RECT 128.550 153.600 129.750 161.850 ;
        RECT 137.100 160.050 138.900 161.850 ;
        RECT 139.950 158.850 142.050 160.950 ;
        RECT 143.250 160.050 145.050 161.850 ;
        RECT 140.100 157.050 141.900 158.850 ;
        RECT 146.700 154.800 147.750 163.050 ;
        RECT 149.550 162.450 150.450 173.550 ;
        RECT 153.000 173.400 154.800 179.250 ;
        RECT 157.200 175.050 159.000 179.250 ;
        RECT 160.500 176.400 162.300 179.250 ;
        RECT 157.200 173.400 162.900 175.050 ;
        RECT 152.100 168.150 153.900 169.950 ;
        RECT 151.950 166.050 154.050 168.150 ;
        RECT 154.950 167.850 157.050 169.950 ;
        RECT 158.100 168.150 159.900 169.950 ;
        RECT 155.100 166.050 156.900 167.850 ;
        RECT 157.950 166.050 160.050 168.150 ;
        RECT 161.700 166.950 162.900 173.400 ;
        RECT 173.550 174.300 175.350 179.250 ;
        RECT 176.550 175.200 178.350 179.250 ;
        RECT 179.550 174.300 181.350 179.250 ;
        RECT 173.550 172.950 181.350 174.300 ;
        RECT 182.550 173.400 184.350 179.250 ;
        RECT 189.000 173.400 190.800 179.250 ;
        RECT 193.200 175.050 195.000 179.250 ;
        RECT 196.500 176.400 198.300 179.250 ;
        RECT 193.200 173.400 198.900 175.050 ;
        RECT 182.550 171.300 183.750 173.400 ;
        RECT 180.000 170.250 183.750 171.300 ;
        RECT 166.950 166.950 169.050 169.050 ;
        RECT 176.100 168.150 177.900 169.950 ;
        RECT 160.950 164.850 163.050 166.950 ;
        RECT 167.550 165.450 168.450 166.950 ;
        RECT 169.950 165.450 172.050 166.050 ;
        RECT 154.950 162.450 157.050 163.050 ;
        RECT 149.550 161.550 157.050 162.450 ;
        RECT 154.950 160.950 157.050 161.550 ;
        RECT 161.700 159.600 162.900 164.850 ;
        RECT 167.550 164.550 172.050 165.450 ;
        RECT 172.950 164.850 175.050 166.950 ;
        RECT 175.950 166.050 178.050 168.150 ;
        RECT 179.850 166.950 181.050 170.250 ;
        RECT 188.100 168.150 189.900 169.950 ;
        RECT 178.950 164.850 181.050 166.950 ;
        RECT 187.950 166.050 190.050 168.150 ;
        RECT 190.950 167.850 193.050 169.950 ;
        RECT 194.100 168.150 195.900 169.950 ;
        RECT 191.100 166.050 192.900 167.850 ;
        RECT 193.950 166.050 196.050 168.150 ;
        RECT 197.700 166.950 198.900 173.400 ;
        RECT 203.550 174.300 205.350 179.250 ;
        RECT 206.550 175.200 208.350 179.250 ;
        RECT 209.550 174.300 211.350 179.250 ;
        RECT 203.550 172.950 211.350 174.300 ;
        RECT 212.550 173.400 214.350 179.250 ;
        RECT 220.650 176.400 222.450 179.250 ;
        RECT 223.650 176.400 225.450 179.250 ;
        RECT 226.650 176.400 228.450 179.250 ;
        RECT 233.550 176.400 235.350 179.250 ;
        RECT 236.550 176.400 238.350 179.250 ;
        RECT 212.550 171.300 213.750 173.400 ;
        RECT 210.000 170.250 213.750 171.300 ;
        RECT 206.100 168.150 207.900 169.950 ;
        RECT 196.950 164.850 199.050 166.950 ;
        RECT 202.950 164.850 205.050 166.950 ;
        RECT 205.950 166.050 208.050 168.150 ;
        RECT 209.850 166.950 211.050 170.250 ;
        RECT 223.950 169.950 225.000 176.400 ;
        RECT 223.950 167.850 226.050 169.950 ;
        RECT 232.950 167.850 235.050 169.950 ;
        RECT 236.400 168.150 237.600 176.400 ;
        RECT 248.850 172.200 250.650 179.250 ;
        RECT 253.350 173.400 255.150 179.250 ;
        RECT 262.650 176.400 264.450 179.250 ;
        RECT 265.650 176.400 267.450 179.250 ;
        RECT 268.650 176.400 270.450 179.250 ;
        RECT 248.850 171.300 252.450 172.200 ;
        RECT 208.950 164.850 211.050 166.950 ;
        RECT 220.950 164.850 223.050 166.950 ;
        RECT 169.950 163.950 172.050 164.550 ;
        RECT 173.100 163.050 174.900 164.850 ;
        RECT 178.950 159.600 180.150 164.850 ;
        RECT 181.950 161.850 184.050 163.950 ;
        RECT 181.950 160.050 183.750 161.850 ;
        RECT 197.700 159.600 198.900 164.850 ;
        RECT 203.100 163.050 204.900 164.850 ;
        RECT 208.950 159.600 210.150 164.850 ;
        RECT 211.950 161.850 214.050 163.950 ;
        RECT 221.100 163.050 222.900 164.850 ;
        RECT 211.950 160.050 213.750 161.850 ;
        RECT 223.950 160.650 225.000 167.850 ;
        RECT 226.950 164.850 229.050 166.950 ;
        RECT 233.100 166.050 234.900 167.850 ;
        RECT 235.950 166.050 238.050 168.150 ;
        RECT 227.100 163.050 228.900 164.850 ;
        RECT 222.450 159.600 225.000 160.650 ;
        RECT 140.700 153.900 147.750 154.800 ;
        RECT 140.700 153.600 142.350 153.900 ;
        RECT 113.550 147.750 115.350 153.000 ;
        RECT 116.550 147.750 118.350 153.600 ;
        RECT 125.550 147.750 127.350 153.600 ;
        RECT 128.550 147.750 130.350 153.600 ;
        RECT 131.550 147.750 133.350 153.600 ;
        RECT 137.550 147.750 139.350 153.600 ;
        RECT 140.550 147.750 142.350 153.600 ;
        RECT 146.550 153.600 147.750 153.900 ;
        RECT 152.550 158.700 160.350 159.600 ;
        RECT 143.550 147.750 145.350 153.000 ;
        RECT 146.550 147.750 148.350 153.600 ;
        RECT 152.550 147.750 154.350 158.700 ;
        RECT 155.550 147.750 157.350 157.800 ;
        RECT 158.550 147.750 160.350 158.700 ;
        RECT 161.550 147.750 163.350 159.600 ;
        RECT 174.300 147.750 176.100 159.600 ;
        RECT 178.500 147.750 180.300 159.600 ;
        RECT 188.550 158.700 196.350 159.600 ;
        RECT 181.800 147.750 183.600 153.600 ;
        RECT 188.550 147.750 190.350 158.700 ;
        RECT 191.550 147.750 193.350 157.800 ;
        RECT 194.550 147.750 196.350 158.700 ;
        RECT 197.550 147.750 199.350 159.600 ;
        RECT 204.300 147.750 206.100 159.600 ;
        RECT 208.500 147.750 210.300 159.600 ;
        RECT 211.800 147.750 213.600 153.600 ;
        RECT 222.450 147.750 224.250 159.600 ;
        RECT 226.650 147.750 228.450 159.600 ;
        RECT 236.400 153.600 237.600 166.050 ;
        RECT 248.100 165.150 249.900 166.950 ;
        RECT 247.950 163.050 250.050 165.150 ;
        RECT 251.250 163.950 252.450 171.300 ;
        RECT 265.950 169.950 267.000 176.400 ;
        RECT 275.850 173.400 277.650 179.250 ;
        RECT 280.350 172.200 282.150 179.250 ;
        RECT 293.550 174.300 295.350 179.250 ;
        RECT 296.550 175.200 298.350 179.250 ;
        RECT 299.550 174.300 301.350 179.250 ;
        RECT 293.550 172.950 301.350 174.300 ;
        RECT 302.550 173.400 304.350 179.250 ;
        RECT 278.550 171.300 282.150 172.200 ;
        RECT 302.550 171.300 303.750 173.400 ;
        RECT 314.850 172.200 316.650 179.250 ;
        RECT 319.350 173.400 321.150 179.250 ;
        RECT 326.550 176.400 328.350 179.250 ;
        RECT 329.550 176.400 331.350 179.250 ;
        RECT 314.850 171.300 318.450 172.200 ;
        RECT 265.950 167.850 268.050 169.950 ;
        RECT 254.100 165.150 255.900 166.950 ;
        RECT 250.950 161.850 253.050 163.950 ;
        RECT 253.950 163.050 256.050 165.150 ;
        RECT 262.950 164.850 265.050 166.950 ;
        RECT 263.100 163.050 264.900 164.850 ;
        RECT 251.250 153.600 252.450 161.850 ;
        RECT 265.950 160.650 267.000 167.850 ;
        RECT 268.950 164.850 271.050 166.950 ;
        RECT 275.100 165.150 276.900 166.950 ;
        RECT 269.100 163.050 270.900 164.850 ;
        RECT 274.950 163.050 277.050 165.150 ;
        RECT 278.550 163.950 279.750 171.300 ;
        RECT 300.000 170.250 303.750 171.300 ;
        RECT 296.100 168.150 297.900 169.950 ;
        RECT 281.100 165.150 282.900 166.950 ;
        RECT 277.950 161.850 280.050 163.950 ;
        RECT 280.950 163.050 283.050 165.150 ;
        RECT 292.950 164.850 295.050 166.950 ;
        RECT 295.950 166.050 298.050 168.150 ;
        RECT 299.850 166.950 301.050 170.250 ;
        RECT 298.950 164.850 301.050 166.950 ;
        RECT 314.100 165.150 315.900 166.950 ;
        RECT 293.100 163.050 294.900 164.850 ;
        RECT 264.450 159.600 267.000 160.650 ;
        RECT 233.550 147.750 235.350 153.600 ;
        RECT 236.550 147.750 238.350 153.600 ;
        RECT 247.650 147.750 249.450 153.600 ;
        RECT 250.650 147.750 252.450 153.600 ;
        RECT 253.650 147.750 255.450 153.600 ;
        RECT 264.450 147.750 266.250 159.600 ;
        RECT 268.650 147.750 270.450 159.600 ;
        RECT 278.550 153.600 279.750 161.850 ;
        RECT 298.950 159.600 300.150 164.850 ;
        RECT 301.950 161.850 304.050 163.950 ;
        RECT 313.950 163.050 316.050 165.150 ;
        RECT 317.250 163.950 318.450 171.300 ;
        RECT 319.950 171.450 322.050 172.050 ;
        RECT 319.950 170.550 324.450 171.450 ;
        RECT 319.950 169.950 322.050 170.550 ;
        RECT 320.100 165.150 321.900 166.950 ;
        RECT 316.950 161.850 319.050 163.950 ;
        RECT 319.950 163.050 322.050 165.150 ;
        RECT 323.550 162.450 324.450 170.550 ;
        RECT 325.950 167.850 328.050 169.950 ;
        RECT 329.400 168.150 330.600 176.400 ;
        RECT 334.950 172.950 337.050 175.050 ;
        RECT 339.000 173.400 340.800 179.250 ;
        RECT 343.200 175.050 345.000 179.250 ;
        RECT 346.500 176.400 348.300 179.250 ;
        RECT 343.200 173.400 348.900 175.050 ;
        RECT 326.100 166.050 327.900 167.850 ;
        RECT 328.950 166.050 331.050 168.150 ;
        RECT 325.950 162.450 328.050 163.050 ;
        RECT 301.950 160.050 303.750 161.850 ;
        RECT 275.550 147.750 277.350 153.600 ;
        RECT 278.550 147.750 280.350 153.600 ;
        RECT 281.550 147.750 283.350 153.600 ;
        RECT 294.300 147.750 296.100 159.600 ;
        RECT 298.500 147.750 300.300 159.600 ;
        RECT 317.250 153.600 318.450 161.850 ;
        RECT 323.550 161.550 328.050 162.450 ;
        RECT 325.950 160.950 328.050 161.550 ;
        RECT 319.950 157.950 322.050 160.050 ;
        RECT 320.550 156.450 321.450 157.950 ;
        RECT 325.950 156.450 328.050 157.050 ;
        RECT 320.550 155.550 328.050 156.450 ;
        RECT 325.950 154.950 328.050 155.550 ;
        RECT 329.400 153.600 330.600 166.050 ;
        RECT 331.950 162.450 334.050 163.050 ;
        RECT 335.550 162.450 336.450 172.950 ;
        RECT 338.100 168.150 339.900 169.950 ;
        RECT 337.950 166.050 340.050 168.150 ;
        RECT 340.950 167.850 343.050 169.950 ;
        RECT 344.100 168.150 345.900 169.950 ;
        RECT 341.100 166.050 342.900 167.850 ;
        RECT 343.950 166.050 346.050 168.150 ;
        RECT 347.700 166.950 348.900 173.400 ;
        RECT 362.100 171.000 363.900 179.250 ;
        RECT 359.400 169.350 363.900 171.000 ;
        RECT 367.500 170.400 369.300 179.250 ;
        RECT 376.800 173.400 378.600 179.250 ;
        RECT 381.000 173.400 382.800 179.250 ;
        RECT 385.200 173.400 387.000 179.250 ;
        RECT 346.950 164.850 349.050 166.950 ;
        RECT 359.400 165.150 360.600 169.350 ;
        RECT 377.250 168.150 379.050 169.950 ;
        RECT 331.950 161.550 336.450 162.450 ;
        RECT 331.950 160.950 334.050 161.550 ;
        RECT 347.700 159.600 348.900 164.850 ;
        RECT 358.950 163.050 361.050 165.150 ;
        RECT 373.950 164.850 376.050 166.950 ;
        RECT 376.950 166.050 379.050 168.150 ;
        RECT 381.000 166.950 382.050 173.400 ;
        RECT 398.850 172.200 400.650 179.250 ;
        RECT 403.350 173.400 405.150 179.250 ;
        RECT 415.650 173.400 417.450 179.250 ;
        RECT 398.850 171.300 402.450 172.200 ;
        RECT 379.950 164.850 382.050 166.950 ;
        RECT 382.950 168.150 384.750 169.950 ;
        RECT 382.950 166.050 385.050 168.150 ;
        RECT 385.950 164.850 388.050 166.950 ;
        RECT 398.100 165.150 399.900 166.950 ;
        RECT 338.550 158.700 346.350 159.600 ;
        RECT 301.800 147.750 303.600 153.600 ;
        RECT 313.650 147.750 315.450 153.600 ;
        RECT 316.650 147.750 318.450 153.600 ;
        RECT 319.650 147.750 321.450 153.600 ;
        RECT 326.550 147.750 328.350 153.600 ;
        RECT 329.550 147.750 331.350 153.600 ;
        RECT 338.550 147.750 340.350 158.700 ;
        RECT 341.550 147.750 343.350 157.800 ;
        RECT 344.550 147.750 346.350 158.700 ;
        RECT 347.550 147.750 349.350 159.600 ;
        RECT 359.250 154.800 360.300 163.050 ;
        RECT 361.950 161.850 364.050 163.950 ;
        RECT 367.950 161.850 370.050 163.950 ;
        RECT 374.100 163.050 375.900 164.850 ;
        RECT 361.950 160.050 363.750 161.850 ;
        RECT 364.950 158.850 367.050 160.950 ;
        RECT 368.100 160.050 369.900 161.850 ;
        RECT 379.950 161.400 380.850 164.850 ;
        RECT 385.950 163.050 387.750 164.850 ;
        RECT 397.950 163.050 400.050 165.150 ;
        RECT 401.250 163.950 402.450 171.300 ;
        RECT 403.950 171.450 406.050 172.050 ;
        RECT 403.950 170.550 408.450 171.450 ;
        RECT 403.950 169.950 406.050 170.550 ;
        RECT 404.100 165.150 405.900 166.950 ;
        RECT 400.950 161.850 403.050 163.950 ;
        RECT 403.950 163.050 406.050 165.150 ;
        RECT 407.550 163.050 408.450 170.550 ;
        RECT 416.250 171.300 417.450 173.400 ;
        RECT 418.650 174.300 420.450 179.250 ;
        RECT 421.650 175.200 423.450 179.250 ;
        RECT 424.650 174.300 426.450 179.250 ;
        RECT 418.650 172.950 426.450 174.300 ;
        RECT 433.650 178.500 441.450 179.250 ;
        RECT 433.650 173.400 435.450 178.500 ;
        RECT 436.650 173.400 438.450 177.600 ;
        RECT 439.650 174.000 441.450 178.500 ;
        RECT 442.650 174.900 444.450 179.250 ;
        RECT 445.650 174.000 447.450 179.250 ;
        RECT 424.950 171.450 427.050 172.050 ;
        RECT 433.950 171.450 436.050 172.050 ;
        RECT 416.250 170.250 420.000 171.300 ;
        RECT 424.950 170.550 429.450 171.450 ;
        RECT 418.950 166.950 420.150 170.250 ;
        RECT 424.950 169.950 427.050 170.550 ;
        RECT 422.100 168.150 423.900 169.950 ;
        RECT 418.950 164.850 421.050 166.950 ;
        RECT 421.950 166.050 424.050 168.150 ;
        RECT 424.950 164.850 427.050 166.950 ;
        RECT 376.800 160.500 380.850 161.400 ;
        RECT 376.800 159.600 378.600 160.500 ;
        RECT 365.100 157.050 366.900 158.850 ;
        RECT 359.250 153.900 366.300 154.800 ;
        RECT 359.250 153.600 360.450 153.900 ;
        RECT 358.650 147.750 360.450 153.600 ;
        RECT 364.650 153.600 366.300 153.900 ;
        RECT 361.650 147.750 363.450 153.000 ;
        RECT 364.650 147.750 366.450 153.600 ;
        RECT 367.650 147.750 369.450 153.600 ;
        RECT 373.650 148.500 375.450 159.600 ;
        RECT 376.650 149.400 378.450 159.600 ;
        RECT 379.650 158.400 387.450 159.300 ;
        RECT 379.650 148.500 381.450 158.400 ;
        RECT 373.650 147.750 381.450 148.500 ;
        RECT 382.650 147.750 384.450 157.500 ;
        RECT 385.650 147.750 387.450 158.400 ;
        RECT 401.250 153.600 402.450 161.850 ;
        RECT 406.950 160.950 409.050 163.050 ;
        RECT 415.950 161.850 418.050 163.950 ;
        RECT 416.250 160.050 418.050 161.850 ;
        RECT 419.850 159.600 421.050 164.850 ;
        RECT 425.100 163.050 426.900 164.850 ;
        RECT 397.650 147.750 399.450 153.600 ;
        RECT 400.650 147.750 402.450 153.600 ;
        RECT 403.650 147.750 405.450 153.600 ;
        RECT 416.400 147.750 418.200 153.600 ;
        RECT 419.700 147.750 421.500 159.600 ;
        RECT 423.900 147.750 425.700 159.600 ;
        RECT 428.550 156.450 429.450 170.550 ;
        RECT 431.550 170.550 436.050 171.450 ;
        RECT 437.250 171.900 438.150 173.400 ;
        RECT 439.650 173.100 447.450 174.000 ;
        RECT 452.550 174.300 454.350 179.250 ;
        RECT 455.550 175.200 457.350 179.250 ;
        RECT 458.550 174.300 460.350 179.250 ;
        RECT 452.550 172.950 460.350 174.300 ;
        RECT 461.550 173.400 463.350 179.250 ;
        RECT 437.250 170.850 441.600 171.900 ;
        RECT 461.550 171.300 462.750 173.400 ;
        RECT 431.550 160.050 432.450 170.550 ;
        RECT 433.950 169.950 436.050 170.550 ;
        RECT 437.700 168.150 439.500 169.950 ;
        RECT 433.950 164.850 436.050 166.950 ;
        RECT 436.950 166.050 439.050 168.150 ;
        RECT 440.400 166.950 441.600 170.850 ;
        RECT 459.000 170.250 462.750 171.300 ;
        RECT 467.700 170.400 469.500 179.250 ;
        RECT 473.100 171.000 474.900 179.250 ;
        RECT 488.550 171.900 490.350 179.250 ;
        RECT 493.050 173.400 494.850 179.250 ;
        RECT 496.050 174.900 497.850 179.250 ;
        RECT 496.050 173.400 499.350 174.900 ;
        RECT 494.250 171.900 496.050 172.500 ;
        RECT 443.100 168.150 444.900 169.950 ;
        RECT 455.100 168.150 456.900 169.950 ;
        RECT 439.950 164.850 442.050 166.950 ;
        RECT 442.950 166.050 445.050 168.150 ;
        RECT 445.950 164.850 448.050 166.950 ;
        RECT 451.950 164.850 454.050 166.950 ;
        RECT 454.950 166.050 457.050 168.150 ;
        RECT 458.850 166.950 460.050 170.250 ;
        RECT 473.100 169.350 477.600 171.000 ;
        RECT 488.550 170.700 496.050 171.900 ;
        RECT 457.950 164.850 460.050 166.950 ;
        RECT 476.400 165.150 477.600 169.350 ;
        RECT 434.250 163.050 436.050 164.850 ;
        RECT 430.950 157.950 433.050 160.050 ;
        RECT 440.250 159.600 441.450 164.850 ;
        RECT 446.100 163.050 447.900 164.850 ;
        RECT 452.100 163.050 453.900 164.850 ;
        RECT 457.950 159.600 459.150 164.850 ;
        RECT 460.950 161.850 463.050 163.950 ;
        RECT 466.950 161.850 469.050 163.950 ;
        RECT 472.950 161.850 475.050 163.950 ;
        RECT 475.950 163.050 478.050 165.150 ;
        RECT 487.950 164.850 490.050 166.950 ;
        RECT 488.100 163.050 489.900 164.850 ;
        RECT 460.950 160.050 462.750 161.850 ;
        RECT 467.100 160.050 468.900 161.850 ;
        RECT 430.950 156.450 433.050 157.050 ;
        RECT 428.550 155.550 433.050 156.450 ;
        RECT 430.950 154.950 433.050 155.550 ;
        RECT 435.150 147.750 436.950 159.600 ;
        RECT 439.650 147.750 442.950 159.600 ;
        RECT 445.650 147.750 447.450 159.600 ;
        RECT 453.300 147.750 455.100 159.600 ;
        RECT 457.500 147.750 459.300 159.600 ;
        RECT 469.950 158.850 472.050 160.950 ;
        RECT 473.250 160.050 475.050 161.850 ;
        RECT 470.100 157.050 471.900 158.850 ;
        RECT 476.700 154.800 477.750 163.050 ;
        RECT 470.700 153.900 477.750 154.800 ;
        RECT 470.700 153.600 472.350 153.900 ;
        RECT 460.800 147.750 462.600 153.600 ;
        RECT 467.550 147.750 469.350 153.600 ;
        RECT 470.550 147.750 472.350 153.600 ;
        RECT 476.550 153.600 477.750 153.900 ;
        RECT 491.700 153.600 492.900 170.700 ;
        RECT 498.150 166.950 499.350 173.400 ;
        RECT 506.550 174.300 508.350 179.250 ;
        RECT 509.550 175.200 511.350 179.250 ;
        RECT 512.550 174.300 514.350 179.250 ;
        RECT 506.550 172.950 514.350 174.300 ;
        RECT 515.550 173.400 517.350 179.250 ;
        RECT 524.850 173.400 526.650 179.250 ;
        RECT 515.550 171.300 516.750 173.400 ;
        RECT 529.350 172.200 531.150 179.250 ;
        RECT 541.650 173.400 543.450 179.250 ;
        RECT 513.000 170.250 516.750 171.300 ;
        RECT 527.550 171.300 531.150 172.200 ;
        RECT 542.250 171.300 543.450 173.400 ;
        RECT 544.650 174.300 546.450 179.250 ;
        RECT 547.650 175.200 549.450 179.250 ;
        RECT 550.650 174.300 552.450 179.250 ;
        RECT 568.650 176.400 570.450 179.250 ;
        RECT 571.650 176.400 573.450 179.250 ;
        RECT 574.650 176.400 576.450 179.250 ;
        RECT 577.650 176.400 579.750 179.250 ;
        RECT 568.650 175.500 569.700 176.400 ;
        RECT 574.650 175.500 575.700 176.400 ;
        RECT 544.650 172.950 552.450 174.300 ;
        RECT 564.900 174.600 575.700 175.500 ;
        RECT 591.150 174.900 592.950 179.250 ;
        RECT 509.100 168.150 510.900 169.950 ;
        RECT 494.100 165.150 495.900 166.950 ;
        RECT 493.950 163.050 496.050 165.150 ;
        RECT 496.950 164.850 499.350 166.950 ;
        RECT 505.950 164.850 508.050 166.950 ;
        RECT 508.950 166.050 511.050 168.150 ;
        RECT 512.850 166.950 514.050 170.250 ;
        RECT 511.950 164.850 514.050 166.950 ;
        RECT 524.100 165.150 525.900 166.950 ;
        RECT 498.150 159.600 499.350 164.850 ;
        RECT 506.100 163.050 507.900 164.850 ;
        RECT 511.950 159.600 513.150 164.850 ;
        RECT 514.950 161.850 517.050 163.950 ;
        RECT 523.950 163.050 526.050 165.150 ;
        RECT 527.550 163.950 528.750 171.300 ;
        RECT 542.250 170.250 546.000 171.300 ;
        RECT 544.950 166.950 546.150 170.250 ;
        RECT 548.100 168.150 549.900 169.950 ;
        RECT 564.900 168.150 566.100 174.600 ;
        RECT 589.650 173.400 592.950 174.900 ;
        RECT 594.150 173.400 595.950 179.250 ;
        RECT 572.100 168.150 573.900 169.950 ;
        RECT 530.100 165.150 531.900 166.950 ;
        RECT 526.950 161.850 529.050 163.950 ;
        RECT 529.950 163.050 532.050 165.150 ;
        RECT 544.950 164.850 547.050 166.950 ;
        RECT 547.950 166.050 550.050 168.150 ;
        RECT 550.950 164.850 553.050 166.950 ;
        RECT 562.950 166.050 566.100 168.150 ;
        RECT 541.950 161.850 544.050 163.950 ;
        RECT 514.950 160.050 516.750 161.850 ;
        RECT 473.550 147.750 475.350 153.000 ;
        RECT 476.550 147.750 478.350 153.600 ;
        RECT 488.550 147.750 490.350 153.600 ;
        RECT 491.550 147.750 493.350 153.600 ;
        RECT 495.150 147.750 496.950 159.600 ;
        RECT 498.150 147.750 499.950 159.600 ;
        RECT 507.300 147.750 509.100 159.600 ;
        RECT 511.500 147.750 513.300 159.600 ;
        RECT 514.950 156.450 517.050 157.050 ;
        RECT 520.950 156.450 523.050 157.050 ;
        RECT 514.950 155.550 523.050 156.450 ;
        RECT 514.950 154.950 517.050 155.550 ;
        RECT 520.950 154.950 523.050 155.550 ;
        RECT 527.550 153.600 528.750 161.850 ;
        RECT 542.250 160.050 544.050 161.850 ;
        RECT 545.850 159.600 547.050 164.850 ;
        RECT 551.100 163.050 552.900 164.850 ;
        RECT 564.900 160.800 566.100 166.050 ;
        RECT 568.950 164.850 571.050 166.950 ;
        RECT 571.950 166.050 574.050 168.150 ;
        RECT 589.650 166.950 590.850 173.400 ;
        RECT 592.950 171.900 594.750 172.500 ;
        RECT 598.650 171.900 600.450 179.250 ;
        RECT 610.650 173.400 612.450 179.250 ;
        RECT 592.950 170.700 600.450 171.900 ;
        RECT 607.950 171.450 610.050 172.050 ;
        RECT 577.950 164.850 580.050 166.950 ;
        RECT 589.650 164.850 592.050 166.950 ;
        RECT 593.100 165.150 594.900 166.950 ;
        RECT 569.100 163.050 570.900 164.850 ;
        RECT 578.100 163.050 579.900 164.850 ;
        RECT 562.650 159.600 566.100 160.800 ;
        RECT 589.650 159.600 590.850 164.850 ;
        RECT 592.950 163.050 595.050 165.150 ;
        RECT 514.800 147.750 516.600 153.600 ;
        RECT 524.550 147.750 526.350 153.600 ;
        RECT 527.550 147.750 529.350 153.600 ;
        RECT 530.550 147.750 532.350 153.600 ;
        RECT 542.400 147.750 544.200 153.600 ;
        RECT 545.700 147.750 547.500 159.600 ;
        RECT 549.900 147.750 551.700 159.600 ;
        RECT 559.050 148.500 560.850 157.800 ;
        RECT 562.650 157.200 563.850 159.600 ;
        RECT 562.050 149.400 563.850 157.200 ;
        RECT 565.050 157.200 573.450 158.100 ;
        RECT 565.050 148.500 566.850 157.200 ;
        RECT 559.050 147.750 566.850 148.500 ;
        RECT 568.650 148.500 570.450 156.300 ;
        RECT 571.650 149.400 573.450 157.200 ;
        RECT 574.650 157.500 582.450 158.400 ;
        RECT 574.650 148.500 576.450 157.500 ;
        RECT 568.650 147.750 576.450 148.500 ;
        RECT 577.650 147.750 579.450 156.600 ;
        RECT 580.650 147.750 582.450 157.500 ;
        RECT 589.050 147.750 590.850 159.600 ;
        RECT 592.050 147.750 593.850 159.600 ;
        RECT 596.100 153.600 597.300 170.700 ;
        RECT 605.550 170.550 610.050 171.450 ;
        RECT 598.950 164.850 601.050 166.950 ;
        RECT 605.550 166.050 606.450 170.550 ;
        RECT 607.950 169.950 610.050 170.550 ;
        RECT 611.250 171.300 612.450 173.400 ;
        RECT 613.650 174.300 615.450 179.250 ;
        RECT 616.650 175.200 618.450 179.250 ;
        RECT 619.650 174.300 621.450 179.250 ;
        RECT 613.650 172.950 621.450 174.300 ;
        RECT 623.550 174.300 625.350 179.250 ;
        RECT 626.550 175.200 628.350 179.250 ;
        RECT 629.550 174.300 631.350 179.250 ;
        RECT 623.550 172.950 631.350 174.300 ;
        RECT 632.550 173.400 634.350 179.250 ;
        RECT 638.850 173.400 640.650 179.250 ;
        RECT 632.550 171.300 633.750 173.400 ;
        RECT 643.350 172.200 645.150 179.250 ;
        RECT 656.550 176.400 658.350 179.250 ;
        RECT 659.550 176.400 661.350 179.250 ;
        RECT 662.550 176.400 664.350 179.250 ;
        RECT 611.250 170.250 615.000 171.300 ;
        RECT 630.000 170.250 633.750 171.300 ;
        RECT 641.550 171.300 645.150 172.200 ;
        RECT 610.950 168.450 613.050 169.050 ;
        RECT 608.550 167.550 613.050 168.450 ;
        RECT 599.100 163.050 600.900 164.850 ;
        RECT 604.950 163.950 607.050 166.050 ;
        RECT 608.550 162.450 609.450 167.550 ;
        RECT 610.950 166.950 613.050 167.550 ;
        RECT 613.950 166.950 615.150 170.250 ;
        RECT 617.100 168.150 618.900 169.950 ;
        RECT 626.100 168.150 627.900 169.950 ;
        RECT 613.950 164.850 616.050 166.950 ;
        RECT 616.950 166.050 619.050 168.150 ;
        RECT 619.950 164.850 622.050 166.950 ;
        RECT 622.950 164.850 625.050 166.950 ;
        RECT 625.950 166.050 628.050 168.150 ;
        RECT 629.850 166.950 631.050 170.250 ;
        RECT 628.950 164.850 631.050 166.950 ;
        RECT 638.100 165.150 639.900 166.950 ;
        RECT 605.550 161.550 609.450 162.450 ;
        RECT 610.950 161.850 613.050 163.950 ;
        RECT 605.550 160.050 606.450 161.550 ;
        RECT 611.250 160.050 613.050 161.850 ;
        RECT 604.950 157.950 607.050 160.050 ;
        RECT 614.850 159.600 616.050 164.850 ;
        RECT 620.100 163.050 621.900 164.850 ;
        RECT 623.100 163.050 624.900 164.850 ;
        RECT 628.950 159.600 630.150 164.850 ;
        RECT 631.950 161.850 634.050 163.950 ;
        RECT 637.950 163.050 640.050 165.150 ;
        RECT 641.550 163.950 642.750 171.300 ;
        RECT 660.000 169.950 661.050 176.400 ;
        RECT 674.700 170.400 676.500 179.250 ;
        RECT 680.100 171.000 681.900 179.250 ;
        RECT 658.950 167.850 661.050 169.950 ;
        RECT 680.100 169.350 684.600 171.000 ;
        RECT 692.700 170.400 694.500 179.250 ;
        RECT 698.100 171.000 699.900 179.250 ;
        RECT 698.100 169.350 702.600 171.000 ;
        RECT 710.700 170.400 712.500 179.250 ;
        RECT 716.100 171.000 717.900 179.250 ;
        RECT 731.550 174.300 733.350 179.250 ;
        RECT 734.550 175.200 736.350 179.250 ;
        RECT 737.550 174.300 739.350 179.250 ;
        RECT 731.550 172.950 739.350 174.300 ;
        RECT 740.550 173.400 742.350 179.250 ;
        RECT 751.650 176.400 753.450 179.250 ;
        RECT 754.650 176.400 756.450 179.250 ;
        RECT 757.650 176.400 759.450 179.250 ;
        RECT 766.650 176.400 768.450 179.250 ;
        RECT 769.650 176.400 771.450 179.250 ;
        RECT 772.650 176.400 774.450 179.250 ;
        RECT 777.750 176.400 779.550 179.250 ;
        RECT 780.750 176.400 782.550 179.250 ;
        RECT 740.550 171.300 741.750 173.400 ;
        RECT 716.100 169.350 720.600 171.000 ;
        RECT 738.000 170.250 741.750 171.300 ;
        RECT 644.100 165.150 645.900 166.950 ;
        RECT 640.950 161.850 643.050 163.950 ;
        RECT 643.950 163.050 646.050 165.150 ;
        RECT 655.950 164.850 658.050 166.950 ;
        RECT 656.100 163.050 657.900 164.850 ;
        RECT 631.950 160.050 633.750 161.850 ;
        RECT 595.650 147.750 597.450 153.600 ;
        RECT 598.650 147.750 600.450 153.600 ;
        RECT 611.400 147.750 613.200 153.600 ;
        RECT 614.700 147.750 616.500 159.600 ;
        RECT 618.900 147.750 620.700 159.600 ;
        RECT 624.300 147.750 626.100 159.600 ;
        RECT 628.500 147.750 630.300 159.600 ;
        RECT 641.550 153.600 642.750 161.850 ;
        RECT 660.000 160.650 661.050 167.850 ;
        RECT 670.950 166.950 673.050 169.050 ;
        RECT 661.950 164.850 664.050 166.950 ;
        RECT 662.100 163.050 663.900 164.850 ;
        RECT 660.000 159.600 662.550 160.650 ;
        RECT 631.800 147.750 633.600 153.600 ;
        RECT 638.550 147.750 640.350 153.600 ;
        RECT 641.550 147.750 643.350 153.600 ;
        RECT 644.550 147.750 646.350 153.600 ;
        RECT 656.550 147.750 658.350 159.600 ;
        RECT 660.750 147.750 662.550 159.600 ;
        RECT 671.550 156.450 672.450 166.950 ;
        RECT 683.400 165.150 684.600 169.350 ;
        RECT 701.400 165.150 702.600 169.350 ;
        RECT 719.400 165.150 720.600 169.350 ;
        RECT 734.100 168.150 735.900 169.950 ;
        RECT 673.950 161.850 676.050 163.950 ;
        RECT 679.950 161.850 682.050 163.950 ;
        RECT 682.950 163.050 685.050 165.150 ;
        RECT 674.100 160.050 675.900 161.850 ;
        RECT 676.950 158.850 679.050 160.950 ;
        RECT 680.250 160.050 682.050 161.850 ;
        RECT 677.100 157.050 678.900 158.850 ;
        RECT 673.950 156.450 676.050 157.050 ;
        RECT 671.550 155.550 676.050 156.450 ;
        RECT 673.950 154.950 676.050 155.550 ;
        RECT 683.700 154.800 684.750 163.050 ;
        RECT 691.950 161.850 694.050 163.950 ;
        RECT 697.950 161.850 700.050 163.950 ;
        RECT 700.950 163.050 703.050 165.150 ;
        RECT 692.100 160.050 693.900 161.850 ;
        RECT 694.950 158.850 697.050 160.950 ;
        RECT 698.250 160.050 700.050 161.850 ;
        RECT 695.100 157.050 696.900 158.850 ;
        RECT 701.700 154.800 702.750 163.050 ;
        RECT 709.950 161.850 712.050 163.950 ;
        RECT 715.950 161.850 718.050 163.950 ;
        RECT 718.950 163.050 721.050 165.150 ;
        RECT 730.950 164.850 733.050 166.950 ;
        RECT 733.950 166.050 736.050 168.150 ;
        RECT 737.850 166.950 739.050 170.250 ;
        RECT 754.950 169.950 756.000 176.400 ;
        RECT 769.950 169.950 771.000 176.400 ;
        RECT 754.950 167.850 757.050 169.950 ;
        RECT 769.950 167.850 772.050 169.950 ;
        RECT 781.050 168.150 782.550 176.400 ;
        RECT 736.950 164.850 739.050 166.950 ;
        RECT 751.950 164.850 754.050 166.950 ;
        RECT 731.100 163.050 732.900 164.850 ;
        RECT 710.100 160.050 711.900 161.850 ;
        RECT 712.950 158.850 715.050 160.950 ;
        RECT 716.250 160.050 718.050 161.850 ;
        RECT 713.100 157.050 714.900 158.850 ;
        RECT 719.700 154.800 720.750 163.050 ;
        RECT 736.950 159.600 738.150 164.850 ;
        RECT 739.950 161.850 742.050 163.950 ;
        RECT 752.100 163.050 753.900 164.850 ;
        RECT 739.950 160.050 741.750 161.850 ;
        RECT 754.950 160.650 756.000 167.850 ;
        RECT 757.950 164.850 760.050 166.950 ;
        RECT 766.950 164.850 769.050 166.950 ;
        RECT 758.100 163.050 759.900 164.850 ;
        RECT 767.100 163.050 768.900 164.850 ;
        RECT 769.950 160.650 771.000 167.850 ;
        RECT 772.950 164.850 775.050 166.950 ;
        RECT 778.950 166.050 782.550 168.150 ;
        RECT 773.100 163.050 774.900 164.850 ;
        RECT 753.450 159.600 756.000 160.650 ;
        RECT 768.450 159.600 771.000 160.650 ;
        RECT 677.700 153.900 684.750 154.800 ;
        RECT 677.700 153.600 679.350 153.900 ;
        RECT 674.550 147.750 676.350 153.600 ;
        RECT 677.550 147.750 679.350 153.600 ;
        RECT 683.550 153.600 684.750 153.900 ;
        RECT 695.700 153.900 702.750 154.800 ;
        RECT 695.700 153.600 697.350 153.900 ;
        RECT 680.550 147.750 682.350 153.000 ;
        RECT 683.550 147.750 685.350 153.600 ;
        RECT 692.550 147.750 694.350 153.600 ;
        RECT 695.550 147.750 697.350 153.600 ;
        RECT 701.550 153.600 702.750 153.900 ;
        RECT 713.700 153.900 720.750 154.800 ;
        RECT 713.700 153.600 715.350 153.900 ;
        RECT 698.550 147.750 700.350 153.000 ;
        RECT 701.550 147.750 703.350 153.600 ;
        RECT 710.550 147.750 712.350 153.600 ;
        RECT 713.550 147.750 715.350 153.600 ;
        RECT 719.550 153.600 720.750 153.900 ;
        RECT 716.550 147.750 718.350 153.000 ;
        RECT 719.550 147.750 721.350 153.600 ;
        RECT 732.300 147.750 734.100 159.600 ;
        RECT 736.500 147.750 738.300 159.600 ;
        RECT 739.800 147.750 741.600 153.600 ;
        RECT 753.450 147.750 755.250 159.600 ;
        RECT 757.650 147.750 759.450 159.600 ;
        RECT 768.450 147.750 770.250 159.600 ;
        RECT 772.650 147.750 774.450 159.600 ;
        RECT 781.050 153.600 782.550 166.050 ;
        RECT 784.650 173.400 786.450 179.250 ;
        RECT 790.050 173.400 791.850 179.250 ;
        RECT 795.600 174.600 797.400 179.250 ;
        RECT 800.250 175.500 802.050 179.250 ;
        RECT 803.250 175.500 805.050 179.250 ;
        RECT 806.250 175.500 808.050 179.250 ;
        RECT 793.200 173.400 797.400 174.600 ;
        RECT 799.950 173.400 802.050 175.500 ;
        RECT 802.950 173.400 805.050 175.500 ;
        RECT 805.950 173.400 808.050 175.500 ;
        RECT 810.000 175.500 811.800 179.250 ;
        RECT 813.000 176.400 814.800 179.250 ;
        RECT 816.000 175.500 817.800 179.250 ;
        RECT 820.500 176.400 822.300 179.250 ;
        RECT 823.500 176.400 825.300 179.250 ;
        RECT 826.500 176.400 828.300 179.250 ;
        RECT 829.500 176.400 831.300 179.250 ;
        RECT 810.000 173.700 812.850 175.500 ;
        RECT 810.750 173.400 812.850 173.700 ;
        RECT 814.950 173.700 817.800 175.500 ;
        RECT 818.700 174.750 820.500 175.200 ;
        RECT 823.950 175.050 825.300 176.400 ;
        RECT 826.950 175.050 828.300 176.400 ;
        RECT 829.950 175.050 831.300 176.400 ;
        RECT 814.950 173.400 817.050 173.700 ;
        RECT 818.700 173.400 822.750 174.750 ;
        RECT 784.650 158.550 785.850 173.400 ;
        RECT 793.200 169.800 794.700 173.400 ;
        RECT 799.350 170.700 806.100 172.500 ;
        RECT 807.000 170.700 813.900 172.500 ;
        RECT 821.850 172.050 822.750 173.400 ;
        RECT 823.950 172.950 826.050 175.050 ;
        RECT 826.950 172.950 829.050 175.050 ;
        RECT 829.950 172.950 832.050 175.050 ;
        RECT 821.850 171.900 826.950 172.050 ;
        RECT 821.850 171.150 829.500 171.900 ;
        RECT 825.150 170.700 829.500 171.150 ;
        RECT 807.000 169.800 808.050 170.700 ;
        RECT 825.150 170.250 826.950 170.700 ;
        RECT 786.900 168.000 794.700 169.800 ;
        RECT 798.150 168.750 808.050 169.800 ;
        RECT 798.150 166.950 799.200 168.750 ;
        RECT 808.950 168.450 816.600 169.800 ;
        RECT 808.950 167.700 809.850 168.450 ;
        RECT 790.950 165.900 799.200 166.950 ;
        RECT 800.250 166.650 809.850 167.700 ;
        RECT 790.950 161.850 793.050 165.900 ;
        RECT 800.250 165.000 801.150 166.650 ;
        RECT 810.750 165.750 814.650 167.550 ;
        RECT 815.550 166.950 816.600 168.450 ;
        RECT 817.950 169.650 820.050 169.950 ;
        RECT 817.950 167.850 821.850 169.650 ;
        RECT 828.450 167.250 829.500 170.700 ;
        RECT 831.000 169.800 832.050 172.950 ;
        RECT 833.700 173.400 835.500 179.250 ;
        RECT 839.100 173.400 840.900 179.250 ;
        RECT 844.500 173.400 846.300 179.250 ;
        RECT 850.650 173.400 852.450 179.250 ;
        RECT 853.650 176.400 855.450 179.250 ;
        RECT 856.650 176.400 858.450 179.250 ;
        RECT 859.650 176.400 861.450 179.250 ;
        RECT 833.700 172.500 835.200 173.400 ;
        RECT 833.700 171.300 842.100 172.500 ;
        RECT 840.300 170.700 842.100 171.300 ;
        RECT 845.100 169.800 846.300 173.400 ;
        RECT 831.000 168.900 846.300 169.800 ;
        RECT 815.550 166.050 827.550 166.950 ;
        RECT 794.100 163.200 801.150 165.000 ;
        RECT 802.500 163.950 804.300 165.750 ;
        RECT 810.750 165.450 812.850 165.750 ;
        RECT 814.950 164.550 817.050 164.850 ;
        RECT 823.800 164.550 825.600 165.150 ;
        RECT 814.950 163.950 825.600 164.550 ;
        RECT 802.500 163.350 825.600 163.950 ;
        RECT 826.500 164.550 827.550 166.050 ;
        RECT 828.450 165.450 830.250 167.250 ;
        RECT 832.050 166.950 843.900 168.000 ;
        RECT 832.050 164.550 833.250 166.950 ;
        RECT 842.100 165.150 843.900 166.950 ;
        RECT 826.500 163.650 833.250 164.550 ;
        RECT 835.950 163.650 838.050 163.950 ;
        RECT 802.500 162.750 817.050 163.350 ;
        RECT 834.150 162.450 838.050 163.650 ;
        RECT 841.950 163.050 844.050 165.150 ;
        RECT 824.100 161.850 838.050 162.450 ;
        RECT 798.000 161.550 837.750 161.850 ;
        RECT 786.750 160.650 788.550 161.250 ;
        RECT 798.000 160.650 826.050 161.550 ;
        RECT 786.750 159.450 799.050 160.650 ;
        RECT 826.950 160.050 829.050 160.350 ;
        RECT 836.700 160.050 838.500 160.650 ;
        RECT 799.950 158.550 802.050 159.750 ;
        RECT 784.650 157.650 802.050 158.550 ;
        RECT 805.950 158.400 826.050 159.750 ;
        RECT 805.950 157.650 808.050 158.400 ;
        RECT 787.500 153.600 788.700 157.650 ;
        RECT 789.600 155.700 791.400 156.300 ;
        RECT 796.350 156.150 798.150 156.300 ;
        RECT 789.600 154.500 795.300 155.700 ;
        RECT 796.350 154.950 805.050 156.150 ;
        RECT 796.350 154.500 798.150 154.950 ;
        RECT 777.750 147.750 779.550 153.600 ;
        RECT 780.750 147.750 782.550 153.600 ;
        RECT 784.500 147.750 786.300 153.600 ;
        RECT 787.500 147.750 789.300 153.600 ;
        RECT 790.500 147.750 792.300 153.600 ;
        RECT 793.500 147.750 795.300 154.500 ;
        RECT 802.950 154.050 805.050 154.950 ;
        RECT 796.500 147.750 798.300 153.600 ;
        RECT 799.800 151.800 801.900 153.900 ;
        RECT 800.400 150.600 801.900 151.800 ;
        RECT 800.250 147.750 802.050 150.600 ;
        RECT 803.250 147.750 805.050 154.050 ;
        RECT 806.550 150.600 807.900 157.650 ;
        RECT 824.100 157.350 826.050 158.400 ;
        RECT 826.950 158.850 838.500 160.050 ;
        RECT 826.950 158.250 829.050 158.850 ;
        RECT 840.000 157.350 841.800 158.100 ;
        RECT 809.100 154.800 813.000 156.600 ;
        RECT 810.000 154.500 813.000 154.800 ;
        RECT 814.950 156.150 817.050 156.600 ;
        RECT 824.100 156.300 841.800 157.350 ;
        RECT 814.950 154.500 817.350 156.150 ;
        RECT 806.250 147.750 808.050 150.600 ;
        RECT 810.000 147.750 811.800 154.500 ;
        RECT 816.000 153.600 817.350 154.500 ;
        RECT 823.950 153.600 826.050 154.050 ;
        RECT 813.000 147.750 814.800 153.600 ;
        RECT 816.000 147.750 817.800 153.600 ;
        RECT 819.750 147.750 821.550 153.600 ;
        RECT 823.500 151.950 826.050 153.600 ;
        RECT 826.950 151.950 829.050 154.050 ;
        RECT 829.950 151.950 832.050 154.050 ;
        RECT 823.500 150.600 824.700 151.950 ;
        RECT 826.950 150.600 827.850 151.950 ;
        RECT 829.950 150.600 831.150 151.950 ;
        RECT 822.750 147.750 824.700 150.600 ;
        RECT 825.750 147.750 827.850 150.600 ;
        RECT 828.750 147.750 831.150 150.600 ;
        RECT 832.500 147.750 834.300 151.050 ;
        RECT 835.500 147.750 837.300 156.300 ;
        RECT 845.100 155.400 846.300 168.900 ;
        RECT 850.950 168.150 852.000 173.400 ;
        RECT 856.650 172.200 857.550 176.400 ;
        RECT 854.250 171.300 857.550 172.200 ;
        RECT 854.250 170.400 856.050 171.300 ;
        RECT 850.950 166.050 853.050 168.150 ;
        RECT 851.550 159.450 852.900 166.050 ;
        RECT 854.400 162.150 855.300 170.400 ;
        RECT 859.950 167.850 862.050 169.950 ;
        RECT 856.950 164.850 859.050 166.950 ;
        RECT 860.100 166.050 861.900 167.850 ;
        RECT 857.100 163.050 858.900 164.850 ;
        RECT 854.250 162.000 856.050 162.150 ;
        RECT 854.250 160.800 861.450 162.000 ;
        RECT 854.250 160.350 856.050 160.800 ;
        RECT 860.250 159.600 861.450 160.800 ;
        RECT 851.550 158.100 853.950 159.450 ;
        RECT 842.250 154.500 846.300 155.400 ;
        RECT 842.250 153.600 843.300 154.500 ;
        RECT 838.500 147.750 840.300 153.600 ;
        RECT 841.500 147.750 843.300 153.600 ;
        RECT 844.500 147.750 846.300 153.600 ;
        RECT 852.150 147.750 853.950 158.100 ;
        RECT 855.150 147.750 856.950 159.450 ;
        RECT 859.650 147.750 861.450 159.600 ;
        RECT 2.700 137.400 4.500 143.250 ;
        RECT 5.700 137.400 7.500 143.250 ;
        RECT 8.700 137.400 10.500 143.250 ;
        RECT 5.700 136.500 6.750 137.400 ;
        RECT 2.700 135.600 6.750 136.500 ;
        RECT 2.700 122.100 3.900 135.600 ;
        RECT 11.700 134.700 13.500 143.250 ;
        RECT 14.700 139.950 16.500 143.250 ;
        RECT 17.850 140.400 20.250 143.250 ;
        RECT 21.150 140.400 23.250 143.250 ;
        RECT 24.300 140.400 26.250 143.250 ;
        RECT 17.850 139.050 19.050 140.400 ;
        RECT 21.150 139.050 22.050 140.400 ;
        RECT 24.300 139.050 25.500 140.400 ;
        RECT 16.950 136.950 19.050 139.050 ;
        RECT 19.950 136.950 22.050 139.050 ;
        RECT 22.950 137.400 25.500 139.050 ;
        RECT 27.450 137.400 29.250 143.250 ;
        RECT 31.200 137.400 33.000 143.250 ;
        RECT 34.200 137.400 36.000 143.250 ;
        RECT 22.950 136.950 25.050 137.400 ;
        RECT 31.650 136.500 33.000 137.400 ;
        RECT 37.200 136.500 39.000 143.250 ;
        RECT 40.950 140.400 42.750 143.250 ;
        RECT 31.650 134.850 34.050 136.500 ;
        RECT 7.200 133.650 24.900 134.700 ;
        RECT 31.950 134.400 34.050 134.850 ;
        RECT 36.000 136.200 39.000 136.500 ;
        RECT 36.000 134.400 39.900 136.200 ;
        RECT 7.200 132.900 9.000 133.650 ;
        RECT 19.950 132.150 22.050 132.750 ;
        RECT 10.500 130.950 22.050 132.150 ;
        RECT 22.950 132.600 24.900 133.650 ;
        RECT 41.100 133.350 42.450 140.400 ;
        RECT 43.950 136.950 45.750 143.250 ;
        RECT 46.950 140.400 48.750 143.250 ;
        RECT 47.100 139.200 48.600 140.400 ;
        RECT 47.100 137.100 49.200 139.200 ;
        RECT 50.700 137.400 52.500 143.250 ;
        RECT 43.950 136.050 46.050 136.950 ;
        RECT 53.700 136.500 55.500 143.250 ;
        RECT 56.700 137.400 58.500 143.250 ;
        RECT 59.700 137.400 61.500 143.250 ;
        RECT 62.700 137.400 64.500 143.250 ;
        RECT 66.450 137.400 68.250 143.250 ;
        RECT 69.450 137.400 71.250 143.250 ;
        RECT 82.650 137.400 84.450 143.250 ;
        RECT 85.650 137.400 87.450 143.250 ;
        RECT 88.650 137.400 90.450 143.250 ;
        RECT 92.550 137.400 94.350 143.250 ;
        RECT 95.550 137.400 97.350 143.250 ;
        RECT 50.850 136.050 52.650 136.500 ;
        RECT 43.950 134.850 52.650 136.050 ;
        RECT 53.700 135.300 59.400 136.500 ;
        RECT 50.850 134.700 52.650 134.850 ;
        RECT 57.600 134.700 59.400 135.300 ;
        RECT 60.300 133.350 61.500 137.400 ;
        RECT 40.950 132.600 43.050 133.350 ;
        RECT 22.950 131.250 43.050 132.600 ;
        RECT 46.950 132.450 64.350 133.350 ;
        RECT 46.950 131.250 49.050 132.450 ;
        RECT 10.500 130.350 12.300 130.950 ;
        RECT 19.950 130.650 22.050 130.950 ;
        RECT 49.950 130.350 62.250 131.550 ;
        RECT 22.950 129.450 51.000 130.350 ;
        RECT 60.450 129.750 62.250 130.350 ;
        RECT 11.250 129.150 51.000 129.450 ;
        RECT 10.950 128.550 24.900 129.150 ;
        RECT 4.950 125.850 7.050 127.950 ;
        RECT 10.950 127.350 14.850 128.550 ;
        RECT 31.950 127.650 46.500 128.250 ;
        RECT 10.950 127.050 13.050 127.350 ;
        RECT 15.750 126.450 22.500 127.350 ;
        RECT 5.100 124.050 6.900 125.850 ;
        RECT 15.750 124.050 16.950 126.450 ;
        RECT 5.100 123.000 16.950 124.050 ;
        RECT 18.750 123.750 20.550 125.550 ;
        RECT 21.450 124.950 22.500 126.450 ;
        RECT 23.400 127.050 46.500 127.650 ;
        RECT 23.400 126.450 34.050 127.050 ;
        RECT 23.400 125.850 25.200 126.450 ;
        RECT 31.950 126.150 34.050 126.450 ;
        RECT 36.150 125.250 38.250 125.550 ;
        RECT 44.700 125.250 46.500 127.050 ;
        RECT 47.850 126.000 54.900 127.800 ;
        RECT 21.450 124.050 33.450 124.950 ;
        RECT 2.700 121.200 18.000 122.100 ;
        RECT 2.700 117.600 3.900 121.200 ;
        RECT 6.900 119.700 8.700 120.300 ;
        RECT 6.900 118.500 15.300 119.700 ;
        RECT 13.800 117.600 15.300 118.500 ;
        RECT 2.700 111.750 4.500 117.600 ;
        RECT 8.100 111.750 9.900 117.600 ;
        RECT 13.500 111.750 15.300 117.600 ;
        RECT 16.950 118.050 18.000 121.200 ;
        RECT 19.500 120.300 20.550 123.750 ;
        RECT 27.150 121.350 31.050 123.150 ;
        RECT 28.950 121.050 31.050 121.350 ;
        RECT 32.400 122.550 33.450 124.050 ;
        RECT 34.350 123.450 38.250 125.250 ;
        RECT 47.850 124.350 48.750 126.000 ;
        RECT 55.950 125.100 58.050 129.150 ;
        RECT 39.150 123.300 48.750 124.350 ;
        RECT 49.800 124.050 58.050 125.100 ;
        RECT 39.150 122.550 40.050 123.300 ;
        RECT 32.400 121.200 40.050 122.550 ;
        RECT 49.800 122.250 50.850 124.050 ;
        RECT 40.950 121.200 50.850 122.250 ;
        RECT 54.300 121.200 62.100 123.000 ;
        RECT 22.050 120.300 23.850 120.750 ;
        RECT 40.950 120.300 42.000 121.200 ;
        RECT 19.500 119.850 23.850 120.300 ;
        RECT 19.500 119.100 27.150 119.850 ;
        RECT 22.050 118.950 27.150 119.100 ;
        RECT 16.950 115.950 19.050 118.050 ;
        RECT 19.950 115.950 22.050 118.050 ;
        RECT 22.950 115.950 25.050 118.050 ;
        RECT 26.250 117.600 27.150 118.950 ;
        RECT 35.100 118.500 42.000 120.300 ;
        RECT 42.900 118.500 49.650 120.300 ;
        RECT 54.300 117.600 55.800 121.200 ;
        RECT 63.150 117.600 64.350 132.450 ;
        RECT 26.250 116.250 30.300 117.600 ;
        RECT 31.950 117.300 34.050 117.600 ;
        RECT 17.700 114.600 19.050 115.950 ;
        RECT 20.700 114.600 22.050 115.950 ;
        RECT 23.700 114.600 25.050 115.950 ;
        RECT 28.500 115.800 30.300 116.250 ;
        RECT 31.200 115.500 34.050 117.300 ;
        RECT 36.150 117.300 38.250 117.600 ;
        RECT 36.150 115.500 39.000 117.300 ;
        RECT 17.700 111.750 19.500 114.600 ;
        RECT 20.700 111.750 22.500 114.600 ;
        RECT 23.700 111.750 25.500 114.600 ;
        RECT 26.700 111.750 28.500 114.600 ;
        RECT 31.200 111.750 33.000 115.500 ;
        RECT 34.200 111.750 36.000 114.600 ;
        RECT 37.200 111.750 39.000 115.500 ;
        RECT 40.950 115.500 43.050 117.600 ;
        RECT 43.950 115.500 46.050 117.600 ;
        RECT 46.950 115.500 49.050 117.600 ;
        RECT 51.600 116.400 55.800 117.600 ;
        RECT 40.950 111.750 42.750 115.500 ;
        RECT 43.950 111.750 45.750 115.500 ;
        RECT 46.950 111.750 48.750 115.500 ;
        RECT 51.600 111.750 53.400 116.400 ;
        RECT 57.150 111.750 58.950 117.600 ;
        RECT 62.550 111.750 64.350 117.600 ;
        RECT 66.450 124.950 67.950 137.400 ;
        RECT 86.250 129.150 87.450 137.400 ;
        RECT 82.950 125.850 85.050 127.950 ;
        RECT 85.950 127.050 88.050 129.150 ;
        RECT 66.450 122.850 70.050 124.950 ;
        RECT 83.100 124.050 84.900 125.850 ;
        RECT 66.450 114.600 67.950 122.850 ;
        RECT 86.250 119.700 87.450 127.050 ;
        RECT 88.950 125.850 91.050 127.950 ;
        RECT 89.100 124.050 90.900 125.850 ;
        RECT 95.400 124.950 96.600 137.400 ;
        RECT 101.550 131.400 103.350 143.250 ;
        RECT 105.750 131.400 107.550 143.250 ;
        RECT 117.300 131.400 119.100 143.250 ;
        RECT 121.500 131.400 123.300 143.250 ;
        RECT 124.800 137.400 126.600 143.250 ;
        RECT 135.300 131.400 137.100 143.250 ;
        RECT 139.500 131.400 141.300 143.250 ;
        RECT 142.800 137.400 144.600 143.250 ;
        RECT 157.650 137.400 159.450 143.250 ;
        RECT 160.650 138.000 162.450 143.250 ;
        RECT 158.250 137.100 159.450 137.400 ;
        RECT 163.650 137.400 165.450 143.250 ;
        RECT 166.650 137.400 168.450 143.250 ;
        RECT 163.650 137.100 165.300 137.400 ;
        RECT 158.250 136.200 165.300 137.100 ;
        RECT 105.000 130.350 107.550 131.400 ;
        RECT 101.100 126.150 102.900 127.950 ;
        RECT 92.100 123.150 93.900 124.950 ;
        RECT 91.950 121.050 94.050 123.150 ;
        RECT 94.950 122.850 97.050 124.950 ;
        RECT 100.950 124.050 103.050 126.150 ;
        RECT 105.000 123.150 106.050 130.350 ;
        RECT 107.100 126.150 108.900 127.950 ;
        RECT 116.100 126.150 117.900 127.950 ;
        RECT 121.950 126.150 123.150 131.400 ;
        RECT 124.950 129.150 126.750 130.950 ;
        RECT 124.950 127.050 127.050 129.150 ;
        RECT 134.100 126.150 135.900 127.950 ;
        RECT 139.950 126.150 141.150 131.400 ;
        RECT 142.950 129.150 144.750 130.950 ;
        RECT 142.950 127.050 145.050 129.150 ;
        RECT 158.250 127.950 159.300 136.200 ;
        RECT 164.100 132.150 165.900 133.950 ;
        RECT 160.950 129.150 162.750 130.950 ;
        RECT 163.950 130.050 166.050 132.150 ;
        RECT 172.650 131.400 174.450 143.250 ;
        RECT 175.650 132.300 177.450 143.250 ;
        RECT 178.650 133.200 180.450 143.250 ;
        RECT 181.650 132.300 183.450 143.250 ;
        RECT 193.650 137.400 195.450 143.250 ;
        RECT 196.650 138.000 198.450 143.250 ;
        RECT 175.650 131.400 183.450 132.300 ;
        RECT 194.250 137.100 195.450 137.400 ;
        RECT 199.650 137.400 201.450 143.250 ;
        RECT 202.650 137.400 204.450 143.250 ;
        RECT 211.650 137.400 213.450 143.250 ;
        RECT 214.650 137.400 216.450 143.250 ;
        RECT 217.650 137.400 219.450 143.250 ;
        RECT 221.550 137.400 223.350 143.250 ;
        RECT 224.550 137.400 226.350 143.250 ;
        RECT 227.550 138.000 229.350 143.250 ;
        RECT 199.650 137.100 201.300 137.400 ;
        RECT 194.250 136.200 201.300 137.100 ;
        RECT 167.100 129.150 168.900 130.950 ;
        RECT 106.950 124.050 109.050 126.150 ;
        RECT 115.950 124.050 118.050 126.150 ;
        RECT 83.850 118.800 87.450 119.700 ;
        RECT 66.450 111.750 68.250 114.600 ;
        RECT 69.450 111.750 71.250 114.600 ;
        RECT 83.850 111.750 85.650 118.800 ;
        RECT 88.350 111.750 90.150 117.600 ;
        RECT 95.400 114.600 96.600 122.850 ;
        RECT 103.950 121.050 106.050 123.150 ;
        RECT 118.950 122.850 121.050 124.950 ;
        RECT 121.950 124.050 124.050 126.150 ;
        RECT 133.950 124.050 136.050 126.150 ;
        RECT 119.100 121.050 120.900 122.850 ;
        RECT 105.000 114.600 106.050 121.050 ;
        RECT 122.850 120.750 124.050 124.050 ;
        RECT 136.950 122.850 139.050 124.950 ;
        RECT 139.950 124.050 142.050 126.150 ;
        RECT 157.950 125.850 160.050 127.950 ;
        RECT 160.950 127.050 163.050 129.150 ;
        RECT 166.950 127.050 169.050 129.150 ;
        RECT 173.100 126.150 174.300 131.400 ;
        RECT 194.250 127.950 195.300 136.200 ;
        RECT 200.100 132.150 201.900 133.950 ;
        RECT 196.950 129.150 198.750 130.950 ;
        RECT 199.950 130.050 202.050 132.150 ;
        RECT 203.100 129.150 204.900 130.950 ;
        RECT 215.250 129.150 216.450 137.400 ;
        RECT 224.700 137.100 226.350 137.400 ;
        RECT 230.550 137.400 232.350 143.250 ;
        RECT 241.650 137.400 243.450 143.250 ;
        RECT 244.650 137.400 246.450 143.250 ;
        RECT 247.650 137.400 249.450 143.250 ;
        RECT 254.550 137.400 256.350 143.250 ;
        RECT 257.550 137.400 259.350 143.250 ;
        RECT 260.550 137.400 262.350 143.250 ;
        RECT 271.650 137.400 273.450 143.250 ;
        RECT 274.650 137.400 276.450 143.250 ;
        RECT 277.650 137.400 279.450 143.250 ;
        RECT 283.650 137.400 285.450 143.250 ;
        RECT 286.650 137.400 288.450 143.250 ;
        RECT 289.650 137.400 291.450 143.250 ;
        RECT 299.550 137.400 301.350 143.250 ;
        RECT 302.550 137.400 304.350 143.250 ;
        RECT 230.550 137.100 231.750 137.400 ;
        RECT 224.700 136.200 231.750 137.100 ;
        RECT 224.100 132.150 225.900 133.950 ;
        RECT 221.100 129.150 222.900 130.950 ;
        RECT 223.950 130.050 226.050 132.150 ;
        RECT 227.250 129.150 229.050 130.950 ;
        RECT 137.100 121.050 138.900 122.850 ;
        RECT 140.850 120.750 142.050 124.050 ;
        RECT 158.400 121.650 159.600 125.850 ;
        RECT 172.950 124.050 175.050 126.150 ;
        RECT 193.950 125.850 196.050 127.950 ;
        RECT 196.950 127.050 199.050 129.150 ;
        RECT 202.950 127.050 205.050 129.150 ;
        RECT 211.950 125.850 214.050 127.950 ;
        RECT 214.950 127.050 217.050 129.150 ;
        RECT 123.000 119.700 126.750 120.750 ;
        RECT 141.000 119.700 144.750 120.750 ;
        RECT 158.400 120.000 162.900 121.650 ;
        RECT 116.550 116.700 124.350 118.050 ;
        RECT 92.550 111.750 94.350 114.600 ;
        RECT 95.550 111.750 97.350 114.600 ;
        RECT 101.550 111.750 103.350 114.600 ;
        RECT 104.550 111.750 106.350 114.600 ;
        RECT 107.550 111.750 109.350 114.600 ;
        RECT 116.550 111.750 118.350 116.700 ;
        RECT 119.550 111.750 121.350 115.800 ;
        RECT 122.550 111.750 124.350 116.700 ;
        RECT 125.550 117.600 126.750 119.700 ;
        RECT 125.550 111.750 127.350 117.600 ;
        RECT 134.550 116.700 142.350 118.050 ;
        RECT 134.550 111.750 136.350 116.700 ;
        RECT 137.550 111.750 139.350 115.800 ;
        RECT 140.550 111.750 142.350 116.700 ;
        RECT 143.550 117.600 144.750 119.700 ;
        RECT 143.550 111.750 145.350 117.600 ;
        RECT 161.100 111.750 162.900 120.000 ;
        RECT 166.500 111.750 168.300 120.600 ;
        RECT 173.100 117.600 174.300 124.050 ;
        RECT 175.950 122.850 178.050 124.950 ;
        RECT 179.100 123.150 180.900 124.950 ;
        RECT 176.100 121.050 177.900 122.850 ;
        RECT 178.950 121.050 181.050 123.150 ;
        RECT 181.950 122.850 184.050 124.950 ;
        RECT 182.100 121.050 183.900 122.850 ;
        RECT 194.400 121.650 195.600 125.850 ;
        RECT 212.100 124.050 213.900 125.850 ;
        RECT 194.400 120.000 198.900 121.650 ;
        RECT 173.100 115.950 178.800 117.600 ;
        RECT 173.700 111.750 175.500 114.600 ;
        RECT 177.000 111.750 178.800 115.950 ;
        RECT 181.200 111.750 183.000 117.600 ;
        RECT 197.100 111.750 198.900 120.000 ;
        RECT 202.500 111.750 204.300 120.600 ;
        RECT 215.250 119.700 216.450 127.050 ;
        RECT 217.950 125.850 220.050 127.950 ;
        RECT 220.950 127.050 223.050 129.150 ;
        RECT 226.950 127.050 229.050 129.150 ;
        RECT 230.700 127.950 231.750 136.200 ;
        RECT 245.250 129.150 246.450 137.400 ;
        RECT 257.550 129.150 258.750 137.400 ;
        RECT 275.250 129.150 276.450 137.400 ;
        RECT 287.250 129.150 288.450 137.400 ;
        RECT 229.950 125.850 232.050 127.950 ;
        RECT 241.950 125.850 244.050 127.950 ;
        RECT 244.950 127.050 247.050 129.150 ;
        RECT 218.100 124.050 219.900 125.850 ;
        RECT 230.400 121.650 231.600 125.850 ;
        RECT 242.100 124.050 243.900 125.850 ;
        RECT 212.850 118.800 216.450 119.700 ;
        RECT 212.850 111.750 214.650 118.800 ;
        RECT 217.350 111.750 219.150 117.600 ;
        RECT 221.700 111.750 223.500 120.600 ;
        RECT 227.100 120.000 231.600 121.650 ;
        RECT 227.100 111.750 228.900 120.000 ;
        RECT 245.250 119.700 246.450 127.050 ;
        RECT 247.950 125.850 250.050 127.950 ;
        RECT 253.950 125.850 256.050 127.950 ;
        RECT 256.950 127.050 259.050 129.150 ;
        RECT 248.100 124.050 249.900 125.850 ;
        RECT 254.100 124.050 255.900 125.850 ;
        RECT 242.850 118.800 246.450 119.700 ;
        RECT 257.550 119.700 258.750 127.050 ;
        RECT 259.950 125.850 262.050 127.950 ;
        RECT 271.950 125.850 274.050 127.950 ;
        RECT 274.950 127.050 277.050 129.150 ;
        RECT 260.100 124.050 261.900 125.850 ;
        RECT 272.100 124.050 273.900 125.850 ;
        RECT 275.250 119.700 276.450 127.050 ;
        RECT 277.950 125.850 280.050 127.950 ;
        RECT 283.950 125.850 286.050 127.950 ;
        RECT 286.950 127.050 289.050 129.150 ;
        RECT 278.100 124.050 279.900 125.850 ;
        RECT 284.100 124.050 285.900 125.850 ;
        RECT 287.250 119.700 288.450 127.050 ;
        RECT 289.950 125.850 292.050 127.950 ;
        RECT 299.100 126.150 300.900 127.950 ;
        RECT 290.100 124.050 291.900 125.850 ;
        RECT 298.950 124.050 301.050 126.150 ;
        RECT 302.700 120.300 303.900 137.400 ;
        RECT 306.150 131.400 307.950 143.250 ;
        RECT 309.150 131.400 310.950 143.250 ;
        RECT 317.550 137.400 319.350 143.250 ;
        RECT 320.550 137.400 322.350 143.250 ;
        RECT 335.400 137.400 337.200 143.250 ;
        RECT 304.950 125.850 307.050 127.950 ;
        RECT 309.150 126.150 310.350 131.400 ;
        RECT 305.100 124.050 306.900 125.850 ;
        RECT 307.950 124.050 310.350 126.150 ;
        RECT 320.400 124.950 321.600 137.400 ;
        RECT 331.950 130.950 334.050 133.050 ;
        RECT 338.700 131.400 340.500 143.250 ;
        RECT 342.900 131.400 344.700 143.250 ;
        RECT 348.300 131.400 350.100 143.250 ;
        RECT 352.500 131.400 354.300 143.250 ;
        RECT 355.800 137.400 357.600 143.250 ;
        RECT 371.400 137.400 373.200 143.250 ;
        RECT 358.950 133.950 361.050 136.050 ;
        RECT 257.550 118.800 261.150 119.700 ;
        RECT 242.850 111.750 244.650 118.800 ;
        RECT 247.350 111.750 249.150 117.600 ;
        RECT 254.850 111.750 256.650 117.600 ;
        RECT 259.350 111.750 261.150 118.800 ;
        RECT 272.850 118.800 276.450 119.700 ;
        RECT 284.850 118.800 288.450 119.700 ;
        RECT 299.550 119.100 307.050 120.300 ;
        RECT 272.850 111.750 274.650 118.800 ;
        RECT 277.350 111.750 279.150 117.600 ;
        RECT 284.850 111.750 286.650 118.800 ;
        RECT 289.350 111.750 291.150 117.600 ;
        RECT 299.550 111.750 301.350 119.100 ;
        RECT 305.250 118.500 307.050 119.100 ;
        RECT 309.150 117.600 310.350 124.050 ;
        RECT 317.100 123.150 318.900 124.950 ;
        RECT 316.950 121.050 319.050 123.150 ;
        RECT 319.950 122.850 322.050 124.950 ;
        RECT 332.550 123.450 333.450 130.950 ;
        RECT 335.250 129.150 337.050 130.950 ;
        RECT 334.950 127.050 337.050 129.150 ;
        RECT 338.850 126.150 340.050 131.400 ;
        RECT 344.100 126.150 345.900 127.950 ;
        RECT 347.100 126.150 348.900 127.950 ;
        RECT 352.950 126.150 354.150 131.400 ;
        RECT 355.950 129.150 357.750 130.950 ;
        RECT 355.950 127.050 358.050 129.150 ;
        RECT 337.950 124.050 340.050 126.150 ;
        RECT 334.950 123.450 337.050 124.050 ;
        RECT 304.050 111.750 305.850 117.600 ;
        RECT 307.050 116.100 310.350 117.600 ;
        RECT 307.050 111.750 308.850 116.100 ;
        RECT 320.400 114.600 321.600 122.850 ;
        RECT 332.550 122.550 337.050 123.450 ;
        RECT 334.950 121.950 337.050 122.550 ;
        RECT 337.950 120.750 339.150 124.050 ;
        RECT 340.950 122.850 343.050 124.950 ;
        RECT 343.950 124.050 346.050 126.150 ;
        RECT 346.950 124.050 349.050 126.150 ;
        RECT 349.950 122.850 352.050 124.950 ;
        RECT 352.950 124.050 355.050 126.150 ;
        RECT 341.100 121.050 342.900 122.850 ;
        RECT 350.100 121.050 351.900 122.850 ;
        RECT 353.850 120.750 355.050 124.050 ;
        RECT 355.950 123.450 358.050 124.050 ;
        RECT 359.550 123.450 360.450 133.950 ;
        RECT 374.700 131.400 376.500 143.250 ;
        RECT 378.900 131.400 380.700 143.250 ;
        RECT 383.550 137.400 385.350 143.250 ;
        RECT 386.550 137.400 388.350 143.250 ;
        RECT 389.550 138.000 391.350 143.250 ;
        RECT 386.700 137.100 388.350 137.400 ;
        RECT 392.550 137.400 394.350 143.250 ;
        RECT 400.650 137.400 402.450 143.250 ;
        RECT 403.650 138.000 405.450 143.250 ;
        RECT 392.550 137.100 393.750 137.400 ;
        RECT 386.700 136.200 393.750 137.100 ;
        RECT 386.100 132.150 387.900 133.950 ;
        RECT 364.950 129.450 367.050 130.050 ;
        RECT 364.950 128.550 369.450 129.450 ;
        RECT 371.250 129.150 373.050 130.950 ;
        RECT 364.950 127.950 367.050 128.550 ;
        RECT 355.950 122.550 360.450 123.450 ;
        RECT 368.550 123.450 369.450 128.550 ;
        RECT 370.950 127.050 373.050 129.150 ;
        RECT 374.850 126.150 376.050 131.400 ;
        RECT 383.100 129.150 384.900 130.950 ;
        RECT 385.950 130.050 388.050 132.150 ;
        RECT 389.250 129.150 391.050 130.950 ;
        RECT 380.100 126.150 381.900 127.950 ;
        RECT 382.950 127.050 385.050 129.150 ;
        RECT 388.950 127.050 391.050 129.150 ;
        RECT 392.700 127.950 393.750 136.200 ;
        RECT 401.250 137.100 402.450 137.400 ;
        RECT 406.650 137.400 408.450 143.250 ;
        RECT 409.650 137.400 411.450 143.250 ;
        RECT 406.650 137.100 408.300 137.400 ;
        RECT 401.250 136.200 408.300 137.100 ;
        RECT 401.250 127.950 402.300 136.200 ;
        RECT 407.100 132.150 408.900 133.950 ;
        RECT 403.950 129.150 405.750 130.950 ;
        RECT 406.950 130.050 409.050 132.150 ;
        RECT 419.550 131.400 421.350 143.250 ;
        RECT 423.750 131.400 425.550 143.250 ;
        RECT 439.650 131.400 441.450 143.250 ;
        RECT 442.650 131.400 444.450 143.250 ;
        RECT 455.400 137.400 457.200 143.250 ;
        RECT 458.700 131.400 460.500 143.250 ;
        RECT 462.900 131.400 464.700 143.250 ;
        RECT 471.300 131.400 473.100 143.250 ;
        RECT 475.500 131.400 477.300 143.250 ;
        RECT 478.800 137.400 480.600 143.250 ;
        RECT 488.400 137.400 490.200 143.250 ;
        RECT 410.100 129.150 411.900 130.950 ;
        RECT 423.000 130.350 425.550 131.400 ;
        RECT 373.950 124.050 376.050 126.150 ;
        RECT 370.950 123.450 373.050 124.050 ;
        RECT 368.550 122.550 373.050 123.450 ;
        RECT 355.950 121.950 358.050 122.550 ;
        RECT 370.950 121.950 373.050 122.550 ;
        RECT 373.950 120.750 375.150 124.050 ;
        RECT 376.950 122.850 379.050 124.950 ;
        RECT 379.950 124.050 382.050 126.150 ;
        RECT 391.950 125.850 394.050 127.950 ;
        RECT 400.950 125.850 403.050 127.950 ;
        RECT 403.950 127.050 406.050 129.150 ;
        RECT 409.950 127.050 412.050 129.150 ;
        RECT 419.100 126.150 420.900 127.950 ;
        RECT 377.100 121.050 378.900 122.850 ;
        RECT 392.400 121.650 393.600 125.850 ;
        RECT 335.250 119.700 339.000 120.750 ;
        RECT 354.000 119.700 357.750 120.750 ;
        RECT 335.250 117.600 336.450 119.700 ;
        RECT 317.550 111.750 319.350 114.600 ;
        RECT 320.550 111.750 322.350 114.600 ;
        RECT 334.650 111.750 336.450 117.600 ;
        RECT 337.650 116.700 345.450 118.050 ;
        RECT 337.650 111.750 339.450 116.700 ;
        RECT 340.650 111.750 342.450 115.800 ;
        RECT 343.650 111.750 345.450 116.700 ;
        RECT 347.550 116.700 355.350 118.050 ;
        RECT 347.550 111.750 349.350 116.700 ;
        RECT 350.550 111.750 352.350 115.800 ;
        RECT 353.550 111.750 355.350 116.700 ;
        RECT 356.550 117.600 357.750 119.700 ;
        RECT 371.250 119.700 375.000 120.750 ;
        RECT 371.250 117.600 372.450 119.700 ;
        RECT 356.550 111.750 358.350 117.600 ;
        RECT 370.650 111.750 372.450 117.600 ;
        RECT 373.650 116.700 381.450 118.050 ;
        RECT 373.650 111.750 375.450 116.700 ;
        RECT 376.650 111.750 378.450 115.800 ;
        RECT 379.650 111.750 381.450 116.700 ;
        RECT 383.700 111.750 385.500 120.600 ;
        RECT 389.100 120.000 393.600 121.650 ;
        RECT 401.400 121.650 402.600 125.850 ;
        RECT 418.950 124.050 421.050 126.150 ;
        RECT 423.000 123.150 424.050 130.350 ;
        RECT 425.100 126.150 426.900 127.950 ;
        RECT 440.400 126.150 441.600 131.400 ;
        RECT 455.250 129.150 457.050 130.950 ;
        RECT 454.950 127.050 457.050 129.150 ;
        RECT 458.850 126.150 460.050 131.400 ;
        RECT 464.100 126.150 465.900 127.950 ;
        RECT 470.100 126.150 471.900 127.950 ;
        RECT 475.950 126.150 477.150 131.400 ;
        RECT 484.950 130.950 487.050 133.050 ;
        RECT 491.700 131.400 493.500 143.250 ;
        RECT 495.900 131.400 497.700 143.250 ;
        RECT 503.550 137.400 505.350 143.250 ;
        RECT 506.550 137.400 508.350 143.250 ;
        RECT 509.550 137.400 511.350 143.250 ;
        RECT 518.550 137.400 520.350 143.250 ;
        RECT 521.550 137.400 523.350 143.250 ;
        RECT 524.550 137.400 526.350 143.250 ;
        RECT 536.400 137.400 538.200 143.250 ;
        RECT 478.950 129.150 480.750 130.950 ;
        RECT 478.950 127.050 481.050 129.150 ;
        RECT 424.950 124.050 427.050 126.150 ;
        RECT 439.950 124.050 442.050 126.150 ;
        RECT 401.400 120.000 405.900 121.650 ;
        RECT 421.950 121.050 424.050 123.150 ;
        RECT 389.100 111.750 390.900 120.000 ;
        RECT 404.100 111.750 405.900 120.000 ;
        RECT 409.500 111.750 411.300 120.600 ;
        RECT 423.000 114.600 424.050 121.050 ;
        RECT 440.400 117.600 441.600 124.050 ;
        RECT 442.950 122.850 445.050 124.950 ;
        RECT 457.950 124.050 460.050 126.150 ;
        RECT 443.100 121.050 444.900 122.850 ;
        RECT 457.950 120.750 459.150 124.050 ;
        RECT 460.950 122.850 463.050 124.950 ;
        RECT 463.950 124.050 466.050 126.150 ;
        RECT 469.950 124.050 472.050 126.150 ;
        RECT 472.950 122.850 475.050 124.950 ;
        RECT 475.950 124.050 478.050 126.150 ;
        RECT 461.100 121.050 462.900 122.850 ;
        RECT 473.100 121.050 474.900 122.850 ;
        RECT 455.250 119.700 459.000 120.750 ;
        RECT 463.950 120.450 466.050 121.050 ;
        RECT 469.950 120.450 472.050 121.050 ;
        RECT 476.850 120.750 478.050 124.050 ;
        RECT 478.950 123.450 481.050 124.050 ;
        RECT 485.550 123.450 486.450 130.950 ;
        RECT 488.250 129.150 490.050 130.950 ;
        RECT 487.950 127.050 490.050 129.150 ;
        RECT 491.850 126.150 493.050 131.400 ;
        RECT 506.550 129.150 507.750 137.400 ;
        RECT 521.550 129.150 522.750 137.400 ;
        RECT 539.700 131.400 541.500 143.250 ;
        RECT 543.900 131.400 545.700 143.250 ;
        RECT 548.550 137.400 550.350 143.250 ;
        RECT 551.550 137.400 553.350 143.250 ;
        RECT 554.550 138.000 556.350 143.250 ;
        RECT 551.700 137.100 553.350 137.400 ;
        RECT 557.550 137.400 559.350 143.250 ;
        RECT 569.550 137.400 571.350 143.250 ;
        RECT 572.550 137.400 574.350 143.250 ;
        RECT 557.550 137.100 558.750 137.400 ;
        RECT 551.700 136.200 558.750 137.100 ;
        RECT 551.100 132.150 552.900 133.950 ;
        RECT 536.250 129.150 538.050 130.950 ;
        RECT 497.100 126.150 498.900 127.950 ;
        RECT 478.950 122.550 486.450 123.450 ;
        RECT 490.950 124.050 493.050 126.150 ;
        RECT 478.950 121.950 481.050 122.550 ;
        RECT 490.950 120.750 492.150 124.050 ;
        RECT 493.950 122.850 496.050 124.950 ;
        RECT 496.950 124.050 499.050 126.150 ;
        RECT 502.950 125.850 505.050 127.950 ;
        RECT 505.950 127.050 508.050 129.150 ;
        RECT 503.100 124.050 504.900 125.850 ;
        RECT 494.100 121.050 495.900 122.850 ;
        RECT 455.250 117.600 456.450 119.700 ;
        RECT 463.950 119.550 472.050 120.450 ;
        RECT 477.000 119.700 480.750 120.750 ;
        RECT 463.950 118.950 466.050 119.550 ;
        RECT 469.950 118.950 472.050 119.550 ;
        RECT 419.550 111.750 421.350 114.600 ;
        RECT 422.550 111.750 424.350 114.600 ;
        RECT 425.550 111.750 427.350 114.600 ;
        RECT 439.650 111.750 441.450 117.600 ;
        RECT 442.650 111.750 444.450 117.600 ;
        RECT 454.650 111.750 456.450 117.600 ;
        RECT 457.650 116.700 465.450 118.050 ;
        RECT 457.650 111.750 459.450 116.700 ;
        RECT 460.650 111.750 462.450 115.800 ;
        RECT 463.650 111.750 465.450 116.700 ;
        RECT 470.550 116.700 478.350 118.050 ;
        RECT 470.550 111.750 472.350 116.700 ;
        RECT 473.550 111.750 475.350 115.800 ;
        RECT 476.550 111.750 478.350 116.700 ;
        RECT 479.550 117.600 480.750 119.700 ;
        RECT 488.250 119.700 492.000 120.750 ;
        RECT 506.550 119.700 507.750 127.050 ;
        RECT 508.950 125.850 511.050 127.950 ;
        RECT 517.950 125.850 520.050 127.950 ;
        RECT 520.950 127.050 523.050 129.150 ;
        RECT 509.100 124.050 510.900 125.850 ;
        RECT 518.100 124.050 519.900 125.850 ;
        RECT 521.550 119.700 522.750 127.050 ;
        RECT 523.950 125.850 526.050 127.950 ;
        RECT 535.950 127.050 538.050 129.150 ;
        RECT 539.850 126.150 541.050 131.400 ;
        RECT 548.100 129.150 549.900 130.950 ;
        RECT 550.950 130.050 553.050 132.150 ;
        RECT 554.250 129.150 556.050 130.950 ;
        RECT 545.100 126.150 546.900 127.950 ;
        RECT 547.950 127.050 550.050 129.150 ;
        RECT 553.950 127.050 556.050 129.150 ;
        RECT 557.700 127.950 558.750 136.200 ;
        RECT 559.950 132.450 562.050 133.050 ;
        RECT 568.950 132.450 571.050 133.050 ;
        RECT 559.950 131.550 571.050 132.450 ;
        RECT 559.950 130.950 562.050 131.550 ;
        RECT 568.950 130.950 571.050 131.550 ;
        RECT 524.100 124.050 525.900 125.850 ;
        RECT 538.950 124.050 541.050 126.150 ;
        RECT 538.950 120.750 540.150 124.050 ;
        RECT 541.950 122.850 544.050 124.950 ;
        RECT 544.950 124.050 547.050 126.150 ;
        RECT 556.950 125.850 559.050 127.950 ;
        RECT 569.100 126.150 570.900 127.950 ;
        RECT 542.100 121.050 543.900 122.850 ;
        RECT 557.400 121.650 558.600 125.850 ;
        RECT 568.950 124.050 571.050 126.150 ;
        RECT 536.250 119.700 540.000 120.750 ;
        RECT 488.250 117.600 489.450 119.700 ;
        RECT 506.550 118.800 510.150 119.700 ;
        RECT 521.550 118.800 525.150 119.700 ;
        RECT 479.550 111.750 481.350 117.600 ;
        RECT 487.650 111.750 489.450 117.600 ;
        RECT 490.650 116.700 498.450 118.050 ;
        RECT 490.650 111.750 492.450 116.700 ;
        RECT 493.650 111.750 495.450 115.800 ;
        RECT 496.650 111.750 498.450 116.700 ;
        RECT 503.850 111.750 505.650 117.600 ;
        RECT 508.350 111.750 510.150 118.800 ;
        RECT 518.850 111.750 520.650 117.600 ;
        RECT 523.350 111.750 525.150 118.800 ;
        RECT 536.250 117.600 537.450 119.700 ;
        RECT 535.650 111.750 537.450 117.600 ;
        RECT 538.650 116.700 546.450 118.050 ;
        RECT 538.650 111.750 540.450 116.700 ;
        RECT 541.650 111.750 543.450 115.800 ;
        RECT 544.650 111.750 546.450 116.700 ;
        RECT 548.700 111.750 550.500 120.600 ;
        RECT 554.100 120.000 558.600 121.650 ;
        RECT 572.700 120.300 573.900 137.400 ;
        RECT 576.150 131.400 577.950 143.250 ;
        RECT 579.150 131.400 580.950 143.250 ;
        RECT 590.550 137.400 592.350 143.250 ;
        RECT 593.550 137.400 595.350 143.250 ;
        RECT 596.550 138.000 598.350 143.250 ;
        RECT 593.700 137.100 595.350 137.400 ;
        RECT 599.550 137.400 601.350 143.250 ;
        RECT 607.650 137.400 609.450 143.250 ;
        RECT 610.650 137.400 612.450 143.250 ;
        RECT 613.650 137.400 615.450 143.250 ;
        RECT 620.550 137.400 622.350 143.250 ;
        RECT 623.550 137.400 625.350 143.250 ;
        RECT 599.550 137.100 600.750 137.400 ;
        RECT 593.700 136.200 600.750 137.100 ;
        RECT 593.100 132.150 594.900 133.950 ;
        RECT 574.950 125.850 577.050 127.950 ;
        RECT 579.150 126.150 580.350 131.400 ;
        RECT 590.100 129.150 591.900 130.950 ;
        RECT 592.950 130.050 595.050 132.150 ;
        RECT 596.250 129.150 598.050 130.950 ;
        RECT 589.950 127.050 592.050 129.150 ;
        RECT 595.950 127.050 598.050 129.150 ;
        RECT 599.700 127.950 600.750 136.200 ;
        RECT 611.250 129.150 612.450 137.400 ;
        RECT 575.100 124.050 576.900 125.850 ;
        RECT 577.950 124.050 580.350 126.150 ;
        RECT 598.950 125.850 601.050 127.950 ;
        RECT 607.950 125.850 610.050 127.950 ;
        RECT 610.950 127.050 613.050 129.150 ;
        RECT 554.100 111.750 555.900 120.000 ;
        RECT 569.550 119.100 577.050 120.300 ;
        RECT 569.550 111.750 571.350 119.100 ;
        RECT 575.250 118.500 577.050 119.100 ;
        RECT 579.150 117.600 580.350 124.050 ;
        RECT 599.400 121.650 600.600 125.850 ;
        RECT 608.100 124.050 609.900 125.850 ;
        RECT 574.050 111.750 575.850 117.600 ;
        RECT 577.050 116.100 580.350 117.600 ;
        RECT 577.050 111.750 578.850 116.100 ;
        RECT 590.700 111.750 592.500 120.600 ;
        RECT 596.100 120.000 600.600 121.650 ;
        RECT 596.100 111.750 597.900 120.000 ;
        RECT 611.250 119.700 612.450 127.050 ;
        RECT 613.950 125.850 616.050 127.950 ;
        RECT 620.100 126.150 621.900 127.950 ;
        RECT 614.100 124.050 615.900 125.850 ;
        RECT 619.950 124.050 622.050 126.150 ;
        RECT 623.700 120.300 624.900 137.400 ;
        RECT 627.150 131.400 628.950 143.250 ;
        RECT 630.150 131.400 631.950 143.250 ;
        RECT 640.650 137.400 642.450 143.250 ;
        RECT 643.650 138.000 645.450 143.250 ;
        RECT 641.250 137.100 642.450 137.400 ;
        RECT 646.650 137.400 648.450 143.250 ;
        RECT 649.650 137.400 651.450 143.250 ;
        RECT 656.550 137.400 658.350 143.250 ;
        RECT 659.550 137.400 661.350 143.250 ;
        RECT 662.550 138.000 664.350 143.250 ;
        RECT 646.650 137.100 648.300 137.400 ;
        RECT 641.250 136.200 648.300 137.100 ;
        RECT 659.700 137.100 661.350 137.400 ;
        RECT 665.550 137.400 667.350 143.250 ;
        RECT 665.550 137.100 666.750 137.400 ;
        RECT 659.700 136.200 666.750 137.100 ;
        RECT 625.950 125.850 628.050 127.950 ;
        RECT 630.150 126.150 631.350 131.400 ;
        RECT 641.250 127.950 642.300 136.200 ;
        RECT 647.100 132.150 648.900 133.950 ;
        RECT 659.100 132.150 660.900 133.950 ;
        RECT 643.950 129.150 645.750 130.950 ;
        RECT 646.950 130.050 649.050 132.150 ;
        RECT 650.100 129.150 651.900 130.950 ;
        RECT 656.100 129.150 657.900 130.950 ;
        RECT 658.950 130.050 661.050 132.150 ;
        RECT 662.250 129.150 664.050 130.950 ;
        RECT 626.100 124.050 627.900 125.850 ;
        RECT 628.950 124.050 631.350 126.150 ;
        RECT 640.950 125.850 643.050 127.950 ;
        RECT 643.950 127.050 646.050 129.150 ;
        RECT 649.950 127.050 652.050 129.150 ;
        RECT 655.950 127.050 658.050 129.150 ;
        RECT 661.950 127.050 664.050 129.150 ;
        RECT 665.700 127.950 666.750 136.200 ;
        RECT 676.650 131.400 678.450 143.250 ;
        RECT 679.650 132.300 681.450 143.250 ;
        RECT 682.650 133.200 684.450 143.250 ;
        RECT 685.650 132.300 687.450 143.250 ;
        RECT 692.550 137.400 694.350 143.250 ;
        RECT 695.550 137.400 697.350 143.250 ;
        RECT 698.550 137.400 700.350 143.250 ;
        RECT 706.650 137.400 708.450 143.250 ;
        RECT 709.650 137.400 711.450 143.250 ;
        RECT 712.650 137.400 714.450 143.250 ;
        RECT 721.650 137.400 723.450 143.250 ;
        RECT 724.650 137.400 726.450 143.250 ;
        RECT 727.650 137.400 729.450 143.250 ;
        RECT 737.550 137.400 739.350 143.250 ;
        RECT 740.550 137.400 742.350 143.250 ;
        RECT 743.550 137.400 745.350 143.250 ;
        RECT 679.650 131.400 687.450 132.300 ;
        RECT 664.950 125.850 667.050 127.950 ;
        RECT 677.100 126.150 678.300 131.400 ;
        RECT 695.550 129.150 696.750 137.400 ;
        RECT 710.250 129.150 711.450 137.400 ;
        RECT 718.950 130.950 721.050 133.050 ;
        RECT 608.850 118.800 612.450 119.700 ;
        RECT 620.550 119.100 628.050 120.300 ;
        RECT 608.850 111.750 610.650 118.800 ;
        RECT 613.350 111.750 615.150 117.600 ;
        RECT 620.550 111.750 622.350 119.100 ;
        RECT 626.250 118.500 628.050 119.100 ;
        RECT 630.150 117.600 631.350 124.050 ;
        RECT 641.400 121.650 642.600 125.850 ;
        RECT 665.400 121.650 666.600 125.850 ;
        RECT 676.950 124.050 679.050 126.150 ;
        RECT 691.950 125.850 694.050 127.950 ;
        RECT 694.950 127.050 697.050 129.150 ;
        RECT 641.400 120.000 645.900 121.650 ;
        RECT 625.050 111.750 626.850 117.600 ;
        RECT 628.050 116.100 631.350 117.600 ;
        RECT 628.050 111.750 629.850 116.100 ;
        RECT 644.100 111.750 645.900 120.000 ;
        RECT 649.500 111.750 651.300 120.600 ;
        RECT 656.700 111.750 658.500 120.600 ;
        RECT 662.100 120.000 666.600 121.650 ;
        RECT 662.100 111.750 663.900 120.000 ;
        RECT 677.100 117.600 678.300 124.050 ;
        RECT 679.950 122.850 682.050 124.950 ;
        RECT 683.100 123.150 684.900 124.950 ;
        RECT 680.100 121.050 681.900 122.850 ;
        RECT 682.950 121.050 685.050 123.150 ;
        RECT 685.950 122.850 688.050 124.950 ;
        RECT 692.100 124.050 693.900 125.850 ;
        RECT 686.100 121.050 687.900 122.850 ;
        RECT 695.550 119.700 696.750 127.050 ;
        RECT 697.950 125.850 700.050 127.950 ;
        RECT 706.950 125.850 709.050 127.950 ;
        RECT 709.950 127.050 712.050 129.150 ;
        RECT 698.100 124.050 699.900 125.850 ;
        RECT 707.100 124.050 708.900 125.850 ;
        RECT 710.250 119.700 711.450 127.050 ;
        RECT 712.950 125.850 715.050 127.950 ;
        RECT 713.100 124.050 714.900 125.850 ;
        RECT 719.550 121.050 720.450 130.950 ;
        RECT 725.250 129.150 726.450 137.400 ;
        RECT 740.550 129.150 741.750 137.400 ;
        RECT 759.450 131.400 761.250 143.250 ;
        RECT 763.650 131.400 765.450 143.250 ;
        RECT 774.300 131.400 776.100 143.250 ;
        RECT 778.500 131.400 780.300 143.250 ;
        RECT 781.800 137.400 783.600 143.250 ;
        RECT 796.650 137.400 798.450 143.250 ;
        RECT 799.650 138.000 801.450 143.250 ;
        RECT 797.250 137.100 798.450 137.400 ;
        RECT 802.650 137.400 804.450 143.250 ;
        RECT 805.650 137.400 807.450 143.250 ;
        RECT 802.650 137.100 804.300 137.400 ;
        RECT 797.250 136.200 804.300 137.100 ;
        RECT 759.450 130.350 762.000 131.400 ;
        RECT 721.950 125.850 724.050 127.950 ;
        RECT 724.950 127.050 727.050 129.150 ;
        RECT 722.100 124.050 723.900 125.850 ;
        RECT 695.550 118.800 699.150 119.700 ;
        RECT 677.100 115.950 682.800 117.600 ;
        RECT 677.700 111.750 679.500 114.600 ;
        RECT 681.000 111.750 682.800 115.950 ;
        RECT 685.200 111.750 687.000 117.600 ;
        RECT 692.850 111.750 694.650 117.600 ;
        RECT 697.350 111.750 699.150 118.800 ;
        RECT 707.850 118.800 711.450 119.700 ;
        RECT 718.950 118.950 721.050 121.050 ;
        RECT 725.250 119.700 726.450 127.050 ;
        RECT 727.950 125.850 730.050 127.950 ;
        RECT 736.950 125.850 739.050 127.950 ;
        RECT 739.950 127.050 742.050 129.150 ;
        RECT 728.100 124.050 729.900 125.850 ;
        RECT 737.100 124.050 738.900 125.850 ;
        RECT 722.850 118.800 726.450 119.700 ;
        RECT 740.550 119.700 741.750 127.050 ;
        RECT 742.950 125.850 745.050 127.950 ;
        RECT 758.100 126.150 759.900 127.950 ;
        RECT 743.100 124.050 744.900 125.850 ;
        RECT 757.950 124.050 760.050 126.150 ;
        RECT 760.950 123.150 762.000 130.350 ;
        RECT 764.100 126.150 765.900 127.950 ;
        RECT 773.100 126.150 774.900 127.950 ;
        RECT 778.950 126.150 780.150 131.400 ;
        RECT 781.950 129.150 783.750 130.950 ;
        RECT 781.950 127.050 784.050 129.150 ;
        RECT 797.250 127.950 798.300 136.200 ;
        RECT 803.100 132.150 804.900 133.950 ;
        RECT 799.950 129.150 801.750 130.950 ;
        RECT 802.950 130.050 805.050 132.150 ;
        RECT 809.550 131.400 811.350 143.250 ;
        RECT 813.750 131.400 815.550 143.250 ;
        RECT 806.100 129.150 807.900 130.950 ;
        RECT 813.000 130.350 815.550 131.400 ;
        RECT 821.550 131.400 823.350 143.250 ;
        RECT 826.050 131.550 827.850 143.250 ;
        RECT 829.050 132.900 830.850 143.250 ;
        RECT 842.550 137.400 844.350 143.250 ;
        RECT 845.550 137.400 847.350 143.250 ;
        RECT 829.050 131.550 831.450 132.900 ;
        RECT 763.950 124.050 766.050 126.150 ;
        RECT 772.950 124.050 775.050 126.150 ;
        RECT 760.950 121.050 763.050 123.150 ;
        RECT 775.950 122.850 778.050 124.950 ;
        RECT 778.950 124.050 781.050 126.150 ;
        RECT 796.950 125.850 799.050 127.950 ;
        RECT 799.950 127.050 802.050 129.150 ;
        RECT 805.950 127.050 808.050 129.150 ;
        RECT 809.100 126.150 810.900 127.950 ;
        RECT 776.100 121.050 777.900 122.850 ;
        RECT 740.550 118.800 744.150 119.700 ;
        RECT 707.850 111.750 709.650 118.800 ;
        RECT 712.350 111.750 714.150 117.600 ;
        RECT 722.850 111.750 724.650 118.800 ;
        RECT 727.350 111.750 729.150 117.600 ;
        RECT 737.850 111.750 739.650 117.600 ;
        RECT 742.350 111.750 744.150 118.800 ;
        RECT 760.950 114.600 762.000 121.050 ;
        RECT 779.850 120.750 781.050 124.050 ;
        RECT 797.400 121.650 798.600 125.850 ;
        RECT 808.950 124.050 811.050 126.150 ;
        RECT 813.000 123.150 814.050 130.350 ;
        RECT 821.550 130.200 822.750 131.400 ;
        RECT 826.950 130.200 828.750 130.650 ;
        RECT 821.550 129.000 828.750 130.200 ;
        RECT 826.950 128.850 828.750 129.000 ;
        RECT 815.100 126.150 816.900 127.950 ;
        RECT 824.100 126.150 825.900 127.950 ;
        RECT 814.950 124.050 817.050 126.150 ;
        RECT 821.100 123.150 822.900 124.950 ;
        RECT 823.950 124.050 826.050 126.150 ;
        RECT 780.000 119.700 783.750 120.750 ;
        RECT 797.400 120.000 801.900 121.650 ;
        RECT 811.950 121.050 814.050 123.150 ;
        RECT 820.950 121.050 823.050 123.150 ;
        RECT 773.550 116.700 781.350 118.050 ;
        RECT 757.650 111.750 759.450 114.600 ;
        RECT 760.650 111.750 762.450 114.600 ;
        RECT 763.650 111.750 765.450 114.600 ;
        RECT 773.550 111.750 775.350 116.700 ;
        RECT 776.550 111.750 778.350 115.800 ;
        RECT 779.550 111.750 781.350 116.700 ;
        RECT 782.550 117.600 783.750 119.700 ;
        RECT 782.550 111.750 784.350 117.600 ;
        RECT 800.100 111.750 801.900 120.000 ;
        RECT 805.500 111.750 807.300 120.600 ;
        RECT 813.000 114.600 814.050 121.050 ;
        RECT 827.700 120.600 828.600 128.850 ;
        RECT 830.100 124.950 831.450 131.550 ;
        RECT 845.400 124.950 846.600 137.400 ;
        RECT 829.950 122.850 832.050 124.950 ;
        RECT 842.100 123.150 843.900 124.950 ;
        RECT 826.950 119.700 828.750 120.600 ;
        RECT 825.450 118.800 828.750 119.700 ;
        RECT 825.450 114.600 826.350 118.800 ;
        RECT 831.000 117.600 832.050 122.850 ;
        RECT 841.950 121.050 844.050 123.150 ;
        RECT 844.950 122.850 847.050 124.950 ;
        RECT 809.550 111.750 811.350 114.600 ;
        RECT 812.550 111.750 814.350 114.600 ;
        RECT 815.550 111.750 817.350 114.600 ;
        RECT 821.550 111.750 823.350 114.600 ;
        RECT 824.550 111.750 826.350 114.600 ;
        RECT 827.550 111.750 829.350 114.600 ;
        RECT 830.550 111.750 832.350 117.600 ;
        RECT 845.400 114.600 846.600 122.850 ;
        RECT 842.550 111.750 844.350 114.600 ;
        RECT 845.550 111.750 847.350 114.600 ;
        RECT 11.850 100.200 13.650 107.250 ;
        RECT 16.350 101.400 18.150 107.250 ;
        RECT 23.850 100.200 25.650 107.250 ;
        RECT 28.350 101.400 30.150 107.250 ;
        RECT 38.850 101.400 40.650 107.250 ;
        RECT 43.350 100.200 45.150 107.250 ;
        RECT 11.850 99.300 15.450 100.200 ;
        RECT 23.850 99.300 27.450 100.200 ;
        RECT 11.100 93.150 12.900 94.950 ;
        RECT 10.950 91.050 13.050 93.150 ;
        RECT 14.250 91.950 15.450 99.300 ;
        RECT 17.100 93.150 18.900 94.950 ;
        RECT 23.100 93.150 24.900 94.950 ;
        RECT 13.950 89.850 16.050 91.950 ;
        RECT 16.950 91.050 19.050 93.150 ;
        RECT 22.950 91.050 25.050 93.150 ;
        RECT 26.250 91.950 27.450 99.300 ;
        RECT 41.550 99.300 45.150 100.200 ;
        RECT 29.100 93.150 30.900 94.950 ;
        RECT 38.100 93.150 39.900 94.950 ;
        RECT 25.950 89.850 28.050 91.950 ;
        RECT 28.950 91.050 31.050 93.150 ;
        RECT 37.950 91.050 40.050 93.150 ;
        RECT 41.550 91.950 42.750 99.300 ;
        RECT 59.100 99.000 60.900 107.250 ;
        RECT 56.400 97.350 60.900 99.000 ;
        RECT 64.500 98.400 66.300 107.250 ;
        RECT 68.550 102.300 70.350 107.250 ;
        RECT 71.550 103.200 73.350 107.250 ;
        RECT 74.550 102.300 76.350 107.250 ;
        RECT 68.550 100.950 76.350 102.300 ;
        RECT 77.550 101.400 79.350 107.250 ;
        RECT 83.550 104.400 85.350 107.250 ;
        RECT 86.550 104.400 88.350 107.250 ;
        RECT 89.550 104.400 91.350 107.250 ;
        RECT 77.550 99.300 78.750 101.400 ;
        RECT 75.000 98.250 78.750 99.300 ;
        RECT 44.100 93.150 45.900 94.950 ;
        RECT 56.400 93.150 57.600 97.350 ;
        RECT 71.100 96.150 72.900 97.950 ;
        RECT 40.950 89.850 43.050 91.950 ;
        RECT 43.950 91.050 46.050 93.150 ;
        RECT 55.950 91.050 58.050 93.150 ;
        RECT 67.950 92.850 70.050 94.950 ;
        RECT 70.950 94.050 73.050 96.150 ;
        RECT 74.850 94.950 76.050 98.250 ;
        RECT 87.000 97.950 88.050 104.400 ;
        RECT 101.550 102.300 103.350 107.250 ;
        RECT 104.550 103.200 106.350 107.250 ;
        RECT 107.550 102.300 109.350 107.250 ;
        RECT 101.550 100.950 109.350 102.300 ;
        RECT 110.550 101.400 112.350 107.250 ;
        RECT 124.650 104.400 126.450 107.250 ;
        RECT 127.650 104.400 129.450 107.250 ;
        RECT 110.550 99.300 111.750 101.400 ;
        RECT 108.000 98.250 111.750 99.300 ;
        RECT 85.950 95.850 88.050 97.950 ;
        RECT 104.100 96.150 105.900 97.950 ;
        RECT 73.950 92.850 76.050 94.950 ;
        RECT 82.950 92.850 85.050 94.950 ;
        RECT 14.250 81.600 15.450 89.850 ;
        RECT 26.250 81.600 27.450 89.850 ;
        RECT 41.550 81.600 42.750 89.850 ;
        RECT 56.250 82.800 57.300 91.050 ;
        RECT 58.950 89.850 61.050 91.950 ;
        RECT 64.950 89.850 67.050 91.950 ;
        RECT 68.100 91.050 69.900 92.850 ;
        RECT 58.950 88.050 60.750 89.850 ;
        RECT 61.950 86.850 64.050 88.950 ;
        RECT 65.100 88.050 66.900 89.850 ;
        RECT 73.950 87.600 75.150 92.850 ;
        RECT 76.950 89.850 79.050 91.950 ;
        RECT 83.100 91.050 84.900 92.850 ;
        RECT 76.950 88.050 78.750 89.850 ;
        RECT 87.000 88.650 88.050 95.850 ;
        RECT 88.950 92.850 91.050 94.950 ;
        RECT 100.950 92.850 103.050 94.950 ;
        RECT 103.950 94.050 106.050 96.150 ;
        RECT 107.850 94.950 109.050 98.250 ;
        RECT 125.400 96.150 126.600 104.400 ;
        RECT 134.550 102.300 136.350 107.250 ;
        RECT 137.550 103.200 139.350 107.250 ;
        RECT 140.550 102.300 142.350 107.250 ;
        RECT 134.550 100.950 142.350 102.300 ;
        RECT 143.550 101.400 145.350 107.250 ;
        RECT 155.550 102.300 157.350 107.250 ;
        RECT 158.550 103.200 160.350 107.250 ;
        RECT 161.550 102.300 163.350 107.250 ;
        RECT 143.550 99.300 144.750 101.400 ;
        RECT 155.550 100.950 163.350 102.300 ;
        RECT 164.550 101.400 166.350 107.250 ;
        RECT 175.650 101.400 177.450 107.250 ;
        RECT 178.650 101.400 180.450 107.250 ;
        RECT 190.650 101.400 192.450 107.250 ;
        RECT 164.550 99.300 165.750 101.400 ;
        RECT 141.000 98.250 144.750 99.300 ;
        RECT 162.000 98.250 165.750 99.300 ;
        RECT 106.950 92.850 109.050 94.950 ;
        RECT 124.950 94.050 127.050 96.150 ;
        RECT 127.950 95.850 130.050 97.950 ;
        RECT 137.100 96.150 138.900 97.950 ;
        RECT 128.100 94.050 129.900 95.850 ;
        RECT 89.100 91.050 90.900 92.850 ;
        RECT 101.100 91.050 102.900 92.850 ;
        RECT 87.000 87.600 89.550 88.650 ;
        RECT 106.950 87.600 108.150 92.850 ;
        RECT 109.950 89.850 112.050 91.950 ;
        RECT 109.950 88.050 111.750 89.850 ;
        RECT 62.100 85.050 63.900 86.850 ;
        RECT 56.250 81.900 63.300 82.800 ;
        RECT 56.250 81.600 57.450 81.900 ;
        RECT 10.650 75.750 12.450 81.600 ;
        RECT 13.650 75.750 15.450 81.600 ;
        RECT 16.650 75.750 18.450 81.600 ;
        RECT 22.650 75.750 24.450 81.600 ;
        RECT 25.650 75.750 27.450 81.600 ;
        RECT 28.650 75.750 30.450 81.600 ;
        RECT 38.550 75.750 40.350 81.600 ;
        RECT 41.550 75.750 43.350 81.600 ;
        RECT 44.550 75.750 46.350 81.600 ;
        RECT 55.650 75.750 57.450 81.600 ;
        RECT 61.650 81.600 63.300 81.900 ;
        RECT 58.650 75.750 60.450 81.000 ;
        RECT 61.650 75.750 63.450 81.600 ;
        RECT 64.650 75.750 66.450 81.600 ;
        RECT 69.300 75.750 71.100 87.600 ;
        RECT 73.500 75.750 75.300 87.600 ;
        RECT 76.800 75.750 78.600 81.600 ;
        RECT 83.550 75.750 85.350 87.600 ;
        RECT 87.750 75.750 89.550 87.600 ;
        RECT 102.300 75.750 104.100 87.600 ;
        RECT 106.500 75.750 108.300 87.600 ;
        RECT 125.400 81.600 126.600 94.050 ;
        RECT 133.950 92.850 136.050 94.950 ;
        RECT 136.950 94.050 139.050 96.150 ;
        RECT 140.850 94.950 142.050 98.250 ;
        RECT 158.100 96.150 159.900 97.950 ;
        RECT 139.950 92.850 142.050 94.950 ;
        RECT 154.950 92.850 157.050 94.950 ;
        RECT 157.950 94.050 160.050 96.150 ;
        RECT 161.850 94.950 163.050 98.250 ;
        RECT 176.400 94.950 177.600 101.400 ;
        RECT 191.250 99.300 192.450 101.400 ;
        RECT 193.650 102.300 195.450 107.250 ;
        RECT 196.650 103.200 198.450 107.250 ;
        RECT 199.650 102.300 201.450 107.250 ;
        RECT 193.650 100.950 201.450 102.300 ;
        RECT 210.000 101.400 211.800 107.250 ;
        RECT 214.200 103.050 216.000 107.250 ;
        RECT 217.500 104.400 219.300 107.250 ;
        RECT 214.200 101.400 219.900 103.050 ;
        RECT 191.250 98.250 195.000 99.300 ;
        RECT 179.100 96.150 180.900 97.950 ;
        RECT 190.950 96.450 193.050 97.050 ;
        RECT 160.950 92.850 163.050 94.950 ;
        RECT 175.950 92.850 178.050 94.950 ;
        RECT 178.950 94.050 181.050 96.150 ;
        RECT 188.550 95.550 193.050 96.450 ;
        RECT 134.100 91.050 135.900 92.850 ;
        RECT 139.950 87.600 141.150 92.850 ;
        RECT 142.950 89.850 145.050 91.950 ;
        RECT 155.100 91.050 156.900 92.850 ;
        RECT 142.950 88.050 144.750 89.850 ;
        RECT 160.950 87.600 162.150 92.850 ;
        RECT 163.950 89.850 166.050 91.950 ;
        RECT 163.950 88.050 165.750 89.850 ;
        RECT 176.400 87.600 177.600 92.850 ;
        RECT 109.800 75.750 111.600 81.600 ;
        RECT 124.650 75.750 126.450 81.600 ;
        RECT 127.650 75.750 129.450 81.600 ;
        RECT 135.300 75.750 137.100 87.600 ;
        RECT 139.500 75.750 141.300 87.600 ;
        RECT 142.800 75.750 144.600 81.600 ;
        RECT 156.300 75.750 158.100 87.600 ;
        RECT 160.500 75.750 162.300 87.600 ;
        RECT 163.800 75.750 165.600 81.600 ;
        RECT 175.650 75.750 177.450 87.600 ;
        RECT 178.650 75.750 180.450 87.600 ;
        RECT 188.550 84.450 189.450 95.550 ;
        RECT 190.950 94.950 193.050 95.550 ;
        RECT 193.950 94.950 195.150 98.250 ;
        RECT 197.100 96.150 198.900 97.950 ;
        RECT 209.100 96.150 210.900 97.950 ;
        RECT 193.950 92.850 196.050 94.950 ;
        RECT 196.950 94.050 199.050 96.150 ;
        RECT 199.950 92.850 202.050 94.950 ;
        RECT 208.950 94.050 211.050 96.150 ;
        RECT 211.950 95.850 214.050 97.950 ;
        RECT 215.100 96.150 216.900 97.950 ;
        RECT 212.100 94.050 213.900 95.850 ;
        RECT 214.950 94.050 217.050 96.150 ;
        RECT 218.700 94.950 219.900 101.400 ;
        RECT 233.850 100.200 235.650 107.250 ;
        RECT 238.350 101.400 240.150 107.250 ;
        RECT 233.850 99.300 237.450 100.200 ;
        RECT 217.950 92.850 220.050 94.950 ;
        RECT 233.100 93.150 234.900 94.950 ;
        RECT 190.950 89.850 193.050 91.950 ;
        RECT 191.250 88.050 193.050 89.850 ;
        RECT 194.850 87.600 196.050 92.850 ;
        RECT 200.100 91.050 201.900 92.850 ;
        RECT 218.700 87.600 219.900 92.850 ;
        RECT 232.950 91.050 235.050 93.150 ;
        RECT 236.250 91.950 237.450 99.300 ;
        RECT 248.100 99.000 249.900 107.250 ;
        RECT 245.400 97.350 249.900 99.000 ;
        RECT 253.500 98.400 255.300 107.250 ;
        RECT 260.850 101.400 262.650 107.250 ;
        RECT 265.350 100.200 267.150 107.250 ;
        RECT 263.550 99.300 267.150 100.200 ;
        RECT 239.100 93.150 240.900 94.950 ;
        RECT 245.400 93.150 246.600 97.350 ;
        RECT 260.100 93.150 261.900 94.950 ;
        RECT 235.950 89.850 238.050 91.950 ;
        RECT 238.950 91.050 241.050 93.150 ;
        RECT 244.950 91.050 247.050 93.150 ;
        RECT 190.950 84.450 193.050 85.050 ;
        RECT 188.550 83.550 193.050 84.450 ;
        RECT 190.950 82.950 193.050 83.550 ;
        RECT 191.400 75.750 193.200 81.600 ;
        RECT 194.700 75.750 196.500 87.600 ;
        RECT 198.900 75.750 200.700 87.600 ;
        RECT 209.550 86.700 217.350 87.600 ;
        RECT 209.550 75.750 211.350 86.700 ;
        RECT 212.550 75.750 214.350 85.800 ;
        RECT 215.550 75.750 217.350 86.700 ;
        RECT 218.550 75.750 220.350 87.600 ;
        RECT 236.250 81.600 237.450 89.850 ;
        RECT 245.250 82.800 246.300 91.050 ;
        RECT 247.950 89.850 250.050 91.950 ;
        RECT 253.950 89.850 256.050 91.950 ;
        RECT 259.950 91.050 262.050 93.150 ;
        RECT 263.550 91.950 264.750 99.300 ;
        RECT 272.700 98.400 274.500 107.250 ;
        RECT 278.100 99.000 279.900 107.250 ;
        RECT 290.550 102.300 292.350 107.250 ;
        RECT 293.550 103.200 295.350 107.250 ;
        RECT 296.550 102.300 298.350 107.250 ;
        RECT 290.550 100.950 298.350 102.300 ;
        RECT 299.550 101.400 301.350 107.250 ;
        RECT 308.550 102.300 310.350 107.250 ;
        RECT 311.550 103.200 313.350 107.250 ;
        RECT 314.550 102.300 316.350 107.250 ;
        RECT 299.550 99.300 300.750 101.400 ;
        RECT 308.550 100.950 316.350 102.300 ;
        RECT 317.550 101.400 319.350 107.250 ;
        RECT 325.650 104.400 327.450 107.250 ;
        RECT 328.650 104.400 330.450 107.250 ;
        RECT 331.650 104.400 333.450 107.250 ;
        RECT 317.550 99.300 318.750 101.400 ;
        RECT 278.100 97.350 282.600 99.000 ;
        RECT 297.000 98.250 300.750 99.300 ;
        RECT 315.000 98.250 318.750 99.300 ;
        RECT 266.100 93.150 267.900 94.950 ;
        RECT 281.400 93.150 282.600 97.350 ;
        RECT 293.100 96.150 294.900 97.950 ;
        RECT 262.950 89.850 265.050 91.950 ;
        RECT 265.950 91.050 268.050 93.150 ;
        RECT 271.950 89.850 274.050 91.950 ;
        RECT 277.950 89.850 280.050 91.950 ;
        RECT 280.950 91.050 283.050 93.150 ;
        RECT 289.950 92.850 292.050 94.950 ;
        RECT 292.950 94.050 295.050 96.150 ;
        RECT 296.850 94.950 298.050 98.250 ;
        RECT 311.100 96.150 312.900 97.950 ;
        RECT 295.950 92.850 298.050 94.950 ;
        RECT 307.950 92.850 310.050 94.950 ;
        RECT 310.950 94.050 313.050 96.150 ;
        RECT 314.850 94.950 316.050 98.250 ;
        RECT 328.950 97.950 330.000 104.400 ;
        RECT 335.550 99.900 337.350 107.250 ;
        RECT 340.050 101.400 341.850 107.250 ;
        RECT 343.050 102.900 344.850 107.250 ;
        RECT 343.050 101.400 346.350 102.900 ;
        RECT 351.000 101.400 352.800 107.250 ;
        RECT 355.200 103.050 357.000 107.250 ;
        RECT 358.500 104.400 360.300 107.250 ;
        RECT 355.200 101.400 360.900 103.050 ;
        RECT 341.250 99.900 343.050 100.500 ;
        RECT 335.550 98.700 343.050 99.900 ;
        RECT 328.950 95.850 331.050 97.950 ;
        RECT 313.950 92.850 316.050 94.950 ;
        RECT 325.950 92.850 328.050 94.950 ;
        RECT 290.100 91.050 291.900 92.850 ;
        RECT 247.950 88.050 249.750 89.850 ;
        RECT 250.950 86.850 253.050 88.950 ;
        RECT 254.100 88.050 255.900 89.850 ;
        RECT 251.100 85.050 252.900 86.850 ;
        RECT 245.250 81.900 252.300 82.800 ;
        RECT 245.250 81.600 246.450 81.900 ;
        RECT 232.650 75.750 234.450 81.600 ;
        RECT 235.650 75.750 237.450 81.600 ;
        RECT 238.650 75.750 240.450 81.600 ;
        RECT 244.650 75.750 246.450 81.600 ;
        RECT 250.650 81.600 252.300 81.900 ;
        RECT 263.550 81.600 264.750 89.850 ;
        RECT 272.100 88.050 273.900 89.850 ;
        RECT 274.950 86.850 277.050 88.950 ;
        RECT 278.250 88.050 280.050 89.850 ;
        RECT 275.100 85.050 276.900 86.850 ;
        RECT 281.700 82.800 282.750 91.050 ;
        RECT 295.950 87.600 297.150 92.850 ;
        RECT 298.950 89.850 301.050 91.950 ;
        RECT 308.100 91.050 309.900 92.850 ;
        RECT 298.950 88.050 300.750 89.850 ;
        RECT 313.950 87.600 315.150 92.850 ;
        RECT 316.950 89.850 319.050 91.950 ;
        RECT 326.100 91.050 327.900 92.850 ;
        RECT 316.950 88.050 318.750 89.850 ;
        RECT 328.950 88.650 330.000 95.850 ;
        RECT 331.950 92.850 334.050 94.950 ;
        RECT 334.950 92.850 337.050 94.950 ;
        RECT 332.100 91.050 333.900 92.850 ;
        RECT 335.100 91.050 336.900 92.850 ;
        RECT 327.450 87.600 330.000 88.650 ;
        RECT 275.700 81.900 282.750 82.800 ;
        RECT 275.700 81.600 277.350 81.900 ;
        RECT 247.650 75.750 249.450 81.000 ;
        RECT 250.650 75.750 252.450 81.600 ;
        RECT 253.650 75.750 255.450 81.600 ;
        RECT 260.550 75.750 262.350 81.600 ;
        RECT 263.550 75.750 265.350 81.600 ;
        RECT 266.550 75.750 268.350 81.600 ;
        RECT 272.550 75.750 274.350 81.600 ;
        RECT 275.550 75.750 277.350 81.600 ;
        RECT 281.550 81.600 282.750 81.900 ;
        RECT 278.550 75.750 280.350 81.000 ;
        RECT 281.550 75.750 283.350 81.600 ;
        RECT 291.300 75.750 293.100 87.600 ;
        RECT 295.500 75.750 297.300 87.600 ;
        RECT 298.800 75.750 300.600 81.600 ;
        RECT 309.300 75.750 311.100 87.600 ;
        RECT 313.500 75.750 315.300 87.600 ;
        RECT 316.800 75.750 318.600 81.600 ;
        RECT 327.450 75.750 329.250 87.600 ;
        RECT 331.650 75.750 333.450 87.600 ;
        RECT 338.700 81.600 339.900 98.700 ;
        RECT 345.150 94.950 346.350 101.400 ;
        RECT 350.100 96.150 351.900 97.950 ;
        RECT 341.100 93.150 342.900 94.950 ;
        RECT 340.950 91.050 343.050 93.150 ;
        RECT 343.950 92.850 346.350 94.950 ;
        RECT 349.950 94.050 352.050 96.150 ;
        RECT 352.950 95.850 355.050 97.950 ;
        RECT 356.100 96.150 357.900 97.950 ;
        RECT 353.100 94.050 354.900 95.850 ;
        RECT 355.950 94.050 358.050 96.150 ;
        RECT 359.700 94.950 360.900 101.400 ;
        RECT 374.850 100.200 376.650 107.250 ;
        RECT 379.350 101.400 381.150 107.250 ;
        RECT 390.000 101.400 391.800 107.250 ;
        RECT 394.200 101.400 396.000 107.250 ;
        RECT 398.400 101.400 400.200 107.250 ;
        RECT 407.550 102.300 409.350 107.250 ;
        RECT 410.550 103.200 412.350 107.250 ;
        RECT 413.550 102.300 415.350 107.250 ;
        RECT 374.850 99.300 378.450 100.200 ;
        RECT 358.950 92.850 361.050 94.950 ;
        RECT 374.100 93.150 375.900 94.950 ;
        RECT 345.150 87.600 346.350 92.850 ;
        RECT 359.700 87.600 360.900 92.850 ;
        RECT 373.950 91.050 376.050 93.150 ;
        RECT 377.250 91.950 378.450 99.300 ;
        RECT 392.250 96.150 394.050 97.950 ;
        RECT 380.100 93.150 381.900 94.950 ;
        RECT 376.950 89.850 379.050 91.950 ;
        RECT 379.950 91.050 382.050 93.150 ;
        RECT 388.950 92.850 391.050 94.950 ;
        RECT 391.950 94.050 394.050 96.150 ;
        RECT 394.950 94.950 396.000 101.400 ;
        RECT 407.550 100.950 415.350 102.300 ;
        RECT 416.550 101.400 418.350 107.250 ;
        RECT 416.550 99.300 417.750 101.400 ;
        RECT 414.000 98.250 417.750 99.300 ;
        RECT 428.700 98.400 430.500 107.250 ;
        RECT 434.100 99.000 435.900 107.250 ;
        RECT 449.550 102.300 451.350 107.250 ;
        RECT 452.550 103.200 454.350 107.250 ;
        RECT 455.550 102.300 457.350 107.250 ;
        RECT 449.550 100.950 457.350 102.300 ;
        RECT 458.550 101.400 460.350 107.250 ;
        RECT 467.550 102.300 469.350 107.250 ;
        RECT 470.550 103.200 472.350 107.250 ;
        RECT 473.550 102.300 475.350 107.250 ;
        RECT 458.550 99.300 459.750 101.400 ;
        RECT 467.550 100.950 475.350 102.300 ;
        RECT 476.550 101.400 478.350 107.250 ;
        RECT 485.550 102.300 487.350 107.250 ;
        RECT 488.550 103.200 490.350 107.250 ;
        RECT 491.550 102.300 493.350 107.250 ;
        RECT 476.550 99.300 477.750 101.400 ;
        RECT 485.550 100.950 493.350 102.300 ;
        RECT 494.550 101.400 496.350 107.250 ;
        RECT 506.700 104.400 508.500 107.250 ;
        RECT 510.000 103.050 511.800 107.250 ;
        RECT 506.100 101.400 511.800 103.050 ;
        RECT 514.200 101.400 516.000 107.250 ;
        RECT 494.550 99.300 495.750 101.400 ;
        RECT 397.950 96.150 399.750 97.950 ;
        RECT 410.100 96.150 411.900 97.950 ;
        RECT 394.950 92.850 397.050 94.950 ;
        RECT 397.950 94.050 400.050 96.150 ;
        RECT 400.950 92.850 403.050 94.950 ;
        RECT 406.950 92.850 409.050 94.950 ;
        RECT 409.950 94.050 412.050 96.150 ;
        RECT 413.850 94.950 415.050 98.250 ;
        RECT 434.100 97.350 438.600 99.000 ;
        RECT 456.000 98.250 459.750 99.300 ;
        RECT 474.000 98.250 477.750 99.300 ;
        RECT 492.000 98.250 495.750 99.300 ;
        RECT 412.950 92.850 415.050 94.950 ;
        RECT 437.400 93.150 438.600 97.350 ;
        RECT 452.100 96.150 453.900 97.950 ;
        RECT 389.250 91.050 391.050 92.850 ;
        RECT 335.550 75.750 337.350 81.600 ;
        RECT 338.550 75.750 340.350 81.600 ;
        RECT 342.150 75.750 343.950 87.600 ;
        RECT 345.150 75.750 346.950 87.600 ;
        RECT 350.550 86.700 358.350 87.600 ;
        RECT 350.550 75.750 352.350 86.700 ;
        RECT 353.550 75.750 355.350 85.800 ;
        RECT 356.550 75.750 358.350 86.700 ;
        RECT 359.550 75.750 361.350 87.600 ;
        RECT 377.250 81.600 378.450 89.850 ;
        RECT 396.150 89.400 397.050 92.850 ;
        RECT 401.100 91.050 402.900 92.850 ;
        RECT 407.100 91.050 408.900 92.850 ;
        RECT 396.150 88.500 400.200 89.400 ;
        RECT 398.400 87.600 400.200 88.500 ;
        RECT 412.950 87.600 414.150 92.850 ;
        RECT 415.950 89.850 418.050 91.950 ;
        RECT 427.950 89.850 430.050 91.950 ;
        RECT 433.950 89.850 436.050 91.950 ;
        RECT 436.950 91.050 439.050 93.150 ;
        RECT 448.950 92.850 451.050 94.950 ;
        RECT 451.950 94.050 454.050 96.150 ;
        RECT 455.850 94.950 457.050 98.250 ;
        RECT 470.100 96.150 471.900 97.950 ;
        RECT 454.950 92.850 457.050 94.950 ;
        RECT 466.950 92.850 469.050 94.950 ;
        RECT 469.950 94.050 472.050 96.150 ;
        RECT 473.850 94.950 475.050 98.250 ;
        RECT 488.100 96.150 489.900 97.950 ;
        RECT 472.950 92.850 475.050 94.950 ;
        RECT 484.950 92.850 487.050 94.950 ;
        RECT 487.950 94.050 490.050 96.150 ;
        RECT 491.850 94.950 493.050 98.250 ;
        RECT 506.100 94.950 507.300 101.400 ;
        RECT 524.700 98.400 526.500 107.250 ;
        RECT 530.100 99.000 531.900 107.250 ;
        RECT 542.850 100.200 544.650 107.250 ;
        RECT 547.350 101.400 549.150 107.250 ;
        RECT 542.850 99.300 546.450 100.200 ;
        RECT 509.100 96.150 510.900 97.950 ;
        RECT 490.950 92.850 493.050 94.950 ;
        RECT 505.950 92.850 508.050 94.950 ;
        RECT 508.950 94.050 511.050 96.150 ;
        RECT 511.950 95.850 514.050 97.950 ;
        RECT 515.100 96.150 516.900 97.950 ;
        RECT 530.100 97.350 534.600 99.000 ;
        RECT 526.950 96.450 529.050 97.050 ;
        RECT 512.100 94.050 513.900 95.850 ;
        RECT 514.950 94.050 517.050 96.150 ;
        RECT 518.550 95.550 529.050 96.450 ;
        RECT 449.100 91.050 450.900 92.850 ;
        RECT 415.950 88.050 417.750 89.850 ;
        RECT 428.100 88.050 429.900 89.850 ;
        RECT 389.550 86.400 397.350 87.300 ;
        RECT 373.650 75.750 375.450 81.600 ;
        RECT 376.650 75.750 378.450 81.600 ;
        RECT 379.650 75.750 381.450 81.600 ;
        RECT 389.550 75.750 391.350 86.400 ;
        RECT 392.550 75.750 394.350 85.500 ;
        RECT 395.550 76.500 397.350 86.400 ;
        RECT 398.550 77.400 400.350 87.600 ;
        RECT 401.550 76.500 403.350 87.600 ;
        RECT 395.550 75.750 403.350 76.500 ;
        RECT 408.300 75.750 410.100 87.600 ;
        RECT 412.500 75.750 414.300 87.600 ;
        RECT 430.950 86.850 433.050 88.950 ;
        RECT 434.250 88.050 436.050 89.850 ;
        RECT 431.100 85.050 432.900 86.850 ;
        RECT 437.700 82.800 438.750 91.050 ;
        RECT 454.950 87.600 456.150 92.850 ;
        RECT 457.950 89.850 460.050 91.950 ;
        RECT 467.100 91.050 468.900 92.850 ;
        RECT 457.950 88.050 459.750 89.850 ;
        RECT 472.950 87.600 474.150 92.850 ;
        RECT 475.950 89.850 478.050 91.950 ;
        RECT 485.100 91.050 486.900 92.850 ;
        RECT 475.950 88.050 477.750 89.850 ;
        RECT 490.950 87.600 492.150 92.850 ;
        RECT 493.950 89.850 496.050 91.950 ;
        RECT 493.950 88.050 495.750 89.850 ;
        RECT 506.100 87.600 507.300 92.850 ;
        RECT 514.950 90.450 517.050 91.050 ;
        RECT 518.550 90.450 519.450 95.550 ;
        RECT 526.950 94.950 529.050 95.550 ;
        RECT 533.400 93.150 534.600 97.350 ;
        RECT 542.100 93.150 543.900 94.950 ;
        RECT 514.950 89.550 519.450 90.450 ;
        RECT 523.950 89.850 526.050 91.950 ;
        RECT 529.950 89.850 532.050 91.950 ;
        RECT 532.950 91.050 535.050 93.150 ;
        RECT 541.950 91.050 544.050 93.150 ;
        RECT 545.250 91.950 546.450 99.300 ;
        RECT 554.550 99.900 556.350 107.250 ;
        RECT 559.050 101.400 560.850 107.250 ;
        RECT 562.050 102.900 563.850 107.250 ;
        RECT 562.050 101.400 565.350 102.900 ;
        RECT 560.250 99.900 562.050 100.500 ;
        RECT 554.550 98.700 562.050 99.900 ;
        RECT 548.100 93.150 549.900 94.950 ;
        RECT 514.950 88.950 517.050 89.550 ;
        RECT 524.100 88.050 525.900 89.850 ;
        RECT 431.700 81.900 438.750 82.800 ;
        RECT 431.700 81.600 433.350 81.900 ;
        RECT 415.800 75.750 417.600 81.600 ;
        RECT 428.550 75.750 430.350 81.600 ;
        RECT 431.550 75.750 433.350 81.600 ;
        RECT 437.550 81.600 438.750 81.900 ;
        RECT 434.550 75.750 436.350 81.000 ;
        RECT 437.550 75.750 439.350 81.600 ;
        RECT 450.300 75.750 452.100 87.600 ;
        RECT 454.500 75.750 456.300 87.600 ;
        RECT 457.800 75.750 459.600 81.600 ;
        RECT 468.300 75.750 470.100 87.600 ;
        RECT 472.500 75.750 474.300 87.600 ;
        RECT 475.800 75.750 477.600 81.600 ;
        RECT 486.300 75.750 488.100 87.600 ;
        RECT 490.500 75.750 492.300 87.600 ;
        RECT 493.800 75.750 495.600 81.600 ;
        RECT 505.650 75.750 507.450 87.600 ;
        RECT 508.650 86.700 516.450 87.600 ;
        RECT 526.950 86.850 529.050 88.950 ;
        RECT 530.250 88.050 532.050 89.850 ;
        RECT 508.650 75.750 510.450 86.700 ;
        RECT 511.650 75.750 513.450 85.800 ;
        RECT 514.650 75.750 516.450 86.700 ;
        RECT 527.100 85.050 528.900 86.850 ;
        RECT 533.700 82.800 534.750 91.050 ;
        RECT 544.950 89.850 547.050 91.950 ;
        RECT 547.950 91.050 550.050 93.150 ;
        RECT 553.950 92.850 556.050 94.950 ;
        RECT 554.100 91.050 555.900 92.850 ;
        RECT 527.700 81.900 534.750 82.800 ;
        RECT 527.700 81.600 529.350 81.900 ;
        RECT 524.550 75.750 526.350 81.600 ;
        RECT 527.550 75.750 529.350 81.600 ;
        RECT 533.550 81.600 534.750 81.900 ;
        RECT 545.250 81.600 546.450 89.850 ;
        RECT 557.700 81.600 558.900 98.700 ;
        RECT 564.150 94.950 565.350 101.400 ;
        RECT 575.700 98.400 577.500 107.250 ;
        RECT 581.100 99.000 582.900 107.250 ;
        RECT 593.700 104.400 595.500 107.250 ;
        RECT 597.000 103.050 598.800 107.250 ;
        RECT 593.100 101.400 598.800 103.050 ;
        RECT 601.200 101.400 603.000 107.250 ;
        RECT 608.850 101.400 610.650 107.250 ;
        RECT 581.100 97.350 585.600 99.000 ;
        RECT 560.100 93.150 561.900 94.950 ;
        RECT 559.950 91.050 562.050 93.150 ;
        RECT 562.950 92.850 565.350 94.950 ;
        RECT 584.400 93.150 585.600 97.350 ;
        RECT 593.100 94.950 594.300 101.400 ;
        RECT 613.350 100.200 615.150 107.250 ;
        RECT 611.550 99.300 615.150 100.200 ;
        RECT 596.100 96.150 597.900 97.950 ;
        RECT 564.150 87.600 565.350 92.850 ;
        RECT 574.950 89.850 577.050 91.950 ;
        RECT 580.950 89.850 583.050 91.950 ;
        RECT 583.950 91.050 586.050 93.150 ;
        RECT 592.950 92.850 595.050 94.950 ;
        RECT 595.950 94.050 598.050 96.150 ;
        RECT 598.950 95.850 601.050 97.950 ;
        RECT 602.100 96.150 603.900 97.950 ;
        RECT 599.100 94.050 600.900 95.850 ;
        RECT 601.950 94.050 604.050 96.150 ;
        RECT 608.100 93.150 609.900 94.950 ;
        RECT 575.100 88.050 576.900 89.850 ;
        RECT 530.550 75.750 532.350 81.000 ;
        RECT 533.550 75.750 535.350 81.600 ;
        RECT 541.650 75.750 543.450 81.600 ;
        RECT 544.650 75.750 546.450 81.600 ;
        RECT 547.650 75.750 549.450 81.600 ;
        RECT 554.550 75.750 556.350 81.600 ;
        RECT 557.550 75.750 559.350 81.600 ;
        RECT 561.150 75.750 562.950 87.600 ;
        RECT 564.150 75.750 565.950 87.600 ;
        RECT 577.950 86.850 580.050 88.950 ;
        RECT 581.250 88.050 583.050 89.850 ;
        RECT 578.100 85.050 579.900 86.850 ;
        RECT 584.700 82.800 585.750 91.050 ;
        RECT 593.100 87.600 594.300 92.850 ;
        RECT 607.950 91.050 610.050 93.150 ;
        RECT 611.550 91.950 612.750 99.300 ;
        RECT 623.700 98.400 625.500 107.250 ;
        RECT 629.100 99.000 630.900 107.250 ;
        RECT 642.000 101.400 643.800 107.250 ;
        RECT 646.200 103.050 648.000 107.250 ;
        RECT 649.500 104.400 651.300 107.250 ;
        RECT 646.200 101.400 651.900 103.050 ;
        RECT 661.650 101.400 663.450 107.250 ;
        RECT 629.100 97.350 633.600 99.000 ;
        RECT 614.100 93.150 615.900 94.950 ;
        RECT 632.400 93.150 633.600 97.350 ;
        RECT 641.100 96.150 642.900 97.950 ;
        RECT 640.950 94.050 643.050 96.150 ;
        RECT 643.950 95.850 646.050 97.950 ;
        RECT 647.100 96.150 648.900 97.950 ;
        RECT 644.100 94.050 645.900 95.850 ;
        RECT 646.950 94.050 649.050 96.150 ;
        RECT 650.700 94.950 651.900 101.400 ;
        RECT 662.250 99.300 663.450 101.400 ;
        RECT 664.650 102.300 666.450 107.250 ;
        RECT 667.650 103.200 669.450 107.250 ;
        RECT 670.650 102.300 672.450 107.250 ;
        RECT 664.650 100.950 672.450 102.300 ;
        RECT 677.550 99.900 679.350 107.250 ;
        RECT 682.050 101.400 683.850 107.250 ;
        RECT 685.050 102.900 686.850 107.250 ;
        RECT 692.550 104.400 694.350 107.250 ;
        RECT 695.550 104.400 697.350 107.250 ;
        RECT 698.550 104.400 700.350 107.250 ;
        RECT 710.250 104.400 712.350 107.250 ;
        RECT 713.550 104.400 715.350 107.250 ;
        RECT 716.550 104.400 718.350 107.250 ;
        RECT 719.550 104.400 721.350 107.250 ;
        RECT 685.050 101.400 688.350 102.900 ;
        RECT 683.250 99.900 685.050 100.500 ;
        RECT 662.250 98.250 666.000 99.300 ;
        RECT 677.550 98.700 685.050 99.900 ;
        RECT 664.950 94.950 666.150 98.250 ;
        RECT 668.100 96.150 669.900 97.950 ;
        RECT 610.950 89.850 613.050 91.950 ;
        RECT 613.950 91.050 616.050 93.150 ;
        RECT 622.950 89.850 625.050 91.950 ;
        RECT 628.950 89.850 631.050 91.950 ;
        RECT 631.950 91.050 634.050 93.150 ;
        RECT 649.950 92.850 652.050 94.950 ;
        RECT 664.950 92.850 667.050 94.950 ;
        RECT 667.950 94.050 670.050 96.150 ;
        RECT 670.950 92.850 673.050 94.950 ;
        RECT 676.950 92.850 679.050 94.950 ;
        RECT 578.700 81.900 585.750 82.800 ;
        RECT 578.700 81.600 580.350 81.900 ;
        RECT 575.550 75.750 577.350 81.600 ;
        RECT 578.550 75.750 580.350 81.600 ;
        RECT 584.550 81.600 585.750 81.900 ;
        RECT 581.550 75.750 583.350 81.000 ;
        RECT 584.550 75.750 586.350 81.600 ;
        RECT 592.650 75.750 594.450 87.600 ;
        RECT 595.650 86.700 603.450 87.600 ;
        RECT 595.650 75.750 597.450 86.700 ;
        RECT 598.650 75.750 600.450 85.800 ;
        RECT 601.650 75.750 603.450 86.700 ;
        RECT 611.550 81.600 612.750 89.850 ;
        RECT 623.100 88.050 624.900 89.850 ;
        RECT 625.950 86.850 628.050 88.950 ;
        RECT 629.250 88.050 631.050 89.850 ;
        RECT 626.100 85.050 627.900 86.850 ;
        RECT 632.700 82.800 633.750 91.050 ;
        RECT 650.700 87.600 651.900 92.850 ;
        RECT 661.950 89.850 664.050 91.950 ;
        RECT 662.250 88.050 664.050 89.850 ;
        RECT 665.850 87.600 667.050 92.850 ;
        RECT 671.100 91.050 672.900 92.850 ;
        RECT 677.100 91.050 678.900 92.850 ;
        RECT 626.700 81.900 633.750 82.800 ;
        RECT 626.700 81.600 628.350 81.900 ;
        RECT 608.550 75.750 610.350 81.600 ;
        RECT 611.550 75.750 613.350 81.600 ;
        RECT 614.550 75.750 616.350 81.600 ;
        RECT 623.550 75.750 625.350 81.600 ;
        RECT 626.550 75.750 628.350 81.600 ;
        RECT 632.550 81.600 633.750 81.900 ;
        RECT 641.550 86.700 649.350 87.600 ;
        RECT 629.550 75.750 631.350 81.000 ;
        RECT 632.550 75.750 634.350 81.600 ;
        RECT 641.550 75.750 643.350 86.700 ;
        RECT 644.550 75.750 646.350 85.800 ;
        RECT 647.550 75.750 649.350 86.700 ;
        RECT 650.550 75.750 652.350 87.600 ;
        RECT 662.400 75.750 664.200 81.600 ;
        RECT 665.700 75.750 667.500 87.600 ;
        RECT 669.900 75.750 671.700 87.600 ;
        RECT 680.700 81.600 681.900 98.700 ;
        RECT 687.150 94.950 688.350 101.400 ;
        RECT 696.000 97.950 697.050 104.400 ;
        RECT 714.300 103.500 715.350 104.400 ;
        RECT 720.300 103.500 721.350 104.400 ;
        RECT 714.300 102.600 725.100 103.500 ;
        RECT 694.950 95.850 697.050 97.950 ;
        RECT 716.100 96.150 717.900 97.950 ;
        RECT 723.900 96.150 725.100 102.600 ;
        RECT 737.850 100.200 739.650 107.250 ;
        RECT 742.350 101.400 744.150 107.250 ;
        RECT 751.650 104.400 753.450 107.250 ;
        RECT 754.650 104.400 756.450 107.250 ;
        RECT 737.850 99.300 741.450 100.200 ;
        RECT 683.100 93.150 684.900 94.950 ;
        RECT 682.950 91.050 685.050 93.150 ;
        RECT 685.950 92.850 688.350 94.950 ;
        RECT 691.950 92.850 694.050 94.950 ;
        RECT 687.150 87.600 688.350 92.850 ;
        RECT 692.100 91.050 693.900 92.850 ;
        RECT 696.000 88.650 697.050 95.850 ;
        RECT 697.950 92.850 700.050 94.950 ;
        RECT 709.950 92.850 712.050 94.950 ;
        RECT 715.950 94.050 718.050 96.150 ;
        RECT 718.950 92.850 721.050 94.950 ;
        RECT 723.900 94.050 727.050 96.150 ;
        RECT 698.100 91.050 699.900 92.850 ;
        RECT 710.100 91.050 711.900 92.850 ;
        RECT 719.100 91.050 720.900 92.850 ;
        RECT 723.900 88.800 725.100 94.050 ;
        RECT 737.100 93.150 738.900 94.950 ;
        RECT 736.950 91.050 739.050 93.150 ;
        RECT 740.250 91.950 741.450 99.300 ;
        RECT 752.400 96.150 753.600 104.400 ;
        RECT 761.550 102.300 763.350 107.250 ;
        RECT 764.550 103.200 766.350 107.250 ;
        RECT 767.550 102.300 769.350 107.250 ;
        RECT 761.550 100.950 769.350 102.300 ;
        RECT 770.550 101.400 772.350 107.250 ;
        RECT 776.550 102.300 778.350 107.250 ;
        RECT 779.550 103.200 781.350 107.250 ;
        RECT 782.550 102.300 784.350 107.250 ;
        RECT 760.950 99.450 763.050 100.050 ;
        RECT 758.550 98.550 763.050 99.450 ;
        RECT 770.550 99.300 771.750 101.400 ;
        RECT 776.550 100.950 784.350 102.300 ;
        RECT 785.550 101.400 787.350 107.250 ;
        RECT 796.650 101.400 798.450 107.250 ;
        RECT 785.550 99.300 786.750 101.400 ;
        RECT 743.100 93.150 744.900 94.950 ;
        RECT 751.950 94.050 754.050 96.150 ;
        RECT 754.950 95.850 757.050 97.950 ;
        RECT 755.100 94.050 756.900 95.850 ;
        RECT 739.950 89.850 742.050 91.950 ;
        RECT 742.950 91.050 745.050 93.150 ;
        RECT 696.000 87.600 698.550 88.650 ;
        RECT 723.900 87.600 727.350 88.800 ;
        RECT 677.550 75.750 679.350 81.600 ;
        RECT 680.550 75.750 682.350 81.600 ;
        RECT 684.150 75.750 685.950 87.600 ;
        RECT 687.150 75.750 688.950 87.600 ;
        RECT 692.550 75.750 694.350 87.600 ;
        RECT 696.750 75.750 698.550 87.600 ;
        RECT 707.550 85.500 715.350 86.400 ;
        RECT 707.550 75.750 709.350 85.500 ;
        RECT 710.550 75.750 712.350 84.600 ;
        RECT 713.550 76.500 715.350 85.500 ;
        RECT 716.550 85.200 724.950 86.100 ;
        RECT 716.550 77.400 718.350 85.200 ;
        RECT 719.550 76.500 721.350 84.300 ;
        RECT 713.550 75.750 721.350 76.500 ;
        RECT 723.150 76.500 724.950 85.200 ;
        RECT 726.150 85.200 727.350 87.600 ;
        RECT 726.150 77.400 727.950 85.200 ;
        RECT 729.150 76.500 730.950 85.800 ;
        RECT 740.250 81.600 741.450 89.850 ;
        RECT 752.400 81.600 753.600 94.050 ;
        RECT 758.550 91.050 759.450 98.550 ;
        RECT 760.950 97.950 763.050 98.550 ;
        RECT 768.000 98.250 771.750 99.300 ;
        RECT 783.000 98.250 786.750 99.300 ;
        RECT 797.250 99.300 798.450 101.400 ;
        RECT 799.650 102.300 801.450 107.250 ;
        RECT 802.650 103.200 804.450 107.250 ;
        RECT 805.650 102.300 807.450 107.250 ;
        RECT 812.550 104.400 814.350 107.250 ;
        RECT 815.550 104.400 817.350 107.250 ;
        RECT 818.550 104.400 820.350 107.250 ;
        RECT 799.650 100.950 807.450 102.300 ;
        RECT 797.250 98.250 801.000 99.300 ;
        RECT 764.100 96.150 765.900 97.950 ;
        RECT 760.950 92.850 763.050 94.950 ;
        RECT 763.950 94.050 766.050 96.150 ;
        RECT 767.850 94.950 769.050 98.250 ;
        RECT 779.100 96.150 780.900 97.950 ;
        RECT 766.950 92.850 769.050 94.950 ;
        RECT 775.950 92.850 778.050 94.950 ;
        RECT 778.950 94.050 781.050 96.150 ;
        RECT 782.850 94.950 784.050 98.250 ;
        RECT 784.950 96.450 787.050 97.050 ;
        RECT 793.950 96.450 796.050 97.050 ;
        RECT 784.950 95.550 796.050 96.450 ;
        RECT 784.950 94.950 787.050 95.550 ;
        RECT 793.950 94.950 796.050 95.550 ;
        RECT 799.950 94.950 801.150 98.250 ;
        RECT 816.000 97.950 817.050 104.400 ;
        RECT 827.550 99.900 829.350 107.250 ;
        RECT 832.050 101.400 833.850 107.250 ;
        RECT 835.050 102.900 836.850 107.250 ;
        RECT 845.550 104.400 847.350 107.250 ;
        RECT 848.550 104.400 850.350 107.250 ;
        RECT 851.550 104.400 853.350 107.250 ;
        RECT 835.050 101.400 838.350 102.900 ;
        RECT 833.250 99.900 835.050 100.500 ;
        RECT 827.550 98.700 835.050 99.900 ;
        RECT 803.100 96.150 804.900 97.950 ;
        RECT 781.950 92.850 784.050 94.950 ;
        RECT 799.950 92.850 802.050 94.950 ;
        RECT 802.950 94.050 805.050 96.150 ;
        RECT 814.950 95.850 817.050 97.950 ;
        RECT 805.950 92.850 808.050 94.950 ;
        RECT 811.950 92.850 814.050 94.950 ;
        RECT 761.100 91.050 762.900 92.850 ;
        RECT 757.950 88.950 760.050 91.050 ;
        RECT 766.950 87.600 768.150 92.850 ;
        RECT 769.950 89.850 772.050 91.950 ;
        RECT 776.100 91.050 777.900 92.850 ;
        RECT 769.950 88.050 771.750 89.850 ;
        RECT 781.950 87.600 783.150 92.850 ;
        RECT 784.950 89.850 787.050 91.950 ;
        RECT 796.950 89.850 799.050 91.950 ;
        RECT 784.950 88.050 786.750 89.850 ;
        RECT 797.250 88.050 799.050 89.850 ;
        RECT 800.850 87.600 802.050 92.850 ;
        RECT 806.100 91.050 807.900 92.850 ;
        RECT 812.100 91.050 813.900 92.850 ;
        RECT 816.000 88.650 817.050 95.850 ;
        RECT 817.950 92.850 820.050 94.950 ;
        RECT 826.950 92.850 829.050 94.950 ;
        RECT 818.100 91.050 819.900 92.850 ;
        RECT 827.100 91.050 828.900 92.850 ;
        RECT 816.000 87.600 818.550 88.650 ;
        RECT 723.150 75.750 730.950 76.500 ;
        RECT 736.650 75.750 738.450 81.600 ;
        RECT 739.650 75.750 741.450 81.600 ;
        RECT 742.650 75.750 744.450 81.600 ;
        RECT 751.650 75.750 753.450 81.600 ;
        RECT 754.650 75.750 756.450 81.600 ;
        RECT 762.300 75.750 764.100 87.600 ;
        RECT 766.500 75.750 768.300 87.600 ;
        RECT 769.800 75.750 771.600 81.600 ;
        RECT 777.300 75.750 779.100 87.600 ;
        RECT 781.500 75.750 783.300 87.600 ;
        RECT 784.800 75.750 786.600 81.600 ;
        RECT 797.400 75.750 799.200 81.600 ;
        RECT 800.700 75.750 802.500 87.600 ;
        RECT 804.900 75.750 806.700 87.600 ;
        RECT 812.550 75.750 814.350 87.600 ;
        RECT 816.750 75.750 818.550 87.600 ;
        RECT 830.700 81.600 831.900 98.700 ;
        RECT 837.150 94.950 838.350 101.400 ;
        RECT 849.000 97.950 850.050 104.400 ;
        RECT 847.950 95.850 850.050 97.950 ;
        RECT 833.100 93.150 834.900 94.950 ;
        RECT 832.950 91.050 835.050 93.150 ;
        RECT 835.950 92.850 838.350 94.950 ;
        RECT 844.950 92.850 847.050 94.950 ;
        RECT 837.150 87.600 838.350 92.850 ;
        RECT 845.100 91.050 846.900 92.850 ;
        RECT 849.000 88.650 850.050 95.850 ;
        RECT 850.950 92.850 853.050 94.950 ;
        RECT 851.100 91.050 852.900 92.850 ;
        RECT 849.000 87.600 851.550 88.650 ;
        RECT 827.550 75.750 829.350 81.600 ;
        RECT 830.550 75.750 832.350 81.600 ;
        RECT 834.150 75.750 835.950 87.600 ;
        RECT 837.150 75.750 838.950 87.600 ;
        RECT 845.550 75.750 847.350 87.600 ;
        RECT 849.750 75.750 851.550 87.600 ;
        RECT 2.700 65.400 4.500 71.250 ;
        RECT 5.700 65.400 7.500 71.250 ;
        RECT 8.700 65.400 10.500 71.250 ;
        RECT 5.700 64.500 6.750 65.400 ;
        RECT 2.700 63.600 6.750 64.500 ;
        RECT 2.700 50.100 3.900 63.600 ;
        RECT 11.700 62.700 13.500 71.250 ;
        RECT 14.700 67.950 16.500 71.250 ;
        RECT 17.850 68.400 20.250 71.250 ;
        RECT 21.150 68.400 23.250 71.250 ;
        RECT 24.300 68.400 26.250 71.250 ;
        RECT 17.850 67.050 19.050 68.400 ;
        RECT 21.150 67.050 22.050 68.400 ;
        RECT 24.300 67.050 25.500 68.400 ;
        RECT 16.950 64.950 19.050 67.050 ;
        RECT 19.950 64.950 22.050 67.050 ;
        RECT 22.950 65.400 25.500 67.050 ;
        RECT 27.450 65.400 29.250 71.250 ;
        RECT 31.200 65.400 33.000 71.250 ;
        RECT 34.200 65.400 36.000 71.250 ;
        RECT 22.950 64.950 25.050 65.400 ;
        RECT 31.650 64.500 33.000 65.400 ;
        RECT 37.200 64.500 39.000 71.250 ;
        RECT 40.950 68.400 42.750 71.250 ;
        RECT 31.650 62.850 34.050 64.500 ;
        RECT 7.200 61.650 24.900 62.700 ;
        RECT 31.950 62.400 34.050 62.850 ;
        RECT 36.000 64.200 39.000 64.500 ;
        RECT 36.000 62.400 39.900 64.200 ;
        RECT 7.200 60.900 9.000 61.650 ;
        RECT 19.950 60.150 22.050 60.750 ;
        RECT 10.500 58.950 22.050 60.150 ;
        RECT 22.950 60.600 24.900 61.650 ;
        RECT 41.100 61.350 42.450 68.400 ;
        RECT 43.950 64.950 45.750 71.250 ;
        RECT 46.950 68.400 48.750 71.250 ;
        RECT 47.100 67.200 48.600 68.400 ;
        RECT 47.100 65.100 49.200 67.200 ;
        RECT 50.700 65.400 52.500 71.250 ;
        RECT 43.950 64.050 46.050 64.950 ;
        RECT 53.700 64.500 55.500 71.250 ;
        RECT 56.700 65.400 58.500 71.250 ;
        RECT 59.700 65.400 61.500 71.250 ;
        RECT 62.700 65.400 64.500 71.250 ;
        RECT 66.450 65.400 68.250 71.250 ;
        RECT 69.450 65.400 71.250 71.250 ;
        RECT 80.400 65.400 82.200 71.250 ;
        RECT 50.850 64.050 52.650 64.500 ;
        RECT 43.950 62.850 52.650 64.050 ;
        RECT 53.700 63.300 59.400 64.500 ;
        RECT 50.850 62.700 52.650 62.850 ;
        RECT 57.600 62.700 59.400 63.300 ;
        RECT 60.300 61.350 61.500 65.400 ;
        RECT 40.950 60.600 43.050 61.350 ;
        RECT 22.950 59.250 43.050 60.600 ;
        RECT 46.950 60.450 64.350 61.350 ;
        RECT 46.950 59.250 49.050 60.450 ;
        RECT 10.500 58.350 12.300 58.950 ;
        RECT 19.950 58.650 22.050 58.950 ;
        RECT 49.950 58.350 62.250 59.550 ;
        RECT 22.950 57.450 51.000 58.350 ;
        RECT 60.450 57.750 62.250 58.350 ;
        RECT 11.250 57.150 51.000 57.450 ;
        RECT 10.950 56.550 24.900 57.150 ;
        RECT 4.950 53.850 7.050 55.950 ;
        RECT 10.950 55.350 14.850 56.550 ;
        RECT 31.950 55.650 46.500 56.250 ;
        RECT 10.950 55.050 13.050 55.350 ;
        RECT 15.750 54.450 22.500 55.350 ;
        RECT 5.100 52.050 6.900 53.850 ;
        RECT 15.750 52.050 16.950 54.450 ;
        RECT 5.100 51.000 16.950 52.050 ;
        RECT 18.750 51.750 20.550 53.550 ;
        RECT 21.450 52.950 22.500 54.450 ;
        RECT 23.400 55.050 46.500 55.650 ;
        RECT 23.400 54.450 34.050 55.050 ;
        RECT 23.400 53.850 25.200 54.450 ;
        RECT 31.950 54.150 34.050 54.450 ;
        RECT 36.150 53.250 38.250 53.550 ;
        RECT 44.700 53.250 46.500 55.050 ;
        RECT 47.850 54.000 54.900 55.800 ;
        RECT 21.450 52.050 33.450 52.950 ;
        RECT 2.700 49.200 18.000 50.100 ;
        RECT 2.700 45.600 3.900 49.200 ;
        RECT 6.900 47.700 8.700 48.300 ;
        RECT 6.900 46.500 15.300 47.700 ;
        RECT 13.800 45.600 15.300 46.500 ;
        RECT 2.700 39.750 4.500 45.600 ;
        RECT 8.100 39.750 9.900 45.600 ;
        RECT 13.500 39.750 15.300 45.600 ;
        RECT 16.950 46.050 18.000 49.200 ;
        RECT 19.500 48.300 20.550 51.750 ;
        RECT 27.150 49.350 31.050 51.150 ;
        RECT 28.950 49.050 31.050 49.350 ;
        RECT 32.400 50.550 33.450 52.050 ;
        RECT 34.350 51.450 38.250 53.250 ;
        RECT 47.850 52.350 48.750 54.000 ;
        RECT 55.950 53.100 58.050 57.150 ;
        RECT 39.150 51.300 48.750 52.350 ;
        RECT 49.800 52.050 58.050 53.100 ;
        RECT 39.150 50.550 40.050 51.300 ;
        RECT 32.400 49.200 40.050 50.550 ;
        RECT 49.800 50.250 50.850 52.050 ;
        RECT 40.950 49.200 50.850 50.250 ;
        RECT 54.300 49.200 62.100 51.000 ;
        RECT 22.050 48.300 23.850 48.750 ;
        RECT 40.950 48.300 42.000 49.200 ;
        RECT 19.500 47.850 23.850 48.300 ;
        RECT 19.500 47.100 27.150 47.850 ;
        RECT 22.050 46.950 27.150 47.100 ;
        RECT 16.950 43.950 19.050 46.050 ;
        RECT 19.950 43.950 22.050 46.050 ;
        RECT 22.950 43.950 25.050 46.050 ;
        RECT 26.250 45.600 27.150 46.950 ;
        RECT 35.100 46.500 42.000 48.300 ;
        RECT 42.900 46.500 49.650 48.300 ;
        RECT 54.300 45.600 55.800 49.200 ;
        RECT 63.150 45.600 64.350 60.450 ;
        RECT 26.250 44.250 30.300 45.600 ;
        RECT 31.950 45.300 34.050 45.600 ;
        RECT 17.700 42.600 19.050 43.950 ;
        RECT 20.700 42.600 22.050 43.950 ;
        RECT 23.700 42.600 25.050 43.950 ;
        RECT 28.500 43.800 30.300 44.250 ;
        RECT 31.200 43.500 34.050 45.300 ;
        RECT 36.150 45.300 38.250 45.600 ;
        RECT 36.150 43.500 39.000 45.300 ;
        RECT 17.700 39.750 19.500 42.600 ;
        RECT 20.700 39.750 22.500 42.600 ;
        RECT 23.700 39.750 25.500 42.600 ;
        RECT 26.700 39.750 28.500 42.600 ;
        RECT 31.200 39.750 33.000 43.500 ;
        RECT 34.200 39.750 36.000 42.600 ;
        RECT 37.200 39.750 39.000 43.500 ;
        RECT 40.950 43.500 43.050 45.600 ;
        RECT 43.950 43.500 46.050 45.600 ;
        RECT 46.950 43.500 49.050 45.600 ;
        RECT 51.600 44.400 55.800 45.600 ;
        RECT 40.950 39.750 42.750 43.500 ;
        RECT 43.950 39.750 45.750 43.500 ;
        RECT 46.950 39.750 48.750 43.500 ;
        RECT 51.600 39.750 53.400 44.400 ;
        RECT 57.150 39.750 58.950 45.600 ;
        RECT 62.550 39.750 64.350 45.600 ;
        RECT 66.450 52.950 67.950 65.400 ;
        RECT 83.700 59.400 85.500 71.250 ;
        RECT 87.900 59.400 89.700 71.250 ;
        RECT 97.650 65.400 99.450 71.250 ;
        RECT 100.650 65.400 102.450 71.250 ;
        RECT 103.650 65.400 105.450 71.250 ;
        RECT 109.650 65.400 111.450 71.250 ;
        RECT 112.650 65.400 114.450 71.250 ;
        RECT 115.650 65.400 117.450 71.250 ;
        RECT 80.250 57.150 82.050 58.950 ;
        RECT 79.950 55.050 82.050 57.150 ;
        RECT 83.850 54.150 85.050 59.400 ;
        RECT 101.250 57.150 102.450 65.400 ;
        RECT 113.250 57.150 114.450 65.400 ;
        RECT 123.450 59.400 125.250 71.250 ;
        RECT 127.650 59.400 129.450 71.250 ;
        RECT 141.450 59.400 143.250 71.250 ;
        RECT 145.650 59.400 147.450 71.250 ;
        RECT 154.650 65.400 156.450 71.250 ;
        RECT 157.650 66.000 159.450 71.250 ;
        RECT 155.250 65.100 156.450 65.400 ;
        RECT 160.650 65.400 162.450 71.250 ;
        RECT 163.650 65.400 165.450 71.250 ;
        RECT 167.550 65.400 169.350 71.250 ;
        RECT 170.550 65.400 172.350 71.250 ;
        RECT 160.650 65.100 162.300 65.400 ;
        RECT 155.250 64.200 162.300 65.100 ;
        RECT 123.450 58.350 126.000 59.400 ;
        RECT 141.450 58.350 144.000 59.400 ;
        RECT 89.100 54.150 90.900 55.950 ;
        RECT 66.450 50.850 70.050 52.950 ;
        RECT 82.950 52.050 85.050 54.150 ;
        RECT 66.450 42.600 67.950 50.850 ;
        RECT 82.950 48.750 84.150 52.050 ;
        RECT 85.950 50.850 88.050 52.950 ;
        RECT 88.950 52.050 91.050 54.150 ;
        RECT 97.950 53.850 100.050 55.950 ;
        RECT 100.950 55.050 103.050 57.150 ;
        RECT 98.100 52.050 99.900 53.850 ;
        RECT 86.100 49.050 87.900 50.850 ;
        RECT 80.250 47.700 84.000 48.750 ;
        RECT 101.250 47.700 102.450 55.050 ;
        RECT 103.950 53.850 106.050 55.950 ;
        RECT 109.950 53.850 112.050 55.950 ;
        RECT 112.950 55.050 115.050 57.150 ;
        RECT 104.100 52.050 105.900 53.850 ;
        RECT 110.100 52.050 111.900 53.850 ;
        RECT 113.250 47.700 114.450 55.050 ;
        RECT 115.950 53.850 118.050 55.950 ;
        RECT 122.100 54.150 123.900 55.950 ;
        RECT 116.100 52.050 117.900 53.850 ;
        RECT 121.950 52.050 124.050 54.150 ;
        RECT 80.250 45.600 81.450 47.700 ;
        RECT 98.850 46.800 102.450 47.700 ;
        RECT 110.850 46.800 114.450 47.700 ;
        RECT 124.950 51.150 126.000 58.350 ;
        RECT 128.100 54.150 129.900 55.950 ;
        RECT 140.100 54.150 141.900 55.950 ;
        RECT 127.950 52.050 130.050 54.150 ;
        RECT 139.950 52.050 142.050 54.150 ;
        RECT 142.950 51.150 144.000 58.350 ;
        RECT 155.250 55.950 156.300 64.200 ;
        RECT 161.100 60.150 162.900 61.950 ;
        RECT 157.950 57.150 159.750 58.950 ;
        RECT 160.950 58.050 163.050 60.150 ;
        RECT 164.100 57.150 165.900 58.950 ;
        RECT 146.100 54.150 147.900 55.950 ;
        RECT 145.950 52.050 148.050 54.150 ;
        RECT 154.950 53.850 157.050 55.950 ;
        RECT 157.950 55.050 160.050 57.150 ;
        RECT 163.950 55.050 166.050 57.150 ;
        RECT 124.950 49.050 127.050 51.150 ;
        RECT 142.950 49.050 145.050 51.150 ;
        RECT 155.400 49.650 156.600 53.850 ;
        RECT 170.400 52.950 171.600 65.400 ;
        RECT 183.450 59.400 185.250 71.250 ;
        RECT 187.650 59.400 189.450 71.250 ;
        RECT 195.450 59.400 197.250 71.250 ;
        RECT 199.650 59.400 201.450 71.250 ;
        RECT 205.650 65.400 207.450 71.250 ;
        RECT 208.650 65.400 210.450 71.250 ;
        RECT 211.650 65.400 213.450 71.250 ;
        RECT 183.450 58.350 186.000 59.400 ;
        RECT 195.450 58.350 198.000 59.400 ;
        RECT 182.100 54.150 183.900 55.950 ;
        RECT 167.100 51.150 168.900 52.950 ;
        RECT 66.450 39.750 68.250 42.600 ;
        RECT 69.450 39.750 71.250 42.600 ;
        RECT 79.650 39.750 81.450 45.600 ;
        RECT 82.650 44.700 90.450 46.050 ;
        RECT 82.650 39.750 84.450 44.700 ;
        RECT 85.650 39.750 87.450 43.800 ;
        RECT 88.650 39.750 90.450 44.700 ;
        RECT 98.850 39.750 100.650 46.800 ;
        RECT 103.350 39.750 105.150 45.600 ;
        RECT 110.850 39.750 112.650 46.800 ;
        RECT 115.350 39.750 117.150 45.600 ;
        RECT 124.950 42.600 126.000 49.050 ;
        RECT 142.950 42.600 144.000 49.050 ;
        RECT 155.400 48.000 159.900 49.650 ;
        RECT 166.950 49.050 169.050 51.150 ;
        RECT 169.950 50.850 172.050 52.950 ;
        RECT 181.950 52.050 184.050 54.150 ;
        RECT 184.950 51.150 186.000 58.350 ;
        RECT 188.100 54.150 189.900 55.950 ;
        RECT 194.100 54.150 195.900 55.950 ;
        RECT 187.950 52.050 190.050 54.150 ;
        RECT 193.950 52.050 196.050 54.150 ;
        RECT 196.950 51.150 198.000 58.350 ;
        RECT 209.250 57.150 210.450 65.400 ;
        RECT 221.550 60.300 223.350 71.250 ;
        RECT 224.550 61.200 226.350 71.250 ;
        RECT 227.550 60.300 229.350 71.250 ;
        RECT 221.550 59.400 229.350 60.300 ;
        RECT 230.550 59.400 232.350 71.250 ;
        RECT 239.550 65.400 241.350 71.250 ;
        RECT 242.550 65.400 244.350 71.250 ;
        RECT 245.550 66.000 247.350 71.250 ;
        RECT 242.700 65.100 244.350 65.400 ;
        RECT 248.550 65.400 250.350 71.250 ;
        RECT 259.650 65.400 261.450 71.250 ;
        RECT 262.650 65.400 264.450 71.250 ;
        RECT 269.550 65.400 271.350 71.250 ;
        RECT 272.550 65.400 274.350 71.250 ;
        RECT 275.550 65.400 277.350 71.250 ;
        RECT 283.650 65.400 285.450 71.250 ;
        RECT 286.650 66.000 288.450 71.250 ;
        RECT 248.550 65.100 249.750 65.400 ;
        RECT 242.700 64.200 249.750 65.100 ;
        RECT 242.100 60.150 243.900 61.950 ;
        RECT 200.100 54.150 201.900 55.950 ;
        RECT 199.950 52.050 202.050 54.150 ;
        RECT 205.950 53.850 208.050 55.950 ;
        RECT 208.950 55.050 211.050 57.150 ;
        RECT 206.100 52.050 207.900 53.850 ;
        RECT 121.650 39.750 123.450 42.600 ;
        RECT 124.650 39.750 126.450 42.600 ;
        RECT 127.650 39.750 129.450 42.600 ;
        RECT 139.650 39.750 141.450 42.600 ;
        RECT 142.650 39.750 144.450 42.600 ;
        RECT 145.650 39.750 147.450 42.600 ;
        RECT 158.100 39.750 159.900 48.000 ;
        RECT 163.500 39.750 165.300 48.600 ;
        RECT 170.400 42.600 171.600 50.850 ;
        RECT 184.950 49.050 187.050 51.150 ;
        RECT 196.950 49.050 199.050 51.150 ;
        RECT 184.950 42.600 186.000 49.050 ;
        RECT 196.950 42.600 198.000 49.050 ;
        RECT 209.250 47.700 210.450 55.050 ;
        RECT 211.950 53.850 214.050 55.950 ;
        RECT 230.700 54.150 231.900 59.400 ;
        RECT 239.100 57.150 240.900 58.950 ;
        RECT 241.950 58.050 244.050 60.150 ;
        RECT 245.250 57.150 247.050 58.950 ;
        RECT 238.950 55.050 241.050 57.150 ;
        RECT 244.950 55.050 247.050 57.150 ;
        RECT 248.700 55.950 249.750 64.200 ;
        RECT 212.100 52.050 213.900 53.850 ;
        RECT 220.950 50.850 223.050 52.950 ;
        RECT 224.100 51.150 225.900 52.950 ;
        RECT 221.100 49.050 222.900 50.850 ;
        RECT 223.950 49.050 226.050 51.150 ;
        RECT 226.950 50.850 229.050 52.950 ;
        RECT 229.950 52.050 232.050 54.150 ;
        RECT 247.950 53.850 250.050 55.950 ;
        RECT 227.100 49.050 228.900 50.850 ;
        RECT 206.850 46.800 210.450 47.700 ;
        RECT 167.550 39.750 169.350 42.600 ;
        RECT 170.550 39.750 172.350 42.600 ;
        RECT 181.650 39.750 183.450 42.600 ;
        RECT 184.650 39.750 186.450 42.600 ;
        RECT 187.650 39.750 189.450 42.600 ;
        RECT 193.650 39.750 195.450 42.600 ;
        RECT 196.650 39.750 198.450 42.600 ;
        RECT 199.650 39.750 201.450 42.600 ;
        RECT 206.850 39.750 208.650 46.800 ;
        RECT 230.700 45.600 231.900 52.050 ;
        RECT 248.400 49.650 249.600 53.850 ;
        RECT 260.400 52.950 261.600 65.400 ;
        RECT 272.550 57.150 273.750 65.400 ;
        RECT 284.250 65.100 285.450 65.400 ;
        RECT 289.650 65.400 291.450 71.250 ;
        RECT 292.650 65.400 294.450 71.250 ;
        RECT 299.550 65.400 301.350 71.250 ;
        RECT 302.550 65.400 304.350 71.250 ;
        RECT 289.650 65.100 291.300 65.400 ;
        RECT 284.250 64.200 291.300 65.100 ;
        RECT 268.950 53.850 271.050 55.950 ;
        RECT 271.950 55.050 274.050 57.150 ;
        RECT 284.250 55.950 285.300 64.200 ;
        RECT 290.100 60.150 291.900 61.950 ;
        RECT 286.950 57.150 288.750 58.950 ;
        RECT 289.950 58.050 292.050 60.150 ;
        RECT 293.100 57.150 294.900 58.950 ;
        RECT 259.950 50.850 262.050 52.950 ;
        RECT 263.100 51.150 264.900 52.950 ;
        RECT 269.100 52.050 270.900 53.850 ;
        RECT 211.350 39.750 213.150 45.600 ;
        RECT 222.000 39.750 223.800 45.600 ;
        RECT 226.200 43.950 231.900 45.600 ;
        RECT 226.200 39.750 228.000 43.950 ;
        RECT 229.500 39.750 231.300 42.600 ;
        RECT 239.700 39.750 241.500 48.600 ;
        RECT 245.100 48.000 249.600 49.650 ;
        RECT 245.100 39.750 246.900 48.000 ;
        RECT 260.400 42.600 261.600 50.850 ;
        RECT 262.950 49.050 265.050 51.150 ;
        RECT 272.550 47.700 273.750 55.050 ;
        RECT 274.950 53.850 277.050 55.950 ;
        RECT 283.950 53.850 286.050 55.950 ;
        RECT 286.950 55.050 289.050 57.150 ;
        RECT 292.950 55.050 295.050 57.150 ;
        RECT 275.100 52.050 276.900 53.850 ;
        RECT 284.400 49.650 285.600 53.850 ;
        RECT 302.400 52.950 303.600 65.400 ;
        RECT 315.300 59.400 317.100 71.250 ;
        RECT 319.500 59.400 321.300 71.250 ;
        RECT 322.800 65.400 324.600 71.250 ;
        RECT 332.550 59.400 334.350 71.250 ;
        RECT 336.750 59.400 338.550 71.250 ;
        RECT 347.550 59.400 349.350 71.250 ;
        RECT 351.750 59.400 353.550 71.250 ;
        RECT 367.650 59.400 369.450 71.250 ;
        RECT 370.650 60.300 372.450 71.250 ;
        RECT 373.650 61.200 375.450 71.250 ;
        RECT 376.650 60.300 378.450 71.250 ;
        RECT 384.150 60.900 385.950 71.250 ;
        RECT 370.650 59.400 378.450 60.300 ;
        RECT 383.550 59.550 385.950 60.900 ;
        RECT 387.150 59.550 388.950 71.250 ;
        RECT 314.100 54.150 315.900 55.950 ;
        RECT 319.950 54.150 321.150 59.400 ;
        RECT 322.950 57.150 324.750 58.950 ;
        RECT 336.000 58.350 338.550 59.400 ;
        RECT 351.000 58.350 353.550 59.400 ;
        RECT 322.950 55.050 325.050 57.150 ;
        RECT 332.100 54.150 333.900 55.950 ;
        RECT 299.100 51.150 300.900 52.950 ;
        RECT 284.400 48.000 288.900 49.650 ;
        RECT 298.950 49.050 301.050 51.150 ;
        RECT 301.950 50.850 304.050 52.950 ;
        RECT 313.950 52.050 316.050 54.150 ;
        RECT 316.950 50.850 319.050 52.950 ;
        RECT 319.950 52.050 322.050 54.150 ;
        RECT 331.950 52.050 334.050 54.150 ;
        RECT 272.550 46.800 276.150 47.700 ;
        RECT 259.650 39.750 261.450 42.600 ;
        RECT 262.650 39.750 264.450 42.600 ;
        RECT 269.850 39.750 271.650 45.600 ;
        RECT 274.350 39.750 276.150 46.800 ;
        RECT 287.100 39.750 288.900 48.000 ;
        RECT 292.500 39.750 294.300 48.600 ;
        RECT 302.400 42.600 303.600 50.850 ;
        RECT 317.100 49.050 318.900 50.850 ;
        RECT 320.850 48.750 322.050 52.050 ;
        RECT 336.000 51.150 337.050 58.350 ;
        RECT 338.100 54.150 339.900 55.950 ;
        RECT 347.100 54.150 348.900 55.950 ;
        RECT 337.950 52.050 340.050 54.150 ;
        RECT 346.950 52.050 349.050 54.150 ;
        RECT 351.000 51.150 352.050 58.350 ;
        RECT 353.100 54.150 354.900 55.950 ;
        RECT 368.100 54.150 369.300 59.400 ;
        RECT 352.950 52.050 355.050 54.150 ;
        RECT 367.950 52.050 370.050 54.150 ;
        RECT 383.550 52.950 384.900 59.550 ;
        RECT 391.650 59.400 393.450 71.250 ;
        RECT 399.300 59.400 401.100 71.250 ;
        RECT 403.500 59.400 405.300 71.250 ;
        RECT 406.800 65.400 408.600 71.250 ;
        RECT 419.400 65.400 421.200 71.250 ;
        RECT 422.700 59.400 424.500 71.250 ;
        RECT 426.900 59.400 428.700 71.250 ;
        RECT 431.550 65.400 433.350 71.250 ;
        RECT 434.550 65.400 436.350 71.250 ;
        RECT 437.550 65.400 439.350 71.250 ;
        RECT 451.650 65.400 453.450 71.250 ;
        RECT 454.650 66.000 456.450 71.250 ;
        RECT 386.250 58.200 388.050 58.650 ;
        RECT 392.250 58.200 393.450 59.400 ;
        RECT 386.250 57.000 393.450 58.200 ;
        RECT 386.250 56.850 388.050 57.000 ;
        RECT 334.950 49.050 337.050 51.150 ;
        RECT 349.950 49.050 352.050 51.150 ;
        RECT 321.000 47.700 324.750 48.750 ;
        RECT 314.550 44.700 322.350 46.050 ;
        RECT 299.550 39.750 301.350 42.600 ;
        RECT 302.550 39.750 304.350 42.600 ;
        RECT 314.550 39.750 316.350 44.700 ;
        RECT 317.550 39.750 319.350 43.800 ;
        RECT 320.550 39.750 322.350 44.700 ;
        RECT 323.550 45.600 324.750 47.700 ;
        RECT 323.550 39.750 325.350 45.600 ;
        RECT 336.000 42.600 337.050 49.050 ;
        RECT 337.950 48.450 340.050 49.050 ;
        RECT 346.950 48.450 349.050 49.050 ;
        RECT 337.950 47.550 349.050 48.450 ;
        RECT 337.950 46.950 340.050 47.550 ;
        RECT 346.950 46.950 349.050 47.550 ;
        RECT 351.000 42.600 352.050 49.050 ;
        RECT 368.100 45.600 369.300 52.050 ;
        RECT 370.950 50.850 373.050 52.950 ;
        RECT 374.100 51.150 375.900 52.950 ;
        RECT 371.100 49.050 372.900 50.850 ;
        RECT 373.950 49.050 376.050 51.150 ;
        RECT 376.950 50.850 379.050 52.950 ;
        RECT 382.950 50.850 385.050 52.950 ;
        RECT 377.100 49.050 378.900 50.850 ;
        RECT 382.950 45.600 384.000 50.850 ;
        RECT 386.400 48.600 387.300 56.850 ;
        RECT 389.100 54.150 390.900 55.950 ;
        RECT 398.100 54.150 399.900 55.950 ;
        RECT 403.950 54.150 405.150 59.400 ;
        RECT 406.950 57.150 408.750 58.950 ;
        RECT 419.250 57.150 421.050 58.950 ;
        RECT 406.950 55.050 409.050 57.150 ;
        RECT 418.950 55.050 421.050 57.150 ;
        RECT 422.850 54.150 424.050 59.400 ;
        RECT 434.550 57.150 435.750 65.400 ;
        RECT 452.250 65.100 453.450 65.400 ;
        RECT 457.650 65.400 459.450 71.250 ;
        RECT 460.650 65.400 462.450 71.250 ;
        RECT 473.400 65.400 475.200 71.250 ;
        RECT 457.650 65.100 459.300 65.400 ;
        RECT 452.250 64.200 459.300 65.100 ;
        RECT 428.100 54.150 429.900 55.950 ;
        RECT 388.950 52.050 391.050 54.150 ;
        RECT 392.100 51.150 393.900 52.950 ;
        RECT 397.950 52.050 400.050 54.150 ;
        RECT 391.950 49.050 394.050 51.150 ;
        RECT 400.950 50.850 403.050 52.950 ;
        RECT 403.950 52.050 406.050 54.150 ;
        RECT 401.100 49.050 402.900 50.850 ;
        RECT 404.850 48.750 406.050 52.050 ;
        RECT 421.950 52.050 424.050 54.150 ;
        RECT 421.950 48.750 423.150 52.050 ;
        RECT 424.950 50.850 427.050 52.950 ;
        RECT 427.950 52.050 430.050 54.150 ;
        RECT 430.950 53.850 433.050 55.950 ;
        RECT 433.950 55.050 436.050 57.150 ;
        RECT 452.250 55.950 453.300 64.200 ;
        RECT 458.100 60.150 459.900 61.950 ;
        RECT 454.950 57.150 456.750 58.950 ;
        RECT 457.950 58.050 460.050 60.150 ;
        RECT 476.700 59.400 478.500 71.250 ;
        RECT 480.900 59.400 482.700 71.250 ;
        RECT 491.550 59.400 493.350 71.250 ;
        RECT 494.550 59.400 496.350 71.250 ;
        RECT 508.650 59.400 510.450 71.250 ;
        RECT 511.650 59.400 513.450 71.250 ;
        RECT 515.550 59.400 517.350 71.250 ;
        RECT 461.100 57.150 462.900 58.950 ;
        RECT 473.250 57.150 475.050 58.950 ;
        RECT 431.100 52.050 432.900 53.850 ;
        RECT 425.100 49.050 426.900 50.850 ;
        RECT 386.250 47.700 388.050 48.600 ;
        RECT 405.000 47.700 408.750 48.750 ;
        RECT 386.250 46.800 389.550 47.700 ;
        RECT 368.100 43.950 373.800 45.600 ;
        RECT 332.550 39.750 334.350 42.600 ;
        RECT 335.550 39.750 337.350 42.600 ;
        RECT 338.550 39.750 340.350 42.600 ;
        RECT 347.550 39.750 349.350 42.600 ;
        RECT 350.550 39.750 352.350 42.600 ;
        RECT 353.550 39.750 355.350 42.600 ;
        RECT 368.700 39.750 370.500 42.600 ;
        RECT 372.000 39.750 373.800 43.950 ;
        RECT 376.200 39.750 378.000 45.600 ;
        RECT 382.650 39.750 384.450 45.600 ;
        RECT 388.650 42.600 389.550 46.800 ;
        RECT 398.550 44.700 406.350 46.050 ;
        RECT 385.650 39.750 387.450 42.600 ;
        RECT 388.650 39.750 390.450 42.600 ;
        RECT 391.650 39.750 393.450 42.600 ;
        RECT 398.550 39.750 400.350 44.700 ;
        RECT 401.550 39.750 403.350 43.800 ;
        RECT 404.550 39.750 406.350 44.700 ;
        RECT 407.550 45.600 408.750 47.700 ;
        RECT 419.250 47.700 423.000 48.750 ;
        RECT 434.550 47.700 435.750 55.050 ;
        RECT 436.950 53.850 439.050 55.950 ;
        RECT 451.950 53.850 454.050 55.950 ;
        RECT 454.950 55.050 457.050 57.150 ;
        RECT 460.950 55.050 463.050 57.150 ;
        RECT 472.950 55.050 475.050 57.150 ;
        RECT 476.850 54.150 478.050 59.400 ;
        RECT 482.100 54.150 483.900 55.950 ;
        RECT 494.400 54.150 495.600 59.400 ;
        RECT 509.400 54.150 510.600 59.400 ;
        RECT 518.550 58.500 520.350 71.250 ;
        RECT 521.550 59.400 523.350 71.250 ;
        RECT 524.550 58.500 526.350 71.250 ;
        RECT 527.550 59.400 529.350 71.250 ;
        RECT 530.550 58.500 532.350 71.250 ;
        RECT 533.550 59.400 535.350 71.250 ;
        RECT 536.550 58.500 538.350 71.250 ;
        RECT 539.550 59.400 541.350 71.250 ;
        RECT 546.750 65.400 548.550 71.250 ;
        RECT 549.750 65.400 551.550 71.250 ;
        RECT 553.500 65.400 555.300 71.250 ;
        RECT 556.500 65.400 558.300 71.250 ;
        RECT 559.500 65.400 561.300 71.250 ;
        RECT 518.550 57.300 522.450 58.500 ;
        RECT 524.550 57.300 528.300 58.500 ;
        RECT 530.550 57.300 534.300 58.500 ;
        RECT 536.550 57.300 539.250 58.500 ;
        RECT 437.100 52.050 438.900 53.850 ;
        RECT 452.400 49.650 453.600 53.850 ;
        RECT 475.950 52.050 478.050 54.150 ;
        RECT 452.400 48.000 456.900 49.650 ;
        RECT 475.950 48.750 477.150 52.050 ;
        RECT 478.950 50.850 481.050 52.950 ;
        RECT 481.950 52.050 484.050 54.150 ;
        RECT 490.950 50.850 493.050 52.950 ;
        RECT 493.950 52.050 496.050 54.150 ;
        RECT 508.950 52.050 511.050 54.150 ;
        RECT 479.100 49.050 480.900 50.850 ;
        RECT 491.100 49.050 492.900 50.850 ;
        RECT 419.250 45.600 420.450 47.700 ;
        RECT 434.550 46.800 438.150 47.700 ;
        RECT 407.550 39.750 409.350 45.600 ;
        RECT 418.650 39.750 420.450 45.600 ;
        RECT 421.650 44.700 429.450 46.050 ;
        RECT 421.650 39.750 423.450 44.700 ;
        RECT 424.650 39.750 426.450 43.800 ;
        RECT 427.650 39.750 429.450 44.700 ;
        RECT 431.850 39.750 433.650 45.600 ;
        RECT 436.350 39.750 438.150 46.800 ;
        RECT 455.100 39.750 456.900 48.000 ;
        RECT 460.500 39.750 462.300 48.600 ;
        RECT 473.250 47.700 477.000 48.750 ;
        RECT 473.250 45.600 474.450 47.700 ;
        RECT 472.650 39.750 474.450 45.600 ;
        RECT 475.650 44.700 483.450 46.050 ;
        RECT 494.400 45.600 495.600 52.050 ;
        RECT 509.400 45.600 510.600 52.050 ;
        RECT 511.950 50.850 514.050 52.950 ;
        RECT 517.950 50.850 520.050 52.950 ;
        RECT 512.100 49.050 513.900 50.850 ;
        RECT 518.100 49.050 519.900 50.850 ;
        RECT 521.250 50.400 522.450 57.300 ;
        RECT 527.100 50.400 528.300 57.300 ;
        RECT 533.100 50.400 534.300 57.300 ;
        RECT 538.200 52.950 539.250 57.300 ;
        RECT 550.050 52.950 551.550 65.400 ;
        RECT 556.500 61.350 557.700 65.400 ;
        RECT 562.500 64.500 564.300 71.250 ;
        RECT 565.500 65.400 567.300 71.250 ;
        RECT 569.250 68.400 571.050 71.250 ;
        RECT 569.400 67.200 570.900 68.400 ;
        RECT 568.800 65.100 570.900 67.200 ;
        RECT 572.250 64.950 574.050 71.250 ;
        RECT 575.250 68.400 577.050 71.250 ;
        RECT 558.600 63.300 564.300 64.500 ;
        RECT 565.350 64.050 567.150 64.500 ;
        RECT 571.950 64.050 574.050 64.950 ;
        RECT 558.600 62.700 560.400 63.300 ;
        RECT 565.350 62.850 574.050 64.050 ;
        RECT 565.350 62.700 567.150 62.850 ;
        RECT 575.550 61.350 576.900 68.400 ;
        RECT 579.000 64.500 580.800 71.250 ;
        RECT 582.000 65.400 583.800 71.250 ;
        RECT 585.000 65.400 586.800 71.250 ;
        RECT 588.750 65.400 590.550 71.250 ;
        RECT 591.750 68.400 593.700 71.250 ;
        RECT 594.750 68.400 596.850 71.250 ;
        RECT 597.750 68.400 600.150 71.250 ;
        RECT 592.500 67.050 593.700 68.400 ;
        RECT 595.950 67.050 596.850 68.400 ;
        RECT 598.950 67.050 600.150 68.400 ;
        RECT 601.500 67.950 603.300 71.250 ;
        RECT 592.500 65.400 595.050 67.050 ;
        RECT 585.000 64.500 586.350 65.400 ;
        RECT 592.950 64.950 595.050 65.400 ;
        RECT 595.950 64.950 598.050 67.050 ;
        RECT 598.950 64.950 601.050 67.050 ;
        RECT 579.000 64.200 582.000 64.500 ;
        RECT 578.100 62.400 582.000 64.200 ;
        RECT 583.950 62.850 586.350 64.500 ;
        RECT 583.950 62.400 586.050 62.850 ;
        RECT 604.500 62.700 606.300 71.250 ;
        RECT 607.500 65.400 609.300 71.250 ;
        RECT 610.500 65.400 612.300 71.250 ;
        RECT 613.500 65.400 615.300 71.250 ;
        RECT 618.750 65.400 620.550 71.250 ;
        RECT 621.750 65.400 623.550 71.250 ;
        RECT 625.500 65.400 627.300 71.250 ;
        RECT 628.500 65.400 630.300 71.250 ;
        RECT 631.500 65.400 633.300 71.250 ;
        RECT 611.250 64.500 612.300 65.400 ;
        RECT 611.250 63.600 615.300 64.500 ;
        RECT 593.100 61.650 610.800 62.700 ;
        RECT 538.200 50.850 541.050 52.950 ;
        RECT 547.950 50.850 551.550 52.950 ;
        RECT 521.250 48.600 525.300 50.400 ;
        RECT 527.100 48.600 531.300 50.400 ;
        RECT 533.100 48.600 537.300 50.400 ;
        RECT 521.250 47.700 522.450 48.600 ;
        RECT 527.100 47.700 528.300 48.600 ;
        RECT 533.100 47.700 534.300 48.600 ;
        RECT 538.200 47.700 539.250 50.850 ;
        RECT 518.400 46.500 522.450 47.700 ;
        RECT 524.550 46.500 528.300 47.700 ;
        RECT 530.400 46.500 534.300 47.700 ;
        RECT 536.400 46.650 539.250 47.700 ;
        RECT 536.400 46.500 539.100 46.650 ;
        RECT 518.400 45.600 520.200 46.500 ;
        RECT 475.650 39.750 477.450 44.700 ;
        RECT 478.650 39.750 480.450 43.800 ;
        RECT 481.650 39.750 483.450 44.700 ;
        RECT 491.550 39.750 493.350 45.600 ;
        RECT 494.550 39.750 496.350 45.600 ;
        RECT 508.650 39.750 510.450 45.600 ;
        RECT 511.650 39.750 513.450 45.600 ;
        RECT 515.550 39.750 517.350 45.600 ;
        RECT 518.550 39.750 520.350 45.600 ;
        RECT 521.550 39.750 523.350 45.600 ;
        RECT 524.550 39.750 526.350 46.500 ;
        RECT 530.400 45.600 532.200 46.500 ;
        RECT 536.400 45.600 538.200 46.500 ;
        RECT 527.550 39.750 529.350 45.600 ;
        RECT 530.550 39.750 532.350 45.600 ;
        RECT 533.550 39.750 535.350 45.600 ;
        RECT 536.550 39.750 538.350 45.600 ;
        RECT 539.550 39.750 541.350 45.600 ;
        RECT 550.050 42.600 551.550 50.850 ;
        RECT 546.750 39.750 548.550 42.600 ;
        RECT 549.750 39.750 551.550 42.600 ;
        RECT 553.650 60.450 571.050 61.350 ;
        RECT 553.650 45.600 554.850 60.450 ;
        RECT 555.750 58.350 568.050 59.550 ;
        RECT 568.950 59.250 571.050 60.450 ;
        RECT 574.950 60.600 577.050 61.350 ;
        RECT 593.100 60.600 595.050 61.650 ;
        RECT 609.000 60.900 610.800 61.650 ;
        RECT 574.950 59.250 595.050 60.600 ;
        RECT 595.950 60.150 598.050 60.750 ;
        RECT 595.950 58.950 607.500 60.150 ;
        RECT 595.950 58.650 598.050 58.950 ;
        RECT 605.700 58.350 607.500 58.950 ;
        RECT 555.750 57.750 557.550 58.350 ;
        RECT 567.000 57.450 595.050 58.350 ;
        RECT 567.000 57.150 606.750 57.450 ;
        RECT 559.950 53.100 562.050 57.150 ;
        RECT 593.100 56.550 607.050 57.150 ;
        RECT 563.100 54.000 570.150 55.800 ;
        RECT 559.950 52.050 568.200 53.100 ;
        RECT 555.900 49.200 563.700 51.000 ;
        RECT 567.150 50.250 568.200 52.050 ;
        RECT 569.250 52.350 570.150 54.000 ;
        RECT 571.500 55.650 586.050 56.250 ;
        RECT 571.500 55.050 594.600 55.650 ;
        RECT 603.150 55.350 607.050 56.550 ;
        RECT 571.500 53.250 573.300 55.050 ;
        RECT 583.950 54.450 594.600 55.050 ;
        RECT 583.950 54.150 586.050 54.450 ;
        RECT 592.800 53.850 594.600 54.450 ;
        RECT 595.500 54.450 602.250 55.350 ;
        RECT 604.950 55.050 607.050 55.350 ;
        RECT 579.750 53.250 581.850 53.550 ;
        RECT 569.250 51.300 578.850 52.350 ;
        RECT 579.750 51.450 583.650 53.250 ;
        RECT 595.500 52.950 596.550 54.450 ;
        RECT 584.550 52.050 596.550 52.950 ;
        RECT 577.950 50.550 578.850 51.300 ;
        RECT 584.550 50.550 585.600 52.050 ;
        RECT 597.450 51.750 599.250 53.550 ;
        RECT 601.050 52.050 602.250 54.450 ;
        RECT 610.950 53.850 613.050 55.950 ;
        RECT 611.100 52.050 612.900 53.850 ;
        RECT 567.150 49.200 577.050 50.250 ;
        RECT 577.950 49.200 585.600 50.550 ;
        RECT 586.950 49.350 590.850 51.150 ;
        RECT 562.200 45.600 563.700 49.200 ;
        RECT 576.000 48.300 577.050 49.200 ;
        RECT 586.950 49.050 589.050 49.350 ;
        RECT 594.150 48.300 595.950 48.750 ;
        RECT 597.450 48.300 598.500 51.750 ;
        RECT 601.050 51.000 612.900 52.050 ;
        RECT 614.100 50.100 615.300 63.600 ;
        RECT 622.050 52.950 623.550 65.400 ;
        RECT 628.500 61.350 629.700 65.400 ;
        RECT 634.500 64.500 636.300 71.250 ;
        RECT 637.500 65.400 639.300 71.250 ;
        RECT 641.250 68.400 643.050 71.250 ;
        RECT 641.400 67.200 642.900 68.400 ;
        RECT 640.800 65.100 642.900 67.200 ;
        RECT 644.250 64.950 646.050 71.250 ;
        RECT 647.250 68.400 649.050 71.250 ;
        RECT 630.600 63.300 636.300 64.500 ;
        RECT 637.350 64.050 639.150 64.500 ;
        RECT 643.950 64.050 646.050 64.950 ;
        RECT 630.600 62.700 632.400 63.300 ;
        RECT 637.350 62.850 646.050 64.050 ;
        RECT 637.350 62.700 639.150 62.850 ;
        RECT 647.550 61.350 648.900 68.400 ;
        RECT 651.000 64.500 652.800 71.250 ;
        RECT 654.000 65.400 655.800 71.250 ;
        RECT 657.000 65.400 658.800 71.250 ;
        RECT 660.750 65.400 662.550 71.250 ;
        RECT 663.750 68.400 665.700 71.250 ;
        RECT 666.750 68.400 668.850 71.250 ;
        RECT 669.750 68.400 672.150 71.250 ;
        RECT 664.500 67.050 665.700 68.400 ;
        RECT 667.950 67.050 668.850 68.400 ;
        RECT 670.950 67.050 672.150 68.400 ;
        RECT 673.500 67.950 675.300 71.250 ;
        RECT 664.500 65.400 667.050 67.050 ;
        RECT 657.000 64.500 658.350 65.400 ;
        RECT 664.950 64.950 667.050 65.400 ;
        RECT 667.950 64.950 670.050 67.050 ;
        RECT 670.950 64.950 673.050 67.050 ;
        RECT 651.000 64.200 654.000 64.500 ;
        RECT 650.100 62.400 654.000 64.200 ;
        RECT 655.950 62.850 658.350 64.500 ;
        RECT 655.950 62.400 658.050 62.850 ;
        RECT 676.500 62.700 678.300 71.250 ;
        RECT 679.500 65.400 681.300 71.250 ;
        RECT 682.500 65.400 684.300 71.250 ;
        RECT 685.500 65.400 687.300 71.250 ;
        RECT 697.650 65.400 699.450 71.250 ;
        RECT 700.650 65.400 702.450 71.250 ;
        RECT 703.650 65.400 705.450 71.250 ;
        RECT 715.650 65.400 717.450 71.250 ;
        RECT 718.650 66.000 720.450 71.250 ;
        RECT 683.250 64.500 684.300 65.400 ;
        RECT 683.250 63.600 687.300 64.500 ;
        RECT 665.100 61.650 682.800 62.700 ;
        RECT 619.950 50.850 623.550 52.950 ;
        RECT 568.350 46.500 575.100 48.300 ;
        RECT 576.000 46.500 582.900 48.300 ;
        RECT 594.150 47.850 598.500 48.300 ;
        RECT 590.850 47.100 598.500 47.850 ;
        RECT 600.000 49.200 615.300 50.100 ;
        RECT 590.850 46.950 595.950 47.100 ;
        RECT 590.850 45.600 591.750 46.950 ;
        RECT 600.000 46.050 601.050 49.200 ;
        RECT 609.300 47.700 611.100 48.300 ;
        RECT 553.650 39.750 555.450 45.600 ;
        RECT 559.050 39.750 560.850 45.600 ;
        RECT 562.200 44.400 566.400 45.600 ;
        RECT 564.600 39.750 566.400 44.400 ;
        RECT 568.950 43.500 571.050 45.600 ;
        RECT 571.950 43.500 574.050 45.600 ;
        RECT 574.950 43.500 577.050 45.600 ;
        RECT 579.750 45.300 581.850 45.600 ;
        RECT 569.250 39.750 571.050 43.500 ;
        RECT 572.250 39.750 574.050 43.500 ;
        RECT 575.250 39.750 577.050 43.500 ;
        RECT 579.000 43.500 581.850 45.300 ;
        RECT 583.950 45.300 586.050 45.600 ;
        RECT 583.950 43.500 586.800 45.300 ;
        RECT 587.700 44.250 591.750 45.600 ;
        RECT 587.700 43.800 589.500 44.250 ;
        RECT 592.950 43.950 595.050 46.050 ;
        RECT 595.950 43.950 598.050 46.050 ;
        RECT 598.950 43.950 601.050 46.050 ;
        RECT 602.700 46.500 611.100 47.700 ;
        RECT 602.700 45.600 604.200 46.500 ;
        RECT 614.100 45.600 615.300 49.200 ;
        RECT 579.000 39.750 580.800 43.500 ;
        RECT 582.000 39.750 583.800 42.600 ;
        RECT 585.000 39.750 586.800 43.500 ;
        RECT 592.950 42.600 594.300 43.950 ;
        RECT 595.950 42.600 597.300 43.950 ;
        RECT 598.950 42.600 600.300 43.950 ;
        RECT 589.500 39.750 591.300 42.600 ;
        RECT 592.500 39.750 594.300 42.600 ;
        RECT 595.500 39.750 597.300 42.600 ;
        RECT 598.500 39.750 600.300 42.600 ;
        RECT 602.700 39.750 604.500 45.600 ;
        RECT 608.100 39.750 609.900 45.600 ;
        RECT 613.500 39.750 615.300 45.600 ;
        RECT 622.050 42.600 623.550 50.850 ;
        RECT 618.750 39.750 620.550 42.600 ;
        RECT 621.750 39.750 623.550 42.600 ;
        RECT 625.650 60.450 643.050 61.350 ;
        RECT 625.650 45.600 626.850 60.450 ;
        RECT 627.750 58.350 640.050 59.550 ;
        RECT 640.950 59.250 643.050 60.450 ;
        RECT 646.950 60.600 649.050 61.350 ;
        RECT 665.100 60.600 667.050 61.650 ;
        RECT 681.000 60.900 682.800 61.650 ;
        RECT 646.950 59.250 667.050 60.600 ;
        RECT 667.950 60.150 670.050 60.750 ;
        RECT 667.950 58.950 679.500 60.150 ;
        RECT 667.950 58.650 670.050 58.950 ;
        RECT 677.700 58.350 679.500 58.950 ;
        RECT 627.750 57.750 629.550 58.350 ;
        RECT 639.000 57.450 667.050 58.350 ;
        RECT 639.000 57.150 678.750 57.450 ;
        RECT 631.950 53.100 634.050 57.150 ;
        RECT 665.100 56.550 679.050 57.150 ;
        RECT 635.100 54.000 642.150 55.800 ;
        RECT 631.950 52.050 640.200 53.100 ;
        RECT 627.900 49.200 635.700 51.000 ;
        RECT 639.150 50.250 640.200 52.050 ;
        RECT 641.250 52.350 642.150 54.000 ;
        RECT 643.500 55.650 658.050 56.250 ;
        RECT 643.500 55.050 666.600 55.650 ;
        RECT 675.150 55.350 679.050 56.550 ;
        RECT 643.500 53.250 645.300 55.050 ;
        RECT 655.950 54.450 666.600 55.050 ;
        RECT 655.950 54.150 658.050 54.450 ;
        RECT 664.800 53.850 666.600 54.450 ;
        RECT 667.500 54.450 674.250 55.350 ;
        RECT 676.950 55.050 679.050 55.350 ;
        RECT 651.750 53.250 653.850 53.550 ;
        RECT 641.250 51.300 650.850 52.350 ;
        RECT 651.750 51.450 655.650 53.250 ;
        RECT 667.500 52.950 668.550 54.450 ;
        RECT 656.550 52.050 668.550 52.950 ;
        RECT 649.950 50.550 650.850 51.300 ;
        RECT 656.550 50.550 657.600 52.050 ;
        RECT 669.450 51.750 671.250 53.550 ;
        RECT 673.050 52.050 674.250 54.450 ;
        RECT 682.950 53.850 685.050 55.950 ;
        RECT 683.100 52.050 684.900 53.850 ;
        RECT 639.150 49.200 649.050 50.250 ;
        RECT 649.950 49.200 657.600 50.550 ;
        RECT 658.950 49.350 662.850 51.150 ;
        RECT 634.200 45.600 635.700 49.200 ;
        RECT 648.000 48.300 649.050 49.200 ;
        RECT 658.950 49.050 661.050 49.350 ;
        RECT 666.150 48.300 667.950 48.750 ;
        RECT 669.450 48.300 670.500 51.750 ;
        RECT 673.050 51.000 684.900 52.050 ;
        RECT 686.100 50.100 687.300 63.600 ;
        RECT 701.250 57.150 702.450 65.400 ;
        RECT 716.250 65.100 717.450 65.400 ;
        RECT 721.650 65.400 723.450 71.250 ;
        RECT 724.650 65.400 726.450 71.250 ;
        RECT 721.650 65.100 723.300 65.400 ;
        RECT 716.250 64.200 723.300 65.100 ;
        RECT 703.950 60.450 706.050 61.050 ;
        RECT 712.950 60.450 715.050 61.050 ;
        RECT 703.950 59.550 715.050 60.450 ;
        RECT 703.950 58.950 706.050 59.550 ;
        RECT 712.950 58.950 715.050 59.550 ;
        RECT 697.950 53.850 700.050 55.950 ;
        RECT 700.950 55.050 703.050 57.150 ;
        RECT 716.250 55.950 717.300 64.200 ;
        RECT 722.100 60.150 723.900 61.950 ;
        RECT 718.950 57.150 720.750 58.950 ;
        RECT 721.950 58.050 724.050 60.150 ;
        RECT 734.550 59.400 736.350 71.250 ;
        RECT 725.100 57.150 726.900 58.950 ;
        RECT 737.550 58.500 739.350 71.250 ;
        RECT 740.550 59.400 742.350 71.250 ;
        RECT 743.550 58.500 745.350 71.250 ;
        RECT 746.550 59.400 748.350 71.250 ;
        RECT 749.550 58.500 751.350 71.250 ;
        RECT 752.550 59.400 754.350 71.250 ;
        RECT 755.550 58.500 757.350 71.250 ;
        RECT 758.550 59.400 760.350 71.250 ;
        RECT 767.550 59.400 769.350 71.250 ;
        RECT 770.550 59.400 772.350 71.250 ;
        RECT 777.750 65.400 779.550 71.250 ;
        RECT 780.750 65.400 782.550 71.250 ;
        RECT 784.500 65.400 786.300 71.250 ;
        RECT 787.500 65.400 789.300 71.250 ;
        RECT 790.500 65.400 792.300 71.250 ;
        RECT 737.550 57.300 741.450 58.500 ;
        RECT 743.550 57.300 747.300 58.500 ;
        RECT 749.550 57.300 753.300 58.500 ;
        RECT 755.550 57.300 758.250 58.500 ;
        RECT 698.100 52.050 699.900 53.850 ;
        RECT 640.350 46.500 647.100 48.300 ;
        RECT 648.000 46.500 654.900 48.300 ;
        RECT 666.150 47.850 670.500 48.300 ;
        RECT 662.850 47.100 670.500 47.850 ;
        RECT 672.000 49.200 687.300 50.100 ;
        RECT 662.850 46.950 667.950 47.100 ;
        RECT 662.850 45.600 663.750 46.950 ;
        RECT 672.000 46.050 673.050 49.200 ;
        RECT 681.300 47.700 683.100 48.300 ;
        RECT 625.650 39.750 627.450 45.600 ;
        RECT 631.050 39.750 632.850 45.600 ;
        RECT 634.200 44.400 638.400 45.600 ;
        RECT 636.600 39.750 638.400 44.400 ;
        RECT 640.950 43.500 643.050 45.600 ;
        RECT 643.950 43.500 646.050 45.600 ;
        RECT 646.950 43.500 649.050 45.600 ;
        RECT 651.750 45.300 653.850 45.600 ;
        RECT 641.250 39.750 643.050 43.500 ;
        RECT 644.250 39.750 646.050 43.500 ;
        RECT 647.250 39.750 649.050 43.500 ;
        RECT 651.000 43.500 653.850 45.300 ;
        RECT 655.950 45.300 658.050 45.600 ;
        RECT 655.950 43.500 658.800 45.300 ;
        RECT 659.700 44.250 663.750 45.600 ;
        RECT 659.700 43.800 661.500 44.250 ;
        RECT 664.950 43.950 667.050 46.050 ;
        RECT 667.950 43.950 670.050 46.050 ;
        RECT 670.950 43.950 673.050 46.050 ;
        RECT 674.700 46.500 683.100 47.700 ;
        RECT 674.700 45.600 676.200 46.500 ;
        RECT 686.100 45.600 687.300 49.200 ;
        RECT 701.250 47.700 702.450 55.050 ;
        RECT 703.950 53.850 706.050 55.950 ;
        RECT 715.950 53.850 718.050 55.950 ;
        RECT 718.950 55.050 721.050 57.150 ;
        RECT 724.950 55.050 727.050 57.150 ;
        RECT 704.100 52.050 705.900 53.850 ;
        RECT 716.400 49.650 717.600 53.850 ;
        RECT 736.950 50.850 739.050 52.950 ;
        RECT 716.400 48.000 720.900 49.650 ;
        RECT 737.100 49.050 738.900 50.850 ;
        RECT 740.250 50.400 741.450 57.300 ;
        RECT 746.100 50.400 747.300 57.300 ;
        RECT 752.100 50.400 753.300 57.300 ;
        RECT 757.200 52.950 758.250 57.300 ;
        RECT 770.400 54.150 771.600 59.400 ;
        RECT 757.200 50.850 760.050 52.950 ;
        RECT 766.950 50.850 769.050 52.950 ;
        RECT 769.950 52.050 772.050 54.150 ;
        RECT 781.050 52.950 782.550 65.400 ;
        RECT 787.500 61.350 788.700 65.400 ;
        RECT 793.500 64.500 795.300 71.250 ;
        RECT 796.500 65.400 798.300 71.250 ;
        RECT 800.250 68.400 802.050 71.250 ;
        RECT 800.400 67.200 801.900 68.400 ;
        RECT 799.800 65.100 801.900 67.200 ;
        RECT 803.250 64.950 805.050 71.250 ;
        RECT 806.250 68.400 808.050 71.250 ;
        RECT 789.600 63.300 795.300 64.500 ;
        RECT 796.350 64.050 798.150 64.500 ;
        RECT 802.950 64.050 805.050 64.950 ;
        RECT 789.600 62.700 791.400 63.300 ;
        RECT 796.350 62.850 805.050 64.050 ;
        RECT 796.350 62.700 798.150 62.850 ;
        RECT 806.550 61.350 807.900 68.400 ;
        RECT 810.000 64.500 811.800 71.250 ;
        RECT 813.000 65.400 814.800 71.250 ;
        RECT 816.000 65.400 817.800 71.250 ;
        RECT 819.750 65.400 821.550 71.250 ;
        RECT 822.750 68.400 824.700 71.250 ;
        RECT 825.750 68.400 827.850 71.250 ;
        RECT 828.750 68.400 831.150 71.250 ;
        RECT 823.500 67.050 824.700 68.400 ;
        RECT 826.950 67.050 827.850 68.400 ;
        RECT 829.950 67.050 831.150 68.400 ;
        RECT 832.500 67.950 834.300 71.250 ;
        RECT 823.500 65.400 826.050 67.050 ;
        RECT 816.000 64.500 817.350 65.400 ;
        RECT 823.950 64.950 826.050 65.400 ;
        RECT 826.950 64.950 829.050 67.050 ;
        RECT 829.950 64.950 832.050 67.050 ;
        RECT 810.000 64.200 813.000 64.500 ;
        RECT 809.100 62.400 813.000 64.200 ;
        RECT 814.950 62.850 817.350 64.500 ;
        RECT 814.950 62.400 817.050 62.850 ;
        RECT 835.500 62.700 837.300 71.250 ;
        RECT 838.500 65.400 840.300 71.250 ;
        RECT 841.500 65.400 843.300 71.250 ;
        RECT 844.500 65.400 846.300 71.250 ;
        RECT 842.250 64.500 843.300 65.400 ;
        RECT 842.250 63.600 846.300 64.500 ;
        RECT 824.100 61.650 841.800 62.700 ;
        RECT 740.250 48.600 744.300 50.400 ;
        RECT 746.100 48.600 750.300 50.400 ;
        RECT 752.100 48.600 756.300 50.400 ;
        RECT 651.000 39.750 652.800 43.500 ;
        RECT 654.000 39.750 655.800 42.600 ;
        RECT 657.000 39.750 658.800 43.500 ;
        RECT 664.950 42.600 666.300 43.950 ;
        RECT 667.950 42.600 669.300 43.950 ;
        RECT 670.950 42.600 672.300 43.950 ;
        RECT 661.500 39.750 663.300 42.600 ;
        RECT 664.500 39.750 666.300 42.600 ;
        RECT 667.500 39.750 669.300 42.600 ;
        RECT 670.500 39.750 672.300 42.600 ;
        RECT 674.700 39.750 676.500 45.600 ;
        RECT 680.100 39.750 681.900 45.600 ;
        RECT 685.500 39.750 687.300 45.600 ;
        RECT 698.850 46.800 702.450 47.700 ;
        RECT 698.850 39.750 700.650 46.800 ;
        RECT 703.350 39.750 705.150 45.600 ;
        RECT 719.100 39.750 720.900 48.000 ;
        RECT 724.500 39.750 726.300 48.600 ;
        RECT 740.250 47.700 741.450 48.600 ;
        RECT 746.100 47.700 747.300 48.600 ;
        RECT 752.100 47.700 753.300 48.600 ;
        RECT 757.200 47.700 758.250 50.850 ;
        RECT 767.100 49.050 768.900 50.850 ;
        RECT 737.400 46.500 741.450 47.700 ;
        RECT 743.550 46.500 747.300 47.700 ;
        RECT 749.400 46.500 753.300 47.700 ;
        RECT 755.400 46.650 758.250 47.700 ;
        RECT 755.400 46.500 758.100 46.650 ;
        RECT 737.400 45.600 739.200 46.500 ;
        RECT 734.550 39.750 736.350 45.600 ;
        RECT 737.550 39.750 739.350 45.600 ;
        RECT 740.550 39.750 742.350 45.600 ;
        RECT 743.550 39.750 745.350 46.500 ;
        RECT 749.400 45.600 751.200 46.500 ;
        RECT 755.400 45.600 757.200 46.500 ;
        RECT 770.400 45.600 771.600 52.050 ;
        RECT 778.950 50.850 782.550 52.950 ;
        RECT 746.550 39.750 748.350 45.600 ;
        RECT 749.550 39.750 751.350 45.600 ;
        RECT 752.550 39.750 754.350 45.600 ;
        RECT 755.550 39.750 757.350 45.600 ;
        RECT 758.550 39.750 760.350 45.600 ;
        RECT 767.550 39.750 769.350 45.600 ;
        RECT 770.550 39.750 772.350 45.600 ;
        RECT 781.050 42.600 782.550 50.850 ;
        RECT 777.750 39.750 779.550 42.600 ;
        RECT 780.750 39.750 782.550 42.600 ;
        RECT 784.650 60.450 802.050 61.350 ;
        RECT 784.650 45.600 785.850 60.450 ;
        RECT 786.750 58.350 799.050 59.550 ;
        RECT 799.950 59.250 802.050 60.450 ;
        RECT 805.950 60.600 808.050 61.350 ;
        RECT 824.100 60.600 826.050 61.650 ;
        RECT 840.000 60.900 841.800 61.650 ;
        RECT 805.950 59.250 826.050 60.600 ;
        RECT 826.950 60.150 829.050 60.750 ;
        RECT 826.950 58.950 838.500 60.150 ;
        RECT 826.950 58.650 829.050 58.950 ;
        RECT 836.700 58.350 838.500 58.950 ;
        RECT 786.750 57.750 788.550 58.350 ;
        RECT 798.000 57.450 826.050 58.350 ;
        RECT 798.000 57.150 837.750 57.450 ;
        RECT 790.950 53.100 793.050 57.150 ;
        RECT 824.100 56.550 838.050 57.150 ;
        RECT 794.100 54.000 801.150 55.800 ;
        RECT 790.950 52.050 799.200 53.100 ;
        RECT 786.900 49.200 794.700 51.000 ;
        RECT 798.150 50.250 799.200 52.050 ;
        RECT 800.250 52.350 801.150 54.000 ;
        RECT 802.500 55.650 817.050 56.250 ;
        RECT 802.500 55.050 825.600 55.650 ;
        RECT 834.150 55.350 838.050 56.550 ;
        RECT 802.500 53.250 804.300 55.050 ;
        RECT 814.950 54.450 825.600 55.050 ;
        RECT 814.950 54.150 817.050 54.450 ;
        RECT 823.800 53.850 825.600 54.450 ;
        RECT 826.500 54.450 833.250 55.350 ;
        RECT 835.950 55.050 838.050 55.350 ;
        RECT 810.750 53.250 812.850 53.550 ;
        RECT 800.250 51.300 809.850 52.350 ;
        RECT 810.750 51.450 814.650 53.250 ;
        RECT 826.500 52.950 827.550 54.450 ;
        RECT 815.550 52.050 827.550 52.950 ;
        RECT 808.950 50.550 809.850 51.300 ;
        RECT 815.550 50.550 816.600 52.050 ;
        RECT 828.450 51.750 830.250 53.550 ;
        RECT 832.050 52.050 833.250 54.450 ;
        RECT 841.950 53.850 844.050 55.950 ;
        RECT 842.100 52.050 843.900 53.850 ;
        RECT 798.150 49.200 808.050 50.250 ;
        RECT 808.950 49.200 816.600 50.550 ;
        RECT 817.950 49.350 821.850 51.150 ;
        RECT 793.200 45.600 794.700 49.200 ;
        RECT 807.000 48.300 808.050 49.200 ;
        RECT 817.950 49.050 820.050 49.350 ;
        RECT 825.150 48.300 826.950 48.750 ;
        RECT 828.450 48.300 829.500 51.750 ;
        RECT 832.050 51.000 843.900 52.050 ;
        RECT 845.100 50.100 846.300 63.600 ;
        RECT 799.350 46.500 806.100 48.300 ;
        RECT 807.000 46.500 813.900 48.300 ;
        RECT 825.150 47.850 829.500 48.300 ;
        RECT 821.850 47.100 829.500 47.850 ;
        RECT 831.000 49.200 846.300 50.100 ;
        RECT 821.850 46.950 826.950 47.100 ;
        RECT 821.850 45.600 822.750 46.950 ;
        RECT 831.000 46.050 832.050 49.200 ;
        RECT 840.300 47.700 842.100 48.300 ;
        RECT 784.650 39.750 786.450 45.600 ;
        RECT 790.050 39.750 791.850 45.600 ;
        RECT 793.200 44.400 797.400 45.600 ;
        RECT 795.600 39.750 797.400 44.400 ;
        RECT 799.950 43.500 802.050 45.600 ;
        RECT 802.950 43.500 805.050 45.600 ;
        RECT 805.950 43.500 808.050 45.600 ;
        RECT 810.750 45.300 812.850 45.600 ;
        RECT 800.250 39.750 802.050 43.500 ;
        RECT 803.250 39.750 805.050 43.500 ;
        RECT 806.250 39.750 808.050 43.500 ;
        RECT 810.000 43.500 812.850 45.300 ;
        RECT 814.950 45.300 817.050 45.600 ;
        RECT 814.950 43.500 817.800 45.300 ;
        RECT 818.700 44.250 822.750 45.600 ;
        RECT 818.700 43.800 820.500 44.250 ;
        RECT 823.950 43.950 826.050 46.050 ;
        RECT 826.950 43.950 829.050 46.050 ;
        RECT 829.950 43.950 832.050 46.050 ;
        RECT 833.700 46.500 842.100 47.700 ;
        RECT 833.700 45.600 835.200 46.500 ;
        RECT 845.100 45.600 846.300 49.200 ;
        RECT 810.000 39.750 811.800 43.500 ;
        RECT 813.000 39.750 814.800 42.600 ;
        RECT 816.000 39.750 817.800 43.500 ;
        RECT 823.950 42.600 825.300 43.950 ;
        RECT 826.950 42.600 828.300 43.950 ;
        RECT 829.950 42.600 831.300 43.950 ;
        RECT 820.500 39.750 822.300 42.600 ;
        RECT 823.500 39.750 825.300 42.600 ;
        RECT 826.500 39.750 828.300 42.600 ;
        RECT 829.500 39.750 831.300 42.600 ;
        RECT 833.700 39.750 835.500 45.600 ;
        RECT 839.100 39.750 840.900 45.600 ;
        RECT 844.500 39.750 846.300 45.600 ;
        RECT 2.700 29.400 4.500 35.250 ;
        RECT 8.100 29.400 9.900 35.250 ;
        RECT 13.500 29.400 15.300 35.250 ;
        RECT 17.700 32.400 19.500 35.250 ;
        RECT 20.700 32.400 22.500 35.250 ;
        RECT 23.700 32.400 25.500 35.250 ;
        RECT 26.700 32.400 28.500 35.250 ;
        RECT 17.700 31.050 19.050 32.400 ;
        RECT 20.700 31.050 22.050 32.400 ;
        RECT 23.700 31.050 25.050 32.400 ;
        RECT 31.200 31.500 33.000 35.250 ;
        RECT 34.200 32.400 36.000 35.250 ;
        RECT 37.200 31.500 39.000 35.250 ;
        RECT 2.700 25.800 3.900 29.400 ;
        RECT 13.800 28.500 15.300 29.400 ;
        RECT 6.900 27.300 15.300 28.500 ;
        RECT 16.950 28.950 19.050 31.050 ;
        RECT 19.950 28.950 22.050 31.050 ;
        RECT 22.950 28.950 25.050 31.050 ;
        RECT 28.500 30.750 30.300 31.200 ;
        RECT 26.250 29.400 30.300 30.750 ;
        RECT 31.200 29.700 34.050 31.500 ;
        RECT 31.950 29.400 34.050 29.700 ;
        RECT 36.150 29.700 39.000 31.500 ;
        RECT 40.950 31.500 42.750 35.250 ;
        RECT 43.950 31.500 45.750 35.250 ;
        RECT 46.950 31.500 48.750 35.250 ;
        RECT 36.150 29.400 38.250 29.700 ;
        RECT 40.950 29.400 43.050 31.500 ;
        RECT 43.950 29.400 46.050 31.500 ;
        RECT 46.950 29.400 49.050 31.500 ;
        RECT 51.600 30.600 53.400 35.250 ;
        RECT 51.600 29.400 55.800 30.600 ;
        RECT 57.150 29.400 58.950 35.250 ;
        RECT 62.550 29.400 64.350 35.250 ;
        RECT 6.900 26.700 8.700 27.300 ;
        RECT 16.950 25.800 18.000 28.950 ;
        RECT 26.250 28.050 27.150 29.400 ;
        RECT 22.050 27.900 27.150 28.050 ;
        RECT 2.700 24.900 18.000 25.800 ;
        RECT 19.500 27.150 27.150 27.900 ;
        RECT 19.500 26.700 23.850 27.150 ;
        RECT 35.100 26.700 42.000 28.500 ;
        RECT 42.900 26.700 49.650 28.500 ;
        RECT 2.700 11.400 3.900 24.900 ;
        RECT 5.100 22.950 16.950 24.000 ;
        RECT 19.500 23.250 20.550 26.700 ;
        RECT 22.050 26.250 23.850 26.700 ;
        RECT 28.950 25.650 31.050 25.950 ;
        RECT 40.950 25.800 42.000 26.700 ;
        RECT 54.300 25.800 55.800 29.400 ;
        RECT 27.150 23.850 31.050 25.650 ;
        RECT 32.400 24.450 40.050 25.800 ;
        RECT 40.950 24.750 50.850 25.800 ;
        RECT 5.100 21.150 6.900 22.950 ;
        RECT 4.950 19.050 7.050 21.150 ;
        RECT 15.750 20.550 16.950 22.950 ;
        RECT 18.750 21.450 20.550 23.250 ;
        RECT 32.400 22.950 33.450 24.450 ;
        RECT 39.150 23.700 40.050 24.450 ;
        RECT 21.450 22.050 33.450 22.950 ;
        RECT 21.450 20.550 22.500 22.050 ;
        RECT 34.350 21.750 38.250 23.550 ;
        RECT 39.150 22.650 48.750 23.700 ;
        RECT 36.150 21.450 38.250 21.750 ;
        RECT 10.950 19.650 13.050 19.950 ;
        RECT 15.750 19.650 22.500 20.550 ;
        RECT 23.400 20.550 25.200 21.150 ;
        RECT 31.950 20.550 34.050 20.850 ;
        RECT 23.400 19.950 34.050 20.550 ;
        RECT 44.700 19.950 46.500 21.750 ;
        RECT 10.950 18.450 14.850 19.650 ;
        RECT 23.400 19.350 46.500 19.950 ;
        RECT 31.950 18.750 46.500 19.350 ;
        RECT 47.850 21.000 48.750 22.650 ;
        RECT 49.800 22.950 50.850 24.750 ;
        RECT 54.300 24.000 62.100 25.800 ;
        RECT 49.800 21.900 58.050 22.950 ;
        RECT 47.850 19.200 54.900 21.000 ;
        RECT 10.950 17.850 24.900 18.450 ;
        RECT 55.950 17.850 58.050 21.900 ;
        RECT 11.250 17.550 51.000 17.850 ;
        RECT 22.950 16.650 51.000 17.550 ;
        RECT 60.450 16.650 62.250 17.250 ;
        RECT 10.500 16.050 12.300 16.650 ;
        RECT 19.950 16.050 22.050 16.350 ;
        RECT 10.500 14.850 22.050 16.050 ;
        RECT 19.950 14.250 22.050 14.850 ;
        RECT 22.950 14.400 43.050 15.750 ;
        RECT 7.200 13.350 9.000 14.100 ;
        RECT 22.950 13.350 24.900 14.400 ;
        RECT 40.950 13.650 43.050 14.400 ;
        RECT 46.950 14.550 49.050 15.750 ;
        RECT 49.950 15.450 62.250 16.650 ;
        RECT 63.150 14.550 64.350 29.400 ;
        RECT 46.950 13.650 64.350 14.550 ;
        RECT 66.450 32.400 68.250 35.250 ;
        RECT 69.450 32.400 71.250 35.250 ;
        RECT 66.450 24.150 67.950 32.400 ;
        RECT 74.550 29.400 76.350 35.250 ;
        RECT 77.550 29.400 79.350 35.250 ;
        RECT 89.850 29.400 91.650 35.250 ;
        RECT 74.100 24.150 75.900 25.950 ;
        RECT 66.450 22.050 70.050 24.150 ;
        RECT 73.950 22.050 76.050 24.150 ;
        RECT 77.400 22.950 78.600 29.400 ;
        RECT 94.350 28.200 96.150 35.250 ;
        RECT 103.650 29.400 105.450 35.250 ;
        RECT 92.550 27.300 96.150 28.200 ;
        RECT 104.250 27.300 105.450 29.400 ;
        RECT 106.650 30.300 108.450 35.250 ;
        RECT 109.650 31.200 111.450 35.250 ;
        RECT 112.650 30.300 114.450 35.250 ;
        RECT 106.650 28.950 114.450 30.300 ;
        RECT 116.550 30.300 118.350 35.250 ;
        RECT 119.550 31.200 121.350 35.250 ;
        RECT 122.550 30.300 124.350 35.250 ;
        RECT 116.550 28.950 124.350 30.300 ;
        RECT 125.550 29.400 127.350 35.250 ;
        RECT 137.550 30.300 139.350 35.250 ;
        RECT 140.550 31.200 142.350 35.250 ;
        RECT 143.550 30.300 145.350 35.250 ;
        RECT 125.550 27.300 126.750 29.400 ;
        RECT 137.550 28.950 145.350 30.300 ;
        RECT 146.550 29.400 148.350 35.250 ;
        RECT 160.650 32.400 162.450 35.250 ;
        RECT 163.650 32.400 165.450 35.250 ;
        RECT 173.550 32.400 175.350 35.250 ;
        RECT 176.550 32.400 178.350 35.250 ;
        RECT 146.550 27.300 147.750 29.400 ;
        RECT 7.200 12.300 24.900 13.350 ;
        RECT 2.700 10.500 6.750 11.400 ;
        RECT 5.700 9.600 6.750 10.500 ;
        RECT 2.700 3.750 4.500 9.600 ;
        RECT 5.700 3.750 7.500 9.600 ;
        RECT 8.700 3.750 10.500 9.600 ;
        RECT 11.700 3.750 13.500 12.300 ;
        RECT 31.950 12.150 34.050 12.600 ;
        RECT 31.650 10.500 34.050 12.150 ;
        RECT 36.000 10.800 39.900 12.600 ;
        RECT 36.000 10.500 39.000 10.800 ;
        RECT 16.950 7.950 19.050 10.050 ;
        RECT 19.950 7.950 22.050 10.050 ;
        RECT 22.950 9.600 25.050 10.050 ;
        RECT 31.650 9.600 33.000 10.500 ;
        RECT 22.950 7.950 25.500 9.600 ;
        RECT 14.700 3.750 16.500 7.050 ;
        RECT 17.850 6.600 19.050 7.950 ;
        RECT 21.150 6.600 22.050 7.950 ;
        RECT 24.300 6.600 25.500 7.950 ;
        RECT 17.850 3.750 20.250 6.600 ;
        RECT 21.150 3.750 23.250 6.600 ;
        RECT 24.300 3.750 26.250 6.600 ;
        RECT 27.450 3.750 29.250 9.600 ;
        RECT 31.200 3.750 33.000 9.600 ;
        RECT 34.200 3.750 36.000 9.600 ;
        RECT 37.200 3.750 39.000 10.500 ;
        RECT 41.100 6.600 42.450 13.650 ;
        RECT 50.850 12.150 52.650 12.300 ;
        RECT 43.950 10.950 52.650 12.150 ;
        RECT 57.600 11.700 59.400 12.300 ;
        RECT 43.950 10.050 46.050 10.950 ;
        RECT 50.850 10.500 52.650 10.950 ;
        RECT 53.700 10.500 59.400 11.700 ;
        RECT 40.950 3.750 42.750 6.600 ;
        RECT 43.950 3.750 45.750 10.050 ;
        RECT 47.100 7.800 49.200 9.900 ;
        RECT 47.100 6.600 48.600 7.800 ;
        RECT 46.950 3.750 48.750 6.600 ;
        RECT 50.700 3.750 52.500 9.600 ;
        RECT 53.700 3.750 55.500 10.500 ;
        RECT 60.300 9.600 61.500 13.650 ;
        RECT 66.450 9.600 67.950 22.050 ;
        RECT 76.950 20.850 79.050 22.950 ;
        RECT 89.100 21.150 90.900 22.950 ;
        RECT 77.400 15.600 78.600 20.850 ;
        RECT 88.950 19.050 91.050 21.150 ;
        RECT 92.550 19.950 93.750 27.300 ;
        RECT 104.250 26.250 108.000 27.300 ;
        RECT 123.000 26.250 126.750 27.300 ;
        RECT 144.000 26.250 147.750 27.300 ;
        RECT 106.950 22.950 108.150 26.250 ;
        RECT 110.100 24.150 111.900 25.950 ;
        RECT 119.100 24.150 120.900 25.950 ;
        RECT 95.100 21.150 96.900 22.950 ;
        RECT 91.950 17.850 94.050 19.950 ;
        RECT 94.950 19.050 97.050 21.150 ;
        RECT 106.950 20.850 109.050 22.950 ;
        RECT 109.950 22.050 112.050 24.150 ;
        RECT 112.950 20.850 115.050 22.950 ;
        RECT 115.950 20.850 118.050 22.950 ;
        RECT 118.950 22.050 121.050 24.150 ;
        RECT 122.850 22.950 124.050 26.250 ;
        RECT 124.950 24.450 127.050 25.050 ;
        RECT 130.950 24.450 133.050 25.050 ;
        RECT 124.950 23.550 133.050 24.450 ;
        RECT 140.100 24.150 141.900 25.950 ;
        RECT 124.950 22.950 127.050 23.550 ;
        RECT 130.950 22.950 133.050 23.550 ;
        RECT 121.950 20.850 124.050 22.950 ;
        RECT 136.950 20.850 139.050 22.950 ;
        RECT 139.950 22.050 142.050 24.150 ;
        RECT 143.850 22.950 145.050 26.250 ;
        RECT 161.400 24.150 162.600 32.400 ;
        RECT 142.950 20.850 145.050 22.950 ;
        RECT 160.950 22.050 163.050 24.150 ;
        RECT 163.950 23.850 166.050 25.950 ;
        RECT 172.950 23.850 175.050 25.950 ;
        RECT 176.400 24.150 177.600 32.400 ;
        RECT 182.700 29.400 184.500 35.250 ;
        RECT 188.100 29.400 189.900 35.250 ;
        RECT 193.500 29.400 195.300 35.250 ;
        RECT 197.700 32.400 199.500 35.250 ;
        RECT 200.700 32.400 202.500 35.250 ;
        RECT 203.700 32.400 205.500 35.250 ;
        RECT 206.700 32.400 208.500 35.250 ;
        RECT 197.700 31.050 199.050 32.400 ;
        RECT 200.700 31.050 202.050 32.400 ;
        RECT 203.700 31.050 205.050 32.400 ;
        RECT 211.200 31.500 213.000 35.250 ;
        RECT 214.200 32.400 216.000 35.250 ;
        RECT 217.200 31.500 219.000 35.250 ;
        RECT 182.700 25.800 183.900 29.400 ;
        RECT 193.800 28.500 195.300 29.400 ;
        RECT 186.900 27.300 195.300 28.500 ;
        RECT 196.950 28.950 199.050 31.050 ;
        RECT 199.950 28.950 202.050 31.050 ;
        RECT 202.950 28.950 205.050 31.050 ;
        RECT 208.500 30.750 210.300 31.200 ;
        RECT 206.250 29.400 210.300 30.750 ;
        RECT 211.200 29.700 214.050 31.500 ;
        RECT 211.950 29.400 214.050 29.700 ;
        RECT 216.150 29.700 219.000 31.500 ;
        RECT 220.950 31.500 222.750 35.250 ;
        RECT 223.950 31.500 225.750 35.250 ;
        RECT 226.950 31.500 228.750 35.250 ;
        RECT 216.150 29.400 218.250 29.700 ;
        RECT 220.950 29.400 223.050 31.500 ;
        RECT 223.950 29.400 226.050 31.500 ;
        RECT 226.950 29.400 229.050 31.500 ;
        RECT 231.600 30.600 233.400 35.250 ;
        RECT 231.600 29.400 235.800 30.600 ;
        RECT 237.150 29.400 238.950 35.250 ;
        RECT 242.550 29.400 244.350 35.250 ;
        RECT 186.900 26.700 188.700 27.300 ;
        RECT 196.950 25.800 198.000 28.950 ;
        RECT 206.250 28.050 207.150 29.400 ;
        RECT 202.050 27.900 207.150 28.050 ;
        RECT 182.700 24.900 198.000 25.800 ;
        RECT 199.500 27.150 207.150 27.900 ;
        RECT 199.500 26.700 203.850 27.150 ;
        RECT 215.100 26.700 222.000 28.500 ;
        RECT 222.900 26.700 229.650 28.500 ;
        RECT 164.100 22.050 165.900 23.850 ;
        RECT 173.100 22.050 174.900 23.850 ;
        RECT 175.950 22.050 178.050 24.150 ;
        RECT 103.950 17.850 106.050 19.950 ;
        RECT 56.700 3.750 58.500 9.600 ;
        RECT 59.700 3.750 61.500 9.600 ;
        RECT 62.700 3.750 64.500 9.600 ;
        RECT 66.450 3.750 68.250 9.600 ;
        RECT 69.450 3.750 71.250 9.600 ;
        RECT 74.550 3.750 76.350 15.600 ;
        RECT 77.550 3.750 79.350 15.600 ;
        RECT 92.550 9.600 93.750 17.850 ;
        RECT 104.250 16.050 106.050 17.850 ;
        RECT 107.850 15.600 109.050 20.850 ;
        RECT 113.100 19.050 114.900 20.850 ;
        RECT 116.100 19.050 117.900 20.850 ;
        RECT 121.950 15.600 123.150 20.850 ;
        RECT 124.950 17.850 127.050 19.950 ;
        RECT 137.100 19.050 138.900 20.850 ;
        RECT 124.950 16.050 126.750 17.850 ;
        RECT 142.950 15.600 144.150 20.850 ;
        RECT 145.950 17.850 148.050 19.950 ;
        RECT 145.950 16.050 147.750 17.850 ;
        RECT 89.550 3.750 91.350 9.600 ;
        RECT 92.550 3.750 94.350 9.600 ;
        RECT 95.550 3.750 97.350 9.600 ;
        RECT 104.400 3.750 106.200 9.600 ;
        RECT 107.700 3.750 109.500 15.600 ;
        RECT 111.900 3.750 113.700 15.600 ;
        RECT 117.300 3.750 119.100 15.600 ;
        RECT 121.500 3.750 123.300 15.600 ;
        RECT 124.800 3.750 126.600 9.600 ;
        RECT 138.300 3.750 140.100 15.600 ;
        RECT 142.500 3.750 144.300 15.600 ;
        RECT 161.400 9.600 162.600 22.050 ;
        RECT 176.400 9.600 177.600 22.050 ;
        RECT 182.700 11.400 183.900 24.900 ;
        RECT 185.100 22.950 196.950 24.000 ;
        RECT 199.500 23.250 200.550 26.700 ;
        RECT 202.050 26.250 203.850 26.700 ;
        RECT 208.950 25.650 211.050 25.950 ;
        RECT 220.950 25.800 222.000 26.700 ;
        RECT 234.300 25.800 235.800 29.400 ;
        RECT 207.150 23.850 211.050 25.650 ;
        RECT 212.400 24.450 220.050 25.800 ;
        RECT 220.950 24.750 230.850 25.800 ;
        RECT 185.100 21.150 186.900 22.950 ;
        RECT 184.950 19.050 187.050 21.150 ;
        RECT 195.750 20.550 196.950 22.950 ;
        RECT 198.750 21.450 200.550 23.250 ;
        RECT 212.400 22.950 213.450 24.450 ;
        RECT 219.150 23.700 220.050 24.450 ;
        RECT 201.450 22.050 213.450 22.950 ;
        RECT 201.450 20.550 202.500 22.050 ;
        RECT 214.350 21.750 218.250 23.550 ;
        RECT 219.150 22.650 228.750 23.700 ;
        RECT 216.150 21.450 218.250 21.750 ;
        RECT 190.950 19.650 193.050 19.950 ;
        RECT 195.750 19.650 202.500 20.550 ;
        RECT 203.400 20.550 205.200 21.150 ;
        RECT 211.950 20.550 214.050 20.850 ;
        RECT 203.400 19.950 214.050 20.550 ;
        RECT 224.700 19.950 226.500 21.750 ;
        RECT 190.950 18.450 194.850 19.650 ;
        RECT 203.400 19.350 226.500 19.950 ;
        RECT 211.950 18.750 226.500 19.350 ;
        RECT 227.850 21.000 228.750 22.650 ;
        RECT 229.800 22.950 230.850 24.750 ;
        RECT 234.300 24.000 242.100 25.800 ;
        RECT 229.800 21.900 238.050 22.950 ;
        RECT 227.850 19.200 234.900 21.000 ;
        RECT 190.950 17.850 204.900 18.450 ;
        RECT 235.950 17.850 238.050 21.900 ;
        RECT 191.250 17.550 231.000 17.850 ;
        RECT 202.950 16.650 231.000 17.550 ;
        RECT 240.450 16.650 242.250 17.250 ;
        RECT 190.500 16.050 192.300 16.650 ;
        RECT 199.950 16.050 202.050 16.350 ;
        RECT 190.500 14.850 202.050 16.050 ;
        RECT 199.950 14.250 202.050 14.850 ;
        RECT 202.950 14.400 223.050 15.750 ;
        RECT 187.200 13.350 189.000 14.100 ;
        RECT 202.950 13.350 204.900 14.400 ;
        RECT 220.950 13.650 223.050 14.400 ;
        RECT 226.950 14.550 229.050 15.750 ;
        RECT 229.950 15.450 242.250 16.650 ;
        RECT 243.150 14.550 244.350 29.400 ;
        RECT 226.950 13.650 244.350 14.550 ;
        RECT 246.450 32.400 248.250 35.250 ;
        RECT 249.450 32.400 251.250 35.250 ;
        RECT 246.450 24.150 247.950 32.400 ;
        RECT 257.550 30.300 259.350 35.250 ;
        RECT 260.550 31.200 262.350 35.250 ;
        RECT 263.550 30.300 265.350 35.250 ;
        RECT 257.550 28.950 265.350 30.300 ;
        RECT 266.550 29.400 268.350 35.250 ;
        RECT 266.550 27.300 267.750 29.400 ;
        RECT 278.850 28.200 280.650 35.250 ;
        RECT 283.350 29.400 285.150 35.250 ;
        RECT 292.650 32.400 294.450 35.250 ;
        RECT 295.650 32.400 297.450 35.250 ;
        RECT 298.650 32.400 300.450 35.250 ;
        RECT 278.850 27.300 282.450 28.200 ;
        RECT 264.000 26.250 267.750 27.300 ;
        RECT 260.100 24.150 261.900 25.950 ;
        RECT 246.450 22.050 250.050 24.150 ;
        RECT 187.200 12.300 204.900 13.350 ;
        RECT 182.700 10.500 186.750 11.400 ;
        RECT 185.700 9.600 186.750 10.500 ;
        RECT 145.800 3.750 147.600 9.600 ;
        RECT 160.650 3.750 162.450 9.600 ;
        RECT 163.650 3.750 165.450 9.600 ;
        RECT 173.550 3.750 175.350 9.600 ;
        RECT 176.550 3.750 178.350 9.600 ;
        RECT 182.700 3.750 184.500 9.600 ;
        RECT 185.700 3.750 187.500 9.600 ;
        RECT 188.700 3.750 190.500 9.600 ;
        RECT 191.700 3.750 193.500 12.300 ;
        RECT 211.950 12.150 214.050 12.600 ;
        RECT 211.650 10.500 214.050 12.150 ;
        RECT 216.000 10.800 219.900 12.600 ;
        RECT 216.000 10.500 219.000 10.800 ;
        RECT 196.950 7.950 199.050 10.050 ;
        RECT 199.950 7.950 202.050 10.050 ;
        RECT 202.950 9.600 205.050 10.050 ;
        RECT 211.650 9.600 213.000 10.500 ;
        RECT 202.950 7.950 205.500 9.600 ;
        RECT 194.700 3.750 196.500 7.050 ;
        RECT 197.850 6.600 199.050 7.950 ;
        RECT 201.150 6.600 202.050 7.950 ;
        RECT 204.300 6.600 205.500 7.950 ;
        RECT 197.850 3.750 200.250 6.600 ;
        RECT 201.150 3.750 203.250 6.600 ;
        RECT 204.300 3.750 206.250 6.600 ;
        RECT 207.450 3.750 209.250 9.600 ;
        RECT 211.200 3.750 213.000 9.600 ;
        RECT 214.200 3.750 216.000 9.600 ;
        RECT 217.200 3.750 219.000 10.500 ;
        RECT 221.100 6.600 222.450 13.650 ;
        RECT 230.850 12.150 232.650 12.300 ;
        RECT 223.950 10.950 232.650 12.150 ;
        RECT 237.600 11.700 239.400 12.300 ;
        RECT 223.950 10.050 226.050 10.950 ;
        RECT 230.850 10.500 232.650 10.950 ;
        RECT 233.700 10.500 239.400 11.700 ;
        RECT 220.950 3.750 222.750 6.600 ;
        RECT 223.950 3.750 225.750 10.050 ;
        RECT 227.100 7.800 229.200 9.900 ;
        RECT 227.100 6.600 228.600 7.800 ;
        RECT 226.950 3.750 228.750 6.600 ;
        RECT 230.700 3.750 232.500 9.600 ;
        RECT 233.700 3.750 235.500 10.500 ;
        RECT 240.300 9.600 241.500 13.650 ;
        RECT 246.450 9.600 247.950 22.050 ;
        RECT 256.950 20.850 259.050 22.950 ;
        RECT 259.950 22.050 262.050 24.150 ;
        RECT 263.850 22.950 265.050 26.250 ;
        RECT 262.950 20.850 265.050 22.950 ;
        RECT 278.100 21.150 279.900 22.950 ;
        RECT 257.100 19.050 258.900 20.850 ;
        RECT 262.950 15.600 264.150 20.850 ;
        RECT 265.950 17.850 268.050 19.950 ;
        RECT 277.950 19.050 280.050 21.150 ;
        RECT 281.250 19.950 282.450 27.300 ;
        RECT 295.950 25.950 297.000 32.400 ;
        RECT 305.550 30.300 307.350 35.250 ;
        RECT 308.550 31.200 310.350 35.250 ;
        RECT 311.550 30.300 313.350 35.250 ;
        RECT 305.550 28.950 313.350 30.300 ;
        RECT 314.550 29.400 316.350 35.250 ;
        RECT 325.650 29.400 327.450 35.250 ;
        RECT 314.550 27.300 315.750 29.400 ;
        RECT 312.000 26.250 315.750 27.300 ;
        RECT 326.250 27.300 327.450 29.400 ;
        RECT 328.650 30.300 330.450 35.250 ;
        RECT 331.650 31.200 333.450 35.250 ;
        RECT 334.650 30.300 336.450 35.250 ;
        RECT 328.650 28.950 336.450 30.300 ;
        RECT 344.850 28.200 346.650 35.250 ;
        RECT 349.350 29.400 351.150 35.250 ;
        RECT 359.550 32.400 361.350 35.250 ;
        RECT 362.550 32.400 364.350 35.250 ;
        RECT 365.550 32.400 367.350 35.250 ;
        RECT 344.850 27.300 348.450 28.200 ;
        RECT 326.250 26.250 330.000 27.300 ;
        RECT 295.950 23.850 298.050 25.950 ;
        RECT 308.100 24.150 309.900 25.950 ;
        RECT 284.100 21.150 285.900 22.950 ;
        RECT 280.950 17.850 283.050 19.950 ;
        RECT 283.950 19.050 286.050 21.150 ;
        RECT 292.950 20.850 295.050 22.950 ;
        RECT 293.100 19.050 294.900 20.850 ;
        RECT 265.950 16.050 267.750 17.850 ;
        RECT 236.700 3.750 238.500 9.600 ;
        RECT 239.700 3.750 241.500 9.600 ;
        RECT 242.700 3.750 244.500 9.600 ;
        RECT 246.450 3.750 248.250 9.600 ;
        RECT 249.450 3.750 251.250 9.600 ;
        RECT 258.300 3.750 260.100 15.600 ;
        RECT 262.500 3.750 264.300 15.600 ;
        RECT 281.250 9.600 282.450 17.850 ;
        RECT 295.950 16.650 297.000 23.850 ;
        RECT 298.950 20.850 301.050 22.950 ;
        RECT 304.950 20.850 307.050 22.950 ;
        RECT 307.950 22.050 310.050 24.150 ;
        RECT 311.850 22.950 313.050 26.250 ;
        RECT 310.950 20.850 313.050 22.950 ;
        RECT 328.950 22.950 330.150 26.250 ;
        RECT 332.100 24.150 333.900 25.950 ;
        RECT 328.950 20.850 331.050 22.950 ;
        RECT 331.950 22.050 334.050 24.150 ;
        RECT 334.950 20.850 337.050 22.950 ;
        RECT 344.100 21.150 345.900 22.950 ;
        RECT 299.100 19.050 300.900 20.850 ;
        RECT 305.100 19.050 306.900 20.850 ;
        RECT 294.450 15.600 297.000 16.650 ;
        RECT 310.950 15.600 312.150 20.850 ;
        RECT 313.950 17.850 316.050 19.950 ;
        RECT 325.950 17.850 328.050 19.950 ;
        RECT 313.950 16.050 315.750 17.850 ;
        RECT 326.250 16.050 328.050 17.850 ;
        RECT 329.850 15.600 331.050 20.850 ;
        RECT 335.100 19.050 336.900 20.850 ;
        RECT 343.950 19.050 346.050 21.150 ;
        RECT 347.250 19.950 348.450 27.300 ;
        RECT 363.000 25.950 364.050 32.400 ;
        RECT 375.000 29.400 376.800 35.250 ;
        RECT 379.200 31.050 381.000 35.250 ;
        RECT 382.500 32.400 384.300 35.250 ;
        RECT 379.200 29.400 384.900 31.050 ;
        RECT 389.550 29.400 391.350 35.250 ;
        RECT 392.550 29.400 394.350 35.250 ;
        RECT 401.550 30.300 403.350 35.250 ;
        RECT 404.550 31.200 406.350 35.250 ;
        RECT 407.550 30.300 409.350 35.250 ;
        RECT 361.950 23.850 364.050 25.950 ;
        RECT 374.100 24.150 375.900 25.950 ;
        RECT 350.100 21.150 351.900 22.950 ;
        RECT 346.950 17.850 349.050 19.950 ;
        RECT 349.950 19.050 352.050 21.150 ;
        RECT 358.950 20.850 361.050 22.950 ;
        RECT 359.100 19.050 360.900 20.850 ;
        RECT 265.800 3.750 267.600 9.600 ;
        RECT 277.650 3.750 279.450 9.600 ;
        RECT 280.650 3.750 282.450 9.600 ;
        RECT 283.650 3.750 285.450 9.600 ;
        RECT 294.450 3.750 296.250 15.600 ;
        RECT 298.650 3.750 300.450 15.600 ;
        RECT 306.300 3.750 308.100 15.600 ;
        RECT 310.500 3.750 312.300 15.600 ;
        RECT 313.800 3.750 315.600 9.600 ;
        RECT 326.400 3.750 328.200 9.600 ;
        RECT 329.700 3.750 331.500 15.600 ;
        RECT 333.900 3.750 335.700 15.600 ;
        RECT 347.250 9.600 348.450 17.850 ;
        RECT 363.000 16.650 364.050 23.850 ;
        RECT 364.950 20.850 367.050 22.950 ;
        RECT 373.950 22.050 376.050 24.150 ;
        RECT 376.950 23.850 379.050 25.950 ;
        RECT 380.100 24.150 381.900 25.950 ;
        RECT 377.100 22.050 378.900 23.850 ;
        RECT 379.950 22.050 382.050 24.150 ;
        RECT 383.700 22.950 384.900 29.400 ;
        RECT 389.100 24.150 390.900 25.950 ;
        RECT 382.950 20.850 385.050 22.950 ;
        RECT 388.950 22.050 391.050 24.150 ;
        RECT 392.400 22.950 393.600 29.400 ;
        RECT 401.550 28.950 409.350 30.300 ;
        RECT 410.550 29.400 412.350 35.250 ;
        RECT 410.550 27.300 411.750 29.400 ;
        RECT 422.850 28.200 424.650 35.250 ;
        RECT 427.350 29.400 429.150 35.250 ;
        RECT 436.650 32.400 438.450 35.250 ;
        RECT 439.650 32.400 441.450 35.250 ;
        RECT 442.650 32.400 444.450 35.250 ;
        RECT 422.850 27.300 426.450 28.200 ;
        RECT 408.000 26.250 411.750 27.300 ;
        RECT 404.100 24.150 405.900 25.950 ;
        RECT 391.950 20.850 394.050 22.950 ;
        RECT 400.950 20.850 403.050 22.950 ;
        RECT 403.950 22.050 406.050 24.150 ;
        RECT 407.850 22.950 409.050 26.250 ;
        RECT 406.950 20.850 409.050 22.950 ;
        RECT 422.100 21.150 423.900 22.950 ;
        RECT 365.100 19.050 366.900 20.850 ;
        RECT 363.000 15.600 365.550 16.650 ;
        RECT 383.700 15.600 384.900 20.850 ;
        RECT 392.400 15.600 393.600 20.850 ;
        RECT 401.100 19.050 402.900 20.850 ;
        RECT 406.950 15.600 408.150 20.850 ;
        RECT 409.950 17.850 412.050 19.950 ;
        RECT 421.950 19.050 424.050 21.150 ;
        RECT 425.250 19.950 426.450 27.300 ;
        RECT 439.950 25.950 441.000 32.400 ;
        RECT 454.800 29.400 456.600 35.250 ;
        RECT 459.000 29.400 460.800 35.250 ;
        RECT 463.200 29.400 465.000 35.250 ;
        RECT 470.850 29.400 472.650 35.250 ;
        RECT 439.950 23.850 442.050 25.950 ;
        RECT 455.250 24.150 457.050 25.950 ;
        RECT 428.100 21.150 429.900 22.950 ;
        RECT 424.950 17.850 427.050 19.950 ;
        RECT 427.950 19.050 430.050 21.150 ;
        RECT 436.950 20.850 439.050 22.950 ;
        RECT 437.100 19.050 438.900 20.850 ;
        RECT 409.950 16.050 411.750 17.850 ;
        RECT 343.650 3.750 345.450 9.600 ;
        RECT 346.650 3.750 348.450 9.600 ;
        RECT 349.650 3.750 351.450 9.600 ;
        RECT 359.550 3.750 361.350 15.600 ;
        RECT 363.750 3.750 365.550 15.600 ;
        RECT 374.550 14.700 382.350 15.600 ;
        RECT 374.550 3.750 376.350 14.700 ;
        RECT 377.550 3.750 379.350 13.800 ;
        RECT 380.550 3.750 382.350 14.700 ;
        RECT 383.550 3.750 385.350 15.600 ;
        RECT 389.550 3.750 391.350 15.600 ;
        RECT 392.550 3.750 394.350 15.600 ;
        RECT 402.300 3.750 404.100 15.600 ;
        RECT 406.500 3.750 408.300 15.600 ;
        RECT 425.250 9.600 426.450 17.850 ;
        RECT 439.950 16.650 441.000 23.850 ;
        RECT 442.950 20.850 445.050 22.950 ;
        RECT 451.950 20.850 454.050 22.950 ;
        RECT 454.950 22.050 457.050 24.150 ;
        RECT 459.000 22.950 460.050 29.400 ;
        RECT 475.350 28.200 477.150 35.250 ;
        RECT 485.550 32.400 487.350 35.250 ;
        RECT 488.550 32.400 490.350 35.250 ;
        RECT 473.550 27.300 477.150 28.200 ;
        RECT 457.950 20.850 460.050 22.950 ;
        RECT 460.950 24.150 462.750 25.950 ;
        RECT 460.950 22.050 463.050 24.150 ;
        RECT 463.950 20.850 466.050 22.950 ;
        RECT 470.100 21.150 471.900 22.950 ;
        RECT 443.100 19.050 444.900 20.850 ;
        RECT 452.100 19.050 453.900 20.850 ;
        RECT 457.950 17.400 458.850 20.850 ;
        RECT 463.950 19.050 465.750 20.850 ;
        RECT 469.950 19.050 472.050 21.150 ;
        RECT 473.550 19.950 474.750 27.300 ;
        RECT 484.950 23.850 487.050 25.950 ;
        RECT 488.400 24.150 489.600 32.400 ;
        RECT 497.550 30.300 499.350 35.250 ;
        RECT 500.550 31.200 502.350 35.250 ;
        RECT 503.550 30.300 505.350 35.250 ;
        RECT 497.550 28.950 505.350 30.300 ;
        RECT 506.550 29.400 508.350 35.250 ;
        RECT 512.550 32.400 514.350 35.250 ;
        RECT 515.550 32.400 517.350 35.250 ;
        RECT 518.550 32.400 520.350 35.250 ;
        RECT 506.550 27.300 507.750 29.400 ;
        RECT 504.000 26.250 507.750 27.300 ;
        RECT 500.100 24.150 501.900 25.950 ;
        RECT 476.100 21.150 477.900 22.950 ;
        RECT 485.100 22.050 486.900 23.850 ;
        RECT 487.950 22.050 490.050 24.150 ;
        RECT 472.950 17.850 475.050 19.950 ;
        RECT 475.950 19.050 478.050 21.150 ;
        RECT 438.450 15.600 441.000 16.650 ;
        RECT 454.800 16.500 458.850 17.400 ;
        RECT 454.800 15.600 456.600 16.500 ;
        RECT 409.800 3.750 411.600 9.600 ;
        RECT 421.650 3.750 423.450 9.600 ;
        RECT 424.650 3.750 426.450 9.600 ;
        RECT 427.650 3.750 429.450 9.600 ;
        RECT 438.450 3.750 440.250 15.600 ;
        RECT 442.650 3.750 444.450 15.600 ;
        RECT 451.650 4.500 453.450 15.600 ;
        RECT 454.650 5.400 456.450 15.600 ;
        RECT 457.650 14.400 465.450 15.300 ;
        RECT 457.650 4.500 459.450 14.400 ;
        RECT 451.650 3.750 459.450 4.500 ;
        RECT 460.650 3.750 462.450 13.500 ;
        RECT 463.650 3.750 465.450 14.400 ;
        RECT 473.550 9.600 474.750 17.850 ;
        RECT 488.400 9.600 489.600 22.050 ;
        RECT 496.950 20.850 499.050 22.950 ;
        RECT 499.950 22.050 502.050 24.150 ;
        RECT 503.850 22.950 505.050 26.250 ;
        RECT 516.000 25.950 517.050 32.400 ;
        RECT 530.850 28.200 532.650 35.250 ;
        RECT 535.350 29.400 537.150 35.250 ;
        RECT 530.850 27.300 534.450 28.200 ;
        RECT 514.950 23.850 517.050 25.950 ;
        RECT 502.950 20.850 505.050 22.950 ;
        RECT 511.950 20.850 514.050 22.950 ;
        RECT 497.100 19.050 498.900 20.850 ;
        RECT 502.950 15.600 504.150 20.850 ;
        RECT 505.950 17.850 508.050 19.950 ;
        RECT 512.100 19.050 513.900 20.850 ;
        RECT 505.950 16.050 507.750 17.850 ;
        RECT 516.000 16.650 517.050 23.850 ;
        RECT 517.950 20.850 520.050 22.950 ;
        RECT 530.100 21.150 531.900 22.950 ;
        RECT 518.100 19.050 519.900 20.850 ;
        RECT 529.950 19.050 532.050 21.150 ;
        RECT 533.250 19.950 534.450 27.300 ;
        RECT 542.700 26.400 544.500 35.250 ;
        RECT 548.100 27.000 549.900 35.250 ;
        RECT 563.850 28.200 565.650 35.250 ;
        RECT 568.350 29.400 570.150 35.250 ;
        RECT 575.850 29.400 577.650 35.250 ;
        RECT 580.350 28.200 582.150 35.250 ;
        RECT 588.750 32.400 590.550 35.250 ;
        RECT 591.750 32.400 593.550 35.250 ;
        RECT 563.850 27.300 567.450 28.200 ;
        RECT 548.100 25.350 552.600 27.000 ;
        RECT 536.100 21.150 537.900 22.950 ;
        RECT 551.400 21.150 552.600 25.350 ;
        RECT 563.100 21.150 564.900 22.950 ;
        RECT 532.950 17.850 535.050 19.950 ;
        RECT 535.950 19.050 538.050 21.150 ;
        RECT 541.950 17.850 544.050 19.950 ;
        RECT 547.950 17.850 550.050 19.950 ;
        RECT 550.950 19.050 553.050 21.150 ;
        RECT 562.950 19.050 565.050 21.150 ;
        RECT 566.250 19.950 567.450 27.300 ;
        RECT 578.550 27.300 582.150 28.200 ;
        RECT 569.100 21.150 570.900 22.950 ;
        RECT 575.100 21.150 576.900 22.950 ;
        RECT 516.000 15.600 518.550 16.650 ;
        RECT 470.550 3.750 472.350 9.600 ;
        RECT 473.550 3.750 475.350 9.600 ;
        RECT 476.550 3.750 478.350 9.600 ;
        RECT 485.550 3.750 487.350 9.600 ;
        RECT 488.550 3.750 490.350 9.600 ;
        RECT 498.300 3.750 500.100 15.600 ;
        RECT 502.500 3.750 504.300 15.600 ;
        RECT 505.800 3.750 507.600 9.600 ;
        RECT 512.550 3.750 514.350 15.600 ;
        RECT 516.750 3.750 518.550 15.600 ;
        RECT 533.250 9.600 534.450 17.850 ;
        RECT 542.100 16.050 543.900 17.850 ;
        RECT 544.950 14.850 547.050 16.950 ;
        RECT 548.250 16.050 550.050 17.850 ;
        RECT 545.100 13.050 546.900 14.850 ;
        RECT 551.700 10.800 552.750 19.050 ;
        RECT 565.950 17.850 568.050 19.950 ;
        RECT 568.950 19.050 571.050 21.150 ;
        RECT 574.950 19.050 577.050 21.150 ;
        RECT 578.550 19.950 579.750 27.300 ;
        RECT 592.050 24.150 593.550 32.400 ;
        RECT 581.100 21.150 582.900 22.950 ;
        RECT 589.950 22.050 593.550 24.150 ;
        RECT 577.950 17.850 580.050 19.950 ;
        RECT 580.950 19.050 583.050 21.150 ;
        RECT 545.700 9.900 552.750 10.800 ;
        RECT 545.700 9.600 547.350 9.900 ;
        RECT 529.650 3.750 531.450 9.600 ;
        RECT 532.650 3.750 534.450 9.600 ;
        RECT 535.650 3.750 537.450 9.600 ;
        RECT 542.550 3.750 544.350 9.600 ;
        RECT 545.550 3.750 547.350 9.600 ;
        RECT 551.550 9.600 552.750 9.900 ;
        RECT 566.250 9.600 567.450 17.850 ;
        RECT 578.550 9.600 579.750 17.850 ;
        RECT 592.050 9.600 593.550 22.050 ;
        RECT 595.650 29.400 597.450 35.250 ;
        RECT 601.050 29.400 602.850 35.250 ;
        RECT 606.600 30.600 608.400 35.250 ;
        RECT 611.250 31.500 613.050 35.250 ;
        RECT 614.250 31.500 616.050 35.250 ;
        RECT 617.250 31.500 619.050 35.250 ;
        RECT 604.200 29.400 608.400 30.600 ;
        RECT 610.950 29.400 613.050 31.500 ;
        RECT 613.950 29.400 616.050 31.500 ;
        RECT 616.950 29.400 619.050 31.500 ;
        RECT 621.000 31.500 622.800 35.250 ;
        RECT 624.000 32.400 625.800 35.250 ;
        RECT 627.000 31.500 628.800 35.250 ;
        RECT 631.500 32.400 633.300 35.250 ;
        RECT 634.500 32.400 636.300 35.250 ;
        RECT 637.500 32.400 639.300 35.250 ;
        RECT 640.500 32.400 642.300 35.250 ;
        RECT 621.000 29.700 623.850 31.500 ;
        RECT 621.750 29.400 623.850 29.700 ;
        RECT 625.950 29.700 628.800 31.500 ;
        RECT 629.700 30.750 631.500 31.200 ;
        RECT 634.950 31.050 636.300 32.400 ;
        RECT 637.950 31.050 639.300 32.400 ;
        RECT 640.950 31.050 642.300 32.400 ;
        RECT 625.950 29.400 628.050 29.700 ;
        RECT 629.700 29.400 633.750 30.750 ;
        RECT 595.650 14.550 596.850 29.400 ;
        RECT 604.200 25.800 605.700 29.400 ;
        RECT 610.350 26.700 617.100 28.500 ;
        RECT 618.000 26.700 624.900 28.500 ;
        RECT 632.850 28.050 633.750 29.400 ;
        RECT 634.950 28.950 637.050 31.050 ;
        RECT 637.950 28.950 640.050 31.050 ;
        RECT 640.950 28.950 643.050 31.050 ;
        RECT 632.850 27.900 637.950 28.050 ;
        RECT 632.850 27.150 640.500 27.900 ;
        RECT 636.150 26.700 640.500 27.150 ;
        RECT 618.000 25.800 619.050 26.700 ;
        RECT 636.150 26.250 637.950 26.700 ;
        RECT 597.900 24.000 605.700 25.800 ;
        RECT 609.150 24.750 619.050 25.800 ;
        RECT 609.150 22.950 610.200 24.750 ;
        RECT 619.950 24.450 627.600 25.800 ;
        RECT 619.950 23.700 620.850 24.450 ;
        RECT 601.950 21.900 610.200 22.950 ;
        RECT 611.250 22.650 620.850 23.700 ;
        RECT 601.950 17.850 604.050 21.900 ;
        RECT 611.250 21.000 612.150 22.650 ;
        RECT 621.750 21.750 625.650 23.550 ;
        RECT 626.550 22.950 627.600 24.450 ;
        RECT 628.950 25.650 631.050 25.950 ;
        RECT 628.950 23.850 632.850 25.650 ;
        RECT 639.450 23.250 640.500 26.700 ;
        RECT 642.000 25.800 643.050 28.950 ;
        RECT 644.700 29.400 646.500 35.250 ;
        RECT 650.100 29.400 651.900 35.250 ;
        RECT 655.500 29.400 657.300 35.250 ;
        RECT 663.000 29.400 664.800 35.250 ;
        RECT 667.200 31.050 669.000 35.250 ;
        RECT 670.500 32.400 672.300 35.250 ;
        RECT 680.550 32.400 682.350 35.250 ;
        RECT 683.550 32.400 685.350 35.250 ;
        RECT 686.550 32.400 688.350 35.250 ;
        RECT 695.550 32.400 697.350 35.250 ;
        RECT 698.550 32.400 700.350 35.250 ;
        RECT 701.550 32.400 703.350 35.250 ;
        RECT 667.200 29.400 672.900 31.050 ;
        RECT 644.700 28.500 646.200 29.400 ;
        RECT 644.700 27.300 653.100 28.500 ;
        RECT 651.300 26.700 653.100 27.300 ;
        RECT 656.100 25.800 657.300 29.400 ;
        RECT 642.000 24.900 657.300 25.800 ;
        RECT 626.550 22.050 638.550 22.950 ;
        RECT 605.100 19.200 612.150 21.000 ;
        RECT 613.500 19.950 615.300 21.750 ;
        RECT 621.750 21.450 623.850 21.750 ;
        RECT 625.950 20.550 628.050 20.850 ;
        RECT 634.800 20.550 636.600 21.150 ;
        RECT 625.950 19.950 636.600 20.550 ;
        RECT 613.500 19.350 636.600 19.950 ;
        RECT 637.500 20.550 638.550 22.050 ;
        RECT 639.450 21.450 641.250 23.250 ;
        RECT 643.050 22.950 654.900 24.000 ;
        RECT 643.050 20.550 644.250 22.950 ;
        RECT 653.100 21.150 654.900 22.950 ;
        RECT 637.500 19.650 644.250 20.550 ;
        RECT 646.950 19.650 649.050 19.950 ;
        RECT 613.500 18.750 628.050 19.350 ;
        RECT 645.150 18.450 649.050 19.650 ;
        RECT 652.950 19.050 655.050 21.150 ;
        RECT 635.100 17.850 649.050 18.450 ;
        RECT 609.000 17.550 648.750 17.850 ;
        RECT 597.750 16.650 599.550 17.250 ;
        RECT 609.000 16.650 637.050 17.550 ;
        RECT 597.750 15.450 610.050 16.650 ;
        RECT 637.950 16.050 640.050 16.350 ;
        RECT 647.700 16.050 649.500 16.650 ;
        RECT 610.950 14.550 613.050 15.750 ;
        RECT 595.650 13.650 613.050 14.550 ;
        RECT 616.950 14.400 637.050 15.750 ;
        RECT 616.950 13.650 619.050 14.400 ;
        RECT 598.500 9.600 599.700 13.650 ;
        RECT 600.600 11.700 602.400 12.300 ;
        RECT 607.350 12.150 609.150 12.300 ;
        RECT 600.600 10.500 606.300 11.700 ;
        RECT 607.350 10.950 616.050 12.150 ;
        RECT 607.350 10.500 609.150 10.950 ;
        RECT 548.550 3.750 550.350 9.000 ;
        RECT 551.550 3.750 553.350 9.600 ;
        RECT 562.650 3.750 564.450 9.600 ;
        RECT 565.650 3.750 567.450 9.600 ;
        RECT 568.650 3.750 570.450 9.600 ;
        RECT 575.550 3.750 577.350 9.600 ;
        RECT 578.550 3.750 580.350 9.600 ;
        RECT 581.550 3.750 583.350 9.600 ;
        RECT 588.750 3.750 590.550 9.600 ;
        RECT 591.750 3.750 593.550 9.600 ;
        RECT 595.500 3.750 597.300 9.600 ;
        RECT 598.500 3.750 600.300 9.600 ;
        RECT 601.500 3.750 603.300 9.600 ;
        RECT 604.500 3.750 606.300 10.500 ;
        RECT 613.950 10.050 616.050 10.950 ;
        RECT 607.500 3.750 609.300 9.600 ;
        RECT 610.800 7.800 612.900 9.900 ;
        RECT 611.400 6.600 612.900 7.800 ;
        RECT 611.250 3.750 613.050 6.600 ;
        RECT 614.250 3.750 616.050 10.050 ;
        RECT 617.550 6.600 618.900 13.650 ;
        RECT 635.100 13.350 637.050 14.400 ;
        RECT 637.950 14.850 649.500 16.050 ;
        RECT 637.950 14.250 640.050 14.850 ;
        RECT 651.000 13.350 652.800 14.100 ;
        RECT 620.100 10.800 624.000 12.600 ;
        RECT 621.000 10.500 624.000 10.800 ;
        RECT 625.950 12.150 628.050 12.600 ;
        RECT 635.100 12.300 652.800 13.350 ;
        RECT 625.950 10.500 628.350 12.150 ;
        RECT 617.250 3.750 619.050 6.600 ;
        RECT 621.000 3.750 622.800 10.500 ;
        RECT 627.000 9.600 628.350 10.500 ;
        RECT 634.950 9.600 637.050 10.050 ;
        RECT 624.000 3.750 625.800 9.600 ;
        RECT 627.000 3.750 628.800 9.600 ;
        RECT 630.750 3.750 632.550 9.600 ;
        RECT 634.500 7.950 637.050 9.600 ;
        RECT 637.950 7.950 640.050 10.050 ;
        RECT 640.950 7.950 643.050 10.050 ;
        RECT 634.500 6.600 635.700 7.950 ;
        RECT 637.950 6.600 638.850 7.950 ;
        RECT 640.950 6.600 642.150 7.950 ;
        RECT 633.750 3.750 635.700 6.600 ;
        RECT 636.750 3.750 638.850 6.600 ;
        RECT 639.750 3.750 642.150 6.600 ;
        RECT 643.500 3.750 645.300 7.050 ;
        RECT 646.500 3.750 648.300 12.300 ;
        RECT 656.100 11.400 657.300 24.900 ;
        RECT 662.100 24.150 663.900 25.950 ;
        RECT 661.950 22.050 664.050 24.150 ;
        RECT 664.950 23.850 667.050 25.950 ;
        RECT 668.100 24.150 669.900 25.950 ;
        RECT 665.100 22.050 666.900 23.850 ;
        RECT 667.950 22.050 670.050 24.150 ;
        RECT 671.700 22.950 672.900 29.400 ;
        RECT 684.000 25.950 685.050 32.400 ;
        RECT 699.000 25.950 700.050 32.400 ;
        RECT 710.850 29.400 712.650 35.250 ;
        RECT 715.350 28.200 717.150 35.250 ;
        RECT 725.850 29.400 727.650 35.250 ;
        RECT 730.350 28.200 732.150 35.250 ;
        RECT 737.850 29.400 739.650 35.250 ;
        RECT 742.350 28.200 744.150 35.250 ;
        RECT 682.950 23.850 685.050 25.950 ;
        RECT 697.950 23.850 700.050 25.950 ;
        RECT 670.950 20.850 673.050 22.950 ;
        RECT 679.950 20.850 682.050 22.950 ;
        RECT 671.700 15.600 672.900 20.850 ;
        RECT 680.100 19.050 681.900 20.850 ;
        RECT 684.000 16.650 685.050 23.850 ;
        RECT 685.950 20.850 688.050 22.950 ;
        RECT 694.950 20.850 697.050 22.950 ;
        RECT 686.100 19.050 687.900 20.850 ;
        RECT 695.100 19.050 696.900 20.850 ;
        RECT 699.000 16.650 700.050 23.850 ;
        RECT 713.550 27.300 717.150 28.200 ;
        RECT 728.550 27.300 732.150 28.200 ;
        RECT 740.550 27.300 744.150 28.200 ;
        RECT 700.950 20.850 703.050 22.950 ;
        RECT 710.100 21.150 711.900 22.950 ;
        RECT 701.100 19.050 702.900 20.850 ;
        RECT 709.950 19.050 712.050 21.150 ;
        RECT 713.550 19.950 714.750 27.300 ;
        RECT 716.100 21.150 717.900 22.950 ;
        RECT 725.100 21.150 726.900 22.950 ;
        RECT 712.950 17.850 715.050 19.950 ;
        RECT 715.950 19.050 718.050 21.150 ;
        RECT 724.950 19.050 727.050 21.150 ;
        RECT 728.550 19.950 729.750 27.300 ;
        RECT 731.100 21.150 732.900 22.950 ;
        RECT 737.100 21.150 738.900 22.950 ;
        RECT 727.950 17.850 730.050 19.950 ;
        RECT 730.950 19.050 733.050 21.150 ;
        RECT 736.950 19.050 739.050 21.150 ;
        RECT 740.550 19.950 741.750 27.300 ;
        RECT 752.700 26.400 754.500 35.250 ;
        RECT 758.100 27.000 759.900 35.250 ;
        RECT 770.850 29.400 772.650 35.250 ;
        RECT 775.350 28.200 777.150 35.250 ;
        RECT 783.750 32.400 785.550 35.250 ;
        RECT 786.750 32.400 788.550 35.250 ;
        RECT 773.550 27.300 777.150 28.200 ;
        RECT 758.100 25.350 762.600 27.000 ;
        RECT 743.100 21.150 744.900 22.950 ;
        RECT 761.400 21.150 762.600 25.350 ;
        RECT 770.100 21.150 771.900 22.950 ;
        RECT 739.950 17.850 742.050 19.950 ;
        RECT 742.950 19.050 745.050 21.150 ;
        RECT 751.950 17.850 754.050 19.950 ;
        RECT 757.950 17.850 760.050 19.950 ;
        RECT 760.950 19.050 763.050 21.150 ;
        RECT 769.950 19.050 772.050 21.150 ;
        RECT 773.550 19.950 774.750 27.300 ;
        RECT 787.050 24.150 788.550 32.400 ;
        RECT 776.100 21.150 777.900 22.950 ;
        RECT 784.950 22.050 788.550 24.150 ;
        RECT 684.000 15.600 686.550 16.650 ;
        RECT 699.000 15.600 701.550 16.650 ;
        RECT 653.250 10.500 657.300 11.400 ;
        RECT 662.550 14.700 670.350 15.600 ;
        RECT 653.250 9.600 654.300 10.500 ;
        RECT 649.500 3.750 651.300 9.600 ;
        RECT 652.500 3.750 654.300 9.600 ;
        RECT 655.500 3.750 657.300 9.600 ;
        RECT 662.550 3.750 664.350 14.700 ;
        RECT 665.550 3.750 667.350 13.800 ;
        RECT 668.550 3.750 670.350 14.700 ;
        RECT 671.550 3.750 673.350 15.600 ;
        RECT 680.550 3.750 682.350 15.600 ;
        RECT 684.750 3.750 686.550 15.600 ;
        RECT 695.550 3.750 697.350 15.600 ;
        RECT 699.750 3.750 701.550 15.600 ;
        RECT 713.550 9.600 714.750 17.850 ;
        RECT 728.550 9.600 729.750 17.850 ;
        RECT 740.550 9.600 741.750 17.850 ;
        RECT 752.100 16.050 753.900 17.850 ;
        RECT 754.950 14.850 757.050 16.950 ;
        RECT 758.250 16.050 760.050 17.850 ;
        RECT 755.100 13.050 756.900 14.850 ;
        RECT 761.700 10.800 762.750 19.050 ;
        RECT 772.950 17.850 775.050 19.950 ;
        RECT 775.950 19.050 778.050 21.150 ;
        RECT 755.700 9.900 762.750 10.800 ;
        RECT 755.700 9.600 757.350 9.900 ;
        RECT 710.550 3.750 712.350 9.600 ;
        RECT 713.550 3.750 715.350 9.600 ;
        RECT 716.550 3.750 718.350 9.600 ;
        RECT 725.550 3.750 727.350 9.600 ;
        RECT 728.550 3.750 730.350 9.600 ;
        RECT 731.550 3.750 733.350 9.600 ;
        RECT 737.550 3.750 739.350 9.600 ;
        RECT 740.550 3.750 742.350 9.600 ;
        RECT 743.550 3.750 745.350 9.600 ;
        RECT 752.550 3.750 754.350 9.600 ;
        RECT 755.550 3.750 757.350 9.600 ;
        RECT 761.550 9.600 762.750 9.900 ;
        RECT 773.550 9.600 774.750 17.850 ;
        RECT 787.050 9.600 788.550 22.050 ;
        RECT 790.650 29.400 792.450 35.250 ;
        RECT 796.050 29.400 797.850 35.250 ;
        RECT 801.600 30.600 803.400 35.250 ;
        RECT 806.250 31.500 808.050 35.250 ;
        RECT 809.250 31.500 811.050 35.250 ;
        RECT 812.250 31.500 814.050 35.250 ;
        RECT 799.200 29.400 803.400 30.600 ;
        RECT 805.950 29.400 808.050 31.500 ;
        RECT 808.950 29.400 811.050 31.500 ;
        RECT 811.950 29.400 814.050 31.500 ;
        RECT 816.000 31.500 817.800 35.250 ;
        RECT 819.000 32.400 820.800 35.250 ;
        RECT 822.000 31.500 823.800 35.250 ;
        RECT 826.500 32.400 828.300 35.250 ;
        RECT 829.500 32.400 831.300 35.250 ;
        RECT 832.500 32.400 834.300 35.250 ;
        RECT 835.500 32.400 837.300 35.250 ;
        RECT 816.000 29.700 818.850 31.500 ;
        RECT 816.750 29.400 818.850 29.700 ;
        RECT 820.950 29.700 823.800 31.500 ;
        RECT 824.700 30.750 826.500 31.200 ;
        RECT 829.950 31.050 831.300 32.400 ;
        RECT 832.950 31.050 834.300 32.400 ;
        RECT 835.950 31.050 837.300 32.400 ;
        RECT 820.950 29.400 823.050 29.700 ;
        RECT 824.700 29.400 828.750 30.750 ;
        RECT 790.650 14.550 791.850 29.400 ;
        RECT 799.200 25.800 800.700 29.400 ;
        RECT 805.350 26.700 812.100 28.500 ;
        RECT 813.000 26.700 819.900 28.500 ;
        RECT 827.850 28.050 828.750 29.400 ;
        RECT 829.950 28.950 832.050 31.050 ;
        RECT 832.950 28.950 835.050 31.050 ;
        RECT 835.950 28.950 838.050 31.050 ;
        RECT 827.850 27.900 832.950 28.050 ;
        RECT 827.850 27.150 835.500 27.900 ;
        RECT 831.150 26.700 835.500 27.150 ;
        RECT 813.000 25.800 814.050 26.700 ;
        RECT 831.150 26.250 832.950 26.700 ;
        RECT 792.900 24.000 800.700 25.800 ;
        RECT 804.150 24.750 814.050 25.800 ;
        RECT 804.150 22.950 805.200 24.750 ;
        RECT 814.950 24.450 822.600 25.800 ;
        RECT 814.950 23.700 815.850 24.450 ;
        RECT 796.950 21.900 805.200 22.950 ;
        RECT 806.250 22.650 815.850 23.700 ;
        RECT 796.950 17.850 799.050 21.900 ;
        RECT 806.250 21.000 807.150 22.650 ;
        RECT 816.750 21.750 820.650 23.550 ;
        RECT 821.550 22.950 822.600 24.450 ;
        RECT 823.950 25.650 826.050 25.950 ;
        RECT 823.950 23.850 827.850 25.650 ;
        RECT 834.450 23.250 835.500 26.700 ;
        RECT 837.000 25.800 838.050 28.950 ;
        RECT 839.700 29.400 841.500 35.250 ;
        RECT 845.100 29.400 846.900 35.250 ;
        RECT 850.500 29.400 852.300 35.250 ;
        RECT 839.700 28.500 841.200 29.400 ;
        RECT 839.700 27.300 848.100 28.500 ;
        RECT 846.300 26.700 848.100 27.300 ;
        RECT 851.100 25.800 852.300 29.400 ;
        RECT 837.000 24.900 852.300 25.800 ;
        RECT 821.550 22.050 833.550 22.950 ;
        RECT 800.100 19.200 807.150 21.000 ;
        RECT 808.500 19.950 810.300 21.750 ;
        RECT 816.750 21.450 818.850 21.750 ;
        RECT 820.950 20.550 823.050 20.850 ;
        RECT 829.800 20.550 831.600 21.150 ;
        RECT 820.950 19.950 831.600 20.550 ;
        RECT 808.500 19.350 831.600 19.950 ;
        RECT 832.500 20.550 833.550 22.050 ;
        RECT 834.450 21.450 836.250 23.250 ;
        RECT 838.050 22.950 849.900 24.000 ;
        RECT 838.050 20.550 839.250 22.950 ;
        RECT 848.100 21.150 849.900 22.950 ;
        RECT 832.500 19.650 839.250 20.550 ;
        RECT 841.950 19.650 844.050 19.950 ;
        RECT 808.500 18.750 823.050 19.350 ;
        RECT 840.150 18.450 844.050 19.650 ;
        RECT 847.950 19.050 850.050 21.150 ;
        RECT 830.100 17.850 844.050 18.450 ;
        RECT 804.000 17.550 843.750 17.850 ;
        RECT 792.750 16.650 794.550 17.250 ;
        RECT 804.000 16.650 832.050 17.550 ;
        RECT 792.750 15.450 805.050 16.650 ;
        RECT 832.950 16.050 835.050 16.350 ;
        RECT 842.700 16.050 844.500 16.650 ;
        RECT 805.950 14.550 808.050 15.750 ;
        RECT 790.650 13.650 808.050 14.550 ;
        RECT 811.950 14.400 832.050 15.750 ;
        RECT 811.950 13.650 814.050 14.400 ;
        RECT 793.500 9.600 794.700 13.650 ;
        RECT 795.600 11.700 797.400 12.300 ;
        RECT 802.350 12.150 804.150 12.300 ;
        RECT 795.600 10.500 801.300 11.700 ;
        RECT 802.350 10.950 811.050 12.150 ;
        RECT 802.350 10.500 804.150 10.950 ;
        RECT 758.550 3.750 760.350 9.000 ;
        RECT 761.550 3.750 763.350 9.600 ;
        RECT 770.550 3.750 772.350 9.600 ;
        RECT 773.550 3.750 775.350 9.600 ;
        RECT 776.550 3.750 778.350 9.600 ;
        RECT 783.750 3.750 785.550 9.600 ;
        RECT 786.750 3.750 788.550 9.600 ;
        RECT 790.500 3.750 792.300 9.600 ;
        RECT 793.500 3.750 795.300 9.600 ;
        RECT 796.500 3.750 798.300 9.600 ;
        RECT 799.500 3.750 801.300 10.500 ;
        RECT 808.950 10.050 811.050 10.950 ;
        RECT 802.500 3.750 804.300 9.600 ;
        RECT 805.800 7.800 807.900 9.900 ;
        RECT 806.400 6.600 807.900 7.800 ;
        RECT 806.250 3.750 808.050 6.600 ;
        RECT 809.250 3.750 811.050 10.050 ;
        RECT 812.550 6.600 813.900 13.650 ;
        RECT 830.100 13.350 832.050 14.400 ;
        RECT 832.950 14.850 844.500 16.050 ;
        RECT 832.950 14.250 835.050 14.850 ;
        RECT 846.000 13.350 847.800 14.100 ;
        RECT 815.100 10.800 819.000 12.600 ;
        RECT 816.000 10.500 819.000 10.800 ;
        RECT 820.950 12.150 823.050 12.600 ;
        RECT 830.100 12.300 847.800 13.350 ;
        RECT 820.950 10.500 823.350 12.150 ;
        RECT 812.250 3.750 814.050 6.600 ;
        RECT 816.000 3.750 817.800 10.500 ;
        RECT 822.000 9.600 823.350 10.500 ;
        RECT 829.950 9.600 832.050 10.050 ;
        RECT 819.000 3.750 820.800 9.600 ;
        RECT 822.000 3.750 823.800 9.600 ;
        RECT 825.750 3.750 827.550 9.600 ;
        RECT 829.500 7.950 832.050 9.600 ;
        RECT 832.950 7.950 835.050 10.050 ;
        RECT 835.950 7.950 838.050 10.050 ;
        RECT 829.500 6.600 830.700 7.950 ;
        RECT 832.950 6.600 833.850 7.950 ;
        RECT 835.950 6.600 837.150 7.950 ;
        RECT 828.750 3.750 830.700 6.600 ;
        RECT 831.750 3.750 833.850 6.600 ;
        RECT 834.750 3.750 837.150 6.600 ;
        RECT 838.500 3.750 840.300 7.050 ;
        RECT 841.500 3.750 843.300 12.300 ;
        RECT 851.100 11.400 852.300 24.900 ;
        RECT 848.250 10.500 852.300 11.400 ;
        RECT 848.250 9.600 849.300 10.500 ;
        RECT 844.500 3.750 846.300 9.600 ;
        RECT 847.500 3.750 849.300 9.600 ;
        RECT 850.500 3.750 852.300 9.600 ;
      LAYER metal2 ;
        RECT 64.950 820.950 67.050 823.050 ;
        RECT 67.950 820.950 70.050 823.050 ;
        RECT 70.950 820.950 73.050 823.050 ;
        RECT 79.950 821.400 82.050 823.500 ;
        RECT 84.150 821.400 86.250 823.500 ;
        RECT 88.950 821.400 91.050 823.500 ;
        RECT 91.950 821.400 94.050 823.500 ;
        RECT 94.950 821.400 97.050 823.500 ;
        RECT 10.950 817.950 13.050 820.050 ;
        RECT 22.950 817.950 25.050 820.050 ;
        RECT 28.950 817.950 31.050 820.050 ;
        RECT 37.950 817.950 40.050 820.050 ;
        RECT 40.950 817.950 43.050 820.050 ;
        RECT 11.400 817.050 12.450 817.950 ;
        RECT 7.950 814.950 10.050 817.050 ;
        RECT 10.950 814.950 13.050 817.050 ;
        RECT 16.950 816.450 19.050 817.050 ;
        RECT 14.250 815.250 15.750 816.150 ;
        RECT 16.950 815.400 21.450 816.450 ;
        RECT 16.950 814.950 19.050 815.400 ;
        RECT 8.400 814.050 9.450 814.950 ;
        RECT 7.950 811.950 10.050 814.050 ;
        RECT 11.250 812.850 12.750 813.750 ;
        RECT 13.950 811.950 16.050 814.050 ;
        RECT 17.250 812.850 19.050 813.750 ;
        RECT 7.950 809.850 10.050 810.750 ;
        RECT 14.400 808.050 15.450 811.950 ;
        RECT 20.400 810.450 21.450 815.400 ;
        RECT 23.400 811.050 24.450 817.950 ;
        RECT 29.400 814.050 30.450 817.950 ;
        RECT 38.400 817.050 39.450 817.950 ;
        RECT 37.950 814.950 40.050 817.050 ;
        RECT 41.250 815.850 42.750 816.750 ;
        RECT 43.950 816.450 46.050 817.050 ;
        RECT 43.950 815.400 51.450 816.450 ;
        RECT 43.950 814.950 46.050 815.400 ;
        RECT 25.950 812.250 27.750 813.150 ;
        RECT 28.950 811.950 31.050 814.050 ;
        RECT 32.250 812.250 34.050 813.150 ;
        RECT 37.950 812.850 40.050 813.750 ;
        RECT 43.950 812.850 46.050 813.750 ;
        RECT 17.400 809.400 21.450 810.450 ;
        RECT 7.950 805.950 10.050 808.050 ;
        RECT 13.950 805.950 16.050 808.050 ;
        RECT 8.400 778.050 9.450 805.950 ;
        RECT 7.950 777.450 10.050 778.050 ;
        RECT 5.400 776.400 10.050 777.450 ;
        RECT 13.950 777.450 16.050 778.050 ;
        RECT 17.400 777.450 18.450 809.400 ;
        RECT 22.950 808.950 25.050 811.050 ;
        RECT 25.950 808.950 28.050 811.050 ;
        RECT 29.250 809.850 30.750 810.750 ;
        RECT 31.950 808.950 34.050 811.050 ;
        RECT 26.400 805.050 27.450 808.950 ;
        RECT 25.950 802.950 28.050 805.050 ;
        RECT 5.400 769.050 6.450 776.400 ;
        RECT 7.950 775.950 10.050 776.400 ;
        RECT 11.250 776.250 12.750 777.150 ;
        RECT 13.950 776.400 18.450 777.450 ;
        RECT 13.950 775.950 16.050 776.400 ;
        RECT 7.950 773.850 9.750 774.750 ;
        RECT 10.950 772.950 13.050 775.050 ;
        RECT 14.250 773.850 16.050 774.750 ;
        RECT 4.950 766.950 7.050 769.050 ;
        RECT 17.400 763.050 18.450 776.400 ;
        RECT 28.950 775.950 31.050 778.050 ;
        RECT 40.950 775.950 43.050 778.050 ;
        RECT 44.250 776.250 45.750 777.150 ;
        RECT 46.950 775.950 49.050 778.050 ;
        RECT 29.400 775.050 30.450 775.950 ;
        RECT 22.950 773.250 25.050 774.150 ;
        RECT 28.950 772.950 31.050 775.050 ;
        RECT 40.950 773.850 42.750 774.750 ;
        RECT 43.950 772.950 46.050 775.050 ;
        RECT 47.250 773.850 49.050 774.750 ;
        RECT 19.950 770.250 21.750 771.150 ;
        RECT 22.950 769.950 25.050 772.050 ;
        RECT 28.950 770.850 31.050 771.750 ;
        RECT 19.950 766.950 22.050 769.050 ;
        RECT 23.400 763.050 24.450 769.950 ;
        RECT 44.400 769.050 45.450 772.950 ;
        RECT 50.400 772.050 51.450 815.400 ;
        RECT 52.950 812.250 55.050 813.150 ;
        RECT 52.950 808.950 55.050 811.050 ;
        RECT 58.950 809.850 61.050 810.750 ;
        RECT 53.400 799.050 54.450 808.950 ;
        RECT 65.550 802.050 66.750 820.950 ;
        RECT 68.550 808.350 69.750 820.950 ;
        RECT 67.950 806.250 70.050 808.350 ;
        RECT 68.550 802.050 69.750 806.250 ;
        RECT 71.550 802.050 72.750 820.950 ;
        RECT 76.950 817.950 79.050 820.050 ;
        RECT 76.950 815.850 79.050 816.750 ;
        RECT 80.250 812.850 81.450 821.400 ;
        RECT 84.450 815.550 85.650 821.400 ;
        RECT 84.150 813.450 86.250 815.550 ;
        RECT 79.950 810.750 82.050 812.850 ;
        RECT 80.250 804.600 81.450 810.750 ;
        RECT 84.450 804.600 85.650 813.450 ;
        RECT 89.400 807.750 90.600 821.400 ;
        RECT 88.950 805.650 91.050 807.750 ;
        RECT 79.950 802.500 82.050 804.600 ;
        RECT 84.000 802.500 86.100 804.600 ;
        RECT 92.550 804.150 93.750 821.400 ;
        RECT 95.250 807.750 96.450 821.400 ;
        RECT 181.950 820.950 184.050 823.050 ;
        RECT 241.950 820.950 244.050 823.050 ;
        RECT 274.950 820.950 277.050 823.050 ;
        RECT 283.950 820.950 286.050 823.050 ;
        RECT 286.950 820.950 289.050 823.050 ;
        RECT 289.950 820.950 292.050 823.050 ;
        RECT 298.950 821.400 301.050 823.500 ;
        RECT 303.150 821.400 305.250 823.500 ;
        RECT 307.950 821.400 310.050 823.500 ;
        RECT 310.950 821.400 313.050 823.500 ;
        RECT 313.950 821.400 316.050 823.500 ;
        RECT 118.950 817.950 121.050 820.050 ;
        RECT 130.950 817.950 133.050 820.050 ;
        RECT 136.950 817.950 139.050 820.050 ;
        RECT 115.950 815.250 118.050 816.150 ;
        RECT 103.950 811.950 106.050 814.050 ;
        RECT 115.950 813.450 118.050 814.050 ;
        RECT 119.400 813.450 120.450 817.950 ;
        RECT 127.950 815.250 130.050 816.150 ;
        RECT 130.950 815.850 133.050 816.750 ;
        RECT 115.950 812.400 120.450 813.450 ;
        RECT 115.950 811.950 118.050 812.400 ;
        RECT 121.950 811.950 124.050 814.050 ;
        RECT 127.950 811.950 130.050 814.050 ;
        RECT 103.950 809.850 106.050 810.750 ;
        RECT 94.950 805.650 97.050 807.750 ;
        RECT 91.950 802.050 94.050 804.150 ;
        RECT 64.950 799.950 67.050 802.050 ;
        RECT 67.950 799.950 70.050 802.050 ;
        RECT 70.950 799.950 73.050 802.050 ;
        RECT 95.250 801.900 96.450 805.650 ;
        RECT 95.100 799.800 97.200 801.900 ;
        RECT 52.950 796.950 55.050 799.050 ;
        RECT 67.950 796.950 70.050 799.050 ;
        RECT 68.400 778.050 69.450 796.950 ;
        RECT 79.950 784.950 82.050 787.050 ;
        RECT 82.950 784.950 85.050 787.050 ;
        RECT 85.950 784.950 88.050 787.050 ;
        RECT 110.100 785.100 112.200 787.200 ;
        RECT 67.950 777.450 70.050 778.050 ;
        RECT 67.950 776.400 72.450 777.450 ;
        RECT 67.950 775.950 70.050 776.400 ;
        RECT 52.950 773.250 55.050 774.150 ;
        RECT 58.950 773.250 61.050 774.150 ;
        RECT 67.950 773.850 70.050 774.750 ;
        RECT 49.950 769.950 52.050 772.050 ;
        RECT 52.950 769.950 55.050 772.050 ;
        RECT 56.250 770.250 57.750 771.150 ;
        RECT 58.950 769.950 61.050 772.050 ;
        RECT 53.400 769.050 54.450 769.950 ;
        RECT 25.950 766.950 28.050 769.050 ;
        RECT 43.950 766.950 46.050 769.050 ;
        RECT 52.950 766.950 55.050 769.050 ;
        RECT 55.950 766.950 58.050 769.050 ;
        RECT 16.950 760.950 19.050 763.050 ;
        RECT 22.950 760.950 25.050 763.050 ;
        RECT 16.950 748.950 19.050 751.050 ;
        RECT 19.950 748.950 22.050 751.050 ;
        RECT 22.950 748.950 25.050 751.050 ;
        RECT 4.950 740.250 7.050 741.150 ;
        RECT 4.950 736.950 7.050 739.050 ;
        RECT 10.950 737.850 13.050 738.750 ;
        RECT 5.400 715.050 6.450 736.950 ;
        RECT 17.550 730.050 18.750 748.950 ;
        RECT 20.550 736.350 21.750 748.950 ;
        RECT 19.950 734.250 22.050 736.350 ;
        RECT 20.550 730.050 21.750 734.250 ;
        RECT 23.550 730.050 24.750 748.950 ;
        RECT 16.950 727.950 19.050 730.050 ;
        RECT 19.950 727.950 22.050 730.050 ;
        RECT 22.950 727.950 25.050 730.050 ;
        RECT 4.950 712.950 7.050 715.050 ;
        RECT 26.400 709.050 27.450 766.950 ;
        RECT 56.400 757.050 57.450 766.950 ;
        RECT 28.950 754.950 31.050 757.050 ;
        RECT 55.950 754.950 58.050 757.050 ;
        RECT 29.400 748.050 30.450 754.950 ;
        RECT 55.950 751.950 58.050 754.050 ;
        RECT 31.950 749.400 34.050 751.500 ;
        RECT 36.150 749.400 38.250 751.500 ;
        RECT 40.950 749.400 43.050 751.500 ;
        RECT 43.950 749.400 46.050 751.500 ;
        RECT 46.950 749.400 49.050 751.500 ;
        RECT 28.950 745.950 31.050 748.050 ;
        RECT 28.950 743.850 31.050 744.750 ;
        RECT 32.250 740.850 33.450 749.400 ;
        RECT 36.450 743.550 37.650 749.400 ;
        RECT 36.150 741.450 38.250 743.550 ;
        RECT 31.950 738.750 34.050 740.850 ;
        RECT 32.250 732.600 33.450 738.750 ;
        RECT 36.450 732.600 37.650 741.450 ;
        RECT 41.400 735.750 42.600 749.400 ;
        RECT 40.950 733.650 43.050 735.750 ;
        RECT 31.950 730.500 34.050 732.600 ;
        RECT 36.000 730.500 38.100 732.600 ;
        RECT 44.550 732.150 45.750 749.400 ;
        RECT 47.250 735.750 48.450 749.400 ;
        RECT 56.400 742.050 57.450 751.950 ;
        RECT 59.400 748.050 60.450 769.950 ;
        RECT 58.950 745.950 61.050 748.050 ;
        RECT 55.950 739.950 58.050 742.050 ;
        RECT 55.950 737.850 58.050 738.750 ;
        RECT 46.950 733.650 49.050 735.750 ;
        RECT 43.950 730.050 46.050 732.150 ;
        RECT 47.250 729.900 48.450 733.650 ;
        RECT 47.100 727.800 49.200 729.900 ;
        RECT 59.400 718.050 60.450 745.950 ;
        RECT 67.950 743.250 70.050 744.150 ;
        RECT 67.950 739.950 70.050 742.050 ;
        RECT 68.400 739.050 69.450 739.950 ;
        RECT 67.950 736.950 70.050 739.050 ;
        RECT 28.950 715.950 31.050 718.050 ;
        RECT 58.950 715.950 61.050 718.050 ;
        RECT 13.950 706.950 16.050 709.050 ;
        RECT 25.950 706.950 28.050 709.050 ;
        RECT 14.400 706.050 15.450 706.950 ;
        RECT 7.950 703.950 10.050 706.050 ;
        RECT 11.250 704.250 12.750 705.150 ;
        RECT 13.950 703.950 16.050 706.050 ;
        RECT 7.950 701.850 9.750 702.750 ;
        RECT 10.950 700.950 13.050 703.050 ;
        RECT 14.250 701.850 16.050 702.750 ;
        RECT 19.950 701.250 22.050 702.150 ;
        RECT 25.950 701.250 28.050 702.150 ;
        RECT 19.950 697.950 22.050 700.050 ;
        RECT 25.950 699.450 28.050 700.050 ;
        RECT 29.400 699.450 30.450 715.950 ;
        RECT 71.400 715.050 72.450 776.400 ;
        RECT 73.950 776.250 76.050 777.150 ;
        RECT 80.550 766.050 81.750 784.950 ;
        RECT 83.550 780.750 84.750 784.950 ;
        RECT 82.950 778.650 85.050 780.750 ;
        RECT 83.550 766.050 84.750 778.650 ;
        RECT 86.550 766.050 87.750 784.950 ;
        RECT 94.950 782.400 97.050 784.500 ;
        RECT 99.000 782.400 101.100 784.500 ;
        RECT 106.950 782.850 109.050 784.950 ;
        RECT 95.250 776.250 96.450 782.400 ;
        RECT 94.950 774.150 97.050 776.250 ;
        RECT 91.950 770.250 94.050 771.150 ;
        RECT 91.950 766.950 94.050 769.050 ;
        RECT 79.950 763.950 82.050 766.050 ;
        RECT 82.950 763.950 85.050 766.050 ;
        RECT 85.950 763.950 88.050 766.050 ;
        RECT 92.400 760.050 93.450 766.950 ;
        RECT 95.250 765.600 96.450 774.150 ;
        RECT 99.450 773.550 100.650 782.400 ;
        RECT 103.950 779.250 106.050 781.350 ;
        RECT 99.150 771.450 101.250 773.550 ;
        RECT 99.450 765.600 100.650 771.450 ;
        RECT 104.400 765.600 105.600 779.250 ;
        RECT 107.550 765.600 108.750 782.850 ;
        RECT 110.250 781.350 111.450 785.100 ;
        RECT 109.950 779.250 112.050 781.350 ;
        RECT 110.250 765.600 111.450 779.250 ;
        RECT 118.950 776.250 121.050 777.150 ;
        RECT 118.950 774.450 121.050 775.050 ;
        RECT 122.400 774.450 123.450 811.950 ;
        RECT 124.950 808.950 127.050 811.050 ;
        RECT 118.950 773.400 123.450 774.450 ;
        RECT 118.950 772.950 121.050 773.400 ;
        RECT 115.950 766.950 118.050 769.050 ;
        RECT 94.950 763.500 97.050 765.600 ;
        RECT 99.150 763.500 101.250 765.600 ;
        RECT 103.950 763.500 106.050 765.600 ;
        RECT 106.950 763.500 109.050 765.600 ;
        RECT 109.950 763.500 112.050 765.600 ;
        RECT 76.950 757.950 79.050 760.050 ;
        RECT 91.950 757.950 94.050 760.050 ;
        RECT 77.400 748.050 78.450 757.950 ;
        RECT 91.950 748.950 94.050 751.050 ;
        RECT 73.950 745.950 76.050 748.050 ;
        RECT 76.950 745.950 79.050 748.050 ;
        RECT 74.400 745.050 75.450 745.950 ;
        RECT 73.950 742.950 76.050 745.050 ;
        RECT 77.250 743.850 78.750 744.750 ;
        RECT 79.950 742.950 82.050 745.050 ;
        RECT 73.950 740.850 76.050 741.750 ;
        RECT 79.950 740.850 82.050 741.750 ;
        RECT 92.400 738.450 93.450 748.950 ;
        RECT 116.400 745.050 117.450 766.950 ;
        RECT 119.400 757.050 120.450 772.950 ;
        RECT 125.400 763.050 126.450 808.950 ;
        RECT 130.950 772.950 133.050 775.050 ;
        RECT 133.950 772.950 136.050 775.050 ;
        RECT 130.950 770.850 133.050 771.750 ;
        RECT 124.950 760.950 127.050 763.050 ;
        RECT 118.950 754.950 121.050 757.050 ;
        RECT 119.400 754.050 120.450 754.950 ;
        RECT 118.950 751.950 121.050 754.050 ;
        RECT 118.950 745.950 121.050 748.050 ;
        RECT 97.950 742.950 100.050 745.050 ;
        RECT 103.950 742.950 106.050 745.050 ;
        RECT 109.950 742.950 112.050 745.050 ;
        RECT 113.250 743.250 114.750 744.150 ;
        RECT 115.950 742.950 118.050 745.050 ;
        RECT 98.400 742.050 99.450 742.950 ;
        RECT 94.950 740.250 96.750 741.150 ;
        RECT 97.950 739.950 100.050 742.050 ;
        RECT 101.250 740.250 103.050 741.150 ;
        RECT 94.950 738.450 97.050 739.050 ;
        RECT 92.400 737.400 97.050 738.450 ;
        RECT 98.250 737.850 99.750 738.750 ;
        RECT 100.950 738.450 103.050 739.050 ;
        RECT 104.400 738.450 105.450 742.950 ;
        RECT 106.950 739.950 109.050 742.050 ;
        RECT 110.250 740.850 111.750 741.750 ;
        RECT 112.950 739.950 115.050 742.050 ;
        RECT 116.250 740.850 118.050 741.750 ;
        RECT 94.950 736.950 97.050 737.400 ;
        RECT 100.950 737.400 105.450 738.450 ;
        RECT 106.950 737.850 109.050 738.750 ;
        RECT 100.950 736.950 103.050 737.400 ;
        RECT 109.950 733.950 112.050 736.050 ;
        RECT 34.950 712.950 37.050 715.050 ;
        RECT 46.950 712.950 49.050 715.050 ;
        RECT 49.950 712.950 52.050 715.050 ;
        RECT 52.950 712.950 55.050 715.050 ;
        RECT 70.950 712.950 73.050 715.050 ;
        RECT 77.100 713.100 79.200 715.200 ;
        RECT 35.400 706.050 36.450 712.950 ;
        RECT 34.950 703.950 37.050 706.050 ;
        RECT 40.950 704.250 43.050 705.150 ;
        RECT 34.950 701.850 37.050 702.750 ;
        RECT 23.250 698.250 24.750 699.150 ;
        RECT 25.950 698.400 30.450 699.450 ;
        RECT 25.950 697.950 28.050 698.400 ;
        RECT 20.400 697.050 21.450 697.950 ;
        RECT 19.950 694.950 22.050 697.050 ;
        RECT 22.950 694.950 25.050 697.050 ;
        RECT 16.950 676.950 19.050 679.050 ;
        RECT 19.950 676.950 22.050 679.050 ;
        RECT 22.950 676.950 25.050 679.050 ;
        RECT 4.950 668.250 7.050 669.150 ;
        RECT 4.950 664.950 7.050 667.050 ;
        RECT 10.950 665.850 13.050 666.750 ;
        RECT 5.400 634.050 6.450 664.950 ;
        RECT 17.550 658.050 18.750 676.950 ;
        RECT 20.550 664.350 21.750 676.950 ;
        RECT 19.950 662.250 22.050 664.350 ;
        RECT 20.550 658.050 21.750 662.250 ;
        RECT 23.550 658.050 24.750 676.950 ;
        RECT 16.950 655.950 19.050 658.050 ;
        RECT 19.950 655.950 22.050 658.050 ;
        RECT 22.950 655.950 25.050 658.050 ;
        RECT 16.950 640.950 19.050 643.050 ;
        RECT 19.950 640.950 22.050 643.050 ;
        RECT 22.950 640.950 25.050 643.050 ;
        RECT 4.950 633.450 7.050 634.050 ;
        RECT 4.950 632.400 9.450 633.450 ;
        RECT 4.950 631.950 7.050 632.400 ;
        RECT 4.950 629.850 7.050 630.750 ;
        RECT 8.400 601.050 9.450 632.400 ;
        RECT 10.950 632.250 13.050 633.150 ;
        RECT 17.550 622.050 18.750 640.950 ;
        RECT 20.550 636.750 21.750 640.950 ;
        RECT 19.950 634.650 22.050 636.750 ;
        RECT 20.550 622.050 21.750 634.650 ;
        RECT 23.550 622.050 24.750 640.950 ;
        RECT 26.400 628.050 27.450 697.950 ;
        RECT 47.550 694.050 48.750 712.950 ;
        RECT 50.550 708.750 51.750 712.950 ;
        RECT 49.950 706.650 52.050 708.750 ;
        RECT 50.550 694.050 51.750 706.650 ;
        RECT 53.550 694.050 54.750 712.950 ;
        RECT 61.950 710.400 64.050 712.500 ;
        RECT 66.000 710.400 68.100 712.500 ;
        RECT 73.950 710.850 76.050 712.950 ;
        RECT 62.250 704.250 63.450 710.400 ;
        RECT 61.950 702.150 64.050 704.250 ;
        RECT 58.950 698.250 61.050 699.150 ;
        RECT 58.950 694.950 61.050 697.050 ;
        RECT 46.950 691.950 49.050 694.050 ;
        RECT 49.950 691.950 52.050 694.050 ;
        RECT 52.950 691.950 55.050 694.050 ;
        RECT 62.250 693.600 63.450 702.150 ;
        RECT 66.450 701.550 67.650 710.400 ;
        RECT 70.950 707.250 73.050 709.350 ;
        RECT 66.150 699.450 68.250 701.550 ;
        RECT 66.450 693.600 67.650 699.450 ;
        RECT 71.400 693.600 72.600 707.250 ;
        RECT 74.550 693.600 75.750 710.850 ;
        RECT 77.250 709.350 78.450 713.100 ;
        RECT 76.950 707.250 79.050 709.350 ;
        RECT 77.250 693.600 78.450 707.250 ;
        RECT 82.950 703.950 85.050 706.050 ;
        RECT 85.950 704.250 88.050 705.150 ;
        RECT 97.950 703.950 100.050 706.050 ;
        RECT 61.950 691.500 64.050 693.600 ;
        RECT 66.150 691.500 68.250 693.600 ;
        RECT 70.950 691.500 73.050 693.600 ;
        RECT 73.950 691.500 76.050 693.600 ;
        RECT 76.950 691.500 79.050 693.600 ;
        RECT 31.950 677.400 34.050 679.500 ;
        RECT 36.150 677.400 38.250 679.500 ;
        RECT 40.950 677.400 43.050 679.500 ;
        RECT 43.950 677.400 46.050 679.500 ;
        RECT 46.950 677.400 49.050 679.500 ;
        RECT 28.950 673.950 31.050 676.050 ;
        RECT 28.950 671.850 31.050 672.750 ;
        RECT 32.250 668.850 33.450 677.400 ;
        RECT 36.450 671.550 37.650 677.400 ;
        RECT 36.150 669.450 38.250 671.550 ;
        RECT 31.950 666.750 34.050 668.850 ;
        RECT 32.250 660.600 33.450 666.750 ;
        RECT 36.450 660.600 37.650 669.450 ;
        RECT 41.400 663.750 42.600 677.400 ;
        RECT 40.950 661.650 43.050 663.750 ;
        RECT 31.950 658.500 34.050 660.600 ;
        RECT 36.000 658.500 38.100 660.600 ;
        RECT 44.550 660.150 45.750 677.400 ;
        RECT 47.250 663.750 48.450 677.400 ;
        RECT 83.400 676.050 84.450 703.950 ;
        RECT 98.400 703.050 99.450 703.950 ;
        RECT 110.400 703.050 111.450 733.950 ;
        RECT 113.400 718.050 114.450 739.950 ;
        RECT 115.950 736.950 118.050 739.050 ;
        RECT 112.950 715.950 115.050 718.050 ;
        RECT 85.950 700.950 88.050 703.050 ;
        RECT 94.950 700.950 97.050 703.050 ;
        RECT 97.950 700.950 100.050 703.050 ;
        RECT 109.950 700.950 112.050 703.050 ;
        RECT 86.400 691.050 87.450 700.950 ;
        RECT 85.950 688.950 88.050 691.050 ;
        RECT 82.950 673.950 85.050 676.050 ;
        RECT 67.950 671.250 70.050 672.150 ;
        RECT 79.950 671.250 82.050 672.150 ;
        RECT 82.950 671.850 85.050 672.750 ;
        RECT 86.400 670.050 87.450 688.950 ;
        RECT 95.400 673.050 96.450 700.950 ;
        RECT 97.950 698.850 100.050 699.750 ;
        RECT 109.950 698.850 112.050 699.750 ;
        RECT 112.950 698.250 115.050 699.150 ;
        RECT 112.950 696.450 115.050 697.050 ;
        RECT 116.400 696.450 117.450 736.950 ;
        RECT 119.400 733.050 120.450 745.950 ;
        RECT 125.400 736.050 126.450 760.950 ;
        RECT 130.950 747.450 133.050 748.050 ;
        RECT 134.400 747.450 135.450 772.950 ;
        RECT 130.950 746.400 135.450 747.450 ;
        RECT 130.950 745.950 133.050 746.400 ;
        RECT 127.950 743.250 130.050 744.150 ;
        RECT 130.950 743.850 133.050 744.750 ;
        RECT 127.950 739.950 130.050 742.050 ;
        RECT 124.950 733.950 127.050 736.050 ;
        RECT 118.950 730.950 121.050 733.050 ;
        RECT 121.950 706.950 124.050 709.050 ;
        RECT 127.950 707.250 130.050 708.150 ;
        RECT 122.400 706.050 123.450 706.950 ;
        RECT 137.400 706.050 138.450 817.950 ;
        RECT 139.950 814.950 142.050 817.050 ;
        RECT 148.950 816.450 151.050 817.050 ;
        RECT 145.950 815.250 147.750 816.150 ;
        RECT 148.950 815.400 153.450 816.450 ;
        RECT 148.950 814.950 151.050 815.400 ;
        RECT 139.950 812.850 142.050 813.750 ;
        RECT 145.950 811.950 148.050 814.050 ;
        RECT 149.250 812.850 151.050 813.750 ;
        RECT 146.400 811.050 147.450 811.950 ;
        RECT 145.950 808.950 148.050 811.050 ;
        RECT 152.400 808.050 153.450 815.400 ;
        RECT 154.950 815.250 157.050 816.150 ;
        RECT 154.950 811.950 157.050 814.050 ;
        RECT 172.950 812.250 174.750 813.150 ;
        RECT 175.950 811.950 178.050 814.050 ;
        RECT 179.250 812.250 181.050 813.150 ;
        RECT 155.400 811.050 156.450 811.950 ;
        RECT 154.950 808.950 157.050 811.050 ;
        RECT 163.950 808.950 166.050 811.050 ;
        RECT 172.950 808.950 175.050 811.050 ;
        RECT 176.250 809.850 177.750 810.750 ;
        RECT 178.950 810.450 181.050 811.050 ;
        RECT 182.400 810.450 183.450 820.950 ;
        RECT 242.400 820.050 243.450 820.950 ;
        RECT 187.950 817.950 190.050 820.050 ;
        RECT 229.950 819.450 232.050 820.050 ;
        RECT 212.400 818.400 222.450 819.450 ;
        RECT 188.400 814.050 189.450 817.950 ;
        RECT 193.950 814.950 196.050 817.050 ;
        RECT 199.950 814.950 202.050 817.050 ;
        RECT 184.950 812.250 186.750 813.150 ;
        RECT 187.950 811.950 190.050 814.050 ;
        RECT 191.250 812.250 193.050 813.150 ;
        RECT 178.950 809.400 183.450 810.450 ;
        RECT 178.950 808.950 181.050 809.400 ;
        RECT 184.950 808.950 187.050 811.050 ;
        RECT 188.250 809.850 189.750 810.750 ;
        RECT 190.950 810.450 193.050 811.050 ;
        RECT 194.400 810.450 195.450 814.950 ;
        RECT 200.400 814.050 201.450 814.950 ;
        RECT 196.950 812.250 198.750 813.150 ;
        RECT 199.950 811.950 202.050 814.050 ;
        RECT 203.250 812.250 205.050 813.150 ;
        RECT 190.950 809.400 195.450 810.450 ;
        RECT 190.950 808.950 193.050 809.400 ;
        RECT 196.950 808.950 199.050 811.050 ;
        RECT 200.250 809.850 201.750 810.750 ;
        RECT 202.950 808.950 205.050 811.050 ;
        RECT 151.950 805.950 154.050 808.050 ;
        RECT 154.950 779.250 157.050 780.150 ;
        RECT 139.950 775.950 142.050 778.050 ;
        RECT 145.950 775.950 148.050 778.050 ;
        RECT 148.950 775.950 151.050 778.050 ;
        RECT 151.950 776.250 153.750 777.150 ;
        RECT 154.950 775.950 157.050 778.050 ;
        RECT 158.250 776.250 159.750 777.150 ;
        RECT 160.950 775.950 163.050 778.050 ;
        RECT 140.400 772.050 141.450 775.950 ;
        RECT 146.400 775.050 147.450 775.950 ;
        RECT 145.950 772.950 148.050 775.050 ;
        RECT 139.950 769.950 142.050 772.050 ;
        RECT 142.950 770.250 145.050 771.150 ;
        RECT 145.950 770.850 148.050 771.750 ;
        RECT 142.950 766.950 145.050 769.050 ;
        RECT 149.400 751.050 150.450 775.950 ;
        RECT 151.950 772.950 154.050 775.050 ;
        RECT 152.400 751.050 153.450 772.950 ;
        RECT 155.400 772.050 156.450 775.950 ;
        RECT 164.400 775.050 165.450 808.950 ;
        RECT 169.950 787.950 172.050 790.050 ;
        RECT 170.400 778.050 171.450 787.950 ;
        RECT 169.950 775.950 172.050 778.050 ;
        RECT 175.950 777.450 178.050 778.050 ;
        RECT 179.400 777.450 180.450 808.950 ;
        RECT 203.400 805.050 204.450 808.950 ;
        RECT 208.950 805.950 211.050 808.050 ;
        RECT 202.950 802.950 205.050 805.050 ;
        RECT 173.250 776.250 174.750 777.150 ;
        RECT 175.950 776.400 180.450 777.450 ;
        RECT 175.950 775.950 178.050 776.400 ;
        RECT 157.950 772.950 160.050 775.050 ;
        RECT 161.250 773.850 163.050 774.750 ;
        RECT 163.950 772.950 166.050 775.050 ;
        RECT 169.950 773.850 171.750 774.750 ;
        RECT 172.950 772.950 175.050 775.050 ;
        RECT 176.250 773.850 178.050 774.750 ;
        RECT 154.950 769.950 157.050 772.050 ;
        RECT 173.400 769.050 174.450 772.950 ;
        RECT 172.950 766.950 175.050 769.050 ;
        RECT 179.400 762.450 180.450 776.400 ;
        RECT 193.950 776.250 196.050 777.150 ;
        RECT 184.950 773.250 186.750 774.150 ;
        RECT 187.950 772.950 190.050 775.050 ;
        RECT 191.250 773.250 192.750 774.150 ;
        RECT 193.950 772.950 196.050 775.050 ;
        RECT 199.950 773.250 202.050 774.150 ;
        RECT 205.950 773.250 208.050 774.150 ;
        RECT 184.950 769.950 187.050 772.050 ;
        RECT 188.250 770.850 189.750 771.750 ;
        RECT 190.950 769.950 193.050 772.050 ;
        RECT 199.950 769.950 202.050 772.050 ;
        RECT 205.950 771.450 208.050 772.050 ;
        RECT 209.400 771.450 210.450 805.950 ;
        RECT 212.400 775.050 213.450 818.400 ;
        RECT 221.400 817.050 222.450 818.400 ;
        RECT 227.400 818.400 232.050 819.450 ;
        RECT 214.950 814.950 217.050 817.050 ;
        RECT 218.250 815.250 219.750 816.150 ;
        RECT 220.950 814.950 223.050 817.050 ;
        RECT 223.950 814.950 226.050 817.050 ;
        RECT 224.400 814.050 225.450 814.950 ;
        RECT 214.950 812.850 216.750 813.750 ;
        RECT 217.950 811.950 220.050 814.050 ;
        RECT 221.250 812.850 222.750 813.750 ;
        RECT 223.950 811.950 226.050 814.050 ;
        RECT 218.400 811.050 219.450 811.950 ;
        RECT 217.950 808.950 220.050 811.050 ;
        RECT 223.950 809.850 226.050 810.750 ;
        RECT 214.950 775.950 217.050 778.050 ;
        RECT 211.950 772.950 214.050 775.050 ;
        RECT 214.950 773.850 217.050 774.750 ;
        RECT 203.250 770.250 204.750 771.150 ;
        RECT 205.950 770.400 210.450 771.450 ;
        RECT 205.950 769.950 208.050 770.400 ;
        RECT 185.400 766.050 186.450 769.950 ;
        RECT 202.950 766.950 205.050 769.050 ;
        RECT 184.950 763.950 187.050 766.050 ;
        RECT 179.400 761.400 183.450 762.450 ;
        RECT 178.950 754.950 181.050 757.050 ;
        RECT 148.950 748.950 151.050 751.050 ;
        RECT 151.950 748.950 154.050 751.050 ;
        RECT 145.950 745.950 148.050 748.050 ;
        RECT 149.400 747.450 150.450 748.950 ;
        RECT 151.950 747.450 154.050 748.050 ;
        RECT 149.400 746.400 154.050 747.450 ;
        RECT 151.950 745.950 154.050 746.400 ;
        RECT 157.950 745.950 160.050 748.050 ;
        RECT 158.400 745.050 159.450 745.950 ;
        RECT 142.950 743.250 145.050 744.150 ;
        RECT 145.950 743.850 148.050 744.750 ;
        RECT 148.950 743.250 151.050 744.150 ;
        RECT 151.950 743.850 154.050 744.750 ;
        RECT 154.950 743.250 156.750 744.150 ;
        RECT 157.950 742.950 160.050 745.050 ;
        RECT 163.950 742.950 166.050 745.050 ;
        RECT 166.950 743.250 169.050 744.150 ;
        RECT 142.950 739.950 145.050 742.050 ;
        RECT 148.950 739.950 151.050 742.050 ;
        RECT 154.950 739.950 157.050 742.050 ;
        RECT 158.250 740.850 160.050 741.750 ;
        RECT 164.400 741.450 165.450 742.950 ;
        RECT 179.400 742.050 180.450 754.950 ;
        RECT 166.950 741.450 169.050 742.050 ;
        RECT 164.400 740.400 169.050 741.450 ;
        RECT 166.950 739.950 169.050 740.400 ;
        RECT 178.950 739.950 181.050 742.050 ;
        RECT 148.950 733.950 151.050 736.050 ;
        RECT 142.950 706.950 145.050 709.050 ;
        RECT 143.400 706.050 144.450 706.950 ;
        RECT 121.950 703.950 124.050 706.050 ;
        RECT 125.250 704.250 126.750 705.150 ;
        RECT 127.950 703.950 130.050 706.050 ;
        RECT 131.250 704.250 133.050 705.150 ;
        RECT 136.950 703.950 139.050 706.050 ;
        RECT 142.950 703.950 145.050 706.050 ;
        RECT 118.950 700.950 121.050 703.050 ;
        RECT 121.950 701.850 123.750 702.750 ;
        RECT 124.950 700.950 127.050 703.050 ;
        RECT 112.950 695.400 117.450 696.450 ;
        RECT 112.950 694.950 115.050 695.400 ;
        RECT 113.400 679.050 114.450 694.950 ;
        RECT 112.950 676.950 115.050 679.050 ;
        RECT 94.950 670.950 97.050 673.050 ;
        RECT 98.250 671.250 99.750 672.150 ;
        RECT 100.950 670.950 103.050 673.050 ;
        RECT 106.950 670.950 109.050 673.050 ;
        RECT 112.950 670.950 115.050 673.050 ;
        RECT 55.950 669.450 58.050 670.050 ;
        RECT 53.400 668.400 58.050 669.450 ;
        RECT 46.950 661.650 49.050 663.750 ;
        RECT 43.950 658.050 46.050 660.150 ;
        RECT 47.250 657.900 48.450 661.650 ;
        RECT 47.100 655.800 49.200 657.900 ;
        RECT 47.100 641.100 49.200 643.200 ;
        RECT 31.950 638.400 34.050 640.500 ;
        RECT 36.000 638.400 38.100 640.500 ;
        RECT 43.950 638.850 46.050 640.950 ;
        RECT 32.250 632.250 33.450 638.400 ;
        RECT 31.950 630.150 34.050 632.250 ;
        RECT 25.950 625.950 28.050 628.050 ;
        RECT 28.950 626.250 31.050 627.150 ;
        RECT 28.950 622.950 31.050 625.050 ;
        RECT 29.400 622.050 30.450 622.950 ;
        RECT 16.950 619.950 19.050 622.050 ;
        RECT 19.950 619.950 22.050 622.050 ;
        RECT 22.950 619.950 25.050 622.050 ;
        RECT 28.950 619.950 31.050 622.050 ;
        RECT 32.250 621.600 33.450 630.150 ;
        RECT 36.450 629.550 37.650 638.400 ;
        RECT 40.950 635.250 43.050 637.350 ;
        RECT 36.150 627.450 38.250 629.550 ;
        RECT 36.450 621.600 37.650 627.450 ;
        RECT 41.400 621.600 42.600 635.250 ;
        RECT 44.550 621.600 45.750 638.850 ;
        RECT 47.250 637.350 48.450 641.100 ;
        RECT 46.950 635.250 49.050 637.350 ;
        RECT 47.250 621.600 48.450 635.250 ;
        RECT 53.400 630.450 54.450 668.400 ;
        RECT 55.950 667.950 58.050 668.400 ;
        RECT 67.950 667.950 70.050 670.050 ;
        RECT 79.950 667.950 82.050 670.050 ;
        RECT 85.950 667.950 88.050 670.050 ;
        RECT 91.950 669.450 94.050 670.050 ;
        RECT 89.400 668.400 94.050 669.450 ;
        RECT 95.250 668.850 96.750 669.750 ;
        RECT 55.950 665.850 58.050 666.750 ;
        RECT 68.400 664.050 69.450 667.950 ;
        RECT 80.400 667.050 81.450 667.950 ;
        RECT 89.400 667.050 90.450 668.400 ;
        RECT 91.950 667.950 94.050 668.400 ;
        RECT 97.950 667.950 100.050 670.050 ;
        RECT 101.250 668.850 103.050 669.750 ;
        RECT 79.950 664.950 82.050 667.050 ;
        RECT 88.950 664.950 91.050 667.050 ;
        RECT 91.950 665.850 94.050 666.750 ;
        RECT 67.950 661.950 70.050 664.050 ;
        RECT 98.400 661.050 99.450 667.950 ;
        RECT 107.400 666.450 108.450 670.950 ;
        RECT 113.400 670.050 114.450 670.950 ;
        RECT 109.950 668.250 111.750 669.150 ;
        RECT 112.950 667.950 115.050 670.050 ;
        RECT 116.250 668.250 118.050 669.150 ;
        RECT 109.950 666.450 112.050 667.050 ;
        RECT 107.400 665.400 112.050 666.450 ;
        RECT 113.250 665.850 114.750 666.750 ;
        RECT 115.950 666.450 118.050 667.050 ;
        RECT 119.400 666.450 120.450 700.950 ;
        RECT 128.400 700.050 129.450 703.950 ;
        RECT 130.950 700.950 133.050 703.050 ;
        RECT 136.950 701.250 139.050 702.150 ;
        RECT 142.950 701.850 145.050 702.750 ;
        RECT 145.950 701.250 148.050 702.150 ;
        RECT 127.950 697.950 130.050 700.050 ;
        RECT 131.400 696.450 132.450 700.950 ;
        RECT 136.950 697.950 139.050 700.050 ;
        RECT 145.950 697.950 148.050 700.050 ;
        RECT 133.950 696.450 136.050 697.050 ;
        RECT 131.400 695.400 136.050 696.450 ;
        RECT 133.950 694.950 136.050 695.400 ;
        RECT 127.950 673.950 130.050 676.050 ;
        RECT 128.400 673.050 129.450 673.950 ;
        RECT 121.950 670.950 124.050 673.050 ;
        RECT 125.250 671.250 126.750 672.150 ;
        RECT 127.950 670.950 130.050 673.050 ;
        RECT 121.950 668.850 123.750 669.750 ;
        RECT 124.950 667.950 127.050 670.050 ;
        RECT 128.250 668.850 129.750 669.750 ;
        RECT 130.950 667.950 133.050 670.050 ;
        RECT 97.950 658.950 100.050 661.050 ;
        RECT 55.950 632.250 58.050 633.150 ;
        RECT 107.400 631.050 108.450 665.400 ;
        RECT 109.950 664.950 112.050 665.400 ;
        RECT 115.950 665.400 120.450 666.450 ;
        RECT 115.950 664.950 118.050 665.400 ;
        RECT 116.400 637.050 117.450 664.950 ;
        RECT 118.950 661.950 121.050 664.050 ;
        RECT 115.950 634.950 118.050 637.050 ;
        RECT 55.950 630.450 58.050 631.050 ;
        RECT 53.400 629.400 58.050 630.450 ;
        RECT 55.950 628.950 58.050 629.400 ;
        RECT 67.950 630.450 70.050 631.050 ;
        RECT 67.950 629.400 72.450 630.450 ;
        RECT 67.950 628.950 70.050 629.400 ;
        RECT 31.950 619.500 34.050 621.600 ;
        RECT 36.150 619.500 38.250 621.600 ;
        RECT 40.950 619.500 43.050 621.600 ;
        RECT 43.950 619.500 46.050 621.600 ;
        RECT 46.950 619.500 49.050 621.600 ;
        RECT 16.950 604.950 19.050 607.050 ;
        RECT 19.950 604.950 22.050 607.050 ;
        RECT 22.950 604.950 25.050 607.050 ;
        RECT 31.950 605.400 34.050 607.500 ;
        RECT 36.150 605.400 38.250 607.500 ;
        RECT 40.950 605.400 43.050 607.500 ;
        RECT 43.950 605.400 46.050 607.500 ;
        RECT 46.950 605.400 49.050 607.500 ;
        RECT 7.950 598.950 10.050 601.050 ;
        RECT 4.950 596.250 7.050 597.150 ;
        RECT 4.950 594.450 7.050 595.050 ;
        RECT 8.400 594.450 9.450 598.950 ;
        RECT 4.950 593.400 9.450 594.450 ;
        RECT 10.950 593.850 13.050 594.750 ;
        RECT 4.950 592.950 7.050 593.400 ;
        RECT 17.550 586.050 18.750 604.950 ;
        RECT 20.550 592.350 21.750 604.950 ;
        RECT 19.950 590.250 22.050 592.350 ;
        RECT 20.550 586.050 21.750 590.250 ;
        RECT 23.550 586.050 24.750 604.950 ;
        RECT 28.950 601.950 31.050 604.050 ;
        RECT 28.950 599.850 31.050 600.750 ;
        RECT 32.250 596.850 33.450 605.400 ;
        RECT 36.450 599.550 37.650 605.400 ;
        RECT 36.150 597.450 38.250 599.550 ;
        RECT 31.950 594.750 34.050 596.850 ;
        RECT 32.250 588.600 33.450 594.750 ;
        RECT 36.450 588.600 37.650 597.450 ;
        RECT 41.400 591.750 42.600 605.400 ;
        RECT 40.950 589.650 43.050 591.750 ;
        RECT 31.950 586.500 34.050 588.600 ;
        RECT 36.000 586.500 38.100 588.600 ;
        RECT 44.550 588.150 45.750 605.400 ;
        RECT 47.250 591.750 48.450 605.400 ;
        RECT 56.400 598.050 57.450 628.950 ;
        RECT 67.950 626.850 70.050 627.750 ;
        RECT 71.400 625.050 72.450 629.400 ;
        RECT 79.950 629.250 82.050 630.150 ;
        RECT 85.950 629.250 88.050 630.150 ;
        RECT 94.950 628.950 97.050 631.050 ;
        RECT 106.950 628.950 109.050 631.050 ;
        RECT 115.950 628.950 118.050 631.050 ;
        RECT 79.950 625.950 82.050 628.050 ;
        RECT 83.250 626.250 84.750 627.150 ;
        RECT 85.950 625.950 88.050 628.050 ;
        RECT 94.950 626.850 97.050 627.750 ;
        RECT 97.950 626.250 100.050 627.150 ;
        RECT 106.950 626.850 109.050 627.750 ;
        RECT 109.950 626.250 112.050 627.150 ;
        RECT 112.950 626.250 115.050 627.150 ;
        RECT 115.950 626.850 118.050 627.750 ;
        RECT 70.950 622.950 73.050 625.050 ;
        RECT 80.400 601.050 81.450 625.950 ;
        RECT 119.400 625.050 120.450 661.950 ;
        RECT 125.400 655.050 126.450 667.950 ;
        RECT 134.400 667.050 135.450 694.950 ;
        RECT 137.400 673.050 138.450 697.950 ;
        RECT 136.950 670.950 139.050 673.050 ;
        RECT 139.950 668.250 141.750 669.150 ;
        RECT 142.950 667.950 145.050 670.050 ;
        RECT 146.250 668.250 148.050 669.150 ;
        RECT 130.950 665.850 133.050 666.750 ;
        RECT 133.950 664.950 136.050 667.050 ;
        RECT 139.950 664.950 142.050 667.050 ;
        RECT 143.250 665.850 144.750 666.750 ;
        RECT 145.950 666.450 148.050 667.050 ;
        RECT 149.400 666.450 150.450 733.950 ;
        RECT 155.400 733.050 156.450 739.950 ;
        RECT 157.950 736.950 160.050 739.050 ;
        RECT 154.950 730.950 157.050 733.050 ;
        RECT 158.400 718.050 159.450 736.950 ;
        RECT 167.400 721.050 168.450 739.950 ;
        RECT 178.950 737.850 181.050 738.750 ;
        RECT 166.950 718.950 169.050 721.050 ;
        RECT 157.950 715.950 160.050 718.050 ;
        RECT 158.400 706.050 159.450 715.950 ;
        RECT 169.950 709.950 172.050 712.050 ;
        RECT 178.950 709.950 181.050 712.050 ;
        RECT 163.950 707.250 166.050 708.150 ;
        RECT 157.950 703.950 160.050 706.050 ;
        RECT 161.250 704.250 162.750 705.150 ;
        RECT 163.950 703.950 166.050 706.050 ;
        RECT 167.250 704.250 169.050 705.150 ;
        RECT 157.950 701.850 159.750 702.750 ;
        RECT 160.950 700.950 163.050 703.050 ;
        RECT 161.400 700.050 162.450 700.950 ;
        RECT 164.400 700.050 165.450 703.950 ;
        RECT 166.950 700.950 169.050 703.050 ;
        RECT 160.950 697.950 163.050 700.050 ;
        RECT 163.950 697.950 166.050 700.050 ;
        RECT 167.400 685.050 168.450 700.950 ;
        RECT 166.950 682.950 169.050 685.050 ;
        RECT 170.400 679.050 171.450 709.950 ;
        RECT 179.400 706.050 180.450 709.950 ;
        RECT 178.950 703.950 181.050 706.050 ;
        RECT 175.950 701.250 178.050 702.150 ;
        RECT 178.950 701.850 181.050 702.750 ;
        RECT 182.400 700.050 183.450 761.400 ;
        RECT 185.400 739.050 186.450 763.950 ;
        RECT 187.950 749.400 190.050 751.500 ;
        RECT 190.950 749.400 193.050 751.500 ;
        RECT 193.950 749.400 196.050 751.500 ;
        RECT 198.750 749.400 200.850 751.500 ;
        RECT 202.950 749.400 205.050 751.500 ;
        RECT 184.950 736.950 187.050 739.050 ;
        RECT 188.550 735.750 189.750 749.400 ;
        RECT 187.950 733.650 190.050 735.750 ;
        RECT 188.550 729.900 189.750 733.650 ;
        RECT 191.250 732.150 192.450 749.400 ;
        RECT 194.400 735.750 195.600 749.400 ;
        RECT 199.350 743.550 200.550 749.400 ;
        RECT 198.750 741.450 200.850 743.550 ;
        RECT 193.950 733.650 196.050 735.750 ;
        RECT 199.350 732.600 200.550 741.450 ;
        RECT 203.550 740.850 204.750 749.400 ;
        RECT 205.950 745.950 208.050 748.050 ;
        RECT 205.950 743.850 208.050 744.750 ;
        RECT 202.950 738.750 205.050 740.850 ;
        RECT 203.550 732.600 204.750 738.750 ;
        RECT 209.400 733.050 210.450 770.400 ;
        RECT 218.400 766.050 219.450 808.950 ;
        RECT 227.400 790.050 228.450 818.400 ;
        RECT 229.950 817.950 232.050 818.400 ;
        RECT 241.950 817.950 244.050 820.050 ;
        RECT 256.950 817.950 259.050 820.050 ;
        RECT 259.950 817.950 262.050 820.050 ;
        RECT 257.400 817.050 258.450 817.950 ;
        RECT 229.950 815.850 232.050 816.750 ;
        RECT 232.950 815.250 235.050 816.150 ;
        RECT 235.950 814.950 238.050 817.050 ;
        RECT 241.950 815.850 244.050 816.750 ;
        RECT 244.950 815.250 247.050 816.150 ;
        RECT 256.950 814.950 259.050 817.050 ;
        RECT 260.250 815.850 261.750 816.750 ;
        RECT 262.950 816.450 265.050 817.050 ;
        RECT 262.950 815.400 267.450 816.450 ;
        RECT 262.950 814.950 265.050 815.400 ;
        RECT 232.950 813.450 235.050 814.050 ;
        RECT 236.400 813.450 237.450 814.950 ;
        RECT 232.950 812.400 237.450 813.450 ;
        RECT 232.950 811.950 235.050 812.400 ;
        RECT 244.950 811.950 247.050 814.050 ;
        RECT 256.950 812.850 259.050 813.750 ;
        RECT 262.950 812.850 265.050 813.750 ;
        RECT 266.400 808.050 267.450 815.400 ;
        RECT 275.400 814.050 276.450 820.950 ;
        RECT 271.950 812.250 274.050 813.150 ;
        RECT 274.950 811.950 277.050 814.050 ;
        RECT 271.950 808.950 274.050 811.050 ;
        RECT 272.400 808.050 273.450 808.950 ;
        RECT 265.950 805.950 268.050 808.050 ;
        RECT 271.950 805.950 274.050 808.050 ;
        RECT 226.950 787.950 229.050 790.050 ;
        RECT 235.950 787.950 238.050 790.050 ;
        RECT 226.950 784.950 229.050 787.050 ;
        RECT 229.950 784.950 232.050 787.050 ;
        RECT 232.950 784.950 235.050 787.050 ;
        RECT 220.950 776.250 223.050 777.150 ;
        RECT 223.950 775.950 226.050 778.050 ;
        RECT 217.950 763.950 220.050 766.050 ;
        RECT 211.950 748.950 214.050 751.050 ;
        RECT 214.950 748.950 217.050 751.050 ;
        RECT 217.950 748.950 220.050 751.050 ;
        RECT 190.950 730.050 193.050 732.150 ;
        RECT 198.900 730.500 201.000 732.600 ;
        RECT 202.950 730.500 205.050 732.600 ;
        RECT 208.950 730.950 211.050 733.050 ;
        RECT 212.250 730.050 213.450 748.950 ;
        RECT 215.250 736.350 216.450 748.950 ;
        RECT 214.950 734.250 217.050 736.350 ;
        RECT 215.250 730.050 216.450 734.250 ;
        RECT 218.250 730.050 219.450 748.950 ;
        RECT 224.400 742.050 225.450 775.950 ;
        RECT 227.550 766.050 228.750 784.950 ;
        RECT 230.550 780.750 231.750 784.950 ;
        RECT 229.950 778.650 232.050 780.750 ;
        RECT 230.550 766.050 231.750 778.650 ;
        RECT 233.550 766.050 234.750 784.950 ;
        RECT 226.950 763.950 229.050 766.050 ;
        RECT 229.950 763.950 232.050 766.050 ;
        RECT 232.950 763.950 235.050 766.050 ;
        RECT 236.400 745.050 237.450 787.950 ;
        RECT 257.100 785.100 259.200 787.200 ;
        RECT 241.950 782.400 244.050 784.500 ;
        RECT 246.000 782.400 248.100 784.500 ;
        RECT 253.950 782.850 256.050 784.950 ;
        RECT 242.250 776.250 243.450 782.400 ;
        RECT 241.950 774.150 244.050 776.250 ;
        RECT 238.950 770.250 241.050 771.150 ;
        RECT 238.950 766.950 241.050 769.050 ;
        RECT 242.250 765.600 243.450 774.150 ;
        RECT 246.450 773.550 247.650 782.400 ;
        RECT 250.950 779.250 253.050 781.350 ;
        RECT 246.150 771.450 248.250 773.550 ;
        RECT 246.450 765.600 247.650 771.450 ;
        RECT 251.400 765.600 252.600 779.250 ;
        RECT 254.550 765.600 255.750 782.850 ;
        RECT 257.250 781.350 258.450 785.100 ;
        RECT 256.950 779.250 259.050 781.350 ;
        RECT 257.250 765.600 258.450 779.250 ;
        RECT 272.400 778.050 273.450 805.950 ;
        RECT 265.950 776.250 268.050 777.150 ;
        RECT 271.950 775.950 274.050 778.050 ;
        RECT 265.950 772.950 268.050 775.050 ;
        RECT 266.400 772.050 267.450 772.950 ;
        RECT 265.950 769.950 268.050 772.050 ;
        RECT 241.950 763.500 244.050 765.600 ;
        RECT 246.150 763.500 248.250 765.600 ;
        RECT 250.950 763.500 253.050 765.600 ;
        RECT 253.950 763.500 256.050 765.600 ;
        RECT 256.950 763.500 259.050 765.600 ;
        RECT 266.400 757.050 267.450 769.950 ;
        RECT 265.950 754.950 268.050 757.050 ;
        RECT 238.950 751.950 241.050 754.050 ;
        RECT 244.950 751.950 247.050 754.050 ;
        RECT 235.950 742.950 238.050 745.050 ;
        RECT 223.950 739.950 226.050 742.050 ;
        RECT 229.950 740.250 232.050 741.150 ;
        RECT 223.950 737.850 226.050 738.750 ;
        RECT 187.800 727.800 189.900 729.900 ;
        RECT 211.950 727.950 214.050 730.050 ;
        RECT 214.950 727.950 217.050 730.050 ;
        RECT 217.950 727.950 220.050 730.050 ;
        RECT 220.950 718.950 223.050 721.050 ;
        RECT 187.950 715.950 190.050 718.050 ;
        RECT 188.400 709.050 189.450 715.950 ;
        RECT 208.950 712.950 211.050 715.050 ;
        RECT 214.950 712.950 217.050 715.050 ;
        RECT 187.950 706.950 190.050 709.050 ;
        RECT 184.950 701.250 187.050 702.150 ;
        RECT 175.950 697.950 178.050 700.050 ;
        RECT 181.950 697.950 184.050 700.050 ;
        RECT 184.950 697.950 187.050 700.050 ;
        RECT 188.400 699.450 189.450 706.950 ;
        RECT 209.400 706.050 210.450 712.950 ;
        RECT 208.950 703.950 211.050 706.050 ;
        RECT 190.950 701.250 193.050 702.150 ;
        RECT 196.950 701.250 199.050 702.150 ;
        RECT 205.950 701.250 208.050 702.150 ;
        RECT 190.950 699.450 193.050 700.050 ;
        RECT 188.400 698.400 193.050 699.450 ;
        RECT 185.400 697.050 186.450 697.950 ;
        RECT 184.950 694.950 187.050 697.050 ;
        RECT 188.400 690.450 189.450 698.400 ;
        RECT 190.950 697.950 193.050 698.400 ;
        RECT 194.250 698.250 195.750 699.150 ;
        RECT 196.950 697.950 199.050 700.050 ;
        RECT 205.950 699.450 208.050 700.050 ;
        RECT 209.400 699.450 210.450 703.950 ;
        RECT 211.950 701.250 214.050 702.150 ;
        RECT 205.950 698.400 210.450 699.450 ;
        RECT 211.950 699.450 214.050 700.050 ;
        RECT 215.400 699.450 216.450 712.950 ;
        RECT 217.950 703.950 220.050 706.050 ;
        RECT 217.950 701.850 220.050 702.750 ;
        RECT 211.950 698.400 216.450 699.450 ;
        RECT 205.950 697.950 208.050 698.400 ;
        RECT 211.950 697.950 214.050 698.400 ;
        RECT 217.950 697.950 220.050 700.050 ;
        RECT 193.950 694.950 196.050 697.050 ;
        RECT 185.400 689.400 189.450 690.450 ;
        RECT 157.950 676.950 160.050 679.050 ;
        RECT 169.950 676.950 172.050 679.050 ;
        RECT 158.400 673.050 159.450 676.950 ;
        RECT 160.950 673.950 163.050 676.050 ;
        RECT 169.950 673.950 172.050 676.050 ;
        RECT 181.950 673.950 184.050 676.050 ;
        RECT 157.950 670.950 160.050 673.050 ;
        RECT 161.250 671.850 162.750 672.750 ;
        RECT 163.950 670.950 166.050 673.050 ;
        RECT 166.950 670.950 169.050 673.050 ;
        RECT 157.950 668.850 160.050 669.750 ;
        RECT 163.950 668.850 166.050 669.750 ;
        RECT 145.950 665.400 150.450 666.450 ;
        RECT 145.950 664.950 148.050 665.400 ;
        RECT 134.400 664.050 135.450 664.950 ;
        RECT 133.950 661.950 136.050 664.050 ;
        RECT 146.400 663.450 147.450 664.950 ;
        RECT 143.400 662.400 147.450 663.450 ;
        RECT 143.400 661.050 144.450 662.400 ;
        RECT 142.950 658.950 145.050 661.050 ;
        RECT 124.950 652.950 127.050 655.050 ;
        RECT 124.950 649.950 127.050 652.050 ;
        RECT 82.950 622.950 85.050 625.050 ;
        RECT 97.950 622.950 100.050 625.050 ;
        RECT 109.950 622.950 112.050 625.050 ;
        RECT 112.950 622.950 115.050 625.050 ;
        RECT 118.950 622.950 121.050 625.050 ;
        RECT 83.400 622.050 84.450 622.950 ;
        RECT 82.950 619.950 85.050 622.050 ;
        RECT 82.950 601.950 85.050 604.050 ;
        RECT 85.950 601.950 88.050 604.050 ;
        RECT 91.950 603.450 94.050 604.050 ;
        RECT 89.400 602.400 94.050 603.450 ;
        RECT 86.400 601.050 87.450 601.950 ;
        RECT 67.950 599.250 70.050 600.150 ;
        RECT 79.950 598.950 82.050 601.050 ;
        RECT 83.250 599.850 84.750 600.750 ;
        RECT 85.950 598.950 88.050 601.050 ;
        RECT 89.400 598.050 90.450 602.400 ;
        RECT 91.950 601.950 94.050 602.400 ;
        RECT 91.950 599.850 94.050 600.750 ;
        RECT 94.950 599.250 97.050 600.150 ;
        RECT 55.950 595.950 58.050 598.050 ;
        RECT 67.950 595.950 70.050 598.050 ;
        RECT 79.950 596.850 82.050 597.750 ;
        RECT 85.950 596.850 88.050 597.750 ;
        RECT 88.950 595.950 91.050 598.050 ;
        RECT 94.950 595.950 97.050 598.050 ;
        RECT 55.950 593.850 58.050 594.750 ;
        RECT 91.950 594.450 94.050 595.050 ;
        RECT 95.400 594.450 96.450 595.950 ;
        RECT 91.950 593.400 96.450 594.450 ;
        RECT 91.950 592.950 94.050 593.400 ;
        RECT 46.950 589.650 49.050 591.750 ;
        RECT 43.950 586.050 46.050 588.150 ;
        RECT 16.950 583.950 19.050 586.050 ;
        RECT 19.950 583.950 22.050 586.050 ;
        RECT 22.950 583.950 25.050 586.050 ;
        RECT 47.250 585.900 48.450 589.650 ;
        RECT 47.100 583.800 49.200 585.900 ;
        RECT 82.950 565.950 85.050 568.050 ;
        RECT 94.950 565.950 97.050 568.050 ;
        RECT 19.950 563.250 22.050 564.150 ;
        RECT 34.950 563.250 37.050 564.150 ;
        RECT 16.950 560.250 18.750 561.150 ;
        RECT 19.950 559.950 22.050 562.050 ;
        RECT 25.950 561.450 28.050 562.050 ;
        RECT 23.250 560.250 24.750 561.150 ;
        RECT 25.950 560.400 30.450 561.450 ;
        RECT 25.950 559.950 28.050 560.400 ;
        RECT 4.950 558.450 7.050 559.050 ;
        RECT 2.400 557.400 7.050 558.450 ;
        RECT 2.400 553.050 3.450 557.400 ;
        RECT 4.950 556.950 7.050 557.400 ;
        RECT 16.950 556.950 19.050 559.050 ;
        RECT 22.950 556.950 25.050 559.050 ;
        RECT 26.250 557.850 28.050 558.750 ;
        RECT 4.950 554.850 7.050 555.750 ;
        RECT 7.950 554.250 10.050 555.150 ;
        RECT 1.950 550.950 4.050 553.050 ;
        RECT 7.950 550.950 10.050 553.050 ;
        RECT 8.400 544.050 9.450 550.950 ;
        RECT 17.400 544.050 18.450 556.950 ;
        RECT 29.400 556.050 30.450 560.400 ;
        RECT 31.950 560.250 33.750 561.150 ;
        RECT 34.950 559.950 37.050 562.050 ;
        RECT 38.250 560.250 39.750 561.150 ;
        RECT 40.950 559.950 43.050 562.050 ;
        RECT 31.950 556.950 34.050 559.050 ;
        RECT 28.950 553.950 31.050 556.050 ;
        RECT 32.400 553.050 33.450 556.950 ;
        RECT 31.950 550.950 34.050 553.050 ;
        RECT 32.400 550.050 33.450 550.950 ;
        RECT 31.950 547.950 34.050 550.050 ;
        RECT 7.950 541.950 10.050 544.050 ;
        RECT 16.950 541.950 19.050 544.050 ;
        RECT 25.950 529.950 28.050 532.050 ;
        RECT 10.950 526.950 13.050 529.050 ;
        RECT 11.400 526.050 12.450 526.950 ;
        RECT 7.950 524.250 9.750 525.150 ;
        RECT 10.950 523.950 13.050 526.050 ;
        RECT 14.250 524.250 16.050 525.150 ;
        RECT 16.950 523.950 19.050 526.050 ;
        RECT 19.950 524.250 21.750 525.150 ;
        RECT 22.950 523.950 25.050 526.050 ;
        RECT 7.950 520.950 10.050 523.050 ;
        RECT 11.250 521.850 12.750 522.750 ;
        RECT 13.950 520.950 16.050 523.050 ;
        RECT 8.400 514.050 9.450 520.950 ;
        RECT 14.400 517.050 15.450 520.950 ;
        RECT 13.950 514.950 16.050 517.050 ;
        RECT 7.950 511.950 10.050 514.050 ;
        RECT 13.950 511.950 16.050 514.050 ;
        RECT 7.950 487.950 10.050 490.050 ;
        RECT 8.400 487.050 9.450 487.950 ;
        RECT 7.950 484.950 10.050 487.050 ;
        RECT 7.950 482.850 10.050 483.750 ;
        RECT 10.950 482.250 13.050 483.150 ;
        RECT 10.950 478.950 13.050 481.050 ;
        RECT 14.400 480.450 15.450 511.950 ;
        RECT 17.400 505.050 18.450 523.950 ;
        RECT 26.400 523.050 27.450 529.950 ;
        RECT 28.950 526.950 31.050 529.050 ;
        RECT 29.400 526.050 30.450 526.950 ;
        RECT 28.950 523.950 31.050 526.050 ;
        RECT 35.400 523.050 36.450 559.950 ;
        RECT 37.950 556.950 40.050 559.050 ;
        RECT 41.250 557.850 43.050 558.750 ;
        RECT 46.950 558.450 49.050 559.050 ;
        RECT 44.400 557.400 49.050 558.450 ;
        RECT 38.400 526.050 39.450 556.950 ;
        RECT 44.400 556.050 45.450 557.400 ;
        RECT 46.950 556.950 49.050 557.400 ;
        RECT 52.950 556.950 55.050 559.050 ;
        RECT 56.250 557.250 58.050 558.150 ;
        RECT 70.950 556.950 73.050 559.050 ;
        RECT 76.950 557.250 79.050 558.150 ;
        RECT 43.950 553.950 46.050 556.050 ;
        RECT 46.950 554.850 49.050 555.750 ;
        RECT 49.950 554.250 52.050 555.150 ;
        RECT 52.950 554.850 54.750 555.750 ;
        RECT 55.950 553.950 58.050 556.050 ;
        RECT 70.950 554.850 73.050 555.750 ;
        RECT 76.950 553.950 79.050 556.050 ;
        RECT 80.250 554.250 82.050 555.150 ;
        RECT 49.950 550.950 52.050 553.050 ;
        RECT 43.950 529.950 46.050 532.050 ;
        RECT 44.400 526.050 45.450 529.950 ;
        RECT 37.950 523.950 40.050 526.050 ;
        RECT 40.950 524.250 42.750 525.150 ;
        RECT 43.950 523.950 46.050 526.050 ;
        RECT 47.250 524.250 49.050 525.150 ;
        RECT 19.950 520.950 22.050 523.050 ;
        RECT 23.250 521.850 24.750 522.750 ;
        RECT 25.950 520.950 28.050 523.050 ;
        RECT 29.250 521.850 31.050 522.750 ;
        RECT 34.950 520.950 37.050 523.050 ;
        RECT 40.950 520.950 43.050 523.050 ;
        RECT 44.250 521.850 45.750 522.750 ;
        RECT 46.950 520.950 49.050 523.050 ;
        RECT 41.400 520.050 42.450 520.950 ;
        RECT 25.950 518.850 28.050 519.750 ;
        RECT 40.950 517.950 43.050 520.050 ;
        RECT 22.950 514.950 25.050 517.050 ;
        RECT 16.950 502.950 19.050 505.050 ;
        RECT 19.950 485.250 22.050 486.150 ;
        RECT 23.400 484.050 24.450 514.950 ;
        RECT 25.950 502.950 28.050 505.050 ;
        RECT 26.400 487.050 27.450 502.950 ;
        RECT 47.400 502.050 48.450 520.950 ;
        RECT 50.400 517.050 51.450 550.950 ;
        RECT 56.400 535.050 57.450 553.950 ;
        RECT 77.400 553.050 78.450 553.950 ;
        RECT 76.950 550.950 79.050 553.050 ;
        RECT 79.950 552.450 82.050 553.050 ;
        RECT 83.400 552.450 84.450 565.950 ;
        RECT 95.400 562.050 96.450 565.950 ;
        RECT 88.950 561.450 91.050 562.050 ;
        RECT 86.400 560.400 91.050 561.450 ;
        RECT 86.400 553.050 87.450 560.400 ;
        RECT 88.950 559.950 91.050 560.400 ;
        RECT 92.250 560.250 93.750 561.150 ;
        RECT 94.950 559.950 97.050 562.050 ;
        RECT 88.950 557.850 90.750 558.750 ;
        RECT 91.950 556.950 94.050 559.050 ;
        RECT 95.250 557.850 97.050 558.750 ;
        RECT 79.950 551.400 84.450 552.450 ;
        RECT 79.950 550.950 82.050 551.400 ;
        RECT 85.950 550.950 88.050 553.050 ;
        RECT 55.950 532.950 58.050 535.050 ;
        RECT 92.400 532.050 93.450 556.950 ;
        RECT 98.400 541.050 99.450 622.950 ;
        RECT 100.950 619.950 103.050 622.050 ;
        RECT 101.400 568.050 102.450 619.950 ;
        RECT 125.400 619.050 126.450 649.950 ;
        RECT 139.950 631.950 142.050 634.050 ;
        RECT 127.950 628.950 130.050 631.050 ;
        RECT 130.950 629.250 133.050 630.150 ;
        RECT 136.950 629.250 139.050 630.150 ;
        RECT 128.400 627.450 129.450 628.950 ;
        RECT 130.950 627.450 133.050 628.050 ;
        RECT 128.400 626.400 133.050 627.450 ;
        RECT 136.950 627.450 139.050 628.050 ;
        RECT 140.400 627.450 141.450 631.950 ;
        RECT 143.400 631.050 144.450 658.950 ;
        RECT 160.950 652.950 163.050 655.050 ;
        RECT 161.400 634.050 162.450 652.950 ;
        RECT 167.400 636.450 168.450 670.950 ;
        RECT 170.400 667.050 171.450 673.950 ;
        RECT 182.400 673.050 183.450 673.950 ;
        RECT 172.950 670.950 175.050 673.050 ;
        RECT 178.950 670.950 181.050 673.050 ;
        RECT 181.950 670.950 184.050 673.050 ;
        RECT 172.950 668.850 175.050 669.750 ;
        RECT 175.950 668.250 178.050 669.150 ;
        RECT 169.950 664.950 172.050 667.050 ;
        RECT 175.950 664.950 178.050 667.050 ;
        RECT 175.950 661.950 178.050 664.050 ;
        RECT 164.400 635.400 168.450 636.450 ;
        RECT 148.950 631.950 151.050 634.050 ;
        RECT 154.950 632.250 157.050 633.150 ;
        RECT 157.950 631.950 160.050 634.050 ;
        RECT 160.950 631.950 163.050 634.050 ;
        RECT 149.400 631.050 150.450 631.950 ;
        RECT 142.950 628.950 145.050 631.050 ;
        RECT 145.950 629.250 147.750 630.150 ;
        RECT 148.950 628.950 151.050 631.050 ;
        RECT 152.250 629.250 153.750 630.150 ;
        RECT 154.950 628.950 157.050 631.050 ;
        RECT 130.950 625.950 133.050 626.400 ;
        RECT 134.250 626.250 135.750 627.150 ;
        RECT 136.950 626.400 141.450 627.450 ;
        RECT 136.950 625.950 139.050 626.400 ;
        RECT 145.950 625.950 148.050 628.050 ;
        RECT 149.250 626.850 150.750 627.750 ;
        RECT 151.950 625.950 154.050 628.050 ;
        RECT 127.950 622.950 130.050 625.050 ;
        RECT 133.950 622.950 136.050 625.050 ;
        RECT 128.400 619.050 129.450 622.950 ;
        RECT 109.950 616.950 112.050 619.050 ;
        RECT 124.950 616.950 127.050 619.050 ;
        RECT 127.950 616.950 130.050 619.050 ;
        RECT 110.400 601.050 111.450 616.950 ;
        RECT 112.950 613.950 115.050 616.050 ;
        RECT 113.400 604.050 114.450 613.950 ;
        RECT 134.400 613.050 135.450 622.950 ;
        RECT 151.950 616.950 154.050 619.050 ;
        RECT 152.400 613.050 153.450 616.950 ;
        RECT 124.950 610.950 127.050 613.050 ;
        RECT 133.950 610.950 136.050 613.050 ;
        RECT 151.950 610.950 154.050 613.050 ;
        RECT 118.950 607.950 121.050 610.050 ;
        RECT 112.950 601.950 115.050 604.050 ;
        RECT 103.950 598.950 106.050 601.050 ;
        RECT 106.950 598.950 109.050 601.050 ;
        RECT 109.950 598.950 112.050 601.050 ;
        RECT 103.950 596.850 106.050 597.750 ;
        RECT 100.950 565.950 103.050 568.050 ;
        RECT 107.400 565.050 108.450 598.950 ;
        RECT 109.950 596.850 112.050 597.750 ;
        RECT 106.950 562.950 109.050 565.050 ;
        RECT 109.950 559.950 112.050 562.050 ;
        RECT 100.950 557.250 103.050 558.150 ;
        RECT 106.950 557.250 109.050 558.150 ;
        RECT 100.950 553.950 103.050 556.050 ;
        RECT 104.250 554.250 105.750 555.150 ;
        RECT 106.950 553.950 109.050 556.050 ;
        RECT 101.400 547.050 102.450 553.950 ;
        RECT 103.950 550.950 106.050 553.050 ;
        RECT 103.950 547.950 106.050 550.050 ;
        RECT 100.950 544.950 103.050 547.050 ;
        RECT 97.950 538.950 100.050 541.050 ;
        RECT 91.950 529.950 94.050 532.050 ;
        RECT 85.950 526.950 88.050 529.050 ;
        RECT 88.950 526.950 91.050 529.050 ;
        RECT 55.950 523.950 58.050 526.050 ;
        RECT 58.950 524.250 60.750 525.150 ;
        RECT 61.950 523.950 64.050 526.050 ;
        RECT 67.950 525.450 70.050 526.050 ;
        RECT 67.950 524.400 72.450 525.450 ;
        RECT 67.950 523.950 70.050 524.400 ;
        RECT 56.400 522.450 57.450 523.950 ;
        RECT 58.950 522.450 61.050 523.050 ;
        RECT 56.400 521.400 61.050 522.450 ;
        RECT 62.250 521.850 63.750 522.750 ;
        RECT 58.950 520.950 61.050 521.400 ;
        RECT 64.950 520.950 67.050 523.050 ;
        RECT 68.250 521.850 70.050 522.750 ;
        RECT 71.400 520.050 72.450 524.400 ;
        RECT 73.950 524.250 75.750 525.150 ;
        RECT 76.950 523.950 79.050 526.050 ;
        RECT 80.250 524.250 82.050 525.150 ;
        RECT 82.950 523.950 85.050 526.050 ;
        RECT 73.950 520.950 76.050 523.050 ;
        RECT 77.250 521.850 78.750 522.750 ;
        RECT 79.950 520.950 82.050 523.050 ;
        RECT 80.400 520.050 81.450 520.950 ;
        RECT 64.950 518.850 67.050 519.750 ;
        RECT 70.950 517.950 73.050 520.050 ;
        RECT 79.950 517.950 82.050 520.050 ;
        RECT 49.950 514.950 52.050 517.050 ;
        RECT 46.950 499.950 49.050 502.050 ;
        RECT 64.950 499.950 67.050 502.050 ;
        RECT 37.950 488.250 40.050 489.150 ;
        RECT 55.950 487.950 58.050 490.050 ;
        RECT 61.950 488.250 64.050 489.150 ;
        RECT 56.400 487.050 57.450 487.950 ;
        RECT 25.950 484.950 28.050 487.050 ;
        RECT 37.950 484.950 40.050 487.050 ;
        RECT 41.250 485.250 42.750 486.150 ;
        RECT 43.950 484.950 46.050 487.050 ;
        RECT 47.250 485.250 49.050 486.150 ;
        RECT 49.950 484.950 52.050 487.050 ;
        RECT 52.950 485.250 54.750 486.150 ;
        RECT 55.950 484.950 58.050 487.050 ;
        RECT 59.250 485.250 60.750 486.150 ;
        RECT 61.950 484.950 64.050 487.050 ;
        RECT 16.950 482.250 18.750 483.150 ;
        RECT 19.950 481.950 22.050 484.050 ;
        RECT 22.950 481.950 25.050 484.050 ;
        RECT 25.950 482.850 28.050 483.750 ;
        RECT 16.950 480.450 19.050 481.050 ;
        RECT 14.400 479.400 19.050 480.450 ;
        RECT 16.950 478.950 19.050 479.400 ;
        RECT 11.400 457.050 12.450 478.950 ;
        RECT 10.950 454.950 13.050 457.050 ;
        RECT 11.400 454.050 12.450 454.950 ;
        RECT 7.950 452.250 9.750 453.150 ;
        RECT 10.950 451.950 13.050 454.050 ;
        RECT 14.250 452.250 16.050 453.150 ;
        RECT 7.950 448.950 10.050 451.050 ;
        RECT 11.250 449.850 12.750 450.750 ;
        RECT 13.950 448.950 16.050 451.050 ;
        RECT 8.400 448.050 9.450 448.950 ;
        RECT 7.950 445.950 10.050 448.050 ;
        RECT 7.950 439.950 10.050 442.050 ;
        RECT 8.400 415.050 9.450 439.950 ;
        RECT 7.950 412.950 10.050 415.050 ;
        RECT 14.400 412.050 15.450 448.950 ;
        RECT 17.400 442.050 18.450 478.950 ;
        RECT 25.950 475.950 28.050 478.050 ;
        RECT 26.400 460.050 27.450 475.950 ;
        RECT 25.950 457.950 28.050 460.050 ;
        RECT 38.400 457.050 39.450 484.950 ;
        RECT 40.950 481.950 43.050 484.050 ;
        RECT 44.250 482.850 45.750 483.750 ;
        RECT 46.950 481.950 49.050 484.050 ;
        RECT 47.400 481.050 48.450 481.950 ;
        RECT 46.950 478.950 49.050 481.050 ;
        RECT 50.400 478.050 51.450 484.950 ;
        RECT 52.950 481.950 55.050 484.050 ;
        RECT 56.250 482.850 57.750 483.750 ;
        RECT 58.950 481.950 61.050 484.050 ;
        RECT 53.400 478.050 54.450 481.950 ;
        RECT 62.400 481.050 63.450 484.950 ;
        RECT 65.400 484.050 66.450 499.950 ;
        RECT 71.400 487.050 72.450 517.950 ;
        RECT 80.400 505.050 81.450 517.950 ;
        RECT 79.950 502.950 82.050 505.050 ;
        RECT 83.400 493.050 84.450 523.950 ;
        RECT 86.400 523.050 87.450 526.950 ;
        RECT 89.400 526.050 90.450 526.950 ;
        RECT 104.400 526.050 105.450 547.950 ;
        RECT 110.400 529.050 111.450 559.950 ;
        RECT 113.400 547.050 114.450 601.950 ;
        RECT 119.400 601.050 120.450 607.950 ;
        RECT 121.950 604.950 124.050 607.050 ;
        RECT 122.400 604.050 123.450 604.950 ;
        RECT 121.950 601.950 124.050 604.050 ;
        RECT 125.400 601.050 126.450 610.950 ;
        RECT 134.400 607.050 135.450 610.950 ;
        RECT 136.950 607.950 139.050 610.050 ;
        RECT 145.950 607.950 148.050 610.050 ;
        RECT 127.950 604.950 130.050 607.050 ;
        RECT 133.950 604.950 136.050 607.050 ;
        RECT 118.950 600.450 121.050 601.050 ;
        RECT 116.400 599.400 121.050 600.450 ;
        RECT 122.250 599.850 123.750 600.750 ;
        RECT 116.400 562.050 117.450 599.400 ;
        RECT 118.950 598.950 121.050 599.400 ;
        RECT 124.950 598.950 127.050 601.050 ;
        RECT 118.950 596.850 121.050 597.750 ;
        RECT 124.950 596.850 127.050 597.750 ;
        RECT 128.400 592.050 129.450 604.950 ;
        RECT 137.400 604.050 138.450 607.950 ;
        RECT 139.950 604.950 142.050 607.050 ;
        RECT 140.400 604.050 141.450 604.950 ;
        RECT 133.950 601.950 136.050 604.050 ;
        RECT 136.950 601.950 139.050 604.050 ;
        RECT 139.950 601.950 142.050 604.050 ;
        RECT 137.400 601.050 138.450 601.950 ;
        RECT 146.400 601.050 147.450 607.950 ;
        RECT 152.400 601.050 153.450 610.950 ;
        RECT 155.400 610.050 156.450 628.950 ;
        RECT 158.400 625.050 159.450 631.950 ;
        RECT 160.950 628.950 163.050 631.050 ;
        RECT 157.950 622.950 160.050 625.050 ;
        RECT 154.950 607.950 157.050 610.050 ;
        RECT 154.950 601.950 157.050 604.050 ;
        RECT 130.950 598.950 133.050 601.050 ;
        RECT 134.250 599.850 135.750 600.750 ;
        RECT 136.950 598.950 139.050 601.050 ;
        RECT 139.950 599.850 142.050 600.750 ;
        RECT 142.950 599.250 145.050 600.150 ;
        RECT 145.950 598.950 148.050 601.050 ;
        RECT 151.950 598.950 154.050 601.050 ;
        RECT 155.250 599.850 156.750 600.750 ;
        RECT 157.950 598.950 160.050 601.050 ;
        RECT 130.950 596.850 133.050 597.750 ;
        RECT 136.950 596.850 139.050 597.750 ;
        RECT 142.950 595.950 145.050 598.050 ;
        RECT 136.950 592.950 139.050 595.050 ;
        RECT 127.950 589.950 130.050 592.050 ;
        RECT 118.950 562.950 121.050 565.050 ;
        RECT 115.950 559.950 118.050 562.050 ;
        RECT 112.950 544.950 115.050 547.050 ;
        RECT 109.950 526.950 112.050 529.050 ;
        RECT 88.950 523.950 91.050 526.050 ;
        RECT 94.950 523.950 97.050 526.050 ;
        RECT 98.250 524.250 100.050 525.150 ;
        RECT 100.950 523.950 103.050 526.050 ;
        RECT 103.950 523.950 106.050 526.050 ;
        RECT 109.950 523.950 112.050 526.050 ;
        RECT 113.250 524.250 115.050 525.150 ;
        RECT 115.950 523.950 118.050 526.050 ;
        RECT 85.950 520.950 88.050 523.050 ;
        RECT 88.950 521.850 90.750 522.750 ;
        RECT 91.950 520.950 94.050 523.050 ;
        RECT 95.250 521.850 96.750 522.750 ;
        RECT 97.950 520.950 100.050 523.050 ;
        RECT 91.950 518.850 94.050 519.750 ;
        RECT 101.400 519.450 102.450 523.950 ;
        RECT 103.950 521.850 105.750 522.750 ;
        RECT 106.950 520.950 109.050 523.050 ;
        RECT 110.250 521.850 111.750 522.750 ;
        RECT 112.950 520.950 115.050 523.050 ;
        RECT 98.400 518.400 102.450 519.450 ;
        RECT 106.950 518.850 109.050 519.750 ;
        RECT 82.950 490.950 85.050 493.050 ;
        RECT 91.950 491.250 94.050 492.150 ;
        RECT 98.400 490.050 99.450 518.400 ;
        RECT 113.400 517.050 114.450 520.950 ;
        RECT 112.950 514.950 115.050 517.050 ;
        RECT 116.400 499.050 117.450 523.950 ;
        RECT 115.950 496.950 118.050 499.050 ;
        RECT 119.400 496.050 120.450 562.950 ;
        RECT 124.950 559.950 127.050 562.050 ;
        RECT 121.950 557.250 124.050 558.150 ;
        RECT 124.950 557.850 127.050 558.750 ;
        RECT 121.950 553.950 124.050 556.050 ;
        RECT 128.400 544.050 129.450 589.950 ;
        RECT 137.400 559.050 138.450 592.950 ;
        RECT 143.400 580.050 144.450 595.950 ;
        RECT 142.950 577.950 145.050 580.050 ;
        RECT 130.950 557.250 133.050 558.150 ;
        RECT 136.950 556.950 139.050 559.050 ;
        RECT 130.950 553.950 133.050 556.050 ;
        RECT 136.950 554.850 139.050 555.750 ;
        RECT 131.400 553.050 132.450 553.950 ;
        RECT 146.400 553.050 147.450 598.950 ;
        RECT 151.950 596.850 154.050 597.750 ;
        RECT 154.950 595.950 157.050 598.050 ;
        RECT 157.950 596.850 160.050 597.750 ;
        RECT 151.950 556.950 154.050 559.050 ;
        RECT 130.950 550.950 133.050 553.050 ;
        RECT 145.950 550.950 148.050 553.050 ;
        RECT 127.950 541.950 130.050 544.050 ;
        RECT 124.950 525.450 127.050 526.050 ;
        RECT 128.400 525.450 129.450 541.950 ;
        RECT 142.950 531.450 145.050 532.050 ;
        RECT 137.400 530.400 145.050 531.450 ;
        RECT 124.950 524.400 129.450 525.450 ;
        RECT 124.950 523.950 127.050 524.400 ;
        RECT 130.950 523.950 133.050 526.050 ;
        RECT 134.250 524.250 136.050 525.150 ;
        RECT 124.950 521.850 126.750 522.750 ;
        RECT 127.950 520.950 130.050 523.050 ;
        RECT 131.250 521.850 132.750 522.750 ;
        RECT 133.950 522.450 136.050 523.050 ;
        RECT 137.400 522.450 138.450 530.400 ;
        RECT 142.950 529.950 145.050 530.400 ;
        RECT 139.950 527.250 142.050 528.150 ;
        RECT 142.950 527.850 145.050 528.750 ;
        RECT 145.950 527.250 147.750 528.150 ;
        RECT 148.950 526.950 151.050 529.050 ;
        RECT 139.950 523.950 142.050 526.050 ;
        RECT 145.950 523.950 148.050 526.050 ;
        RECT 149.250 524.850 151.050 525.750 ;
        RECT 133.950 521.400 138.450 522.450 ;
        RECT 133.950 520.950 136.050 521.400 ;
        RECT 127.950 518.850 130.050 519.750 ;
        RECT 152.400 505.050 153.450 556.950 ;
        RECT 155.400 514.050 156.450 595.950 ;
        RECT 157.950 554.850 160.050 555.750 ;
        RECT 161.400 550.050 162.450 628.950 ;
        RECT 164.400 604.050 165.450 635.400 ;
        RECT 172.950 634.950 175.050 637.050 ;
        RECT 173.400 634.050 174.450 634.950 ;
        RECT 166.950 631.950 169.050 634.050 ;
        RECT 170.250 632.250 171.750 633.150 ;
        RECT 172.950 631.950 175.050 634.050 ;
        RECT 166.950 629.850 168.750 630.750 ;
        RECT 169.950 628.950 172.050 631.050 ;
        RECT 173.250 629.850 175.050 630.750 ;
        RECT 170.400 627.450 171.450 628.950 ;
        RECT 167.400 626.400 171.450 627.450 ;
        RECT 163.950 601.950 166.050 604.050 ;
        RECT 160.950 547.950 163.050 550.050 ;
        RECT 164.400 547.050 165.450 601.950 ;
        RECT 163.950 544.950 166.050 547.050 ;
        RECT 160.950 532.950 163.050 535.050 ;
        RECT 161.400 526.050 162.450 532.950 ;
        RECT 163.950 526.950 166.050 529.050 ;
        RECT 160.950 523.950 163.050 526.050 ;
        RECT 163.950 524.850 166.050 525.750 ;
        RECT 154.950 511.950 157.050 514.050 ;
        RECT 167.400 511.050 168.450 626.400 ;
        RECT 176.400 598.050 177.450 661.950 ;
        RECT 179.400 655.050 180.450 670.950 ;
        RECT 181.950 668.850 184.050 669.750 ;
        RECT 178.950 652.950 181.050 655.050 ;
        RECT 185.400 639.450 186.450 689.400 ;
        RECT 190.950 685.950 193.050 688.050 ;
        RECT 191.400 670.050 192.450 685.950 ;
        RECT 194.400 676.050 195.450 694.950 ;
        RECT 193.950 673.950 196.050 676.050 ;
        RECT 193.950 670.950 196.050 673.050 ;
        RECT 199.950 672.450 202.050 673.050 ;
        RECT 212.400 672.450 213.450 697.950 ;
        RECT 218.400 678.450 219.450 697.950 ;
        RECT 221.400 697.050 222.450 718.950 ;
        RECT 229.950 712.950 232.050 715.050 ;
        RECT 232.950 712.950 235.050 715.050 ;
        RECT 235.950 712.950 238.050 715.050 ;
        RECT 223.950 704.250 226.050 705.150 ;
        RECT 226.950 700.950 229.050 703.050 ;
        RECT 220.950 694.950 223.050 697.050 ;
        RECT 197.250 671.250 198.750 672.150 ;
        RECT 199.950 671.400 204.450 672.450 ;
        RECT 199.950 670.950 202.050 671.400 ;
        RECT 190.950 667.950 193.050 670.050 ;
        RECT 194.250 668.850 195.750 669.750 ;
        RECT 196.950 667.950 199.050 670.050 ;
        RECT 200.250 668.850 202.050 669.750 ;
        RECT 203.400 667.050 204.450 671.400 ;
        RECT 209.400 671.400 213.450 672.450 ;
        RECT 215.400 677.400 219.450 678.450 ;
        RECT 190.950 665.850 193.050 666.750 ;
        RECT 202.950 664.950 205.050 667.050 ;
        RECT 209.400 652.050 210.450 671.400 ;
        RECT 215.400 670.050 216.450 677.400 ;
        RECT 217.950 673.950 220.050 676.050 ;
        RECT 211.950 668.250 213.750 669.150 ;
        RECT 214.950 667.950 217.050 670.050 ;
        RECT 218.400 667.050 219.450 673.950 ;
        RECT 221.400 670.050 222.450 694.950 ;
        RECT 227.400 691.050 228.450 700.950 ;
        RECT 230.550 694.050 231.750 712.950 ;
        RECT 233.550 708.750 234.750 712.950 ;
        RECT 232.950 706.650 235.050 708.750 ;
        RECT 233.550 694.050 234.750 706.650 ;
        RECT 236.550 694.050 237.750 712.950 ;
        RECT 239.400 700.050 240.450 751.950 ;
        RECT 245.400 748.050 246.450 751.950 ;
        RECT 247.950 748.950 250.050 751.050 ;
        RECT 244.950 745.950 247.050 748.050 ;
        RECT 248.400 745.050 249.450 748.950 ;
        RECT 275.400 745.050 276.450 811.950 ;
        RECT 277.950 809.850 280.050 810.750 ;
        RECT 284.550 802.050 285.750 820.950 ;
        RECT 287.550 808.350 288.750 820.950 ;
        RECT 286.950 806.250 289.050 808.350 ;
        RECT 287.550 802.050 288.750 806.250 ;
        RECT 290.550 802.050 291.750 820.950 ;
        RECT 295.950 817.950 298.050 820.050 ;
        RECT 295.950 815.850 298.050 816.750 ;
        RECT 299.250 812.850 300.450 821.400 ;
        RECT 303.450 815.550 304.650 821.400 ;
        RECT 303.150 813.450 305.250 815.550 ;
        RECT 295.950 808.950 298.050 811.050 ;
        RECT 298.950 810.750 301.050 812.850 ;
        RECT 283.950 799.950 286.050 802.050 ;
        RECT 286.950 799.950 289.050 802.050 ;
        RECT 289.950 799.950 292.050 802.050 ;
        RECT 277.950 787.950 280.050 790.050 ;
        RECT 278.400 775.050 279.450 787.950 ;
        RECT 277.950 772.950 280.050 775.050 ;
        RECT 286.950 774.450 289.050 775.050 ;
        RECT 284.400 773.400 289.050 774.450 ;
        RECT 277.950 770.850 280.050 771.750 ;
        RECT 284.400 765.450 285.450 773.400 ;
        RECT 286.950 772.950 289.050 773.400 ;
        RECT 296.400 774.450 297.450 808.950 ;
        RECT 299.250 804.600 300.450 810.750 ;
        RECT 303.450 804.600 304.650 813.450 ;
        RECT 308.400 807.750 309.600 821.400 ;
        RECT 307.950 805.650 310.050 807.750 ;
        RECT 298.950 802.500 301.050 804.600 ;
        RECT 303.000 802.500 305.100 804.600 ;
        RECT 311.550 804.150 312.750 821.400 ;
        RECT 314.250 807.750 315.450 821.400 ;
        RECT 442.950 820.950 445.050 823.050 ;
        RECT 451.950 820.950 454.050 823.050 ;
        RECT 502.950 820.950 505.050 823.050 ;
        RECT 508.950 820.950 511.050 823.050 ;
        RECT 523.950 820.950 526.050 823.050 ;
        RECT 787.950 820.950 790.050 823.050 ;
        RECT 796.950 820.950 799.050 823.050 ;
        RECT 340.950 817.950 343.050 820.050 ;
        RECT 421.950 817.950 424.050 820.050 ;
        RECT 328.950 814.950 331.050 817.050 ;
        RECT 334.950 815.250 337.050 816.150 ;
        RECT 322.950 813.450 325.050 814.050 ;
        RECT 322.950 812.400 327.450 813.450 ;
        RECT 322.950 811.950 325.050 812.400 ;
        RECT 326.400 811.050 327.450 812.400 ;
        RECT 322.950 809.850 325.050 810.750 ;
        RECT 325.950 808.950 328.050 811.050 ;
        RECT 313.950 805.650 316.050 807.750 ;
        RECT 310.950 802.050 313.050 804.150 ;
        RECT 314.250 801.900 315.450 805.650 ;
        RECT 314.100 799.800 316.200 801.900 ;
        RECT 307.800 785.100 309.900 787.200 ;
        RECT 308.550 781.350 309.750 785.100 ;
        RECT 310.950 782.850 313.050 784.950 ;
        RECT 307.950 779.250 310.050 781.350 ;
        RECT 298.950 776.250 301.050 777.150 ;
        RECT 298.950 774.450 301.050 775.050 ;
        RECT 296.400 773.400 301.050 774.450 ;
        RECT 296.400 772.050 297.450 773.400 ;
        RECT 298.950 772.950 301.050 773.400 ;
        RECT 286.950 770.850 289.050 771.750 ;
        RECT 295.950 769.950 298.050 772.050 ;
        RECT 308.550 765.600 309.750 779.250 ;
        RECT 311.250 765.600 312.450 782.850 ;
        RECT 318.900 782.400 321.000 784.500 ;
        RECT 322.950 782.400 325.050 784.500 ;
        RECT 313.950 779.250 316.050 781.350 ;
        RECT 314.400 765.600 315.600 779.250 ;
        RECT 319.350 773.550 320.550 782.400 ;
        RECT 323.550 776.250 324.750 782.400 ;
        RECT 322.950 774.150 325.050 776.250 ;
        RECT 318.750 771.450 320.850 773.550 ;
        RECT 319.350 765.600 320.550 771.450 ;
        RECT 323.550 765.600 324.750 774.150 ;
        RECT 325.950 770.250 328.050 771.150 ;
        RECT 325.950 766.950 328.050 769.050 ;
        RECT 284.400 764.400 288.450 765.450 ;
        RECT 283.950 757.950 286.050 760.050 ;
        RECT 277.950 754.950 280.050 757.050 ;
        RECT 278.400 748.050 279.450 754.950 ;
        RECT 277.950 745.950 280.050 748.050 ;
        RECT 280.950 745.950 283.050 748.050 ;
        RECT 281.400 745.050 282.450 745.950 ;
        RECT 241.950 742.950 244.050 745.050 ;
        RECT 245.250 743.850 246.750 744.750 ;
        RECT 247.950 742.950 250.050 745.050 ;
        RECT 262.950 743.250 265.050 744.150 ;
        RECT 268.950 743.250 271.050 744.150 ;
        RECT 274.950 742.950 277.050 745.050 ;
        RECT 278.250 743.850 279.750 744.750 ;
        RECT 280.950 742.950 283.050 745.050 ;
        RECT 241.950 740.850 244.050 741.750 ;
        RECT 247.950 740.850 250.050 741.750 ;
        RECT 262.950 739.950 265.050 742.050 ;
        RECT 268.950 739.950 271.050 742.050 ;
        RECT 274.950 740.850 277.050 741.750 ;
        RECT 280.950 740.850 283.050 741.750 ;
        RECT 263.400 736.050 264.450 739.950 ;
        RECT 262.950 733.950 265.050 736.050 ;
        RECT 260.100 713.100 262.200 715.200 ;
        RECT 244.950 710.400 247.050 712.500 ;
        RECT 249.000 710.400 251.100 712.500 ;
        RECT 256.950 710.850 259.050 712.950 ;
        RECT 245.250 704.250 246.450 710.400 ;
        RECT 244.950 702.150 247.050 704.250 ;
        RECT 238.950 697.950 241.050 700.050 ;
        RECT 241.950 698.250 244.050 699.150 ;
        RECT 241.950 694.950 244.050 697.050 ;
        RECT 229.950 691.950 232.050 694.050 ;
        RECT 232.950 691.950 235.050 694.050 ;
        RECT 235.950 691.950 238.050 694.050 ;
        RECT 238.950 691.950 241.050 694.050 ;
        RECT 226.950 688.950 229.050 691.050 ;
        RECT 235.950 688.950 238.050 691.050 ;
        RECT 236.400 676.050 237.450 688.950 ;
        RECT 239.400 685.050 240.450 691.950 ;
        RECT 242.400 691.050 243.450 694.950 ;
        RECT 245.250 693.600 246.450 702.150 ;
        RECT 249.450 701.550 250.650 710.400 ;
        RECT 253.950 707.250 256.050 709.350 ;
        RECT 249.150 699.450 251.250 701.550 ;
        RECT 249.450 693.600 250.650 699.450 ;
        RECT 254.400 693.600 255.600 707.250 ;
        RECT 257.550 693.600 258.750 710.850 ;
        RECT 260.250 709.350 261.450 713.100 ;
        RECT 259.950 707.250 262.050 709.350 ;
        RECT 269.400 709.050 270.450 739.950 ;
        RECT 260.250 693.600 261.450 707.250 ;
        RECT 262.950 706.950 265.050 709.050 ;
        RECT 268.950 706.950 271.050 709.050 ;
        RECT 263.400 694.050 264.450 706.950 ;
        RECT 268.950 704.250 271.050 705.150 ;
        RECT 268.950 700.950 271.050 703.050 ;
        RECT 271.950 700.950 274.050 703.050 ;
        RECT 280.950 700.950 283.050 703.050 ;
        RECT 244.950 691.500 247.050 693.600 ;
        RECT 249.150 691.500 251.250 693.600 ;
        RECT 253.950 691.500 256.050 693.600 ;
        RECT 256.950 691.500 259.050 693.600 ;
        RECT 259.950 691.500 262.050 693.600 ;
        RECT 262.950 691.950 265.050 694.050 ;
        RECT 241.950 688.950 244.050 691.050 ;
        RECT 238.950 682.950 241.050 685.050 ;
        RECT 232.950 673.950 235.050 676.050 ;
        RECT 235.950 673.950 238.050 676.050 ;
        RECT 233.400 673.050 234.450 673.950 ;
        RECT 239.400 673.050 240.450 682.950 ;
        RECT 256.950 679.950 259.050 682.050 ;
        RECT 247.950 676.950 250.050 679.050 ;
        RECT 248.400 676.050 249.450 676.950 ;
        RECT 241.950 673.950 244.050 676.050 ;
        RECT 247.950 673.950 250.050 676.050 ;
        RECT 232.950 670.950 235.050 673.050 ;
        RECT 236.250 671.850 237.750 672.750 ;
        RECT 238.950 670.950 241.050 673.050 ;
        RECT 220.950 667.950 223.050 670.050 ;
        RECT 232.950 668.850 235.050 669.750 ;
        RECT 235.950 667.950 238.050 670.050 ;
        RECT 238.950 668.850 241.050 669.750 ;
        RECT 242.400 669.450 243.450 673.950 ;
        RECT 257.400 673.050 258.450 679.950 ;
        RECT 272.400 679.050 273.450 700.950 ;
        RECT 280.950 698.850 283.050 699.750 ;
        RECT 271.950 676.950 274.050 679.050 ;
        RECT 262.950 673.950 265.050 676.050 ;
        RECT 268.950 675.450 271.050 676.050 ;
        RECT 268.950 674.400 276.450 675.450 ;
        RECT 268.950 673.950 271.050 674.400 ;
        RECT 244.950 671.250 247.050 672.150 ;
        RECT 247.950 671.850 250.050 672.750 ;
        RECT 250.950 670.950 253.050 673.050 ;
        RECT 254.250 671.250 255.750 672.150 ;
        RECT 256.950 670.950 259.050 673.050 ;
        RECT 244.950 669.450 247.050 670.050 ;
        RECT 242.400 668.400 247.050 669.450 ;
        RECT 250.950 668.850 252.750 669.750 ;
        RECT 244.950 667.950 247.050 668.400 ;
        RECT 253.950 667.950 256.050 670.050 ;
        RECT 257.250 668.850 258.750 669.750 ;
        RECT 259.950 669.450 262.050 670.050 ;
        RECT 263.400 669.450 264.450 673.950 ;
        RECT 275.400 673.050 276.450 674.400 ;
        RECT 280.950 673.950 283.050 676.050 ;
        RECT 281.400 673.050 282.450 673.950 ;
        RECT 268.950 670.950 271.050 673.050 ;
        RECT 272.250 671.250 273.750 672.150 ;
        RECT 274.950 670.950 277.050 673.050 ;
        RECT 278.250 671.250 279.750 672.150 ;
        RECT 280.950 670.950 283.050 673.050 ;
        RECT 259.950 668.400 264.450 669.450 ;
        RECT 268.950 668.850 270.750 669.750 ;
        RECT 259.950 667.950 262.050 668.400 ;
        RECT 271.950 667.950 274.050 670.050 ;
        RECT 275.250 668.850 276.750 669.750 ;
        RECT 277.950 667.950 280.050 670.050 ;
        RECT 281.250 668.850 283.050 669.750 ;
        RECT 211.950 664.950 214.050 667.050 ;
        RECT 215.250 665.850 216.750 666.750 ;
        RECT 217.950 664.950 220.050 667.050 ;
        RECT 221.250 665.850 223.050 666.750 ;
        RECT 217.950 662.850 220.050 663.750 ;
        RECT 208.950 649.950 211.050 652.050 ;
        RECT 185.400 638.400 189.450 639.450 ;
        RECT 184.950 634.950 187.050 637.050 ;
        RECT 185.400 634.050 186.450 634.950 ;
        RECT 178.950 631.950 181.050 634.050 ;
        RECT 182.250 632.250 183.750 633.150 ;
        RECT 184.950 631.950 187.050 634.050 ;
        RECT 178.950 629.850 180.750 630.750 ;
        RECT 181.950 628.950 184.050 631.050 ;
        RECT 185.250 629.850 187.050 630.750 ;
        RECT 182.400 622.050 183.450 628.950 ;
        RECT 181.950 619.950 184.050 622.050 ;
        RECT 181.950 601.950 184.050 604.050 ;
        RECT 181.950 599.850 184.050 600.750 ;
        RECT 184.950 599.250 187.050 600.150 ;
        RECT 172.950 596.250 174.750 597.150 ;
        RECT 175.950 595.950 178.050 598.050 ;
        RECT 179.250 596.250 181.050 597.150 ;
        RECT 184.950 595.950 187.050 598.050 ;
        RECT 172.950 592.950 175.050 595.050 ;
        RECT 176.250 593.850 177.750 594.750 ;
        RECT 178.950 592.950 181.050 595.050 ;
        RECT 173.400 592.050 174.450 592.950 ;
        RECT 172.950 589.950 175.050 592.050 ;
        RECT 188.400 562.050 189.450 638.400 ;
        RECT 190.950 634.950 193.050 637.050 ;
        RECT 223.950 635.250 226.050 636.150 ;
        RECT 191.400 628.050 192.450 634.950 ;
        RECT 236.400 634.050 237.450 667.950 ;
        RECT 254.400 664.050 255.450 667.950 ;
        RECT 259.950 665.850 262.050 666.750 ;
        RECT 253.950 661.950 256.050 664.050 ;
        RECT 247.950 658.950 250.050 661.050 ;
        RECT 241.950 635.250 244.050 636.150 ;
        RECT 248.400 634.050 249.450 658.950 ;
        RECT 272.400 658.050 273.450 667.950 ;
        RECT 278.400 664.050 279.450 667.950 ;
        RECT 277.950 661.950 280.050 664.050 ;
        RECT 253.950 655.950 256.050 658.050 ;
        RECT 271.950 655.950 274.050 658.050 ;
        RECT 250.950 649.950 253.050 652.050 ;
        RECT 202.950 632.250 205.050 633.150 ;
        RECT 217.950 631.950 220.050 634.050 ;
        RECT 221.250 632.250 222.750 633.150 ;
        RECT 223.950 631.950 226.050 634.050 ;
        RECT 227.250 632.250 229.050 633.150 ;
        RECT 232.950 631.950 235.050 634.050 ;
        RECT 235.950 631.950 238.050 634.050 ;
        RECT 238.950 632.250 240.750 633.150 ;
        RECT 241.950 631.950 244.050 634.050 ;
        RECT 245.250 632.250 246.750 633.150 ;
        RECT 247.950 631.950 250.050 634.050 ;
        RECT 233.400 631.050 234.450 631.950 ;
        RECT 193.950 629.250 195.750 630.150 ;
        RECT 196.950 628.950 199.050 631.050 ;
        RECT 202.950 630.450 205.050 631.050 ;
        RECT 200.250 629.250 201.750 630.150 ;
        RECT 202.950 629.400 207.450 630.450 ;
        RECT 202.950 628.950 205.050 629.400 ;
        RECT 190.950 625.950 193.050 628.050 ;
        RECT 193.950 625.950 196.050 628.050 ;
        RECT 197.250 626.850 198.750 627.750 ;
        RECT 199.950 625.950 202.050 628.050 ;
        RECT 202.950 625.950 205.050 628.050 ;
        RECT 193.950 624.450 196.050 625.050 ;
        RECT 200.400 624.450 201.450 625.950 ;
        RECT 193.950 623.400 201.450 624.450 ;
        RECT 193.950 622.950 196.050 623.400 ;
        RECT 190.950 610.950 193.050 613.050 ;
        RECT 178.950 559.950 181.050 562.050 ;
        RECT 187.950 559.950 190.050 562.050 ;
        RECT 169.950 557.250 172.050 558.150 ;
        RECT 175.950 557.250 178.050 558.150 ;
        RECT 169.950 553.950 172.050 556.050 ;
        RECT 175.950 555.450 178.050 556.050 ;
        RECT 179.400 555.450 180.450 559.950 ;
        RECT 181.950 557.250 184.050 558.150 ;
        RECT 187.950 557.250 190.050 558.150 ;
        RECT 191.400 556.050 192.450 610.950 ;
        RECT 203.400 604.050 204.450 625.950 ;
        RECT 206.400 622.050 207.450 629.400 ;
        RECT 208.950 628.950 211.050 631.050 ;
        RECT 217.950 629.850 219.750 630.750 ;
        RECT 220.950 628.950 223.050 631.050 ;
        RECT 226.950 628.950 229.050 631.050 ;
        RECT 232.950 628.950 235.050 631.050 ;
        RECT 238.950 628.950 241.050 631.050 ;
        RECT 244.950 628.950 247.050 631.050 ;
        RECT 248.250 629.850 250.050 630.750 ;
        RECT 205.950 619.950 208.050 622.050 ;
        RECT 209.400 616.050 210.450 628.950 ;
        RECT 221.400 619.050 222.450 628.950 ;
        RECT 223.950 622.950 226.050 625.050 ;
        RECT 220.950 616.950 223.050 619.050 ;
        RECT 208.950 613.950 211.050 616.050 ;
        RECT 217.950 604.950 220.050 607.050 ;
        RECT 202.950 601.950 205.050 604.050 ;
        RECT 211.950 601.950 214.050 604.050 ;
        RECT 214.950 601.950 217.050 604.050 ;
        RECT 212.400 601.050 213.450 601.950 ;
        RECT 218.400 601.050 219.450 604.950 ;
        RECT 220.950 601.950 223.050 604.050 ;
        RECT 199.950 600.450 202.050 601.050 ;
        RECT 197.400 599.400 202.050 600.450 ;
        RECT 203.250 599.850 204.750 600.750 ;
        RECT 205.950 600.450 208.050 601.050 ;
        RECT 197.400 598.050 198.450 599.400 ;
        RECT 199.950 598.950 202.050 599.400 ;
        RECT 205.950 599.400 210.450 600.450 ;
        RECT 205.950 598.950 208.050 599.400 ;
        RECT 196.950 595.950 199.050 598.050 ;
        RECT 199.950 596.850 202.050 597.750 ;
        RECT 205.950 596.850 208.050 597.750 ;
        RECT 197.400 565.050 198.450 595.950 ;
        RECT 209.400 583.050 210.450 599.400 ;
        RECT 211.950 598.950 214.050 601.050 ;
        RECT 215.250 599.850 216.750 600.750 ;
        RECT 217.950 598.950 220.050 601.050 ;
        RECT 211.950 596.850 214.050 597.750 ;
        RECT 217.950 596.850 220.050 597.750 ;
        RECT 221.400 595.050 222.450 601.950 ;
        RECT 220.950 592.950 223.050 595.050 ;
        RECT 224.400 592.050 225.450 622.950 ;
        RECT 227.400 595.050 228.450 628.950 ;
        RECT 232.950 626.850 235.050 627.750 ;
        RECT 235.950 626.250 238.050 627.150 ;
        RECT 235.950 622.950 238.050 625.050 ;
        RECT 236.400 622.050 237.450 622.950 ;
        RECT 235.950 619.950 238.050 622.050 ;
        RECT 245.400 619.050 246.450 628.950 ;
        RECT 232.950 616.950 235.050 619.050 ;
        RECT 244.950 616.950 247.050 619.050 ;
        RECT 229.950 601.950 232.050 604.050 ;
        RECT 230.400 598.050 231.450 601.950 ;
        RECT 233.400 601.050 234.450 616.950 ;
        RECT 238.950 610.950 241.050 613.050 ;
        RECT 241.950 610.950 244.050 613.050 ;
        RECT 239.400 610.050 240.450 610.950 ;
        RECT 238.950 607.950 241.050 610.050 ;
        RECT 239.400 601.050 240.450 607.950 ;
        RECT 242.400 601.050 243.450 610.950 ;
        RECT 232.950 598.950 235.050 601.050 ;
        RECT 236.250 599.250 237.750 600.150 ;
        RECT 238.950 598.950 241.050 601.050 ;
        RECT 241.950 598.950 244.050 601.050 ;
        RECT 251.400 600.450 252.450 649.950 ;
        RECT 254.400 601.050 255.450 655.950 ;
        RECT 284.400 655.050 285.450 757.950 ;
        RECT 287.400 742.050 288.450 764.400 ;
        RECT 307.950 763.500 310.050 765.600 ;
        RECT 310.950 763.500 313.050 765.600 ;
        RECT 313.950 763.500 316.050 765.600 ;
        RECT 318.750 763.500 320.850 765.600 ;
        RECT 322.950 763.500 325.050 765.600 ;
        RECT 301.950 760.950 304.050 763.050 ;
        RECT 295.950 754.950 298.050 757.050 ;
        RECT 292.950 751.950 295.050 754.050 ;
        RECT 289.950 745.950 292.050 748.050 ;
        RECT 290.400 742.050 291.450 745.950 ;
        RECT 286.950 739.950 289.050 742.050 ;
        RECT 289.950 739.950 292.050 742.050 ;
        RECT 293.400 739.050 294.450 751.950 ;
        RECT 296.400 742.050 297.450 754.950 ;
        RECT 295.950 739.950 298.050 742.050 ;
        RECT 299.250 740.250 301.050 741.150 ;
        RECT 286.950 736.950 289.050 739.050 ;
        RECT 289.950 737.850 291.750 738.750 ;
        RECT 292.950 736.950 295.050 739.050 ;
        RECT 296.250 737.850 297.750 738.750 ;
        RECT 298.950 736.950 301.050 739.050 ;
        RECT 287.400 712.050 288.450 736.950 ;
        RECT 292.950 734.850 295.050 735.750 ;
        RECT 295.950 733.950 298.050 736.050 ;
        RECT 289.950 730.950 292.050 733.050 ;
        RECT 286.950 709.950 289.050 712.050 ;
        RECT 290.400 699.450 291.450 730.950 ;
        RECT 296.400 703.050 297.450 733.950 ;
        RECT 299.400 709.050 300.450 736.950 ;
        RECT 302.400 736.050 303.450 760.950 ;
        RECT 304.950 757.950 307.050 760.050 ;
        RECT 305.400 745.050 306.450 757.950 ;
        RECT 322.950 751.950 325.050 754.050 ;
        RECT 323.400 751.050 324.450 751.950 ;
        RECT 322.950 748.950 325.050 751.050 ;
        RECT 307.950 745.950 310.050 748.050 ;
        RECT 319.950 745.950 322.050 748.050 ;
        RECT 323.400 745.050 324.450 748.950 ;
        RECT 329.400 747.450 330.450 814.950 ;
        RECT 334.950 811.950 337.050 814.050 ;
        RECT 341.400 790.050 342.450 817.950 ;
        RECT 346.950 814.950 349.050 817.050 ;
        RECT 352.950 816.450 355.050 817.050 ;
        RECT 350.400 815.400 355.050 816.450 ;
        RECT 346.950 812.850 349.050 813.750 ;
        RECT 350.400 808.050 351.450 815.400 ;
        RECT 352.950 814.950 355.050 815.400 ;
        RECT 370.950 814.950 373.050 817.050 ;
        RECT 391.950 815.250 394.050 816.150 ;
        RECT 412.950 815.250 415.050 816.150 ;
        RECT 421.950 815.850 424.050 816.750 ;
        RECT 424.950 815.250 427.050 816.150 ;
        RECT 352.950 812.850 355.050 813.750 ;
        RECT 370.950 812.850 373.050 813.750 ;
        RECT 376.950 812.850 379.050 813.750 ;
        RECT 391.950 811.950 394.050 814.050 ;
        RECT 415.950 811.950 418.050 814.050 ;
        RECT 424.950 811.950 427.050 814.050 ;
        RECT 433.950 812.250 435.750 813.150 ;
        RECT 436.950 811.950 439.050 814.050 ;
        RECT 440.250 812.250 442.050 813.150 ;
        RECT 392.400 811.050 393.450 811.950 ;
        RECT 391.950 808.950 394.050 811.050 ;
        RECT 349.950 805.950 352.050 808.050 ;
        RECT 340.950 787.950 343.050 790.050 ;
        RECT 331.950 784.950 334.050 787.050 ;
        RECT 334.950 784.950 337.050 787.050 ;
        RECT 337.950 784.950 340.050 787.050 ;
        RECT 332.250 766.050 333.450 784.950 ;
        RECT 335.250 780.750 336.450 784.950 ;
        RECT 334.950 778.650 337.050 780.750 ;
        RECT 335.250 766.050 336.450 778.650 ;
        RECT 338.250 766.050 339.450 784.950 ;
        RECT 341.400 768.450 342.450 787.950 ;
        RECT 346.950 781.950 349.050 784.050 ;
        RECT 343.950 776.250 346.050 777.150 ;
        RECT 341.400 767.400 345.450 768.450 ;
        RECT 331.950 763.950 334.050 766.050 ;
        RECT 334.950 763.950 337.050 766.050 ;
        RECT 337.950 763.950 340.050 766.050 ;
        RECT 331.950 748.950 334.050 751.050 ;
        RECT 326.400 746.400 330.450 747.450 ;
        RECT 304.950 742.950 307.050 745.050 ;
        RECT 308.250 743.850 309.750 744.750 ;
        RECT 310.950 744.450 313.050 745.050 ;
        RECT 310.950 743.400 315.450 744.450 ;
        RECT 319.950 743.850 321.750 744.750 ;
        RECT 310.950 742.950 313.050 743.400 ;
        RECT 304.950 740.850 307.050 741.750 ;
        RECT 310.950 740.850 313.050 741.750 ;
        RECT 301.950 733.950 304.050 736.050 ;
        RECT 314.400 718.050 315.450 743.400 ;
        RECT 322.950 742.950 325.050 745.050 ;
        RECT 322.950 740.850 325.050 741.750 ;
        RECT 313.950 715.950 316.050 718.050 ;
        RECT 326.400 715.050 327.450 746.400 ;
        RECT 332.400 745.050 333.450 748.950 ;
        RECT 344.400 748.050 345.450 767.400 ;
        RECT 347.400 751.050 348.450 781.950 ;
        RECT 350.400 778.050 351.450 805.950 ;
        RECT 412.950 781.950 415.050 784.050 ;
        RECT 413.400 781.050 414.450 781.950 ;
        RECT 409.950 779.250 412.050 780.150 ;
        RECT 412.950 778.950 415.050 781.050 ;
        RECT 349.950 775.950 352.050 778.050 ;
        RECT 388.950 775.950 391.050 778.050 ;
        RECT 403.950 775.950 406.050 778.050 ;
        RECT 407.250 776.250 408.750 777.150 ;
        RECT 409.950 775.950 412.050 778.050 ;
        RECT 413.250 776.250 415.050 777.150 ;
        RECT 349.950 773.850 352.050 774.750 ;
        RECT 358.950 773.250 361.050 774.150 ;
        RECT 361.950 773.850 364.050 774.750 ;
        RECT 367.950 773.250 370.050 774.150 ;
        RECT 379.950 773.250 382.050 774.150 ;
        RECT 385.950 773.250 388.050 774.150 ;
        RECT 358.950 769.950 361.050 772.050 ;
        RECT 367.950 769.950 370.050 772.050 ;
        RECT 385.950 771.450 388.050 772.050 ;
        RECT 383.400 770.400 388.050 771.450 ;
        RECT 359.400 769.050 360.450 769.950 ;
        RECT 358.950 766.950 361.050 769.050 ;
        RECT 364.950 766.950 367.050 769.050 ;
        RECT 355.950 763.950 358.050 766.050 ;
        RECT 346.950 748.950 349.050 751.050 ;
        RECT 347.400 748.050 348.450 748.950 ;
        RECT 340.950 747.450 343.050 748.050 ;
        RECT 335.400 746.400 343.050 747.450 ;
        RECT 328.950 743.250 331.050 744.150 ;
        RECT 331.950 742.950 334.050 745.050 ;
        RECT 328.950 739.950 331.050 742.050 ;
        RECT 325.950 712.950 328.050 715.050 ;
        RECT 316.950 709.950 319.050 712.050 ;
        RECT 298.950 706.950 301.050 709.050 ;
        RECT 313.950 706.950 316.050 709.050 ;
        RECT 314.400 706.050 315.450 706.950 ;
        RECT 307.950 703.950 310.050 706.050 ;
        RECT 311.250 704.250 312.750 705.150 ;
        RECT 313.950 703.950 316.050 706.050 ;
        RECT 292.950 701.250 294.750 702.150 ;
        RECT 295.950 700.950 298.050 703.050 ;
        RECT 301.950 702.450 304.050 703.050 ;
        RECT 301.950 701.400 306.450 702.450 ;
        RECT 307.950 701.850 309.750 702.750 ;
        RECT 301.950 700.950 304.050 701.400 ;
        RECT 305.400 700.050 306.450 701.400 ;
        RECT 310.950 700.950 313.050 703.050 ;
        RECT 314.250 701.850 316.050 702.750 ;
        RECT 311.400 700.050 312.450 700.950 ;
        RECT 292.950 699.450 295.050 700.050 ;
        RECT 290.400 698.400 295.050 699.450 ;
        RECT 296.250 698.850 298.050 699.750 ;
        RECT 292.950 697.950 295.050 698.400 ;
        RECT 298.950 698.250 301.050 699.150 ;
        RECT 301.950 698.850 304.050 699.750 ;
        RECT 304.950 697.950 307.050 700.050 ;
        RECT 310.950 697.950 313.050 700.050 ;
        RECT 298.950 694.950 301.050 697.050 ;
        RECT 289.950 688.950 292.050 691.050 ;
        RECT 286.950 673.950 289.050 676.050 ;
        RECT 271.950 652.950 274.050 655.050 ;
        RECT 283.950 652.950 286.050 655.050 ;
        RECT 268.950 643.950 271.050 646.050 ;
        RECT 262.950 634.950 265.050 637.050 ;
        RECT 263.400 634.050 264.450 634.950 ;
        RECT 269.400 634.050 270.450 643.950 ;
        RECT 262.950 631.950 265.050 634.050 ;
        RECT 266.250 632.250 267.750 633.150 ;
        RECT 268.950 631.950 271.050 634.050 ;
        RECT 262.950 629.850 264.750 630.750 ;
        RECT 265.950 628.950 268.050 631.050 ;
        RECT 269.250 629.850 271.050 630.750 ;
        RECT 266.400 625.050 267.450 628.950 ;
        RECT 265.950 622.950 268.050 625.050 ;
        RECT 272.400 619.050 273.450 652.950 ;
        RECT 287.400 646.050 288.450 673.950 ;
        RECT 286.950 643.950 289.050 646.050 ;
        RECT 274.950 640.950 277.050 643.050 ;
        RECT 265.950 616.950 268.050 619.050 ;
        RECT 271.950 616.950 274.050 619.050 ;
        RECT 259.950 604.950 262.050 607.050 ;
        RECT 260.400 604.050 261.450 604.950 ;
        RECT 259.950 601.950 262.050 604.050 ;
        RECT 260.400 601.050 261.450 601.950 ;
        RECT 266.400 601.050 267.450 616.950 ;
        RECT 275.400 607.050 276.450 640.950 ;
        RECT 290.400 634.050 291.450 688.950 ;
        RECT 299.400 676.050 300.450 694.950 ;
        RECT 304.950 676.950 307.050 679.050 ;
        RECT 313.950 676.950 316.050 679.050 ;
        RECT 298.950 673.950 301.050 676.050 ;
        RECT 305.400 673.050 306.450 676.950 ;
        RECT 307.950 673.950 310.050 676.050 ;
        RECT 295.950 670.950 298.050 673.050 ;
        RECT 299.250 671.250 300.750 672.150 ;
        RECT 301.950 670.950 304.050 673.050 ;
        RECT 304.950 670.950 307.050 673.050 ;
        RECT 308.250 671.850 309.750 672.750 ;
        RECT 310.950 670.950 313.050 673.050 ;
        RECT 292.950 667.950 295.050 670.050 ;
        RECT 296.250 668.850 297.750 669.750 ;
        RECT 298.950 667.950 301.050 670.050 ;
        RECT 302.250 668.850 304.050 669.750 ;
        RECT 304.950 668.850 307.050 669.750 ;
        RECT 307.950 667.950 310.050 670.050 ;
        RECT 310.950 668.850 313.050 669.750 ;
        RECT 292.950 665.850 295.050 666.750 ;
        RECT 299.400 640.050 300.450 667.950 ;
        RECT 308.400 664.050 309.450 667.950 ;
        RECT 307.950 661.950 310.050 664.050 ;
        RECT 314.400 640.050 315.450 676.950 ;
        RECT 298.950 637.950 301.050 640.050 ;
        RECT 313.950 637.950 316.050 640.050 ;
        RECT 317.400 637.050 318.450 709.950 ;
        RECT 319.950 703.950 322.050 706.050 ;
        RECT 329.400 705.450 330.450 739.950 ;
        RECT 335.400 706.050 336.450 746.400 ;
        RECT 340.950 745.950 343.050 746.400 ;
        RECT 343.950 745.950 346.050 748.050 ;
        RECT 346.950 745.950 349.050 748.050 ;
        RECT 344.400 745.050 345.450 745.950 ;
        RECT 337.950 742.950 340.050 745.050 ;
        RECT 341.250 743.850 342.750 744.750 ;
        RECT 343.950 742.950 346.050 745.050 ;
        RECT 346.950 743.850 349.050 744.750 ;
        RECT 349.950 743.250 352.050 744.150 ;
        RECT 337.950 740.850 340.050 741.750 ;
        RECT 343.950 740.850 346.050 741.750 ;
        RECT 349.950 739.950 352.050 742.050 ;
        RECT 337.950 706.950 340.050 709.050 ;
        RECT 329.400 704.400 333.450 705.450 ;
        RECT 320.400 697.050 321.450 703.950 ;
        RECT 322.950 700.950 325.050 703.050 ;
        RECT 325.950 701.250 327.750 702.150 ;
        RECT 328.950 700.950 331.050 703.050 ;
        RECT 332.400 702.450 333.450 704.400 ;
        RECT 334.950 703.950 337.050 706.050 ;
        RECT 338.400 703.050 339.450 706.950 ;
        RECT 334.950 702.450 337.050 703.050 ;
        RECT 332.400 701.400 337.050 702.450 ;
        RECT 334.950 700.950 337.050 701.400 ;
        RECT 337.950 700.950 340.050 703.050 ;
        RECT 343.950 700.950 346.050 703.050 ;
        RECT 347.250 701.250 349.050 702.150 ;
        RECT 319.950 694.950 322.050 697.050 ;
        RECT 323.400 676.050 324.450 700.950 ;
        RECT 350.400 700.050 351.450 739.950 ;
        RECT 325.950 697.950 328.050 700.050 ;
        RECT 329.250 698.850 331.050 699.750 ;
        RECT 331.950 698.250 334.050 699.150 ;
        RECT 334.950 698.850 337.050 699.750 ;
        RECT 337.950 698.850 340.050 699.750 ;
        RECT 340.950 698.250 343.050 699.150 ;
        RECT 343.950 698.850 345.750 699.750 ;
        RECT 346.950 697.950 349.050 700.050 ;
        RECT 349.950 697.950 352.050 700.050 ;
        RECT 326.400 688.050 327.450 697.950 ;
        RECT 331.950 694.950 334.050 697.050 ;
        RECT 340.950 694.950 343.050 697.050 ;
        RECT 334.950 691.950 337.050 694.050 ;
        RECT 325.950 685.950 328.050 688.050 ;
        RECT 331.950 682.950 334.050 685.050 ;
        RECT 322.950 673.950 325.050 676.050 ;
        RECT 322.950 667.950 325.050 670.050 ;
        RECT 325.950 668.250 327.750 669.150 ;
        RECT 328.950 667.950 331.050 670.050 ;
        RECT 323.400 658.050 324.450 667.950 ;
        RECT 332.400 667.050 333.450 682.950 ;
        RECT 335.400 670.050 336.450 691.950 ;
        RECT 347.400 688.050 348.450 697.950 ;
        RECT 349.950 694.950 352.050 697.050 ;
        RECT 350.400 694.050 351.450 694.950 ;
        RECT 349.950 691.950 352.050 694.050 ;
        RECT 352.950 691.950 355.050 694.050 ;
        RECT 346.950 685.950 349.050 688.050 ;
        RECT 346.950 676.950 349.050 679.050 ;
        RECT 347.400 676.050 348.450 676.950 ;
        RECT 346.950 673.950 349.050 676.050 ;
        RECT 353.400 673.050 354.450 691.950 ;
        RECT 356.400 682.050 357.450 763.950 ;
        RECT 361.950 739.950 364.050 742.050 ;
        RECT 365.400 739.050 366.450 766.950 ;
        RECT 368.400 763.050 369.450 769.950 ;
        RECT 367.950 760.950 370.050 763.050 ;
        RECT 379.950 754.950 382.050 757.050 ;
        RECT 367.950 748.950 370.050 751.050 ;
        RECT 368.400 742.050 369.450 748.950 ;
        RECT 373.950 745.950 376.050 748.050 ;
        RECT 367.950 739.950 370.050 742.050 ;
        RECT 371.250 740.250 373.050 741.150 ;
        RECT 361.950 737.850 363.750 738.750 ;
        RECT 364.950 736.950 367.050 739.050 ;
        RECT 368.250 737.850 369.750 738.750 ;
        RECT 370.950 736.950 373.050 739.050 ;
        RECT 364.950 734.850 367.050 735.750 ;
        RECT 371.400 709.050 372.450 736.950 ;
        RECT 370.950 706.950 373.050 709.050 ;
        RECT 374.400 706.050 375.450 745.950 ;
        RECT 380.400 720.450 381.450 754.950 ;
        RECT 383.400 739.050 384.450 770.400 ;
        RECT 385.950 769.950 388.050 770.400 ;
        RECT 389.400 747.450 390.450 775.950 ;
        RECT 403.950 773.850 405.750 774.750 ;
        RECT 406.950 772.950 409.050 775.050 ;
        RECT 410.400 772.050 411.450 775.950 ;
        RECT 416.400 775.050 417.450 811.950 ;
        RECT 425.400 811.050 426.450 811.950 ;
        RECT 424.950 808.950 427.050 811.050 ;
        RECT 433.950 808.950 436.050 811.050 ;
        RECT 437.250 809.850 438.750 810.750 ;
        RECT 439.950 810.450 442.050 811.050 ;
        RECT 443.400 810.450 444.450 820.950 ;
        RECT 452.400 820.050 453.450 820.950 ;
        RECT 445.950 817.950 448.050 820.050 ;
        RECT 451.950 817.950 454.050 820.050 ;
        RECT 475.950 817.950 478.050 820.050 ;
        RECT 484.950 817.950 487.050 820.050 ;
        RECT 439.950 809.400 444.450 810.450 ;
        RECT 439.950 808.950 442.050 809.400 ;
        RECT 446.400 808.050 447.450 817.950 ;
        RECT 485.400 817.050 486.450 817.950 ;
        RECT 503.400 817.050 504.450 820.950 ;
        RECT 448.950 815.250 451.050 816.150 ;
        RECT 451.950 815.850 454.050 816.750 ;
        RECT 457.950 816.450 460.050 817.050 ;
        RECT 469.950 816.450 472.050 817.050 ;
        RECT 454.950 815.250 456.750 816.150 ;
        RECT 457.950 815.400 462.450 816.450 ;
        RECT 457.950 814.950 460.050 815.400 ;
        RECT 448.950 811.950 451.050 814.050 ;
        RECT 451.950 811.950 454.050 814.050 ;
        RECT 454.950 811.950 457.050 814.050 ;
        RECT 458.250 812.850 460.050 813.750 ;
        RECT 449.400 811.050 450.450 811.950 ;
        RECT 448.950 808.950 451.050 811.050 ;
        RECT 445.950 805.950 448.050 808.050 ;
        RECT 452.400 781.050 453.450 811.950 ;
        RECT 455.400 805.050 456.450 811.950 ;
        RECT 461.400 811.050 462.450 815.400 ;
        RECT 467.400 815.400 472.050 816.450 ;
        RECT 460.950 808.950 463.050 811.050 ;
        RECT 454.950 802.950 457.050 805.050 ;
        RECT 463.950 802.950 466.050 805.050 ;
        RECT 460.950 781.950 463.050 784.050 ;
        RECT 424.950 778.950 427.050 781.050 ;
        RECT 451.950 778.950 454.050 781.050 ;
        RECT 454.950 778.950 457.050 781.050 ;
        RECT 425.400 778.050 426.450 778.950 ;
        RECT 455.400 778.050 456.450 778.950 ;
        RECT 461.400 778.050 462.450 781.950 ;
        RECT 424.950 775.950 427.050 778.050 ;
        RECT 439.950 777.450 442.050 778.050 ;
        RECT 437.400 776.400 442.050 777.450 ;
        RECT 445.950 777.450 448.050 778.050 ;
        RECT 412.950 772.950 415.050 775.050 ;
        RECT 415.950 772.950 418.050 775.050 ;
        RECT 421.950 773.250 424.050 774.150 ;
        RECT 424.950 773.850 427.050 774.750 ;
        RECT 430.950 773.250 433.050 774.150 ;
        RECT 413.400 772.050 414.450 772.950 ;
        RECT 409.950 769.950 412.050 772.050 ;
        RECT 412.950 769.950 415.050 772.050 ;
        RECT 406.950 754.950 409.050 757.050 ;
        RECT 409.950 754.950 412.050 757.050 ;
        RECT 397.950 751.950 400.050 754.050 ;
        RECT 400.950 751.950 403.050 754.050 ;
        RECT 398.400 748.050 399.450 751.950 ;
        RECT 386.400 746.400 390.450 747.450 ;
        RECT 386.400 745.050 387.450 746.400 ;
        RECT 397.950 745.950 400.050 748.050 ;
        RECT 398.400 745.050 399.450 745.950 ;
        RECT 385.950 742.950 388.050 745.050 ;
        RECT 389.250 743.250 390.750 744.150 ;
        RECT 391.950 742.950 394.050 745.050 ;
        RECT 395.250 743.250 396.750 744.150 ;
        RECT 397.950 742.950 400.050 745.050 ;
        RECT 385.950 740.850 387.750 741.750 ;
        RECT 388.950 739.950 391.050 742.050 ;
        RECT 392.250 740.850 393.750 741.750 ;
        RECT 394.950 739.950 397.050 742.050 ;
        RECT 398.250 740.850 400.050 741.750 ;
        RECT 382.950 736.950 385.050 739.050 ;
        RECT 389.400 738.450 390.450 739.950 ;
        RECT 386.400 737.400 390.450 738.450 ;
        RECT 380.400 719.400 384.450 720.450 ;
        RECT 379.950 715.950 382.050 718.050 ;
        RECT 380.400 706.050 381.450 715.950 ;
        RECT 370.950 703.950 373.050 706.050 ;
        RECT 373.950 703.950 376.050 706.050 ;
        RECT 377.250 704.250 378.750 705.150 ;
        RECT 379.950 703.950 382.050 706.050 ;
        RECT 358.950 701.250 361.050 702.150 ;
        RECT 364.950 701.250 367.050 702.150 ;
        RECT 358.950 697.950 361.050 700.050 ;
        RECT 362.250 698.250 363.750 699.150 ;
        RECT 364.950 697.950 367.050 700.050 ;
        RECT 359.400 697.050 360.450 697.950 ;
        RECT 358.950 694.950 361.050 697.050 ;
        RECT 361.950 694.950 364.050 697.050 ;
        RECT 358.950 693.450 361.050 694.050 ;
        RECT 362.400 693.450 363.450 694.950 ;
        RECT 358.950 692.400 363.450 693.450 ;
        RECT 358.950 691.950 361.050 692.400 ;
        RECT 367.950 685.950 370.050 688.050 ;
        RECT 361.950 682.950 364.050 685.050 ;
        RECT 355.950 679.950 358.050 682.050 ;
        RECT 362.400 676.050 363.450 682.950 ;
        RECT 358.950 673.950 361.050 676.050 ;
        RECT 361.950 673.950 364.050 676.050 ;
        RECT 359.400 673.050 360.450 673.950 ;
        RECT 343.950 671.250 346.050 672.150 ;
        RECT 346.950 671.850 349.050 672.750 ;
        RECT 349.950 671.250 351.750 672.150 ;
        RECT 352.950 670.950 355.050 673.050 ;
        RECT 358.950 670.950 361.050 673.050 ;
        RECT 362.250 671.850 363.750 672.750 ;
        RECT 364.950 670.950 367.050 673.050 ;
        RECT 334.950 667.950 337.050 670.050 ;
        RECT 343.950 667.950 346.050 670.050 ;
        RECT 349.950 667.950 352.050 670.050 ;
        RECT 353.250 668.850 355.050 669.750 ;
        RECT 358.950 668.850 361.050 669.750 ;
        RECT 364.950 668.850 367.050 669.750 ;
        RECT 344.400 667.050 345.450 667.950 ;
        RECT 325.950 664.950 328.050 667.050 ;
        RECT 329.250 665.850 330.750 666.750 ;
        RECT 331.950 664.950 334.050 667.050 ;
        RECT 335.250 665.850 337.050 666.750 ;
        RECT 343.950 664.950 346.050 667.050 ;
        RECT 322.950 655.950 325.050 658.050 ;
        RECT 326.400 643.050 327.450 664.950 ;
        RECT 331.950 662.850 334.050 663.750 ;
        RECT 337.950 655.950 340.050 658.050 ;
        RECT 325.950 640.950 328.050 643.050 ;
        RECT 295.950 634.950 298.050 637.050 ;
        RECT 304.950 634.950 307.050 637.050 ;
        RECT 316.950 634.950 319.050 637.050 ;
        RECT 331.950 634.950 334.050 637.050 ;
        RECT 277.950 631.950 280.050 634.050 ;
        RECT 280.950 632.250 283.050 633.150 ;
        RECT 286.950 631.950 289.050 634.050 ;
        RECT 289.950 631.950 292.050 634.050 ;
        RECT 292.950 631.950 295.050 634.050 ;
        RECT 274.950 604.950 277.050 607.050 ;
        RECT 278.400 601.050 279.450 631.950 ;
        RECT 287.400 631.050 288.450 631.950 ;
        RECT 280.950 628.950 283.050 631.050 ;
        RECT 284.250 629.250 285.750 630.150 ;
        RECT 286.950 628.950 289.050 631.050 ;
        RECT 290.250 629.250 292.050 630.150 ;
        RECT 281.400 622.050 282.450 628.950 ;
        RECT 283.950 625.950 286.050 628.050 ;
        RECT 287.250 626.850 288.750 627.750 ;
        RECT 289.950 627.450 292.050 628.050 ;
        RECT 293.400 627.450 294.450 631.950 ;
        RECT 296.400 628.050 297.450 634.950 ;
        RECT 298.950 631.950 301.050 634.050 ;
        RECT 299.400 631.050 300.450 631.950 ;
        RECT 298.950 628.950 301.050 631.050 ;
        RECT 289.950 626.400 294.450 627.450 ;
        RECT 289.950 625.950 292.050 626.400 ;
        RECT 295.950 625.950 298.050 628.050 ;
        RECT 298.950 626.850 301.050 627.750 ;
        RECT 301.950 626.250 304.050 627.150 ;
        RECT 301.950 622.950 304.050 625.050 ;
        RECT 280.950 619.950 283.050 622.050 ;
        RECT 289.950 610.950 292.050 613.050 ;
        RECT 305.400 612.450 306.450 634.950 ;
        RECT 317.400 634.050 318.450 634.950 ;
        RECT 307.950 631.950 310.050 634.050 ;
        RECT 313.950 633.450 316.050 634.050 ;
        RECT 316.950 633.450 319.050 634.050 ;
        RECT 311.250 632.250 312.750 633.150 ;
        RECT 313.950 632.400 319.050 633.450 ;
        RECT 322.950 633.450 325.050 634.050 ;
        RECT 313.950 631.950 316.050 632.400 ;
        RECT 316.950 631.950 319.050 632.400 ;
        RECT 320.250 632.250 321.750 633.150 ;
        RECT 322.950 632.400 327.450 633.450 ;
        RECT 322.950 631.950 325.050 632.400 ;
        RECT 307.950 629.850 309.750 630.750 ;
        RECT 310.950 628.950 313.050 631.050 ;
        RECT 314.250 629.850 316.050 630.750 ;
        RECT 316.950 629.850 318.750 630.750 ;
        RECT 319.950 628.950 322.050 631.050 ;
        RECT 323.250 629.850 325.050 630.750 ;
        RECT 320.400 628.050 321.450 628.950 ;
        RECT 319.950 625.950 322.050 628.050 ;
        RECT 310.950 622.950 313.050 625.050 ;
        RECT 305.400 611.400 309.450 612.450 ;
        RECT 248.400 599.400 252.450 600.450 ;
        RECT 242.400 598.050 243.450 598.950 ;
        RECT 229.950 595.950 232.050 598.050 ;
        RECT 233.250 596.850 234.750 597.750 ;
        RECT 235.950 595.950 238.050 598.050 ;
        RECT 239.250 596.850 241.050 597.750 ;
        RECT 241.950 595.950 244.050 598.050 ;
        RECT 226.950 592.950 229.050 595.050 ;
        RECT 229.950 593.850 232.050 594.750 ;
        RECT 223.950 589.950 226.050 592.050 ;
        RECT 202.950 580.950 205.050 583.050 ;
        RECT 208.950 580.950 211.050 583.050 ;
        RECT 199.950 565.950 202.050 568.050 ;
        RECT 196.950 562.950 199.050 565.050 ;
        RECT 200.400 562.050 201.450 565.950 ;
        RECT 203.400 562.050 204.450 580.950 ;
        RECT 211.950 565.950 214.050 568.050 ;
        RECT 208.950 562.950 211.050 565.050 ;
        RECT 209.400 562.050 210.450 562.950 ;
        RECT 193.950 559.950 196.050 562.050 ;
        RECT 197.250 560.250 198.750 561.150 ;
        RECT 199.950 559.950 202.050 562.050 ;
        RECT 202.950 559.950 205.050 562.050 ;
        RECT 206.250 560.250 207.750 561.150 ;
        RECT 208.950 559.950 211.050 562.050 ;
        RECT 212.400 559.050 213.450 565.950 ;
        RECT 227.400 562.050 228.450 592.950 ;
        RECT 229.950 586.950 232.050 589.050 ;
        RECT 226.950 559.950 229.050 562.050 ;
        RECT 193.950 557.850 195.750 558.750 ;
        RECT 196.950 556.950 199.050 559.050 ;
        RECT 200.250 557.850 202.050 558.750 ;
        RECT 202.950 557.850 204.750 558.750 ;
        RECT 205.950 556.950 208.050 559.050 ;
        RECT 209.250 557.850 211.050 558.750 ;
        RECT 211.950 556.950 214.050 559.050 ;
        RECT 220.950 557.250 223.050 558.150 ;
        RECT 226.950 557.250 229.050 558.150 ;
        RECT 173.250 554.250 174.750 555.150 ;
        RECT 175.950 554.400 180.450 555.450 ;
        RECT 175.950 553.950 178.050 554.400 ;
        RECT 181.950 553.950 184.050 556.050 ;
        RECT 185.250 554.250 186.750 555.150 ;
        RECT 187.950 553.950 190.050 556.050 ;
        RECT 190.950 553.950 193.050 556.050 ;
        RECT 170.400 544.050 171.450 553.950 ;
        RECT 172.950 550.950 175.050 553.050 ;
        RECT 184.950 550.950 187.050 553.050 ;
        RECT 169.950 541.950 172.050 544.050 ;
        RECT 173.400 532.050 174.450 550.950 ;
        RECT 181.950 547.950 184.050 550.050 ;
        RECT 172.950 529.950 175.050 532.050 ;
        RECT 172.950 528.450 175.050 529.050 ;
        RECT 169.950 527.250 171.750 528.150 ;
        RECT 172.950 527.400 177.450 528.450 ;
        RECT 172.950 526.950 175.050 527.400 ;
        RECT 169.950 523.950 172.050 526.050 ;
        RECT 173.250 524.850 175.050 525.750 ;
        RECT 166.950 508.950 169.050 511.050 ;
        RECT 176.400 505.050 177.450 527.400 ;
        RECT 178.950 527.250 181.050 528.150 ;
        RECT 178.950 523.950 181.050 526.050 ;
        RECT 179.400 508.050 180.450 523.950 ;
        RECT 178.950 505.950 181.050 508.050 ;
        RECT 151.950 502.950 154.050 505.050 ;
        RECT 172.950 502.950 175.050 505.050 ;
        RECT 175.950 502.950 178.050 505.050 ;
        RECT 121.950 496.950 124.050 499.050 ;
        RECT 136.950 496.950 139.050 499.050 ;
        RECT 139.950 496.950 142.050 499.050 ;
        RECT 142.950 496.950 145.050 499.050 ;
        RECT 167.100 497.100 169.200 499.200 ;
        RECT 118.950 493.950 121.050 496.050 ;
        RECT 118.950 490.950 121.050 493.050 ;
        RECT 88.950 488.250 90.750 489.150 ;
        RECT 91.950 487.950 94.050 490.050 ;
        RECT 95.250 488.250 96.750 489.150 ;
        RECT 97.950 487.950 100.050 490.050 ;
        RECT 115.950 488.250 118.050 489.150 ;
        RECT 70.950 484.950 73.050 487.050 ;
        RECT 79.950 486.450 82.050 487.050 ;
        RECT 73.950 485.250 76.050 486.150 ;
        RECT 79.950 485.400 84.450 486.450 ;
        RECT 79.950 484.950 82.050 485.400 ;
        RECT 83.400 484.050 84.450 485.400 ;
        RECT 88.950 484.950 91.050 487.050 ;
        RECT 89.400 484.050 90.450 484.950 ;
        RECT 92.400 484.050 93.450 487.950 ;
        RECT 94.950 484.950 97.050 487.050 ;
        RECT 98.250 485.850 100.050 486.750 ;
        RECT 100.950 484.950 103.050 487.050 ;
        RECT 106.950 485.250 108.750 486.150 ;
        RECT 109.950 484.950 112.050 487.050 ;
        RECT 115.950 486.450 118.050 487.050 ;
        RECT 119.400 486.450 120.450 490.950 ;
        RECT 113.250 485.250 114.750 486.150 ;
        RECT 115.950 485.400 120.450 486.450 ;
        RECT 115.950 484.950 118.050 485.400 ;
        RECT 64.950 481.950 67.050 484.050 ;
        RECT 70.950 482.250 72.750 483.150 ;
        RECT 73.950 481.950 76.050 484.050 ;
        RECT 79.950 482.850 82.050 483.750 ;
        RECT 82.950 481.950 85.050 484.050 ;
        RECT 88.950 481.950 91.050 484.050 ;
        RECT 91.950 481.950 94.050 484.050 ;
        RECT 74.400 481.050 75.450 481.950 ;
        RECT 61.950 478.950 64.050 481.050 ;
        RECT 70.950 478.950 73.050 481.050 ;
        RECT 73.950 478.950 76.050 481.050 ;
        RECT 49.950 475.950 52.050 478.050 ;
        RECT 52.950 475.950 55.050 478.050 ;
        RECT 71.400 477.450 72.450 478.950 ;
        RECT 71.400 476.400 75.450 477.450 ;
        RECT 64.950 472.950 67.050 475.050 ;
        RECT 58.950 457.950 61.050 460.050 ;
        RECT 59.400 457.050 60.450 457.950 ;
        RECT 65.400 457.050 66.450 472.950 ;
        RECT 74.400 460.050 75.450 476.400 ;
        RECT 95.400 472.050 96.450 484.950 ;
        RECT 101.400 481.050 102.450 484.950 ;
        RECT 122.400 484.050 123.450 496.950 ;
        RECT 124.950 493.950 127.050 496.050 ;
        RECT 127.950 493.950 130.050 496.050 ;
        RECT 125.400 490.050 126.450 493.950 ;
        RECT 124.950 487.950 127.050 490.050 ;
        RECT 124.950 485.850 127.050 486.750 ;
        RECT 106.950 481.950 109.050 484.050 ;
        RECT 110.250 482.850 111.750 483.750 ;
        RECT 112.950 481.950 115.050 484.050 ;
        RECT 121.950 481.950 124.050 484.050 ;
        RECT 100.950 478.950 103.050 481.050 ;
        RECT 88.950 469.950 91.050 472.050 ;
        RECT 94.950 469.950 97.050 472.050 ;
        RECT 89.400 460.050 90.450 469.950 ;
        RECT 101.400 460.050 102.450 478.950 ;
        RECT 107.400 472.050 108.450 481.950 ;
        RECT 106.950 469.950 109.050 472.050 ;
        RECT 73.950 457.950 76.050 460.050 ;
        RECT 88.950 457.950 91.050 460.050 ;
        RECT 91.950 457.950 94.050 460.050 ;
        RECT 94.950 457.950 97.050 460.050 ;
        RECT 100.950 457.950 103.050 460.050 ;
        RECT 109.950 457.950 112.050 460.050 ;
        RECT 121.950 459.450 124.050 460.050 ;
        RECT 119.400 458.400 124.050 459.450 ;
        RECT 89.400 457.050 90.450 457.950 ;
        RECT 95.400 457.050 96.450 457.950 ;
        RECT 22.950 456.450 25.050 457.050 ;
        RECT 20.400 455.400 25.050 456.450 ;
        RECT 26.250 455.850 27.750 456.750 ;
        RECT 28.950 456.450 31.050 457.050 ;
        RECT 20.400 448.050 21.450 455.400 ;
        RECT 22.950 454.950 25.050 455.400 ;
        RECT 28.950 455.400 33.450 456.450 ;
        RECT 28.950 454.950 31.050 455.400 ;
        RECT 22.950 452.850 25.050 453.750 ;
        RECT 28.950 452.850 31.050 453.750 ;
        RECT 32.400 451.050 33.450 455.400 ;
        RECT 34.950 454.950 37.050 457.050 ;
        RECT 37.950 454.950 40.050 457.050 ;
        RECT 43.950 454.950 46.050 457.050 ;
        RECT 55.950 454.950 58.050 457.050 ;
        RECT 58.950 454.950 61.050 457.050 ;
        RECT 62.250 455.250 63.750 456.150 ;
        RECT 64.950 454.950 67.050 457.050 ;
        RECT 70.950 454.950 73.050 457.050 ;
        RECT 74.250 455.850 75.750 456.750 ;
        RECT 76.950 456.450 79.050 457.050 ;
        RECT 76.950 455.400 81.450 456.450 ;
        RECT 76.950 454.950 79.050 455.400 ;
        RECT 56.400 454.050 57.450 454.950 ;
        RECT 80.400 454.050 81.450 455.400 ;
        RECT 85.950 454.950 88.050 457.050 ;
        RECT 88.950 454.950 91.050 457.050 ;
        RECT 92.250 455.850 93.750 456.750 ;
        RECT 94.950 454.950 97.050 457.050 ;
        RECT 34.950 452.850 37.050 453.750 ;
        RECT 40.950 452.250 43.050 453.150 ;
        RECT 43.950 452.850 46.050 453.750 ;
        RECT 55.950 451.950 58.050 454.050 ;
        RECT 59.250 452.850 60.750 453.750 ;
        RECT 61.950 451.950 64.050 454.050 ;
        RECT 65.250 452.850 67.050 453.750 ;
        RECT 70.950 452.850 73.050 453.750 ;
        RECT 76.950 452.850 79.050 453.750 ;
        RECT 79.950 451.950 82.050 454.050 ;
        RECT 31.950 448.950 34.050 451.050 ;
        RECT 40.950 448.950 43.050 451.050 ;
        RECT 49.950 448.950 52.050 451.050 ;
        RECT 55.950 449.850 58.050 450.750 ;
        RECT 19.950 445.950 22.050 448.050 ;
        RECT 22.950 445.950 25.050 448.050 ;
        RECT 16.950 439.950 19.050 442.050 ;
        RECT 23.400 415.050 24.450 445.950 ;
        RECT 31.950 424.950 34.050 427.050 ;
        RECT 28.950 416.250 31.050 417.150 ;
        RECT 19.950 413.250 21.750 414.150 ;
        RECT 22.950 412.950 25.050 415.050 ;
        RECT 28.950 414.450 31.050 415.050 ;
        RECT 32.400 414.450 33.450 424.950 ;
        RECT 50.400 424.050 51.450 448.950 ;
        RECT 49.950 421.950 52.050 424.050 ;
        RECT 40.950 417.450 43.050 418.050 ;
        RECT 38.400 416.400 43.050 417.450 ;
        RECT 26.250 413.250 27.750 414.150 ;
        RECT 28.950 413.400 33.450 414.450 ;
        RECT 28.950 412.950 31.050 413.400 ;
        RECT 34.950 412.950 37.050 415.050 ;
        RECT 7.950 410.850 10.050 411.750 ;
        RECT 10.950 410.250 13.050 411.150 ;
        RECT 13.950 409.950 16.050 412.050 ;
        RECT 19.950 409.950 22.050 412.050 ;
        RECT 23.250 410.850 24.750 411.750 ;
        RECT 25.950 409.950 28.050 412.050 ;
        RECT 10.950 406.950 13.050 409.050 ;
        RECT 11.400 394.050 12.450 406.950 ;
        RECT 10.950 391.950 13.050 394.050 ;
        RECT 20.400 391.050 21.450 409.950 ;
        RECT 25.950 406.950 28.050 409.050 ;
        RECT 16.950 388.950 19.050 391.050 ;
        RECT 19.950 388.950 22.050 391.050 ;
        RECT 10.950 385.950 13.050 388.050 ;
        RECT 11.400 382.050 12.450 385.950 ;
        RECT 7.950 380.250 9.750 381.150 ;
        RECT 10.950 379.950 13.050 382.050 ;
        RECT 14.250 380.250 16.050 381.150 ;
        RECT 7.950 376.950 10.050 379.050 ;
        RECT 11.250 377.850 12.750 378.750 ;
        RECT 13.950 376.950 16.050 379.050 ;
        RECT 8.400 375.450 9.450 376.950 ;
        RECT 14.400 376.050 15.450 376.950 ;
        RECT 8.400 374.400 12.450 375.450 ;
        RECT 1.950 355.950 4.050 358.050 ;
        RECT 2.400 307.050 3.450 355.950 ;
        RECT 7.950 342.450 10.050 343.050 ;
        RECT 5.400 341.400 10.050 342.450 ;
        RECT 5.400 312.450 6.450 341.400 ;
        RECT 7.950 340.950 10.050 341.400 ;
        RECT 7.950 338.850 10.050 339.750 ;
        RECT 11.400 331.050 12.450 374.400 ;
        RECT 13.950 373.950 16.050 376.050 ;
        RECT 17.400 342.450 18.450 388.950 ;
        RECT 19.950 385.950 22.050 388.050 ;
        RECT 19.950 383.850 22.050 384.750 ;
        RECT 22.950 383.250 25.050 384.150 ;
        RECT 22.950 379.950 25.050 382.050 ;
        RECT 23.400 343.050 24.450 379.950 ;
        RECT 26.400 346.050 27.450 406.950 ;
        RECT 35.400 406.050 36.450 412.950 ;
        RECT 38.400 409.050 39.450 416.400 ;
        RECT 40.950 415.950 43.050 416.400 ;
        RECT 44.250 416.250 45.750 417.150 ;
        RECT 46.950 415.950 49.050 418.050 ;
        RECT 50.400 415.050 51.450 421.950 ;
        RECT 62.400 421.050 63.450 451.950 ;
        RECT 64.950 436.950 67.050 439.050 ;
        RECT 61.950 418.950 64.050 421.050 ;
        RECT 52.950 416.250 55.050 417.150 ;
        RECT 58.950 415.950 61.050 418.050 ;
        RECT 59.400 415.050 60.450 415.950 ;
        RECT 40.950 413.850 42.750 414.750 ;
        RECT 43.950 412.950 46.050 415.050 ;
        RECT 47.250 413.850 49.050 414.750 ;
        RECT 49.950 412.950 52.050 415.050 ;
        RECT 52.950 412.950 55.050 415.050 ;
        RECT 56.250 413.250 57.750 414.150 ;
        RECT 58.950 412.950 61.050 415.050 ;
        RECT 62.250 413.250 64.050 414.150 ;
        RECT 53.400 412.050 54.450 412.950 ;
        RECT 52.950 409.950 55.050 412.050 ;
        RECT 55.950 409.950 58.050 412.050 ;
        RECT 59.250 410.850 60.750 411.750 ;
        RECT 61.950 409.950 64.050 412.050 ;
        RECT 62.400 409.050 63.450 409.950 ;
        RECT 37.950 406.950 40.050 409.050 ;
        RECT 61.950 406.950 64.050 409.050 ;
        RECT 34.950 403.950 37.050 406.050 ;
        RECT 62.400 403.050 63.450 406.950 ;
        RECT 61.950 400.950 64.050 403.050 ;
        RECT 37.950 391.950 40.050 394.050 ;
        RECT 38.400 382.050 39.450 391.950 ;
        RECT 65.400 385.050 66.450 436.950 ;
        RECT 67.950 418.950 70.050 421.050 ;
        RECT 68.400 408.450 69.450 418.950 ;
        RECT 73.950 415.950 76.050 418.050 ;
        RECT 79.950 416.250 82.050 417.150 ;
        RECT 82.950 415.950 85.050 418.050 ;
        RECT 74.400 415.050 75.450 415.950 ;
        RECT 70.950 413.250 72.750 414.150 ;
        RECT 73.950 412.950 76.050 415.050 ;
        RECT 77.250 413.250 78.750 414.150 ;
        RECT 79.950 412.950 82.050 415.050 ;
        RECT 70.950 409.950 73.050 412.050 ;
        RECT 74.250 410.850 75.750 411.750 ;
        RECT 76.950 409.950 79.050 412.050 ;
        RECT 68.400 407.400 72.450 408.450 ;
        RECT 43.950 382.950 46.050 385.050 ;
        RECT 52.950 382.950 55.050 385.050 ;
        RECT 58.950 382.950 61.050 385.050 ;
        RECT 64.950 382.950 67.050 385.050 ;
        RECT 34.950 380.250 36.750 381.150 ;
        RECT 37.950 379.950 40.050 382.050 ;
        RECT 41.250 380.250 43.050 381.150 ;
        RECT 34.950 376.950 37.050 379.050 ;
        RECT 38.250 377.850 39.750 378.750 ;
        RECT 40.950 378.450 43.050 379.050 ;
        RECT 44.400 378.450 45.450 382.950 ;
        RECT 53.400 382.050 54.450 382.950 ;
        RECT 49.950 380.250 51.750 381.150 ;
        RECT 52.950 379.950 55.050 382.050 ;
        RECT 56.250 380.250 58.050 381.150 ;
        RECT 40.950 377.400 45.450 378.450 ;
        RECT 40.950 376.950 43.050 377.400 ;
        RECT 49.950 376.950 52.050 379.050 ;
        RECT 53.250 377.850 54.750 378.750 ;
        RECT 55.950 378.450 58.050 379.050 ;
        RECT 59.400 378.450 60.450 382.950 ;
        RECT 61.950 380.250 63.750 381.150 ;
        RECT 64.950 379.950 67.050 382.050 ;
        RECT 68.250 380.250 70.050 381.150 ;
        RECT 71.400 379.050 72.450 407.400 ;
        RECT 77.400 397.050 78.450 409.950 ;
        RECT 76.950 394.950 79.050 397.050 ;
        RECT 80.400 388.050 81.450 412.950 ;
        RECT 83.400 412.050 84.450 415.950 ;
        RECT 82.950 409.950 85.050 412.050 ;
        RECT 79.950 385.950 82.050 388.050 ;
        RECT 82.950 385.950 85.050 388.050 ;
        RECT 83.400 385.050 84.450 385.950 ;
        RECT 76.950 382.950 79.050 385.050 ;
        RECT 80.250 383.850 81.750 384.750 ;
        RECT 82.950 382.950 85.050 385.050 ;
        RECT 76.950 380.850 79.050 381.750 ;
        RECT 82.950 380.850 85.050 381.750 ;
        RECT 55.950 377.400 60.450 378.450 ;
        RECT 55.950 376.950 58.050 377.400 ;
        RECT 61.950 376.950 64.050 379.050 ;
        RECT 65.250 377.850 66.750 378.750 ;
        RECT 67.950 376.950 70.050 379.050 ;
        RECT 70.950 376.950 73.050 379.050 ;
        RECT 50.400 355.050 51.450 376.950 ;
        RECT 62.400 370.050 63.450 376.950 ;
        RECT 64.950 373.950 67.050 376.050 ;
        RECT 61.950 367.950 64.050 370.050 ;
        RECT 49.950 352.950 52.050 355.050 ;
        RECT 31.950 346.950 34.050 349.050 ;
        RECT 37.950 346.950 40.050 349.050 ;
        RECT 32.400 346.050 33.450 346.950 ;
        RECT 25.950 343.950 28.050 346.050 ;
        RECT 29.250 344.250 30.750 345.150 ;
        RECT 31.950 343.950 34.050 346.050 ;
        RECT 34.950 343.950 37.050 346.050 ;
        RECT 13.950 341.250 16.050 342.150 ;
        RECT 17.400 341.400 21.450 342.450 ;
        RECT 13.950 337.950 16.050 340.050 ;
        RECT 17.250 338.250 19.050 339.150 ;
        RECT 16.950 334.950 19.050 337.050 ;
        RECT 10.950 328.950 13.050 331.050 ;
        RECT 13.950 316.950 16.050 319.050 ;
        RECT 14.400 313.050 15.450 316.950 ;
        RECT 20.400 313.050 21.450 341.400 ;
        RECT 22.950 340.950 25.050 343.050 ;
        RECT 25.950 341.850 27.750 342.750 ;
        RECT 28.950 340.950 31.050 343.050 ;
        RECT 32.250 341.850 34.050 342.750 ;
        RECT 23.400 337.050 24.450 340.950 ;
        RECT 29.400 340.050 30.450 340.950 ;
        RECT 35.400 340.050 36.450 343.950 ;
        RECT 28.950 337.950 31.050 340.050 ;
        RECT 34.950 337.950 37.050 340.050 ;
        RECT 22.950 334.950 25.050 337.050 ;
        RECT 29.400 334.050 30.450 337.950 ;
        RECT 38.400 337.050 39.450 346.950 ;
        RECT 40.950 341.250 43.050 342.150 ;
        RECT 46.950 341.250 49.050 342.150 ;
        RECT 40.950 337.950 43.050 340.050 ;
        RECT 44.250 338.250 45.750 339.150 ;
        RECT 46.950 337.950 49.050 340.050 ;
        RECT 34.950 334.950 37.050 337.050 ;
        RECT 37.950 334.950 40.050 337.050 ;
        RECT 28.950 331.950 31.050 334.050 ;
        RECT 28.950 313.950 31.050 316.050 ;
        RECT 31.950 313.950 34.050 316.050 ;
        RECT 29.400 313.050 30.450 313.950 ;
        RECT 7.950 312.450 10.050 313.050 ;
        RECT 5.400 311.400 10.050 312.450 ;
        RECT 7.950 310.950 10.050 311.400 ;
        RECT 11.250 311.250 12.750 312.150 ;
        RECT 13.950 310.950 16.050 313.050 ;
        RECT 19.950 312.450 22.050 313.050 ;
        RECT 17.250 311.250 18.750 312.150 ;
        RECT 19.950 311.400 24.450 312.450 ;
        RECT 19.950 310.950 22.050 311.400 ;
        RECT 7.950 308.850 9.750 309.750 ;
        RECT 10.950 307.950 13.050 310.050 ;
        RECT 14.250 308.850 15.750 309.750 ;
        RECT 16.950 307.950 19.050 310.050 ;
        RECT 20.250 308.850 22.050 309.750 ;
        RECT 23.400 309.450 24.450 311.400 ;
        RECT 25.950 311.250 27.750 312.150 ;
        RECT 28.950 310.950 31.050 313.050 ;
        RECT 25.950 309.450 28.050 310.050 ;
        RECT 23.400 308.400 28.050 309.450 ;
        RECT 29.250 308.850 31.050 309.750 ;
        RECT 25.950 307.950 28.050 308.400 ;
        RECT 1.950 304.950 4.050 307.050 ;
        RECT 7.950 304.950 10.050 307.050 ;
        RECT 1.950 286.950 4.050 289.050 ;
        RECT 2.400 223.050 3.450 286.950 ;
        RECT 4.950 283.950 7.050 286.050 ;
        RECT 5.400 274.050 6.450 283.950 ;
        RECT 4.950 271.950 7.050 274.050 ;
        RECT 4.950 269.850 7.050 270.750 ;
        RECT 8.400 265.050 9.450 304.950 ;
        RECT 11.400 292.050 12.450 307.950 ;
        RECT 10.950 289.950 13.050 292.050 ;
        RECT 13.950 283.950 16.050 286.050 ;
        RECT 10.950 272.250 13.050 273.150 ;
        RECT 7.950 262.950 10.050 265.050 ;
        RECT 8.400 241.050 9.450 262.950 ;
        RECT 14.400 247.050 15.450 283.950 ;
        RECT 16.950 280.950 19.050 283.050 ;
        RECT 19.950 280.950 22.050 283.050 ;
        RECT 22.950 280.950 25.050 283.050 ;
        RECT 17.550 262.050 18.750 280.950 ;
        RECT 20.550 276.750 21.750 280.950 ;
        RECT 19.950 274.650 22.050 276.750 ;
        RECT 20.550 262.050 21.750 274.650 ;
        RECT 23.550 262.050 24.750 280.950 ;
        RECT 26.400 271.050 27.450 307.950 ;
        RECT 32.400 307.050 33.450 313.950 ;
        RECT 31.950 304.950 34.050 307.050 ;
        RECT 35.400 295.050 36.450 334.950 ;
        RECT 37.950 328.950 40.050 331.050 ;
        RECT 38.400 301.050 39.450 328.950 ;
        RECT 41.400 316.050 42.450 337.950 ;
        RECT 47.400 337.050 48.450 337.950 ;
        RECT 43.950 334.950 46.050 337.050 ;
        RECT 46.950 334.950 49.050 337.050 ;
        RECT 44.400 328.050 45.450 334.950 ;
        RECT 43.950 325.950 46.050 328.050 ;
        RECT 43.950 319.950 46.050 322.050 ;
        RECT 40.950 313.950 43.050 316.050 ;
        RECT 44.400 313.050 45.450 319.950 ;
        RECT 43.950 310.950 46.050 313.050 ;
        RECT 40.950 308.250 42.750 309.150 ;
        RECT 43.950 307.950 46.050 310.050 ;
        RECT 47.250 308.250 49.050 309.150 ;
        RECT 40.950 304.950 43.050 307.050 ;
        RECT 44.250 305.850 45.750 306.750 ;
        RECT 46.950 304.950 49.050 307.050 ;
        RECT 37.950 298.950 40.050 301.050 ;
        RECT 47.400 298.050 48.450 304.950 ;
        RECT 46.950 295.950 49.050 298.050 ;
        RECT 34.950 292.950 37.050 295.050 ;
        RECT 50.400 289.050 51.450 352.950 ;
        RECT 58.950 343.950 61.050 346.050 ;
        RECT 59.400 343.050 60.450 343.950 ;
        RECT 52.950 340.950 55.050 343.050 ;
        RECT 58.950 340.950 61.050 343.050 ;
        RECT 62.250 341.250 64.050 342.150 ;
        RECT 65.400 340.050 66.450 373.950 ;
        RECT 68.400 373.050 69.450 376.950 ;
        RECT 67.950 370.950 70.050 373.050 ;
        RECT 67.950 343.950 70.050 346.050 ;
        RECT 52.950 338.850 55.050 339.750 ;
        RECT 55.950 338.250 58.050 339.150 ;
        RECT 58.950 338.850 60.750 339.750 ;
        RECT 61.950 337.950 64.050 340.050 ;
        RECT 64.950 337.950 67.050 340.050 ;
        RECT 55.950 334.950 58.050 337.050 ;
        RECT 56.400 334.050 57.450 334.950 ;
        RECT 55.950 331.950 58.050 334.050 ;
        RECT 62.400 325.050 63.450 337.950 ;
        RECT 61.950 322.950 64.050 325.050 ;
        RECT 65.400 322.050 66.450 337.950 ;
        RECT 68.400 328.050 69.450 343.950 ;
        RECT 67.950 325.950 70.050 328.050 ;
        RECT 64.950 319.950 67.050 322.050 ;
        RECT 71.400 319.050 72.450 376.950 ;
        RECT 86.400 376.050 87.450 454.950 ;
        RECT 88.950 452.850 91.050 453.750 ;
        RECT 94.950 452.850 97.050 453.750 ;
        RECT 97.950 451.950 100.050 454.050 ;
        RECT 94.950 448.950 97.050 451.050 ;
        RECT 88.950 439.950 91.050 442.050 ;
        RECT 89.400 418.050 90.450 439.950 ;
        RECT 95.400 421.050 96.450 448.950 ;
        RECT 98.400 442.050 99.450 451.950 ;
        RECT 97.950 439.950 100.050 442.050 ;
        RECT 101.400 427.050 102.450 457.950 ;
        RECT 110.400 454.050 111.450 457.950 ;
        RECT 103.950 451.950 106.050 454.050 ;
        RECT 109.950 451.950 112.050 454.050 ;
        RECT 113.250 452.250 115.050 453.150 ;
        RECT 103.950 449.850 105.750 450.750 ;
        RECT 106.950 448.950 109.050 451.050 ;
        RECT 110.250 449.850 111.750 450.750 ;
        RECT 112.950 448.950 115.050 451.050 ;
        RECT 106.950 446.850 109.050 447.750 ;
        RECT 100.950 424.950 103.050 427.050 ;
        RECT 97.950 421.950 100.050 424.050 ;
        RECT 94.950 418.950 97.050 421.050 ;
        RECT 95.400 418.050 96.450 418.950 ;
        RECT 88.950 415.950 91.050 418.050 ;
        RECT 92.250 416.250 93.750 417.150 ;
        RECT 94.950 415.950 97.050 418.050 ;
        RECT 88.950 413.850 90.750 414.750 ;
        RECT 91.950 412.950 94.050 415.050 ;
        RECT 95.250 413.850 97.050 414.750 ;
        RECT 92.400 412.050 93.450 412.950 ;
        RECT 91.950 409.950 94.050 412.050 ;
        RECT 98.400 411.450 99.450 421.950 ;
        RECT 101.400 421.050 102.450 424.950 ;
        RECT 100.950 418.950 103.050 421.050 ;
        RECT 103.950 418.950 106.050 421.050 ;
        RECT 104.400 415.050 105.450 418.950 ;
        RECT 109.950 416.250 112.050 417.150 ;
        RECT 100.950 413.250 102.750 414.150 ;
        RECT 103.950 412.950 106.050 415.050 ;
        RECT 107.250 413.250 108.750 414.150 ;
        RECT 109.950 412.950 112.050 415.050 ;
        RECT 100.950 411.450 103.050 412.050 ;
        RECT 98.400 410.400 103.050 411.450 ;
        RECT 104.250 410.850 105.750 411.750 ;
        RECT 100.950 409.950 103.050 410.400 ;
        RECT 106.950 409.950 109.050 412.050 ;
        RECT 97.950 406.950 100.050 409.050 ;
        RECT 98.400 394.050 99.450 406.950 ;
        RECT 110.400 400.050 111.450 412.950 ;
        RECT 109.950 397.950 112.050 400.050 ;
        RECT 113.400 397.050 114.450 448.950 ;
        RECT 119.400 439.050 120.450 458.400 ;
        RECT 121.950 457.950 124.050 458.400 ;
        RECT 121.950 455.850 124.050 456.750 ;
        RECT 124.950 455.250 127.050 456.150 ;
        RECT 124.950 451.950 127.050 454.050 ;
        RECT 118.950 436.950 121.050 439.050 ;
        RECT 125.400 418.050 126.450 451.950 ;
        RECT 128.400 451.050 129.450 493.950 ;
        RECT 130.950 488.250 133.050 489.150 ;
        RECT 133.950 487.950 136.050 490.050 ;
        RECT 134.400 477.450 135.450 487.950 ;
        RECT 137.550 478.050 138.750 496.950 ;
        RECT 140.550 492.750 141.750 496.950 ;
        RECT 139.950 490.650 142.050 492.750 ;
        RECT 140.550 478.050 141.750 490.650 ;
        RECT 143.550 478.050 144.750 496.950 ;
        RECT 151.950 494.400 154.050 496.500 ;
        RECT 156.000 494.400 158.100 496.500 ;
        RECT 163.950 494.850 166.050 496.950 ;
        RECT 152.250 488.250 153.450 494.400 ;
        RECT 151.950 486.150 154.050 488.250 ;
        RECT 148.950 482.250 151.050 483.150 ;
        RECT 148.950 478.950 151.050 481.050 ;
        RECT 149.400 478.050 150.450 478.950 ;
        RECT 131.400 476.400 135.450 477.450 ;
        RECT 127.950 448.950 130.050 451.050 ;
        RECT 127.950 421.950 130.050 424.050 ;
        RECT 118.950 415.950 121.050 418.050 ;
        RECT 121.950 416.250 124.050 417.150 ;
        RECT 124.950 415.950 127.050 418.050 ;
        RECT 103.950 394.950 106.050 397.050 ;
        RECT 112.950 394.950 115.050 397.050 ;
        RECT 97.950 391.950 100.050 394.050 ;
        RECT 94.950 387.450 97.050 388.050 ;
        RECT 89.400 386.400 97.050 387.450 ;
        RECT 89.400 385.050 90.450 386.400 ;
        RECT 94.950 385.950 97.050 386.400 ;
        RECT 97.950 385.950 100.050 388.050 ;
        RECT 98.400 385.050 99.450 385.950 ;
        RECT 88.950 382.950 91.050 385.050 ;
        RECT 91.950 382.950 94.050 385.050 ;
        RECT 95.250 383.850 96.750 384.750 ;
        RECT 97.950 382.950 100.050 385.050 ;
        RECT 91.950 380.850 94.050 381.750 ;
        RECT 97.950 380.850 100.050 381.750 ;
        RECT 85.950 373.950 88.050 376.050 ;
        RECT 94.950 373.950 97.050 376.050 ;
        RECT 73.950 340.950 76.050 343.050 ;
        RECT 76.950 341.250 79.050 342.150 ;
        RECT 82.950 341.250 85.050 342.150 ;
        RECT 85.950 341.250 88.050 342.150 ;
        RECT 91.950 341.250 94.050 342.150 ;
        RECT 74.400 339.450 75.450 340.950 ;
        RECT 76.950 339.450 79.050 340.050 ;
        RECT 74.400 338.400 79.050 339.450 ;
        RECT 76.950 337.950 79.050 338.400 ;
        RECT 80.250 338.250 81.750 339.150 ;
        RECT 82.950 337.950 85.050 340.050 ;
        RECT 85.950 337.950 88.050 340.050 ;
        RECT 89.250 338.250 90.750 339.150 ;
        RECT 91.950 337.950 94.050 340.050 ;
        RECT 76.950 334.950 79.050 337.050 ;
        RECT 79.950 334.950 82.050 337.050 ;
        RECT 83.400 336.450 84.450 337.950 ;
        RECT 88.950 336.450 91.050 337.050 ;
        RECT 83.400 335.400 91.050 336.450 ;
        RECT 88.950 334.950 91.050 335.400 ;
        RECT 67.950 316.950 70.050 319.050 ;
        RECT 70.950 316.950 73.050 319.050 ;
        RECT 55.950 313.950 58.050 316.050 ;
        RECT 68.400 313.050 69.450 316.950 ;
        RECT 73.950 313.950 76.050 316.050 ;
        RECT 74.400 313.050 75.450 313.950 ;
        RECT 77.400 313.050 78.450 334.950 ;
        RECT 88.950 331.950 91.050 334.050 ;
        RECT 89.400 321.450 90.450 331.950 ;
        RECT 92.400 331.050 93.450 337.950 ;
        RECT 91.950 328.950 94.050 331.050 ;
        RECT 89.400 320.400 93.450 321.450 ;
        RECT 79.950 316.950 82.050 319.050 ;
        RECT 88.950 316.950 91.050 319.050 ;
        RECT 52.950 311.250 55.050 312.150 ;
        RECT 55.950 311.850 58.050 312.750 ;
        RECT 61.950 312.450 64.050 313.050 ;
        RECT 58.950 311.250 60.750 312.150 ;
        RECT 61.950 311.400 66.450 312.450 ;
        RECT 61.950 310.950 64.050 311.400 ;
        RECT 52.950 307.950 55.050 310.050 ;
        RECT 58.950 307.950 61.050 310.050 ;
        RECT 62.250 308.850 64.050 309.750 ;
        RECT 58.950 304.950 61.050 307.050 ;
        RECT 49.950 286.950 52.050 289.050 ;
        RECT 47.100 281.100 49.200 283.200 ;
        RECT 31.950 278.400 34.050 280.500 ;
        RECT 36.000 278.400 38.100 280.500 ;
        RECT 43.950 278.850 46.050 280.950 ;
        RECT 32.250 272.250 33.450 278.400 ;
        RECT 25.950 268.950 28.050 271.050 ;
        RECT 31.950 270.150 34.050 272.250 ;
        RECT 25.950 265.950 28.050 268.050 ;
        RECT 28.950 266.250 31.050 267.150 ;
        RECT 16.950 259.950 19.050 262.050 ;
        RECT 19.950 259.950 22.050 262.050 ;
        RECT 22.950 259.950 25.050 262.050 ;
        RECT 26.400 256.050 27.450 265.950 ;
        RECT 28.950 262.950 31.050 265.050 ;
        RECT 25.950 253.950 28.050 256.050 ;
        RECT 25.950 250.950 28.050 253.050 ;
        RECT 16.950 247.950 19.050 250.050 ;
        RECT 13.950 244.950 16.050 247.050 ;
        RECT 7.950 240.450 10.050 241.050 ;
        RECT 5.400 239.400 10.050 240.450 ;
        RECT 1.950 220.950 4.050 223.050 ;
        RECT 1.950 199.950 4.050 202.050 ;
        RECT 2.400 129.450 3.450 199.950 ;
        RECT 5.400 162.450 6.450 239.400 ;
        RECT 7.950 238.950 10.050 239.400 ;
        RECT 11.250 239.250 13.050 240.150 ;
        RECT 7.950 236.850 9.750 237.750 ;
        RECT 10.950 235.950 13.050 238.050 ;
        RECT 7.950 232.950 10.050 235.050 ;
        RECT 17.400 234.450 18.450 247.950 ;
        RECT 26.400 241.050 27.450 250.950 ;
        RECT 29.400 250.050 30.450 262.950 ;
        RECT 32.250 261.600 33.450 270.150 ;
        RECT 36.450 269.550 37.650 278.400 ;
        RECT 40.950 275.250 43.050 277.350 ;
        RECT 36.150 267.450 38.250 269.550 ;
        RECT 36.450 261.600 37.650 267.450 ;
        RECT 41.400 261.600 42.600 275.250 ;
        RECT 44.550 261.600 45.750 278.850 ;
        RECT 47.250 277.350 48.450 281.100 ;
        RECT 46.950 275.250 49.050 277.350 ;
        RECT 47.250 261.600 48.450 275.250 ;
        RECT 55.950 272.250 58.050 273.150 ;
        RECT 52.950 268.950 55.050 271.050 ;
        RECT 55.950 268.950 58.050 271.050 ;
        RECT 31.950 259.500 34.050 261.600 ;
        RECT 36.150 259.500 38.250 261.600 ;
        RECT 40.950 259.500 43.050 261.600 ;
        RECT 43.950 259.500 46.050 261.600 ;
        RECT 46.950 259.500 49.050 261.600 ;
        RECT 49.950 256.950 52.050 259.050 ;
        RECT 34.950 253.950 37.050 256.050 ;
        RECT 28.950 247.950 31.050 250.050 ;
        RECT 31.950 247.950 34.050 250.050 ;
        RECT 28.950 244.950 31.050 247.050 ;
        RECT 19.950 238.950 22.050 241.050 ;
        RECT 23.250 239.250 24.750 240.150 ;
        RECT 25.950 238.950 28.050 241.050 ;
        RECT 29.400 238.050 30.450 244.950 ;
        RECT 19.950 236.850 21.750 237.750 ;
        RECT 22.950 235.950 25.050 238.050 ;
        RECT 26.250 236.850 27.750 237.750 ;
        RECT 28.950 235.950 31.050 238.050 ;
        RECT 17.400 233.400 21.450 234.450 ;
        RECT 8.400 202.050 9.450 232.950 ;
        RECT 16.950 229.950 19.050 232.050 ;
        RECT 7.950 199.950 10.050 202.050 ;
        RECT 10.950 199.950 13.050 202.050 ;
        RECT 11.400 199.050 12.450 199.950 ;
        RECT 7.950 197.250 9.750 198.150 ;
        RECT 10.950 196.950 13.050 199.050 ;
        RECT 7.950 193.950 10.050 196.050 ;
        RECT 11.250 194.850 13.050 195.750 ;
        RECT 8.400 169.050 9.450 193.950 ;
        RECT 17.400 169.050 18.450 229.950 ;
        RECT 7.950 166.950 10.050 169.050 ;
        RECT 16.950 166.950 19.050 169.050 ;
        RECT 7.950 164.250 9.750 165.150 ;
        RECT 10.950 163.950 13.050 166.050 ;
        RECT 14.250 164.250 16.050 165.150 ;
        RECT 7.950 162.450 10.050 163.050 ;
        RECT 5.400 161.400 10.050 162.450 ;
        RECT 11.250 161.850 12.750 162.750 ;
        RECT 13.950 162.450 16.050 163.050 ;
        RECT 17.400 162.450 18.450 166.950 ;
        RECT 7.950 160.950 10.050 161.400 ;
        RECT 13.950 161.400 18.450 162.450 ;
        RECT 13.950 160.950 16.050 161.400 ;
        RECT 4.950 129.450 7.050 130.050 ;
        RECT 2.400 128.400 7.050 129.450 ;
        RECT 2.400 57.450 3.450 128.400 ;
        RECT 4.950 127.950 7.050 128.400 ;
        RECT 4.950 125.850 7.050 126.750 ;
        RECT 8.400 100.050 9.450 160.950 ;
        RECT 10.950 128.250 13.050 129.150 ;
        RECT 7.950 97.950 10.050 100.050 ;
        RECT 14.400 97.050 15.450 160.950 ;
        RECT 20.400 160.050 21.450 233.400 ;
        RECT 23.400 208.050 24.450 235.950 ;
        RECT 28.950 233.850 31.050 234.750 ;
        RECT 32.400 211.050 33.450 247.950 ;
        RECT 31.950 208.950 34.050 211.050 ;
        RECT 35.400 208.050 36.450 253.950 ;
        RECT 43.950 247.950 46.050 250.050 ;
        RECT 50.400 249.450 51.450 256.950 ;
        RECT 47.400 248.400 51.450 249.450 ;
        RECT 37.950 241.950 40.050 244.050 ;
        RECT 38.400 241.050 39.450 241.950 ;
        RECT 44.400 241.050 45.450 247.950 ;
        RECT 37.950 238.950 40.050 241.050 ;
        RECT 41.250 239.250 42.750 240.150 ;
        RECT 43.950 238.950 46.050 241.050 ;
        RECT 47.400 238.050 48.450 248.400 ;
        RECT 49.950 244.950 52.050 247.050 ;
        RECT 37.950 236.850 39.750 237.750 ;
        RECT 40.950 235.950 43.050 238.050 ;
        RECT 44.250 236.850 45.750 237.750 ;
        RECT 46.950 235.950 49.050 238.050 ;
        RECT 41.400 208.050 42.450 235.950 ;
        RECT 43.950 232.950 46.050 235.050 ;
        RECT 46.950 233.850 49.050 234.750 ;
        RECT 22.950 205.950 25.050 208.050 ;
        RECT 25.950 205.950 28.050 208.050 ;
        RECT 34.950 205.950 37.050 208.050 ;
        RECT 40.950 205.950 43.050 208.050 ;
        RECT 26.400 199.050 27.450 205.950 ;
        RECT 35.400 202.050 36.450 205.950 ;
        RECT 44.400 202.050 45.450 232.950 ;
        RECT 50.400 220.050 51.450 244.950 ;
        RECT 53.400 237.450 54.450 268.950 ;
        RECT 56.400 241.050 57.450 268.950 ;
        RECT 59.400 241.050 60.450 304.950 ;
        RECT 61.950 298.950 64.050 301.050 ;
        RECT 62.400 277.050 63.450 298.950 ;
        RECT 61.950 274.950 64.050 277.050 ;
        RECT 62.400 256.050 63.450 274.950 ;
        RECT 65.400 262.050 66.450 311.400 ;
        RECT 67.950 310.950 70.050 313.050 ;
        RECT 71.250 311.250 72.750 312.150 ;
        RECT 73.950 310.950 76.050 313.050 ;
        RECT 76.950 310.950 79.050 313.050 ;
        RECT 67.950 308.850 69.750 309.750 ;
        RECT 70.950 307.950 73.050 310.050 ;
        RECT 74.250 308.850 75.750 309.750 ;
        RECT 76.950 307.950 79.050 310.050 ;
        RECT 71.400 295.050 72.450 307.950 ;
        RECT 76.950 305.850 79.050 306.750 ;
        RECT 73.950 295.950 76.050 298.050 ;
        RECT 67.950 292.950 70.050 295.050 ;
        RECT 70.950 292.950 73.050 295.050 ;
        RECT 68.400 271.050 69.450 292.950 ;
        RECT 70.950 289.950 73.050 292.050 ;
        RECT 67.950 268.950 70.050 271.050 ;
        RECT 67.950 266.850 70.050 267.750 ;
        RECT 64.950 259.950 67.050 262.050 ;
        RECT 61.950 253.950 64.050 256.050 ;
        RECT 67.950 253.950 70.050 256.050 ;
        RECT 55.950 238.950 58.050 241.050 ;
        RECT 58.950 238.950 61.050 241.050 ;
        RECT 62.250 239.250 63.750 240.150 ;
        RECT 64.950 238.950 67.050 241.050 ;
        RECT 55.950 237.450 58.050 238.050 ;
        RECT 53.400 236.400 58.050 237.450 ;
        RECT 59.250 236.850 60.750 237.750 ;
        RECT 55.950 235.950 58.050 236.400 ;
        RECT 61.950 235.950 64.050 238.050 ;
        RECT 65.250 236.850 67.050 237.750 ;
        RECT 52.950 232.950 55.050 235.050 ;
        RECT 55.950 233.850 58.050 234.750 ;
        RECT 58.950 232.950 61.050 235.050 ;
        RECT 49.950 217.950 52.050 220.050 ;
        RECT 53.400 216.450 54.450 232.950 ;
        RECT 50.400 215.400 54.450 216.450 ;
        RECT 46.950 205.950 49.050 208.050 ;
        RECT 47.400 202.050 48.450 205.950 ;
        RECT 50.400 205.050 51.450 215.400 ;
        RECT 49.950 202.950 52.050 205.050 ;
        RECT 52.950 203.250 55.050 204.150 ;
        RECT 31.950 199.950 34.050 202.050 ;
        RECT 34.950 199.950 37.050 202.050 ;
        RECT 38.250 200.250 39.750 201.150 ;
        RECT 40.950 199.950 43.050 202.050 ;
        RECT 43.950 199.950 46.050 202.050 ;
        RECT 46.950 199.950 49.050 202.050 ;
        RECT 50.250 200.250 51.750 201.150 ;
        RECT 52.950 199.950 55.050 202.050 ;
        RECT 56.250 200.250 58.050 201.150 ;
        RECT 22.950 197.250 25.050 198.150 ;
        RECT 25.950 196.950 28.050 199.050 ;
        RECT 28.950 197.250 31.050 198.150 ;
        RECT 22.950 193.950 25.050 196.050 ;
        RECT 28.950 195.450 31.050 196.050 ;
        RECT 32.400 195.450 33.450 199.950 ;
        RECT 34.950 197.850 36.750 198.750 ;
        RECT 37.950 196.950 40.050 199.050 ;
        RECT 41.250 197.850 43.050 198.750 ;
        RECT 26.250 194.250 27.750 195.150 ;
        RECT 28.950 194.400 33.450 195.450 ;
        RECT 28.950 193.950 31.050 194.400 ;
        RECT 25.950 190.950 28.050 193.050 ;
        RECT 26.400 184.050 27.450 190.950 ;
        RECT 28.950 187.950 31.050 190.050 ;
        RECT 25.950 181.950 28.050 184.050 ;
        RECT 29.400 172.050 30.450 187.950 ;
        RECT 31.950 172.950 34.050 175.050 ;
        RECT 22.950 169.950 25.050 172.050 ;
        RECT 28.950 169.950 31.050 172.050 ;
        RECT 23.400 165.450 24.450 169.950 ;
        RECT 25.950 167.250 28.050 168.150 ;
        RECT 28.950 167.850 31.050 168.750 ;
        RECT 32.400 166.050 33.450 172.950 ;
        RECT 38.400 171.450 39.450 196.950 ;
        RECT 44.400 172.050 45.450 199.950 ;
        RECT 46.950 197.850 48.750 198.750 ;
        RECT 49.950 198.450 52.050 199.050 ;
        RECT 49.950 197.400 54.450 198.450 ;
        RECT 49.950 196.950 52.050 197.400 ;
        RECT 53.400 196.050 54.450 197.400 ;
        RECT 55.950 196.950 58.050 199.050 ;
        RECT 52.950 193.950 55.050 196.050 ;
        RECT 55.950 193.950 58.050 196.050 ;
        RECT 46.950 175.950 49.050 178.050 ;
        RECT 35.400 170.400 39.450 171.450 ;
        RECT 25.950 165.450 28.050 166.050 ;
        RECT 23.400 164.400 28.050 165.450 ;
        RECT 25.950 163.950 28.050 164.400 ;
        RECT 28.950 163.950 31.050 166.050 ;
        RECT 31.950 163.950 34.050 166.050 ;
        RECT 19.950 157.950 22.050 160.050 ;
        RECT 16.950 136.950 19.050 139.050 ;
        RECT 19.950 136.950 22.050 139.050 ;
        RECT 22.950 136.950 25.050 139.050 ;
        RECT 17.550 118.050 18.750 136.950 ;
        RECT 20.550 132.750 21.750 136.950 ;
        RECT 19.950 130.650 22.050 132.750 ;
        RECT 20.550 118.050 21.750 130.650 ;
        RECT 23.550 118.050 24.750 136.950 ;
        RECT 29.400 133.050 30.450 163.950 ;
        RECT 35.400 145.050 36.450 170.400 ;
        RECT 40.950 169.950 43.050 172.050 ;
        RECT 43.950 169.950 46.050 172.050 ;
        RECT 47.400 169.050 48.450 175.950 ;
        RECT 49.950 169.950 52.050 172.050 ;
        RECT 37.950 167.250 40.050 168.150 ;
        RECT 40.950 167.850 43.050 168.750 ;
        RECT 43.950 167.250 45.750 168.150 ;
        RECT 46.950 166.950 49.050 169.050 ;
        RECT 37.950 163.950 40.050 166.050 ;
        RECT 40.950 163.950 43.050 166.050 ;
        RECT 43.950 163.950 46.050 166.050 ;
        RECT 47.250 164.850 49.050 165.750 ;
        RECT 41.400 151.050 42.450 163.950 ;
        RECT 44.400 154.050 45.450 163.950 ;
        RECT 43.950 151.950 46.050 154.050 ;
        RECT 40.950 148.950 43.050 151.050 ;
        RECT 34.950 142.950 37.050 145.050 ;
        RECT 50.400 142.050 51.450 169.950 ;
        RECT 53.400 148.050 54.450 193.950 ;
        RECT 52.950 145.950 55.050 148.050 ;
        RECT 49.950 139.950 52.050 142.050 ;
        RECT 47.100 137.100 49.200 139.200 ;
        RECT 31.950 134.400 34.050 136.500 ;
        RECT 36.000 134.400 38.100 136.500 ;
        RECT 43.950 134.850 46.050 136.950 ;
        RECT 28.950 130.950 31.050 133.050 ;
        RECT 32.250 128.250 33.450 134.400 ;
        RECT 31.950 126.150 34.050 128.250 ;
        RECT 28.950 122.250 31.050 123.150 ;
        RECT 28.950 120.450 31.050 121.050 ;
        RECT 26.400 119.400 31.050 120.450 ;
        RECT 16.950 115.950 19.050 118.050 ;
        RECT 19.950 115.950 22.050 118.050 ;
        RECT 22.950 115.950 25.050 118.050 ;
        RECT 13.950 94.950 16.050 97.050 ;
        RECT 19.950 94.950 22.050 97.050 ;
        RECT 20.400 94.050 21.450 94.950 ;
        RECT 26.400 94.050 27.450 119.400 ;
        RECT 28.950 118.950 31.050 119.400 ;
        RECT 32.250 117.600 33.450 126.150 ;
        RECT 36.450 125.550 37.650 134.400 ;
        RECT 40.950 131.250 43.050 133.350 ;
        RECT 36.150 123.450 38.250 125.550 ;
        RECT 36.450 117.600 37.650 123.450 ;
        RECT 41.400 117.600 42.600 131.250 ;
        RECT 44.550 117.600 45.750 134.850 ;
        RECT 47.250 133.350 48.450 137.100 ;
        RECT 46.950 131.250 49.050 133.350 ;
        RECT 56.400 132.450 57.450 193.950 ;
        RECT 59.400 187.050 60.450 232.950 ;
        RECT 62.400 226.050 63.450 235.950 ;
        RECT 64.950 232.950 67.050 235.050 ;
        RECT 61.950 223.950 64.050 226.050 ;
        RECT 65.400 223.050 66.450 232.950 ;
        RECT 68.400 232.050 69.450 253.950 ;
        RECT 71.400 244.050 72.450 289.950 ;
        RECT 70.950 241.950 73.050 244.050 ;
        RECT 74.400 240.450 75.450 295.950 ;
        RECT 80.400 283.050 81.450 316.950 ;
        RECT 89.400 316.050 90.450 316.950 ;
        RECT 88.950 313.950 91.050 316.050 ;
        RECT 92.400 313.050 93.450 320.400 ;
        RECT 85.950 312.450 88.050 313.050 ;
        RECT 83.400 311.400 88.050 312.450 ;
        RECT 89.250 311.850 90.750 312.750 ;
        RECT 83.400 289.050 84.450 311.400 ;
        RECT 85.950 310.950 88.050 311.400 ;
        RECT 91.950 310.950 94.050 313.050 ;
        RECT 85.950 308.850 88.050 309.750 ;
        RECT 91.950 308.850 94.050 309.750 ;
        RECT 82.950 286.950 85.050 289.050 ;
        RECT 79.950 280.950 82.050 283.050 ;
        RECT 95.400 277.050 96.450 373.950 ;
        RECT 100.950 340.950 103.050 343.050 ;
        RECT 97.950 338.250 100.050 339.150 ;
        RECT 100.950 338.850 103.050 339.750 ;
        RECT 97.950 334.950 100.050 337.050 ;
        RECT 98.400 328.050 99.450 334.950 ;
        RECT 104.400 328.050 105.450 394.950 ;
        RECT 112.950 391.950 115.050 394.050 ;
        RECT 113.400 388.050 114.450 391.950 ;
        RECT 109.950 385.950 112.050 388.050 ;
        RECT 112.950 385.950 115.050 388.050 ;
        RECT 110.400 385.050 111.450 385.950 ;
        RECT 106.950 382.950 109.050 385.050 ;
        RECT 109.950 382.950 112.050 385.050 ;
        RECT 113.250 383.850 114.750 384.750 ;
        RECT 115.950 382.950 118.050 385.050 ;
        RECT 97.950 325.950 100.050 328.050 ;
        RECT 103.950 325.950 106.050 328.050 ;
        RECT 107.400 319.050 108.450 382.950 ;
        RECT 119.400 382.050 120.450 415.950 ;
        RECT 128.400 415.050 129.450 421.950 ;
        RECT 131.400 418.050 132.450 476.400 ;
        RECT 136.950 475.950 139.050 478.050 ;
        RECT 139.950 475.950 142.050 478.050 ;
        RECT 142.950 475.950 145.050 478.050 ;
        RECT 148.950 475.950 151.050 478.050 ;
        RECT 152.250 477.600 153.450 486.150 ;
        RECT 156.450 485.550 157.650 494.400 ;
        RECT 160.950 491.250 163.050 493.350 ;
        RECT 156.150 483.450 158.250 485.550 ;
        RECT 156.450 477.600 157.650 483.450 ;
        RECT 161.400 477.600 162.600 491.250 ;
        RECT 164.550 477.600 165.750 494.850 ;
        RECT 167.250 493.350 168.450 497.100 ;
        RECT 166.950 491.250 169.050 493.350 ;
        RECT 167.250 477.600 168.450 491.250 ;
        RECT 173.400 486.450 174.450 502.950 ;
        RECT 182.400 499.050 183.450 547.950 ;
        RECT 185.400 529.050 186.450 550.950 ;
        RECT 188.400 547.050 189.450 553.950 ;
        RECT 197.400 553.050 198.450 556.950 ;
        RECT 220.950 553.950 223.050 556.050 ;
        RECT 226.950 553.950 229.050 556.050 ;
        RECT 196.950 550.950 199.050 553.050 ;
        RECT 227.400 550.050 228.450 553.950 ;
        RECT 226.950 547.950 229.050 550.050 ;
        RECT 187.950 544.950 190.050 547.050 ;
        RECT 199.950 535.950 202.050 538.050 ;
        RECT 190.950 529.950 193.050 532.050 ;
        RECT 193.950 529.950 196.050 532.050 ;
        RECT 191.400 529.050 192.450 529.950 ;
        RECT 184.950 526.950 187.050 529.050 ;
        RECT 190.950 526.950 193.050 529.050 ;
        RECT 185.400 523.050 186.450 526.950 ;
        RECT 190.950 524.850 193.050 525.750 ;
        RECT 184.950 520.950 187.050 523.050 ;
        RECT 190.950 502.950 193.050 505.050 ;
        RECT 181.950 496.950 184.050 499.050 ;
        RECT 175.950 488.250 178.050 489.150 ;
        RECT 175.950 486.450 178.050 487.050 ;
        RECT 173.400 485.400 178.050 486.450 ;
        RECT 175.950 484.950 178.050 485.400 ;
        RECT 187.950 484.950 190.050 487.050 ;
        RECT 176.400 481.050 177.450 484.950 ;
        RECT 187.950 482.850 190.050 483.750 ;
        RECT 175.950 478.950 178.050 481.050 ;
        RECT 151.950 475.500 154.050 477.600 ;
        RECT 156.150 475.500 158.250 477.600 ;
        RECT 160.950 475.500 163.050 477.600 ;
        RECT 163.950 475.500 166.050 477.600 ;
        RECT 166.950 475.500 169.050 477.600 ;
        RECT 133.950 472.950 136.050 475.050 ;
        RECT 134.400 460.050 135.450 472.950 ;
        RECT 157.950 460.950 160.050 463.050 ;
        RECT 160.950 460.950 163.050 463.050 ;
        RECT 163.950 460.950 166.050 463.050 ;
        RECT 169.950 460.950 172.050 463.050 ;
        RECT 172.950 461.400 175.050 463.500 ;
        RECT 177.150 461.400 179.250 463.500 ;
        RECT 181.950 461.400 184.050 463.500 ;
        RECT 184.950 461.400 187.050 463.500 ;
        RECT 187.950 461.400 190.050 463.500 ;
        RECT 133.950 457.950 136.050 460.050 ;
        RECT 133.950 455.850 136.050 456.750 ;
        RECT 136.950 455.250 139.050 456.150 ;
        RECT 136.950 451.950 139.050 454.050 ;
        RECT 145.950 452.250 148.050 453.150 ;
        RECT 137.400 445.050 138.450 451.950 ;
        RECT 145.950 448.950 148.050 451.050 ;
        RECT 151.950 449.850 154.050 450.750 ;
        RECT 136.950 442.950 139.050 445.050 ;
        RECT 137.400 424.050 138.450 442.950 ;
        RECT 158.550 442.050 159.750 460.950 ;
        RECT 161.550 448.350 162.750 460.950 ;
        RECT 160.950 446.250 163.050 448.350 ;
        RECT 161.550 442.050 162.750 446.250 ;
        RECT 164.550 442.050 165.750 460.950 ;
        RECT 170.400 460.050 171.450 460.950 ;
        RECT 169.950 457.950 172.050 460.050 ;
        RECT 169.950 455.850 172.050 456.750 ;
        RECT 173.250 452.850 174.450 461.400 ;
        RECT 177.450 455.550 178.650 461.400 ;
        RECT 177.150 453.450 179.250 455.550 ;
        RECT 172.950 450.750 175.050 452.850 ;
        RECT 173.250 444.600 174.450 450.750 ;
        RECT 177.450 444.600 178.650 453.450 ;
        RECT 182.400 447.750 183.600 461.400 ;
        RECT 181.950 445.650 184.050 447.750 ;
        RECT 172.950 442.500 175.050 444.600 ;
        RECT 177.000 442.500 179.100 444.600 ;
        RECT 185.550 444.150 186.750 461.400 ;
        RECT 188.250 447.750 189.450 461.400 ;
        RECT 191.400 448.050 192.450 502.950 ;
        RECT 194.400 484.050 195.450 529.950 ;
        RECT 200.400 529.050 201.450 535.950 ;
        RECT 220.950 532.950 223.050 535.050 ;
        RECT 214.950 529.950 217.050 532.050 ;
        RECT 199.950 526.950 202.050 529.050 ;
        RECT 215.400 526.050 216.450 529.950 ;
        RECT 196.950 524.250 199.050 525.150 ;
        RECT 199.950 524.850 202.050 525.750 ;
        RECT 211.950 524.250 213.750 525.150 ;
        RECT 214.950 523.950 217.050 526.050 ;
        RECT 218.250 524.250 220.050 525.150 ;
        RECT 196.950 520.950 199.050 523.050 ;
        RECT 211.950 520.950 214.050 523.050 ;
        RECT 215.250 521.850 216.750 522.750 ;
        RECT 217.950 522.450 220.050 523.050 ;
        RECT 221.400 522.450 222.450 532.950 ;
        RECT 230.400 532.050 231.450 586.950 ;
        RECT 244.950 583.950 247.050 586.050 ;
        RECT 238.950 571.950 241.050 574.050 ;
        RECT 239.400 562.050 240.450 571.950 ;
        RECT 245.400 562.050 246.450 583.950 ;
        RECT 238.950 561.450 241.050 562.050 ;
        RECT 236.400 560.400 241.050 561.450 ;
        RECT 236.400 553.050 237.450 560.400 ;
        RECT 238.950 559.950 241.050 560.400 ;
        RECT 242.250 560.250 243.750 561.150 ;
        RECT 244.950 559.950 247.050 562.050 ;
        RECT 238.950 557.850 240.750 558.750 ;
        RECT 241.950 556.950 244.050 559.050 ;
        RECT 245.250 557.850 247.050 558.750 ;
        RECT 248.400 556.050 249.450 599.400 ;
        RECT 253.950 598.950 256.050 601.050 ;
        RECT 257.250 599.250 258.750 600.150 ;
        RECT 259.950 598.950 262.050 601.050 ;
        RECT 265.950 598.950 268.050 601.050 ;
        RECT 271.950 600.450 274.050 601.050 ;
        RECT 269.400 599.400 274.050 600.450 ;
        RECT 250.950 595.950 253.050 598.050 ;
        RECT 254.250 596.850 255.750 597.750 ;
        RECT 256.950 595.950 259.050 598.050 ;
        RECT 260.250 596.850 262.050 597.750 ;
        RECT 250.950 593.850 253.050 594.750 ;
        RECT 257.400 580.050 258.450 595.950 ;
        RECT 256.950 577.950 259.050 580.050 ;
        RECT 256.950 574.950 259.050 577.050 ;
        RECT 250.950 568.950 253.050 571.050 ;
        RECT 247.950 553.950 250.050 556.050 ;
        RECT 235.950 550.950 238.050 553.050 ;
        RECT 236.400 547.050 237.450 550.950 ;
        RECT 235.950 544.950 238.050 547.050 ;
        RECT 238.950 544.950 241.050 547.050 ;
        RECT 239.400 535.050 240.450 544.950 ;
        RECT 251.400 538.050 252.450 568.950 ;
        RECT 257.400 559.050 258.450 574.950 ;
        RECT 266.400 574.050 267.450 598.950 ;
        RECT 269.400 580.050 270.450 599.400 ;
        RECT 271.950 598.950 274.050 599.400 ;
        RECT 275.250 599.250 276.750 600.150 ;
        RECT 277.950 598.950 280.050 601.050 ;
        RECT 283.950 600.450 286.050 601.050 ;
        RECT 281.250 599.250 282.750 600.150 ;
        RECT 283.950 599.400 288.450 600.450 ;
        RECT 283.950 598.950 286.050 599.400 ;
        RECT 271.950 596.850 273.750 597.750 ;
        RECT 274.950 595.950 277.050 598.050 ;
        RECT 278.250 596.850 279.750 597.750 ;
        RECT 280.950 595.950 283.050 598.050 ;
        RECT 284.250 596.850 286.050 597.750 ;
        RECT 287.400 586.050 288.450 599.400 ;
        RECT 290.400 598.050 291.450 610.950 ;
        RECT 304.950 607.950 307.050 610.050 ;
        RECT 295.950 601.950 298.050 604.050 ;
        RECT 292.950 598.950 295.050 601.050 ;
        RECT 296.250 599.850 297.750 600.750 ;
        RECT 298.950 600.450 301.050 601.050 ;
        RECT 298.950 599.400 303.450 600.450 ;
        RECT 298.950 598.950 301.050 599.400 ;
        RECT 289.950 595.950 292.050 598.050 ;
        RECT 292.950 596.850 295.050 597.750 ;
        RECT 295.950 595.950 298.050 598.050 ;
        RECT 298.950 596.850 301.050 597.750 ;
        RECT 286.950 583.950 289.050 586.050 ;
        RECT 268.950 577.950 271.050 580.050 ;
        RECT 265.950 571.950 268.050 574.050 ;
        RECT 296.400 565.050 297.450 595.950 ;
        RECT 302.400 586.050 303.450 599.400 ;
        RECT 305.400 595.050 306.450 607.950 ;
        RECT 308.400 601.050 309.450 611.400 ;
        RECT 307.950 598.950 310.050 601.050 ;
        RECT 311.400 598.050 312.450 622.950 ;
        RECT 326.400 619.050 327.450 632.400 ;
        RECT 332.400 627.450 333.450 634.950 ;
        RECT 338.400 631.050 339.450 655.950 ;
        RECT 344.400 637.050 345.450 664.950 ;
        RECT 350.400 661.050 351.450 667.950 ;
        RECT 368.400 666.450 369.450 685.950 ;
        RECT 371.400 670.050 372.450 703.950 ;
        RECT 373.950 701.850 375.750 702.750 ;
        RECT 376.950 700.950 379.050 703.050 ;
        RECT 380.250 701.850 382.050 702.750 ;
        RECT 373.950 673.950 376.050 676.050 ;
        RECT 370.950 667.950 373.050 670.050 ;
        RECT 365.400 665.400 369.450 666.450 ;
        RECT 349.950 658.950 352.050 661.050 ;
        RECT 346.950 652.950 349.050 655.050 ;
        RECT 343.950 634.950 346.050 637.050 ;
        RECT 343.950 632.250 346.050 633.150 ;
        RECT 334.950 629.250 336.750 630.150 ;
        RECT 337.950 628.950 340.050 631.050 ;
        RECT 341.250 629.250 342.750 630.150 ;
        RECT 343.950 628.950 346.050 631.050 ;
        RECT 334.950 627.450 337.050 628.050 ;
        RECT 332.400 626.400 337.050 627.450 ;
        RECT 338.250 626.850 339.750 627.750 ;
        RECT 334.950 625.950 337.050 626.400 ;
        RECT 340.950 625.950 343.050 628.050 ;
        RECT 325.950 616.950 328.050 619.050 ;
        RECT 335.400 610.050 336.450 625.950 ;
        RECT 341.400 616.050 342.450 625.950 ;
        RECT 344.400 625.050 345.450 628.950 ;
        RECT 343.950 622.950 346.050 625.050 ;
        RECT 340.950 613.950 343.050 616.050 ;
        RECT 347.400 610.050 348.450 652.950 ;
        RECT 361.950 646.950 364.050 649.050 ;
        RECT 349.950 631.950 352.050 634.050 ;
        RECT 355.950 633.450 358.050 634.050 ;
        RECT 353.250 632.250 354.750 633.150 ;
        RECT 355.950 632.400 360.450 633.450 ;
        RECT 355.950 631.950 358.050 632.400 ;
        RECT 359.400 631.050 360.450 632.400 ;
        RECT 349.950 629.850 351.750 630.750 ;
        RECT 352.950 628.950 355.050 631.050 ;
        RECT 356.250 629.850 358.050 630.750 ;
        RECT 358.950 628.950 361.050 631.050 ;
        RECT 353.400 622.050 354.450 628.950 ;
        RECT 358.950 625.950 361.050 628.050 ;
        RECT 352.950 619.950 355.050 622.050 ;
        RECT 334.950 607.950 337.050 610.050 ;
        RECT 343.950 607.950 346.050 610.050 ;
        RECT 346.950 607.950 349.050 610.050 ;
        RECT 316.950 604.950 319.050 607.050 ;
        RECT 319.950 604.950 322.050 607.050 ;
        RECT 307.950 596.250 309.750 597.150 ;
        RECT 310.950 595.950 313.050 598.050 ;
        RECT 314.250 596.250 316.050 597.150 ;
        RECT 304.950 592.950 307.050 595.050 ;
        RECT 307.950 592.950 310.050 595.050 ;
        RECT 311.250 593.850 312.750 594.750 ;
        RECT 313.950 592.950 316.050 595.050 ;
        RECT 301.950 583.950 304.050 586.050 ;
        RECT 308.400 574.050 309.450 592.950 ;
        RECT 310.950 577.950 313.050 580.050 ;
        RECT 307.950 571.950 310.050 574.050 ;
        RECT 265.950 562.950 268.050 565.050 ;
        RECT 295.950 562.950 298.050 565.050 ;
        RECT 298.950 563.250 301.050 564.150 ;
        RECT 266.400 559.050 267.450 562.950 ;
        RECT 311.400 562.050 312.450 577.950 ;
        RECT 314.400 562.050 315.450 592.950 ;
        RECT 271.950 560.250 274.050 561.150 ;
        RECT 295.950 560.250 297.750 561.150 ;
        RECT 298.950 559.950 301.050 562.050 ;
        RECT 304.950 561.450 307.050 562.050 ;
        RECT 302.250 560.250 303.750 561.150 ;
        RECT 304.950 560.400 309.450 561.450 ;
        RECT 304.950 559.950 307.050 560.400 ;
        RECT 253.950 556.950 256.050 559.050 ;
        RECT 256.950 556.950 259.050 559.050 ;
        RECT 262.950 557.250 264.750 558.150 ;
        RECT 265.950 556.950 268.050 559.050 ;
        RECT 271.950 558.450 274.050 559.050 ;
        RECT 269.250 557.250 270.750 558.150 ;
        RECT 271.950 557.400 276.450 558.450 ;
        RECT 271.950 556.950 274.050 557.400 ;
        RECT 254.400 553.050 255.450 556.950 ;
        RECT 256.950 554.850 259.050 555.750 ;
        RECT 259.950 554.250 262.050 555.150 ;
        RECT 262.950 553.950 265.050 556.050 ;
        RECT 266.250 554.850 267.750 555.750 ;
        RECT 268.950 553.950 271.050 556.050 ;
        RECT 253.950 550.950 256.050 553.050 ;
        RECT 259.950 550.950 262.050 553.050 ;
        RECT 254.400 544.050 255.450 550.950 ;
        RECT 271.950 547.950 274.050 550.050 ;
        RECT 253.950 541.950 256.050 544.050 ;
        RECT 265.950 541.950 268.050 544.050 ;
        RECT 256.950 538.950 259.050 541.050 ;
        RECT 250.950 535.950 253.050 538.050 ;
        RECT 238.950 532.950 241.050 535.050 ;
        RECT 226.950 529.950 229.050 532.050 ;
        RECT 229.950 529.950 232.050 532.050 ;
        RECT 244.950 529.950 247.050 532.050 ;
        RECT 227.400 529.050 228.450 529.950 ;
        RECT 226.950 526.950 229.050 529.050 ;
        RECT 230.250 527.850 231.750 528.750 ;
        RECT 232.950 528.450 235.050 529.050 ;
        RECT 232.950 527.400 237.450 528.450 ;
        RECT 232.950 526.950 235.050 527.400 ;
        RECT 226.950 524.850 229.050 525.750 ;
        RECT 232.950 524.850 235.050 525.750 ;
        RECT 217.950 521.400 222.450 522.450 ;
        RECT 217.950 520.950 220.050 521.400 ;
        RECT 223.950 520.950 226.050 523.050 ;
        RECT 236.400 522.450 237.450 527.400 ;
        RECT 238.950 524.250 240.750 525.150 ;
        RECT 241.950 523.950 244.050 526.050 ;
        RECT 245.400 523.050 246.450 529.950 ;
        RECT 257.400 529.050 258.450 538.950 ;
        RECT 266.400 534.450 267.450 541.950 ;
        RECT 263.400 533.400 267.450 534.450 ;
        RECT 259.950 529.950 262.050 532.050 ;
        RECT 263.400 529.050 264.450 533.400 ;
        RECT 272.400 532.050 273.450 547.950 ;
        RECT 275.400 532.050 276.450 557.400 ;
        RECT 277.950 557.250 280.050 558.150 ;
        RECT 283.950 557.250 286.050 558.150 ;
        RECT 286.950 556.950 289.050 559.050 ;
        RECT 295.950 556.950 298.050 559.050 ;
        RECT 301.950 556.950 304.050 559.050 ;
        RECT 305.250 557.850 307.050 558.750 ;
        RECT 277.950 553.950 280.050 556.050 ;
        RECT 283.950 555.450 286.050 556.050 ;
        RECT 287.400 555.450 288.450 556.950 ;
        RECT 281.250 554.250 282.750 555.150 ;
        RECT 283.950 554.400 288.450 555.450 ;
        RECT 283.950 553.950 286.050 554.400 ;
        RECT 280.950 550.950 283.050 553.050 ;
        RECT 281.400 538.050 282.450 550.950 ;
        RECT 280.950 535.950 283.050 538.050 ;
        RECT 280.950 532.950 283.050 535.050 ;
        RECT 265.950 529.950 268.050 532.050 ;
        RECT 271.950 529.950 274.050 532.050 ;
        RECT 274.950 529.950 277.050 532.050 ;
        RECT 247.950 526.950 250.050 529.050 ;
        RECT 256.950 528.450 259.050 529.050 ;
        RECT 254.400 527.400 259.050 528.450 ;
        RECT 260.250 527.850 261.750 528.750 ;
        RECT 248.400 526.050 249.450 526.950 ;
        RECT 247.950 523.950 250.050 526.050 ;
        RECT 238.950 522.450 241.050 523.050 ;
        RECT 236.400 521.400 241.050 522.450 ;
        RECT 242.250 521.850 243.750 522.750 ;
        RECT 238.950 520.950 241.050 521.400 ;
        RECT 244.950 520.950 247.050 523.050 ;
        RECT 248.250 521.850 250.050 522.750 ;
        RECT 211.950 499.950 214.050 502.050 ;
        RECT 199.950 491.250 202.050 492.150 ;
        RECT 196.950 488.250 198.750 489.150 ;
        RECT 199.950 487.950 202.050 490.050 ;
        RECT 205.950 489.450 208.050 490.050 ;
        RECT 203.250 488.250 204.750 489.150 ;
        RECT 205.950 488.400 210.450 489.450 ;
        RECT 205.950 487.950 208.050 488.400 ;
        RECT 196.950 484.950 199.050 487.050 ;
        RECT 193.950 481.950 196.050 484.050 ;
        RECT 193.950 478.950 196.050 481.050 ;
        RECT 194.400 453.450 195.450 478.950 ;
        RECT 197.400 475.050 198.450 484.950 ;
        RECT 196.950 472.950 199.050 475.050 ;
        RECT 200.400 454.050 201.450 487.950 ;
        RECT 202.950 484.950 205.050 487.050 ;
        RECT 206.250 485.850 208.050 486.750 ;
        RECT 203.400 484.050 204.450 484.950 ;
        RECT 209.400 484.050 210.450 488.400 ;
        RECT 202.950 481.950 205.050 484.050 ;
        RECT 208.950 481.950 211.050 484.050 ;
        RECT 212.400 475.050 213.450 499.950 ;
        RECT 214.950 485.250 217.050 486.150 ;
        RECT 220.950 485.250 223.050 486.150 ;
        RECT 214.950 481.950 217.050 484.050 ;
        RECT 218.250 482.250 219.750 483.150 ;
        RECT 220.950 481.950 223.050 484.050 ;
        RECT 211.950 472.950 214.050 475.050 ;
        RECT 208.950 455.250 211.050 456.150 ;
        RECT 196.950 453.450 199.050 454.050 ;
        RECT 194.400 452.400 199.050 453.450 ;
        RECT 187.950 445.650 190.050 447.750 ;
        RECT 190.950 445.950 193.050 448.050 ;
        RECT 184.950 442.050 187.050 444.150 ;
        RECT 157.950 439.950 160.050 442.050 ;
        RECT 160.950 439.950 163.050 442.050 ;
        RECT 163.950 439.950 166.050 442.050 ;
        RECT 188.250 441.900 189.450 445.650 ;
        RECT 188.100 439.800 190.200 441.900 ;
        RECT 181.950 436.950 184.050 439.050 ;
        RECT 184.950 436.950 187.050 439.050 ;
        RECT 175.950 433.950 178.050 436.050 ;
        RECT 133.950 421.950 136.050 424.050 ;
        RECT 136.950 421.950 139.050 424.050 ;
        RECT 130.950 415.950 133.050 418.050 ;
        RECT 121.950 412.950 124.050 415.050 ;
        RECT 125.250 413.250 126.750 414.150 ;
        RECT 127.950 412.950 130.050 415.050 ;
        RECT 131.250 413.250 133.050 414.150 ;
        RECT 122.400 412.050 123.450 412.950 ;
        RECT 134.400 412.050 135.450 421.950 ;
        RECT 136.950 418.950 139.050 421.050 ;
        RECT 166.950 419.250 169.050 420.150 ;
        RECT 121.950 409.950 124.050 412.050 ;
        RECT 124.950 409.950 127.050 412.050 ;
        RECT 128.250 410.850 129.750 411.750 ;
        RECT 130.950 409.950 133.050 412.050 ;
        RECT 133.950 409.950 136.050 412.050 ;
        RECT 125.400 409.050 126.450 409.950 ;
        RECT 124.950 406.950 127.050 409.050 ;
        RECT 131.400 403.050 132.450 409.950 ;
        RECT 137.400 408.450 138.450 418.950 ;
        RECT 163.950 416.250 165.750 417.150 ;
        RECT 166.950 415.950 169.050 418.050 ;
        RECT 170.250 416.250 171.750 417.150 ;
        RECT 172.950 415.950 175.050 418.050 ;
        RECT 139.950 413.250 142.050 414.150 ;
        RECT 145.950 413.250 148.050 414.150 ;
        RECT 148.950 412.950 151.050 415.050 ;
        RECT 151.950 412.950 154.050 415.050 ;
        RECT 155.250 413.250 157.050 414.150 ;
        RECT 163.950 412.950 166.050 415.050 ;
        RECT 139.950 409.950 142.050 412.050 ;
        RECT 143.250 410.250 144.750 411.150 ;
        RECT 145.950 409.950 148.050 412.050 ;
        RECT 146.400 409.050 147.450 409.950 ;
        RECT 142.950 408.450 145.050 409.050 ;
        RECT 137.400 407.400 145.050 408.450 ;
        RECT 142.950 406.950 145.050 407.400 ;
        RECT 145.950 406.950 148.050 409.050 ;
        RECT 121.950 400.950 124.050 403.050 ;
        RECT 130.950 400.950 133.050 403.050 ;
        RECT 109.950 380.850 112.050 381.750 ;
        RECT 115.950 380.850 118.050 381.750 ;
        RECT 118.950 379.950 121.050 382.050 ;
        RECT 119.400 373.050 120.450 379.950 ;
        RECT 122.400 373.050 123.450 400.950 ;
        RECT 142.950 397.950 145.050 400.050 ;
        RECT 127.950 385.950 130.050 388.050 ;
        RECT 124.950 382.950 127.050 385.050 ;
        RECT 128.250 383.850 129.750 384.750 ;
        RECT 130.950 384.450 133.050 385.050 ;
        RECT 130.950 383.400 135.450 384.450 ;
        RECT 130.950 382.950 133.050 383.400 ;
        RECT 124.950 380.850 127.050 381.750 ;
        RECT 130.950 380.850 133.050 381.750 ;
        RECT 118.950 370.950 121.050 373.050 ;
        RECT 121.950 370.950 124.050 373.050 ;
        RECT 121.950 361.950 124.050 364.050 ;
        RECT 115.950 347.250 118.050 348.150 ;
        RECT 122.400 346.050 123.450 361.950 ;
        RECT 127.950 349.950 130.050 352.050 ;
        RECT 124.950 346.950 127.050 349.050 ;
        RECT 112.950 344.250 114.750 345.150 ;
        RECT 115.950 343.950 118.050 346.050 ;
        RECT 119.250 344.250 120.750 345.150 ;
        RECT 121.950 343.950 124.050 346.050 ;
        RECT 116.400 343.050 117.450 343.950 ;
        RECT 112.950 340.950 115.050 343.050 ;
        RECT 115.950 340.950 118.050 343.050 ;
        RECT 118.950 340.950 121.050 343.050 ;
        RECT 122.250 341.850 124.050 342.750 ;
        RECT 113.400 337.050 114.450 340.950 ;
        RECT 112.950 334.950 115.050 337.050 ;
        RECT 115.950 319.950 118.050 322.050 ;
        RECT 106.950 316.950 109.050 319.050 ;
        RECT 97.950 313.950 100.050 316.050 ;
        RECT 109.950 313.950 112.050 316.050 ;
        RECT 82.950 275.250 85.050 276.150 ;
        RECT 88.950 274.950 91.050 277.050 ;
        RECT 94.950 274.950 97.050 277.050 ;
        RECT 76.950 271.950 79.050 274.050 ;
        RECT 80.250 272.250 81.750 273.150 ;
        RECT 82.950 271.950 85.050 274.050 ;
        RECT 86.250 272.250 88.050 273.150 ;
        RECT 76.950 269.850 78.750 270.750 ;
        RECT 79.950 270.450 82.050 271.050 ;
        RECT 79.950 269.400 84.450 270.450 ;
        RECT 79.950 268.950 82.050 269.400 ;
        RECT 79.950 265.950 82.050 268.050 ;
        RECT 76.950 253.950 79.050 256.050 ;
        RECT 71.400 239.400 75.450 240.450 ;
        RECT 71.400 238.050 72.450 239.400 ;
        RECT 77.400 238.050 78.450 253.950 ;
        RECT 80.400 238.050 81.450 265.950 ;
        RECT 83.400 265.050 84.450 269.400 ;
        RECT 85.950 268.950 88.050 271.050 ;
        RECT 82.950 262.950 85.050 265.050 ;
        RECT 86.400 259.050 87.450 268.950 ;
        RECT 85.950 256.950 88.050 259.050 ;
        RECT 85.950 238.950 88.050 241.050 ;
        RECT 70.950 235.950 73.050 238.050 ;
        RECT 73.950 235.950 76.050 238.050 ;
        RECT 76.950 235.950 79.050 238.050 ;
        RECT 79.950 235.950 82.050 238.050 ;
        RECT 83.250 236.250 85.050 237.150 ;
        RECT 70.950 232.950 73.050 235.050 ;
        RECT 73.950 233.850 75.750 234.750 ;
        RECT 76.950 232.950 79.050 235.050 ;
        RECT 80.250 233.850 81.750 234.750 ;
        RECT 82.950 232.950 85.050 235.050 ;
        RECT 67.950 229.950 70.050 232.050 ;
        RECT 71.400 229.050 72.450 232.950 ;
        RECT 76.950 230.850 79.050 231.750 ;
        RECT 70.950 226.950 73.050 229.050 ;
        RECT 76.950 226.950 79.050 229.050 ;
        RECT 64.950 220.950 67.050 223.050 ;
        RECT 61.950 217.950 64.050 220.050 ;
        RECT 64.950 217.950 67.050 220.050 ;
        RECT 58.950 184.950 61.050 187.050 ;
        RECT 62.400 172.050 63.450 217.950 ;
        RECT 65.400 205.050 66.450 217.950 ;
        RECT 70.950 208.950 73.050 211.050 ;
        RECT 73.950 208.950 76.050 211.050 ;
        RECT 71.400 205.050 72.450 208.950 ;
        RECT 64.950 202.950 67.050 205.050 ;
        RECT 70.950 202.950 73.050 205.050 ;
        RECT 65.400 202.050 66.450 202.950 ;
        RECT 71.400 202.050 72.450 202.950 ;
        RECT 74.400 202.050 75.450 208.950 ;
        RECT 64.950 199.950 67.050 202.050 ;
        RECT 68.250 200.250 69.750 201.150 ;
        RECT 70.950 199.950 73.050 202.050 ;
        RECT 73.950 199.950 76.050 202.050 ;
        RECT 64.950 197.850 66.750 198.750 ;
        RECT 67.950 196.950 70.050 199.050 ;
        RECT 71.250 197.850 73.050 198.750 ;
        RECT 68.400 193.050 69.450 196.950 ;
        RECT 77.400 196.050 78.450 226.950 ;
        RECT 79.950 205.950 82.050 208.050 ;
        RECT 80.400 201.450 81.450 205.950 ;
        RECT 83.400 205.050 84.450 232.950 ;
        RECT 86.400 214.050 87.450 238.950 ;
        RECT 89.400 223.050 90.450 274.950 ;
        RECT 91.950 268.950 94.050 271.050 ;
        RECT 95.250 269.250 97.050 270.150 ;
        RECT 91.950 266.850 93.750 267.750 ;
        RECT 94.950 265.950 97.050 268.050 ;
        RECT 91.950 247.950 94.050 250.050 ;
        RECT 92.400 243.450 93.450 247.950 ;
        RECT 95.400 247.050 96.450 265.950 ;
        RECT 98.400 256.050 99.450 313.950 ;
        RECT 116.400 313.050 117.450 319.950 ;
        RECT 125.400 316.050 126.450 346.950 ;
        RECT 128.400 343.050 129.450 349.950 ;
        RECT 134.400 349.050 135.450 383.400 ;
        RECT 143.400 382.050 144.450 397.950 ;
        RECT 139.950 380.250 141.750 381.150 ;
        RECT 142.950 379.950 145.050 382.050 ;
        RECT 146.250 380.250 148.050 381.150 ;
        RECT 139.950 376.950 142.050 379.050 ;
        RECT 143.250 377.850 144.750 378.750 ;
        RECT 145.950 376.950 148.050 379.050 ;
        RECT 140.400 373.050 141.450 376.950 ;
        RECT 146.400 376.050 147.450 376.950 ;
        RECT 145.950 373.950 148.050 376.050 ;
        RECT 139.950 370.950 142.050 373.050 ;
        RECT 142.950 367.950 145.050 370.050 ;
        RECT 130.950 346.950 133.050 349.050 ;
        RECT 133.950 346.950 136.050 349.050 ;
        RECT 139.950 346.950 142.050 349.050 ;
        RECT 127.950 340.950 130.050 343.050 ;
        RECT 131.400 340.050 132.450 346.950 ;
        RECT 140.400 346.050 141.450 346.950 ;
        RECT 133.950 343.950 136.050 346.050 ;
        RECT 137.250 344.250 138.750 345.150 ;
        RECT 139.950 343.950 142.050 346.050 ;
        RECT 133.950 341.850 135.750 342.750 ;
        RECT 136.950 340.950 139.050 343.050 ;
        RECT 140.250 341.850 142.050 342.750 ;
        RECT 137.400 340.050 138.450 340.950 ;
        RECT 130.950 337.950 133.050 340.050 ;
        RECT 136.950 337.950 139.050 340.050 ;
        RECT 118.950 313.950 121.050 316.050 ;
        RECT 124.950 313.950 127.050 316.050 ;
        RECT 103.950 310.950 106.050 313.050 ;
        RECT 107.250 311.250 109.050 312.150 ;
        RECT 109.950 311.850 112.050 312.750 ;
        RECT 112.950 311.250 115.050 312.150 ;
        RECT 115.950 310.950 118.050 313.050 ;
        RECT 119.250 311.850 120.750 312.750 ;
        RECT 121.950 312.450 124.050 313.050 ;
        RECT 121.950 311.400 126.450 312.450 ;
        RECT 121.950 310.950 124.050 311.400 ;
        RECT 103.950 308.850 105.750 309.750 ;
        RECT 106.950 309.450 109.050 310.050 ;
        RECT 109.950 309.450 112.050 310.050 ;
        RECT 106.950 308.400 112.050 309.450 ;
        RECT 106.950 307.950 109.050 308.400 ;
        RECT 109.950 307.950 112.050 308.400 ;
        RECT 112.950 307.950 115.050 310.050 ;
        RECT 115.950 308.850 118.050 309.750 ;
        RECT 118.950 307.950 121.050 310.050 ;
        RECT 121.950 308.850 124.050 309.750 ;
        RECT 113.400 307.050 114.450 307.950 ;
        RECT 103.950 304.950 106.050 307.050 ;
        RECT 112.950 304.950 115.050 307.050 ;
        RECT 100.950 280.950 103.050 283.050 ;
        RECT 101.400 265.050 102.450 280.950 ;
        RECT 100.950 262.950 103.050 265.050 ;
        RECT 104.400 259.050 105.450 304.950 ;
        RECT 113.400 283.050 114.450 304.950 ;
        RECT 112.950 280.950 115.050 283.050 ;
        RECT 112.950 274.950 115.050 277.050 ;
        RECT 113.400 271.050 114.450 274.950 ;
        RECT 119.400 274.050 120.450 307.950 ;
        RECT 125.400 301.050 126.450 311.400 ;
        RECT 136.950 310.950 139.050 313.050 ;
        RECT 137.400 310.050 138.450 310.950 ;
        RECT 143.400 310.050 144.450 367.950 ;
        RECT 146.400 349.050 147.450 373.950 ;
        RECT 149.400 349.050 150.450 412.950 ;
        RECT 164.400 412.050 165.450 412.950 ;
        RECT 167.400 412.050 168.450 415.950 ;
        RECT 169.950 412.950 172.050 415.050 ;
        RECT 173.250 413.850 175.050 414.750 ;
        RECT 151.950 410.850 153.750 411.750 ;
        RECT 154.950 409.950 157.050 412.050 ;
        RECT 163.950 409.950 166.050 412.050 ;
        RECT 166.950 409.950 169.050 412.050 ;
        RECT 172.950 409.950 175.050 412.050 ;
        RECT 151.950 406.950 154.050 409.050 ;
        RECT 152.400 373.050 153.450 406.950 ;
        RECT 155.400 406.050 156.450 409.950 ;
        RECT 154.950 403.950 157.050 406.050 ;
        RECT 155.400 376.050 156.450 403.950 ;
        RECT 163.950 391.950 166.050 394.050 ;
        RECT 166.950 391.950 169.050 394.050 ;
        RECT 164.400 388.050 165.450 391.950 ;
        RECT 163.950 385.950 166.050 388.050 ;
        RECT 157.950 382.950 160.050 385.050 ;
        RECT 160.950 383.250 163.050 384.150 ;
        RECT 163.950 383.850 166.050 384.750 ;
        RECT 158.400 376.050 159.450 382.950 ;
        RECT 160.950 379.950 163.050 382.050 ;
        RECT 163.950 379.950 166.050 382.050 ;
        RECT 154.950 373.950 157.050 376.050 ;
        RECT 157.950 375.450 160.050 376.050 ;
        RECT 161.400 375.450 162.450 379.950 ;
        RECT 164.400 376.050 165.450 379.950 ;
        RECT 157.950 374.400 162.450 375.450 ;
        RECT 157.950 373.950 160.050 374.400 ;
        RECT 163.950 373.950 166.050 376.050 ;
        RECT 151.950 370.950 154.050 373.050 ;
        RECT 164.400 370.050 165.450 373.950 ;
        RECT 163.950 367.950 166.050 370.050 ;
        RECT 167.400 349.050 168.450 391.950 ;
        RECT 173.400 382.050 174.450 409.950 ;
        RECT 176.400 400.050 177.450 433.950 ;
        RECT 182.400 418.050 183.450 436.950 ;
        RECT 178.950 415.950 181.050 418.050 ;
        RECT 181.950 415.950 184.050 418.050 ;
        RECT 175.950 397.950 178.050 400.050 ;
        RECT 169.950 380.250 171.750 381.150 ;
        RECT 172.950 379.950 175.050 382.050 ;
        RECT 176.250 380.250 178.050 381.150 ;
        RECT 169.950 376.950 172.050 379.050 ;
        RECT 173.250 377.850 174.750 378.750 ;
        RECT 175.950 376.950 178.050 379.050 ;
        RECT 170.400 376.050 171.450 376.950 ;
        RECT 169.950 373.950 172.050 376.050 ;
        RECT 176.400 373.050 177.450 376.950 ;
        RECT 172.950 370.950 175.050 373.050 ;
        RECT 175.950 370.950 178.050 373.050 ;
        RECT 145.950 346.950 148.050 349.050 ;
        RECT 148.950 346.950 151.050 349.050 ;
        RECT 157.950 346.950 160.050 349.050 ;
        RECT 160.950 346.950 163.050 349.050 ;
        RECT 166.950 346.950 169.050 349.050 ;
        RECT 146.400 322.050 147.450 346.950 ;
        RECT 148.950 343.950 151.050 346.050 ;
        RECT 152.250 344.250 153.750 345.150 ;
        RECT 154.950 343.950 157.050 346.050 ;
        RECT 148.950 341.850 150.750 342.750 ;
        RECT 151.950 340.950 154.050 343.050 ;
        RECT 155.250 341.850 157.050 342.750 ;
        RECT 145.950 319.950 148.050 322.050 ;
        RECT 127.950 307.950 130.050 310.050 ;
        RECT 133.950 308.250 135.750 309.150 ;
        RECT 136.950 307.950 139.050 310.050 ;
        RECT 140.250 308.250 142.050 309.150 ;
        RECT 142.950 307.950 145.050 310.050 ;
        RECT 124.950 298.950 127.050 301.050 ;
        RECT 121.950 280.950 124.050 283.050 ;
        RECT 118.950 271.950 121.050 274.050 ;
        RECT 122.400 271.050 123.450 280.950 ;
        RECT 109.950 269.250 112.050 270.150 ;
        RECT 112.950 268.950 115.050 271.050 ;
        RECT 115.950 269.250 118.050 270.150 ;
        RECT 118.950 269.250 121.050 270.150 ;
        RECT 121.950 268.950 124.050 271.050 ;
        RECT 124.950 269.250 127.050 270.150 ;
        RECT 128.400 268.050 129.450 307.950 ;
        RECT 130.950 304.950 133.050 307.050 ;
        RECT 133.950 304.950 136.050 307.050 ;
        RECT 137.250 305.850 138.750 306.750 ;
        RECT 139.950 304.950 142.050 307.050 ;
        RECT 131.400 277.050 132.450 304.950 ;
        RECT 134.400 301.050 135.450 304.950 ;
        RECT 140.400 304.050 141.450 304.950 ;
        RECT 146.400 304.050 147.450 319.950 ;
        RECT 152.400 313.050 153.450 340.950 ;
        RECT 154.950 334.950 157.050 337.050 ;
        RECT 155.400 313.050 156.450 334.950 ;
        RECT 158.400 319.050 159.450 346.950 ;
        RECT 161.400 346.050 162.450 346.950 ;
        RECT 160.950 343.950 163.050 346.050 ;
        RECT 166.950 345.450 169.050 346.050 ;
        RECT 164.250 344.250 165.750 345.150 ;
        RECT 166.950 344.400 171.450 345.450 ;
        RECT 166.950 343.950 169.050 344.400 ;
        RECT 160.950 341.850 162.750 342.750 ;
        RECT 163.950 340.950 166.050 343.050 ;
        RECT 167.250 341.850 169.050 342.750 ;
        RECT 160.950 337.950 163.050 340.050 ;
        RECT 163.950 337.950 166.050 340.050 ;
        RECT 170.400 339.450 171.450 344.400 ;
        RECT 167.400 338.400 171.450 339.450 ;
        RECT 157.950 316.950 160.050 319.050 ;
        RECT 151.950 310.950 154.050 313.050 ;
        RECT 154.950 310.950 157.050 313.050 ;
        RECT 152.400 310.050 153.450 310.950 ;
        RECT 161.400 310.050 162.450 337.950 ;
        RECT 164.400 334.050 165.450 337.950 ;
        RECT 167.400 337.050 168.450 338.400 ;
        RECT 166.950 334.950 169.050 337.050 ;
        RECT 163.950 331.950 166.050 334.050 ;
        RECT 164.400 316.050 165.450 331.950 ;
        RECT 173.400 319.050 174.450 370.950 ;
        RECT 179.400 346.050 180.450 415.950 ;
        RECT 182.400 415.050 183.450 415.950 ;
        RECT 181.950 412.950 184.050 415.050 ;
        RECT 181.950 410.850 184.050 411.750 ;
        RECT 185.400 394.050 186.450 436.950 ;
        RECT 194.400 420.450 195.450 452.400 ;
        RECT 196.950 451.950 199.050 452.400 ;
        RECT 199.950 451.950 202.050 454.050 ;
        RECT 208.950 451.950 211.050 454.050 ;
        RECT 196.950 449.850 199.050 450.750 ;
        RECT 196.950 445.950 199.050 448.050 ;
        RECT 191.400 419.400 195.450 420.450 ;
        RECT 191.400 414.450 192.450 419.400 ;
        RECT 193.950 416.250 196.050 417.150 ;
        RECT 193.950 414.450 196.050 415.050 ;
        RECT 191.400 413.400 196.050 414.450 ;
        RECT 193.950 412.950 196.050 413.400 ;
        RECT 187.950 400.950 190.050 403.050 ;
        RECT 184.950 391.950 187.050 394.050 ;
        RECT 188.400 382.050 189.450 400.950 ;
        RECT 197.400 394.050 198.450 445.950 ;
        RECT 215.400 436.050 216.450 481.950 ;
        RECT 224.400 481.050 225.450 520.950 ;
        RECT 254.400 520.050 255.450 527.400 ;
        RECT 256.950 526.950 259.050 527.400 ;
        RECT 262.950 526.950 265.050 529.050 ;
        RECT 256.950 524.850 259.050 525.750 ;
        RECT 262.950 524.850 265.050 525.750 ;
        RECT 244.950 518.850 247.050 519.750 ;
        RECT 253.950 517.950 256.050 520.050 ;
        RECT 238.950 508.950 241.050 511.050 ;
        RECT 239.400 490.050 240.450 508.950 ;
        RECT 244.950 502.950 247.050 505.050 ;
        RECT 250.950 502.950 253.050 505.050 ;
        RECT 229.950 487.950 232.050 490.050 ;
        RECT 232.950 488.250 235.050 489.150 ;
        RECT 238.950 487.950 241.050 490.050 ;
        RECT 217.950 478.950 220.050 481.050 ;
        RECT 223.950 478.950 226.050 481.050 ;
        RECT 230.400 475.050 231.450 487.950 ;
        RECT 239.400 487.050 240.450 487.950 ;
        RECT 232.950 484.950 235.050 487.050 ;
        RECT 236.250 485.250 237.750 486.150 ;
        RECT 238.950 484.950 241.050 487.050 ;
        RECT 242.250 485.250 244.050 486.150 ;
        RECT 233.400 481.050 234.450 484.950 ;
        RECT 235.950 481.950 238.050 484.050 ;
        RECT 239.250 482.850 240.750 483.750 ;
        RECT 241.950 481.950 244.050 484.050 ;
        RECT 232.950 478.950 235.050 481.050 ;
        RECT 236.400 478.050 237.450 481.950 ;
        RECT 242.400 478.050 243.450 481.950 ;
        RECT 235.950 475.950 238.050 478.050 ;
        RECT 241.950 475.950 244.050 478.050 ;
        RECT 229.950 472.950 232.050 475.050 ;
        RECT 235.950 472.950 238.050 475.050 ;
        RECT 220.950 469.950 223.050 472.050 ;
        RECT 217.950 463.950 220.050 466.050 ;
        RECT 214.950 433.950 217.050 436.050 ;
        RECT 218.400 430.050 219.450 463.950 ;
        RECT 221.400 439.050 222.450 469.950 ;
        RECT 232.950 466.950 235.050 469.050 ;
        RECT 226.950 460.950 229.050 463.050 ;
        RECT 223.950 457.950 226.050 460.050 ;
        RECT 224.400 454.050 225.450 457.950 ;
        RECT 227.400 457.050 228.450 460.950 ;
        RECT 233.400 457.050 234.450 466.950 ;
        RECT 226.950 454.950 229.050 457.050 ;
        RECT 230.250 455.250 231.750 456.150 ;
        RECT 232.950 454.950 235.050 457.050 ;
        RECT 223.950 451.950 226.050 454.050 ;
        RECT 227.250 452.850 228.750 453.750 ;
        RECT 229.950 451.950 232.050 454.050 ;
        RECT 233.250 452.850 235.050 453.750 ;
        RECT 223.950 449.850 226.050 450.750 ;
        RECT 220.950 436.950 223.050 439.050 ;
        RECT 230.400 433.050 231.450 451.950 ;
        RECT 236.400 433.050 237.450 472.950 ;
        RECT 245.400 463.050 246.450 502.950 ;
        RECT 251.400 487.050 252.450 502.950 ;
        RECT 262.950 496.950 265.050 499.050 ;
        RECT 256.950 488.250 259.050 489.150 ;
        RECT 259.950 487.950 262.050 490.050 ;
        RECT 247.950 485.250 249.750 486.150 ;
        RECT 250.950 484.950 253.050 487.050 ;
        RECT 254.250 485.250 255.750 486.150 ;
        RECT 256.950 484.950 259.050 487.050 ;
        RECT 247.950 481.950 250.050 484.050 ;
        RECT 251.250 482.850 252.750 483.750 ;
        RECT 253.950 481.950 256.050 484.050 ;
        RECT 248.400 466.050 249.450 481.950 ;
        RECT 254.400 481.050 255.450 481.950 ;
        RECT 253.950 478.950 256.050 481.050 ;
        RECT 247.950 463.950 250.050 466.050 ;
        RECT 238.950 460.950 241.050 463.050 ;
        RECT 244.950 460.950 247.050 463.050 ;
        RECT 239.400 451.050 240.450 460.950 ;
        RECT 244.950 457.950 247.050 460.050 ;
        RECT 248.400 459.450 249.450 463.950 ;
        RECT 257.400 460.050 258.450 484.950 ;
        RECT 260.400 478.050 261.450 487.950 ;
        RECT 263.400 484.050 264.450 496.950 ;
        RECT 262.950 481.950 265.050 484.050 ;
        RECT 262.950 478.950 265.050 481.050 ;
        RECT 259.950 475.950 262.050 478.050 ;
        RECT 263.400 472.050 264.450 478.950 ;
        RECT 262.950 469.950 265.050 472.050 ;
        RECT 266.400 466.050 267.450 529.950 ;
        RECT 281.400 529.050 282.450 532.950 ;
        RECT 296.400 529.050 297.450 556.950 ;
        RECT 302.400 553.050 303.450 556.950 ;
        RECT 308.400 556.050 309.450 560.400 ;
        RECT 310.950 559.950 313.050 562.050 ;
        RECT 313.950 559.950 316.050 562.050 ;
        RECT 317.400 559.050 318.450 604.950 ;
        RECT 320.400 604.050 321.450 604.950 ;
        RECT 319.950 601.950 322.050 604.050 ;
        RECT 340.950 601.950 343.050 604.050 ;
        RECT 341.400 601.050 342.450 601.950 ;
        RECT 344.400 601.050 345.450 607.950 ;
        RECT 347.400 607.050 348.450 607.950 ;
        RECT 346.950 604.950 349.050 607.050 ;
        RECT 346.950 601.950 349.050 604.050 ;
        RECT 319.950 599.850 322.050 600.750 ;
        RECT 334.950 600.450 337.050 601.050 ;
        RECT 322.950 599.250 325.050 600.150 ;
        RECT 332.400 599.400 337.050 600.450 ;
        RECT 322.950 595.950 325.050 598.050 ;
        RECT 332.400 580.050 333.450 599.400 ;
        RECT 334.950 598.950 337.050 599.400 ;
        RECT 338.250 599.250 339.750 600.150 ;
        RECT 340.950 598.950 343.050 601.050 ;
        RECT 343.950 598.950 346.050 601.050 ;
        RECT 344.400 598.050 345.450 598.950 ;
        RECT 334.950 596.850 336.750 597.750 ;
        RECT 337.950 595.950 340.050 598.050 ;
        RECT 341.250 596.850 342.750 597.750 ;
        RECT 343.950 595.950 346.050 598.050 ;
        RECT 331.950 577.950 334.050 580.050 ;
        RECT 338.400 577.050 339.450 595.950 ;
        RECT 343.950 593.850 346.050 594.750 ;
        RECT 347.400 594.450 348.450 601.950 ;
        RECT 352.950 598.950 355.050 601.050 ;
        RECT 353.400 598.050 354.450 598.950 ;
        RECT 349.950 596.250 351.750 597.150 ;
        RECT 352.950 595.950 355.050 598.050 ;
        RECT 356.250 596.250 358.050 597.150 ;
        RECT 349.950 594.450 352.050 595.050 ;
        RECT 347.400 593.400 352.050 594.450 ;
        RECT 353.250 593.850 354.750 594.750 ;
        RECT 349.950 592.950 352.050 593.400 ;
        RECT 355.950 592.950 358.050 595.050 ;
        RECT 337.950 574.950 340.050 577.050 ;
        RECT 340.950 574.950 343.050 577.050 ;
        RECT 337.950 571.950 340.050 574.050 ;
        RECT 331.950 563.250 334.050 564.150 ;
        RECT 325.950 561.450 328.050 562.050 ;
        RECT 323.400 560.400 328.050 561.450 ;
        RECT 313.950 557.250 316.050 558.150 ;
        RECT 316.950 556.950 319.050 559.050 ;
        RECT 319.950 557.250 322.050 558.150 ;
        RECT 307.950 553.950 310.050 556.050 ;
        RECT 313.950 553.950 316.050 556.050 ;
        RECT 319.950 555.450 322.050 556.050 ;
        RECT 323.400 555.450 324.450 560.400 ;
        RECT 325.950 559.950 328.050 560.400 ;
        RECT 329.250 560.250 330.750 561.150 ;
        RECT 331.950 559.950 334.050 562.050 ;
        RECT 335.250 560.250 337.050 561.150 ;
        RECT 332.400 559.050 333.450 559.950 ;
        RECT 325.950 557.850 327.750 558.750 ;
        RECT 328.950 556.950 331.050 559.050 ;
        RECT 331.950 556.950 334.050 559.050 ;
        RECT 334.950 556.950 337.050 559.050 ;
        RECT 317.250 554.250 318.750 555.150 ;
        RECT 319.950 554.400 324.450 555.450 ;
        RECT 319.950 553.950 322.050 554.400 ;
        RECT 329.400 553.050 330.450 556.950 ;
        RECT 335.400 556.050 336.450 556.950 ;
        RECT 334.950 553.950 337.050 556.050 ;
        RECT 301.950 550.950 304.050 553.050 ;
        RECT 307.950 550.950 310.050 553.050 ;
        RECT 316.950 550.950 319.050 553.050 ;
        RECT 328.950 550.950 331.050 553.050 ;
        RECT 298.950 538.950 301.050 541.050 ;
        RECT 271.950 528.450 274.050 529.050 ;
        RECT 274.950 528.450 277.050 529.050 ;
        RECT 271.950 527.400 277.050 528.450 ;
        RECT 271.950 526.950 274.050 527.400 ;
        RECT 274.950 526.950 277.050 527.400 ;
        RECT 280.950 526.950 283.050 529.050 ;
        RECT 284.400 527.400 291.450 528.450 ;
        RECT 271.950 524.850 274.050 525.750 ;
        RECT 275.400 519.450 276.450 526.950 ;
        RECT 277.950 524.250 280.050 525.150 ;
        RECT 280.950 524.850 283.050 525.750 ;
        RECT 277.950 522.450 280.050 523.050 ;
        RECT 284.400 522.450 285.450 527.400 ;
        RECT 286.950 523.950 289.050 526.050 ;
        RECT 290.400 523.050 291.450 527.400 ;
        RECT 292.950 526.950 295.050 529.050 ;
        RECT 295.950 526.950 298.050 529.050 ;
        RECT 293.400 526.050 294.450 526.950 ;
        RECT 292.950 523.950 295.050 526.050 ;
        RECT 296.250 524.250 298.050 525.150 ;
        RECT 277.950 521.400 285.450 522.450 ;
        RECT 286.950 521.850 288.750 522.750 ;
        RECT 277.950 520.950 280.050 521.400 ;
        RECT 275.400 518.400 279.450 519.450 ;
        RECT 268.950 485.250 271.050 486.150 ;
        RECT 274.950 485.250 277.050 486.150 ;
        RECT 268.950 481.950 271.050 484.050 ;
        RECT 272.250 482.250 273.750 483.150 ;
        RECT 274.950 481.950 277.050 484.050 ;
        RECT 271.950 478.950 274.050 481.050 ;
        RECT 275.400 475.050 276.450 481.950 ;
        RECT 274.950 472.950 277.050 475.050 ;
        RECT 275.400 468.450 276.450 472.950 ;
        RECT 272.400 467.400 276.450 468.450 ;
        RECT 265.950 463.950 268.050 466.050 ;
        RECT 262.950 460.950 265.050 463.050 ;
        RECT 263.400 460.050 264.450 460.950 ;
        RECT 248.400 458.400 252.450 459.450 ;
        RECT 245.400 457.050 246.450 457.950 ;
        RECT 251.400 457.050 252.450 458.400 ;
        RECT 256.950 457.950 259.050 460.050 ;
        RECT 262.950 457.950 265.050 460.050 ;
        RECT 265.950 457.950 268.050 460.050 ;
        RECT 268.950 457.950 271.050 460.050 ;
        RECT 266.400 457.050 267.450 457.950 ;
        RECT 241.950 454.950 244.050 457.050 ;
        RECT 244.950 454.950 247.050 457.050 ;
        RECT 248.250 455.250 249.750 456.150 ;
        RECT 250.950 454.950 253.050 457.050 ;
        RECT 253.950 454.950 256.050 457.050 ;
        RECT 259.950 456.450 262.050 457.050 ;
        RECT 257.400 455.400 262.050 456.450 ;
        RECT 263.250 455.850 264.750 456.750 ;
        RECT 242.400 454.050 243.450 454.950 ;
        RECT 241.950 451.950 244.050 454.050 ;
        RECT 245.250 452.850 246.750 453.750 ;
        RECT 247.950 451.950 250.050 454.050 ;
        RECT 251.250 452.850 253.050 453.750 ;
        RECT 248.400 451.050 249.450 451.950 ;
        RECT 238.950 448.950 241.050 451.050 ;
        RECT 241.950 449.850 244.050 450.750 ;
        RECT 247.950 448.950 250.050 451.050 ;
        RECT 248.400 439.050 249.450 448.950 ;
        RECT 247.950 436.950 250.050 439.050 ;
        RECT 250.950 433.950 253.050 436.050 ;
        RECT 229.950 430.950 232.050 433.050 ;
        RECT 235.950 430.950 238.050 433.050 ;
        RECT 217.950 427.950 220.050 430.050 ;
        RECT 247.950 427.950 250.050 430.050 ;
        RECT 202.800 425.100 204.900 427.200 ;
        RECT 203.550 421.350 204.750 425.100 ;
        RECT 226.950 424.950 229.050 427.050 ;
        RECT 229.950 424.950 232.050 427.050 ;
        RECT 232.950 424.950 235.050 427.050 ;
        RECT 205.950 422.850 208.050 424.950 ;
        RECT 202.950 419.250 205.050 421.350 ;
        RECT 199.950 415.950 202.050 418.050 ;
        RECT 200.400 400.050 201.450 415.950 ;
        RECT 203.550 405.600 204.750 419.250 ;
        RECT 206.250 405.600 207.450 422.850 ;
        RECT 213.900 422.400 216.000 424.500 ;
        RECT 217.950 422.400 220.050 424.500 ;
        RECT 208.950 419.250 211.050 421.350 ;
        RECT 209.400 405.600 210.600 419.250 ;
        RECT 214.350 413.550 215.550 422.400 ;
        RECT 218.550 416.250 219.750 422.400 ;
        RECT 217.950 414.150 220.050 416.250 ;
        RECT 213.750 411.450 215.850 413.550 ;
        RECT 214.350 405.600 215.550 411.450 ;
        RECT 218.550 405.600 219.750 414.150 ;
        RECT 220.950 410.250 223.050 411.150 ;
        RECT 220.950 406.950 223.050 409.050 ;
        RECT 227.250 406.050 228.450 424.950 ;
        RECT 230.250 420.750 231.450 424.950 ;
        RECT 229.950 418.650 232.050 420.750 ;
        RECT 230.250 406.050 231.450 418.650 ;
        RECT 233.250 406.050 234.450 424.950 ;
        RECT 244.950 418.950 247.050 421.050 ;
        RECT 245.400 418.050 246.450 418.950 ;
        RECT 238.950 416.250 241.050 417.150 ;
        RECT 244.950 415.950 247.050 418.050 ;
        RECT 244.950 413.850 247.050 414.750 ;
        RECT 248.400 412.050 249.450 427.950 ;
        RECT 247.950 409.950 250.050 412.050 ;
        RECT 202.950 403.500 205.050 405.600 ;
        RECT 205.950 403.500 208.050 405.600 ;
        RECT 208.950 403.500 211.050 405.600 ;
        RECT 213.750 403.500 215.850 405.600 ;
        RECT 217.950 403.500 220.050 405.600 ;
        RECT 226.950 403.950 229.050 406.050 ;
        RECT 229.950 403.950 232.050 406.050 ;
        RECT 232.950 403.950 235.050 406.050 ;
        RECT 244.950 400.950 247.050 403.050 ;
        RECT 199.950 397.950 202.050 400.050 ;
        RECT 205.950 397.950 208.050 400.050 ;
        RECT 214.950 397.950 217.050 400.050 ;
        RECT 196.950 391.950 199.050 394.050 ;
        RECT 193.950 388.950 196.050 391.050 ;
        RECT 196.950 388.950 199.050 391.050 ;
        RECT 202.950 388.950 205.050 391.050 ;
        RECT 194.400 388.050 195.450 388.950 ;
        RECT 193.950 385.950 196.050 388.050 ;
        RECT 184.950 380.250 186.750 381.150 ;
        RECT 187.950 379.950 190.050 382.050 ;
        RECT 191.250 380.250 193.050 381.150 ;
        RECT 184.950 376.950 187.050 379.050 ;
        RECT 188.250 377.850 189.750 378.750 ;
        RECT 190.950 376.950 193.050 379.050 ;
        RECT 185.400 376.050 186.450 376.950 ;
        RECT 184.950 373.950 187.050 376.050 ;
        RECT 187.950 370.950 190.050 373.050 ;
        RECT 178.950 343.950 181.050 346.050 ;
        RECT 175.950 341.250 177.750 342.150 ;
        RECT 178.950 340.950 181.050 343.050 ;
        RECT 184.950 340.950 187.050 343.050 ;
        RECT 175.950 337.950 178.050 340.050 ;
        RECT 179.250 338.850 181.050 339.750 ;
        RECT 181.950 338.250 184.050 339.150 ;
        RECT 184.950 338.850 187.050 339.750 ;
        RECT 176.400 334.050 177.450 337.950 ;
        RECT 178.950 334.950 181.050 337.050 ;
        RECT 181.950 334.950 184.050 337.050 ;
        RECT 175.950 331.950 178.050 334.050 ;
        RECT 179.400 330.450 180.450 334.950 ;
        RECT 176.400 329.400 180.450 330.450 ;
        RECT 166.950 316.950 169.050 319.050 ;
        RECT 172.950 316.950 175.050 319.050 ;
        RECT 163.950 313.950 166.050 316.050 ;
        RECT 163.950 310.950 166.050 313.050 ;
        RECT 148.950 308.250 150.750 309.150 ;
        RECT 151.950 307.950 154.050 310.050 ;
        RECT 157.950 307.950 160.050 310.050 ;
        RECT 160.950 307.950 163.050 310.050 ;
        RECT 148.950 304.950 151.050 307.050 ;
        RECT 152.250 305.850 153.750 306.750 ;
        RECT 154.950 304.950 157.050 307.050 ;
        RECT 158.250 305.850 160.050 306.750 ;
        RECT 160.950 304.950 163.050 307.050 ;
        RECT 149.400 304.050 150.450 304.950 ;
        RECT 139.950 301.950 142.050 304.050 ;
        RECT 145.950 301.950 148.050 304.050 ;
        RECT 148.950 301.950 151.050 304.050 ;
        RECT 154.950 302.850 157.050 303.750 ;
        RECT 133.950 298.950 136.050 301.050 ;
        RECT 161.400 298.050 162.450 304.950 ;
        RECT 164.400 304.050 165.450 310.950 ;
        RECT 163.950 301.950 166.050 304.050 ;
        RECT 160.950 295.950 163.050 298.050 ;
        RECT 139.950 292.950 142.050 295.050 ;
        RECT 163.950 292.950 166.050 295.050 ;
        RECT 130.950 274.950 133.050 277.050 ;
        RECT 109.950 267.450 112.050 268.050 ;
        RECT 107.400 266.400 112.050 267.450 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 97.950 253.950 100.050 256.050 ;
        RECT 100.950 253.950 103.050 256.050 ;
        RECT 94.950 244.950 97.050 247.050 ;
        RECT 94.950 243.450 97.050 244.050 ;
        RECT 92.400 242.400 97.050 243.450 ;
        RECT 94.950 241.950 97.050 242.400 ;
        RECT 101.400 241.050 102.450 253.950 ;
        RECT 103.950 250.950 106.050 253.050 ;
        RECT 91.950 239.250 94.050 240.150 ;
        RECT 94.950 239.850 97.050 240.750 ;
        RECT 97.950 239.250 99.750 240.150 ;
        RECT 100.950 238.950 103.050 241.050 ;
        RECT 91.950 235.950 94.050 238.050 ;
        RECT 94.950 235.950 97.050 238.050 ;
        RECT 97.950 235.950 100.050 238.050 ;
        RECT 101.250 236.850 103.050 237.750 ;
        RECT 88.950 220.950 91.050 223.050 ;
        RECT 92.400 220.050 93.450 235.950 ;
        RECT 91.950 217.950 94.050 220.050 ;
        RECT 95.400 217.050 96.450 235.950 ;
        RECT 94.950 214.950 97.050 217.050 ;
        RECT 85.950 211.950 88.050 214.050 ;
        RECT 94.950 211.950 97.050 214.050 ;
        RECT 82.950 202.950 85.050 205.050 ;
        RECT 88.950 202.950 91.050 205.050 ;
        RECT 89.400 202.050 90.450 202.950 ;
        RECT 82.950 201.450 85.050 202.050 ;
        RECT 80.400 200.400 85.050 201.450 ;
        RECT 76.950 193.950 79.050 196.050 ;
        RECT 67.950 190.950 70.050 193.050 ;
        RECT 73.950 190.950 76.050 193.050 ;
        RECT 70.950 184.950 73.050 187.050 ;
        RECT 64.950 181.950 67.050 184.050 ;
        RECT 61.950 169.950 64.050 172.050 ;
        RECT 65.400 168.450 66.450 181.950 ;
        RECT 67.950 169.950 70.050 172.050 ;
        RECT 68.400 169.050 69.450 169.950 ;
        RECT 62.400 167.400 66.450 168.450 ;
        RECT 62.400 166.050 63.450 167.400 ;
        RECT 67.950 166.950 70.050 169.050 ;
        RECT 58.950 164.250 60.750 165.150 ;
        RECT 61.950 163.950 64.050 166.050 ;
        RECT 64.950 163.950 67.050 166.050 ;
        RECT 67.950 163.950 70.050 166.050 ;
        RECT 65.400 163.050 66.450 163.950 ;
        RECT 58.950 160.950 61.050 163.050 ;
        RECT 62.250 161.850 63.750 162.750 ;
        RECT 64.950 160.950 67.050 163.050 ;
        RECT 68.250 161.850 70.050 162.750 ;
        RECT 59.400 157.050 60.450 160.950 ;
        RECT 61.950 157.950 64.050 160.050 ;
        RECT 64.950 158.850 67.050 159.750 ;
        RECT 67.950 157.950 70.050 160.050 ;
        RECT 58.950 154.950 61.050 157.050 ;
        RECT 58.950 145.950 61.050 148.050 ;
        RECT 53.400 131.400 57.450 132.450 ;
        RECT 47.250 117.600 48.450 131.250 ;
        RECT 49.950 127.950 52.050 130.050 ;
        RECT 31.950 115.500 34.050 117.600 ;
        RECT 36.150 115.500 38.250 117.600 ;
        RECT 40.950 115.500 43.050 117.600 ;
        RECT 43.950 115.500 46.050 117.600 ;
        RECT 46.950 115.500 49.050 117.600 ;
        RECT 46.950 109.950 49.050 112.050 ;
        RECT 31.950 94.950 34.050 97.050 ;
        RECT 40.950 94.950 43.050 97.050 ;
        RECT 10.950 92.250 12.750 93.150 ;
        RECT 13.950 91.950 16.050 94.050 ;
        RECT 17.250 92.250 19.050 93.150 ;
        RECT 19.950 91.950 22.050 94.050 ;
        RECT 22.950 92.250 24.750 93.150 ;
        RECT 25.950 91.950 28.050 94.050 ;
        RECT 29.250 92.250 31.050 93.150 ;
        RECT 10.950 88.950 13.050 91.050 ;
        RECT 14.250 89.850 15.750 90.750 ;
        RECT 16.950 90.450 19.050 91.050 ;
        RECT 20.400 90.450 21.450 91.950 ;
        RECT 16.950 89.400 21.450 90.450 ;
        RECT 16.950 88.950 19.050 89.400 ;
        RECT 22.950 88.950 25.050 91.050 ;
        RECT 26.250 89.850 27.750 90.750 ;
        RECT 28.950 90.450 31.050 91.050 ;
        RECT 32.400 90.450 33.450 94.950 ;
        RECT 41.400 94.050 42.450 94.950 ;
        RECT 37.950 92.250 39.750 93.150 ;
        RECT 40.950 91.950 43.050 94.050 ;
        RECT 44.250 92.250 46.050 93.150 ;
        RECT 28.950 89.400 33.450 90.450 ;
        RECT 28.950 88.950 31.050 89.400 ;
        RECT 37.950 88.950 40.050 91.050 ;
        RECT 41.250 89.850 42.750 90.750 ;
        RECT 43.950 88.950 46.050 91.050 ;
        RECT 11.400 85.050 12.450 88.950 ;
        RECT 10.950 82.950 13.050 85.050 ;
        RECT 44.400 82.050 45.450 88.950 ;
        RECT 43.950 79.950 46.050 82.050 ;
        RECT 47.400 76.050 48.450 109.950 ;
        RECT 50.400 91.050 51.450 127.950 ;
        RECT 53.400 126.450 54.450 131.400 ;
        RECT 55.950 128.250 58.050 129.150 ;
        RECT 55.950 126.450 58.050 127.050 ;
        RECT 53.400 125.400 58.050 126.450 ;
        RECT 55.950 124.950 58.050 125.400 ;
        RECT 52.950 115.950 55.050 118.050 ;
        RECT 53.400 109.050 54.450 115.950 ;
        RECT 56.400 112.050 57.450 124.950 ;
        RECT 59.400 118.050 60.450 145.950 ;
        RECT 62.400 121.050 63.450 157.950 ;
        RECT 68.400 132.450 69.450 157.950 ;
        RECT 65.400 131.400 69.450 132.450 ;
        RECT 61.950 118.950 64.050 121.050 ;
        RECT 58.950 115.950 61.050 118.050 ;
        RECT 55.950 109.950 58.050 112.050 ;
        RECT 52.950 106.950 55.050 109.050 ;
        RECT 49.950 88.950 52.050 91.050 ;
        RECT 53.400 90.450 54.450 106.950 ;
        RECT 65.400 100.050 66.450 131.400 ;
        RECT 67.950 127.950 70.050 130.050 ;
        RECT 68.400 127.050 69.450 127.950 ;
        RECT 67.950 124.950 70.050 127.050 ;
        RECT 71.400 124.050 72.450 184.950 ;
        RECT 74.400 172.050 75.450 190.950 ;
        RECT 80.400 190.050 81.450 200.400 ;
        RECT 82.950 199.950 85.050 200.400 ;
        RECT 86.250 200.250 87.750 201.150 ;
        RECT 88.950 199.950 91.050 202.050 ;
        RECT 82.950 197.850 84.750 198.750 ;
        RECT 85.950 196.950 88.050 199.050 ;
        RECT 89.250 197.850 91.050 198.750 ;
        RECT 91.950 197.250 94.050 198.150 ;
        RECT 82.950 193.950 85.050 196.050 ;
        RECT 79.950 187.950 82.050 190.050 ;
        RECT 83.400 177.450 84.450 193.950 ;
        RECT 86.400 181.050 87.450 196.950 ;
        RECT 91.950 193.950 94.050 196.050 ;
        RECT 92.400 190.050 93.450 193.950 ;
        RECT 95.400 190.050 96.450 211.950 ;
        RECT 98.400 208.050 99.450 235.950 ;
        RECT 104.400 235.050 105.450 250.950 ;
        RECT 107.400 250.050 108.450 266.400 ;
        RECT 109.950 265.950 112.050 266.400 ;
        RECT 113.250 266.250 114.750 267.150 ;
        RECT 115.950 265.950 118.050 268.050 ;
        RECT 118.950 265.950 121.050 268.050 ;
        RECT 122.250 266.250 123.750 267.150 ;
        RECT 124.950 265.950 127.050 268.050 ;
        RECT 127.950 265.950 130.050 268.050 ;
        RECT 112.950 262.950 115.050 265.050 ;
        RECT 115.950 262.950 118.050 265.050 ;
        RECT 113.400 259.050 114.450 262.950 ;
        RECT 112.950 256.950 115.050 259.050 ;
        RECT 106.950 247.950 109.050 250.050 ;
        RECT 112.950 247.950 115.050 250.050 ;
        RECT 106.950 244.950 109.050 247.050 ;
        RECT 109.950 244.950 112.050 247.050 ;
        RECT 107.400 241.050 108.450 244.950 ;
        RECT 110.400 241.050 111.450 244.950 ;
        RECT 113.400 244.050 114.450 247.950 ;
        RECT 112.950 241.950 115.050 244.050 ;
        RECT 116.400 241.050 117.450 262.950 ;
        RECT 119.400 256.050 120.450 265.950 ;
        RECT 121.950 262.950 124.050 265.050 ;
        RECT 125.400 259.050 126.450 265.950 ;
        RECT 131.400 259.050 132.450 274.950 ;
        RECT 140.400 274.050 141.450 292.950 ;
        RECT 145.950 275.250 148.050 276.150 ;
        RECT 154.950 275.250 157.050 276.150 ;
        RECT 133.950 271.950 136.050 274.050 ;
        RECT 139.950 271.950 142.050 274.050 ;
        RECT 143.250 272.250 144.750 273.150 ;
        RECT 145.950 271.950 148.050 274.050 ;
        RECT 149.250 272.250 151.050 273.150 ;
        RECT 151.950 272.250 153.750 273.150 ;
        RECT 154.950 271.950 157.050 274.050 ;
        RECT 158.250 272.250 159.750 273.150 ;
        RECT 160.950 271.950 163.050 274.050 ;
        RECT 124.950 256.950 127.050 259.050 ;
        RECT 130.950 256.950 133.050 259.050 ;
        RECT 134.400 256.050 135.450 271.950 ;
        RECT 146.400 271.050 147.450 271.950 ;
        RECT 139.950 269.850 141.750 270.750 ;
        RECT 142.950 268.950 145.050 271.050 ;
        RECT 145.950 268.950 148.050 271.050 ;
        RECT 148.950 268.950 151.050 271.050 ;
        RECT 151.950 268.950 154.050 271.050 ;
        RECT 157.950 270.450 160.050 271.050 ;
        RECT 155.400 269.400 160.050 270.450 ;
        RECT 161.250 269.850 163.050 270.750 ;
        RECT 143.400 267.450 144.450 268.950 ;
        RECT 149.400 268.050 150.450 268.950 ;
        RECT 140.400 266.400 144.450 267.450 ;
        RECT 140.400 265.050 141.450 266.400 ;
        RECT 148.950 265.950 151.050 268.050 ;
        RECT 139.950 262.950 142.050 265.050 ;
        RECT 142.950 262.950 145.050 265.050 ;
        RECT 136.950 256.950 139.050 259.050 ;
        RECT 118.950 253.950 121.050 256.050 ;
        RECT 133.950 253.950 136.050 256.050 ;
        RECT 134.400 253.050 135.450 253.950 ;
        RECT 121.950 250.950 124.050 253.050 ;
        RECT 133.950 250.950 136.050 253.050 ;
        RECT 118.950 244.950 121.050 247.050 ;
        RECT 106.950 238.950 109.050 241.050 ;
        RECT 109.950 238.950 112.050 241.050 ;
        RECT 113.250 239.850 114.750 240.750 ;
        RECT 115.950 238.950 118.050 241.050 ;
        RECT 106.950 235.950 109.050 238.050 ;
        RECT 109.950 236.850 112.050 237.750 ;
        RECT 115.950 236.850 118.050 237.750 ;
        RECT 103.950 232.950 106.050 235.050 ;
        RECT 103.950 226.950 106.050 229.050 ;
        RECT 97.950 205.950 100.050 208.050 ;
        RECT 97.950 202.950 100.050 205.050 ;
        RECT 98.400 202.050 99.450 202.950 ;
        RECT 97.950 199.950 100.050 202.050 ;
        RECT 104.400 199.050 105.450 226.950 ;
        RECT 97.950 197.850 100.050 198.750 ;
        RECT 100.950 197.250 103.050 198.150 ;
        RECT 103.950 196.950 106.050 199.050 ;
        RECT 100.950 193.950 103.050 196.050 ;
        RECT 91.950 187.950 94.050 190.050 ;
        RECT 94.950 187.950 97.050 190.050 ;
        RECT 92.400 187.050 93.450 187.950 ;
        RECT 91.950 184.950 94.050 187.050 ;
        RECT 95.400 184.050 96.450 187.950 ;
        RECT 101.400 184.050 102.450 193.950 ;
        RECT 107.400 193.050 108.450 235.950 ;
        RECT 119.400 232.050 120.450 244.950 ;
        RECT 118.950 229.950 121.050 232.050 ;
        RECT 112.950 203.250 115.050 204.150 ;
        RECT 109.950 200.250 111.750 201.150 ;
        RECT 112.950 199.950 115.050 202.050 ;
        RECT 116.250 200.250 117.750 201.150 ;
        RECT 118.950 199.950 121.050 202.050 ;
        RECT 109.950 196.950 112.050 199.050 ;
        RECT 106.950 190.950 109.050 193.050 ;
        RECT 113.400 190.050 114.450 199.950 ;
        RECT 115.950 196.950 118.050 199.050 ;
        RECT 119.250 197.850 121.050 198.750 ;
        RECT 116.400 196.050 117.450 196.950 ;
        RECT 115.950 193.950 118.050 196.050 ;
        RECT 109.950 187.950 112.050 190.050 ;
        RECT 112.950 187.950 115.050 190.050 ;
        RECT 118.950 187.950 121.050 190.050 ;
        RECT 94.950 181.950 97.050 184.050 ;
        RECT 100.950 181.950 103.050 184.050 ;
        RECT 85.950 178.950 88.050 181.050 ;
        RECT 83.400 176.400 87.450 177.450 ;
        RECT 73.950 169.950 76.050 172.050 ;
        RECT 79.950 169.950 82.050 172.050 ;
        RECT 73.950 166.950 76.050 169.050 ;
        RECT 77.250 167.250 79.050 168.150 ;
        RECT 79.950 167.850 82.050 168.750 ;
        RECT 82.950 167.250 85.050 168.150 ;
        RECT 73.950 164.850 75.750 165.750 ;
        RECT 76.950 163.950 79.050 166.050 ;
        RECT 82.950 163.950 85.050 166.050 ;
        RECT 73.950 160.950 76.050 163.050 ;
        RECT 79.950 160.950 82.050 163.050 ;
        RECT 74.400 154.050 75.450 160.950 ;
        RECT 76.950 157.950 79.050 160.050 ;
        RECT 73.950 151.950 76.050 154.050 ;
        RECT 77.400 147.450 78.450 157.950 ;
        RECT 80.400 157.050 81.450 160.950 ;
        RECT 83.400 157.050 84.450 163.950 ;
        RECT 79.950 154.950 82.050 157.050 ;
        RECT 82.950 154.950 85.050 157.050 ;
        RECT 77.400 146.400 81.450 147.450 ;
        RECT 73.950 139.950 76.050 142.050 ;
        RECT 74.400 130.050 75.450 139.950 ;
        RECT 73.950 127.950 76.050 130.050 ;
        RECT 67.950 122.850 70.050 123.750 ;
        RECT 70.950 121.950 73.050 124.050 ;
        RECT 73.950 118.950 76.050 121.050 ;
        RECT 67.950 109.950 70.050 112.050 ;
        RECT 58.950 97.950 61.050 100.050 ;
        RECT 64.950 97.950 67.050 100.050 ;
        RECT 59.400 97.050 60.450 97.950 ;
        RECT 58.950 94.950 61.050 97.050 ;
        RECT 59.400 94.050 60.450 94.950 ;
        RECT 65.400 94.050 66.450 97.950 ;
        RECT 68.400 97.050 69.450 109.950 ;
        RECT 74.400 97.050 75.450 118.950 ;
        RECT 80.400 106.050 81.450 146.400 ;
        RECT 86.400 133.050 87.450 176.400 ;
        RECT 91.950 172.950 94.050 175.050 ;
        RECT 106.950 172.950 109.050 175.050 ;
        RECT 88.950 169.950 91.050 172.050 ;
        RECT 89.400 163.050 90.450 169.950 ;
        RECT 88.950 160.950 91.050 163.050 ;
        RECT 92.400 162.450 93.450 172.950 ;
        RECT 97.950 169.950 100.050 172.050 ;
        RECT 98.400 166.050 99.450 169.950 ;
        RECT 107.400 166.050 108.450 172.950 ;
        RECT 110.400 166.050 111.450 187.950 ;
        RECT 112.950 181.950 115.050 184.050 ;
        RECT 113.400 166.050 114.450 181.950 ;
        RECT 94.950 164.250 96.750 165.150 ;
        RECT 97.950 163.950 100.050 166.050 ;
        RECT 103.950 163.950 106.050 166.050 ;
        RECT 106.950 163.950 109.050 166.050 ;
        RECT 109.950 163.950 112.050 166.050 ;
        RECT 112.950 163.950 115.050 166.050 ;
        RECT 116.250 164.250 118.050 165.150 ;
        RECT 94.950 162.450 97.050 163.050 ;
        RECT 92.400 161.400 97.050 162.450 ;
        RECT 98.250 161.850 99.750 162.750 ;
        RECT 94.950 160.950 97.050 161.400 ;
        RECT 100.950 160.950 103.050 163.050 ;
        RECT 104.250 161.850 106.050 162.750 ;
        RECT 106.950 161.850 108.750 162.750 ;
        RECT 109.950 160.950 112.050 163.050 ;
        RECT 113.250 161.850 114.750 162.750 ;
        RECT 115.950 160.950 118.050 163.050 ;
        RECT 89.400 154.050 90.450 160.950 ;
        RECT 100.950 158.850 103.050 159.750 ;
        RECT 103.950 157.950 106.050 160.050 ;
        RECT 106.950 157.950 109.050 160.050 ;
        RECT 109.950 158.850 112.050 159.750 ;
        RECT 112.950 157.950 115.050 160.050 ;
        RECT 88.950 151.950 91.050 154.050 ;
        RECT 97.950 148.950 100.050 151.050 ;
        RECT 88.950 142.950 91.050 145.050 ;
        RECT 82.950 130.950 85.050 133.050 ;
        RECT 85.950 130.950 88.050 133.050 ;
        RECT 83.400 130.050 84.450 130.950 ;
        RECT 89.400 130.050 90.450 142.950 ;
        RECT 82.950 127.950 85.050 130.050 ;
        RECT 86.250 128.250 87.750 129.150 ;
        RECT 88.950 127.950 91.050 130.050 ;
        RECT 82.950 125.850 84.750 126.750 ;
        RECT 85.950 124.950 88.050 127.050 ;
        RECT 89.250 125.850 91.050 126.750 ;
        RECT 94.950 124.950 97.050 127.050 ;
        RECT 86.400 121.050 87.450 124.950 ;
        RECT 91.950 122.250 94.050 123.150 ;
        RECT 94.950 122.850 97.050 123.750 ;
        RECT 82.950 118.950 85.050 121.050 ;
        RECT 85.950 118.950 88.050 121.050 ;
        RECT 91.950 118.950 94.050 121.050 ;
        RECT 79.950 103.950 82.050 106.050 ;
        RECT 79.950 100.950 82.050 103.050 ;
        RECT 67.950 94.950 70.050 97.050 ;
        RECT 71.250 95.250 72.750 96.150 ;
        RECT 73.950 94.950 76.050 97.050 ;
        RECT 76.950 94.950 79.050 97.050 ;
        RECT 77.400 94.050 78.450 94.950 ;
        RECT 80.400 94.050 81.450 100.950 ;
        RECT 83.400 97.050 84.450 118.950 ;
        RECT 94.950 103.950 97.050 106.050 ;
        RECT 85.950 100.950 88.050 103.050 ;
        RECT 86.400 100.050 87.450 100.950 ;
        RECT 85.950 97.950 88.050 100.050 ;
        RECT 82.950 94.950 85.050 97.050 ;
        RECT 86.250 95.850 87.750 96.750 ;
        RECT 88.950 96.450 91.050 97.050 ;
        RECT 88.950 95.400 93.450 96.450 ;
        RECT 88.950 94.950 91.050 95.400 ;
        RECT 55.950 92.250 57.750 93.150 ;
        RECT 58.950 91.950 61.050 94.050 ;
        RECT 61.950 91.950 64.050 94.050 ;
        RECT 64.950 91.950 67.050 94.050 ;
        RECT 67.950 92.850 69.750 93.750 ;
        RECT 70.950 91.950 73.050 94.050 ;
        RECT 74.250 92.850 75.750 93.750 ;
        RECT 76.950 91.950 79.050 94.050 ;
        RECT 79.950 91.950 82.050 94.050 ;
        RECT 82.950 92.850 85.050 93.750 ;
        RECT 88.950 92.850 91.050 93.750 ;
        RECT 62.400 91.050 63.450 91.950 ;
        RECT 55.950 90.450 58.050 91.050 ;
        RECT 53.400 89.400 58.050 90.450 ;
        RECT 59.250 89.850 60.750 90.750 ;
        RECT 55.950 88.950 58.050 89.400 ;
        RECT 61.950 88.950 64.050 91.050 ;
        RECT 65.250 89.850 67.050 90.750 ;
        RECT 61.950 86.850 64.050 87.750 ;
        RECT 71.400 85.050 72.450 91.950 ;
        RECT 76.950 89.850 79.050 90.750 ;
        RECT 70.950 82.950 73.050 85.050 ;
        RECT 52.950 79.950 55.050 82.050 ;
        RECT 46.950 73.950 49.050 76.050 ;
        RECT 16.950 64.950 19.050 67.050 ;
        RECT 19.950 64.950 22.050 67.050 ;
        RECT 22.950 64.950 25.050 67.050 ;
        RECT 47.100 65.100 49.200 67.200 ;
        RECT 4.950 57.450 7.050 58.050 ;
        RECT 2.400 56.400 7.050 57.450 ;
        RECT 2.400 18.450 3.450 56.400 ;
        RECT 4.950 55.950 7.050 56.400 ;
        RECT 10.950 56.250 13.050 57.150 ;
        RECT 4.950 53.850 7.050 54.750 ;
        RECT 17.550 46.050 18.750 64.950 ;
        RECT 20.550 60.750 21.750 64.950 ;
        RECT 19.950 58.650 22.050 60.750 ;
        RECT 20.550 46.050 21.750 58.650 ;
        RECT 23.550 46.050 24.750 64.950 ;
        RECT 31.950 62.400 34.050 64.500 ;
        RECT 36.000 62.400 38.100 64.500 ;
        RECT 43.950 62.850 46.050 64.950 ;
        RECT 32.250 56.250 33.450 62.400 ;
        RECT 31.950 54.150 34.050 56.250 ;
        RECT 28.950 50.250 31.050 51.150 ;
        RECT 28.950 46.950 31.050 49.050 ;
        RECT 16.950 43.950 19.050 46.050 ;
        RECT 19.950 43.950 22.050 46.050 ;
        RECT 22.950 43.950 25.050 46.050 ;
        RECT 32.250 45.600 33.450 54.150 ;
        RECT 36.450 53.550 37.650 62.400 ;
        RECT 40.950 59.250 43.050 61.350 ;
        RECT 36.150 51.450 38.250 53.550 ;
        RECT 36.450 45.600 37.650 51.450 ;
        RECT 41.400 45.600 42.600 59.250 ;
        RECT 44.550 45.600 45.750 62.850 ;
        RECT 47.250 61.350 48.450 65.100 ;
        RECT 46.950 59.250 49.050 61.350 ;
        RECT 47.250 45.600 48.450 59.250 ;
        RECT 31.950 43.500 34.050 45.600 ;
        RECT 36.150 43.500 38.250 45.600 ;
        RECT 40.950 43.500 43.050 45.600 ;
        RECT 43.950 43.500 46.050 45.600 ;
        RECT 46.950 43.500 49.050 45.600 ;
        RECT 16.950 28.950 19.050 31.050 ;
        RECT 19.950 28.950 22.050 31.050 ;
        RECT 22.950 28.950 25.050 31.050 ;
        RECT 31.950 29.400 34.050 31.500 ;
        RECT 36.150 29.400 38.250 31.500 ;
        RECT 40.950 29.400 43.050 31.500 ;
        RECT 43.950 29.400 46.050 31.500 ;
        RECT 46.950 29.400 49.050 31.500 ;
        RECT 4.950 20.250 7.050 21.150 ;
        RECT 4.950 18.450 7.050 19.050 ;
        RECT 2.400 17.400 7.050 18.450 ;
        RECT 10.950 17.850 13.050 18.750 ;
        RECT 4.950 16.950 7.050 17.400 ;
        RECT 5.400 10.050 6.450 16.950 ;
        RECT 17.550 10.050 18.750 28.950 ;
        RECT 20.550 16.350 21.750 28.950 ;
        RECT 19.950 14.250 22.050 16.350 ;
        RECT 20.550 10.050 21.750 14.250 ;
        RECT 23.550 10.050 24.750 28.950 ;
        RECT 28.950 25.950 31.050 28.050 ;
        RECT 28.950 23.850 31.050 24.750 ;
        RECT 32.250 20.850 33.450 29.400 ;
        RECT 36.450 23.550 37.650 29.400 ;
        RECT 36.150 21.450 38.250 23.550 ;
        RECT 31.950 18.750 34.050 20.850 ;
        RECT 32.250 12.600 33.450 18.750 ;
        RECT 36.450 12.600 37.650 21.450 ;
        RECT 41.400 15.750 42.600 29.400 ;
        RECT 40.950 13.650 43.050 15.750 ;
        RECT 31.950 10.500 34.050 12.600 ;
        RECT 36.000 10.500 38.100 12.600 ;
        RECT 44.550 12.150 45.750 29.400 ;
        RECT 47.250 15.750 48.450 29.400 ;
        RECT 53.400 16.050 54.450 79.950 ;
        RECT 58.950 73.950 61.050 76.050 ;
        RECT 55.950 56.250 58.050 57.150 ;
        RECT 55.950 54.450 58.050 55.050 ;
        RECT 59.400 54.450 60.450 73.950 ;
        RECT 71.400 61.050 72.450 82.950 ;
        RECT 70.950 58.950 73.050 61.050 ;
        RECT 85.950 58.950 88.050 61.050 ;
        RECT 67.950 55.950 70.050 58.050 ;
        RECT 79.950 56.250 82.050 57.150 ;
        RECT 68.400 55.050 69.450 55.950 ;
        RECT 86.400 55.050 87.450 58.950 ;
        RECT 55.950 53.400 60.450 54.450 ;
        RECT 55.950 52.950 58.050 53.400 ;
        RECT 67.950 52.950 70.050 55.050 ;
        RECT 76.950 52.950 79.050 55.050 ;
        RECT 79.950 52.950 82.050 55.050 ;
        RECT 83.250 53.250 84.750 54.150 ;
        RECT 85.950 52.950 88.050 55.050 ;
        RECT 89.250 53.250 91.050 54.150 ;
        RECT 56.400 22.050 57.450 52.950 ;
        RECT 67.950 50.850 70.050 51.750 ;
        RECT 77.400 25.050 78.450 52.950 ;
        RECT 80.400 52.050 81.450 52.950 ;
        RECT 79.950 49.950 82.050 52.050 ;
        RECT 82.950 49.950 85.050 52.050 ;
        RECT 86.250 50.850 87.750 51.750 ;
        RECT 88.950 49.950 91.050 52.050 ;
        RECT 83.400 49.050 84.450 49.950 ;
        RECT 89.400 49.050 90.450 49.950 ;
        RECT 82.950 46.950 85.050 49.050 ;
        RECT 88.950 46.950 91.050 49.050 ;
        RECT 92.400 37.050 93.450 95.400 ;
        RECT 91.950 34.950 94.050 37.050 ;
        RECT 85.950 31.950 88.050 34.050 ;
        RECT 67.950 23.250 70.050 24.150 ;
        RECT 73.950 23.250 75.750 24.150 ;
        RECT 76.950 22.950 79.050 25.050 ;
        RECT 55.950 19.950 58.050 22.050 ;
        RECT 67.950 19.950 70.050 22.050 ;
        RECT 73.950 19.950 76.050 22.050 ;
        RECT 77.250 20.850 79.050 21.750 ;
        RECT 68.400 19.050 69.450 19.950 ;
        RECT 55.950 17.850 58.050 18.750 ;
        RECT 67.950 16.950 70.050 19.050 ;
        RECT 74.400 16.050 75.450 19.950 ;
        RECT 86.400 19.050 87.450 31.950 ;
        RECT 95.400 31.050 96.450 103.950 ;
        RECT 98.400 67.050 99.450 148.950 ;
        RECT 104.400 127.050 105.450 157.950 ;
        RECT 107.400 136.050 108.450 157.950 ;
        RECT 109.950 145.950 112.050 148.050 ;
        RECT 106.950 133.950 109.050 136.050 ;
        RECT 100.950 125.250 103.050 126.150 ;
        RECT 103.950 124.950 106.050 127.050 ;
        RECT 106.950 125.250 109.050 126.150 ;
        RECT 100.950 121.950 103.050 124.050 ;
        RECT 104.250 122.250 105.750 123.150 ;
        RECT 106.950 121.950 109.050 124.050 ;
        RECT 103.950 118.950 106.050 121.050 ;
        RECT 104.400 99.450 105.450 118.950 ;
        RECT 110.400 118.050 111.450 145.950 ;
        RECT 113.400 142.050 114.450 157.950 ;
        RECT 116.400 148.050 117.450 160.950 ;
        RECT 115.950 145.950 118.050 148.050 ;
        RECT 119.400 145.050 120.450 187.950 ;
        RECT 122.400 184.050 123.450 250.950 ;
        RECT 133.950 244.950 136.050 247.050 ;
        RECT 134.400 241.050 135.450 244.950 ;
        RECT 127.950 240.450 130.050 241.050 ;
        RECT 125.400 239.400 130.050 240.450 ;
        RECT 125.400 238.050 126.450 239.400 ;
        RECT 127.950 238.950 130.050 239.400 ;
        RECT 131.250 239.250 132.750 240.150 ;
        RECT 133.950 238.950 136.050 241.050 ;
        RECT 137.400 240.450 138.450 256.950 ;
        RECT 139.950 244.950 142.050 247.050 ;
        RECT 140.400 244.050 141.450 244.950 ;
        RECT 139.950 241.950 142.050 244.050 ;
        RECT 137.400 239.400 141.450 240.450 ;
        RECT 124.950 235.950 127.050 238.050 ;
        RECT 127.950 236.850 129.750 237.750 ;
        RECT 130.950 235.950 133.050 238.050 ;
        RECT 134.250 236.850 135.750 237.750 ;
        RECT 136.950 235.950 139.050 238.050 ;
        RECT 131.400 235.050 132.450 235.950 ;
        RECT 124.950 232.950 127.050 235.050 ;
        RECT 130.950 232.950 133.050 235.050 ;
        RECT 136.950 233.850 139.050 234.750 ;
        RECT 125.400 226.050 126.450 232.950 ;
        RECT 136.950 226.950 139.050 229.050 ;
        RECT 124.950 223.950 127.050 226.050 ;
        RECT 121.950 181.950 124.050 184.050 ;
        RECT 125.400 180.450 126.450 223.950 ;
        RECT 137.400 205.050 138.450 226.950 ;
        RECT 140.400 226.050 141.450 239.400 ;
        RECT 139.950 223.950 142.050 226.050 ;
        RECT 127.950 202.950 130.050 205.050 ;
        RECT 136.950 202.950 139.050 205.050 ;
        RECT 128.400 202.050 129.450 202.950 ;
        RECT 127.950 199.950 130.050 202.050 ;
        RECT 131.250 200.250 132.750 201.150 ;
        RECT 133.950 199.950 136.050 202.050 ;
        RECT 139.950 199.950 142.050 202.050 ;
        RECT 127.950 197.850 129.750 198.750 ;
        RECT 130.950 196.950 133.050 199.050 ;
        RECT 134.250 197.850 136.050 198.750 ;
        RECT 140.400 196.050 141.450 199.950 ;
        RECT 139.950 193.950 142.050 196.050 ;
        RECT 143.400 193.050 144.450 262.950 ;
        RECT 152.400 262.050 153.450 268.950 ;
        RECT 155.400 262.050 156.450 269.400 ;
        RECT 157.950 268.950 160.050 269.400 ;
        RECT 164.400 268.050 165.450 292.950 ;
        RECT 167.400 280.050 168.450 316.950 ;
        RECT 176.400 315.450 177.450 329.400 ;
        RECT 182.400 325.050 183.450 334.950 ;
        RECT 188.400 327.450 189.450 370.950 ;
        RECT 194.400 345.450 195.450 385.950 ;
        RECT 197.400 364.050 198.450 388.950 ;
        RECT 203.400 385.050 204.450 388.950 ;
        RECT 202.950 382.950 205.050 385.050 ;
        RECT 202.950 380.850 205.050 381.750 ;
        RECT 202.950 376.950 205.050 379.050 ;
        RECT 203.400 364.050 204.450 376.950 ;
        RECT 196.950 361.950 199.050 364.050 ;
        RECT 202.950 361.950 205.050 364.050 ;
        RECT 196.950 355.950 199.050 358.050 ;
        RECT 191.400 344.400 195.450 345.450 ;
        RECT 191.400 339.450 192.450 344.400 ;
        RECT 197.400 343.050 198.450 355.950 ;
        RECT 202.950 344.250 205.050 345.150 ;
        RECT 193.950 341.250 195.750 342.150 ;
        RECT 196.950 340.950 199.050 343.050 ;
        RECT 200.250 341.250 201.750 342.150 ;
        RECT 202.950 340.950 205.050 343.050 ;
        RECT 193.950 339.450 196.050 340.050 ;
        RECT 191.400 338.400 196.050 339.450 ;
        RECT 197.250 338.850 198.750 339.750 ;
        RECT 193.950 337.950 196.050 338.400 ;
        RECT 199.950 337.950 202.050 340.050 ;
        RECT 190.950 334.950 193.050 337.050 ;
        RECT 193.950 334.950 196.050 337.050 ;
        RECT 191.400 331.050 192.450 334.950 ;
        RECT 190.950 328.950 193.050 331.050 ;
        RECT 185.400 326.400 189.450 327.450 ;
        RECT 181.950 322.950 184.050 325.050 ;
        RECT 185.400 316.050 186.450 326.400 ;
        RECT 173.400 314.400 177.450 315.450 ;
        RECT 173.400 313.050 174.450 314.400 ;
        RECT 178.950 313.950 181.050 316.050 ;
        RECT 184.950 315.450 187.050 316.050 ;
        RECT 182.400 314.400 187.050 315.450 ;
        RECT 179.400 313.050 180.450 313.950 ;
        RECT 169.950 310.950 172.050 313.050 ;
        RECT 172.950 310.950 175.050 313.050 ;
        RECT 176.250 311.250 177.750 312.150 ;
        RECT 178.950 310.950 181.050 313.050 ;
        RECT 170.400 310.050 171.450 310.950 ;
        RECT 169.950 307.950 172.050 310.050 ;
        RECT 173.250 308.850 174.750 309.750 ;
        RECT 175.950 307.950 178.050 310.050 ;
        RECT 179.250 308.850 181.050 309.750 ;
        RECT 169.950 305.850 172.050 306.750 ;
        RECT 172.950 298.950 175.050 301.050 ;
        RECT 169.950 286.950 172.050 289.050 ;
        RECT 166.950 277.950 169.050 280.050 ;
        RECT 166.950 274.950 169.050 277.050 ;
        RECT 157.950 265.950 160.050 268.050 ;
        RECT 163.950 265.950 166.050 268.050 ;
        RECT 151.950 259.950 154.050 262.050 ;
        RECT 154.950 259.950 157.050 262.050 ;
        RECT 151.950 250.950 154.050 253.050 ;
        RECT 148.950 244.950 151.050 247.050 ;
        RECT 149.400 244.050 150.450 244.950 ;
        RECT 145.950 241.950 148.050 244.050 ;
        RECT 148.950 241.950 151.050 244.050 ;
        RECT 146.400 241.050 147.450 241.950 ;
        RECT 152.400 241.050 153.450 250.950 ;
        RECT 154.950 244.950 157.050 247.050 ;
        RECT 145.950 238.950 148.050 241.050 ;
        RECT 149.250 239.850 150.750 240.750 ;
        RECT 151.950 238.950 154.050 241.050 ;
        RECT 145.950 236.850 148.050 237.750 ;
        RECT 148.950 235.950 151.050 238.050 ;
        RECT 151.950 236.850 154.050 237.750 ;
        RECT 149.400 223.050 150.450 235.950 ;
        RECT 148.950 220.950 151.050 223.050 ;
        RECT 155.400 201.450 156.450 244.950 ;
        RECT 158.400 232.050 159.450 265.950 ;
        RECT 167.400 253.050 168.450 274.950 ;
        RECT 170.400 259.050 171.450 286.950 ;
        RECT 169.950 256.950 172.050 259.050 ;
        RECT 166.950 250.950 169.050 253.050 ;
        RECT 160.950 247.950 163.050 250.050 ;
        RECT 163.950 247.950 166.050 250.050 ;
        RECT 161.400 240.450 162.450 247.950 ;
        RECT 164.400 244.050 165.450 247.950 ;
        RECT 169.950 244.950 172.050 247.050 ;
        RECT 163.950 241.950 166.050 244.050 ;
        RECT 166.950 241.950 169.050 244.050 ;
        RECT 170.400 241.050 171.450 244.950 ;
        RECT 163.950 240.450 166.050 241.050 ;
        RECT 161.400 239.400 166.050 240.450 ;
        RECT 167.250 239.850 168.750 240.750 ;
        RECT 163.950 238.950 166.050 239.400 ;
        RECT 169.950 238.950 172.050 241.050 ;
        RECT 163.950 236.850 166.050 237.750 ;
        RECT 169.950 236.850 172.050 237.750 ;
        RECT 160.950 232.950 163.050 235.050 ;
        RECT 157.950 229.950 160.050 232.050 ;
        RECT 145.950 200.250 148.050 201.150 ;
        RECT 155.400 200.400 159.450 201.450 ;
        RECT 145.950 196.950 148.050 199.050 ;
        RECT 149.250 197.250 150.750 198.150 ;
        RECT 151.950 196.950 154.050 199.050 ;
        RECT 155.250 197.250 157.050 198.150 ;
        RECT 146.400 196.050 147.450 196.950 ;
        RECT 145.950 193.950 148.050 196.050 ;
        RECT 148.950 193.950 151.050 196.050 ;
        RECT 152.250 194.850 153.750 195.750 ;
        RECT 154.950 195.450 157.050 196.050 ;
        RECT 158.400 195.450 159.450 200.400 ;
        RECT 161.400 199.050 162.450 232.950 ;
        RECT 173.400 228.450 174.450 298.950 ;
        RECT 176.400 295.050 177.450 307.950 ;
        RECT 175.950 292.950 178.050 295.050 ;
        RECT 182.400 292.050 183.450 314.400 ;
        RECT 184.950 313.950 187.050 314.400 ;
        RECT 184.950 311.850 187.050 312.750 ;
        RECT 187.950 311.250 190.050 312.150 ;
        RECT 187.950 307.950 190.050 310.050 ;
        RECT 188.400 304.050 189.450 307.950 ;
        RECT 187.950 301.950 190.050 304.050 ;
        RECT 191.400 301.050 192.450 328.950 ;
        RECT 194.400 322.050 195.450 334.950 ;
        RECT 203.400 331.050 204.450 340.950 ;
        RECT 202.950 328.950 205.050 331.050 ;
        RECT 193.950 319.950 196.050 322.050 ;
        RECT 193.950 316.950 196.050 319.050 ;
        RECT 190.950 298.950 193.050 301.050 ;
        RECT 181.950 289.950 184.050 292.050 ;
        RECT 194.400 289.050 195.450 316.950 ;
        RECT 206.400 316.050 207.450 397.950 ;
        RECT 211.950 382.950 214.050 385.050 ;
        RECT 208.950 380.250 211.050 381.150 ;
        RECT 211.950 380.850 214.050 381.750 ;
        RECT 208.950 376.950 211.050 379.050 ;
        RECT 215.400 378.450 216.450 397.950 ;
        RECT 226.950 388.950 229.050 391.050 ;
        RECT 232.950 388.950 235.050 391.050 ;
        RECT 238.950 388.950 241.050 391.050 ;
        RECT 217.950 380.250 219.750 381.150 ;
        RECT 220.950 379.950 223.050 382.050 ;
        RECT 224.250 380.250 226.050 381.150 ;
        RECT 217.950 378.450 220.050 379.050 ;
        RECT 215.400 377.400 220.050 378.450 ;
        RECT 221.250 377.850 222.750 378.750 ;
        RECT 217.950 376.950 220.050 377.400 ;
        RECT 223.950 376.950 226.050 379.050 ;
        RECT 220.950 358.950 223.050 361.050 ;
        RECT 208.950 349.950 211.050 352.050 ;
        RECT 209.400 337.050 210.450 349.950 ;
        RECT 211.950 341.250 214.050 342.150 ;
        RECT 217.950 341.250 220.050 342.150 ;
        RECT 211.950 337.950 214.050 340.050 ;
        RECT 215.250 338.250 216.750 339.150 ;
        RECT 217.950 337.950 220.050 340.050 ;
        RECT 208.950 334.950 211.050 337.050 ;
        RECT 214.950 334.950 217.050 337.050 ;
        RECT 218.400 334.050 219.450 337.950 ;
        RECT 221.400 337.050 222.450 358.950 ;
        RECT 224.400 340.050 225.450 376.950 ;
        RECT 227.400 361.050 228.450 388.950 ;
        RECT 233.400 388.050 234.450 388.950 ;
        RECT 232.950 385.950 235.050 388.050 ;
        RECT 239.400 385.050 240.450 388.950 ;
        RECT 229.950 383.250 232.050 384.150 ;
        RECT 232.950 383.850 235.050 384.750 ;
        RECT 235.950 383.250 237.750 384.150 ;
        RECT 238.950 382.950 241.050 385.050 ;
        RECT 229.950 379.950 232.050 382.050 ;
        RECT 235.950 379.950 238.050 382.050 ;
        RECT 239.250 380.850 241.050 381.750 ;
        RECT 238.950 376.950 241.050 379.050 ;
        RECT 226.950 358.950 229.050 361.050 ;
        RECT 235.950 344.250 238.050 345.150 ;
        RECT 226.950 341.250 228.750 342.150 ;
        RECT 229.950 340.950 232.050 343.050 ;
        RECT 233.250 341.250 234.750 342.150 ;
        RECT 235.950 340.950 238.050 343.050 ;
        RECT 223.950 337.950 226.050 340.050 ;
        RECT 226.950 337.950 229.050 340.050 ;
        RECT 230.250 338.850 231.750 339.750 ;
        RECT 232.950 337.950 235.050 340.050 ;
        RECT 220.950 334.950 223.050 337.050 ;
        RECT 227.400 334.050 228.450 337.950 ;
        RECT 233.400 337.050 234.450 337.950 ;
        RECT 232.950 334.950 235.050 337.050 ;
        RECT 217.950 331.950 220.050 334.050 ;
        RECT 226.950 331.950 229.050 334.050 ;
        RECT 236.400 322.050 237.450 340.950 ;
        RECT 239.400 337.050 240.450 376.950 ;
        RECT 245.400 370.050 246.450 400.950 ;
        RECT 251.400 396.450 252.450 433.950 ;
        RECT 254.400 424.050 255.450 454.950 ;
        RECT 257.400 445.050 258.450 455.400 ;
        RECT 259.950 454.950 262.050 455.400 ;
        RECT 265.950 454.950 268.050 457.050 ;
        RECT 259.950 452.850 262.050 453.750 ;
        RECT 265.950 452.850 268.050 453.750 ;
        RECT 256.950 442.950 259.050 445.050 ;
        RECT 256.950 436.950 259.050 439.050 ;
        RECT 253.950 421.950 256.050 424.050 ;
        RECT 257.400 415.050 258.450 436.950 ;
        RECT 262.950 416.250 265.050 417.150 ;
        RECT 253.950 413.250 255.750 414.150 ;
        RECT 256.950 412.950 259.050 415.050 ;
        RECT 260.250 413.250 261.750 414.150 ;
        RECT 262.950 412.950 265.050 415.050 ;
        RECT 265.950 412.950 268.050 415.050 ;
        RECT 253.950 409.950 256.050 412.050 ;
        RECT 257.250 410.850 258.750 411.750 ;
        RECT 259.950 409.950 262.050 412.050 ;
        RECT 260.400 403.050 261.450 409.950 ;
        RECT 263.400 409.050 264.450 412.950 ;
        RECT 262.950 406.950 265.050 409.050 ;
        RECT 262.950 403.950 265.050 406.050 ;
        RECT 259.950 400.950 262.050 403.050 ;
        RECT 248.400 395.400 252.450 396.450 ;
        RECT 248.400 382.050 249.450 395.400 ;
        RECT 250.950 391.950 253.050 394.050 ;
        RECT 251.400 385.050 252.450 391.950 ;
        RECT 250.950 382.950 253.050 385.050 ;
        RECT 254.250 383.250 255.750 384.150 ;
        RECT 256.950 382.950 259.050 385.050 ;
        RECT 247.950 379.950 250.050 382.050 ;
        RECT 251.250 380.850 252.750 381.750 ;
        RECT 253.950 379.950 256.050 382.050 ;
        RECT 257.250 380.850 259.050 381.750 ;
        RECT 254.400 379.050 255.450 379.950 ;
        RECT 247.950 377.850 250.050 378.750 ;
        RECT 253.950 376.950 256.050 379.050 ;
        RECT 244.950 367.950 247.050 370.050 ;
        RECT 259.950 367.950 262.050 370.050 ;
        RECT 244.950 342.450 247.050 343.050 ;
        RECT 242.400 341.400 247.050 342.450 ;
        RECT 238.950 334.950 241.050 337.050 ;
        RECT 242.400 331.050 243.450 341.400 ;
        RECT 244.950 340.950 247.050 341.400 ;
        RECT 250.950 340.950 253.050 343.050 ;
        RECT 254.250 341.250 256.050 342.150 ;
        RECT 256.950 340.950 259.050 343.050 ;
        RECT 244.950 338.850 247.050 339.750 ;
        RECT 247.950 338.250 250.050 339.150 ;
        RECT 250.950 338.850 252.750 339.750 ;
        RECT 253.950 337.950 256.050 340.050 ;
        RECT 254.400 337.050 255.450 337.950 ;
        RECT 247.950 334.950 250.050 337.050 ;
        RECT 253.950 334.950 256.050 337.050 ;
        RECT 241.950 328.950 244.050 331.050 ;
        RECT 248.400 328.050 249.450 334.950 ;
        RECT 257.400 328.050 258.450 340.950 ;
        RECT 247.950 325.950 250.050 328.050 ;
        RECT 256.950 325.950 259.050 328.050 ;
        RECT 223.950 319.950 226.050 322.050 ;
        RECT 235.950 319.950 238.050 322.050 ;
        RECT 260.400 321.450 261.450 367.950 ;
        RECT 263.400 337.050 264.450 403.950 ;
        RECT 266.400 403.050 267.450 412.950 ;
        RECT 265.950 400.950 268.050 403.050 ;
        RECT 265.950 394.950 268.050 397.050 ;
        RECT 266.400 384.450 267.450 394.950 ;
        RECT 269.400 388.050 270.450 457.950 ;
        RECT 272.400 457.050 273.450 467.400 ;
        RECT 274.950 463.950 277.050 466.050 ;
        RECT 271.950 454.950 274.050 457.050 ;
        RECT 271.950 452.850 274.050 453.750 ;
        RECT 271.950 442.950 274.050 445.050 ;
        RECT 272.400 406.050 273.450 442.950 ;
        RECT 275.400 421.050 276.450 463.950 ;
        RECT 278.400 463.050 279.450 518.400 ;
        RECT 281.400 481.050 282.450 521.400 ;
        RECT 289.950 520.950 292.050 523.050 ;
        RECT 293.250 521.850 294.750 522.750 ;
        RECT 295.950 522.450 298.050 523.050 ;
        RECT 299.400 522.450 300.450 538.950 ;
        RECT 304.950 535.950 307.050 538.050 ;
        RECT 301.950 523.950 304.050 526.050 ;
        RECT 295.950 521.400 300.450 522.450 ;
        RECT 295.950 520.950 298.050 521.400 ;
        RECT 302.400 520.050 303.450 523.950 ;
        RECT 283.950 517.950 286.050 520.050 ;
        RECT 289.950 518.850 292.050 519.750 ;
        RECT 301.950 517.950 304.050 520.050 ;
        RECT 280.950 478.950 283.050 481.050 ;
        RECT 277.950 460.950 280.050 463.050 ;
        RECT 280.950 460.950 283.050 463.050 ;
        RECT 281.400 457.050 282.450 460.950 ;
        RECT 280.950 454.950 283.050 457.050 ;
        RECT 277.950 452.250 280.050 453.150 ;
        RECT 280.950 452.850 283.050 453.750 ;
        RECT 277.950 448.950 280.050 451.050 ;
        RECT 274.950 418.950 277.050 421.050 ;
        RECT 278.400 418.050 279.450 448.950 ;
        RECT 280.950 430.950 283.050 433.050 ;
        RECT 274.950 416.250 277.050 417.150 ;
        RECT 277.950 415.950 280.050 418.050 ;
        RECT 281.400 415.050 282.450 430.950 ;
        RECT 284.400 427.050 285.450 517.950 ;
        RECT 305.400 517.050 306.450 535.950 ;
        RECT 308.400 529.050 309.450 550.950 ;
        RECT 317.400 538.050 318.450 550.950 ;
        RECT 328.950 541.950 331.050 544.050 ;
        RECT 329.400 538.050 330.450 541.950 ;
        RECT 316.950 535.950 319.050 538.050 ;
        RECT 325.950 535.950 328.050 538.050 ;
        RECT 328.950 535.950 331.050 538.050 ;
        RECT 326.400 529.050 327.450 535.950 ;
        RECT 331.950 532.950 334.050 535.050 ;
        RECT 307.950 528.450 310.050 529.050 ;
        RECT 316.950 528.450 319.050 529.050 ;
        RECT 307.950 527.400 312.450 528.450 ;
        RECT 307.950 526.950 310.050 527.400 ;
        RECT 307.950 524.850 310.050 525.750 ;
        RECT 295.950 514.950 298.050 517.050 ;
        RECT 304.950 514.950 307.050 517.050 ;
        RECT 289.950 490.950 292.050 493.050 ;
        RECT 290.400 487.050 291.450 490.950 ;
        RECT 286.950 485.250 289.050 486.150 ;
        RECT 289.950 484.950 292.050 487.050 ;
        RECT 292.950 485.250 295.050 486.150 ;
        RECT 286.950 481.950 289.050 484.050 ;
        RECT 290.250 482.250 291.750 483.150 ;
        RECT 292.950 481.950 295.050 484.050 ;
        RECT 287.400 475.050 288.450 481.950 ;
        RECT 293.400 481.050 294.450 481.950 ;
        RECT 289.950 478.950 292.050 481.050 ;
        RECT 292.950 478.950 295.050 481.050 ;
        RECT 286.950 472.950 289.050 475.050 ;
        RECT 287.400 457.050 288.450 472.950 ;
        RECT 296.400 472.050 297.450 514.950 ;
        RECT 311.400 504.450 312.450 527.400 ;
        RECT 316.950 527.400 321.450 528.450 ;
        RECT 316.950 526.950 319.050 527.400 ;
        RECT 313.950 524.250 316.050 525.150 ;
        RECT 316.950 524.850 319.050 525.750 ;
        RECT 320.400 523.050 321.450 527.400 ;
        RECT 322.950 526.950 325.050 529.050 ;
        RECT 325.950 526.950 328.050 529.050 ;
        RECT 323.400 525.450 324.450 526.950 ;
        RECT 332.400 526.050 333.450 532.950 ;
        RECT 325.950 525.450 328.050 526.050 ;
        RECT 323.400 524.400 328.050 525.450 ;
        RECT 313.950 522.450 316.050 523.050 ;
        RECT 313.950 521.400 318.450 522.450 ;
        RECT 313.950 520.950 316.050 521.400 ;
        RECT 317.400 520.050 318.450 521.400 ;
        RECT 319.950 520.950 322.050 523.050 ;
        RECT 323.400 520.050 324.450 524.400 ;
        RECT 325.950 523.950 328.050 524.400 ;
        RECT 331.950 523.950 334.050 526.050 ;
        RECT 335.250 524.250 337.050 525.150 ;
        RECT 325.950 521.850 327.750 522.750 ;
        RECT 328.950 520.950 331.050 523.050 ;
        RECT 332.250 521.850 333.750 522.750 ;
        RECT 334.950 522.450 337.050 523.050 ;
        RECT 338.400 522.450 339.450 571.950 ;
        RECT 341.400 559.050 342.450 574.950 ;
        RECT 352.950 559.950 355.050 562.050 ;
        RECT 340.950 556.950 343.050 559.050 ;
        RECT 343.950 557.250 346.050 558.150 ;
        RECT 349.950 557.250 352.050 558.150 ;
        RECT 353.400 556.050 354.450 559.950 ;
        RECT 356.400 556.050 357.450 592.950 ;
        RECT 343.950 553.950 346.050 556.050 ;
        RECT 347.250 554.250 348.750 555.150 ;
        RECT 349.950 553.950 352.050 556.050 ;
        RECT 352.950 553.950 355.050 556.050 ;
        RECT 355.950 553.950 358.050 556.050 ;
        RECT 350.400 553.050 351.450 553.950 ;
        RECT 346.950 550.950 349.050 553.050 ;
        RECT 349.950 550.950 352.050 553.050 ;
        RECT 356.400 547.050 357.450 553.950 ;
        RECT 355.950 544.950 358.050 547.050 ;
        RECT 359.400 544.050 360.450 625.950 ;
        RECT 362.400 622.050 363.450 646.950 ;
        RECT 365.400 628.050 366.450 665.400 ;
        RECT 374.400 652.050 375.450 673.950 ;
        RECT 373.950 649.950 376.050 652.050 ;
        RECT 377.400 643.050 378.450 700.950 ;
        RECT 383.400 700.050 384.450 719.400 ;
        RECT 386.400 706.050 387.450 737.400 ;
        RECT 395.400 733.050 396.450 739.950 ;
        RECT 397.950 736.950 400.050 739.050 ;
        RECT 401.400 738.450 402.450 751.950 ;
        RECT 407.400 742.050 408.450 754.950 ;
        RECT 403.950 740.250 405.750 741.150 ;
        RECT 406.950 739.950 409.050 742.050 ;
        RECT 410.400 739.050 411.450 754.950 ;
        RECT 416.400 747.450 417.450 772.950 ;
        RECT 421.950 769.950 424.050 772.050 ;
        RECT 430.950 769.950 433.050 772.050 ;
        RECT 437.400 771.450 438.450 776.400 ;
        RECT 439.950 775.950 442.050 776.400 ;
        RECT 443.250 776.250 444.750 777.150 ;
        RECT 445.950 776.400 450.450 777.450 ;
        RECT 445.950 775.950 448.050 776.400 ;
        RECT 439.950 773.850 441.750 774.750 ;
        RECT 442.950 772.950 445.050 775.050 ;
        RECT 446.250 773.850 448.050 774.750 ;
        RECT 437.400 770.400 441.450 771.450 ;
        RECT 422.400 757.050 423.450 769.950 ;
        RECT 433.950 760.950 436.050 763.050 ;
        RECT 421.950 754.950 424.050 757.050 ;
        RECT 418.950 751.950 421.050 754.050 ;
        RECT 419.400 748.050 420.450 751.950 ;
        RECT 413.400 746.400 417.450 747.450 ;
        RECT 413.400 742.050 414.450 746.400 ;
        RECT 418.950 745.950 421.050 748.050 ;
        RECT 415.950 743.250 418.050 744.150 ;
        RECT 418.950 743.850 421.050 744.750 ;
        RECT 424.950 744.450 427.050 745.050 ;
        RECT 421.950 743.250 423.750 744.150 ;
        RECT 424.950 743.400 429.450 744.450 ;
        RECT 424.950 742.950 427.050 743.400 ;
        RECT 412.950 739.950 415.050 742.050 ;
        RECT 415.950 739.950 418.050 742.050 ;
        RECT 421.950 739.950 424.050 742.050 ;
        RECT 425.250 740.850 427.050 741.750 ;
        RECT 422.400 739.050 423.450 739.950 ;
        RECT 403.950 738.450 406.050 739.050 ;
        RECT 401.400 737.400 406.050 738.450 ;
        RECT 407.250 737.850 408.750 738.750 ;
        RECT 403.950 736.950 406.050 737.400 ;
        RECT 409.950 736.950 412.050 739.050 ;
        RECT 413.250 737.850 415.050 738.750 ;
        RECT 421.950 736.950 424.050 739.050 ;
        RECT 394.950 730.950 397.050 733.050 ;
        RECT 391.950 707.250 394.050 708.150 ;
        RECT 385.950 703.950 388.050 706.050 ;
        RECT 389.250 704.250 390.750 705.150 ;
        RECT 391.950 703.950 394.050 706.050 ;
        RECT 395.250 704.250 397.050 705.150 ;
        RECT 385.950 701.850 387.750 702.750 ;
        RECT 388.950 700.950 391.050 703.050 ;
        RECT 391.950 700.950 394.050 703.050 ;
        RECT 394.950 700.950 397.050 703.050 ;
        RECT 382.950 697.950 385.050 700.050 ;
        RECT 382.950 694.950 385.050 697.050 ;
        RECT 385.950 694.950 388.050 697.050 ;
        RECT 383.400 676.050 384.450 694.950 ;
        RECT 382.950 673.950 385.050 676.050 ;
        RECT 386.400 673.050 387.450 694.950 ;
        RECT 389.400 694.050 390.450 700.950 ;
        RECT 388.950 691.950 391.050 694.050 ;
        RECT 392.400 679.050 393.450 700.950 ;
        RECT 398.400 699.450 399.450 736.950 ;
        RECT 409.950 734.850 412.050 735.750 ;
        RECT 428.400 706.050 429.450 743.400 ;
        RECT 434.400 742.050 435.450 760.950 ;
        RECT 440.400 751.050 441.450 770.400 ;
        RECT 443.400 768.450 444.450 772.950 ;
        RECT 449.400 769.050 450.450 776.400 ;
        RECT 451.950 775.950 454.050 778.050 ;
        RECT 454.950 775.950 457.050 778.050 ;
        RECT 458.250 776.250 459.750 777.150 ;
        RECT 460.950 775.950 463.050 778.050 ;
        RECT 445.950 768.450 448.050 769.050 ;
        RECT 443.400 767.400 448.050 768.450 ;
        RECT 445.950 766.950 448.050 767.400 ;
        RECT 448.950 766.950 451.050 769.050 ;
        RECT 452.400 753.450 453.450 775.950 ;
        RECT 454.950 773.850 456.750 774.750 ;
        RECT 457.950 772.950 460.050 775.050 ;
        RECT 461.250 773.850 463.050 774.750 ;
        RECT 458.400 772.050 459.450 772.950 ;
        RECT 464.400 772.050 465.450 802.950 ;
        RECT 457.950 769.950 460.050 772.050 ;
        RECT 463.950 769.950 466.050 772.050 ;
        RECT 457.950 766.950 460.050 769.050 ;
        RECT 452.400 752.400 456.450 753.450 ;
        RECT 439.950 748.950 442.050 751.050 ;
        RECT 451.950 748.950 454.050 751.050 ;
        RECT 436.950 743.250 439.050 744.150 ;
        RECT 433.950 739.950 436.050 742.050 ;
        RECT 436.950 741.450 439.050 742.050 ;
        RECT 440.400 741.450 441.450 748.950 ;
        RECT 445.950 747.450 448.050 748.050 ;
        RECT 445.950 746.400 450.450 747.450 ;
        RECT 445.950 745.950 448.050 746.400 ;
        RECT 442.950 742.950 445.050 745.050 ;
        RECT 446.250 743.850 448.050 744.750 ;
        RECT 436.950 740.400 441.450 741.450 ;
        RECT 442.950 740.850 445.050 741.750 ;
        RECT 436.950 739.950 439.050 740.400 ;
        RECT 433.950 709.950 436.050 712.050 ;
        RECT 418.950 703.950 421.050 706.050 ;
        RECT 421.950 704.250 424.050 705.150 ;
        RECT 427.950 703.950 430.050 706.050 ;
        RECT 400.950 702.450 403.050 703.050 ;
        RECT 403.950 702.450 406.050 703.050 ;
        RECT 400.950 701.400 406.050 702.450 ;
        RECT 400.950 700.950 403.050 701.400 ;
        RECT 403.950 700.950 406.050 701.400 ;
        RECT 409.950 700.950 412.050 703.050 ;
        RECT 413.250 701.250 415.050 702.150 ;
        RECT 415.950 700.950 418.050 703.050 ;
        RECT 419.400 702.450 420.450 703.950 ;
        RECT 421.950 702.450 424.050 703.050 ;
        RECT 419.400 701.400 424.050 702.450 ;
        RECT 421.950 700.950 424.050 701.400 ;
        RECT 425.250 701.250 426.750 702.150 ;
        RECT 427.950 700.950 430.050 703.050 ;
        RECT 431.250 701.250 433.050 702.150 ;
        RECT 395.400 698.400 399.450 699.450 ;
        RECT 388.950 676.950 391.050 679.050 ;
        RECT 391.950 676.950 394.050 679.050 ;
        RECT 389.400 673.050 390.450 676.950 ;
        RECT 385.950 670.950 388.050 673.050 ;
        RECT 388.950 670.950 391.050 673.050 ;
        RECT 379.950 668.250 381.750 669.150 ;
        RECT 382.950 667.950 385.050 670.050 ;
        RECT 386.400 667.050 387.450 670.950 ;
        RECT 388.950 667.950 391.050 670.050 ;
        RECT 379.950 664.950 382.050 667.050 ;
        RECT 383.250 665.850 384.750 666.750 ;
        RECT 385.950 664.950 388.050 667.050 ;
        RECT 389.250 665.850 391.050 666.750 ;
        RECT 380.400 649.050 381.450 664.950 ;
        RECT 385.950 662.850 388.050 663.750 ;
        RECT 392.400 655.050 393.450 676.950 ;
        RECT 391.950 652.950 394.050 655.050 ;
        RECT 379.950 646.950 382.050 649.050 ;
        RECT 379.950 643.950 382.050 646.050 ;
        RECT 376.950 640.950 379.050 643.050 ;
        RECT 376.950 634.950 379.050 637.050 ;
        RECT 377.400 634.050 378.450 634.950 ;
        RECT 367.950 633.450 370.050 634.050 ;
        RECT 370.950 633.450 373.050 634.050 ;
        RECT 367.950 632.400 373.050 633.450 ;
        RECT 367.950 631.950 370.050 632.400 ;
        RECT 370.950 631.950 373.050 632.400 ;
        RECT 374.250 632.250 375.750 633.150 ;
        RECT 376.950 631.950 379.050 634.050 ;
        RECT 364.950 625.950 367.050 628.050 ;
        RECT 368.400 625.050 369.450 631.950 ;
        RECT 370.950 629.850 372.750 630.750 ;
        RECT 373.950 628.950 376.050 631.050 ;
        RECT 377.250 629.850 379.050 630.750 ;
        RECT 374.400 628.050 375.450 628.950 ;
        RECT 380.400 628.050 381.450 643.950 ;
        RECT 391.950 640.950 394.050 643.050 ;
        RECT 382.950 629.250 385.050 630.150 ;
        RECT 388.950 629.250 391.050 630.150 ;
        RECT 373.950 625.950 376.050 628.050 ;
        RECT 379.950 625.950 382.050 628.050 ;
        RECT 382.950 625.950 385.050 628.050 ;
        RECT 386.250 626.250 387.750 627.150 ;
        RECT 388.950 625.950 391.050 628.050 ;
        RECT 383.400 625.050 384.450 625.950 ;
        RECT 364.950 622.950 367.050 625.050 ;
        RECT 367.950 622.950 370.050 625.050 ;
        RECT 376.950 622.950 379.050 625.050 ;
        RECT 382.950 622.950 385.050 625.050 ;
        RECT 385.950 624.450 388.050 625.050 ;
        RECT 388.950 624.450 391.050 625.050 ;
        RECT 385.950 623.400 391.050 624.450 ;
        RECT 385.950 622.950 388.050 623.400 ;
        RECT 388.950 622.950 391.050 623.400 ;
        RECT 361.950 619.950 364.050 622.050 ;
        RECT 361.950 607.950 364.050 610.050 ;
        RECT 362.400 553.050 363.450 607.950 ;
        RECT 365.400 607.050 366.450 622.950 ;
        RECT 367.950 613.950 370.050 616.050 ;
        RECT 364.950 604.950 367.050 607.050 ;
        RECT 365.400 568.050 366.450 604.950 ;
        RECT 368.400 601.050 369.450 613.950 ;
        RECT 370.950 601.950 373.050 604.050 ;
        RECT 367.950 598.950 370.050 601.050 ;
        RECT 371.250 599.850 372.750 600.750 ;
        RECT 373.950 598.950 376.050 601.050 ;
        RECT 377.400 598.050 378.450 622.950 ;
        RECT 379.950 619.950 382.050 622.050 ;
        RECT 380.400 604.050 381.450 619.950 ;
        RECT 385.950 607.950 388.050 610.050 ;
        RECT 379.950 601.950 382.050 604.050 ;
        RECT 379.950 599.850 382.050 600.750 ;
        RECT 382.950 599.250 385.050 600.150 ;
        RECT 367.950 596.850 370.050 597.750 ;
        RECT 373.950 596.850 376.050 597.750 ;
        RECT 376.950 595.950 379.050 598.050 ;
        RECT 382.950 595.950 385.050 598.050 ;
        RECT 386.400 594.450 387.450 607.950 ;
        RECT 388.950 601.950 391.050 604.050 ;
        RECT 383.400 593.400 387.450 594.450 ;
        RECT 370.950 568.950 373.050 571.050 ;
        RECT 364.950 565.950 367.050 568.050 ;
        RECT 365.400 559.050 366.450 565.950 ;
        RECT 371.400 562.050 372.450 568.950 ;
        RECT 376.950 563.250 379.050 564.150 ;
        RECT 383.400 562.050 384.450 593.400 ;
        RECT 370.950 559.950 373.050 562.050 ;
        RECT 373.950 560.250 375.750 561.150 ;
        RECT 376.950 559.950 379.050 562.050 ;
        RECT 380.250 560.250 381.750 561.150 ;
        RECT 382.950 559.950 385.050 562.050 ;
        RECT 385.950 559.950 388.050 562.050 ;
        RECT 364.950 556.950 367.050 559.050 ;
        RECT 373.950 556.950 376.050 559.050 ;
        RECT 376.950 556.950 379.050 559.050 ;
        RECT 379.950 556.950 382.050 559.050 ;
        RECT 383.250 557.850 385.050 558.750 ;
        RECT 364.950 554.850 367.050 555.750 ;
        RECT 367.950 554.250 370.050 555.150 ;
        RECT 373.950 553.950 376.050 556.050 ;
        RECT 361.950 550.950 364.050 553.050 ;
        RECT 367.950 550.950 370.050 553.050 ;
        RECT 343.950 541.950 346.050 544.050 ;
        RECT 358.950 541.950 361.050 544.050 ;
        RECT 334.950 521.400 339.450 522.450 ;
        RECT 334.950 520.950 337.050 521.400 ;
        RECT 316.950 517.950 319.050 520.050 ;
        RECT 322.950 517.950 325.050 520.050 ;
        RECT 328.950 518.850 331.050 519.750 ;
        RECT 311.400 503.400 315.450 504.450 ;
        RECT 304.950 499.950 307.050 502.050 ;
        RECT 305.400 490.050 306.450 499.950 ;
        RECT 304.950 489.450 307.050 490.050 ;
        RECT 302.400 488.400 307.050 489.450 ;
        RECT 298.950 485.250 301.050 486.150 ;
        RECT 298.950 481.950 301.050 484.050 ;
        RECT 292.950 469.950 295.050 472.050 ;
        RECT 295.950 469.950 298.050 472.050 ;
        RECT 293.400 468.450 294.450 469.950 ;
        RECT 293.400 467.400 297.450 468.450 ;
        RECT 289.950 457.950 292.050 460.050 ;
        RECT 286.950 454.950 289.050 457.050 ;
        RECT 290.400 454.050 291.450 457.950 ;
        RECT 296.400 454.050 297.450 467.400 ;
        RECT 299.400 460.050 300.450 481.950 ;
        RECT 298.950 457.950 301.050 460.050 ;
        RECT 289.950 451.950 292.050 454.050 ;
        RECT 295.950 451.950 298.050 454.050 ;
        RECT 299.250 452.250 301.050 453.150 ;
        RECT 302.400 451.050 303.450 488.400 ;
        RECT 304.950 487.950 307.050 488.400 ;
        RECT 304.950 485.850 307.050 486.750 ;
        RECT 307.950 485.250 310.050 486.150 ;
        RECT 307.950 481.950 310.050 484.050 ;
        RECT 308.400 478.050 309.450 481.950 ;
        RECT 307.950 475.950 310.050 478.050 ;
        RECT 310.950 472.950 313.050 475.050 ;
        RECT 304.950 469.950 307.050 472.050 ;
        RECT 289.950 449.850 291.750 450.750 ;
        RECT 292.950 448.950 295.050 451.050 ;
        RECT 296.250 449.850 297.750 450.750 ;
        RECT 298.950 448.950 301.050 451.050 ;
        RECT 301.950 448.950 304.050 451.050 ;
        RECT 299.400 448.050 300.450 448.950 ;
        RECT 292.950 446.850 295.050 447.750 ;
        RECT 298.950 445.950 301.050 448.050 ;
        RECT 305.400 442.050 306.450 469.950 ;
        RECT 307.950 457.950 310.050 460.050 ;
        RECT 308.400 451.050 309.450 457.950 ;
        RECT 311.400 454.050 312.450 472.950 ;
        RECT 314.400 457.050 315.450 503.400 ;
        RECT 317.400 484.050 318.450 517.950 ;
        RECT 331.950 511.950 334.050 514.050 ;
        RECT 325.950 491.250 328.050 492.150 ;
        RECT 319.950 487.950 322.050 490.050 ;
        RECT 323.250 488.250 324.750 489.150 ;
        RECT 325.950 487.950 328.050 490.050 ;
        RECT 329.250 488.250 331.050 489.150 ;
        RECT 326.400 487.050 327.450 487.950 ;
        RECT 319.950 485.850 321.750 486.750 ;
        RECT 322.950 484.950 325.050 487.050 ;
        RECT 325.950 484.950 328.050 487.050 ;
        RECT 328.950 484.950 331.050 487.050 ;
        RECT 323.400 484.050 324.450 484.950 ;
        RECT 316.950 481.950 319.050 484.050 ;
        RECT 322.950 481.950 325.050 484.050 ;
        RECT 316.950 478.950 319.050 481.050 ;
        RECT 317.400 472.050 318.450 478.950 ;
        RECT 319.950 475.950 322.050 478.050 ;
        RECT 316.950 469.950 319.050 472.050 ;
        RECT 316.950 460.950 319.050 463.050 ;
        RECT 313.950 454.950 316.050 457.050 ;
        RECT 317.400 454.050 318.450 460.950 ;
        RECT 320.400 457.050 321.450 475.950 ;
        RECT 323.400 457.050 324.450 481.950 ;
        RECT 325.950 460.950 328.050 463.050 ;
        RECT 319.950 454.950 322.050 457.050 ;
        RECT 322.950 454.950 325.050 457.050 ;
        RECT 310.950 451.950 313.050 454.050 ;
        RECT 313.950 451.950 316.050 454.050 ;
        RECT 316.950 451.950 319.050 454.050 ;
        RECT 320.250 452.250 322.050 453.150 ;
        RECT 314.400 451.050 315.450 451.950 ;
        RECT 307.950 448.950 310.050 451.050 ;
        RECT 310.950 449.850 312.750 450.750 ;
        RECT 313.950 448.950 316.050 451.050 ;
        RECT 317.250 449.850 318.750 450.750 ;
        RECT 319.950 448.950 322.050 451.050 ;
        RECT 307.950 445.950 310.050 448.050 ;
        RECT 310.950 445.950 313.050 448.050 ;
        RECT 313.950 446.850 316.050 447.750 ;
        RECT 308.400 442.050 309.450 445.950 ;
        RECT 292.950 439.950 295.050 442.050 ;
        RECT 304.950 439.950 307.050 442.050 ;
        RECT 307.950 439.950 310.050 442.050 ;
        RECT 289.950 436.950 292.050 439.050 ;
        RECT 283.950 424.950 286.050 427.050 ;
        RECT 290.400 415.050 291.450 436.950 ;
        RECT 274.950 412.950 277.050 415.050 ;
        RECT 278.250 413.250 279.750 414.150 ;
        RECT 280.950 412.950 283.050 415.050 ;
        RECT 284.250 413.250 286.050 414.150 ;
        RECT 289.950 412.950 292.050 415.050 ;
        RECT 277.950 409.950 280.050 412.050 ;
        RECT 281.250 410.850 282.750 411.750 ;
        RECT 283.950 409.950 286.050 412.050 ;
        RECT 286.950 410.250 289.050 411.150 ;
        RECT 289.950 410.850 292.050 411.750 ;
        RECT 286.950 406.950 289.050 409.050 ;
        RECT 271.950 403.950 274.050 406.050 ;
        RECT 274.950 403.950 277.050 406.050 ;
        RECT 275.400 400.050 276.450 403.950 ;
        RECT 274.950 397.950 277.050 400.050 ;
        RECT 283.950 397.950 286.050 400.050 ;
        RECT 280.950 391.950 283.050 394.050 ;
        RECT 268.950 385.950 271.050 388.050 ;
        RECT 281.400 385.050 282.450 391.950 ;
        RECT 268.950 384.450 271.050 385.050 ;
        RECT 266.400 383.400 271.050 384.450 ;
        RECT 268.950 382.950 271.050 383.400 ;
        RECT 272.250 383.250 273.750 384.150 ;
        RECT 274.950 382.950 277.050 385.050 ;
        RECT 278.250 383.250 279.750 384.150 ;
        RECT 280.950 382.950 283.050 385.050 ;
        RECT 268.950 380.850 270.750 381.750 ;
        RECT 271.950 379.950 274.050 382.050 ;
        RECT 275.250 380.850 276.750 381.750 ;
        RECT 277.950 379.950 280.050 382.050 ;
        RECT 281.250 380.850 283.050 381.750 ;
        RECT 265.950 346.950 268.050 349.050 ;
        RECT 262.950 334.950 265.050 337.050 ;
        RECT 257.400 320.400 261.450 321.450 ;
        RECT 224.400 316.050 225.450 319.950 ;
        RECT 227.400 317.400 246.450 318.450 ;
        RECT 205.950 313.950 208.050 316.050 ;
        RECT 217.950 313.950 220.050 316.050 ;
        RECT 220.950 313.950 223.050 316.050 ;
        RECT 223.950 313.950 226.050 316.050 ;
        RECT 196.950 310.950 199.050 313.050 ;
        RECT 199.950 310.950 202.050 313.050 ;
        RECT 203.250 311.250 204.750 312.150 ;
        RECT 205.950 310.950 208.050 313.050 ;
        RECT 211.950 312.450 214.050 313.050 ;
        RECT 209.250 311.250 210.750 312.150 ;
        RECT 211.950 311.400 216.450 312.450 ;
        RECT 211.950 310.950 214.050 311.400 ;
        RECT 175.950 286.950 178.050 289.050 ;
        RECT 193.950 286.950 196.050 289.050 ;
        RECT 176.400 277.050 177.450 286.950 ;
        RECT 178.950 280.950 181.050 283.050 ;
        RECT 175.950 274.950 178.050 277.050 ;
        RECT 179.400 274.050 180.450 280.950 ;
        RECT 187.950 277.950 190.050 280.050 ;
        RECT 178.950 271.950 181.050 274.050 ;
        RECT 181.950 271.950 184.050 274.050 ;
        RECT 175.950 269.250 178.050 270.150 ;
        RECT 178.950 269.850 181.050 270.750 ;
        RECT 175.950 265.950 178.050 268.050 ;
        RECT 176.400 262.050 177.450 265.950 ;
        RECT 175.950 259.950 178.050 262.050 ;
        RECT 182.400 253.050 183.450 271.950 ;
        RECT 184.950 269.250 187.050 270.150 ;
        RECT 184.950 265.950 187.050 268.050 ;
        RECT 181.950 250.950 184.050 253.050 ;
        RECT 188.400 247.050 189.450 277.950 ;
        RECT 197.400 277.050 198.450 310.950 ;
        RECT 199.950 308.850 201.750 309.750 ;
        RECT 202.950 307.950 205.050 310.050 ;
        RECT 206.250 308.850 207.750 309.750 ;
        RECT 208.950 307.950 211.050 310.050 ;
        RECT 212.250 308.850 214.050 309.750 ;
        RECT 203.400 304.050 204.450 307.950 ;
        RECT 202.950 301.950 205.050 304.050 ;
        RECT 205.950 298.950 208.050 301.050 ;
        RECT 202.950 295.950 205.050 298.050 ;
        RECT 199.950 280.950 202.050 283.050 ;
        RECT 196.950 274.950 199.050 277.050 ;
        RECT 200.400 274.050 201.450 280.950 ;
        RECT 193.950 273.450 196.050 274.050 ;
        RECT 191.400 272.400 196.050 273.450 ;
        RECT 191.400 265.050 192.450 272.400 ;
        RECT 193.950 271.950 196.050 272.400 ;
        RECT 197.250 272.250 198.750 273.150 ;
        RECT 199.950 271.950 202.050 274.050 ;
        RECT 193.950 269.850 195.750 270.750 ;
        RECT 196.950 268.950 199.050 271.050 ;
        RECT 200.250 269.850 202.050 270.750 ;
        RECT 197.400 268.050 198.450 268.950 ;
        RECT 196.950 265.950 199.050 268.050 ;
        RECT 190.950 262.950 193.050 265.050 ;
        RECT 175.950 244.950 178.050 247.050 ;
        RECT 187.950 244.950 190.050 247.050 ;
        RECT 199.950 244.950 202.050 247.050 ;
        RECT 176.400 244.050 177.450 244.950 ;
        RECT 175.950 241.950 178.050 244.050 ;
        RECT 181.950 241.950 184.050 244.050 ;
        RECT 193.950 241.950 196.050 244.050 ;
        RECT 175.950 239.850 178.050 240.750 ;
        RECT 178.950 239.250 181.050 240.150 ;
        RECT 178.950 235.950 181.050 238.050 ;
        RECT 182.400 235.050 183.450 241.950 ;
        RECT 194.400 241.050 195.450 241.950 ;
        RECT 187.950 240.450 190.050 241.050 ;
        RECT 185.400 239.400 190.050 240.450 ;
        RECT 185.400 238.050 186.450 239.400 ;
        RECT 187.950 238.950 190.050 239.400 ;
        RECT 191.250 239.250 192.750 240.150 ;
        RECT 193.950 238.950 196.050 241.050 ;
        RECT 196.950 238.950 199.050 241.050 ;
        RECT 197.400 238.050 198.450 238.950 ;
        RECT 184.950 235.950 187.050 238.050 ;
        RECT 187.950 236.850 189.750 237.750 ;
        RECT 190.950 235.950 193.050 238.050 ;
        RECT 194.250 236.850 195.750 237.750 ;
        RECT 196.950 235.950 199.050 238.050 ;
        RECT 181.950 232.950 184.050 235.050 ;
        RECT 173.400 227.400 177.450 228.450 ;
        RECT 166.950 203.250 169.050 204.150 ;
        RECT 163.950 200.250 165.750 201.150 ;
        RECT 166.950 199.950 169.050 202.050 ;
        RECT 170.250 200.250 171.750 201.150 ;
        RECT 172.950 199.950 175.050 202.050 ;
        RECT 160.950 196.950 163.050 199.050 ;
        RECT 163.950 196.950 166.050 199.050 ;
        RECT 169.950 196.950 172.050 199.050 ;
        RECT 173.250 197.850 175.050 198.750 ;
        RECT 154.950 194.400 159.450 195.450 ;
        RECT 154.950 193.950 157.050 194.400 ;
        RECT 146.400 193.050 147.450 193.950 ;
        RECT 127.950 190.950 130.050 193.050 ;
        RECT 142.950 190.950 145.050 193.050 ;
        RECT 145.950 190.950 148.050 193.050 ;
        RECT 122.400 179.400 126.450 180.450 ;
        RECT 122.400 151.050 123.450 179.400 ;
        RECT 128.400 166.050 129.450 190.950 ;
        RECT 149.400 190.050 150.450 193.950 ;
        RECT 164.400 193.050 165.450 196.950 ;
        RECT 163.950 190.950 166.050 193.050 ;
        RECT 133.950 187.950 136.050 190.050 ;
        RECT 148.950 187.950 151.050 190.050 ;
        RECT 166.950 187.950 169.050 190.050 ;
        RECT 124.950 164.250 126.750 165.150 ;
        RECT 127.950 163.950 130.050 166.050 ;
        RECT 131.250 164.250 133.050 165.150 ;
        RECT 124.950 160.950 127.050 163.050 ;
        RECT 128.250 161.850 129.750 162.750 ;
        RECT 130.950 160.950 133.050 163.050 ;
        RECT 125.400 154.050 126.450 160.950 ;
        RECT 131.400 159.450 132.450 160.950 ;
        RECT 128.400 158.400 132.450 159.450 ;
        RECT 128.400 157.050 129.450 158.400 ;
        RECT 134.400 157.050 135.450 187.950 ;
        RECT 148.950 184.950 151.050 187.050 ;
        RECT 136.950 181.950 139.050 184.050 ;
        RECT 137.400 166.050 138.450 181.950 ;
        RECT 145.950 172.950 148.050 175.050 ;
        RECT 146.400 172.050 147.450 172.950 ;
        RECT 142.950 169.950 145.050 172.050 ;
        RECT 145.950 169.950 148.050 172.050 ;
        RECT 143.400 166.050 144.450 169.950 ;
        RECT 136.950 163.950 139.050 166.050 ;
        RECT 142.950 163.950 145.050 166.050 ;
        RECT 146.250 164.250 148.050 165.150 ;
        RECT 136.950 161.850 138.750 162.750 ;
        RECT 139.950 160.950 142.050 163.050 ;
        RECT 143.250 161.850 144.750 162.750 ;
        RECT 145.950 160.950 148.050 163.050 ;
        RECT 139.950 158.850 142.050 159.750 ;
        RECT 145.950 157.950 148.050 160.050 ;
        RECT 127.950 154.950 130.050 157.050 ;
        RECT 133.950 154.950 136.050 157.050 ;
        RECT 124.950 151.950 127.050 154.050 ;
        RECT 121.950 148.950 124.050 151.050 ;
        RECT 118.950 142.950 121.050 145.050 ;
        RECT 112.950 139.950 115.050 142.050 ;
        RECT 118.950 130.950 121.050 133.050 ;
        RECT 119.400 127.050 120.450 130.950 ;
        RECT 124.950 128.250 127.050 129.150 ;
        RECT 115.950 125.250 117.750 126.150 ;
        RECT 118.950 124.950 121.050 127.050 ;
        RECT 122.250 125.250 123.750 126.150 ;
        RECT 124.950 124.950 127.050 127.050 ;
        RECT 112.950 121.950 115.050 124.050 ;
        RECT 115.950 121.950 118.050 124.050 ;
        RECT 119.250 122.850 120.750 123.750 ;
        RECT 121.950 121.950 124.050 124.050 ;
        RECT 109.950 115.950 112.050 118.050 ;
        RECT 101.400 98.400 105.450 99.450 ;
        RECT 101.400 97.050 102.450 98.400 ;
        RECT 100.950 94.950 103.050 97.050 ;
        RECT 104.250 95.250 105.750 96.150 ;
        RECT 106.950 94.950 109.050 97.050 ;
        RECT 113.400 94.050 114.450 121.950 ;
        RECT 100.950 92.850 102.750 93.750 ;
        RECT 103.950 91.950 106.050 94.050 ;
        RECT 107.250 92.850 108.750 93.750 ;
        RECT 109.950 91.950 112.050 94.050 ;
        RECT 112.950 91.950 115.050 94.050 ;
        RECT 106.950 88.950 109.050 91.050 ;
        RECT 109.950 89.850 112.050 90.750 ;
        RECT 97.950 64.950 100.050 67.050 ;
        RECT 97.950 61.950 100.050 64.050 ;
        RECT 98.400 61.050 99.450 61.950 ;
        RECT 97.950 58.950 100.050 61.050 ;
        RECT 103.950 58.950 106.050 61.050 ;
        RECT 98.400 58.050 99.450 58.950 ;
        RECT 104.400 58.050 105.450 58.950 ;
        RECT 97.950 55.950 100.050 58.050 ;
        RECT 101.250 56.250 102.750 57.150 ;
        RECT 103.950 55.950 106.050 58.050 ;
        RECT 97.950 53.850 99.750 54.750 ;
        RECT 100.950 52.950 103.050 55.050 ;
        RECT 104.250 53.850 106.050 54.750 ;
        RECT 101.400 52.050 102.450 52.950 ;
        RECT 100.950 49.950 103.050 52.050 ;
        RECT 107.400 43.050 108.450 88.950 ;
        RECT 109.950 64.950 112.050 67.050 ;
        RECT 110.400 58.050 111.450 64.950 ;
        RECT 116.400 58.050 117.450 121.950 ;
        RECT 122.400 121.050 123.450 121.950 ;
        RECT 121.950 118.950 124.050 121.050 ;
        RECT 125.400 103.050 126.450 124.950 ;
        RECT 128.400 121.050 129.450 154.950 ;
        RECT 130.950 142.950 133.050 145.050 ;
        RECT 127.950 118.950 130.050 121.050 ;
        RECT 124.950 100.950 127.050 103.050 ;
        RECT 127.950 99.450 130.050 100.050 ;
        RECT 131.400 99.450 132.450 142.950 ;
        RECT 136.950 130.950 139.050 133.050 ;
        RECT 137.400 127.050 138.450 130.950 ;
        RECT 142.950 128.250 145.050 129.150 ;
        RECT 133.950 125.250 135.750 126.150 ;
        RECT 136.950 124.950 139.050 127.050 ;
        RECT 140.250 125.250 141.750 126.150 ;
        RECT 142.950 124.950 145.050 127.050 ;
        RECT 133.950 121.950 136.050 124.050 ;
        RECT 137.250 122.850 138.750 123.750 ;
        RECT 139.950 121.950 142.050 124.050 ;
        RECT 140.400 121.050 141.450 121.950 ;
        RECT 139.950 118.950 142.050 121.050 ;
        RECT 143.400 118.050 144.450 124.950 ;
        RECT 142.950 115.950 145.050 118.050 ;
        RECT 146.400 106.050 147.450 157.950 ;
        RECT 149.400 118.050 150.450 184.950 ;
        RECT 163.950 178.950 166.050 181.050 ;
        RECT 160.950 172.950 163.050 175.050 ;
        RECT 154.950 169.950 157.050 172.050 ;
        RECT 161.400 169.050 162.450 172.950 ;
        RECT 151.950 167.250 154.050 168.150 ;
        RECT 154.950 167.850 157.050 168.750 ;
        RECT 157.950 167.250 159.750 168.150 ;
        RECT 160.950 166.950 163.050 169.050 ;
        RECT 151.950 163.950 154.050 166.050 ;
        RECT 157.950 163.950 160.050 166.050 ;
        RECT 161.250 164.850 163.050 165.750 ;
        RECT 152.400 163.050 153.450 163.950 ;
        RECT 158.400 163.050 159.450 163.950 ;
        RECT 164.400 163.050 165.450 178.950 ;
        RECT 167.400 169.050 168.450 187.950 ;
        RECT 172.950 181.950 175.050 184.050 ;
        RECT 173.400 169.050 174.450 181.950 ;
        RECT 176.400 172.050 177.450 227.400 ;
        RECT 178.950 202.950 181.050 205.050 ;
        RECT 179.400 198.450 180.450 202.950 ;
        RECT 185.400 202.050 186.450 235.950 ;
        RECT 191.400 205.050 192.450 235.950 ;
        RECT 196.950 233.850 199.050 234.750 ;
        RECT 200.400 229.050 201.450 244.950 ;
        RECT 199.950 226.950 202.050 229.050 ;
        RECT 193.950 223.950 196.050 226.050 ;
        RECT 187.950 202.950 190.050 205.050 ;
        RECT 190.950 202.950 193.050 205.050 ;
        RECT 181.950 200.250 184.050 201.150 ;
        RECT 184.950 199.950 187.050 202.050 ;
        RECT 188.400 199.050 189.450 202.950 ;
        RECT 181.950 198.450 184.050 199.050 ;
        RECT 179.400 197.400 184.050 198.450 ;
        RECT 181.950 196.950 184.050 197.400 ;
        RECT 185.250 197.250 186.750 198.150 ;
        RECT 187.950 196.950 190.050 199.050 ;
        RECT 191.250 197.250 193.050 198.150 ;
        RECT 178.950 193.950 181.050 196.050 ;
        RECT 184.950 193.950 187.050 196.050 ;
        RECT 188.250 194.850 189.750 195.750 ;
        RECT 190.950 193.950 193.050 196.050 ;
        RECT 179.400 178.050 180.450 193.950 ;
        RECT 178.950 175.950 181.050 178.050 ;
        RECT 175.950 169.950 178.050 172.050 ;
        RECT 185.400 169.050 186.450 193.950 ;
        RECT 194.400 190.050 195.450 223.950 ;
        RECT 199.950 202.950 202.050 205.050 ;
        RECT 200.400 199.050 201.450 202.950 ;
        RECT 199.950 196.950 202.050 199.050 ;
        RECT 196.950 194.250 199.050 195.150 ;
        RECT 199.950 194.850 202.050 195.750 ;
        RECT 196.950 190.950 199.050 193.050 ;
        RECT 193.950 187.950 196.050 190.050 ;
        RECT 203.400 187.050 204.450 295.950 ;
        RECT 206.400 267.450 207.450 298.950 ;
        RECT 209.400 298.050 210.450 307.950 ;
        RECT 208.950 295.950 211.050 298.050 ;
        RECT 215.400 295.050 216.450 311.400 ;
        RECT 214.950 292.950 217.050 295.050 ;
        RECT 215.400 274.050 216.450 292.950 ;
        RECT 214.950 271.950 217.050 274.050 ;
        RECT 218.400 271.050 219.450 313.950 ;
        RECT 221.400 313.050 222.450 313.950 ;
        RECT 227.400 313.050 228.450 317.400 ;
        RECT 245.400 316.050 246.450 317.400 ;
        RECT 238.950 313.950 241.050 316.050 ;
        RECT 244.950 313.950 247.050 316.050 ;
        RECT 220.950 310.950 223.050 313.050 ;
        RECT 224.250 311.250 225.750 312.150 ;
        RECT 226.950 310.950 229.050 313.050 ;
        RECT 232.950 312.450 235.050 313.050 ;
        RECT 230.250 311.250 231.750 312.150 ;
        RECT 232.950 311.400 237.450 312.450 ;
        RECT 232.950 310.950 235.050 311.400 ;
        RECT 220.950 308.850 222.750 309.750 ;
        RECT 223.950 307.950 226.050 310.050 ;
        RECT 227.250 308.850 228.750 309.750 ;
        RECT 229.950 307.950 232.050 310.050 ;
        RECT 233.250 308.850 235.050 309.750 ;
        RECT 224.400 304.050 225.450 307.950 ;
        RECT 223.950 301.950 226.050 304.050 ;
        RECT 230.400 283.050 231.450 307.950 ;
        RECT 236.400 295.050 237.450 311.400 ;
        RECT 239.400 309.450 240.450 313.950 ;
        RECT 241.950 311.250 244.050 312.150 ;
        RECT 244.950 311.850 247.050 312.750 ;
        RECT 250.950 312.450 253.050 313.050 ;
        RECT 247.950 311.250 249.750 312.150 ;
        RECT 250.950 311.400 255.450 312.450 ;
        RECT 250.950 310.950 253.050 311.400 ;
        RECT 241.950 309.450 244.050 310.050 ;
        RECT 239.400 308.400 244.050 309.450 ;
        RECT 241.950 307.950 244.050 308.400 ;
        RECT 247.950 307.950 250.050 310.050 ;
        RECT 251.250 308.850 253.050 309.750 ;
        RECT 238.950 304.950 241.050 307.050 ;
        RECT 250.950 304.950 253.050 307.050 ;
        RECT 235.950 292.950 238.050 295.050 ;
        RECT 239.400 291.450 240.450 304.950 ;
        RECT 236.400 290.400 240.450 291.450 ;
        RECT 232.950 286.950 235.050 289.050 ;
        RECT 233.400 283.050 234.450 286.950 ;
        RECT 229.950 280.950 232.050 283.050 ;
        RECT 232.950 280.950 235.050 283.050 ;
        RECT 220.950 274.950 223.050 277.050 ;
        RECT 221.400 271.050 222.450 274.950 ;
        RECT 232.950 272.250 235.050 273.150 ;
        RECT 208.950 269.250 210.750 270.150 ;
        RECT 211.950 268.950 214.050 271.050 ;
        RECT 217.950 268.950 220.050 271.050 ;
        RECT 220.950 268.950 223.050 271.050 ;
        RECT 223.950 269.250 225.750 270.150 ;
        RECT 226.950 268.950 229.050 271.050 ;
        RECT 230.250 269.250 231.750 270.150 ;
        RECT 232.950 268.950 235.050 271.050 ;
        RECT 233.400 268.050 234.450 268.950 ;
        RECT 208.950 267.450 211.050 268.050 ;
        RECT 206.400 266.400 211.050 267.450 ;
        RECT 212.250 266.850 214.050 267.750 ;
        RECT 208.950 265.950 211.050 266.400 ;
        RECT 214.950 266.250 217.050 267.150 ;
        RECT 217.950 266.850 220.050 267.750 ;
        RECT 220.950 267.450 223.050 268.050 ;
        RECT 223.950 267.450 226.050 268.050 ;
        RECT 220.950 266.400 226.050 267.450 ;
        RECT 227.250 266.850 228.750 267.750 ;
        RECT 220.950 265.950 223.050 266.400 ;
        RECT 223.950 265.950 226.050 266.400 ;
        RECT 229.950 265.950 232.050 268.050 ;
        RECT 232.950 265.950 235.050 268.050 ;
        RECT 214.950 262.950 217.050 265.050 ;
        RECT 221.400 264.450 222.450 265.950 ;
        RECT 230.400 265.050 231.450 265.950 ;
        RECT 236.400 265.050 237.450 290.400 ;
        RECT 247.950 289.950 250.050 292.050 ;
        RECT 248.400 274.050 249.450 289.950 ;
        RECT 241.950 273.450 244.050 274.050 ;
        RECT 239.400 272.400 244.050 273.450 ;
        RECT 239.400 271.050 240.450 272.400 ;
        RECT 241.950 271.950 244.050 272.400 ;
        RECT 245.250 272.250 246.750 273.150 ;
        RECT 247.950 271.950 250.050 274.050 ;
        RECT 238.950 268.950 241.050 271.050 ;
        RECT 241.950 269.850 243.750 270.750 ;
        RECT 244.950 268.950 247.050 271.050 ;
        RECT 248.250 269.850 250.050 270.750 ;
        RECT 218.400 263.400 222.450 264.450 ;
        RECT 215.400 250.050 216.450 262.950 ;
        RECT 214.950 247.950 217.050 250.050 ;
        RECT 208.950 241.950 211.050 244.050 ;
        RECT 214.950 241.950 217.050 244.050 ;
        RECT 205.950 238.950 208.050 241.050 ;
        RECT 205.950 236.850 208.050 237.750 ;
        RECT 205.950 226.950 208.050 229.050 ;
        RECT 202.950 184.950 205.050 187.050 ;
        RECT 190.950 172.950 193.050 175.050 ;
        RECT 191.400 172.050 192.450 172.950 ;
        RECT 206.400 172.050 207.450 226.950 ;
        RECT 209.400 195.450 210.450 241.950 ;
        RECT 215.400 241.050 216.450 241.950 ;
        RECT 214.950 238.950 217.050 241.050 ;
        RECT 211.950 236.250 214.050 237.150 ;
        RECT 214.950 236.850 217.050 237.750 ;
        RECT 211.950 232.950 214.050 235.050 ;
        RECT 211.950 229.950 214.050 232.050 ;
        RECT 212.400 202.050 213.450 229.950 ;
        RECT 218.400 208.050 219.450 263.400 ;
        RECT 229.950 262.950 232.050 265.050 ;
        RECT 235.950 262.950 238.050 265.050 ;
        RECT 220.950 256.950 223.050 259.050 ;
        RECT 221.400 223.050 222.450 256.950 ;
        RECT 239.400 250.050 240.450 268.950 ;
        RECT 238.950 247.950 241.050 250.050 ;
        RECT 232.950 244.950 235.050 247.050 ;
        RECT 226.950 238.950 229.050 241.050 ;
        RECT 227.400 238.050 228.450 238.950 ;
        RECT 223.950 236.250 225.750 237.150 ;
        RECT 226.950 235.950 229.050 238.050 ;
        RECT 230.250 236.250 232.050 237.150 ;
        RECT 223.950 232.950 226.050 235.050 ;
        RECT 227.250 233.850 228.750 234.750 ;
        RECT 229.950 232.950 232.050 235.050 ;
        RECT 224.400 229.050 225.450 232.950 ;
        RECT 223.950 226.950 226.050 229.050 ;
        RECT 220.950 220.950 223.050 223.050 ;
        RECT 229.950 208.950 232.050 211.050 ;
        RECT 217.950 205.950 220.050 208.050 ;
        RECT 226.950 202.950 229.050 205.050 ;
        RECT 211.950 199.950 214.050 202.050 ;
        RECT 214.950 199.950 217.050 202.050 ;
        RECT 215.400 199.050 216.450 199.950 ;
        RECT 211.950 197.250 213.750 198.150 ;
        RECT 214.950 196.950 217.050 199.050 ;
        RECT 218.250 197.250 219.750 198.150 ;
        RECT 220.950 196.950 223.050 199.050 ;
        RECT 224.250 197.250 226.050 198.150 ;
        RECT 227.400 196.050 228.450 202.950 ;
        RECT 211.950 195.450 214.050 196.050 ;
        RECT 209.400 194.400 214.050 195.450 ;
        RECT 215.250 194.850 216.750 195.750 ;
        RECT 211.950 193.950 214.050 194.400 ;
        RECT 217.950 193.950 220.050 196.050 ;
        RECT 221.250 194.850 222.750 195.750 ;
        RECT 223.950 195.450 226.050 196.050 ;
        RECT 226.950 195.450 229.050 196.050 ;
        RECT 223.950 194.400 229.050 195.450 ;
        RECT 223.950 193.950 226.050 194.400 ;
        RECT 226.950 193.950 229.050 194.400 ;
        RECT 214.950 190.950 217.050 193.050 ;
        RECT 208.950 181.950 211.050 184.050 ;
        RECT 190.950 169.950 193.050 172.050 ;
        RECT 205.950 169.950 208.050 172.050 ;
        RECT 209.400 169.050 210.450 181.950 ;
        RECT 211.950 178.950 214.050 181.050 ;
        RECT 166.950 166.950 169.050 169.050 ;
        RECT 172.950 166.950 175.050 169.050 ;
        RECT 176.250 167.250 177.750 168.150 ;
        RECT 178.950 166.950 181.050 169.050 ;
        RECT 184.950 166.950 187.050 169.050 ;
        RECT 187.950 167.250 190.050 168.150 ;
        RECT 190.950 167.850 193.050 168.750 ;
        RECT 196.950 168.450 199.050 169.050 ;
        RECT 193.950 167.250 195.750 168.150 ;
        RECT 196.950 167.400 201.450 168.450 ;
        RECT 196.950 166.950 199.050 167.400 ;
        RECT 166.950 163.950 169.050 166.050 ;
        RECT 169.950 163.950 172.050 166.050 ;
        RECT 172.950 164.850 174.750 165.750 ;
        RECT 175.950 163.950 178.050 166.050 ;
        RECT 179.250 164.850 180.750 165.750 ;
        RECT 181.950 165.450 184.050 166.050 ;
        RECT 181.950 164.400 186.450 165.450 ;
        RECT 181.950 163.950 184.050 164.400 ;
        RECT 151.950 160.950 154.050 163.050 ;
        RECT 154.950 160.950 157.050 163.050 ;
        RECT 157.950 160.950 160.050 163.050 ;
        RECT 163.950 160.950 166.050 163.050 ;
        RECT 155.400 159.450 156.450 160.950 ;
        RECT 155.400 158.400 159.450 159.450 ;
        RECT 151.950 148.950 154.050 151.050 ;
        RECT 148.950 115.950 151.050 118.050 ;
        RECT 133.950 103.950 136.050 106.050 ;
        RECT 145.950 103.950 148.050 106.050 ;
        RECT 148.950 103.950 151.050 106.050 ;
        RECT 127.950 98.400 132.450 99.450 ;
        RECT 127.950 97.950 130.050 98.400 ;
        RECT 131.400 97.050 132.450 98.400 ;
        RECT 134.400 97.050 135.450 103.950 ;
        RECT 124.950 95.250 127.050 96.150 ;
        RECT 127.950 95.850 130.050 96.750 ;
        RECT 130.950 94.950 133.050 97.050 ;
        RECT 133.950 94.950 136.050 97.050 ;
        RECT 139.950 96.450 142.050 97.050 ;
        RECT 137.250 95.250 138.750 96.150 ;
        RECT 139.950 95.400 147.450 96.450 ;
        RECT 139.950 94.950 142.050 95.400 ;
        RECT 124.950 91.950 127.050 94.050 ;
        RECT 133.950 92.850 135.750 93.750 ;
        RECT 136.950 91.950 139.050 94.050 ;
        RECT 140.250 92.850 141.750 93.750 ;
        RECT 142.950 91.950 145.050 94.050 ;
        RECT 125.400 67.050 126.450 91.950 ;
        RECT 133.950 82.950 136.050 85.050 ;
        RECT 118.950 64.950 121.050 67.050 ;
        RECT 124.950 64.950 127.050 67.050 ;
        RECT 109.950 55.950 112.050 58.050 ;
        RECT 113.250 56.250 114.750 57.150 ;
        RECT 115.950 55.950 118.050 58.050 ;
        RECT 109.950 53.850 111.750 54.750 ;
        RECT 112.950 52.950 115.050 55.050 ;
        RECT 116.250 53.850 118.050 54.750 ;
        RECT 113.400 46.050 114.450 52.950 ;
        RECT 119.400 51.450 120.450 64.950 ;
        RECT 130.950 55.950 133.050 58.050 ;
        RECT 121.950 53.250 124.050 54.150 ;
        RECT 127.950 53.250 130.050 54.150 ;
        RECT 121.950 51.450 124.050 52.050 ;
        RECT 119.400 50.400 124.050 51.450 ;
        RECT 127.950 51.450 130.050 52.050 ;
        RECT 131.400 51.450 132.450 55.950 ;
        RECT 121.950 49.950 124.050 50.400 ;
        RECT 125.250 50.250 126.750 51.150 ;
        RECT 127.950 50.400 132.450 51.450 ;
        RECT 127.950 49.950 130.050 50.400 ;
        RECT 124.950 46.950 127.050 49.050 ;
        RECT 112.950 43.950 115.050 46.050 ;
        RECT 106.950 40.950 109.050 43.050 ;
        RECT 94.950 28.950 97.050 31.050 ;
        RECT 115.950 28.950 118.050 31.050 ;
        RECT 106.950 25.950 109.050 28.050 ;
        RECT 107.400 25.050 108.450 25.950 ;
        RECT 116.400 25.050 117.450 28.950 ;
        RECT 125.400 28.050 126.450 46.950 ;
        RECT 128.400 34.050 129.450 49.950 ;
        RECT 134.400 46.050 135.450 82.950 ;
        RECT 137.400 49.050 138.450 91.950 ;
        RECT 142.950 89.850 145.050 90.750 ;
        RECT 146.400 61.050 147.450 95.400 ;
        RECT 145.950 58.950 148.050 61.050 ;
        RECT 149.400 58.050 150.450 103.950 ;
        RECT 152.400 103.050 153.450 148.950 ;
        RECT 154.950 142.950 157.050 145.050 ;
        RECT 155.400 127.050 156.450 142.950 ;
        RECT 158.400 130.050 159.450 158.400 ;
        RECT 167.400 133.050 168.450 163.950 ;
        RECT 163.950 131.250 166.050 132.150 ;
        RECT 166.950 130.950 169.050 133.050 ;
        RECT 157.950 127.950 160.050 130.050 ;
        RECT 161.250 128.250 162.750 129.150 ;
        RECT 163.950 127.950 166.050 130.050 ;
        RECT 167.250 128.250 169.050 129.150 ;
        RECT 154.950 124.950 157.050 127.050 ;
        RECT 157.950 125.850 159.750 126.750 ;
        RECT 160.950 124.950 163.050 127.050 ;
        RECT 161.400 121.050 162.450 124.950 ;
        RECT 160.950 118.950 163.050 121.050 ;
        RECT 164.400 115.050 165.450 127.950 ;
        RECT 166.950 124.950 169.050 127.050 ;
        RECT 170.400 124.050 171.450 163.950 ;
        RECT 176.400 160.050 177.450 163.950 ;
        RECT 185.400 163.050 186.450 164.400 ;
        RECT 187.950 163.950 190.050 166.050 ;
        RECT 193.950 163.950 196.050 166.050 ;
        RECT 197.250 164.850 199.050 165.750 ;
        RECT 178.950 160.950 181.050 163.050 ;
        RECT 181.950 161.850 184.050 162.750 ;
        RECT 184.950 160.950 187.050 163.050 ;
        RECT 175.950 157.950 178.050 160.050 ;
        RECT 179.400 154.050 180.450 160.950 ;
        RECT 188.400 157.050 189.450 163.950 ;
        RECT 193.950 160.950 196.050 163.050 ;
        RECT 190.950 157.950 193.050 160.050 ;
        RECT 187.950 154.950 190.050 157.050 ;
        RECT 178.950 151.950 181.050 154.050 ;
        RECT 187.950 151.950 190.050 154.050 ;
        RECT 175.950 130.950 178.050 133.050 ;
        RECT 176.400 127.050 177.450 130.950 ;
        RECT 172.950 125.250 174.750 126.150 ;
        RECT 175.950 124.950 178.050 127.050 ;
        RECT 181.950 126.450 184.050 127.050 ;
        RECT 181.950 125.400 186.450 126.450 ;
        RECT 181.950 124.950 184.050 125.400 ;
        RECT 169.950 121.950 172.050 124.050 ;
        RECT 172.950 121.950 175.050 124.050 ;
        RECT 176.250 122.850 178.050 123.750 ;
        RECT 178.950 122.250 181.050 123.150 ;
        RECT 181.950 122.850 184.050 123.750 ;
        RECT 173.400 118.050 174.450 121.950 ;
        RECT 185.400 121.050 186.450 125.400 ;
        RECT 188.400 124.050 189.450 151.950 ;
        RECT 187.950 121.950 190.050 124.050 ;
        RECT 178.950 118.950 181.050 121.050 ;
        RECT 184.950 118.950 187.050 121.050 ;
        RECT 166.950 115.950 169.050 118.050 ;
        RECT 172.950 115.950 175.050 118.050 ;
        RECT 163.950 112.950 166.050 115.050 ;
        RECT 160.950 103.950 163.050 106.050 ;
        RECT 151.950 100.950 154.050 103.050 ;
        RECT 148.950 55.950 151.050 58.050 ;
        RECT 139.950 53.250 142.050 54.150 ;
        RECT 145.950 53.250 148.050 54.150 ;
        RECT 152.400 52.050 153.450 100.950 ;
        RECT 154.950 97.950 157.050 100.050 ;
        RECT 155.400 97.050 156.450 97.950 ;
        RECT 161.400 97.050 162.450 103.950 ;
        RECT 163.950 100.950 166.050 103.050 ;
        RECT 164.400 97.050 165.450 100.950 ;
        RECT 154.950 94.950 157.050 97.050 ;
        RECT 158.250 95.250 159.750 96.150 ;
        RECT 160.950 94.950 163.050 97.050 ;
        RECT 163.950 94.950 166.050 97.050 ;
        RECT 164.400 94.050 165.450 94.950 ;
        RECT 167.400 94.050 168.450 115.950 ;
        RECT 179.400 115.050 180.450 118.950 ;
        RECT 191.400 118.050 192.450 157.950 ;
        RECT 194.400 142.050 195.450 160.950 ;
        RECT 200.400 142.050 201.450 167.400 ;
        RECT 202.950 166.950 205.050 169.050 ;
        RECT 206.250 167.250 207.750 168.150 ;
        RECT 208.950 166.950 211.050 169.050 ;
        RECT 212.400 166.050 213.450 178.950 ;
        RECT 202.950 164.850 204.750 165.750 ;
        RECT 205.950 163.950 208.050 166.050 ;
        RECT 209.250 164.850 210.750 165.750 ;
        RECT 211.950 163.950 214.050 166.050 ;
        RECT 206.400 148.050 207.450 163.950 ;
        RECT 211.950 161.850 214.050 162.750 ;
        RECT 215.400 151.050 216.450 190.950 ;
        RECT 214.950 148.950 217.050 151.050 ;
        RECT 218.400 148.050 219.450 193.950 ;
        RECT 223.950 184.950 226.050 187.050 ;
        RECT 224.400 172.050 225.450 184.950 ;
        RECT 226.950 175.950 229.050 178.050 ;
        RECT 223.950 169.950 226.050 172.050 ;
        RECT 227.400 169.050 228.450 175.950 ;
        RECT 220.950 166.950 223.050 169.050 ;
        RECT 224.250 167.850 225.750 168.750 ;
        RECT 226.950 166.950 229.050 169.050 ;
        RECT 220.950 164.850 223.050 165.750 ;
        RECT 226.950 164.850 229.050 165.750 ;
        RECT 230.400 159.450 231.450 208.950 ;
        RECT 233.400 205.050 234.450 244.950 ;
        RECT 235.950 238.950 238.050 241.050 ;
        RECT 241.950 238.950 244.050 241.050 ;
        RECT 245.400 240.450 246.450 268.950 ;
        RECT 251.400 247.050 252.450 304.950 ;
        RECT 254.400 289.050 255.450 311.400 ;
        RECT 257.400 301.050 258.450 320.400 ;
        RECT 266.400 319.050 267.450 346.950 ;
        RECT 272.400 343.050 273.450 379.950 ;
        RECT 278.400 352.050 279.450 379.950 ;
        RECT 277.950 349.950 280.050 352.050 ;
        RECT 284.400 349.050 285.450 397.950 ;
        RECT 293.400 382.050 294.450 439.950 ;
        RECT 304.950 430.950 307.050 433.050 ;
        RECT 298.950 424.950 301.050 427.050 ;
        RECT 295.950 421.950 298.050 424.050 ;
        RECT 296.400 400.050 297.450 421.950 ;
        RECT 299.400 406.050 300.450 424.950 ;
        RECT 305.400 421.050 306.450 430.950 ;
        RECT 311.400 426.450 312.450 445.950 ;
        RECT 316.950 439.950 319.050 442.050 ;
        RECT 311.400 425.400 315.450 426.450 ;
        RECT 304.950 418.950 307.050 421.050 ;
        RECT 307.950 419.250 310.050 420.150 ;
        RECT 301.950 415.950 304.050 418.050 ;
        RECT 305.250 416.250 306.750 417.150 ;
        RECT 307.950 415.950 310.050 418.050 ;
        RECT 311.250 416.250 313.050 417.150 ;
        RECT 301.950 413.850 303.750 414.750 ;
        RECT 304.950 412.950 307.050 415.050 ;
        RECT 298.950 403.950 301.050 406.050 ;
        RECT 295.950 397.950 298.050 400.050 ;
        RECT 305.400 397.050 306.450 412.950 ;
        RECT 308.400 409.050 309.450 415.950 ;
        RECT 310.950 414.450 313.050 415.050 ;
        RECT 314.400 414.450 315.450 425.400 ;
        RECT 310.950 413.400 315.450 414.450 ;
        RECT 310.950 412.950 313.050 413.400 ;
        RECT 307.950 406.950 310.050 409.050 ;
        RECT 304.950 394.950 307.050 397.050 ;
        RECT 301.950 391.950 304.050 394.050 ;
        RECT 302.400 385.050 303.450 391.950 ;
        RECT 317.400 391.050 318.450 439.950 ;
        RECT 323.400 433.050 324.450 454.950 ;
        RECT 326.400 451.050 327.450 460.950 ;
        RECT 329.400 460.050 330.450 484.950 ;
        RECT 328.950 457.950 331.050 460.050 ;
        RECT 332.400 456.450 333.450 511.950 ;
        RECT 344.400 505.050 345.450 541.950 ;
        RECT 361.950 538.950 364.050 541.050 ;
        RECT 352.950 532.950 355.050 535.050 ;
        RECT 358.950 532.950 361.050 535.050 ;
        RECT 346.950 526.950 349.050 529.050 ;
        RECT 347.400 522.450 348.450 526.950 ;
        RECT 353.400 526.050 354.450 532.950 ;
        RECT 359.400 532.050 360.450 532.950 ;
        RECT 358.950 529.950 361.050 532.050 ;
        RECT 362.400 529.050 363.450 538.950 ;
        RECT 364.950 535.950 367.050 538.050 ;
        RECT 358.950 527.850 360.750 528.750 ;
        RECT 361.950 526.950 364.050 529.050 ;
        RECT 349.950 524.250 351.750 525.150 ;
        RECT 352.950 523.950 355.050 526.050 ;
        RECT 356.250 524.250 358.050 525.150 ;
        RECT 361.950 524.850 364.050 525.750 ;
        RECT 349.950 522.450 352.050 523.050 ;
        RECT 347.400 521.400 352.050 522.450 ;
        RECT 353.250 521.850 354.750 522.750 ;
        RECT 349.950 520.950 352.050 521.400 ;
        RECT 355.950 520.950 358.050 523.050 ;
        RECT 343.950 502.950 346.050 505.050 ;
        RECT 355.950 488.250 358.050 489.150 ;
        RECT 358.950 487.950 361.050 490.050 ;
        RECT 337.950 484.950 340.050 487.050 ;
        RECT 346.950 485.250 348.750 486.150 ;
        RECT 349.950 484.950 352.050 487.050 ;
        RECT 353.250 485.250 354.750 486.150 ;
        RECT 355.950 484.950 358.050 487.050 ;
        RECT 334.950 482.250 337.050 483.150 ;
        RECT 337.950 482.850 340.050 483.750 ;
        RECT 346.950 481.950 349.050 484.050 ;
        RECT 350.250 482.850 351.750 483.750 ;
        RECT 352.950 483.450 355.050 484.050 ;
        RECT 359.400 483.450 360.450 487.950 ;
        RECT 361.950 484.950 364.050 487.050 ;
        RECT 352.950 482.400 360.450 483.450 ;
        RECT 352.950 481.950 355.050 482.400 ;
        RECT 347.400 481.050 348.450 481.950 ;
        RECT 334.950 478.950 337.050 481.050 ;
        RECT 340.950 478.950 343.050 481.050 ;
        RECT 346.950 478.950 349.050 481.050 ;
        RECT 335.400 478.050 336.450 478.950 ;
        RECT 334.950 475.950 337.050 478.050 ;
        RECT 334.950 472.950 337.050 475.050 ;
        RECT 329.400 455.400 333.450 456.450 ;
        RECT 325.950 448.950 328.050 451.050 ;
        RECT 322.950 430.950 325.050 433.050 ;
        RECT 325.950 427.950 328.050 430.050 ;
        RECT 319.950 416.250 322.050 417.150 ;
        RECT 326.400 415.050 327.450 427.950 ;
        RECT 329.400 418.050 330.450 455.400 ;
        RECT 335.400 454.050 336.450 472.950 ;
        RECT 331.950 452.250 333.750 453.150 ;
        RECT 334.950 451.950 337.050 454.050 ;
        RECT 338.250 452.250 340.050 453.150 ;
        RECT 331.950 448.950 334.050 451.050 ;
        RECT 335.250 449.850 336.750 450.750 ;
        RECT 337.950 448.950 340.050 451.050 ;
        RECT 331.950 445.950 334.050 448.050 ;
        RECT 332.400 421.050 333.450 445.950 ;
        RECT 341.400 439.050 342.450 478.950 ;
        RECT 362.400 472.050 363.450 484.950 ;
        RECT 361.950 469.950 364.050 472.050 ;
        RECT 355.950 466.950 358.050 469.050 ;
        RECT 352.950 457.950 355.050 460.050 ;
        RECT 346.950 454.950 349.050 457.050 ;
        RECT 349.950 454.950 352.050 457.050 ;
        RECT 347.400 454.050 348.450 454.950 ;
        RECT 343.950 452.250 345.750 453.150 ;
        RECT 346.950 451.950 349.050 454.050 ;
        RECT 350.400 451.050 351.450 454.950 ;
        RECT 353.400 454.050 354.450 457.950 ;
        RECT 352.950 451.950 355.050 454.050 ;
        RECT 356.400 451.050 357.450 466.950 ;
        RECT 362.400 460.050 363.450 469.950 ;
        RECT 365.400 463.050 366.450 535.950 ;
        RECT 368.400 535.050 369.450 550.950 ;
        RECT 367.950 532.950 370.050 535.050 ;
        RECT 367.950 527.250 370.050 528.150 ;
        RECT 370.950 526.950 373.050 529.050 ;
        RECT 367.950 523.950 370.050 526.050 ;
        RECT 368.400 517.050 369.450 523.950 ;
        RECT 371.400 519.450 372.450 526.950 ;
        RECT 374.400 523.050 375.450 553.950 ;
        RECT 373.950 520.950 376.050 523.050 ;
        RECT 371.400 518.400 375.450 519.450 ;
        RECT 367.950 514.950 370.050 517.050 ;
        RECT 370.950 484.950 373.050 487.050 ;
        RECT 367.950 482.250 370.050 483.150 ;
        RECT 370.950 482.850 373.050 483.750 ;
        RECT 367.950 478.950 370.050 481.050 ;
        RECT 364.950 460.950 367.050 463.050 ;
        RECT 358.950 457.950 361.050 460.050 ;
        RECT 361.950 457.950 364.050 460.050 ;
        RECT 343.950 448.950 346.050 451.050 ;
        RECT 347.250 449.850 348.750 450.750 ;
        RECT 349.950 448.950 352.050 451.050 ;
        RECT 353.250 449.850 355.050 450.750 ;
        RECT 355.950 448.950 358.050 451.050 ;
        RECT 349.950 446.850 352.050 447.750 ;
        RECT 346.950 439.950 349.050 442.050 ;
        RECT 340.950 436.950 343.050 439.050 ;
        RECT 343.950 436.950 346.050 439.050 ;
        RECT 340.950 427.950 343.050 430.050 ;
        RECT 331.950 418.950 334.050 421.050 ;
        RECT 341.400 418.050 342.450 427.950 ;
        RECT 328.950 415.950 331.050 418.050 ;
        RECT 334.950 417.450 337.050 418.050 ;
        RECT 332.400 416.400 337.050 417.450 ;
        RECT 319.950 412.950 322.050 415.050 ;
        RECT 323.250 413.250 324.750 414.150 ;
        RECT 325.950 412.950 328.050 415.050 ;
        RECT 329.250 413.250 331.050 414.150 ;
        RECT 320.400 412.050 321.450 412.950 ;
        RECT 319.950 409.950 322.050 412.050 ;
        RECT 322.950 409.950 325.050 412.050 ;
        RECT 326.250 410.850 327.750 411.750 ;
        RECT 328.950 411.450 331.050 412.050 ;
        RECT 332.400 411.450 333.450 416.400 ;
        RECT 334.950 415.950 337.050 416.400 ;
        RECT 338.250 416.250 339.750 417.150 ;
        RECT 340.950 415.950 343.050 418.050 ;
        RECT 334.950 413.850 336.750 414.750 ;
        RECT 337.950 412.950 340.050 415.050 ;
        RECT 341.250 413.850 343.050 414.750 ;
        RECT 344.400 412.050 345.450 436.950 ;
        RECT 347.400 424.050 348.450 439.950 ;
        RECT 359.400 433.050 360.450 457.950 ;
        RECT 362.400 457.050 363.450 457.950 ;
        RECT 361.950 454.950 364.050 457.050 ;
        RECT 365.250 455.250 366.750 456.150 ;
        RECT 367.950 454.950 370.050 457.050 ;
        RECT 370.950 454.950 373.050 457.050 ;
        RECT 371.400 454.050 372.450 454.950 ;
        RECT 361.950 452.850 363.750 453.750 ;
        RECT 364.950 451.950 367.050 454.050 ;
        RECT 368.250 452.850 369.750 453.750 ;
        RECT 370.950 451.950 373.050 454.050 ;
        RECT 365.400 448.050 366.450 451.950 ;
        RECT 370.950 449.850 373.050 450.750 ;
        RECT 364.950 445.950 367.050 448.050 ;
        RECT 361.950 433.950 364.050 436.050 ;
        RECT 358.950 430.950 361.050 433.050 ;
        RECT 346.950 421.950 349.050 424.050 ;
        RECT 349.950 419.250 352.050 420.150 ;
        RECT 358.950 418.950 361.050 421.050 ;
        RECT 346.950 416.250 348.750 417.150 ;
        RECT 349.950 415.950 352.050 418.050 ;
        RECT 353.250 416.250 354.750 417.150 ;
        RECT 355.950 415.950 358.050 418.050 ;
        RECT 346.950 412.950 349.050 415.050 ;
        RECT 350.400 412.050 351.450 415.950 ;
        RECT 352.950 412.950 355.050 415.050 ;
        RECT 356.250 413.850 358.050 414.750 ;
        RECT 328.950 410.400 333.450 411.450 ;
        RECT 328.950 409.950 331.050 410.400 ;
        RECT 340.950 409.950 343.050 412.050 ;
        RECT 343.950 409.950 346.050 412.050 ;
        RECT 349.950 409.950 352.050 412.050 ;
        RECT 353.400 411.450 354.450 412.950 ;
        RECT 353.400 410.400 357.450 411.450 ;
        RECT 323.400 409.050 324.450 409.950 ;
        RECT 322.950 406.950 325.050 409.050 ;
        RECT 329.400 406.050 330.450 409.950 ;
        RECT 341.400 409.050 342.450 409.950 ;
        RECT 340.950 406.950 343.050 409.050 ;
        RECT 319.950 403.950 322.050 406.050 ;
        RECT 328.950 403.950 331.050 406.050 ;
        RECT 316.950 388.950 319.050 391.050 ;
        RECT 310.950 385.950 313.050 388.050 ;
        RECT 295.950 382.950 298.050 385.050 ;
        RECT 299.250 383.250 300.750 384.150 ;
        RECT 301.950 382.950 304.050 385.050 ;
        RECT 310.950 383.850 313.050 384.750 ;
        RECT 313.950 383.250 316.050 384.150 ;
        RECT 292.950 379.950 295.050 382.050 ;
        RECT 296.250 380.850 297.750 381.750 ;
        RECT 298.950 379.950 301.050 382.050 ;
        RECT 302.250 380.850 304.050 381.750 ;
        RECT 313.950 379.950 316.050 382.050 ;
        RECT 320.400 381.450 321.450 403.950 ;
        RECT 325.950 391.950 328.050 394.050 ;
        RECT 326.400 385.050 327.450 391.950 ;
        RECT 322.950 383.250 324.750 384.150 ;
        RECT 325.950 382.950 328.050 385.050 ;
        RECT 329.400 382.050 330.450 403.950 ;
        RECT 337.950 388.950 340.050 391.050 ;
        RECT 338.400 388.050 339.450 388.950 ;
        RECT 337.950 385.950 340.050 388.050 ;
        RECT 341.400 385.050 342.450 406.950 ;
        RECT 352.950 397.950 355.050 400.050 ;
        RECT 353.400 385.050 354.450 397.950 ;
        RECT 356.400 388.050 357.450 410.400 ;
        RECT 355.950 385.950 358.050 388.050 ;
        RECT 359.400 385.050 360.450 418.950 ;
        RECT 334.950 384.450 337.050 385.050 ;
        RECT 332.400 383.400 337.050 384.450 ;
        RECT 338.250 383.850 339.750 384.750 ;
        RECT 322.950 381.450 325.050 382.050 ;
        RECT 320.400 380.400 325.050 381.450 ;
        RECT 326.250 380.850 328.050 381.750 ;
        RECT 322.950 379.950 325.050 380.400 ;
        RECT 328.950 379.950 331.050 382.050 ;
        RECT 292.950 377.850 295.050 378.750 ;
        RECT 299.400 373.050 300.450 379.950 ;
        RECT 323.400 379.050 324.450 379.950 ;
        RECT 322.950 376.950 325.050 379.050 ;
        RECT 298.950 370.950 301.050 373.050 ;
        RECT 325.950 367.950 328.050 370.050 ;
        RECT 326.400 367.050 327.450 367.950 ;
        RECT 325.950 364.950 328.050 367.050 ;
        RECT 283.950 346.950 286.050 349.050 ;
        RECT 280.950 343.950 283.050 346.050 ;
        RECT 286.950 345.450 289.050 346.050 ;
        RECT 298.950 345.450 301.050 346.050 ;
        RECT 284.250 344.250 285.750 345.150 ;
        RECT 286.950 344.400 291.450 345.450 ;
        RECT 286.950 343.950 289.050 344.400 ;
        RECT 290.400 343.050 291.450 344.400 ;
        RECT 298.950 344.400 303.450 345.450 ;
        RECT 298.950 343.950 301.050 344.400 ;
        RECT 302.400 343.050 303.450 344.400 ;
        RECT 307.950 343.950 310.050 346.050 ;
        RECT 313.950 343.950 316.050 346.050 ;
        RECT 319.950 344.250 322.050 345.150 ;
        RECT 322.950 343.950 325.050 346.050 ;
        RECT 308.400 343.050 309.450 343.950 ;
        RECT 314.400 343.050 315.450 343.950 ;
        RECT 268.950 341.250 271.050 342.150 ;
        RECT 271.950 340.950 274.050 343.050 ;
        RECT 274.950 341.250 277.050 342.150 ;
        RECT 280.950 341.850 282.750 342.750 ;
        RECT 283.950 340.950 286.050 343.050 ;
        RECT 287.250 341.850 289.050 342.750 ;
        RECT 289.950 340.950 292.050 343.050 ;
        RECT 295.950 341.250 298.050 342.150 ;
        RECT 298.950 341.850 301.050 342.750 ;
        RECT 301.950 340.950 304.050 343.050 ;
        RECT 304.950 341.250 307.050 342.150 ;
        RECT 307.950 340.950 310.050 343.050 ;
        RECT 310.950 341.250 312.750 342.150 ;
        RECT 313.950 340.950 316.050 343.050 ;
        RECT 317.250 341.250 318.750 342.150 ;
        RECT 319.950 340.950 322.050 343.050 ;
        RECT 268.950 337.950 271.050 340.050 ;
        RECT 274.950 337.950 277.050 340.050 ;
        RECT 290.400 339.450 291.450 340.950 ;
        RECT 287.400 338.400 291.450 339.450 ;
        RECT 259.950 316.950 262.050 319.050 ;
        RECT 265.950 316.950 268.050 319.050 ;
        RECT 260.400 313.050 261.450 316.950 ;
        RECT 269.400 316.050 270.450 337.950 ;
        RECT 275.400 337.050 276.450 337.950 ;
        RECT 274.950 334.950 277.050 337.050 ;
        RECT 277.950 331.950 280.050 334.050 ;
        RECT 271.950 316.950 274.050 319.050 ;
        RECT 268.950 313.950 271.050 316.050 ;
        RECT 272.400 313.050 273.450 316.950 ;
        RECT 274.950 313.950 277.050 316.050 ;
        RECT 259.950 310.950 262.050 313.050 ;
        RECT 263.250 311.250 264.750 312.150 ;
        RECT 265.950 310.950 268.050 313.050 ;
        RECT 269.250 311.250 270.750 312.150 ;
        RECT 271.950 310.950 274.050 313.050 ;
        RECT 259.950 308.850 261.750 309.750 ;
        RECT 262.950 307.950 265.050 310.050 ;
        RECT 266.250 308.850 267.750 309.750 ;
        RECT 268.950 307.950 271.050 310.050 ;
        RECT 272.250 308.850 274.050 309.750 ;
        RECT 256.950 298.950 259.050 301.050 ;
        RECT 253.950 286.950 256.050 289.050 ;
        RECT 253.950 283.950 256.050 286.050 ;
        RECT 254.400 277.050 255.450 283.950 ;
        RECT 253.950 274.950 256.050 277.050 ;
        RECT 254.400 262.050 255.450 274.950 ;
        RECT 257.400 273.450 258.450 298.950 ;
        RECT 263.400 295.050 264.450 307.950 ;
        RECT 262.950 292.950 265.050 295.050 ;
        RECT 259.950 273.450 262.050 274.050 ;
        RECT 257.400 272.400 262.050 273.450 ;
        RECT 259.950 271.950 262.050 272.400 ;
        RECT 263.250 272.250 264.750 273.150 ;
        RECT 265.950 271.950 268.050 274.050 ;
        RECT 259.950 269.850 261.750 270.750 ;
        RECT 262.950 268.950 265.050 271.050 ;
        RECT 266.250 269.850 268.050 270.750 ;
        RECT 253.950 259.950 256.050 262.050 ;
        RECT 263.400 247.050 264.450 268.950 ;
        RECT 269.400 259.050 270.450 307.950 ;
        RECT 275.400 277.050 276.450 313.950 ;
        RECT 278.400 307.050 279.450 331.950 ;
        RECT 287.400 316.050 288.450 338.400 ;
        RECT 295.950 337.950 298.050 340.050 ;
        RECT 304.950 339.450 307.050 340.050 ;
        RECT 308.400 339.450 309.450 340.950 ;
        RECT 304.950 338.400 309.450 339.450 ;
        RECT 304.950 337.950 307.050 338.400 ;
        RECT 310.950 337.950 313.050 340.050 ;
        RECT 314.250 338.850 315.750 339.750 ;
        RECT 316.950 337.950 319.050 340.050 ;
        RECT 296.400 331.050 297.450 337.950 ;
        RECT 311.400 336.450 312.450 337.950 ;
        RECT 311.400 335.400 315.450 336.450 ;
        RECT 295.950 328.950 298.050 331.050 ;
        RECT 289.950 319.950 292.050 322.050 ;
        RECT 301.950 319.950 304.050 322.050 ;
        RECT 286.950 313.950 289.050 316.050 ;
        RECT 290.400 313.050 291.450 319.950 ;
        RECT 298.950 313.950 301.050 316.050 ;
        RECT 302.400 313.050 303.450 319.950 ;
        RECT 304.950 316.950 307.050 319.050 ;
        RECT 307.950 316.950 310.050 319.050 ;
        RECT 283.950 312.450 286.050 313.050 ;
        RECT 281.400 311.400 286.050 312.450 ;
        RECT 287.250 311.850 288.750 312.750 ;
        RECT 277.950 304.950 280.050 307.050 ;
        RECT 277.950 283.950 280.050 286.050 ;
        RECT 278.400 283.050 279.450 283.950 ;
        RECT 277.950 280.950 280.050 283.050 ;
        RECT 274.950 274.950 277.050 277.050 ;
        RECT 278.400 274.050 279.450 280.950 ;
        RECT 271.950 271.950 274.050 274.050 ;
        RECT 275.250 272.250 276.750 273.150 ;
        RECT 277.950 271.950 280.050 274.050 ;
        RECT 271.950 269.850 273.750 270.750 ;
        RECT 274.950 268.950 277.050 271.050 ;
        RECT 278.250 269.850 280.050 270.750 ;
        RECT 281.400 268.050 282.450 311.400 ;
        RECT 283.950 310.950 286.050 311.400 ;
        RECT 289.950 310.950 292.050 313.050 ;
        RECT 295.950 312.450 298.050 313.050 ;
        RECT 293.400 311.400 298.050 312.450 ;
        RECT 299.250 311.850 300.750 312.750 ;
        RECT 283.950 308.850 286.050 309.750 ;
        RECT 289.950 308.850 292.050 309.750 ;
        RECT 283.950 304.950 286.050 307.050 ;
        RECT 293.400 306.450 294.450 311.400 ;
        RECT 295.950 310.950 298.050 311.400 ;
        RECT 301.950 310.950 304.050 313.050 ;
        RECT 295.950 308.850 298.050 309.750 ;
        RECT 301.950 308.850 304.050 309.750 ;
        RECT 293.400 305.400 297.450 306.450 ;
        RECT 284.400 271.050 285.450 304.950 ;
        RECT 292.950 277.950 295.050 280.050 ;
        RECT 293.400 274.050 294.450 277.950 ;
        RECT 286.950 271.950 289.050 274.050 ;
        RECT 290.250 272.250 291.750 273.150 ;
        RECT 292.950 271.950 295.050 274.050 ;
        RECT 283.950 268.950 286.050 271.050 ;
        RECT 286.950 269.850 288.750 270.750 ;
        RECT 289.950 268.950 292.050 271.050 ;
        RECT 293.250 269.850 295.050 270.750 ;
        RECT 271.950 265.950 274.050 268.050 ;
        RECT 274.950 265.950 277.050 268.050 ;
        RECT 280.950 265.950 283.050 268.050 ;
        RECT 286.950 265.950 289.050 268.050 ;
        RECT 289.950 265.950 292.050 268.050 ;
        RECT 268.950 256.950 271.050 259.050 ;
        RECT 268.950 247.950 271.050 250.050 ;
        RECT 250.950 244.950 253.050 247.050 ;
        RECT 253.950 244.950 256.050 247.050 ;
        RECT 262.950 244.950 265.050 247.050 ;
        RECT 245.400 239.400 249.450 240.450 ;
        RECT 232.950 202.950 235.050 205.050 ;
        RECT 236.400 199.050 237.450 238.950 ;
        RECT 242.400 238.050 243.450 238.950 ;
        RECT 238.950 236.250 240.750 237.150 ;
        RECT 241.950 235.950 244.050 238.050 ;
        RECT 245.250 236.250 247.050 237.150 ;
        RECT 238.950 232.950 241.050 235.050 ;
        RECT 242.250 233.850 243.750 234.750 ;
        RECT 244.950 232.950 247.050 235.050 ;
        RECT 239.400 232.050 240.450 232.950 ;
        RECT 245.400 232.050 246.450 232.950 ;
        RECT 238.950 229.950 241.050 232.050 ;
        RECT 244.950 229.950 247.050 232.050 ;
        RECT 248.400 205.050 249.450 239.400 ;
        RECT 250.950 238.950 253.050 241.050 ;
        RECT 238.950 202.950 241.050 205.050 ;
        RECT 244.950 203.250 247.050 204.150 ;
        RECT 247.950 202.950 250.050 205.050 ;
        RECT 251.400 204.450 252.450 238.950 ;
        RECT 254.400 235.050 255.450 244.950 ;
        RECT 256.950 241.950 259.050 244.050 ;
        RECT 257.400 238.050 258.450 241.950 ;
        RECT 259.950 238.950 262.050 241.050 ;
        RECT 263.250 239.250 264.750 240.150 ;
        RECT 265.950 238.950 268.050 241.050 ;
        RECT 256.950 235.950 259.050 238.050 ;
        RECT 260.250 236.850 261.750 237.750 ;
        RECT 262.950 235.950 265.050 238.050 ;
        RECT 266.250 236.850 268.050 237.750 ;
        RECT 263.400 235.050 264.450 235.950 ;
        RECT 253.950 232.950 256.050 235.050 ;
        RECT 256.950 233.850 259.050 234.750 ;
        RECT 262.950 232.950 265.050 235.050 ;
        RECT 269.400 211.050 270.450 247.950 ;
        RECT 272.400 244.050 273.450 265.950 ;
        RECT 275.400 244.050 276.450 265.950 ;
        RECT 280.950 259.950 283.050 262.050 ;
        RECT 271.950 241.950 274.050 244.050 ;
        RECT 274.950 241.950 277.050 244.050 ;
        RECT 277.950 241.950 280.050 244.050 ;
        RECT 271.950 239.850 274.050 240.750 ;
        RECT 274.950 239.250 277.050 240.150 ;
        RECT 271.950 235.950 274.050 238.050 ;
        RECT 274.950 235.950 277.050 238.050 ;
        RECT 268.950 208.950 271.050 211.050 ;
        RECT 256.950 205.950 259.050 208.050 ;
        RECT 251.400 203.400 255.450 204.450 ;
        RECT 239.400 202.050 240.450 202.950 ;
        RECT 238.950 199.950 241.050 202.050 ;
        RECT 241.950 200.250 243.750 201.150 ;
        RECT 244.950 199.950 247.050 202.050 ;
        RECT 248.250 200.250 249.750 201.150 ;
        RECT 250.950 199.950 253.050 202.050 ;
        RECT 232.950 196.950 235.050 199.050 ;
        RECT 235.950 196.950 238.050 199.050 ;
        RECT 238.950 196.950 241.050 199.050 ;
        RECT 241.950 196.950 244.050 199.050 ;
        RECT 232.950 194.850 235.050 195.750 ;
        RECT 235.950 194.250 238.050 195.150 ;
        RECT 235.950 192.450 238.050 193.050 ;
        RECT 239.400 192.450 240.450 196.950 ;
        RECT 242.400 196.050 243.450 196.950 ;
        RECT 245.400 196.050 246.450 199.950 ;
        RECT 247.950 196.950 250.050 199.050 ;
        RECT 251.250 197.850 253.050 198.750 ;
        RECT 254.400 196.050 255.450 203.400 ;
        RECT 241.950 193.950 244.050 196.050 ;
        RECT 244.950 193.950 247.050 196.050 ;
        RECT 253.950 193.950 256.050 196.050 ;
        RECT 235.950 191.400 240.450 192.450 ;
        RECT 235.950 190.950 238.050 191.400 ;
        RECT 232.950 175.950 235.050 178.050 ;
        RECT 233.400 172.050 234.450 175.950 ;
        RECT 244.950 172.950 247.050 175.050 ;
        RECT 250.950 172.950 253.050 175.050 ;
        RECT 232.950 169.950 235.050 172.050 ;
        RECT 238.950 169.950 241.050 172.050 ;
        RECT 232.950 167.850 235.050 168.750 ;
        RECT 235.950 167.250 238.050 168.150 ;
        RECT 235.950 163.950 238.050 166.050 ;
        RECT 236.400 163.050 237.450 163.950 ;
        RECT 235.950 160.950 238.050 163.050 ;
        RECT 239.400 159.450 240.450 169.950 ;
        RECT 241.950 166.950 244.050 169.050 ;
        RECT 230.400 158.400 234.450 159.450 ;
        RECT 229.950 148.950 232.050 151.050 ;
        RECT 205.950 145.950 208.050 148.050 ;
        RECT 217.950 145.950 220.050 148.050 ;
        RECT 193.950 139.950 196.050 142.050 ;
        RECT 199.950 139.950 202.050 142.050 ;
        RECT 194.400 130.050 195.450 139.950 ;
        RECT 205.950 133.950 208.050 136.050 ;
        RECT 199.950 131.250 202.050 132.150 ;
        RECT 193.950 127.950 196.050 130.050 ;
        RECT 197.250 128.250 198.750 129.150 ;
        RECT 199.950 127.950 202.050 130.050 ;
        RECT 203.250 128.250 205.050 129.150 ;
        RECT 193.950 125.850 195.750 126.750 ;
        RECT 196.950 124.950 199.050 127.050 ;
        RECT 197.400 121.050 198.450 124.950 ;
        RECT 200.400 123.450 201.450 127.950 ;
        RECT 202.950 124.950 205.050 127.050 ;
        RECT 200.400 122.400 204.450 123.450 ;
        RECT 196.950 118.950 199.050 121.050 ;
        RECT 190.950 115.950 193.050 118.050 ;
        RECT 178.950 112.950 181.050 115.050 ;
        RECT 199.950 112.950 202.050 115.050 ;
        RECT 184.950 106.950 187.050 109.050 ;
        RECT 185.400 100.050 186.450 106.950 ;
        RECT 184.950 97.950 187.050 100.050 ;
        RECT 175.950 94.950 178.050 97.050 ;
        RECT 179.250 95.250 181.050 96.150 ;
        RECT 185.400 94.050 186.450 97.950 ;
        RECT 200.400 97.050 201.450 112.950 ;
        RECT 203.400 109.050 204.450 122.400 ;
        RECT 202.950 106.950 205.050 109.050 ;
        RECT 190.950 96.450 193.050 97.050 ;
        RECT 193.950 96.450 196.050 97.050 ;
        RECT 190.950 95.400 196.050 96.450 ;
        RECT 190.950 94.950 193.050 95.400 ;
        RECT 193.950 94.950 196.050 95.400 ;
        RECT 197.250 95.250 198.750 96.150 ;
        RECT 199.950 94.950 202.050 97.050 ;
        RECT 154.950 92.850 156.750 93.750 ;
        RECT 157.950 91.950 160.050 94.050 ;
        RECT 161.250 92.850 162.750 93.750 ;
        RECT 163.950 91.950 166.050 94.050 ;
        RECT 166.950 91.950 169.050 94.050 ;
        RECT 175.950 92.850 177.750 93.750 ;
        RECT 178.950 91.950 181.050 94.050 ;
        RECT 184.950 91.950 187.050 94.050 ;
        RECT 190.950 93.450 193.050 94.050 ;
        RECT 188.400 92.400 193.050 93.450 ;
        RECT 194.250 92.850 195.750 93.750 ;
        RECT 154.950 88.950 157.050 91.050 ;
        RECT 163.950 89.850 166.050 90.750 ;
        RECT 179.400 90.450 180.450 91.950 ;
        RECT 176.400 89.400 180.450 90.450 ;
        RECT 155.400 58.050 156.450 88.950 ;
        RECT 160.950 59.250 163.050 60.150 ;
        RECT 154.950 55.950 157.050 58.050 ;
        RECT 158.250 56.250 159.750 57.150 ;
        RECT 160.950 55.950 163.050 58.050 ;
        RECT 164.250 56.250 166.050 57.150 ;
        RECT 176.400 55.050 177.450 89.400 ;
        RECT 188.400 67.050 189.450 92.400 ;
        RECT 190.950 91.950 193.050 92.400 ;
        RECT 196.950 91.950 199.050 94.050 ;
        RECT 200.250 92.850 202.050 93.750 ;
        RECT 190.950 89.850 193.050 90.750 ;
        RECT 190.950 85.950 193.050 88.050 ;
        RECT 191.400 85.050 192.450 85.950 ;
        RECT 190.950 82.950 193.050 85.050 ;
        RECT 178.950 64.950 181.050 67.050 ;
        RECT 187.950 64.950 190.050 67.050 ;
        RECT 154.950 53.850 156.750 54.750 ;
        RECT 157.950 52.950 160.050 55.050 ;
        RECT 163.950 52.950 166.050 55.050 ;
        RECT 169.950 54.450 172.050 55.050 ;
        RECT 169.950 53.400 174.450 54.450 ;
        RECT 169.950 52.950 172.050 53.400 ;
        RECT 158.400 52.050 159.450 52.950 ;
        RECT 139.950 49.950 142.050 52.050 ;
        RECT 143.250 50.250 144.750 51.150 ;
        RECT 145.950 49.950 148.050 52.050 ;
        RECT 151.950 49.950 154.050 52.050 ;
        RECT 157.950 49.950 160.050 52.050 ;
        RECT 136.950 46.950 139.050 49.050 ;
        RECT 140.400 46.050 141.450 49.950 ;
        RECT 164.400 49.050 165.450 52.950 ;
        RECT 173.400 52.050 174.450 53.400 ;
        RECT 175.950 52.950 178.050 55.050 ;
        RECT 179.400 52.050 180.450 64.950 ;
        RECT 203.400 55.050 204.450 106.950 ;
        RECT 206.400 94.050 207.450 133.950 ;
        RECT 223.950 131.250 226.050 132.150 ;
        RECT 230.400 130.050 231.450 148.950 ;
        RECT 211.950 129.450 214.050 130.050 ;
        RECT 209.400 128.400 214.050 129.450 ;
        RECT 209.400 121.050 210.450 128.400 ;
        RECT 211.950 127.950 214.050 128.400 ;
        RECT 215.250 128.250 216.750 129.150 ;
        RECT 217.950 127.950 220.050 130.050 ;
        RECT 220.950 128.250 222.750 129.150 ;
        RECT 223.950 127.950 226.050 130.050 ;
        RECT 227.250 128.250 228.750 129.150 ;
        RECT 229.950 127.950 232.050 130.050 ;
        RECT 211.950 125.850 213.750 126.750 ;
        RECT 214.950 124.950 217.050 127.050 ;
        RECT 218.250 125.850 220.050 126.750 ;
        RECT 220.950 124.950 223.050 127.050 ;
        RECT 215.400 124.050 216.450 124.950 ;
        RECT 224.400 124.050 225.450 127.950 ;
        RECT 226.950 124.950 229.050 127.050 ;
        RECT 230.250 125.850 232.050 126.750 ;
        RECT 214.950 121.950 217.050 124.050 ;
        RECT 217.950 121.950 220.050 124.050 ;
        RECT 223.950 121.950 226.050 124.050 ;
        RECT 208.950 118.950 211.050 121.050 ;
        RECT 211.950 97.950 214.050 100.050 ;
        RECT 218.400 97.050 219.450 121.950 ;
        RECT 227.400 106.050 228.450 124.950 ;
        RECT 226.950 103.950 229.050 106.050 ;
        RECT 233.400 103.050 234.450 158.400 ;
        RECT 236.400 158.400 240.450 159.450 ;
        RECT 236.400 112.050 237.450 158.400 ;
        RECT 242.400 133.050 243.450 166.950 ;
        RECT 245.400 162.450 246.450 172.950 ;
        RECT 251.400 166.050 252.450 172.950 ;
        RECT 247.950 164.250 249.750 165.150 ;
        RECT 250.950 163.950 253.050 166.050 ;
        RECT 254.250 164.250 256.050 165.150 ;
        RECT 247.950 162.450 250.050 163.050 ;
        RECT 245.400 161.400 250.050 162.450 ;
        RECT 251.250 161.850 252.750 162.750 ;
        RECT 247.950 160.950 250.050 161.400 ;
        RECT 253.950 160.950 256.050 163.050 ;
        RECT 247.950 151.950 250.050 154.050 ;
        RECT 241.950 130.950 244.050 133.050 ;
        RECT 248.400 130.050 249.450 151.950 ;
        RECT 257.400 133.050 258.450 205.950 ;
        RECT 259.950 199.950 262.050 202.050 ;
        RECT 260.400 195.450 261.450 199.950 ;
        RECT 262.950 197.250 265.050 198.150 ;
        RECT 268.950 197.250 271.050 198.150 ;
        RECT 262.950 195.450 265.050 196.050 ;
        RECT 260.400 194.400 265.050 195.450 ;
        RECT 262.950 193.950 265.050 194.400 ;
        RECT 266.250 194.250 267.750 195.150 ;
        RECT 268.950 193.950 271.050 196.050 ;
        RECT 265.950 190.950 268.050 193.050 ;
        RECT 266.400 181.050 267.450 190.950 ;
        RECT 265.950 178.950 268.050 181.050 ;
        RECT 272.400 178.050 273.450 235.950 ;
        RECT 275.400 232.050 276.450 235.950 ;
        RECT 274.950 229.950 277.050 232.050 ;
        RECT 274.950 220.950 277.050 223.050 ;
        RECT 265.950 175.950 268.050 178.050 ;
        RECT 271.950 175.950 274.050 178.050 ;
        RECT 266.400 172.050 267.450 175.950 ;
        RECT 259.950 169.950 262.050 172.050 ;
        RECT 265.950 169.950 268.050 172.050 ;
        RECT 260.400 136.050 261.450 169.950 ;
        RECT 262.950 166.950 265.050 169.050 ;
        RECT 266.250 167.850 267.750 168.750 ;
        RECT 268.950 166.950 271.050 169.050 ;
        RECT 275.400 168.450 276.450 220.950 ;
        RECT 278.400 220.050 279.450 241.950 ;
        RECT 281.400 238.050 282.450 259.950 ;
        RECT 283.950 238.950 286.050 241.050 ;
        RECT 287.400 240.450 288.450 265.950 ;
        RECT 290.400 244.050 291.450 265.950 ;
        RECT 289.950 241.950 292.050 244.050 ;
        RECT 287.400 239.400 291.450 240.450 ;
        RECT 280.950 235.950 283.050 238.050 ;
        RECT 280.950 232.950 283.050 235.050 ;
        RECT 284.400 234.450 285.450 238.950 ;
        RECT 290.400 238.050 291.450 239.400 ;
        RECT 286.950 236.250 288.750 237.150 ;
        RECT 289.950 235.950 292.050 238.050 ;
        RECT 293.250 236.250 295.050 237.150 ;
        RECT 286.950 234.450 289.050 235.050 ;
        RECT 284.400 233.400 289.050 234.450 ;
        RECT 290.250 233.850 291.750 234.750 ;
        RECT 292.950 234.450 295.050 235.050 ;
        RECT 296.400 234.450 297.450 305.400 ;
        RECT 305.400 304.050 306.450 316.950 ;
        RECT 304.950 301.950 307.050 304.050 ;
        RECT 304.950 295.950 307.050 298.050 ;
        RECT 301.950 280.950 304.050 283.050 ;
        RECT 298.950 277.950 301.050 280.050 ;
        RECT 299.400 271.050 300.450 277.950 ;
        RECT 302.400 271.050 303.450 280.950 ;
        RECT 305.400 271.050 306.450 295.950 ;
        RECT 308.400 273.450 309.450 316.950 ;
        RECT 310.950 313.950 313.050 316.050 ;
        RECT 311.400 310.050 312.450 313.950 ;
        RECT 314.400 313.050 315.450 335.400 ;
        RECT 317.400 328.050 318.450 337.950 ;
        RECT 316.950 325.950 319.050 328.050 ;
        RECT 320.400 325.050 321.450 340.950 ;
        RECT 323.400 328.050 324.450 343.950 ;
        RECT 322.950 325.950 325.050 328.050 ;
        RECT 319.950 322.950 322.050 325.050 ;
        RECT 326.400 319.050 327.450 364.950 ;
        RECT 332.400 358.050 333.450 383.400 ;
        RECT 334.950 382.950 337.050 383.400 ;
        RECT 340.950 382.950 343.050 385.050 ;
        RECT 352.950 382.950 355.050 385.050 ;
        RECT 356.250 383.850 357.750 384.750 ;
        RECT 358.950 382.950 361.050 385.050 ;
        RECT 362.400 382.050 363.450 433.950 ;
        RECT 364.950 427.950 367.050 430.050 ;
        RECT 365.400 418.050 366.450 427.950 ;
        RECT 374.400 427.050 375.450 518.400 ;
        RECT 377.400 466.050 378.450 556.950 ;
        RECT 380.400 556.050 381.450 556.950 ;
        RECT 379.950 553.950 382.050 556.050 ;
        RECT 386.400 535.050 387.450 559.950 ;
        RECT 389.400 538.050 390.450 601.950 ;
        RECT 392.400 562.050 393.450 640.950 ;
        RECT 395.400 562.050 396.450 698.400 ;
        RECT 401.400 696.450 402.450 700.950 ;
        RECT 403.950 698.850 406.050 699.750 ;
        RECT 406.950 698.250 409.050 699.150 ;
        RECT 409.950 698.850 411.750 699.750 ;
        RECT 412.950 697.950 415.050 700.050 ;
        RECT 398.400 695.400 402.450 696.450 ;
        RECT 398.400 673.050 399.450 695.400 ;
        RECT 406.950 694.950 409.050 697.050 ;
        RECT 407.400 691.050 408.450 694.950 ;
        RECT 416.400 694.050 417.450 700.950 ;
        RECT 424.950 697.950 427.050 700.050 ;
        RECT 428.250 698.850 429.750 699.750 ;
        RECT 430.950 697.950 433.050 700.050 ;
        RECT 425.400 694.050 426.450 697.950 ;
        RECT 415.950 691.950 418.050 694.050 ;
        RECT 424.950 691.950 427.050 694.050 ;
        RECT 431.400 691.050 432.450 697.950 ;
        RECT 406.950 688.950 409.050 691.050 ;
        RECT 430.950 688.950 433.050 691.050 ;
        RECT 415.950 685.950 418.050 688.050 ;
        RECT 412.950 682.950 415.050 685.050 ;
        RECT 409.950 679.950 412.050 682.050 ;
        RECT 403.950 676.950 406.050 679.050 ;
        RECT 404.400 676.050 405.450 676.950 ;
        RECT 403.950 673.950 406.050 676.050 ;
        RECT 397.950 670.950 400.050 673.050 ;
        RECT 401.250 671.250 403.050 672.150 ;
        RECT 403.950 671.850 406.050 672.750 ;
        RECT 406.950 671.250 409.050 672.150 ;
        RECT 397.950 668.850 399.750 669.750 ;
        RECT 400.950 667.950 403.050 670.050 ;
        RECT 406.950 667.950 409.050 670.050 ;
        RECT 401.400 637.050 402.450 667.950 ;
        RECT 400.950 634.950 403.050 637.050 ;
        RECT 406.950 634.950 409.050 637.050 ;
        RECT 407.400 634.050 408.450 634.950 ;
        RECT 400.950 633.450 403.050 634.050 ;
        RECT 398.400 632.400 403.050 633.450 ;
        RECT 398.400 604.050 399.450 632.400 ;
        RECT 400.950 631.950 403.050 632.400 ;
        RECT 404.250 632.250 405.750 633.150 ;
        RECT 406.950 631.950 409.050 634.050 ;
        RECT 400.950 629.850 402.750 630.750 ;
        RECT 403.950 628.950 406.050 631.050 ;
        RECT 407.250 629.850 409.050 630.750 ;
        RECT 404.400 628.050 405.450 628.950 ;
        RECT 403.950 625.950 406.050 628.050 ;
        RECT 410.400 627.450 411.450 679.950 ;
        RECT 413.400 670.050 414.450 682.950 ;
        RECT 412.950 667.950 415.050 670.050 ;
        RECT 412.950 634.950 415.050 637.050 ;
        RECT 413.400 628.050 414.450 634.950 ;
        RECT 416.400 631.050 417.450 685.950 ;
        RECT 431.400 679.050 432.450 688.950 ;
        RECT 434.400 688.050 435.450 709.950 ;
        RECT 449.400 709.050 450.450 746.400 ;
        RECT 452.400 715.050 453.450 748.950 ;
        RECT 455.400 745.050 456.450 752.400 ;
        RECT 458.400 745.050 459.450 766.950 ;
        RECT 467.400 763.050 468.450 815.400 ;
        RECT 469.950 814.950 472.050 815.400 ;
        RECT 473.250 815.250 475.050 816.150 ;
        RECT 475.950 815.850 478.050 816.750 ;
        RECT 478.950 815.250 481.050 816.150 ;
        RECT 484.950 814.950 487.050 817.050 ;
        RECT 502.950 814.950 505.050 817.050 ;
        RECT 469.950 812.850 471.750 813.750 ;
        RECT 472.950 811.950 475.050 814.050 ;
        RECT 478.950 811.950 481.050 814.050 ;
        RECT 473.400 811.050 474.450 811.950 ;
        RECT 472.950 808.950 475.050 811.050 ;
        RECT 479.400 808.050 480.450 811.950 ;
        RECT 485.400 810.450 486.450 814.950 ;
        RECT 487.950 812.250 489.750 813.150 ;
        RECT 490.950 811.950 493.050 814.050 ;
        RECT 494.250 812.250 496.050 813.150 ;
        RECT 502.950 812.850 505.050 813.750 ;
        RECT 505.950 812.250 508.050 813.150 ;
        RECT 487.950 810.450 490.050 811.050 ;
        RECT 485.400 809.400 490.050 810.450 ;
        RECT 491.250 809.850 492.750 810.750 ;
        RECT 487.950 808.950 490.050 809.400 ;
        RECT 493.950 808.950 496.050 811.050 ;
        RECT 505.950 808.950 508.050 811.050 ;
        RECT 494.400 808.050 495.450 808.950 ;
        RECT 478.950 805.950 481.050 808.050 ;
        RECT 493.950 805.950 496.050 808.050 ;
        RECT 494.400 805.050 495.450 805.950 ;
        RECT 493.950 802.950 496.050 805.050 ;
        RECT 509.400 781.050 510.450 820.950 ;
        RECT 511.950 817.950 514.050 820.050 ;
        RECT 512.400 817.050 513.450 817.950 ;
        RECT 524.400 817.050 525.450 820.950 ;
        RECT 788.400 820.050 789.450 820.950 ;
        RECT 538.950 817.950 541.050 820.050 ;
        RECT 559.950 817.950 562.050 820.050 ;
        RECT 577.950 819.450 580.050 820.050 ;
        RECT 595.950 819.450 598.050 820.050 ;
        RECT 577.950 818.400 582.450 819.450 ;
        RECT 577.950 817.950 580.050 818.400 ;
        RECT 511.950 814.950 514.050 817.050 ;
        RECT 517.950 816.450 520.050 817.050 ;
        RECT 515.400 815.400 520.050 816.450 ;
        RECT 511.950 812.850 514.050 813.750 ;
        RECT 515.400 784.050 516.450 815.400 ;
        RECT 517.950 814.950 520.050 815.400 ;
        RECT 521.250 815.250 522.750 816.150 ;
        RECT 523.950 814.950 526.050 817.050 ;
        RECT 529.950 816.450 532.050 817.050 ;
        RECT 527.250 815.250 528.750 816.150 ;
        RECT 529.950 815.400 534.450 816.450 ;
        RECT 529.950 814.950 532.050 815.400 ;
        RECT 517.950 812.850 519.750 813.750 ;
        RECT 520.950 811.950 523.050 814.050 ;
        RECT 524.250 812.850 525.750 813.750 ;
        RECT 526.950 811.950 529.050 814.050 ;
        RECT 530.250 812.850 532.050 813.750 ;
        RECT 517.950 808.950 520.050 811.050 ;
        RECT 514.950 781.950 517.050 784.050 ;
        RECT 508.950 778.950 511.050 781.050 ;
        RECT 508.950 775.950 511.050 778.050 ;
        RECT 509.400 775.050 510.450 775.950 ;
        RECT 469.950 773.250 472.050 774.150 ;
        RECT 475.950 773.250 478.050 774.150 ;
        RECT 484.950 772.950 487.050 775.050 ;
        RECT 499.950 773.250 501.750 774.150 ;
        RECT 502.950 772.950 505.050 775.050 ;
        RECT 506.250 773.250 507.750 774.150 ;
        RECT 508.950 772.950 511.050 775.050 ;
        RECT 512.250 773.250 514.050 774.150 ;
        RECT 469.950 769.950 472.050 772.050 ;
        RECT 473.250 770.250 474.750 771.150 ;
        RECT 475.950 769.950 478.050 772.050 ;
        RECT 481.950 770.250 484.050 771.150 ;
        RECT 484.950 770.850 487.050 771.750 ;
        RECT 499.950 769.950 502.050 772.050 ;
        RECT 503.250 770.850 504.750 771.750 ;
        RECT 505.950 769.950 508.050 772.050 ;
        RECT 509.250 770.850 510.750 771.750 ;
        RECT 511.950 771.450 514.050 772.050 ;
        RECT 515.400 771.450 516.450 781.950 ;
        RECT 511.950 770.400 516.450 771.450 ;
        RECT 511.950 769.950 514.050 770.400 ;
        RECT 470.400 765.450 471.450 769.950 ;
        RECT 472.950 766.950 475.050 769.050 ;
        RECT 470.400 764.400 474.450 765.450 ;
        RECT 466.950 760.950 469.050 763.050 ;
        RECT 466.950 757.950 469.050 760.050 ;
        RECT 463.950 748.950 466.050 751.050 ;
        RECT 464.400 745.050 465.450 748.950 ;
        RECT 467.400 748.050 468.450 757.950 ;
        RECT 466.950 745.950 469.050 748.050 ;
        RECT 454.950 742.950 457.050 745.050 ;
        RECT 457.950 742.950 460.050 745.050 ;
        RECT 461.250 743.250 462.750 744.150 ;
        RECT 463.950 742.950 466.050 745.050 ;
        RECT 466.950 743.850 469.050 744.750 ;
        RECT 469.950 743.250 472.050 744.150 ;
        RECT 455.400 742.050 456.450 742.950 ;
        RECT 454.950 739.950 457.050 742.050 ;
        RECT 458.250 740.850 459.750 741.750 ;
        RECT 460.950 739.950 463.050 742.050 ;
        RECT 464.250 740.850 466.050 741.750 ;
        RECT 469.950 739.950 472.050 742.050 ;
        RECT 454.950 737.850 457.050 738.750 ;
        RECT 451.950 712.950 454.050 715.050 ;
        RECT 452.400 712.050 453.450 712.950 ;
        RECT 451.950 709.950 454.050 712.050 ;
        RECT 436.950 706.950 439.050 709.050 ;
        RECT 445.950 706.950 448.050 709.050 ;
        RECT 448.950 706.950 451.050 709.050 ;
        RECT 437.400 706.050 438.450 706.950 ;
        RECT 436.950 703.950 439.050 706.050 ;
        RECT 440.250 704.250 441.750 705.150 ;
        RECT 442.950 703.950 445.050 706.050 ;
        RECT 436.950 701.850 438.750 702.750 ;
        RECT 439.950 700.950 442.050 703.050 ;
        RECT 443.250 701.850 445.050 702.750 ;
        RECT 436.950 697.950 439.050 700.050 ;
        RECT 433.950 685.950 436.050 688.050 ;
        RECT 430.950 676.950 433.050 679.050 ;
        RECT 421.950 673.950 424.050 676.050 ;
        RECT 437.400 673.050 438.450 697.950 ;
        RECT 440.400 685.050 441.450 700.950 ;
        RECT 446.400 700.050 447.450 706.950 ;
        RECT 452.400 706.050 453.450 709.950 ;
        RECT 461.400 706.050 462.450 739.950 ;
        RECT 470.400 736.050 471.450 739.950 ;
        RECT 469.950 733.950 472.050 736.050 ;
        RECT 463.950 706.950 466.050 709.050 ;
        RECT 451.950 703.950 454.050 706.050 ;
        RECT 455.250 704.250 456.750 705.150 ;
        RECT 457.950 703.950 460.050 706.050 ;
        RECT 460.950 703.950 463.050 706.050 ;
        RECT 451.950 701.850 453.750 702.750 ;
        RECT 454.950 700.950 457.050 703.050 ;
        RECT 458.250 701.850 460.050 702.750 ;
        RECT 442.950 697.950 445.050 700.050 ;
        RECT 445.950 697.950 448.050 700.050 ;
        RECT 439.950 682.950 442.050 685.050 ;
        RECT 439.950 676.950 442.050 679.050 ;
        RECT 418.950 671.250 421.050 672.150 ;
        RECT 421.950 671.850 424.050 672.750 ;
        RECT 427.950 670.950 430.050 673.050 ;
        RECT 433.950 670.950 436.050 673.050 ;
        RECT 436.950 670.950 439.050 673.050 ;
        RECT 418.950 667.950 421.050 670.050 ;
        RECT 419.400 667.050 420.450 667.950 ;
        RECT 418.950 664.950 421.050 667.050 ;
        RECT 421.950 637.950 424.050 640.050 ;
        RECT 415.950 628.950 418.050 631.050 ;
        RECT 407.400 626.400 411.450 627.450 ;
        RECT 407.400 607.050 408.450 626.400 ;
        RECT 412.950 625.950 415.050 628.050 ;
        RECT 415.950 626.850 418.050 627.750 ;
        RECT 418.950 626.250 421.050 627.150 ;
        RECT 418.950 624.450 421.050 625.050 ;
        RECT 422.400 624.450 423.450 637.950 ;
        RECT 424.950 634.950 427.050 637.050 ;
        RECT 418.950 623.400 423.450 624.450 ;
        RECT 418.950 622.950 421.050 623.400 ;
        RECT 415.950 616.950 418.050 619.050 ;
        RECT 409.950 610.950 412.050 613.050 ;
        RECT 406.950 604.950 409.050 607.050 ;
        RECT 397.950 601.950 400.050 604.050 ;
        RECT 400.950 603.450 403.050 604.050 ;
        RECT 400.950 602.400 405.450 603.450 ;
        RECT 400.950 601.950 403.050 602.400 ;
        RECT 397.950 599.250 400.050 600.150 ;
        RECT 400.950 599.850 403.050 600.750 ;
        RECT 397.950 595.950 400.050 598.050 ;
        RECT 404.400 592.050 405.450 602.400 ;
        RECT 410.400 598.050 411.450 610.950 ;
        RECT 412.950 598.950 415.050 601.050 ;
        RECT 406.950 596.250 408.750 597.150 ;
        RECT 409.950 595.950 412.050 598.050 ;
        RECT 413.400 595.050 414.450 598.950 ;
        RECT 416.400 598.050 417.450 616.950 ;
        RECT 425.400 604.050 426.450 634.950 ;
        RECT 428.400 634.050 429.450 670.950 ;
        RECT 433.950 668.850 436.050 669.750 ;
        RECT 436.950 668.250 439.050 669.150 ;
        RECT 436.950 666.450 439.050 667.050 ;
        RECT 440.400 666.450 441.450 676.950 ;
        RECT 443.400 673.050 444.450 697.950 ;
        RECT 446.400 679.050 447.450 697.950 ;
        RECT 448.950 691.950 451.050 694.050 ;
        RECT 445.950 676.950 448.050 679.050 ;
        RECT 442.950 670.950 445.050 673.050 ;
        RECT 445.950 670.950 448.050 673.050 ;
        RECT 442.950 668.850 445.050 669.750 ;
        RECT 436.950 665.400 441.450 666.450 ;
        RECT 436.950 664.950 439.050 665.400 ;
        RECT 446.400 637.050 447.450 670.950 ;
        RECT 439.950 634.950 442.050 637.050 ;
        RECT 445.950 634.950 448.050 637.050 ;
        RECT 427.950 631.950 430.050 634.050 ;
        RECT 433.950 633.450 436.050 634.050 ;
        RECT 431.250 632.250 432.750 633.150 ;
        RECT 433.950 632.400 438.450 633.450 ;
        RECT 433.950 631.950 436.050 632.400 ;
        RECT 427.950 629.850 429.750 630.750 ;
        RECT 430.950 628.950 433.050 631.050 ;
        RECT 434.250 629.850 436.050 630.750 ;
        RECT 427.950 625.950 430.050 628.050 ;
        RECT 424.950 601.950 427.050 604.050 ;
        RECT 428.400 601.050 429.450 625.950 ;
        RECT 431.400 625.050 432.450 628.950 ;
        RECT 437.400 628.050 438.450 632.400 ;
        RECT 436.950 625.950 439.050 628.050 ;
        RECT 430.950 622.950 433.050 625.050 ;
        RECT 430.950 601.950 433.050 604.050 ;
        RECT 418.950 598.950 421.050 601.050 ;
        RECT 421.950 598.950 424.050 601.050 ;
        RECT 425.250 599.250 426.750 600.150 ;
        RECT 427.950 598.950 430.050 601.050 ;
        RECT 415.950 595.950 418.050 598.050 ;
        RECT 406.950 592.950 409.050 595.050 ;
        RECT 410.250 593.850 411.750 594.750 ;
        RECT 412.950 592.950 415.050 595.050 ;
        RECT 416.250 593.850 418.050 594.750 ;
        RECT 403.950 589.950 406.050 592.050 ;
        RECT 412.950 590.850 415.050 591.750 ;
        RECT 419.400 586.050 420.450 598.950 ;
        RECT 431.400 598.050 432.450 601.950 ;
        RECT 433.950 598.950 436.050 601.050 ;
        RECT 421.950 596.850 423.750 597.750 ;
        RECT 424.950 595.950 427.050 598.050 ;
        RECT 428.250 596.850 429.750 597.750 ;
        RECT 430.950 595.950 433.050 598.050 ;
        RECT 425.400 595.050 426.450 595.950 ;
        RECT 424.950 592.950 427.050 595.050 ;
        RECT 430.950 593.850 433.050 594.750 ;
        RECT 425.400 592.050 426.450 592.950 ;
        RECT 424.950 589.950 427.050 592.050 ;
        RECT 418.950 583.950 421.050 586.050 ;
        RECT 434.400 583.050 435.450 598.950 ;
        RECT 433.950 580.950 436.050 583.050 ;
        RECT 440.400 574.050 441.450 634.950 ;
        RECT 449.400 634.050 450.450 691.950 ;
        RECT 460.950 682.950 463.050 685.050 ;
        RECT 451.950 676.950 454.050 679.050 ;
        RECT 452.400 670.050 453.450 676.950 ;
        RECT 461.400 673.050 462.450 682.950 ;
        RECT 454.950 670.950 457.050 673.050 ;
        RECT 458.250 671.250 459.750 672.150 ;
        RECT 460.950 670.950 463.050 673.050 ;
        RECT 451.950 667.950 454.050 670.050 ;
        RECT 455.250 668.850 456.750 669.750 ;
        RECT 457.950 667.950 460.050 670.050 ;
        RECT 461.250 668.850 463.050 669.750 ;
        RECT 451.950 665.850 454.050 666.750 ;
        RECT 464.400 640.050 465.450 706.950 ;
        RECT 469.950 703.950 472.050 706.050 ;
        RECT 470.400 703.050 471.450 703.950 ;
        RECT 469.950 700.950 472.050 703.050 ;
        RECT 466.950 698.250 469.050 699.150 ;
        RECT 469.950 698.850 472.050 699.750 ;
        RECT 466.950 694.950 469.050 697.050 ;
        RECT 467.400 694.050 468.450 694.950 ;
        RECT 466.950 691.950 469.050 694.050 ;
        RECT 473.400 691.050 474.450 764.400 ;
        RECT 476.400 751.050 477.450 769.950 ;
        RECT 481.950 766.950 484.050 769.050 ;
        RECT 500.400 766.050 501.450 769.950 ;
        RECT 518.400 766.050 519.450 808.950 ;
        RECT 521.400 778.050 522.450 811.950 ;
        RECT 527.400 808.050 528.450 811.950 ;
        RECT 526.950 805.950 529.050 808.050 ;
        RECT 533.400 805.050 534.450 815.400 ;
        RECT 539.400 814.050 540.450 817.950 ;
        RECT 560.400 817.050 561.450 817.950 ;
        RECT 541.950 814.950 544.050 817.050 ;
        RECT 547.950 816.450 550.050 817.050 ;
        RECT 545.250 815.250 546.750 816.150 ;
        RECT 547.950 815.400 552.450 816.450 ;
        RECT 547.950 814.950 550.050 815.400 ;
        RECT 538.950 811.950 541.050 814.050 ;
        RECT 542.250 812.850 543.750 813.750 ;
        RECT 544.950 811.950 547.050 814.050 ;
        RECT 548.250 812.850 550.050 813.750 ;
        RECT 545.400 811.050 546.450 811.950 ;
        RECT 538.950 809.850 541.050 810.750 ;
        RECT 544.950 808.950 547.050 811.050 ;
        RECT 541.950 805.950 544.050 808.050 ;
        RECT 532.950 802.950 535.050 805.050 ;
        RECT 520.950 775.950 523.050 778.050 ;
        RECT 529.950 776.250 532.050 777.150 ;
        RECT 520.950 773.250 522.750 774.150 ;
        RECT 523.950 772.950 526.050 775.050 ;
        RECT 527.250 773.250 528.750 774.150 ;
        RECT 529.950 772.950 532.050 775.050 ;
        RECT 530.400 772.050 531.450 772.950 ;
        RECT 520.950 769.950 523.050 772.050 ;
        RECT 524.250 770.850 525.750 771.750 ;
        RECT 526.950 769.950 529.050 772.050 ;
        RECT 529.950 769.950 532.050 772.050 ;
        RECT 499.950 763.950 502.050 766.050 ;
        RECT 517.950 763.950 520.050 766.050 ;
        RECT 527.400 754.050 528.450 769.950 ;
        RECT 533.400 769.050 534.450 802.950 ;
        RECT 542.400 775.050 543.450 805.950 ;
        RECT 551.400 805.050 552.450 815.400 ;
        RECT 553.950 814.950 556.050 817.050 ;
        RECT 557.250 815.250 558.750 816.150 ;
        RECT 559.950 814.950 562.050 817.050 ;
        RECT 574.950 815.250 577.050 816.150 ;
        RECT 577.950 815.850 580.050 816.750 ;
        RECT 553.950 812.850 555.750 813.750 ;
        RECT 556.950 811.950 559.050 814.050 ;
        RECT 560.250 812.850 561.750 813.750 ;
        RECT 562.950 813.450 565.050 814.050 ;
        RECT 562.950 812.400 567.450 813.450 ;
        RECT 562.950 811.950 565.050 812.400 ;
        RECT 557.400 805.050 558.450 811.950 ;
        RECT 562.950 809.850 565.050 810.750 ;
        RECT 566.400 808.050 567.450 812.400 ;
        RECT 574.950 811.950 577.050 814.050 ;
        RECT 577.950 808.950 580.050 811.050 ;
        RECT 581.400 810.450 582.450 818.400 ;
        RECT 593.400 818.400 598.050 819.450 ;
        RECT 583.950 812.250 585.750 813.150 ;
        RECT 586.950 811.950 589.050 814.050 ;
        RECT 590.250 812.250 592.050 813.150 ;
        RECT 583.950 810.450 586.050 811.050 ;
        RECT 581.400 809.400 586.050 810.450 ;
        RECT 587.250 809.850 588.750 810.750 ;
        RECT 589.950 810.450 592.050 811.050 ;
        RECT 593.400 810.450 594.450 818.400 ;
        RECT 595.950 817.950 598.050 818.400 ;
        RECT 691.950 817.950 694.050 820.050 ;
        RECT 754.950 817.950 757.050 820.050 ;
        RECT 787.950 817.950 790.050 820.050 ;
        RECT 790.950 817.950 793.050 820.050 ;
        RECT 595.950 815.850 598.050 816.750 ;
        RECT 598.950 815.250 601.050 816.150 ;
        RECT 601.950 814.950 604.050 817.050 ;
        RECT 613.950 814.950 616.050 817.050 ;
        RECT 617.250 815.250 618.750 816.150 ;
        RECT 619.950 814.950 622.050 817.050 ;
        RECT 637.950 814.950 640.050 817.050 ;
        RECT 640.950 815.250 642.750 816.150 ;
        RECT 643.950 814.950 646.050 817.050 ;
        RECT 652.950 814.950 655.050 817.050 ;
        RECT 676.950 814.950 679.050 817.050 ;
        RECT 598.950 811.950 601.050 814.050 ;
        RECT 565.950 805.950 568.050 808.050 ;
        RECT 550.950 802.950 553.050 805.050 ;
        RECT 556.950 802.950 559.050 805.050 ;
        RECT 557.400 786.450 558.450 802.950 ;
        RECT 554.400 785.400 558.450 786.450 ;
        RECT 554.400 775.050 555.450 785.400 ;
        RECT 574.950 778.950 577.050 781.050 ;
        RECT 571.950 775.950 574.050 778.050 ;
        RECT 572.400 775.050 573.450 775.950 ;
        RECT 535.950 772.950 538.050 775.050 ;
        RECT 538.950 773.250 540.750 774.150 ;
        RECT 541.950 772.950 544.050 775.050 ;
        RECT 545.250 773.250 546.750 774.150 ;
        RECT 547.950 772.950 550.050 775.050 ;
        RECT 551.250 773.250 553.050 774.150 ;
        RECT 553.950 772.950 556.050 775.050 ;
        RECT 556.950 773.250 559.050 774.150 ;
        RECT 562.950 773.250 565.050 774.150 ;
        RECT 571.950 772.950 574.050 775.050 ;
        RECT 532.950 766.950 535.050 769.050 ;
        RECT 536.400 760.050 537.450 772.950 ;
        RECT 538.950 769.950 541.050 772.050 ;
        RECT 542.250 770.850 543.750 771.750 ;
        RECT 544.950 769.950 547.050 772.050 ;
        RECT 548.250 770.850 549.750 771.750 ;
        RECT 550.950 769.950 553.050 772.050 ;
        RECT 539.400 769.050 540.450 769.950 ;
        RECT 538.950 766.950 541.050 769.050 ;
        RECT 550.950 766.950 553.050 769.050 ;
        RECT 551.400 766.050 552.450 766.950 ;
        RECT 550.950 763.950 553.050 766.050 ;
        RECT 535.950 757.950 538.050 760.050 ;
        RECT 478.950 751.950 481.050 754.050 ;
        RECT 526.950 751.950 529.050 754.050 ;
        RECT 475.950 748.950 478.050 751.050 ;
        RECT 475.950 739.950 478.050 742.050 ;
        RECT 472.950 688.950 475.050 691.050 ;
        RECT 476.400 688.050 477.450 739.950 ;
        RECT 479.400 738.450 480.450 751.950 ;
        RECT 508.950 748.950 511.050 751.050 ;
        RECT 514.950 748.950 517.050 751.050 ;
        RECT 502.950 745.950 505.050 748.050 ;
        RECT 496.950 744.450 499.050 745.050 ;
        RECT 494.400 743.400 499.050 744.450 ;
        RECT 481.950 740.250 483.750 741.150 ;
        RECT 484.950 739.950 487.050 742.050 ;
        RECT 488.250 740.250 490.050 741.150 ;
        RECT 494.400 739.050 495.450 743.400 ;
        RECT 496.950 742.950 499.050 743.400 ;
        RECT 500.250 743.250 502.050 744.150 ;
        RECT 502.950 743.850 505.050 744.750 ;
        RECT 505.950 743.250 508.050 744.150 ;
        RECT 509.400 742.050 510.450 748.950 ;
        RECT 515.400 748.050 516.450 748.950 ;
        RECT 514.950 745.950 517.050 748.050 ;
        RECT 535.950 745.950 538.050 748.050 ;
        RECT 511.950 742.950 514.050 745.050 ;
        RECT 515.250 743.850 516.750 744.750 ;
        RECT 517.950 744.450 520.050 745.050 ;
        RECT 517.950 743.400 522.450 744.450 ;
        RECT 517.950 742.950 520.050 743.400 ;
        RECT 496.950 740.850 498.750 741.750 ;
        RECT 499.950 739.950 502.050 742.050 ;
        RECT 505.950 739.950 508.050 742.050 ;
        RECT 508.950 739.950 511.050 742.050 ;
        RECT 511.950 740.850 514.050 741.750 ;
        RECT 514.950 739.950 517.050 742.050 ;
        RECT 517.950 740.850 520.050 741.750 ;
        RECT 481.950 738.450 484.050 739.050 ;
        RECT 479.400 737.400 484.050 738.450 ;
        RECT 485.250 737.850 486.750 738.750 ;
        RECT 481.950 736.950 484.050 737.400 ;
        RECT 487.950 736.950 490.050 739.050 ;
        RECT 493.950 736.950 496.050 739.050 ;
        RECT 506.400 736.050 507.450 739.950 ;
        RECT 499.950 733.950 502.050 736.050 ;
        RECT 505.950 733.950 508.050 736.050 ;
        RECT 496.950 712.950 499.050 715.050 ;
        RECT 478.950 709.950 481.050 712.050 ;
        RECT 479.400 700.050 480.450 709.950 ;
        RECT 481.950 706.950 484.050 709.050 ;
        RECT 482.400 706.050 483.450 706.950 ;
        RECT 481.950 703.950 484.050 706.050 ;
        RECT 485.250 704.250 486.750 705.150 ;
        RECT 487.950 703.950 490.050 706.050 ;
        RECT 493.950 703.950 496.050 706.050 ;
        RECT 481.950 701.850 483.750 702.750 ;
        RECT 484.950 700.950 487.050 703.050 ;
        RECT 488.250 701.850 490.050 702.750 ;
        RECT 485.400 700.050 486.450 700.950 ;
        RECT 478.950 697.950 481.050 700.050 ;
        RECT 484.950 697.950 487.050 700.050 ;
        RECT 494.400 694.050 495.450 703.950 ;
        RECT 493.950 691.950 496.050 694.050 ;
        RECT 475.950 685.950 478.050 688.050 ;
        RECT 493.950 682.950 496.050 685.050 ;
        RECT 466.950 679.950 469.050 682.050 ;
        RECT 478.950 679.950 481.050 682.050 ;
        RECT 467.400 673.050 468.450 679.950 ;
        RECT 472.950 676.950 475.050 679.050 ;
        RECT 473.400 673.050 474.450 676.950 ;
        RECT 479.400 673.050 480.450 679.950 ;
        RECT 481.950 676.950 484.050 679.050 ;
        RECT 482.400 676.050 483.450 676.950 ;
        RECT 481.950 673.950 484.050 676.050 ;
        RECT 466.950 670.950 469.050 673.050 ;
        RECT 470.250 671.250 471.750 672.150 ;
        RECT 472.950 670.950 475.050 673.050 ;
        RECT 476.250 671.250 477.750 672.150 ;
        RECT 478.950 670.950 481.050 673.050 ;
        RECT 466.950 668.850 468.750 669.750 ;
        RECT 469.950 667.950 472.050 670.050 ;
        RECT 473.250 668.850 474.750 669.750 ;
        RECT 475.950 667.950 478.050 670.050 ;
        RECT 479.250 668.850 481.050 669.750 ;
        RECT 470.400 649.050 471.450 667.950 ;
        RECT 476.400 667.050 477.450 667.950 ;
        RECT 475.950 664.950 478.050 667.050 ;
        RECT 472.950 652.950 475.050 655.050 ;
        RECT 469.950 646.950 472.050 649.050 ;
        RECT 463.950 637.950 466.050 640.050 ;
        RECT 466.950 634.950 469.050 637.050 ;
        RECT 448.950 631.950 451.050 634.050 ;
        RECT 463.950 631.950 466.050 634.050 ;
        RECT 442.950 629.250 444.750 630.150 ;
        RECT 445.950 628.950 448.050 631.050 ;
        RECT 451.950 630.450 454.050 631.050 ;
        RECT 451.950 629.400 456.450 630.450 ;
        RECT 451.950 628.950 454.050 629.400 ;
        RECT 442.950 625.950 445.050 628.050 ;
        RECT 446.250 626.850 448.050 627.750 ;
        RECT 448.950 626.250 451.050 627.150 ;
        RECT 451.950 626.850 454.050 627.750 ;
        RECT 448.950 622.950 451.050 625.050 ;
        RECT 442.950 613.950 445.050 616.050 ;
        RECT 443.400 598.050 444.450 613.950 ;
        RECT 449.400 613.050 450.450 622.950 ;
        RECT 455.400 616.050 456.450 629.400 ;
        RECT 460.950 629.250 463.050 630.150 ;
        RECT 460.950 625.950 463.050 628.050 ;
        RECT 461.400 625.050 462.450 625.950 ;
        RECT 460.950 622.950 463.050 625.050 ;
        RECT 454.950 613.950 457.050 616.050 ;
        RECT 448.950 610.950 451.050 613.050 ;
        RECT 454.950 610.950 457.050 613.050 ;
        RECT 460.950 610.950 463.050 613.050 ;
        RECT 448.950 601.950 451.050 604.050 ;
        RECT 445.950 599.250 448.050 600.150 ;
        RECT 448.950 599.850 451.050 600.750 ;
        RECT 455.400 598.050 456.450 610.950 ;
        RECT 442.950 595.950 445.050 598.050 ;
        RECT 445.950 595.950 448.050 598.050 ;
        RECT 451.950 596.250 453.750 597.150 ;
        RECT 454.950 595.950 457.050 598.050 ;
        RECT 458.250 596.250 460.050 597.150 ;
        RECT 461.400 595.050 462.450 610.950 ;
        RECT 464.400 603.450 465.450 631.950 ;
        RECT 467.400 631.050 468.450 634.950 ;
        RECT 466.950 628.950 469.050 631.050 ;
        RECT 470.250 629.250 472.050 630.150 ;
        RECT 466.950 626.850 468.750 627.750 ;
        RECT 469.950 625.950 472.050 628.050 ;
        RECT 469.950 622.950 472.050 625.050 ;
        RECT 470.400 604.050 471.450 622.950 ;
        RECT 464.400 602.400 468.450 603.450 ;
        RECT 448.950 592.950 451.050 595.050 ;
        RECT 451.950 592.950 454.050 595.050 ;
        RECT 455.250 593.850 456.750 594.750 ;
        RECT 457.950 592.950 460.050 595.050 ;
        RECT 460.950 592.950 463.050 595.050 ;
        RECT 449.400 580.050 450.450 592.950 ;
        RECT 452.400 583.050 453.450 592.950 ;
        RECT 463.950 583.950 466.050 586.050 ;
        RECT 451.950 580.950 454.050 583.050 ;
        RECT 448.950 577.950 451.050 580.050 ;
        RECT 439.950 571.950 442.050 574.050 ;
        RECT 445.950 571.950 448.050 574.050 ;
        RECT 400.950 568.950 403.050 571.050 ;
        RECT 412.800 569.100 414.900 571.200 ;
        RECT 391.950 559.950 394.050 562.050 ;
        RECT 394.950 559.950 397.050 562.050 ;
        RECT 391.950 558.450 394.050 559.050 ;
        RECT 391.950 557.400 396.450 558.450 ;
        RECT 391.950 556.950 394.050 557.400 ;
        RECT 391.950 554.850 394.050 555.750 ;
        RECT 388.950 535.950 391.050 538.050 ;
        RECT 379.950 532.950 382.050 535.050 ;
        RECT 385.950 532.950 388.050 535.050 ;
        RECT 380.400 526.050 381.450 532.950 ;
        RECT 382.950 529.950 385.050 532.050 ;
        RECT 388.950 529.950 391.050 532.050 ;
        RECT 383.400 529.050 384.450 529.950 ;
        RECT 382.950 526.950 385.050 529.050 ;
        RECT 386.250 527.250 388.050 528.150 ;
        RECT 388.950 527.850 391.050 528.750 ;
        RECT 391.950 527.250 394.050 528.150 ;
        RECT 379.950 523.950 382.050 526.050 ;
        RECT 382.950 524.850 384.750 525.750 ;
        RECT 385.950 523.950 388.050 526.050 ;
        RECT 388.950 523.950 391.050 526.050 ;
        RECT 391.950 523.950 394.050 526.050 ;
        RECT 382.950 491.250 385.050 492.150 ;
        RECT 389.400 490.050 390.450 523.950 ;
        RECT 392.400 523.050 393.450 523.950 ;
        RECT 391.950 520.950 394.050 523.050 ;
        RECT 392.400 520.050 393.450 520.950 ;
        RECT 391.950 517.950 394.050 520.050 ;
        RECT 391.950 511.950 394.050 514.050 ;
        RECT 392.400 493.050 393.450 511.950 ;
        RECT 395.400 502.050 396.450 557.400 ;
        RECT 401.400 553.050 402.450 568.950 ;
        RECT 413.550 565.350 414.750 569.100 ;
        RECT 436.950 568.950 439.050 571.050 ;
        RECT 439.950 568.950 442.050 571.050 ;
        RECT 442.950 568.950 445.050 571.050 ;
        RECT 415.950 566.850 418.050 568.950 ;
        RECT 412.950 563.250 415.050 565.350 ;
        RECT 403.950 560.250 406.050 561.150 ;
        RECT 403.950 556.950 406.050 559.050 ;
        RECT 400.950 550.950 403.050 553.050 ;
        RECT 404.400 547.050 405.450 556.950 ;
        RECT 413.550 549.600 414.750 563.250 ;
        RECT 416.250 549.600 417.450 566.850 ;
        RECT 423.900 566.400 426.000 568.500 ;
        RECT 427.950 566.400 430.050 568.500 ;
        RECT 418.950 563.250 421.050 565.350 ;
        RECT 419.400 549.600 420.600 563.250 ;
        RECT 424.350 557.550 425.550 566.400 ;
        RECT 428.550 560.250 429.750 566.400 ;
        RECT 427.950 558.150 430.050 560.250 ;
        RECT 423.750 555.450 425.850 557.550 ;
        RECT 424.350 549.600 425.550 555.450 ;
        RECT 428.550 549.600 429.750 558.150 ;
        RECT 430.950 554.250 433.050 555.150 ;
        RECT 430.950 550.950 433.050 553.050 ;
        RECT 412.950 547.500 415.050 549.600 ;
        RECT 415.950 547.500 418.050 549.600 ;
        RECT 418.950 547.500 421.050 549.600 ;
        RECT 423.750 547.500 425.850 549.600 ;
        RECT 427.950 547.500 430.050 549.600 ;
        RECT 403.950 544.950 406.050 547.050 ;
        RECT 415.950 532.950 418.050 535.050 ;
        RECT 427.950 532.950 430.050 535.050 ;
        RECT 403.950 529.950 406.050 532.050 ;
        RECT 404.400 529.050 405.450 529.950 ;
        RECT 416.400 529.050 417.450 532.950 ;
        RECT 397.950 526.950 400.050 529.050 ;
        RECT 401.250 527.250 402.750 528.150 ;
        RECT 403.950 526.950 406.050 529.050 ;
        RECT 406.950 526.950 409.050 529.050 ;
        RECT 415.950 526.950 418.050 529.050 ;
        RECT 419.250 527.250 420.750 528.150 ;
        RECT 421.950 526.950 424.050 529.050 ;
        RECT 407.400 526.050 408.450 526.950 ;
        RECT 397.950 524.850 399.750 525.750 ;
        RECT 400.950 523.950 403.050 526.050 ;
        RECT 404.250 524.850 405.750 525.750 ;
        RECT 406.950 523.950 409.050 526.050 ;
        RECT 415.950 524.850 417.750 525.750 ;
        RECT 418.950 523.950 421.050 526.050 ;
        RECT 422.250 524.850 423.750 525.750 ;
        RECT 424.950 523.950 427.050 526.050 ;
        RECT 401.400 511.050 402.450 523.950 ;
        RECT 406.950 521.850 409.050 522.750 ;
        RECT 412.950 520.950 415.050 523.050 ;
        RECT 413.400 520.050 414.450 520.950 ;
        RECT 412.950 517.950 415.050 520.050 ;
        RECT 400.950 508.950 403.050 511.050 ;
        RECT 406.950 502.950 409.050 505.050 ;
        RECT 394.950 499.950 397.050 502.050 ;
        RECT 391.950 490.950 394.050 493.050 ;
        RECT 379.950 488.250 381.750 489.150 ;
        RECT 382.950 487.950 385.050 490.050 ;
        RECT 386.250 488.250 387.750 489.150 ;
        RECT 388.950 487.950 391.050 490.050 ;
        RECT 379.950 484.950 382.050 487.050 ;
        RECT 382.950 484.950 385.050 487.050 ;
        RECT 385.950 484.950 388.050 487.050 ;
        RECT 389.250 485.850 391.050 486.750 ;
        RECT 380.400 478.050 381.450 484.950 ;
        RECT 379.950 475.950 382.050 478.050 ;
        RECT 380.400 475.050 381.450 475.950 ;
        RECT 379.950 472.950 382.050 475.050 ;
        RECT 376.950 463.950 379.050 466.050 ;
        RECT 383.400 460.050 384.450 484.950 ;
        RECT 386.400 484.050 387.450 484.950 ;
        RECT 385.950 481.950 388.050 484.050 ;
        RECT 392.400 481.050 393.450 490.950 ;
        RECT 395.400 487.050 396.450 499.950 ;
        RECT 397.950 493.950 400.050 496.050 ;
        RECT 394.950 484.950 397.050 487.050 ;
        RECT 398.400 484.050 399.450 493.950 ;
        RECT 407.400 493.050 408.450 502.950 ;
        RECT 406.950 490.950 409.050 493.050 ;
        RECT 400.950 488.250 403.050 489.150 ;
        RECT 407.400 487.050 408.450 490.950 ;
        RECT 400.950 484.950 403.050 487.050 ;
        RECT 404.250 485.250 405.750 486.150 ;
        RECT 406.950 484.950 409.050 487.050 ;
        RECT 410.250 485.250 412.050 486.150 ;
        RECT 397.950 481.950 400.050 484.050 ;
        RECT 403.950 481.950 406.050 484.050 ;
        RECT 407.250 482.850 408.750 483.750 ;
        RECT 409.950 481.950 412.050 484.050 ;
        RECT 391.950 478.950 394.050 481.050 ;
        RECT 385.950 472.950 388.050 475.050 ;
        RECT 409.950 472.950 412.050 475.050 ;
        RECT 376.950 457.950 379.050 460.050 ;
        RECT 382.950 457.950 385.050 460.050 ;
        RECT 373.950 424.950 376.050 427.050 ;
        RECT 377.400 424.050 378.450 457.950 ;
        RECT 386.400 457.050 387.450 472.950 ;
        RECT 400.950 469.950 403.050 472.050 ;
        RECT 406.950 469.950 409.050 472.050 ;
        RECT 391.950 466.950 394.050 469.050 ;
        RECT 397.950 466.950 400.050 469.050 ;
        RECT 388.950 460.950 391.050 463.050 ;
        RECT 379.950 455.250 382.050 456.150 ;
        RECT 382.950 455.850 385.050 456.750 ;
        RECT 385.950 454.950 388.050 457.050 ;
        RECT 379.950 451.950 382.050 454.050 ;
        RECT 385.950 451.950 388.050 454.050 ;
        RECT 380.400 448.050 381.450 451.950 ;
        RECT 379.950 445.950 382.050 448.050 ;
        RECT 380.400 430.050 381.450 445.950 ;
        RECT 386.400 445.050 387.450 451.950 ;
        RECT 385.950 442.950 388.050 445.050 ;
        RECT 389.400 436.050 390.450 460.950 ;
        RECT 392.400 460.050 393.450 466.950 ;
        RECT 394.950 463.950 397.050 466.050 ;
        RECT 395.400 460.050 396.450 463.950 ;
        RECT 398.400 460.050 399.450 466.950 ;
        RECT 391.950 457.950 394.050 460.050 ;
        RECT 394.950 457.950 397.050 460.050 ;
        RECT 397.950 457.950 400.050 460.050 ;
        RECT 388.950 433.950 391.050 436.050 ;
        RECT 379.950 427.950 382.050 430.050 ;
        RECT 379.950 424.950 382.050 427.050 ;
        RECT 376.950 421.950 379.050 424.050 ;
        RECT 370.950 419.250 373.050 420.150 ;
        RECT 364.950 415.950 367.050 418.050 ;
        RECT 367.950 416.250 369.750 417.150 ;
        RECT 370.950 415.950 373.050 418.050 ;
        RECT 374.250 416.250 375.750 417.150 ;
        RECT 376.950 415.950 379.050 418.050 ;
        RECT 367.950 412.950 370.050 415.050 ;
        RECT 373.950 412.950 376.050 415.050 ;
        RECT 377.250 413.850 379.050 414.750 ;
        RECT 368.400 406.050 369.450 412.950 ;
        RECT 367.950 403.950 370.050 406.050 ;
        RECT 370.950 397.950 373.050 400.050 ;
        RECT 371.400 385.050 372.450 397.950 ;
        RECT 374.400 391.050 375.450 412.950 ;
        RECT 380.400 408.450 381.450 424.950 ;
        RECT 392.400 421.050 393.450 457.950 ;
        RECT 401.400 457.050 402.450 469.950 ;
        RECT 403.950 460.950 406.050 463.050 ;
        RECT 394.950 454.950 397.050 457.050 ;
        RECT 398.250 455.850 399.750 456.750 ;
        RECT 400.950 454.950 403.050 457.050 ;
        RECT 394.950 452.850 397.050 453.750 ;
        RECT 400.950 452.850 403.050 453.750 ;
        RECT 391.950 418.950 394.050 421.050 ;
        RECT 404.400 420.450 405.450 460.950 ;
        RECT 407.400 457.050 408.450 469.950 ;
        RECT 406.950 454.950 409.050 457.050 ;
        RECT 410.400 454.050 411.450 472.950 ;
        RECT 413.400 472.050 414.450 517.950 ;
        RECT 415.950 502.950 418.050 505.050 ;
        RECT 416.400 483.450 417.450 502.950 ;
        RECT 419.400 493.050 420.450 523.950 ;
        RECT 424.950 521.850 427.050 522.750 ;
        RECT 424.950 508.950 427.050 511.050 ;
        RECT 418.950 490.950 421.050 493.050 ;
        RECT 418.950 488.250 421.050 489.150 ;
        RECT 425.400 487.050 426.450 508.950 ;
        RECT 428.400 499.050 429.450 532.950 ;
        RECT 431.400 505.050 432.450 550.950 ;
        RECT 437.250 550.050 438.450 568.950 ;
        RECT 440.250 564.750 441.450 568.950 ;
        RECT 439.950 562.650 442.050 564.750 ;
        RECT 440.250 550.050 441.450 562.650 ;
        RECT 443.250 550.050 444.450 568.950 ;
        RECT 436.950 547.950 439.050 550.050 ;
        RECT 439.950 547.950 442.050 550.050 ;
        RECT 442.950 547.950 445.050 550.050 ;
        RECT 442.950 544.950 445.050 547.050 ;
        RECT 433.950 527.250 436.050 528.150 ;
        RECT 433.950 523.950 436.050 526.050 ;
        RECT 443.400 525.450 444.450 544.950 ;
        RECT 446.400 529.050 447.450 571.950 ;
        RECT 454.950 561.450 457.050 562.050 ;
        RECT 448.950 560.250 451.050 561.150 ;
        RECT 452.400 560.400 457.050 561.450 ;
        RECT 452.400 550.050 453.450 560.400 ;
        RECT 454.950 559.950 457.050 560.400 ;
        RECT 464.400 559.050 465.450 583.950 ;
        RECT 454.950 557.850 457.050 558.750 ;
        RECT 463.950 556.950 466.050 559.050 ;
        RECT 460.950 554.250 463.050 555.150 ;
        RECT 463.950 554.850 466.050 555.750 ;
        RECT 460.950 550.950 463.050 553.050 ;
        RECT 451.950 547.950 454.050 550.050 ;
        RECT 445.950 526.950 448.050 529.050 ;
        RECT 445.950 525.450 448.050 526.050 ;
        RECT 443.400 524.400 448.050 525.450 ;
        RECT 434.400 514.050 435.450 523.950 ;
        RECT 443.400 514.050 444.450 524.400 ;
        RECT 445.950 523.950 448.050 524.400 ;
        RECT 445.950 521.850 448.050 522.750 ;
        RECT 452.400 520.050 453.450 547.950 ;
        RECT 467.400 541.050 468.450 602.400 ;
        RECT 469.950 601.950 472.050 604.050 ;
        RECT 473.400 603.450 474.450 652.950 ;
        RECT 478.950 646.950 481.050 649.050 ;
        RECT 475.950 631.950 478.050 634.050 ;
        RECT 476.400 631.050 477.450 631.950 ;
        RECT 475.950 628.950 478.050 631.050 ;
        RECT 479.400 628.050 480.450 646.950 ;
        RECT 475.950 626.850 478.050 627.750 ;
        RECT 478.950 625.950 481.050 628.050 ;
        RECT 482.400 603.450 483.450 673.950 ;
        RECT 494.400 673.050 495.450 682.950 ;
        RECT 497.400 676.050 498.450 712.950 ;
        RECT 500.400 697.050 501.450 733.950 ;
        RECT 502.950 724.950 505.050 727.050 ;
        RECT 503.400 706.050 504.450 724.950 ;
        RECT 508.950 707.250 511.050 708.150 ;
        RECT 502.950 703.950 505.050 706.050 ;
        RECT 506.250 704.250 507.750 705.150 ;
        RECT 508.950 703.950 511.050 706.050 ;
        RECT 512.250 704.250 514.050 705.150 ;
        RECT 502.950 701.850 504.750 702.750 ;
        RECT 505.950 700.950 508.050 703.050 ;
        RECT 499.950 694.950 502.050 697.050 ;
        RECT 496.950 673.950 499.050 676.050 ;
        RECT 500.400 673.050 501.450 694.950 ;
        RECT 506.400 694.050 507.450 700.950 ;
        RECT 509.400 700.050 510.450 703.950 ;
        RECT 511.950 700.950 514.050 703.050 ;
        RECT 508.950 697.950 511.050 700.050 ;
        RECT 505.950 691.950 508.050 694.050 ;
        RECT 508.950 688.950 511.050 691.050 ;
        RECT 505.950 685.950 508.050 688.050 ;
        RECT 502.950 682.950 505.050 685.050 ;
        RECT 487.950 672.450 490.050 673.050 ;
        RECT 485.400 671.400 490.050 672.450 ;
        RECT 485.400 667.050 486.450 671.400 ;
        RECT 487.950 670.950 490.050 671.400 ;
        RECT 491.250 671.250 492.750 672.150 ;
        RECT 493.950 670.950 496.050 673.050 ;
        RECT 497.250 671.250 498.750 672.150 ;
        RECT 499.950 670.950 502.050 673.050 ;
        RECT 487.950 668.850 489.750 669.750 ;
        RECT 490.950 667.950 493.050 670.050 ;
        RECT 494.250 668.850 495.750 669.750 ;
        RECT 496.950 667.950 499.050 670.050 ;
        RECT 500.250 668.850 502.050 669.750 ;
        RECT 497.400 667.050 498.450 667.950 ;
        RECT 484.950 664.950 487.050 667.050 ;
        RECT 496.950 664.950 499.050 667.050 ;
        RECT 499.950 664.950 502.050 667.050 ;
        RECT 490.950 640.950 493.050 643.050 ;
        RECT 484.950 634.950 487.050 637.050 ;
        RECT 485.400 625.050 486.450 634.950 ;
        RECT 491.400 634.050 492.450 640.950 ;
        RECT 500.400 637.050 501.450 664.950 ;
        RECT 503.400 643.050 504.450 682.950 ;
        RECT 506.400 655.050 507.450 685.950 ;
        RECT 509.400 675.450 510.450 688.950 ;
        RECT 512.400 688.050 513.450 700.950 ;
        RECT 511.950 685.950 514.050 688.050 ;
        RECT 515.400 679.050 516.450 739.950 ;
        RECT 521.400 739.050 522.450 743.400 ;
        RECT 532.950 743.250 535.050 744.150 ;
        RECT 535.950 743.850 538.050 744.750 ;
        RECT 532.950 739.950 535.050 742.050 ;
        RECT 538.950 740.250 540.750 741.150 ;
        RECT 541.950 739.950 544.050 742.050 ;
        RECT 545.250 740.250 547.050 741.150 ;
        RECT 520.950 736.950 523.050 739.050 ;
        RECT 517.950 697.950 520.050 700.050 ;
        RECT 514.950 676.950 517.050 679.050 ;
        RECT 514.950 675.450 517.050 676.050 ;
        RECT 509.400 674.400 517.050 675.450 ;
        RECT 505.950 652.950 508.050 655.050 ;
        RECT 505.950 649.950 508.050 652.050 ;
        RECT 502.950 640.950 505.050 643.050 ;
        RECT 493.950 634.950 496.050 637.050 ;
        RECT 499.950 634.950 502.050 637.050 ;
        RECT 506.400 636.450 507.450 649.950 ;
        RECT 509.400 637.050 510.450 674.400 ;
        RECT 514.950 673.950 517.050 674.400 ;
        RECT 511.950 671.250 514.050 672.150 ;
        RECT 514.950 671.850 517.050 672.750 ;
        RECT 511.950 667.950 514.050 670.050 ;
        RECT 514.950 667.950 517.050 670.050 ;
        RECT 512.400 667.050 513.450 667.950 ;
        RECT 515.400 667.050 516.450 667.950 ;
        RECT 511.950 664.950 514.050 667.050 ;
        RECT 514.950 664.950 517.050 667.050 ;
        RECT 518.400 637.050 519.450 697.950 ;
        RECT 503.400 635.400 507.450 636.450 ;
        RECT 494.400 634.050 495.450 634.950 ;
        RECT 490.950 631.950 493.050 634.050 ;
        RECT 493.950 631.950 496.050 634.050 ;
        RECT 497.250 632.250 498.750 633.150 ;
        RECT 499.950 631.950 502.050 634.050 ;
        RECT 484.950 622.950 487.050 625.050 ;
        RECT 484.950 604.950 487.050 607.050 ;
        RECT 485.400 604.050 486.450 604.950 ;
        RECT 473.400 602.400 477.450 603.450 ;
        RECT 469.950 599.850 472.050 600.750 ;
        RECT 472.950 599.250 475.050 600.150 ;
        RECT 469.950 595.950 472.050 598.050 ;
        RECT 472.950 595.950 475.050 598.050 ;
        RECT 470.400 592.050 471.450 595.950 ;
        RECT 469.950 589.950 472.050 592.050 ;
        RECT 472.950 580.950 475.050 583.050 ;
        RECT 473.400 553.050 474.450 580.950 ;
        RECT 476.400 565.050 477.450 602.400 ;
        RECT 479.400 602.400 483.450 603.450 ;
        RECT 475.950 562.950 478.050 565.050 ;
        RECT 479.400 564.450 480.450 602.400 ;
        RECT 484.950 601.950 487.050 604.050 ;
        RECT 491.400 601.050 492.450 631.950 ;
        RECT 493.950 629.850 495.750 630.750 ;
        RECT 496.950 628.950 499.050 631.050 ;
        RECT 500.250 629.850 502.050 630.750 ;
        RECT 497.400 628.050 498.450 628.950 ;
        RECT 496.950 625.950 499.050 628.050 ;
        RECT 493.950 610.950 496.050 613.050 ;
        RECT 481.950 599.250 484.050 600.150 ;
        RECT 484.950 599.850 487.050 600.750 ;
        RECT 490.950 598.950 493.050 601.050 ;
        RECT 494.400 598.050 495.450 610.950 ;
        RECT 497.400 607.050 498.450 625.950 ;
        RECT 496.950 604.950 499.050 607.050 ;
        RECT 503.400 598.050 504.450 635.400 ;
        RECT 508.950 634.950 511.050 637.050 ;
        RECT 511.950 634.950 514.050 637.050 ;
        RECT 517.950 634.950 520.050 637.050 ;
        RECT 512.400 634.050 513.450 634.950 ;
        RECT 521.400 634.050 522.450 736.950 ;
        RECT 533.400 732.450 534.450 739.950 ;
        RECT 538.950 736.950 541.050 739.050 ;
        RECT 542.250 737.850 543.750 738.750 ;
        RECT 544.950 736.950 547.050 739.050 ;
        RECT 533.400 731.400 537.450 732.450 ;
        RECT 532.950 727.950 535.050 730.050 ;
        RECT 523.950 701.250 526.050 702.150 ;
        RECT 529.950 701.250 532.050 702.150 ;
        RECT 523.950 697.950 526.050 700.050 ;
        RECT 527.250 698.250 528.750 699.150 ;
        RECT 529.950 697.950 532.050 700.050 ;
        RECT 524.400 694.050 525.450 697.950 ;
        RECT 526.950 694.950 529.050 697.050 ;
        RECT 523.950 691.950 526.050 694.050 ;
        RECT 523.950 679.950 526.050 682.050 ;
        RECT 524.400 676.050 525.450 679.950 ;
        RECT 527.400 678.450 528.450 694.950 ;
        RECT 533.400 691.050 534.450 727.950 ;
        RECT 536.400 703.050 537.450 731.400 ;
        RECT 539.400 703.050 540.450 736.950 ;
        RECT 545.400 736.050 546.450 736.950 ;
        RECT 544.950 733.950 547.050 736.050 ;
        RECT 551.400 727.050 552.450 763.950 ;
        RECT 550.950 724.950 553.050 727.050 ;
        RECT 554.400 712.050 555.450 772.950 ;
        RECT 556.950 769.950 559.050 772.050 ;
        RECT 560.250 770.250 561.750 771.150 ;
        RECT 562.950 769.950 565.050 772.050 ;
        RECT 568.950 770.250 571.050 771.150 ;
        RECT 571.950 770.850 574.050 771.750 ;
        RECT 557.400 769.050 558.450 769.950 ;
        RECT 556.950 766.950 559.050 769.050 ;
        RECT 559.950 766.950 562.050 769.050 ;
        RECT 560.400 744.450 561.450 766.950 ;
        RECT 563.400 751.050 564.450 769.950 ;
        RECT 568.950 766.950 571.050 769.050 ;
        RECT 565.950 751.950 568.050 754.050 ;
        RECT 562.950 748.950 565.050 751.050 ;
        RECT 566.400 747.450 567.450 751.950 ;
        RECT 557.400 743.400 561.450 744.450 ;
        RECT 563.400 746.400 567.450 747.450 ;
        RECT 557.400 712.050 558.450 743.400 ;
        RECT 563.400 742.050 564.450 746.400 ;
        RECT 575.400 744.450 576.450 778.950 ;
        RECT 578.400 772.050 579.450 808.950 ;
        RECT 577.950 769.950 580.050 772.050 ;
        RECT 578.400 748.050 579.450 769.950 ;
        RECT 581.400 766.050 582.450 809.400 ;
        RECT 583.950 808.950 586.050 809.400 ;
        RECT 589.950 809.400 594.450 810.450 ;
        RECT 589.950 808.950 592.050 809.400 ;
        RECT 583.950 775.950 586.050 778.050 ;
        RECT 587.250 776.250 588.750 777.150 ;
        RECT 589.950 775.950 592.050 778.050 ;
        RECT 583.950 773.850 585.750 774.750 ;
        RECT 586.950 772.950 589.050 775.050 ;
        RECT 590.250 773.850 592.050 774.750 ;
        RECT 580.950 763.950 583.050 766.050 ;
        RECT 587.400 753.450 588.450 772.950 ;
        RECT 593.400 760.050 594.450 809.400 ;
        RECT 599.400 808.050 600.450 811.950 ;
        RECT 598.950 805.950 601.050 808.050 ;
        RECT 599.400 805.050 600.450 805.950 ;
        RECT 598.950 802.950 601.050 805.050 ;
        RECT 602.400 781.050 603.450 814.950 ;
        RECT 638.400 814.050 639.450 814.950 ;
        RECT 610.950 811.950 613.050 814.050 ;
        RECT 614.250 812.850 615.750 813.750 ;
        RECT 616.950 811.950 619.050 814.050 ;
        RECT 620.250 812.850 622.050 813.750 ;
        RECT 628.950 812.250 630.750 813.150 ;
        RECT 631.950 811.950 634.050 814.050 ;
        RECT 637.950 813.450 640.050 814.050 ;
        RECT 640.950 813.450 643.050 814.050 ;
        RECT 637.950 812.400 643.050 813.450 ;
        RECT 644.250 812.850 646.050 813.750 ;
        RECT 637.950 811.950 640.050 812.400 ;
        RECT 640.950 811.950 643.050 812.400 ;
        RECT 646.950 811.950 649.050 814.050 ;
        RECT 641.400 811.050 642.450 811.950 ;
        RECT 610.950 809.850 613.050 810.750 ;
        RECT 628.950 808.950 631.050 811.050 ;
        RECT 632.250 809.850 633.750 810.750 ;
        RECT 634.950 808.950 637.050 811.050 ;
        RECT 638.250 809.850 640.050 810.750 ;
        RECT 640.950 808.950 643.050 811.050 ;
        RECT 631.950 805.950 634.050 808.050 ;
        RECT 634.950 806.850 637.050 807.750 ;
        RECT 632.400 804.450 633.450 805.950 ;
        RECT 632.400 803.400 636.450 804.450 ;
        RECT 628.950 799.950 631.050 802.050 ;
        RECT 601.950 778.950 604.050 781.050 ;
        RECT 604.950 776.250 607.050 777.150 ;
        RECT 607.950 775.950 610.050 778.050 ;
        RECT 619.950 777.450 622.050 778.050 ;
        RECT 617.400 776.400 622.050 777.450 ;
        RECT 595.950 773.250 597.750 774.150 ;
        RECT 598.950 772.950 601.050 775.050 ;
        RECT 602.250 773.250 603.750 774.150 ;
        RECT 604.950 772.950 607.050 775.050 ;
        RECT 595.950 769.950 598.050 772.050 ;
        RECT 599.250 770.850 600.750 771.750 ;
        RECT 601.950 769.950 604.050 772.050 ;
        RECT 601.950 766.950 604.050 769.050 ;
        RECT 592.950 757.950 595.050 760.050 ;
        RECT 584.400 752.400 588.450 753.450 ;
        RECT 577.950 745.950 580.050 748.050 ;
        RECT 572.400 743.400 576.450 744.450 ;
        RECT 559.950 740.250 561.750 741.150 ;
        RECT 562.950 739.950 565.050 742.050 ;
        RECT 566.250 740.250 568.050 741.150 ;
        RECT 568.950 739.950 571.050 742.050 ;
        RECT 559.950 736.950 562.050 739.050 ;
        RECT 563.250 737.850 564.750 738.750 ;
        RECT 565.950 738.450 568.050 739.050 ;
        RECT 569.400 738.450 570.450 739.950 ;
        RECT 565.950 737.400 570.450 738.450 ;
        RECT 565.950 736.950 568.050 737.400 ;
        RECT 553.950 709.950 556.050 712.050 ;
        RECT 556.950 709.950 559.050 712.050 ;
        RECT 559.950 709.950 562.050 712.050 ;
        RECT 541.950 706.950 544.050 709.050 ;
        RECT 544.950 706.950 547.050 709.050 ;
        RECT 553.950 707.250 556.050 708.150 ;
        RECT 542.400 706.050 543.450 706.950 ;
        RECT 541.950 703.950 544.050 706.050 ;
        RECT 535.950 700.950 538.050 703.050 ;
        RECT 538.950 700.950 541.050 703.050 ;
        RECT 545.400 700.050 546.450 706.950 ;
        RECT 547.950 703.950 550.050 706.050 ;
        RECT 551.250 704.250 552.750 705.150 ;
        RECT 553.950 703.950 556.050 706.050 ;
        RECT 557.250 704.250 559.050 705.150 ;
        RECT 547.950 701.850 549.750 702.750 ;
        RECT 550.950 700.950 553.050 703.050 ;
        RECT 554.400 700.050 555.450 703.950 ;
        RECT 556.950 700.950 559.050 703.050 ;
        RECT 538.950 698.850 541.050 699.750 ;
        RECT 541.950 698.250 544.050 699.150 ;
        RECT 544.950 697.950 547.050 700.050 ;
        RECT 553.950 697.950 556.050 700.050 ;
        RECT 556.950 697.950 559.050 700.050 ;
        RECT 535.950 694.950 538.050 697.050 ;
        RECT 541.950 696.450 544.050 697.050 ;
        RECT 545.400 696.450 546.450 697.950 ;
        RECT 541.950 695.400 546.450 696.450 ;
        RECT 541.950 694.950 544.050 695.400 ;
        RECT 532.950 688.950 535.050 691.050 ;
        RECT 536.400 687.450 537.450 694.950 ;
        RECT 557.400 694.050 558.450 697.950 ;
        RECT 544.950 691.950 547.050 694.050 ;
        RECT 556.950 691.950 559.050 694.050 ;
        RECT 533.400 686.400 537.450 687.450 ;
        RECT 527.400 677.400 531.450 678.450 ;
        RECT 530.400 676.050 531.450 677.400 ;
        RECT 523.950 675.450 526.050 676.050 ;
        RECT 526.950 675.450 529.050 676.050 ;
        RECT 523.950 674.400 529.050 675.450 ;
        RECT 523.950 673.950 526.050 674.400 ;
        RECT 526.950 673.950 529.050 674.400 ;
        RECT 529.950 673.950 532.050 676.050 ;
        RECT 523.950 670.950 526.050 673.050 ;
        RECT 527.250 671.850 528.750 672.750 ;
        RECT 529.950 670.950 532.050 673.050 ;
        RECT 523.950 668.850 526.050 669.750 ;
        RECT 526.950 667.950 529.050 670.050 ;
        RECT 529.950 668.850 532.050 669.750 ;
        RECT 533.400 669.450 534.450 686.400 ;
        RECT 538.950 682.950 541.050 685.050 ;
        RECT 535.950 676.950 538.050 679.050 ;
        RECT 536.400 673.050 537.450 676.950 ;
        RECT 539.400 673.050 540.450 682.950 ;
        RECT 545.400 676.050 546.450 691.950 ;
        RECT 556.950 676.950 559.050 679.050 ;
        RECT 557.400 676.050 558.450 676.950 ;
        RECT 544.950 673.950 547.050 676.050 ;
        RECT 547.950 673.950 550.050 676.050 ;
        RECT 553.950 673.950 556.050 676.050 ;
        RECT 556.950 673.950 559.050 676.050 ;
        RECT 545.400 673.050 546.450 673.950 ;
        RECT 535.950 670.950 538.050 673.050 ;
        RECT 538.950 670.950 541.050 673.050 ;
        RECT 542.250 671.250 543.750 672.150 ;
        RECT 544.950 670.950 547.050 673.050 ;
        RECT 535.950 669.450 538.050 670.050 ;
        RECT 533.400 668.400 538.050 669.450 ;
        RECT 539.250 668.850 540.750 669.750 ;
        RECT 527.400 664.050 528.450 667.950 ;
        RECT 533.400 667.050 534.450 668.400 ;
        RECT 535.950 667.950 538.050 668.400 ;
        RECT 541.950 667.950 544.050 670.050 ;
        RECT 545.250 668.850 547.050 669.750 ;
        RECT 529.950 664.950 532.050 667.050 ;
        RECT 532.950 664.950 535.050 667.050 ;
        RECT 535.950 665.850 538.050 666.750 ;
        RECT 526.950 661.950 529.050 664.050 ;
        RECT 505.950 631.950 508.050 634.050 ;
        RECT 509.250 632.250 510.750 633.150 ;
        RECT 511.950 631.950 514.050 634.050 ;
        RECT 514.950 631.950 517.050 634.050 ;
        RECT 520.950 631.950 523.050 634.050 ;
        RECT 505.950 629.850 507.750 630.750 ;
        RECT 508.950 628.950 511.050 631.050 ;
        RECT 512.250 629.850 514.050 630.750 ;
        RECT 505.950 622.950 508.050 625.050 ;
        RECT 508.950 622.950 511.050 625.050 ;
        RECT 506.400 598.050 507.450 622.950 ;
        RECT 509.400 607.050 510.450 622.950 ;
        RECT 508.950 604.950 511.050 607.050 ;
        RECT 509.400 598.050 510.450 604.950 ;
        RECT 481.950 595.950 484.050 598.050 ;
        RECT 487.950 595.950 490.050 598.050 ;
        RECT 490.950 595.950 493.050 598.050 ;
        RECT 493.950 595.950 496.050 598.050 ;
        RECT 502.950 597.450 505.050 598.050 ;
        RECT 497.250 596.250 499.050 597.150 ;
        RECT 500.400 596.400 505.050 597.450 ;
        RECT 482.400 595.050 483.450 595.950 ;
        RECT 491.400 595.050 492.450 595.950 ;
        RECT 481.950 592.950 484.050 595.050 ;
        RECT 487.950 593.850 489.750 594.750 ;
        RECT 490.950 592.950 493.050 595.050 ;
        RECT 494.250 593.850 495.750 594.750 ;
        RECT 496.950 592.950 499.050 595.050 ;
        RECT 484.950 589.950 487.050 592.050 ;
        RECT 490.950 590.850 493.050 591.750 ;
        RECT 479.400 563.400 483.450 564.450 ;
        RECT 482.400 562.050 483.450 563.400 ;
        RECT 475.950 559.950 478.050 562.050 ;
        RECT 479.250 560.250 480.750 561.150 ;
        RECT 481.950 559.950 484.050 562.050 ;
        RECT 475.950 557.850 477.750 558.750 ;
        RECT 478.950 556.950 481.050 559.050 ;
        RECT 482.250 557.850 484.050 558.750 ;
        RECT 472.950 550.950 475.050 553.050 ;
        RECT 473.400 547.050 474.450 550.950 ;
        RECT 472.950 544.950 475.050 547.050 ;
        RECT 466.950 538.950 469.050 541.050 ;
        RECT 475.950 538.950 478.050 541.050 ;
        RECT 454.950 533.400 457.050 535.500 ;
        RECT 457.950 533.400 460.050 535.500 ;
        RECT 460.950 533.400 463.050 535.500 ;
        RECT 465.750 533.400 467.850 535.500 ;
        RECT 469.950 533.400 472.050 535.500 ;
        RECT 451.950 517.950 454.050 520.050 ;
        RECT 455.550 519.750 456.750 533.400 ;
        RECT 454.950 517.650 457.050 519.750 ;
        RECT 433.950 511.950 436.050 514.050 ;
        RECT 442.950 511.950 445.050 514.050 ;
        RECT 455.550 513.900 456.750 517.650 ;
        RECT 458.250 516.150 459.450 533.400 ;
        RECT 461.400 519.750 462.600 533.400 ;
        RECT 466.350 527.550 467.550 533.400 ;
        RECT 465.750 525.450 467.850 527.550 ;
        RECT 460.950 517.650 463.050 519.750 ;
        RECT 466.350 516.600 467.550 525.450 ;
        RECT 470.550 524.850 471.750 533.400 ;
        RECT 472.950 529.950 475.050 532.050 ;
        RECT 472.950 527.850 475.050 528.750 ;
        RECT 469.950 522.750 472.050 524.850 ;
        RECT 470.550 516.600 471.750 522.750 ;
        RECT 457.950 514.050 460.050 516.150 ;
        RECT 465.900 514.500 468.000 516.600 ;
        RECT 469.950 514.500 472.050 516.600 ;
        RECT 454.800 511.800 456.900 513.900 ;
        RECT 469.950 508.950 472.050 511.050 ;
        RECT 430.950 502.950 433.050 505.050 ;
        RECT 430.950 499.950 433.050 502.050 ;
        RECT 427.950 496.950 430.050 499.050 ;
        RECT 428.400 490.050 429.450 496.950 ;
        RECT 427.950 487.950 430.050 490.050 ;
        RECT 418.950 484.950 421.050 487.050 ;
        RECT 422.250 485.250 423.750 486.150 ;
        RECT 424.950 484.950 427.050 487.050 ;
        RECT 428.250 485.250 430.050 486.150 ;
        RECT 421.950 483.450 424.050 484.050 ;
        RECT 416.400 482.400 424.050 483.450 ;
        RECT 425.250 482.850 426.750 483.750 ;
        RECT 421.950 481.950 424.050 482.400 ;
        RECT 427.950 481.950 430.050 484.050 ;
        RECT 418.950 478.950 421.050 481.050 ;
        RECT 412.950 469.950 415.050 472.050 ;
        RECT 412.950 455.250 414.750 456.150 ;
        RECT 415.950 454.950 418.050 457.050 ;
        RECT 406.950 452.850 409.050 453.750 ;
        RECT 409.950 451.950 412.050 454.050 ;
        RECT 412.950 451.950 415.050 454.050 ;
        RECT 416.250 452.850 418.050 453.750 ;
        RECT 409.950 448.950 412.050 451.050 ;
        RECT 406.950 420.450 409.050 421.050 ;
        RECT 404.400 419.400 409.050 420.450 ;
        RECT 406.950 418.950 409.050 419.400 ;
        RECT 407.400 418.050 408.450 418.950 ;
        RECT 385.950 415.950 388.050 418.050 ;
        RECT 400.950 417.450 403.050 418.050 ;
        RECT 391.950 416.250 394.050 417.150 ;
        RECT 398.400 416.400 403.050 417.450 ;
        RECT 386.400 415.050 387.450 415.950 ;
        RECT 382.950 413.250 384.750 414.150 ;
        RECT 385.950 412.950 388.050 415.050 ;
        RECT 389.250 413.250 390.750 414.150 ;
        RECT 391.950 412.950 394.050 415.050 ;
        RECT 382.950 409.950 385.050 412.050 ;
        RECT 386.250 410.850 387.750 411.750 ;
        RECT 388.950 409.950 391.050 412.050 ;
        RECT 380.400 407.400 384.450 408.450 ;
        RECT 373.950 388.950 376.050 391.050 ;
        RECT 376.950 385.950 379.050 388.050 ;
        RECT 367.950 382.950 370.050 385.050 ;
        RECT 370.950 382.950 373.050 385.050 ;
        RECT 374.250 383.250 376.050 384.150 ;
        RECT 376.950 383.850 379.050 384.750 ;
        RECT 379.950 383.250 382.050 384.150 ;
        RECT 334.950 380.850 337.050 381.750 ;
        RECT 340.950 380.850 343.050 381.750 ;
        RECT 352.950 380.850 355.050 381.750 ;
        RECT 358.950 380.850 361.050 381.750 ;
        RECT 361.950 379.950 364.050 382.050 ;
        RECT 331.950 355.950 334.050 358.050 ;
        RECT 340.950 346.950 343.050 349.050 ;
        RECT 368.400 348.450 369.450 382.950 ;
        RECT 383.400 382.050 384.450 407.400 ;
        RECT 385.950 406.950 388.050 409.050 ;
        RECT 386.400 387.450 387.450 406.950 ;
        RECT 389.400 397.050 390.450 409.950 ;
        RECT 392.400 406.050 393.450 412.950 ;
        RECT 391.950 403.950 394.050 406.050 ;
        RECT 388.950 394.950 391.050 397.050 ;
        RECT 398.400 391.050 399.450 416.400 ;
        RECT 400.950 415.950 403.050 416.400 ;
        RECT 404.250 416.250 405.750 417.150 ;
        RECT 406.950 415.950 409.050 418.050 ;
        RECT 400.950 413.850 402.750 414.750 ;
        RECT 403.950 412.950 406.050 415.050 ;
        RECT 407.250 413.850 409.050 414.750 ;
        RECT 404.400 406.050 405.450 412.950 ;
        RECT 403.950 403.950 406.050 406.050 ;
        RECT 410.400 394.050 411.450 448.950 ;
        RECT 415.950 442.950 418.050 445.050 ;
        RECT 416.400 439.050 417.450 442.950 ;
        RECT 415.950 436.950 418.050 439.050 ;
        RECT 412.950 418.950 415.050 421.050 ;
        RECT 413.400 415.050 414.450 418.950 ;
        RECT 412.950 412.950 415.050 415.050 ;
        RECT 412.950 410.850 415.050 411.750 ;
        RECT 415.950 410.250 418.050 411.150 ;
        RECT 415.950 406.950 418.050 409.050 ;
        RECT 416.400 402.450 417.450 406.950 ;
        RECT 413.400 401.400 417.450 402.450 ;
        RECT 409.950 391.950 412.050 394.050 ;
        RECT 391.950 388.950 394.050 391.050 ;
        RECT 397.950 388.950 400.050 391.050 ;
        RECT 392.400 388.050 393.450 388.950 ;
        RECT 386.400 386.400 390.450 387.450 ;
        RECT 370.950 380.850 372.750 381.750 ;
        RECT 373.950 379.950 376.050 382.050 ;
        RECT 376.950 379.950 379.050 382.050 ;
        RECT 379.950 379.950 382.050 382.050 ;
        RECT 382.950 379.950 385.050 382.050 ;
        RECT 373.950 364.950 376.050 367.050 ;
        RECT 368.400 347.400 372.450 348.450 ;
        RECT 334.950 342.450 337.050 343.050 ;
        RECT 331.950 341.250 333.750 342.150 ;
        RECT 334.950 341.400 339.450 342.450 ;
        RECT 334.950 340.950 337.050 341.400 ;
        RECT 331.950 337.950 334.050 340.050 ;
        RECT 335.250 338.850 337.050 339.750 ;
        RECT 325.950 316.950 328.050 319.050 ;
        RECT 319.950 313.950 322.050 316.050 ;
        RECT 325.950 313.950 328.050 316.050 ;
        RECT 313.950 310.950 316.050 313.050 ;
        RECT 317.250 311.250 319.050 312.150 ;
        RECT 319.950 311.850 322.050 312.750 ;
        RECT 322.950 311.250 325.050 312.150 ;
        RECT 310.950 307.950 313.050 310.050 ;
        RECT 313.950 308.850 315.750 309.750 ;
        RECT 316.950 307.950 319.050 310.050 ;
        RECT 322.950 307.950 325.050 310.050 ;
        RECT 313.950 301.950 316.050 304.050 ;
        RECT 308.400 272.400 312.450 273.450 ;
        RECT 311.400 271.050 312.450 272.400 ;
        RECT 298.950 268.950 301.050 271.050 ;
        RECT 301.950 268.950 304.050 271.050 ;
        RECT 304.950 268.950 307.050 271.050 ;
        RECT 308.250 269.250 310.050 270.150 ;
        RECT 310.950 268.950 313.050 271.050 ;
        RECT 311.400 268.050 312.450 268.950 ;
        RECT 298.950 266.850 301.050 267.750 ;
        RECT 301.950 266.250 304.050 267.150 ;
        RECT 304.950 266.850 306.750 267.750 ;
        RECT 307.950 265.950 310.050 268.050 ;
        RECT 310.950 265.950 313.050 268.050 ;
        RECT 308.400 265.050 309.450 265.950 ;
        RECT 301.950 262.950 304.050 265.050 ;
        RECT 307.950 262.950 310.050 265.050 ;
        RECT 302.400 262.050 303.450 262.950 ;
        RECT 301.950 259.950 304.050 262.050 ;
        RECT 307.950 259.950 310.050 262.050 ;
        RECT 301.950 238.950 304.050 241.050 ;
        RECT 302.400 238.050 303.450 238.950 ;
        RECT 298.950 236.250 300.750 237.150 ;
        RECT 301.950 235.950 304.050 238.050 ;
        RECT 305.250 236.250 307.050 237.150 ;
        RECT 286.950 232.950 289.050 233.400 ;
        RECT 292.950 233.400 297.450 234.450 ;
        RECT 292.950 232.950 295.050 233.400 ;
        RECT 298.950 232.950 301.050 235.050 ;
        RECT 302.250 233.850 303.750 234.750 ;
        RECT 304.950 232.950 307.050 235.050 ;
        RECT 277.950 217.950 280.050 220.050 ;
        RECT 277.950 199.950 280.050 202.050 ;
        RECT 278.400 199.050 279.450 199.950 ;
        RECT 281.400 199.050 282.450 232.950 ;
        RECT 286.950 214.950 289.050 217.050 ;
        RECT 283.950 199.950 286.050 202.050 ;
        RECT 277.950 196.950 280.050 199.050 ;
        RECT 280.950 196.950 283.050 199.050 ;
        RECT 277.950 194.850 280.050 195.750 ;
        RECT 280.950 194.250 283.050 195.150 ;
        RECT 280.950 190.950 283.050 193.050 ;
        RECT 284.400 172.050 285.450 199.950 ;
        RECT 287.400 196.050 288.450 214.950 ;
        RECT 293.400 205.050 294.450 232.950 ;
        RECT 298.950 226.950 301.050 229.050 ;
        RECT 295.950 205.950 298.050 208.050 ;
        RECT 292.950 202.950 295.050 205.050 ;
        RECT 296.400 202.050 297.450 205.950 ;
        RECT 289.950 199.950 292.050 202.050 ;
        RECT 293.250 200.250 294.750 201.150 ;
        RECT 295.950 199.950 298.050 202.050 ;
        RECT 289.950 197.850 291.750 198.750 ;
        RECT 292.950 196.950 295.050 199.050 ;
        RECT 296.250 197.850 298.050 198.750 ;
        RECT 286.950 193.950 289.050 196.050 ;
        RECT 286.950 190.950 289.050 193.050 ;
        RECT 283.950 169.950 286.050 172.050 ;
        RECT 272.400 167.400 276.450 168.450 ;
        RECT 262.950 164.850 265.050 165.750 ;
        RECT 268.950 164.850 271.050 165.750 ;
        RECT 272.400 145.050 273.450 167.400 ;
        RECT 277.950 166.950 280.050 169.050 ;
        RECT 278.400 166.050 279.450 166.950 ;
        RECT 274.950 164.250 276.750 165.150 ;
        RECT 277.950 163.950 280.050 166.050 ;
        RECT 281.250 164.250 283.050 165.150 ;
        RECT 274.950 160.950 277.050 163.050 ;
        RECT 278.250 161.850 279.750 162.750 ;
        RECT 280.950 160.950 283.050 163.050 ;
        RECT 287.400 162.450 288.450 190.950 ;
        RECT 299.400 178.050 300.450 226.950 ;
        RECT 301.950 205.950 304.050 208.050 ;
        RECT 302.400 202.050 303.450 205.950 ;
        RECT 305.400 205.050 306.450 232.950 ;
        RECT 308.400 232.050 309.450 259.950 ;
        RECT 311.400 244.050 312.450 265.950 ;
        RECT 310.950 241.950 313.050 244.050 ;
        RECT 314.400 240.450 315.450 301.950 ;
        RECT 323.400 301.050 324.450 307.950 ;
        RECT 326.400 304.050 327.450 313.950 ;
        RECT 332.400 313.050 333.450 337.950 ;
        RECT 338.400 334.050 339.450 341.400 ;
        RECT 337.950 331.950 340.050 334.050 ;
        RECT 334.950 319.950 337.050 322.050 ;
        RECT 328.950 310.950 331.050 313.050 ;
        RECT 331.950 310.950 334.050 313.050 ;
        RECT 325.950 301.950 328.050 304.050 ;
        RECT 319.950 298.950 322.050 301.050 ;
        RECT 322.950 298.950 325.050 301.050 ;
        RECT 320.400 271.050 321.450 298.950 ;
        RECT 323.400 274.050 324.450 298.950 ;
        RECT 326.400 283.050 327.450 301.950 ;
        RECT 325.950 280.950 328.050 283.050 ;
        RECT 322.950 271.950 325.050 274.050 ;
        RECT 325.950 272.250 328.050 273.150 ;
        RECT 316.950 269.250 318.750 270.150 ;
        RECT 319.950 268.950 322.050 271.050 ;
        RECT 323.250 269.250 324.750 270.150 ;
        RECT 325.950 268.950 328.050 271.050 ;
        RECT 316.950 265.950 319.050 268.050 ;
        RECT 320.250 266.850 321.750 267.750 ;
        RECT 322.950 265.950 325.050 268.050 ;
        RECT 316.950 256.950 319.050 259.050 ;
        RECT 311.400 239.400 315.450 240.450 ;
        RECT 311.400 235.050 312.450 239.400 ;
        RECT 313.950 236.250 316.050 237.150 ;
        RECT 310.950 232.950 313.050 235.050 ;
        RECT 313.950 232.950 316.050 235.050 ;
        RECT 307.950 229.950 310.050 232.050 ;
        RECT 313.950 229.950 316.050 232.050 ;
        RECT 304.950 202.950 307.050 205.050 ;
        RECT 307.950 203.250 310.050 204.150 ;
        RECT 314.400 202.050 315.450 229.950 ;
        RECT 317.400 229.050 318.450 256.950 ;
        RECT 319.950 233.850 322.050 234.750 ;
        RECT 319.950 229.950 322.050 232.050 ;
        RECT 316.950 226.950 319.050 229.050 ;
        RECT 316.950 217.950 319.050 220.050 ;
        RECT 301.950 199.950 304.050 202.050 ;
        RECT 305.250 200.250 306.750 201.150 ;
        RECT 307.950 199.950 310.050 202.050 ;
        RECT 311.250 200.250 313.050 201.150 ;
        RECT 313.950 199.950 316.050 202.050 ;
        RECT 301.950 197.850 303.750 198.750 ;
        RECT 304.950 196.950 307.050 199.050 ;
        RECT 307.950 196.950 310.050 199.050 ;
        RECT 310.950 198.450 313.050 199.050 ;
        RECT 310.950 197.400 315.450 198.450 ;
        RECT 310.950 196.950 313.050 197.400 ;
        RECT 305.400 196.050 306.450 196.950 ;
        RECT 304.950 193.950 307.050 196.050 ;
        RECT 304.950 181.950 307.050 184.050 ;
        RECT 298.950 175.950 301.050 178.050 ;
        RECT 298.950 169.950 301.050 172.050 ;
        RECT 299.400 169.050 300.450 169.950 ;
        RECT 292.950 168.450 295.050 169.050 ;
        RECT 284.400 161.400 288.450 162.450 ;
        RECT 290.400 167.400 295.050 168.450 ;
        RECT 271.950 142.950 274.050 145.050 ;
        RECT 259.950 133.950 262.050 136.050 ;
        RECT 256.950 130.950 259.050 133.050 ;
        RECT 260.400 130.050 261.450 133.950 ;
        RECT 275.400 133.050 276.450 160.950 ;
        RECT 277.950 157.950 280.050 160.050 ;
        RECT 265.950 130.950 268.050 133.050 ;
        RECT 274.950 130.950 277.050 133.050 ;
        RECT 241.950 129.450 244.050 130.050 ;
        RECT 239.400 128.400 244.050 129.450 ;
        RECT 239.400 124.050 240.450 128.400 ;
        RECT 241.950 127.950 244.050 128.400 ;
        RECT 245.250 128.250 246.750 129.150 ;
        RECT 247.950 127.950 250.050 130.050 ;
        RECT 253.950 129.450 256.050 130.050 ;
        RECT 251.400 128.400 256.050 129.450 ;
        RECT 241.950 125.850 243.750 126.750 ;
        RECT 244.950 124.950 247.050 127.050 ;
        RECT 248.250 125.850 250.050 126.750 ;
        RECT 238.950 121.950 241.050 124.050 ;
        RECT 251.400 123.450 252.450 128.400 ;
        RECT 253.950 127.950 256.050 128.400 ;
        RECT 257.250 128.250 258.750 129.150 ;
        RECT 259.950 127.950 262.050 130.050 ;
        RECT 253.950 125.850 255.750 126.750 ;
        RECT 256.950 124.950 259.050 127.050 ;
        RECT 260.250 125.850 262.050 126.750 ;
        RECT 251.400 122.400 255.450 123.450 ;
        RECT 235.950 109.950 238.050 112.050 ;
        RECT 235.950 103.950 238.050 106.050 ;
        RECT 232.950 100.950 235.050 103.050 ;
        RECT 208.950 95.250 211.050 96.150 ;
        RECT 211.950 95.850 214.050 96.750 ;
        RECT 214.950 95.250 216.750 96.150 ;
        RECT 217.950 94.950 220.050 97.050 ;
        RECT 236.400 94.050 237.450 103.950 ;
        RECT 254.400 94.050 255.450 122.400 ;
        RECT 262.950 121.950 265.050 124.050 ;
        RECT 263.400 94.050 264.450 121.950 ;
        RECT 266.400 118.050 267.450 130.950 ;
        RECT 278.400 130.050 279.450 157.950 ;
        RECT 284.400 133.050 285.450 161.400 ;
        RECT 290.400 154.050 291.450 167.400 ;
        RECT 292.950 166.950 295.050 167.400 ;
        RECT 296.250 167.250 297.750 168.150 ;
        RECT 298.950 166.950 301.050 169.050 ;
        RECT 292.950 164.850 294.750 165.750 ;
        RECT 295.950 163.950 298.050 166.050 ;
        RECT 299.250 164.850 300.750 165.750 ;
        RECT 301.950 163.950 304.050 166.050 ;
        RECT 301.950 161.850 304.050 162.750 ;
        RECT 289.950 151.950 292.050 154.050 ;
        RECT 305.400 145.050 306.450 181.950 ;
        RECT 304.950 142.950 307.050 145.050 ;
        RECT 308.400 136.050 309.450 196.950 ;
        RECT 310.950 193.950 313.050 196.050 ;
        RECT 311.400 172.050 312.450 193.950 ;
        RECT 314.400 193.050 315.450 197.400 ;
        RECT 313.950 190.950 316.050 193.050 ;
        RECT 310.950 169.950 313.050 172.050 ;
        RECT 317.400 169.050 318.450 217.950 ;
        RECT 320.400 214.050 321.450 229.950 ;
        RECT 319.950 211.950 322.050 214.050 ;
        RECT 323.400 211.050 324.450 265.950 ;
        RECT 326.400 256.050 327.450 268.950 ;
        RECT 325.950 253.950 328.050 256.050 ;
        RECT 329.400 250.050 330.450 310.950 ;
        RECT 335.400 310.050 336.450 319.950 ;
        RECT 331.950 308.250 333.750 309.150 ;
        RECT 334.950 307.950 337.050 310.050 ;
        RECT 338.250 308.250 340.050 309.150 ;
        RECT 331.950 304.950 334.050 307.050 ;
        RECT 335.250 305.850 336.750 306.750 ;
        RECT 337.950 304.950 340.050 307.050 ;
        RECT 332.400 250.050 333.450 304.950 ;
        RECT 337.950 283.950 340.050 286.050 ;
        RECT 338.400 271.050 339.450 283.950 ;
        RECT 341.400 277.050 342.450 346.950 ;
        RECT 352.950 343.950 355.050 346.050 ;
        RECT 355.950 343.950 358.050 346.050 ;
        RECT 367.950 344.250 370.050 345.150 ;
        RECT 353.400 343.050 354.450 343.950 ;
        RECT 343.950 341.250 345.750 342.150 ;
        RECT 346.950 340.950 349.050 343.050 ;
        RECT 352.950 340.950 355.050 343.050 ;
        RECT 343.950 337.950 346.050 340.050 ;
        RECT 347.250 338.850 349.050 339.750 ;
        RECT 349.950 338.250 352.050 339.150 ;
        RECT 352.950 338.850 355.050 339.750 ;
        RECT 356.400 339.450 357.450 343.950 ;
        RECT 358.950 341.250 360.750 342.150 ;
        RECT 361.950 340.950 364.050 343.050 ;
        RECT 365.250 341.250 366.750 342.150 ;
        RECT 367.950 340.950 370.050 343.050 ;
        RECT 368.400 340.050 369.450 340.950 ;
        RECT 358.950 339.450 361.050 340.050 ;
        RECT 356.400 338.400 361.050 339.450 ;
        RECT 362.250 338.850 363.750 339.750 ;
        RECT 346.950 334.950 349.050 337.050 ;
        RECT 349.950 334.950 352.050 337.050 ;
        RECT 347.400 331.050 348.450 334.950 ;
        RECT 346.950 328.950 349.050 331.050 ;
        RECT 346.950 308.250 348.750 309.150 ;
        RECT 349.950 307.950 352.050 310.050 ;
        RECT 353.250 308.250 355.050 309.150 ;
        RECT 346.950 304.950 349.050 307.050 ;
        RECT 350.250 305.850 351.750 306.750 ;
        RECT 352.950 304.950 355.050 307.050 ;
        RECT 347.400 301.050 348.450 304.950 ;
        RECT 353.400 304.050 354.450 304.950 ;
        RECT 352.950 301.950 355.050 304.050 ;
        RECT 346.950 298.950 349.050 301.050 ;
        RECT 356.400 283.050 357.450 338.400 ;
        RECT 358.950 337.950 361.050 338.400 ;
        RECT 364.950 337.950 367.050 340.050 ;
        RECT 367.950 337.950 370.050 340.050 ;
        RECT 365.400 331.050 366.450 337.950 ;
        RECT 364.950 328.950 367.050 331.050 ;
        RECT 367.950 328.950 370.050 331.050 ;
        RECT 364.950 325.950 367.050 328.050 ;
        RECT 358.950 319.950 361.050 322.050 ;
        RECT 359.400 286.050 360.450 319.950 ;
        RECT 361.950 313.950 364.050 316.050 ;
        RECT 362.400 310.050 363.450 313.950 ;
        RECT 365.400 313.050 366.450 325.950 ;
        RECT 368.400 316.050 369.450 328.950 ;
        RECT 371.400 328.050 372.450 347.400 ;
        RECT 374.400 337.050 375.450 364.950 ;
        RECT 373.950 334.950 376.050 337.050 ;
        RECT 377.400 334.050 378.450 379.950 ;
        RECT 380.400 367.050 381.450 379.950 ;
        RECT 379.950 364.950 382.050 367.050 ;
        RECT 382.950 364.950 385.050 367.050 ;
        RECT 383.400 346.050 384.450 364.950 ;
        RECT 386.400 361.050 387.450 386.400 ;
        RECT 389.400 385.050 390.450 386.400 ;
        RECT 391.950 385.950 394.050 388.050 ;
        RECT 397.950 385.950 400.050 388.050 ;
        RECT 388.950 382.950 391.050 385.050 ;
        RECT 392.250 383.850 393.750 384.750 ;
        RECT 394.950 382.950 397.050 385.050 ;
        RECT 388.950 380.850 391.050 381.750 ;
        RECT 394.950 380.850 397.050 381.750 ;
        RECT 394.950 376.950 397.050 379.050 ;
        RECT 391.950 370.950 394.050 373.050 ;
        RECT 385.950 358.950 388.050 361.050 ;
        RECT 385.950 355.950 388.050 358.050 ;
        RECT 382.950 343.950 385.050 346.050 ;
        RECT 379.950 341.250 382.050 342.150 ;
        RECT 382.950 341.850 385.050 342.750 ;
        RECT 379.950 337.950 382.050 340.050 ;
        RECT 376.950 331.950 379.050 334.050 ;
        RECT 380.400 331.050 381.450 337.950 ;
        RECT 379.950 328.950 382.050 331.050 ;
        RECT 382.950 328.950 385.050 331.050 ;
        RECT 370.950 325.950 373.050 328.050 ;
        RECT 376.950 325.950 379.050 328.050 ;
        RECT 379.950 325.950 382.050 328.050 ;
        RECT 367.950 313.950 370.050 316.050 ;
        RECT 370.950 313.950 373.050 316.050 ;
        RECT 373.950 313.950 376.050 316.050 ;
        RECT 371.400 313.050 372.450 313.950 ;
        RECT 364.950 310.950 367.050 313.050 ;
        RECT 368.250 311.250 369.750 312.150 ;
        RECT 370.950 310.950 373.050 313.050 ;
        RECT 361.950 307.950 364.050 310.050 ;
        RECT 365.250 308.850 366.750 309.750 ;
        RECT 367.950 307.950 370.050 310.050 ;
        RECT 371.250 308.850 373.050 309.750 ;
        RECT 368.400 307.050 369.450 307.950 ;
        RECT 361.950 305.850 364.050 306.750 ;
        RECT 367.950 304.950 370.050 307.050 ;
        RECT 368.400 304.050 369.450 304.950 ;
        RECT 374.400 304.050 375.450 313.950 ;
        RECT 361.950 301.950 364.050 304.050 ;
        RECT 367.950 301.950 370.050 304.050 ;
        RECT 373.950 301.950 376.050 304.050 ;
        RECT 358.950 283.950 361.050 286.050 ;
        RECT 355.950 280.950 358.050 283.050 ;
        RECT 340.950 274.950 343.050 277.050 ;
        RECT 346.950 274.950 349.050 277.050 ;
        RECT 349.950 274.950 352.050 277.050 ;
        RECT 352.950 274.950 355.050 277.050 ;
        RECT 343.950 272.250 346.050 273.150 ;
        RECT 334.950 269.250 336.750 270.150 ;
        RECT 337.950 268.950 340.050 271.050 ;
        RECT 341.250 269.250 342.750 270.150 ;
        RECT 343.950 268.950 346.050 271.050 ;
        RECT 347.400 268.050 348.450 274.950 ;
        RECT 334.950 265.950 337.050 268.050 ;
        RECT 338.250 266.850 339.750 267.750 ;
        RECT 340.950 267.450 343.050 268.050 ;
        RECT 343.950 267.450 346.050 268.050 ;
        RECT 340.950 266.400 346.050 267.450 ;
        RECT 340.950 265.950 343.050 266.400 ;
        RECT 343.950 265.950 346.050 266.400 ;
        RECT 346.950 265.950 349.050 268.050 ;
        RECT 350.400 261.450 351.450 274.950 ;
        RECT 353.400 274.050 354.450 274.950 ;
        RECT 352.950 271.950 355.050 274.050 ;
        RECT 356.250 272.250 357.750 273.150 ;
        RECT 358.950 271.950 361.050 274.050 ;
        RECT 352.950 269.850 354.750 270.750 ;
        RECT 355.950 268.950 358.050 271.050 ;
        RECT 359.250 269.850 361.050 270.750 ;
        RECT 358.950 262.950 361.050 265.050 ;
        RECT 352.950 261.450 355.050 262.050 ;
        RECT 350.400 260.400 355.050 261.450 ;
        RECT 352.950 259.950 355.050 260.400 ;
        RECT 346.950 256.950 349.050 259.050 ;
        RECT 347.400 253.050 348.450 256.950 ;
        RECT 346.950 250.950 349.050 253.050 ;
        RECT 328.950 247.950 331.050 250.050 ;
        RECT 331.950 247.950 334.050 250.050 ;
        RECT 325.950 244.950 328.050 247.050 ;
        RECT 328.950 244.950 331.050 247.050 ;
        RECT 331.950 244.950 334.050 247.050 ;
        RECT 340.950 245.400 343.050 247.500 ;
        RECT 345.150 245.400 347.250 247.500 ;
        RECT 349.950 245.400 352.050 247.500 ;
        RECT 352.950 245.400 355.050 247.500 ;
        RECT 355.950 245.400 358.050 247.500 ;
        RECT 326.550 226.050 327.750 244.950 ;
        RECT 329.550 232.350 330.750 244.950 ;
        RECT 328.950 230.250 331.050 232.350 ;
        RECT 329.550 226.050 330.750 230.250 ;
        RECT 332.550 226.050 333.750 244.950 ;
        RECT 337.950 241.950 340.050 244.050 ;
        RECT 337.950 239.850 340.050 240.750 ;
        RECT 337.950 235.950 340.050 238.050 ;
        RECT 341.250 236.850 342.450 245.400 ;
        RECT 345.450 239.550 346.650 245.400 ;
        RECT 345.150 237.450 347.250 239.550 ;
        RECT 325.950 223.950 328.050 226.050 ;
        RECT 328.950 223.950 331.050 226.050 ;
        RECT 331.950 223.950 334.050 226.050 ;
        RECT 331.950 214.950 334.050 217.050 ;
        RECT 322.950 208.950 325.050 211.050 ;
        RECT 322.950 201.450 325.050 202.050 ;
        RECT 322.950 200.400 327.450 201.450 ;
        RECT 322.950 199.950 325.050 200.400 ;
        RECT 326.400 199.050 327.450 200.400 ;
        RECT 319.950 197.250 322.050 198.150 ;
        RECT 322.950 197.850 325.050 198.750 ;
        RECT 325.950 196.950 328.050 199.050 ;
        RECT 328.950 197.250 331.050 198.150 ;
        RECT 319.950 193.950 322.050 196.050 ;
        RECT 319.950 190.950 322.050 193.050 ;
        RECT 320.400 172.050 321.450 190.950 ;
        RECT 326.400 172.050 327.450 196.950 ;
        RECT 328.950 193.950 331.050 196.050 ;
        RECT 319.950 169.950 322.050 172.050 ;
        RECT 325.950 171.450 328.050 172.050 ;
        RECT 323.400 170.400 328.050 171.450 ;
        RECT 310.950 166.950 313.050 169.050 ;
        RECT 316.950 166.950 319.050 169.050 ;
        RECT 311.400 160.050 312.450 166.950 ;
        RECT 313.950 164.250 315.750 165.150 ;
        RECT 316.950 163.950 319.050 166.050 ;
        RECT 320.250 164.250 322.050 165.150 ;
        RECT 313.950 160.950 316.050 163.050 ;
        RECT 317.250 161.850 318.750 162.750 ;
        RECT 319.950 160.950 322.050 163.050 ;
        RECT 320.400 160.050 321.450 160.950 ;
        RECT 310.950 157.950 313.050 160.050 ;
        RECT 313.950 157.950 316.050 160.050 ;
        RECT 319.950 157.950 322.050 160.050 ;
        RECT 289.950 133.950 292.050 136.050 ;
        RECT 307.950 133.950 310.050 136.050 ;
        RECT 283.950 130.950 286.050 133.050 ;
        RECT 290.400 130.050 291.450 133.950 ;
        RECT 292.950 130.950 295.050 133.050 ;
        RECT 271.950 129.450 274.050 130.050 ;
        RECT 269.400 128.400 274.050 129.450 ;
        RECT 265.950 115.950 268.050 118.050 ;
        RECT 205.950 91.950 208.050 94.050 ;
        RECT 208.950 91.950 211.050 94.050 ;
        RECT 214.950 91.950 217.050 94.050 ;
        RECT 218.250 92.850 220.050 93.750 ;
        RECT 232.950 92.250 234.750 93.150 ;
        RECT 235.950 91.950 238.050 94.050 ;
        RECT 239.250 92.250 241.050 93.150 ;
        RECT 244.950 92.250 246.750 93.150 ;
        RECT 247.950 91.950 250.050 94.050 ;
        RECT 250.950 91.950 253.050 94.050 ;
        RECT 253.950 93.450 256.050 94.050 ;
        RECT 253.950 92.400 258.450 93.450 ;
        RECT 253.950 91.950 256.050 92.400 ;
        RECT 206.400 58.050 207.450 91.950 ;
        RECT 209.400 85.050 210.450 91.950 ;
        RECT 215.400 85.050 216.450 91.950 ;
        RECT 251.400 91.050 252.450 91.950 ;
        RECT 220.950 88.950 223.050 91.050 ;
        RECT 232.950 88.950 235.050 91.050 ;
        RECT 236.250 89.850 237.750 90.750 ;
        RECT 238.950 88.950 241.050 91.050 ;
        RECT 244.950 88.950 247.050 91.050 ;
        RECT 248.250 89.850 249.750 90.750 ;
        RECT 250.950 88.950 253.050 91.050 ;
        RECT 254.250 89.850 256.050 90.750 ;
        RECT 208.950 82.950 211.050 85.050 ;
        RECT 214.950 82.950 217.050 85.050 ;
        RECT 205.950 55.950 208.050 58.050 ;
        RECT 211.950 57.450 214.050 58.050 ;
        RECT 209.250 56.250 210.750 57.150 ;
        RECT 211.950 56.400 216.450 57.450 ;
        RECT 211.950 55.950 214.050 56.400 ;
        RECT 215.400 55.050 216.450 56.400 ;
        RECT 217.950 55.950 220.050 58.050 ;
        RECT 181.950 53.250 184.050 54.150 ;
        RECT 187.950 53.250 190.050 54.150 ;
        RECT 193.950 53.250 196.050 54.150 ;
        RECT 199.950 53.250 202.050 54.150 ;
        RECT 202.950 52.950 205.050 55.050 ;
        RECT 205.950 53.850 207.750 54.750 ;
        RECT 208.950 52.950 211.050 55.050 ;
        RECT 212.250 53.850 214.050 54.750 ;
        RECT 214.950 52.950 217.050 55.050 ;
        RECT 166.950 50.250 169.050 51.150 ;
        RECT 169.950 50.850 172.050 51.750 ;
        RECT 172.950 49.950 175.050 52.050 ;
        RECT 178.950 49.950 181.050 52.050 ;
        RECT 181.950 49.950 184.050 52.050 ;
        RECT 185.250 50.250 186.750 51.150 ;
        RECT 187.950 49.950 190.050 52.050 ;
        RECT 193.950 49.950 196.050 52.050 ;
        RECT 197.250 50.250 198.750 51.150 ;
        RECT 199.950 49.950 202.050 52.050 ;
        RECT 182.400 49.050 183.450 49.950 ;
        RECT 142.950 46.950 145.050 49.050 ;
        RECT 145.950 46.950 148.050 49.050 ;
        RECT 163.950 46.950 166.050 49.050 ;
        RECT 166.950 46.950 169.050 49.050 ;
        RECT 172.950 46.950 175.050 49.050 ;
        RECT 181.950 46.950 184.050 49.050 ;
        RECT 184.950 46.950 187.050 49.050 ;
        RECT 133.950 43.950 136.050 46.050 ;
        RECT 139.950 43.950 142.050 46.050 ;
        RECT 127.950 31.950 130.050 34.050 ;
        RECT 128.400 31.050 129.450 31.950 ;
        RECT 127.950 28.950 130.050 31.050 ;
        RECT 140.400 28.050 141.450 43.950 ;
        RECT 143.400 40.050 144.450 46.950 ;
        RECT 142.950 37.950 145.050 40.050 ;
        RECT 124.950 25.950 127.050 28.050 ;
        RECT 136.950 25.950 139.050 28.050 ;
        RECT 139.950 25.950 142.050 28.050 ;
        RECT 137.400 25.050 138.450 25.950 ;
        RECT 91.950 22.950 94.050 25.050 ;
        RECT 103.950 22.950 106.050 25.050 ;
        RECT 106.950 22.950 109.050 25.050 ;
        RECT 110.250 23.250 111.750 24.150 ;
        RECT 112.950 22.950 115.050 25.050 ;
        RECT 115.950 22.950 118.050 25.050 ;
        RECT 121.950 24.450 124.050 25.050 ;
        RECT 124.950 24.450 127.050 25.050 ;
        RECT 119.250 23.250 120.750 24.150 ;
        RECT 121.950 23.400 127.050 24.450 ;
        RECT 121.950 22.950 124.050 23.400 ;
        RECT 124.950 22.950 127.050 23.400 ;
        RECT 127.950 22.950 130.050 25.050 ;
        RECT 130.950 22.950 133.050 25.050 ;
        RECT 136.950 22.950 139.050 25.050 ;
        RECT 140.250 23.250 141.750 24.150 ;
        RECT 142.950 22.950 145.050 25.050 ;
        RECT 92.400 22.050 93.450 22.950 ;
        RECT 104.400 22.050 105.450 22.950 ;
        RECT 88.950 20.250 90.750 21.150 ;
        RECT 91.950 19.950 94.050 22.050 ;
        RECT 95.250 20.250 97.050 21.150 ;
        RECT 103.950 19.950 106.050 22.050 ;
        RECT 107.250 20.850 108.750 21.750 ;
        RECT 109.950 19.950 112.050 22.050 ;
        RECT 113.250 20.850 115.050 21.750 ;
        RECT 115.950 20.850 117.750 21.750 ;
        RECT 118.950 19.950 121.050 22.050 ;
        RECT 122.250 20.850 123.750 21.750 ;
        RECT 124.950 19.950 127.050 22.050 ;
        RECT 85.950 18.450 88.050 19.050 ;
        RECT 88.950 18.450 91.050 19.050 ;
        RECT 85.950 17.400 91.050 18.450 ;
        RECT 92.250 17.850 93.750 18.750 ;
        RECT 85.950 16.950 88.050 17.400 ;
        RECT 88.950 16.950 91.050 17.400 ;
        RECT 94.950 16.950 97.050 19.050 ;
        RECT 103.950 17.850 106.050 18.750 ;
        RECT 95.400 16.050 96.450 16.950 ;
        RECT 46.950 13.650 49.050 15.750 ;
        RECT 52.950 13.950 55.050 16.050 ;
        RECT 73.950 13.950 76.050 16.050 ;
        RECT 94.950 13.950 97.050 16.050 ;
        RECT 43.950 10.050 46.050 12.150 ;
        RECT 4.950 7.950 7.050 10.050 ;
        RECT 16.950 7.950 19.050 10.050 ;
        RECT 19.950 7.950 22.050 10.050 ;
        RECT 22.950 7.950 25.050 10.050 ;
        RECT 47.250 9.900 48.450 13.650 ;
        RECT 110.400 13.050 111.450 19.950 ;
        RECT 119.400 16.050 120.450 19.950 ;
        RECT 128.400 19.050 129.450 22.950 ;
        RECT 124.950 17.850 127.050 18.750 ;
        RECT 127.950 16.950 130.050 19.050 ;
        RECT 118.950 13.950 121.050 16.050 ;
        RECT 131.400 13.050 132.450 22.950 ;
        RECT 146.400 22.050 147.450 46.950 ;
        RECT 167.400 40.050 168.450 46.950 ;
        RECT 173.400 40.050 174.450 46.950 ;
        RECT 166.950 37.950 169.050 40.050 ;
        RECT 172.950 37.950 175.050 40.050 ;
        RECT 167.400 37.050 168.450 37.950 ;
        RECT 166.950 34.950 169.050 37.050 ;
        RECT 166.950 31.950 169.050 34.050 ;
        RECT 163.950 25.950 166.050 28.050 ;
        RECT 160.950 23.250 163.050 24.150 ;
        RECT 163.950 23.850 166.050 24.750 ;
        RECT 167.400 22.050 168.450 31.950 ;
        RECT 173.400 28.050 174.450 37.950 ;
        RECT 185.400 28.050 186.450 46.950 ;
        RECT 194.400 31.050 195.450 49.950 ;
        RECT 215.400 49.050 216.450 52.950 ;
        RECT 218.400 52.050 219.450 55.950 ;
        RECT 221.400 55.050 222.450 88.950 ;
        RECT 233.400 88.050 234.450 88.950 ;
        RECT 232.950 85.950 235.050 88.050 ;
        RECT 250.950 86.850 253.050 87.750 ;
        RECT 257.400 82.050 258.450 92.400 ;
        RECT 259.950 92.250 261.750 93.150 ;
        RECT 262.950 91.950 265.050 94.050 ;
        RECT 266.250 92.250 268.050 93.150 ;
        RECT 259.950 88.950 262.050 91.050 ;
        RECT 263.250 89.850 264.750 90.750 ;
        RECT 265.950 88.950 268.050 91.050 ;
        RECT 260.400 88.050 261.450 88.950 ;
        RECT 259.950 85.950 262.050 88.050 ;
        RECT 250.950 79.950 253.050 82.050 ;
        RECT 256.950 79.950 259.050 82.050 ;
        RECT 235.950 73.950 238.050 76.050 ;
        RECT 226.950 64.950 229.050 67.050 ;
        RECT 227.400 55.050 228.450 64.950 ;
        RECT 232.950 58.950 235.050 61.050 ;
        RECT 220.950 52.950 223.050 55.050 ;
        RECT 226.950 52.950 229.050 55.050 ;
        RECT 230.250 53.250 232.050 54.150 ;
        RECT 217.950 49.950 220.050 52.050 ;
        RECT 220.950 50.850 223.050 51.750 ;
        RECT 223.950 50.250 226.050 51.150 ;
        RECT 226.950 50.850 228.750 51.750 ;
        RECT 229.950 51.450 232.050 52.050 ;
        RECT 233.400 51.450 234.450 58.950 ;
        RECT 229.950 50.400 234.450 51.450 ;
        RECT 229.950 49.950 232.050 50.400 ;
        RECT 218.400 49.050 219.450 49.950 ;
        RECT 196.950 46.950 199.050 49.050 ;
        RECT 214.950 46.950 217.050 49.050 ;
        RECT 217.950 46.950 220.050 49.050 ;
        RECT 223.950 46.950 226.050 49.050 ;
        RECT 208.950 31.950 211.050 34.050 ;
        RECT 193.950 28.950 196.050 31.050 ;
        RECT 196.950 28.950 199.050 31.050 ;
        RECT 199.950 28.950 202.050 31.050 ;
        RECT 202.950 28.950 205.050 31.050 ;
        RECT 172.950 25.950 175.050 28.050 ;
        RECT 184.950 25.950 187.050 28.050 ;
        RECT 172.950 23.850 175.050 24.750 ;
        RECT 175.950 23.250 178.050 24.150 ;
        RECT 136.950 20.850 138.750 21.750 ;
        RECT 139.950 19.950 142.050 22.050 ;
        RECT 143.250 20.850 144.750 21.750 ;
        RECT 145.950 21.450 148.050 22.050 ;
        RECT 145.950 20.400 150.450 21.450 ;
        RECT 145.950 19.950 148.050 20.400 ;
        RECT 145.950 17.850 148.050 18.750 ;
        RECT 149.400 16.050 150.450 20.400 ;
        RECT 160.950 19.950 163.050 22.050 ;
        RECT 166.950 19.950 169.050 22.050 ;
        RECT 175.950 19.950 178.050 22.050 ;
        RECT 184.950 20.250 187.050 21.150 ;
        RECT 184.950 16.950 187.050 19.050 ;
        RECT 190.950 17.850 193.050 18.750 ;
        RECT 148.950 13.950 151.050 16.050 ;
        RECT 109.950 10.950 112.050 13.050 ;
        RECT 130.950 10.950 133.050 13.050 ;
        RECT 185.400 10.050 186.450 16.950 ;
        RECT 197.550 10.050 198.750 28.950 ;
        RECT 200.550 16.350 201.750 28.950 ;
        RECT 199.950 14.250 202.050 16.350 ;
        RECT 200.550 10.050 201.750 14.250 ;
        RECT 203.550 10.050 204.750 28.950 ;
        RECT 209.400 28.050 210.450 31.950 ;
        RECT 211.950 29.400 214.050 31.500 ;
        RECT 216.150 29.400 218.250 31.500 ;
        RECT 220.950 29.400 223.050 31.500 ;
        RECT 223.950 29.400 226.050 31.500 ;
        RECT 226.950 29.400 229.050 31.500 ;
        RECT 208.950 25.950 211.050 28.050 ;
        RECT 208.950 23.850 211.050 24.750 ;
        RECT 212.250 20.850 213.450 29.400 ;
        RECT 216.450 23.550 217.650 29.400 ;
        RECT 216.150 21.450 218.250 23.550 ;
        RECT 211.950 18.750 214.050 20.850 ;
        RECT 212.250 12.600 213.450 18.750 ;
        RECT 216.450 12.600 217.650 21.450 ;
        RECT 221.400 15.750 222.600 29.400 ;
        RECT 220.950 13.650 223.050 15.750 ;
        RECT 211.950 10.500 214.050 12.600 ;
        RECT 216.000 10.500 218.100 12.600 ;
        RECT 224.550 12.150 225.750 29.400 ;
        RECT 227.250 15.750 228.450 29.400 ;
        RECT 236.400 22.050 237.450 73.950 ;
        RECT 241.950 59.250 244.050 60.150 ;
        RECT 238.950 56.250 240.750 57.150 ;
        RECT 241.950 55.950 244.050 58.050 ;
        RECT 245.250 56.250 246.750 57.150 ;
        RECT 247.950 55.950 250.050 58.050 ;
        RECT 242.400 55.050 243.450 55.950 ;
        RECT 238.950 52.950 241.050 55.050 ;
        RECT 241.950 52.950 244.050 55.050 ;
        RECT 244.950 52.950 247.050 55.050 ;
        RECT 248.250 53.850 250.050 54.750 ;
        RECT 239.400 49.050 240.450 52.950 ;
        RECT 245.400 52.050 246.450 52.950 ;
        RECT 244.950 49.950 247.050 52.050 ;
        RECT 247.950 49.950 250.050 52.050 ;
        RECT 238.950 46.950 241.050 49.050 ;
        RECT 248.400 31.050 249.450 49.950 ;
        RECT 251.400 46.050 252.450 79.950 ;
        RECT 266.400 67.050 267.450 88.950 ;
        RECT 269.400 85.050 270.450 128.400 ;
        RECT 271.950 127.950 274.050 128.400 ;
        RECT 275.250 128.250 276.750 129.150 ;
        RECT 277.950 127.950 280.050 130.050 ;
        RECT 283.950 129.450 286.050 130.050 ;
        RECT 281.400 128.400 286.050 129.450 ;
        RECT 271.950 125.850 273.750 126.750 ;
        RECT 274.950 124.950 277.050 127.050 ;
        RECT 278.250 125.850 280.050 126.750 ;
        RECT 271.950 109.950 274.050 112.050 ;
        RECT 272.400 94.050 273.450 109.950 ;
        RECT 281.400 106.050 282.450 128.400 ;
        RECT 283.950 127.950 286.050 128.400 ;
        RECT 287.250 128.250 288.750 129.150 ;
        RECT 289.950 127.950 292.050 130.050 ;
        RECT 283.950 125.850 285.750 126.750 ;
        RECT 286.950 124.950 289.050 127.050 ;
        RECT 290.250 125.850 292.050 126.750 ;
        RECT 287.400 124.050 288.450 124.950 ;
        RECT 286.950 121.950 289.050 124.050 ;
        RECT 286.950 115.950 289.050 118.050 ;
        RECT 280.950 103.950 283.050 106.050 ;
        RECT 274.950 100.950 277.050 103.050 ;
        RECT 271.950 91.950 274.050 94.050 ;
        RECT 275.400 91.050 276.450 100.950 ;
        RECT 283.950 97.950 286.050 100.050 ;
        RECT 277.950 91.950 280.050 94.050 ;
        RECT 281.250 92.250 283.050 93.150 ;
        RECT 271.950 89.850 273.750 90.750 ;
        RECT 274.950 88.950 277.050 91.050 ;
        RECT 278.250 89.850 279.750 90.750 ;
        RECT 280.950 88.950 283.050 91.050 ;
        RECT 274.950 86.850 277.050 87.750 ;
        RECT 268.950 82.950 271.050 85.050 ;
        RECT 256.950 64.950 259.050 67.050 ;
        RECT 265.950 64.950 268.050 67.050 ;
        RECT 253.950 61.950 256.050 64.050 ;
        RECT 250.950 43.950 253.050 46.050 ;
        RECT 247.950 28.950 250.050 31.050 ;
        RECT 247.950 23.250 250.050 24.150 ;
        RECT 235.950 19.950 238.050 22.050 ;
        RECT 247.950 21.450 250.050 22.050 ;
        RECT 251.400 21.450 252.450 43.950 ;
        RECT 254.400 22.050 255.450 61.950 ;
        RECT 257.400 49.050 258.450 64.950 ;
        RECT 265.950 58.950 268.050 61.050 ;
        RECT 266.400 58.050 267.450 58.950 ;
        RECT 269.400 58.050 270.450 82.950 ;
        RECT 281.400 73.050 282.450 88.950 ;
        RECT 284.400 88.050 285.450 97.950 ;
        RECT 283.950 85.950 286.050 88.050 ;
        RECT 283.950 76.950 286.050 79.050 ;
        RECT 280.950 70.950 283.050 73.050 ;
        RECT 284.400 58.050 285.450 76.950 ;
        RECT 287.400 61.050 288.450 115.950 ;
        RECT 289.950 112.950 292.050 115.050 ;
        RECT 290.400 97.050 291.450 112.950 ;
        RECT 293.400 100.050 294.450 130.950 ;
        RECT 304.950 127.950 307.050 130.050 ;
        RECT 310.950 127.950 313.050 130.050 ;
        RECT 298.950 125.250 301.050 126.150 ;
        RECT 304.950 125.850 307.050 126.750 ;
        RECT 307.950 125.250 310.050 126.150 ;
        RECT 298.950 121.950 301.050 124.050 ;
        RECT 307.950 121.950 310.050 124.050 ;
        RECT 311.400 120.450 312.450 127.950 ;
        RECT 314.400 124.050 315.450 157.950 ;
        RECT 319.950 154.950 322.050 157.050 ;
        RECT 320.400 127.050 321.450 154.950 ;
        RECT 319.950 124.950 322.050 127.050 ;
        RECT 313.950 121.950 316.050 124.050 ;
        RECT 316.950 122.250 319.050 123.150 ;
        RECT 319.950 122.850 322.050 123.750 ;
        RECT 323.400 121.050 324.450 170.400 ;
        RECT 325.950 169.950 328.050 170.400 ;
        RECT 325.950 167.850 328.050 168.750 ;
        RECT 328.950 167.250 331.050 168.150 ;
        RECT 332.400 166.050 333.450 214.950 ;
        RECT 338.400 213.450 339.450 235.950 ;
        RECT 340.950 234.750 343.050 236.850 ;
        RECT 341.250 228.600 342.450 234.750 ;
        RECT 345.450 228.600 346.650 237.450 ;
        RECT 350.400 231.750 351.600 245.400 ;
        RECT 349.950 229.650 352.050 231.750 ;
        RECT 340.950 226.500 343.050 228.600 ;
        RECT 345.000 226.500 347.100 228.600 ;
        RECT 353.550 228.150 354.750 245.400 ;
        RECT 356.250 231.750 357.450 245.400 ;
        RECT 355.950 229.650 358.050 231.750 ;
        RECT 352.950 226.050 355.050 228.150 ;
        RECT 349.950 223.950 352.050 226.050 ;
        RECT 356.250 225.900 357.450 229.650 ;
        RECT 359.400 228.450 360.450 262.950 ;
        RECT 362.400 231.450 363.450 301.950 ;
        RECT 364.950 298.950 367.050 301.050 ;
        RECT 365.400 277.050 366.450 298.950 ;
        RECT 367.950 289.950 370.050 292.050 ;
        RECT 364.950 274.950 367.050 277.050 ;
        RECT 364.950 271.950 367.050 274.050 ;
        RECT 365.400 265.050 366.450 271.950 ;
        RECT 368.400 271.050 369.450 289.950 ;
        RECT 377.400 274.050 378.450 325.950 ;
        RECT 380.400 321.450 381.450 325.950 ;
        RECT 383.400 325.050 384.450 328.950 ;
        RECT 382.950 322.950 385.050 325.050 ;
        RECT 380.400 320.400 384.450 321.450 ;
        RECT 383.400 310.050 384.450 320.400 ;
        RECT 386.400 316.050 387.450 355.950 ;
        RECT 388.950 341.250 391.050 342.150 ;
        RECT 388.950 337.950 391.050 340.050 ;
        RECT 389.400 325.050 390.450 337.950 ;
        RECT 388.950 322.950 391.050 325.050 ;
        RECT 385.950 313.950 388.050 316.050 ;
        RECT 392.400 313.050 393.450 370.950 ;
        RECT 395.400 322.050 396.450 376.950 ;
        RECT 398.400 349.050 399.450 385.950 ;
        RECT 403.950 383.250 406.050 384.150 ;
        RECT 403.950 379.950 406.050 382.050 ;
        RECT 404.400 373.050 405.450 379.950 ;
        RECT 403.950 370.950 406.050 373.050 ;
        RECT 397.950 346.950 400.050 349.050 ;
        RECT 404.400 346.050 405.450 370.950 ;
        RECT 406.950 364.950 409.050 367.050 ;
        RECT 403.950 343.950 406.050 346.050 ;
        RECT 397.950 341.250 400.050 342.150 ;
        RECT 403.950 341.250 406.050 342.150 ;
        RECT 397.950 337.950 400.050 340.050 ;
        RECT 401.250 338.250 402.750 339.150 ;
        RECT 403.950 337.950 406.050 340.050 ;
        RECT 407.400 339.450 408.450 364.950 ;
        RECT 410.400 346.050 411.450 391.950 ;
        RECT 413.400 373.050 414.450 401.400 ;
        RECT 415.950 391.950 418.050 394.050 ;
        RECT 416.400 382.050 417.450 391.950 ;
        RECT 419.400 385.050 420.450 478.950 ;
        RECT 428.400 475.050 429.450 481.950 ;
        RECT 431.400 481.050 432.450 499.950 ;
        RECT 439.950 493.950 442.050 496.050 ;
        RECT 433.950 490.950 436.050 493.050 ;
        RECT 434.400 490.050 435.450 490.950 ;
        RECT 440.400 490.050 441.450 493.950 ;
        RECT 448.950 490.950 451.050 493.050 ;
        RECT 460.950 490.950 463.050 493.050 ;
        RECT 433.950 487.950 436.050 490.050 ;
        RECT 437.250 488.250 438.750 489.150 ;
        RECT 439.950 487.950 442.050 490.050 ;
        RECT 449.400 487.050 450.450 490.950 ;
        RECT 454.950 488.250 457.050 489.150 ;
        RECT 457.950 487.950 460.050 490.050 ;
        RECT 433.950 485.850 435.750 486.750 ;
        RECT 436.950 484.950 439.050 487.050 ;
        RECT 440.250 485.850 442.050 486.750 ;
        RECT 445.950 485.250 447.750 486.150 ;
        RECT 448.950 484.950 451.050 487.050 ;
        RECT 454.950 486.450 457.050 487.050 ;
        RECT 458.400 486.450 459.450 487.950 ;
        RECT 452.250 485.250 453.750 486.150 ;
        RECT 454.950 485.400 459.450 486.450 ;
        RECT 454.950 484.950 457.050 485.400 ;
        RECT 430.950 478.950 433.050 481.050 ;
        RECT 433.950 478.950 436.050 481.050 ;
        RECT 427.950 472.950 430.050 475.050 ;
        RECT 427.950 469.950 430.050 472.050 ;
        RECT 434.400 471.450 435.450 478.950 ;
        RECT 437.400 475.050 438.450 484.950 ;
        RECT 445.950 481.950 448.050 484.050 ;
        RECT 449.250 482.850 450.750 483.750 ;
        RECT 451.950 481.950 454.050 484.050 ;
        RECT 446.400 475.050 447.450 481.950 ;
        RECT 436.950 472.950 439.050 475.050 ;
        RECT 445.950 472.950 448.050 475.050 ;
        RECT 434.400 470.400 438.450 471.450 ;
        RECT 424.950 457.950 427.050 460.050 ;
        RECT 421.950 455.250 424.050 456.150 ;
        RECT 421.950 451.950 424.050 454.050 ;
        RECT 422.400 415.050 423.450 451.950 ;
        RECT 425.400 442.050 426.450 457.950 ;
        RECT 428.400 451.050 429.450 469.950 ;
        RECT 430.950 457.950 433.050 460.050 ;
        RECT 430.950 455.850 433.050 456.750 ;
        RECT 433.950 455.250 436.050 456.150 ;
        RECT 433.950 451.950 436.050 454.050 ;
        RECT 427.950 448.950 430.050 451.050 ;
        RECT 437.400 448.050 438.450 470.400 ;
        RECT 451.950 463.950 454.050 466.050 ;
        RECT 442.950 460.950 445.050 463.050 ;
        RECT 439.950 454.950 442.050 457.050 ;
        RECT 436.950 445.950 439.050 448.050 ;
        RECT 424.950 439.950 427.050 442.050 ;
        RECT 425.400 427.050 426.450 439.950 ;
        RECT 424.950 424.950 427.050 427.050 ;
        RECT 427.950 419.250 430.050 420.150 ;
        RECT 440.400 418.050 441.450 454.950 ;
        RECT 443.400 454.050 444.450 460.950 ;
        RECT 452.400 457.050 453.450 463.950 ;
        RECT 455.400 460.050 456.450 484.950 ;
        RECT 461.400 463.050 462.450 490.950 ;
        RECT 463.950 488.250 466.050 489.150 ;
        RECT 470.400 487.050 471.450 508.950 ;
        RECT 476.400 493.050 477.450 538.950 ;
        RECT 479.400 538.050 480.450 556.950 ;
        RECT 485.400 556.050 486.450 589.950 ;
        RECT 490.950 571.950 493.050 574.050 ;
        RECT 491.400 571.050 492.450 571.950 ;
        RECT 497.400 571.050 498.450 592.950 ;
        RECT 500.400 574.050 501.450 596.400 ;
        RECT 502.950 595.950 505.050 596.400 ;
        RECT 505.950 595.950 508.050 598.050 ;
        RECT 508.950 595.950 511.050 598.050 ;
        RECT 512.250 596.250 514.050 597.150 ;
        RECT 502.950 593.850 504.750 594.750 ;
        RECT 505.950 592.950 508.050 595.050 ;
        RECT 509.250 593.850 510.750 594.750 ;
        RECT 511.950 592.950 514.050 595.050 ;
        RECT 505.950 590.850 508.050 591.750 ;
        RECT 499.950 571.950 502.050 574.050 ;
        RECT 490.950 568.950 493.050 571.050 ;
        RECT 496.950 568.950 499.050 571.050 ;
        RECT 487.950 562.950 490.050 565.050 ;
        RECT 484.950 553.950 487.050 556.050 ;
        RECT 488.400 541.050 489.450 562.950 ;
        RECT 491.400 555.450 492.450 568.950 ;
        RECT 496.950 562.950 499.050 565.050 ;
        RECT 497.400 559.050 498.450 562.950 ;
        RECT 502.950 559.950 505.050 562.050 ;
        RECT 508.950 559.950 511.050 562.050 ;
        RECT 503.400 559.050 504.450 559.950 ;
        RECT 493.950 557.250 495.750 558.150 ;
        RECT 496.950 556.950 499.050 559.050 ;
        RECT 500.250 557.250 501.750 558.150 ;
        RECT 502.950 556.950 505.050 559.050 ;
        RECT 506.250 557.250 508.050 558.150 ;
        RECT 493.950 555.450 496.050 556.050 ;
        RECT 491.400 554.400 496.050 555.450 ;
        RECT 497.250 554.850 498.750 555.750 ;
        RECT 493.950 553.950 496.050 554.400 ;
        RECT 499.950 553.950 502.050 556.050 ;
        RECT 503.250 554.850 504.750 555.750 ;
        RECT 505.950 555.450 508.050 556.050 ;
        RECT 509.400 555.450 510.450 559.950 ;
        RECT 505.950 554.400 510.450 555.450 ;
        RECT 505.950 553.950 508.050 554.400 ;
        RECT 500.400 544.050 501.450 553.950 ;
        RECT 493.950 541.950 496.050 544.050 ;
        RECT 499.950 541.950 502.050 544.050 ;
        RECT 487.950 538.950 490.050 541.050 ;
        RECT 478.950 535.950 481.050 538.050 ;
        RECT 478.950 532.950 481.050 535.050 ;
        RECT 481.950 532.950 484.050 535.050 ;
        RECT 484.950 532.950 487.050 535.050 ;
        RECT 479.250 514.050 480.450 532.950 ;
        RECT 482.250 520.350 483.450 532.950 ;
        RECT 481.950 518.250 484.050 520.350 ;
        RECT 482.250 514.050 483.450 518.250 ;
        RECT 485.250 514.050 486.450 532.950 ;
        RECT 487.950 529.950 490.050 532.050 ;
        RECT 478.950 511.950 481.050 514.050 ;
        RECT 481.950 511.950 484.050 514.050 ;
        RECT 484.950 511.950 487.050 514.050 ;
        RECT 478.950 499.950 481.050 502.050 ;
        RECT 475.950 490.950 478.050 493.050 ;
        RECT 479.400 490.050 480.450 499.950 ;
        RECT 478.950 487.950 481.050 490.050 ;
        RECT 484.950 488.250 487.050 489.150 ;
        RECT 463.950 484.950 466.050 487.050 ;
        RECT 467.250 485.250 468.750 486.150 ;
        RECT 469.950 484.950 472.050 487.050 ;
        RECT 473.250 485.250 475.050 486.150 ;
        RECT 475.950 484.950 478.050 487.050 ;
        RECT 478.950 485.850 481.050 486.750 ;
        RECT 464.400 484.050 465.450 484.950 ;
        RECT 463.950 481.950 466.050 484.050 ;
        RECT 466.950 481.950 469.050 484.050 ;
        RECT 470.250 482.850 471.750 483.750 ;
        RECT 472.950 481.950 475.050 484.050 ;
        RECT 467.400 475.050 468.450 481.950 ;
        RECT 473.400 481.050 474.450 481.950 ;
        RECT 472.950 478.950 475.050 481.050 ;
        RECT 472.950 475.950 475.050 478.050 ;
        RECT 466.950 472.950 469.050 475.050 ;
        RECT 463.950 463.950 466.050 466.050 ;
        RECT 460.950 460.950 463.050 463.050 ;
        RECT 454.950 457.950 457.050 460.050 ;
        RECT 445.950 454.950 448.050 457.050 ;
        RECT 449.250 455.250 450.750 456.150 ;
        RECT 451.950 454.950 454.050 457.050 ;
        RECT 454.950 454.950 457.050 457.050 ;
        RECT 458.250 455.250 459.750 456.150 ;
        RECT 460.950 454.950 463.050 457.050 ;
        RECT 464.400 454.050 465.450 463.950 ;
        RECT 466.950 460.950 469.050 463.050 ;
        RECT 442.950 451.950 445.050 454.050 ;
        RECT 446.250 452.850 447.750 453.750 ;
        RECT 448.950 451.950 451.050 454.050 ;
        RECT 452.250 452.850 454.050 453.750 ;
        RECT 454.950 452.850 456.750 453.750 ;
        RECT 457.950 451.950 460.050 454.050 ;
        RECT 461.250 452.850 462.750 453.750 ;
        RECT 463.950 451.950 466.050 454.050 ;
        RECT 442.950 449.850 445.050 450.750 ;
        RECT 449.400 433.050 450.450 451.950 ;
        RECT 458.400 448.050 459.450 451.950 ;
        RECT 463.950 449.850 466.050 450.750 ;
        RECT 457.950 445.950 460.050 448.050 ;
        RECT 448.950 430.950 451.050 433.050 ;
        RECT 467.400 421.050 468.450 460.950 ;
        RECT 473.400 448.050 474.450 475.950 ;
        RECT 476.400 463.050 477.450 484.950 ;
        RECT 484.950 481.950 487.050 484.050 ;
        RECT 478.950 478.950 481.050 481.050 ;
        RECT 479.400 469.050 480.450 478.950 ;
        RECT 481.950 469.950 484.050 472.050 ;
        RECT 478.950 466.950 481.050 469.050 ;
        RECT 475.950 460.950 478.050 463.050 ;
        RECT 475.950 457.950 478.050 460.050 ;
        RECT 475.950 455.850 478.050 456.750 ;
        RECT 478.950 455.250 481.050 456.150 ;
        RECT 478.950 451.950 481.050 454.050 ;
        RECT 475.950 448.950 478.050 451.050 ;
        RECT 472.950 445.950 475.050 448.050 ;
        RECT 448.950 419.250 451.050 420.150 ;
        RECT 460.950 418.950 463.050 421.050 ;
        RECT 466.950 418.950 469.050 421.050 ;
        RECT 424.950 416.250 426.750 417.150 ;
        RECT 427.950 415.950 430.050 418.050 ;
        RECT 433.950 417.450 436.050 418.050 ;
        RECT 431.250 416.250 432.750 417.150 ;
        RECT 433.950 416.400 438.450 417.450 ;
        RECT 433.950 415.950 436.050 416.400 ;
        RECT 421.950 412.950 424.050 415.050 ;
        RECT 424.950 412.950 427.050 415.050 ;
        RECT 430.950 412.950 433.050 415.050 ;
        RECT 434.250 413.850 436.050 414.750 ;
        RECT 425.400 409.050 426.450 412.950 ;
        RECT 437.400 412.050 438.450 416.400 ;
        RECT 439.950 415.950 442.050 418.050 ;
        RECT 445.950 416.250 447.750 417.150 ;
        RECT 448.950 415.950 451.050 418.050 ;
        RECT 452.250 416.250 453.750 417.150 ;
        RECT 454.950 415.950 457.050 418.050 ;
        RECT 445.950 412.950 448.050 415.050 ;
        RECT 451.950 412.950 454.050 415.050 ;
        RECT 455.250 413.850 457.050 414.750 ;
        RECT 436.950 409.950 439.050 412.050 ;
        RECT 424.950 406.950 427.050 409.050 ;
        RECT 446.400 397.050 447.450 412.950 ;
        RECT 452.400 412.050 453.450 412.950 ;
        RECT 451.950 409.950 454.050 412.050 ;
        RECT 445.950 394.950 448.050 397.050 ;
        RECT 424.950 389.400 427.050 391.500 ;
        RECT 427.950 389.400 430.050 391.500 ;
        RECT 430.950 389.400 433.050 391.500 ;
        RECT 435.750 389.400 437.850 391.500 ;
        RECT 439.950 389.400 442.050 391.500 ;
        RECT 418.950 382.950 421.050 385.050 ;
        RECT 415.950 379.950 418.050 382.050 ;
        RECT 415.950 377.850 418.050 378.750 ;
        RECT 425.550 375.750 426.750 389.400 ;
        RECT 424.950 373.650 427.050 375.750 ;
        RECT 412.950 370.950 415.050 373.050 ;
        RECT 425.550 369.900 426.750 373.650 ;
        RECT 428.250 372.150 429.450 389.400 ;
        RECT 431.400 375.750 432.600 389.400 ;
        RECT 436.350 383.550 437.550 389.400 ;
        RECT 435.750 381.450 437.850 383.550 ;
        RECT 430.950 373.650 433.050 375.750 ;
        RECT 436.350 372.600 437.550 381.450 ;
        RECT 440.550 380.850 441.750 389.400 ;
        RECT 442.950 388.950 445.050 391.050 ;
        RECT 448.950 388.950 451.050 391.050 ;
        RECT 451.950 388.950 454.050 391.050 ;
        RECT 454.950 388.950 457.050 391.050 ;
        RECT 443.400 388.050 444.450 388.950 ;
        RECT 442.950 385.950 445.050 388.050 ;
        RECT 442.950 383.850 445.050 384.750 ;
        RECT 439.950 378.750 442.050 380.850 ;
        RECT 440.550 372.600 441.750 378.750 ;
        RECT 427.950 370.050 430.050 372.150 ;
        RECT 435.900 370.500 438.000 372.600 ;
        RECT 439.950 370.500 442.050 372.600 ;
        RECT 449.250 370.050 450.450 388.950 ;
        RECT 452.250 376.350 453.450 388.950 ;
        RECT 451.950 374.250 454.050 376.350 ;
        RECT 452.250 370.050 453.450 374.250 ;
        RECT 455.250 370.050 456.450 388.950 ;
        RECT 461.400 385.050 462.450 418.950 ;
        RECT 466.950 415.950 469.050 418.050 ;
        RECT 472.950 416.250 475.050 417.150 ;
        RECT 467.400 415.050 468.450 415.950 ;
        RECT 463.950 413.250 465.750 414.150 ;
        RECT 466.950 412.950 469.050 415.050 ;
        RECT 470.250 413.250 471.750 414.150 ;
        RECT 472.950 412.950 475.050 415.050 ;
        RECT 463.950 409.950 466.050 412.050 ;
        RECT 467.250 410.850 468.750 411.750 ;
        RECT 469.950 409.950 472.050 412.050 ;
        RECT 470.400 391.050 471.450 409.950 ;
        RECT 473.400 409.050 474.450 412.950 ;
        RECT 476.400 412.050 477.450 448.950 ;
        RECT 482.400 424.050 483.450 469.950 ;
        RECT 485.400 463.050 486.450 481.950 ;
        RECT 488.400 472.050 489.450 529.950 ;
        RECT 494.400 526.050 495.450 541.950 ;
        RECT 499.950 535.950 502.050 538.050 ;
        RECT 493.950 523.950 496.050 526.050 ;
        RECT 496.950 524.250 499.050 525.150 ;
        RECT 490.950 521.850 493.050 522.750 ;
        RECT 496.950 520.950 499.050 523.050 ;
        RECT 497.400 520.050 498.450 520.950 ;
        RECT 496.950 517.950 499.050 520.050 ;
        RECT 497.400 502.050 498.450 517.950 ;
        RECT 496.950 499.950 499.050 502.050 ;
        RECT 490.950 496.950 493.050 499.050 ;
        RECT 493.950 496.950 496.050 499.050 ;
        RECT 496.950 496.950 499.050 499.050 ;
        RECT 491.550 478.050 492.750 496.950 ;
        RECT 494.550 492.750 495.750 496.950 ;
        RECT 493.950 490.650 496.050 492.750 ;
        RECT 494.550 478.050 495.750 490.650 ;
        RECT 497.550 478.050 498.750 496.950 ;
        RECT 490.950 475.950 493.050 478.050 ;
        RECT 493.950 475.950 496.050 478.050 ;
        RECT 496.950 475.950 499.050 478.050 ;
        RECT 487.950 469.950 490.050 472.050 ;
        RECT 490.950 463.950 493.050 466.050 ;
        RECT 484.950 460.950 487.050 463.050 ;
        RECT 484.950 457.950 487.050 460.050 ;
        RECT 485.400 454.050 486.450 457.950 ;
        RECT 487.950 454.950 490.050 457.050 ;
        RECT 484.950 451.950 487.050 454.050 ;
        RECT 488.400 451.050 489.450 454.950 ;
        RECT 491.400 454.050 492.450 463.950 ;
        RECT 496.950 460.950 499.050 463.050 ;
        RECT 497.400 460.050 498.450 460.950 ;
        RECT 496.950 457.950 499.050 460.050 ;
        RECT 500.400 457.050 501.450 535.950 ;
        RECT 508.950 532.950 511.050 535.050 ;
        RECT 502.950 529.950 505.050 532.050 ;
        RECT 503.400 529.050 504.450 529.950 ;
        RECT 509.400 529.050 510.450 532.950 ;
        RECT 512.400 532.050 513.450 592.950 ;
        RECT 515.400 562.050 516.450 631.950 ;
        RECT 520.950 629.250 523.050 630.150 ;
        RECT 526.950 629.250 529.050 630.150 ;
        RECT 520.950 625.950 523.050 628.050 ;
        RECT 524.250 626.250 525.750 627.150 ;
        RECT 526.950 625.950 529.050 628.050 ;
        RECT 521.400 616.050 522.450 625.950 ;
        RECT 523.950 622.950 526.050 625.050 ;
        RECT 520.950 613.950 523.050 616.050 ;
        RECT 521.400 613.050 522.450 613.950 ;
        RECT 520.950 610.950 523.050 613.050 ;
        RECT 520.950 604.950 523.050 607.050 ;
        RECT 521.400 598.050 522.450 604.950 ;
        RECT 517.950 596.250 519.750 597.150 ;
        RECT 520.950 595.950 523.050 598.050 ;
        RECT 524.250 596.250 526.050 597.150 ;
        RECT 517.950 592.950 520.050 595.050 ;
        RECT 521.250 593.850 522.750 594.750 ;
        RECT 523.950 592.950 526.050 595.050 ;
        RECT 518.400 565.050 519.450 592.950 ;
        RECT 527.400 574.050 528.450 625.950 ;
        RECT 530.400 595.050 531.450 664.950 ;
        RECT 532.950 661.950 535.050 664.050 ;
        RECT 533.400 661.050 534.450 661.950 ;
        RECT 532.950 658.950 535.050 661.050 ;
        RECT 548.400 637.050 549.450 673.950 ;
        RECT 554.400 673.050 555.450 673.950 ;
        RECT 560.400 673.050 561.450 709.950 ;
        RECT 562.950 703.950 565.050 706.050 ;
        RECT 568.950 705.450 571.050 706.050 ;
        RECT 572.400 705.450 573.450 743.400 ;
        RECT 574.950 740.250 576.750 741.150 ;
        RECT 577.950 739.950 580.050 742.050 ;
        RECT 581.250 740.250 583.050 741.150 ;
        RECT 574.950 736.950 577.050 739.050 ;
        RECT 578.250 737.850 579.750 738.750 ;
        RECT 580.950 736.950 583.050 739.050 ;
        RECT 575.400 709.050 576.450 736.950 ;
        RECT 581.400 727.050 582.450 736.950 ;
        RECT 584.400 733.050 585.450 752.400 ;
        RECT 586.950 748.950 589.050 751.050 ;
        RECT 587.400 748.050 588.450 748.950 ;
        RECT 602.400 748.050 603.450 766.950 ;
        RECT 605.400 748.050 606.450 772.950 ;
        RECT 608.400 772.050 609.450 775.950 ;
        RECT 607.950 769.950 610.050 772.050 ;
        RECT 617.400 769.050 618.450 776.400 ;
        RECT 619.950 775.950 622.050 776.400 ;
        RECT 623.250 776.250 624.750 777.150 ;
        RECT 625.950 775.950 628.050 778.050 ;
        RECT 619.950 773.850 621.750 774.750 ;
        RECT 622.950 772.950 625.050 775.050 ;
        RECT 626.250 773.850 628.050 774.750 ;
        RECT 623.400 769.050 624.450 772.950 ;
        RECT 616.950 766.950 619.050 769.050 ;
        RECT 622.950 766.950 625.050 769.050 ;
        RECT 625.950 766.950 628.050 769.050 ;
        RECT 586.950 745.950 589.050 748.050 ;
        RECT 592.950 747.450 595.050 748.050 ;
        RECT 592.950 746.400 597.450 747.450 ;
        RECT 592.950 745.950 595.050 746.400 ;
        RECT 587.400 741.450 588.450 745.950 ;
        RECT 596.400 745.050 597.450 746.400 ;
        RECT 601.950 745.950 604.050 748.050 ;
        RECT 604.950 745.950 607.050 748.050 ;
        RECT 607.950 745.950 610.050 748.050 ;
        RECT 619.950 745.950 622.050 748.050 ;
        RECT 608.400 745.050 609.450 745.950 ;
        RECT 589.950 743.250 592.050 744.150 ;
        RECT 592.950 743.850 595.050 744.750 ;
        RECT 595.950 744.450 598.050 745.050 ;
        RECT 598.950 744.450 601.050 745.050 ;
        RECT 595.950 743.400 601.050 744.450 ;
        RECT 602.250 743.850 603.750 744.750 ;
        RECT 595.950 742.950 598.050 743.400 ;
        RECT 598.950 742.950 601.050 743.400 ;
        RECT 604.950 742.950 607.050 745.050 ;
        RECT 607.950 742.950 610.050 745.050 ;
        RECT 611.250 743.250 612.750 744.150 ;
        RECT 613.950 742.950 616.050 745.050 ;
        RECT 616.950 742.950 619.050 745.050 ;
        RECT 589.950 741.450 592.050 742.050 ;
        RECT 596.400 741.450 597.450 742.950 ;
        RECT 617.400 742.050 618.450 742.950 ;
        RECT 587.400 740.400 592.050 741.450 ;
        RECT 589.950 739.950 592.050 740.400 ;
        RECT 593.400 740.400 597.450 741.450 ;
        RECT 598.950 740.850 601.050 741.750 ;
        RECT 604.950 740.850 607.050 741.750 ;
        RECT 607.950 740.850 609.750 741.750 ;
        RECT 583.950 730.950 586.050 733.050 ;
        RECT 580.950 724.950 583.050 727.050 ;
        RECT 574.950 706.950 577.050 709.050 ;
        RECT 583.950 706.950 586.050 709.050 ;
        RECT 589.950 706.950 592.050 709.050 ;
        RECT 566.250 704.250 567.750 705.150 ;
        RECT 568.950 704.400 576.450 705.450 ;
        RECT 568.950 703.950 571.050 704.400 ;
        RECT 562.950 701.850 564.750 702.750 ;
        RECT 565.950 700.950 568.050 703.050 ;
        RECT 569.250 701.850 571.050 702.750 ;
        RECT 571.950 700.950 574.050 703.050 ;
        RECT 566.400 694.050 567.450 700.950 ;
        RECT 572.400 697.050 573.450 700.950 ;
        RECT 571.950 694.950 574.050 697.050 ;
        RECT 575.400 696.450 576.450 704.400 ;
        RECT 580.950 701.250 583.050 702.150 ;
        RECT 577.950 698.250 579.750 699.150 ;
        RECT 580.950 697.950 583.050 700.050 ;
        RECT 581.400 697.050 582.450 697.950 ;
        RECT 577.950 696.450 580.050 697.050 ;
        RECT 575.400 695.400 580.050 696.450 ;
        RECT 577.950 694.950 580.050 695.400 ;
        RECT 580.950 694.950 583.050 697.050 ;
        RECT 565.950 691.950 568.050 694.050 ;
        RECT 580.950 682.950 583.050 685.050 ;
        RECT 562.950 676.950 565.050 679.050 ;
        RECT 574.950 676.950 577.050 679.050 ;
        RECT 553.950 670.950 556.050 673.050 ;
        RECT 557.250 671.850 558.750 672.750 ;
        RECT 559.950 670.950 562.050 673.050 ;
        RECT 553.950 668.850 556.050 669.750 ;
        RECT 556.950 667.950 559.050 670.050 ;
        RECT 559.950 668.850 562.050 669.750 ;
        RECT 541.950 634.950 544.050 637.050 ;
        RECT 547.950 634.950 550.050 637.050 ;
        RECT 532.950 631.950 535.050 634.050 ;
        RECT 533.400 628.050 534.450 631.950 ;
        RECT 535.950 628.950 538.050 631.050 ;
        RECT 532.950 625.950 535.050 628.050 ;
        RECT 535.950 626.850 538.050 627.750 ;
        RECT 538.950 626.250 541.050 627.150 ;
        RECT 538.950 622.950 541.050 625.050 ;
        RECT 539.400 613.050 540.450 622.950 ;
        RECT 532.950 610.950 535.050 613.050 ;
        RECT 538.950 610.950 541.050 613.050 ;
        RECT 533.400 601.050 534.450 610.950 ;
        RECT 535.950 604.950 538.050 607.050 ;
        RECT 536.400 604.050 537.450 604.950 ;
        RECT 535.950 601.950 538.050 604.050 ;
        RECT 532.950 598.950 535.050 601.050 ;
        RECT 536.250 599.850 537.750 600.750 ;
        RECT 538.950 600.450 541.050 601.050 ;
        RECT 542.400 600.450 543.450 634.950 ;
        RECT 544.950 632.250 547.050 633.150 ;
        RECT 544.950 628.950 547.050 631.050 ;
        RECT 548.250 629.250 549.750 630.150 ;
        RECT 550.950 628.950 553.050 631.050 ;
        RECT 554.250 629.250 556.050 630.150 ;
        RECT 547.950 625.950 550.050 628.050 ;
        RECT 551.250 626.850 552.750 627.750 ;
        RECT 553.950 625.950 556.050 628.050 ;
        RECT 557.400 627.450 558.450 667.950 ;
        RECT 563.400 634.050 564.450 676.950 ;
        RECT 568.950 673.950 571.050 676.050 ;
        RECT 571.950 673.950 574.050 676.050 ;
        RECT 569.400 673.050 570.450 673.950 ;
        RECT 575.400 673.050 576.450 676.950 ;
        RECT 568.950 670.950 571.050 673.050 ;
        RECT 572.250 671.850 573.750 672.750 ;
        RECT 574.950 670.950 577.050 673.050 ;
        RECT 568.950 668.850 571.050 669.750 ;
        RECT 574.950 668.850 577.050 669.750 ;
        RECT 568.950 664.950 571.050 667.050 ;
        RECT 562.950 631.950 565.050 634.050 ;
        RECT 559.950 629.250 562.050 630.150 ;
        RECT 565.950 629.250 568.050 630.150 ;
        RECT 559.950 627.450 562.050 628.050 ;
        RECT 557.400 626.400 562.050 627.450 ;
        RECT 548.400 622.050 549.450 625.950 ;
        RECT 554.400 625.050 555.450 625.950 ;
        RECT 553.950 622.950 556.050 625.050 ;
        RECT 547.950 619.950 550.050 622.050 ;
        RECT 547.950 604.950 550.050 607.050 ;
        RECT 553.950 604.950 556.050 607.050 ;
        RECT 548.400 604.050 549.450 604.950 ;
        RECT 547.950 601.950 550.050 604.050 ;
        RECT 538.950 599.400 543.450 600.450 ;
        RECT 547.950 599.850 550.050 600.750 ;
        RECT 538.950 598.950 541.050 599.400 ;
        RECT 550.950 599.250 553.050 600.150 ;
        RECT 532.950 596.850 535.050 597.750 ;
        RECT 538.950 596.850 541.050 597.750 ;
        RECT 550.950 595.950 553.050 598.050 ;
        RECT 529.950 592.950 532.050 595.050 ;
        RECT 526.950 571.950 529.050 574.050 ;
        RECT 526.950 568.950 529.050 571.050 ;
        RECT 517.950 562.950 520.050 565.050 ;
        RECT 514.950 559.950 517.050 562.050 ;
        RECT 517.950 559.950 520.050 562.050 ;
        RECT 523.950 560.250 526.050 561.150 ;
        RECT 518.400 559.050 519.450 559.950 ;
        RECT 514.950 557.250 516.750 558.150 ;
        RECT 517.950 556.950 520.050 559.050 ;
        RECT 521.250 557.250 522.750 558.150 ;
        RECT 523.950 556.950 526.050 559.050 ;
        RECT 514.950 553.950 517.050 556.050 ;
        RECT 518.250 554.850 519.750 555.750 ;
        RECT 520.950 553.950 523.050 556.050 ;
        RECT 524.400 553.050 525.450 556.950 ;
        RECT 523.950 550.950 526.050 553.050 ;
        RECT 514.950 538.950 517.050 541.050 ;
        RECT 511.950 529.950 514.050 532.050 ;
        RECT 515.400 529.050 516.450 538.950 ;
        RECT 502.950 526.950 505.050 529.050 ;
        RECT 506.250 527.250 507.750 528.150 ;
        RECT 508.950 526.950 511.050 529.050 ;
        RECT 512.250 527.250 513.750 528.150 ;
        RECT 514.950 526.950 517.050 529.050 ;
        RECT 527.400 528.450 528.450 568.950 ;
        RECT 541.950 565.950 544.050 568.050 ;
        RECT 532.950 557.250 535.050 558.150 ;
        RECT 538.950 557.250 541.050 558.150 ;
        RECT 532.950 553.950 535.050 556.050 ;
        RECT 536.250 554.250 537.750 555.150 ;
        RECT 538.950 553.950 541.050 556.050 ;
        RECT 535.950 550.950 538.050 553.050 ;
        RECT 536.400 544.050 537.450 550.950 ;
        RECT 535.950 541.950 538.050 544.050 ;
        RECT 542.400 541.050 543.450 565.950 ;
        RECT 551.400 562.050 552.450 595.950 ;
        RECT 550.950 559.950 553.050 562.050 ;
        RECT 544.950 556.950 547.050 559.050 ;
        RECT 544.950 554.850 547.050 555.750 ;
        RECT 547.950 554.250 550.050 555.150 ;
        RECT 547.950 550.950 550.050 553.050 ;
        RECT 541.950 538.950 544.050 541.050 ;
        RECT 548.400 538.050 549.450 550.950 ;
        RECT 547.950 535.950 550.050 538.050 ;
        RECT 529.950 532.950 532.050 535.050 ;
        RECT 524.400 527.400 528.450 528.450 ;
        RECT 502.950 524.850 504.750 525.750 ;
        RECT 505.950 523.950 508.050 526.050 ;
        RECT 509.250 524.850 510.750 525.750 ;
        RECT 511.950 523.950 514.050 526.050 ;
        RECT 515.250 524.850 517.050 525.750 ;
        RECT 520.950 523.950 523.050 526.050 ;
        RECT 506.400 522.450 507.450 523.950 ;
        RECT 503.400 521.400 507.450 522.450 ;
        RECT 503.400 487.050 504.450 521.400 ;
        RECT 521.400 508.050 522.450 523.950 ;
        RECT 520.950 505.950 523.050 508.050 ;
        RECT 524.400 501.450 525.450 527.400 ;
        RECT 526.950 523.950 529.050 526.050 ;
        RECT 530.400 523.050 531.450 532.950 ;
        RECT 554.400 532.050 555.450 604.950 ;
        RECT 557.400 604.050 558.450 626.400 ;
        RECT 559.950 625.950 562.050 626.400 ;
        RECT 563.250 626.250 564.750 627.150 ;
        RECT 565.950 625.950 568.050 628.050 ;
        RECT 559.950 622.950 562.050 625.050 ;
        RECT 562.950 622.950 565.050 625.050 ;
        RECT 556.950 601.950 559.050 604.050 ;
        RECT 560.400 601.050 561.450 622.950 ;
        RECT 565.950 613.950 568.050 616.050 ;
        RECT 562.950 610.950 565.050 613.050 ;
        RECT 563.400 604.050 564.450 610.950 ;
        RECT 566.400 604.050 567.450 613.950 ;
        RECT 569.400 607.050 570.450 664.950 ;
        RECT 581.400 637.050 582.450 682.950 ;
        RECT 584.400 682.050 585.450 706.950 ;
        RECT 586.950 703.950 589.050 706.050 ;
        RECT 587.400 703.050 588.450 703.950 ;
        RECT 586.950 700.950 589.050 703.050 ;
        RECT 586.950 698.850 589.050 699.750 ;
        RECT 590.400 694.050 591.450 706.950 ;
        RECT 593.400 700.050 594.450 740.400 ;
        RECT 610.950 739.950 613.050 742.050 ;
        RECT 614.250 740.850 615.750 741.750 ;
        RECT 616.950 739.950 619.050 742.050 ;
        RECT 611.400 739.050 612.450 739.950 ;
        RECT 620.400 739.050 621.450 745.950 ;
        RECT 610.950 736.950 613.050 739.050 ;
        RECT 616.950 737.850 619.050 738.750 ;
        RECT 619.950 736.950 622.050 739.050 ;
        RECT 611.400 736.050 612.450 736.950 ;
        RECT 610.950 733.950 613.050 736.050 ;
        RECT 595.950 706.950 598.050 709.050 ;
        RECT 607.950 706.950 610.050 709.050 ;
        RECT 596.400 706.050 597.450 706.950 ;
        RECT 595.950 703.950 598.050 706.050 ;
        RECT 599.250 704.250 600.750 705.150 ;
        RECT 601.950 703.950 604.050 706.050 ;
        RECT 604.950 703.950 607.050 706.050 ;
        RECT 595.950 701.850 597.750 702.750 ;
        RECT 598.950 700.950 601.050 703.050 ;
        RECT 602.250 701.850 604.050 702.750 ;
        RECT 592.950 697.950 595.050 700.050 ;
        RECT 605.400 697.050 606.450 703.950 ;
        RECT 608.400 703.050 609.450 706.950 ;
        RECT 607.950 700.950 610.050 703.050 ;
        RECT 595.950 694.950 598.050 697.050 ;
        RECT 604.950 694.950 607.050 697.050 ;
        RECT 589.950 691.950 592.050 694.050 ;
        RECT 583.950 679.950 586.050 682.050 ;
        RECT 583.950 673.950 586.050 676.050 ;
        RECT 589.950 673.950 592.050 676.050 ;
        RECT 592.950 673.950 595.050 676.050 ;
        RECT 580.950 634.950 583.050 637.050 ;
        RECT 574.950 633.450 577.050 634.050 ;
        RECT 572.400 632.400 577.050 633.450 ;
        RECT 580.950 633.450 583.050 634.050 ;
        RECT 584.400 633.450 585.450 673.950 ;
        RECT 593.400 673.050 594.450 673.950 ;
        RECT 586.950 670.950 589.050 673.050 ;
        RECT 590.250 671.850 591.750 672.750 ;
        RECT 592.950 670.950 595.050 673.050 ;
        RECT 596.400 670.050 597.450 694.950 ;
        RECT 598.950 685.950 601.050 688.050 ;
        RECT 599.400 673.050 600.450 685.950 ;
        RECT 611.400 679.050 612.450 733.950 ;
        RECT 616.950 703.950 619.050 706.050 ;
        RECT 622.950 704.250 625.050 705.150 ;
        RECT 617.400 703.050 618.450 703.950 ;
        RECT 613.950 701.250 615.750 702.150 ;
        RECT 616.950 700.950 619.050 703.050 ;
        RECT 620.250 701.250 621.750 702.150 ;
        RECT 622.950 700.950 625.050 703.050 ;
        RECT 613.950 697.950 616.050 700.050 ;
        RECT 617.250 698.850 618.750 699.750 ;
        RECT 619.950 697.950 622.050 700.050 ;
        RECT 614.400 688.050 615.450 697.950 ;
        RECT 620.400 697.050 621.450 697.950 ;
        RECT 619.950 694.950 622.050 697.050 ;
        RECT 613.950 685.950 616.050 688.050 ;
        RECT 610.950 676.950 613.050 679.050 ;
        RECT 601.950 673.950 604.050 676.050 ;
        RECT 604.950 673.950 607.050 676.050 ;
        RECT 607.950 673.950 610.050 676.050 ;
        RECT 605.400 673.050 606.450 673.950 ;
        RECT 598.950 670.950 601.050 673.050 ;
        RECT 602.250 671.850 603.750 672.750 ;
        RECT 604.950 670.950 607.050 673.050 ;
        RECT 586.950 668.850 589.050 669.750 ;
        RECT 592.950 668.850 595.050 669.750 ;
        RECT 595.950 667.950 598.050 670.050 ;
        RECT 598.950 668.850 601.050 669.750 ;
        RECT 604.950 668.850 607.050 669.750 ;
        RECT 596.400 649.050 597.450 667.950 ;
        RECT 595.950 646.950 598.050 649.050 ;
        RECT 586.950 634.950 589.050 637.050 ;
        RECT 608.400 636.450 609.450 673.950 ;
        RECT 614.400 637.050 615.450 685.950 ;
        RECT 616.950 679.950 619.050 682.050 ;
        RECT 617.400 670.050 618.450 679.950 ;
        RECT 623.400 676.050 624.450 700.950 ;
        RECT 626.400 685.050 627.450 766.950 ;
        RECT 629.400 703.050 630.450 799.950 ;
        RECT 635.400 775.050 636.450 803.400 ;
        RECT 634.950 772.950 637.050 775.050 ;
        RECT 631.950 770.250 634.050 771.150 ;
        RECT 634.950 770.850 637.050 771.750 ;
        RECT 631.950 766.950 634.050 769.050 ;
        RECT 641.400 757.050 642.450 808.950 ;
        RECT 647.400 808.050 648.450 811.950 ;
        RECT 653.400 810.450 654.450 814.950 ;
        RECT 655.950 812.250 657.750 813.150 ;
        RECT 658.950 811.950 661.050 814.050 ;
        RECT 662.250 812.250 664.050 813.150 ;
        RECT 664.950 811.950 667.050 814.050 ;
        RECT 667.950 811.950 670.050 814.050 ;
        RECT 670.950 812.250 672.750 813.150 ;
        RECT 673.950 811.950 676.050 814.050 ;
        RECT 655.950 810.450 658.050 811.050 ;
        RECT 653.400 809.400 658.050 810.450 ;
        RECT 659.250 809.850 660.750 810.750 ;
        RECT 655.950 808.950 658.050 809.400 ;
        RECT 661.950 808.950 664.050 811.050 ;
        RECT 646.950 805.950 649.050 808.050 ;
        RECT 643.950 781.950 646.050 784.050 ;
        RECT 644.400 766.050 645.450 781.950 ;
        RECT 656.400 778.050 657.450 808.950 ;
        RECT 662.400 805.050 663.450 808.950 ;
        RECT 665.400 805.050 666.450 811.950 ;
        RECT 661.950 802.950 664.050 805.050 ;
        RECT 664.950 802.950 667.050 805.050 ;
        RECT 668.400 802.050 669.450 811.950 ;
        RECT 677.400 811.050 678.450 814.950 ;
        RECT 692.400 814.050 693.450 817.950 ;
        RECT 712.950 814.950 715.050 817.050 ;
        RECT 733.950 814.950 736.050 817.050 ;
        RECT 742.950 814.950 745.050 817.050 ;
        RECT 751.950 815.250 754.050 816.150 ;
        RECT 754.950 815.850 757.050 816.750 ;
        RECT 775.950 814.950 778.050 817.050 ;
        RECT 778.950 814.950 781.050 817.050 ;
        RECT 784.950 816.450 787.050 817.050 ;
        RECT 784.950 815.400 789.450 816.450 ;
        RECT 784.950 814.950 787.050 815.400 ;
        RECT 679.950 813.450 682.050 814.050 ;
        RECT 679.950 812.400 684.450 813.450 ;
        RECT 679.950 811.950 682.050 812.400 ;
        RECT 670.950 808.950 673.050 811.050 ;
        RECT 674.250 809.850 675.750 810.750 ;
        RECT 676.950 808.950 679.050 811.050 ;
        RECT 680.250 809.850 682.050 810.750 ;
        RECT 671.400 808.050 672.450 808.950 ;
        RECT 670.950 805.950 673.050 808.050 ;
        RECT 676.950 806.850 679.050 807.750 ;
        RECT 667.950 799.950 670.050 802.050 ;
        RECT 676.950 778.950 679.050 781.050 ;
        RECT 655.950 775.950 658.050 778.050 ;
        RECT 661.950 775.950 664.050 778.050 ;
        RECT 673.950 776.250 676.050 777.150 ;
        RECT 649.950 773.250 652.050 774.150 ;
        RECT 655.950 773.250 658.050 774.150 ;
        RECT 658.950 772.950 661.050 775.050 ;
        RECT 649.950 769.950 652.050 772.050 ;
        RECT 653.250 770.250 654.750 771.150 ;
        RECT 655.950 769.950 658.050 772.050 ;
        RECT 650.400 766.050 651.450 769.950 ;
        RECT 652.950 766.950 655.050 769.050 ;
        RECT 643.950 763.950 646.050 766.050 ;
        RECT 649.950 763.950 652.050 766.050 ;
        RECT 656.400 760.050 657.450 769.950 ;
        RECT 659.400 769.050 660.450 772.950 ;
        RECT 662.400 771.450 663.450 775.950 ;
        RECT 664.950 773.250 666.750 774.150 ;
        RECT 667.950 772.950 670.050 775.050 ;
        RECT 673.950 774.450 676.050 775.050 ;
        RECT 677.400 774.450 678.450 778.950 ;
        RECT 683.400 775.050 684.450 812.400 ;
        RECT 688.950 812.250 690.750 813.150 ;
        RECT 691.950 811.950 694.050 814.050 ;
        RECT 695.250 812.250 697.050 813.150 ;
        RECT 697.950 811.950 700.050 814.050 ;
        RECT 700.950 812.250 702.750 813.150 ;
        RECT 703.950 811.950 706.050 814.050 ;
        RECT 707.250 812.250 709.050 813.150 ;
        RECT 688.950 808.950 691.050 811.050 ;
        RECT 692.250 809.850 693.750 810.750 ;
        RECT 694.950 810.450 697.050 811.050 ;
        RECT 698.400 810.450 699.450 811.950 ;
        RECT 694.950 809.400 699.450 810.450 ;
        RECT 694.950 808.950 697.050 809.400 ;
        RECT 700.950 808.950 703.050 811.050 ;
        RECT 704.250 809.850 705.750 810.750 ;
        RECT 706.950 808.950 709.050 811.050 ;
        RECT 713.400 810.450 714.450 814.950 ;
        RECT 776.400 814.050 777.450 814.950 ;
        RECT 715.950 812.250 717.750 813.150 ;
        RECT 718.950 811.950 721.050 814.050 ;
        RECT 722.250 812.250 724.050 813.150 ;
        RECT 730.950 811.950 733.050 814.050 ;
        RECT 733.950 812.850 736.050 813.750 ;
        RECT 736.950 812.250 739.050 813.150 ;
        RECT 742.950 812.850 745.050 813.750 ;
        RECT 751.950 811.950 754.050 814.050 ;
        RECT 766.950 812.250 768.750 813.150 ;
        RECT 769.950 811.950 772.050 814.050 ;
        RECT 773.250 812.250 775.050 813.150 ;
        RECT 775.950 811.950 778.050 814.050 ;
        RECT 715.950 810.450 718.050 811.050 ;
        RECT 713.400 809.400 718.050 810.450 ;
        RECT 719.250 809.850 720.750 810.750 ;
        RECT 715.950 808.950 718.050 809.400 ;
        RECT 721.950 808.950 724.050 811.050 ;
        RECT 689.400 805.050 690.450 808.950 ;
        RECT 688.950 802.950 691.050 805.050 ;
        RECT 701.400 784.050 702.450 808.950 ;
        RECT 722.400 802.050 723.450 808.950 ;
        RECT 721.950 799.950 724.050 802.050 ;
        RECT 700.950 781.950 703.050 784.050 ;
        RECT 706.950 781.950 709.050 784.050 ;
        RECT 691.950 775.950 694.050 778.050 ;
        RECT 697.950 777.450 700.050 778.050 ;
        RECT 695.250 776.250 696.750 777.150 ;
        RECT 697.950 776.400 702.450 777.450 ;
        RECT 697.950 775.950 700.050 776.400 ;
        RECT 671.250 773.250 672.750 774.150 ;
        RECT 673.950 773.400 678.450 774.450 ;
        RECT 673.950 772.950 676.050 773.400 ;
        RECT 679.950 773.250 682.050 774.150 ;
        RECT 682.950 772.950 685.050 775.050 ;
        RECT 685.950 773.250 688.050 774.150 ;
        RECT 691.950 773.850 693.750 774.750 ;
        RECT 694.950 772.950 697.050 775.050 ;
        RECT 698.250 773.850 700.050 774.750 ;
        RECT 664.950 771.450 667.050 772.050 ;
        RECT 662.400 770.400 667.050 771.450 ;
        RECT 668.250 770.850 669.750 771.750 ;
        RECT 658.950 766.950 661.050 769.050 ;
        RECT 655.950 757.950 658.050 760.050 ;
        RECT 640.950 754.950 643.050 757.050 ;
        RECT 652.950 754.950 655.050 757.050 ;
        RECT 640.950 751.950 643.050 754.050 ;
        RECT 643.950 751.950 646.050 754.050 ;
        RECT 631.950 740.250 633.750 741.150 ;
        RECT 634.950 739.950 637.050 742.050 ;
        RECT 638.250 740.250 640.050 741.150 ;
        RECT 631.950 736.950 634.050 739.050 ;
        RECT 635.250 737.850 636.750 738.750 ;
        RECT 637.950 738.450 640.050 739.050 ;
        RECT 641.400 738.450 642.450 751.950 ;
        RECT 644.400 748.050 645.450 751.950 ;
        RECT 643.950 745.950 646.050 748.050 ;
        RECT 643.950 743.850 646.050 744.750 ;
        RECT 646.950 743.250 649.050 744.150 ;
        RECT 649.950 742.950 652.050 745.050 ;
        RECT 646.950 741.450 649.050 742.050 ;
        RECT 650.400 741.450 651.450 742.950 ;
        RECT 646.950 740.400 651.450 741.450 ;
        RECT 646.950 739.950 649.050 740.400 ;
        RECT 637.950 737.400 642.450 738.450 ;
        RECT 637.950 736.950 640.050 737.400 ;
        RECT 653.400 736.050 654.450 754.950 ;
        RECT 662.400 748.050 663.450 770.400 ;
        RECT 664.950 769.950 667.050 770.400 ;
        RECT 670.950 769.950 673.050 772.050 ;
        RECT 676.950 769.950 679.050 772.050 ;
        RECT 679.950 769.950 682.050 772.050 ;
        RECT 683.250 770.250 684.750 771.150 ;
        RECT 685.950 769.950 688.050 772.050 ;
        RECT 671.400 769.050 672.450 769.950 ;
        RECT 670.950 766.950 673.050 769.050 ;
        RECT 677.400 766.050 678.450 769.950 ;
        RECT 676.950 763.950 679.050 766.050 ;
        RECT 680.400 754.050 681.450 769.950 ;
        RECT 682.950 766.950 685.050 769.050 ;
        RECT 683.400 766.050 684.450 766.950 ;
        RECT 686.400 766.050 687.450 769.950 ;
        RECT 682.950 763.950 685.050 766.050 ;
        RECT 685.950 763.950 688.050 766.050 ;
        RECT 679.950 751.950 682.050 754.050 ;
        RECT 661.950 745.950 664.050 748.050 ;
        RECT 673.950 745.950 676.050 748.050 ;
        RECT 679.950 745.950 682.050 748.050 ;
        RECT 658.950 742.950 661.050 745.050 ;
        RECT 664.950 742.950 667.050 745.050 ;
        RECT 659.400 742.050 660.450 742.950 ;
        RECT 665.400 742.050 666.450 742.950 ;
        RECT 658.950 739.950 661.050 742.050 ;
        RECT 664.950 739.950 667.050 742.050 ;
        RECT 668.250 740.250 670.050 741.150 ;
        RECT 658.950 737.850 660.750 738.750 ;
        RECT 661.950 736.950 664.050 739.050 ;
        RECT 665.250 737.850 666.750 738.750 ;
        RECT 667.950 736.950 670.050 739.050 ;
        RECT 646.950 733.950 649.050 736.050 ;
        RECT 652.950 733.950 655.050 736.050 ;
        RECT 661.950 734.850 664.050 735.750 ;
        RECT 647.400 727.050 648.450 733.950 ;
        RECT 646.950 724.950 649.050 727.050 ;
        RECT 655.950 724.950 658.050 727.050 ;
        RECT 631.950 711.450 634.050 712.050 ;
        RECT 634.950 711.450 637.050 712.050 ;
        RECT 631.950 710.400 637.050 711.450 ;
        RECT 631.950 709.950 634.050 710.400 ;
        RECT 634.950 709.950 637.050 710.400 ;
        RECT 637.950 709.950 640.050 712.050 ;
        RECT 631.950 706.950 634.050 709.050 ;
        RECT 632.400 706.050 633.450 706.950 ;
        RECT 638.400 706.050 639.450 709.950 ;
        RECT 647.400 706.050 648.450 724.950 ;
        RECT 631.950 703.950 634.050 706.050 ;
        RECT 635.250 704.250 636.750 705.150 ;
        RECT 637.950 703.950 640.050 706.050 ;
        RECT 646.950 703.950 649.050 706.050 ;
        RECT 652.950 705.450 655.050 706.050 ;
        RECT 656.400 705.450 657.450 724.950 ;
        RECT 674.400 711.450 675.450 745.950 ;
        RECT 680.400 742.050 681.450 745.950 ;
        RECT 695.400 745.050 696.450 772.950 ;
        RECT 701.400 769.050 702.450 776.400 ;
        RECT 700.950 766.950 703.050 769.050 ;
        RECT 707.400 760.050 708.450 781.950 ;
        RECT 731.400 781.050 732.450 811.950 ;
        RECT 779.400 811.050 780.450 814.950 ;
        RECT 781.950 811.950 784.050 814.050 ;
        RECT 785.250 812.250 787.050 813.150 ;
        RECT 736.950 808.950 739.050 811.050 ;
        RECT 748.950 808.950 751.050 811.050 ;
        RECT 766.950 808.950 769.050 811.050 ;
        RECT 770.250 809.850 771.750 810.750 ;
        RECT 772.950 808.950 775.050 811.050 ;
        RECT 775.950 809.850 777.750 810.750 ;
        RECT 778.950 808.950 781.050 811.050 ;
        RECT 782.250 809.850 783.750 810.750 ;
        RECT 784.950 808.950 787.050 811.050 ;
        RECT 737.400 808.050 738.450 808.950 ;
        RECT 736.950 805.950 739.050 808.050 ;
        RECT 730.950 780.450 733.050 781.050 ;
        RECT 724.950 779.250 727.050 780.150 ;
        RECT 730.950 779.400 735.450 780.450 ;
        RECT 730.950 778.950 733.050 779.400 ;
        RECT 709.950 775.950 712.050 778.050 ;
        RECT 721.950 776.250 723.750 777.150 ;
        RECT 724.950 775.950 727.050 778.050 ;
        RECT 728.250 776.250 729.750 777.150 ;
        RECT 730.950 775.950 733.050 778.050 ;
        RECT 710.400 775.050 711.450 775.950 ;
        RECT 709.950 772.950 712.050 775.050 ;
        RECT 721.950 772.950 724.050 775.050 ;
        RECT 725.400 772.050 726.450 775.950 ;
        RECT 734.400 775.050 735.450 779.400 ;
        RECT 736.950 775.950 739.050 778.050 ;
        RECT 742.950 777.450 745.050 778.050 ;
        RECT 740.250 776.250 741.750 777.150 ;
        RECT 742.950 776.400 747.450 777.450 ;
        RECT 742.950 775.950 745.050 776.400 ;
        RECT 727.950 772.950 730.050 775.050 ;
        RECT 731.250 773.850 733.050 774.750 ;
        RECT 733.950 772.950 736.050 775.050 ;
        RECT 736.950 773.850 738.750 774.750 ;
        RECT 739.950 772.950 742.050 775.050 ;
        RECT 743.250 773.850 745.050 774.750 ;
        RECT 709.950 770.850 712.050 771.750 ;
        RECT 712.950 770.250 715.050 771.150 ;
        RECT 724.950 769.950 727.050 772.050 ;
        RECT 712.950 766.950 715.050 769.050 ;
        RECT 713.400 766.050 714.450 766.950 ;
        RECT 712.950 763.950 715.050 766.050 ;
        RECT 724.950 763.950 727.050 766.050 ;
        RECT 706.950 757.950 709.050 760.050 ;
        RECT 709.950 747.450 712.050 748.050 ;
        RECT 707.400 746.400 712.050 747.450 ;
        RECT 688.950 744.450 691.050 745.050 ;
        RECT 686.400 743.400 691.050 744.450 ;
        RECT 686.400 742.050 687.450 743.400 ;
        RECT 688.950 742.950 691.050 743.400 ;
        RECT 694.950 742.950 697.050 745.050 ;
        RECT 697.950 744.450 700.050 745.050 ;
        RECT 697.950 743.400 702.450 744.450 ;
        RECT 697.950 742.950 700.050 743.400 ;
        RECT 676.950 740.250 678.750 741.150 ;
        RECT 679.950 739.950 682.050 742.050 ;
        RECT 683.250 740.250 685.050 741.150 ;
        RECT 685.950 739.950 688.050 742.050 ;
        RECT 688.950 740.850 691.050 741.750 ;
        RECT 694.950 740.250 697.050 741.150 ;
        RECT 697.950 740.850 700.050 741.750 ;
        RECT 676.950 736.950 679.050 739.050 ;
        RECT 680.250 737.850 681.750 738.750 ;
        RECT 682.950 738.450 685.050 739.050 ;
        RECT 686.400 738.450 687.450 739.950 ;
        RECT 682.950 737.400 687.450 738.450 ;
        RECT 682.950 736.950 685.050 737.400 ;
        RECT 694.950 736.950 697.050 739.050 ;
        RECT 688.950 733.950 691.050 736.050 ;
        RECT 674.400 710.400 678.450 711.450 ;
        RECT 667.950 707.250 670.050 708.150 ;
        RECT 673.950 706.950 676.050 709.050 ;
        RECT 661.950 705.450 664.050 706.050 ;
        RECT 650.250 704.250 651.750 705.150 ;
        RECT 652.950 704.400 657.450 705.450 ;
        RECT 652.950 703.950 655.050 704.400 ;
        RECT 628.950 700.950 631.050 703.050 ;
        RECT 631.950 701.850 633.750 702.750 ;
        RECT 634.950 700.950 637.050 703.050 ;
        RECT 638.250 701.850 640.050 702.750 ;
        RECT 646.950 701.850 648.750 702.750 ;
        RECT 649.950 700.950 652.050 703.050 ;
        RECT 653.250 701.850 655.050 702.750 ;
        RECT 628.950 697.950 631.050 700.050 ;
        RECT 629.400 697.050 630.450 697.950 ;
        RECT 650.400 697.050 651.450 700.950 ;
        RECT 656.400 700.050 657.450 704.400 ;
        RECT 659.400 704.400 664.050 705.450 ;
        RECT 655.950 697.950 658.050 700.050 ;
        RECT 628.950 694.950 631.050 697.050 ;
        RECT 631.950 694.950 634.050 697.050 ;
        RECT 649.950 694.950 652.050 697.050 ;
        RECT 625.950 682.950 628.050 685.050 ;
        RECT 622.950 673.950 625.050 676.050 ;
        RECT 619.950 670.950 622.050 673.050 ;
        RECT 625.950 672.450 628.050 673.050 ;
        RECT 623.250 671.250 624.750 672.150 ;
        RECT 625.950 671.400 630.450 672.450 ;
        RECT 625.950 670.950 628.050 671.400 ;
        RECT 616.950 667.950 619.050 670.050 ;
        RECT 620.250 668.850 621.750 669.750 ;
        RECT 622.950 667.950 625.050 670.050 ;
        RECT 626.250 668.850 628.050 669.750 ;
        RECT 616.950 665.850 619.050 666.750 ;
        RECT 616.950 661.950 619.050 664.050 ;
        RECT 605.400 635.400 609.450 636.450 ;
        RECT 572.400 622.050 573.450 632.400 ;
        RECT 574.950 631.950 577.050 632.400 ;
        RECT 578.250 632.250 579.750 633.150 ;
        RECT 580.950 632.400 585.450 633.450 ;
        RECT 580.950 631.950 583.050 632.400 ;
        RECT 574.950 629.850 576.750 630.750 ;
        RECT 577.950 628.950 580.050 631.050 ;
        RECT 581.250 629.850 583.050 630.750 ;
        RECT 571.950 619.950 574.050 622.050 ;
        RECT 578.400 619.050 579.450 628.950 ;
        RECT 584.400 625.050 585.450 632.400 ;
        RECT 583.950 622.950 586.050 625.050 ;
        RECT 577.950 616.950 580.050 619.050 ;
        RECT 568.950 604.950 571.050 607.050 ;
        RECT 562.950 601.950 565.050 604.050 ;
        RECT 565.950 601.950 568.050 604.050 ;
        RECT 571.950 601.950 574.050 604.050 ;
        RECT 563.400 601.050 564.450 601.950 ;
        RECT 572.400 601.050 573.450 601.950 ;
        RECT 559.950 598.950 562.050 601.050 ;
        RECT 562.950 598.950 565.050 601.050 ;
        RECT 566.250 599.850 567.750 600.750 ;
        RECT 568.950 598.950 571.050 601.050 ;
        RECT 571.950 598.950 574.050 601.050 ;
        RECT 575.250 599.250 576.750 600.150 ;
        RECT 577.950 598.950 580.050 601.050 ;
        RECT 562.950 596.850 565.050 597.750 ;
        RECT 568.950 596.850 571.050 597.750 ;
        RECT 571.950 596.850 573.750 597.750 ;
        RECT 574.950 595.950 577.050 598.050 ;
        RECT 578.250 596.850 579.750 597.750 ;
        RECT 580.950 595.950 583.050 598.050 ;
        RECT 580.950 593.850 583.050 594.750 ;
        RECT 577.950 571.950 580.050 574.050 ;
        RECT 559.950 563.250 562.050 564.150 ;
        RECT 556.950 560.250 558.750 561.150 ;
        RECT 559.950 559.950 562.050 562.050 ;
        RECT 563.250 560.250 564.750 561.150 ;
        RECT 565.950 559.950 568.050 562.050 ;
        RECT 560.400 559.050 561.450 559.950 ;
        RECT 556.950 556.950 559.050 559.050 ;
        RECT 559.950 556.950 562.050 559.050 ;
        RECT 562.950 556.950 565.050 559.050 ;
        RECT 566.250 557.850 568.050 558.750 ;
        RECT 574.950 556.950 577.050 559.050 ;
        RECT 557.400 535.050 558.450 556.950 ;
        RECT 575.400 553.050 576.450 556.950 ;
        RECT 565.950 550.950 568.050 553.050 ;
        RECT 574.950 550.950 577.050 553.050 ;
        RECT 559.950 538.950 562.050 541.050 ;
        RECT 556.950 532.950 559.050 535.050 ;
        RECT 541.950 529.950 544.050 532.050 ;
        RECT 553.950 529.950 556.050 532.050 ;
        RECT 532.950 526.950 535.050 529.050 ;
        RECT 533.400 526.050 534.450 526.950 ;
        RECT 532.950 523.950 535.050 526.050 ;
        RECT 536.250 524.250 538.050 525.150 ;
        RECT 526.950 521.850 528.750 522.750 ;
        RECT 529.950 520.950 532.050 523.050 ;
        RECT 533.250 521.850 534.750 522.750 ;
        RECT 535.950 520.950 538.050 523.050 ;
        RECT 529.950 518.850 532.050 519.750 ;
        RECT 524.400 500.400 528.450 501.450 ;
        RECT 521.100 497.100 523.200 499.200 ;
        RECT 505.950 494.400 508.050 496.500 ;
        RECT 510.000 494.400 512.100 496.500 ;
        RECT 517.950 494.850 520.050 496.950 ;
        RECT 506.250 488.250 507.450 494.400 ;
        RECT 502.950 484.950 505.050 487.050 ;
        RECT 505.950 486.150 508.050 488.250 ;
        RECT 502.950 482.250 505.050 483.150 ;
        RECT 502.950 478.950 505.050 481.050 ;
        RECT 503.400 475.050 504.450 478.950 ;
        RECT 506.250 477.600 507.450 486.150 ;
        RECT 510.450 485.550 511.650 494.400 ;
        RECT 514.950 491.250 517.050 493.350 ;
        RECT 510.150 483.450 512.250 485.550 ;
        RECT 510.450 477.600 511.650 483.450 ;
        RECT 515.400 477.600 516.600 491.250 ;
        RECT 518.550 477.600 519.750 494.850 ;
        RECT 521.250 493.350 522.450 497.100 ;
        RECT 523.950 493.950 526.050 496.050 ;
        RECT 520.950 491.250 523.050 493.350 ;
        RECT 521.250 477.600 522.450 491.250 ;
        RECT 505.950 475.500 508.050 477.600 ;
        RECT 510.150 475.500 512.250 477.600 ;
        RECT 514.950 475.500 517.050 477.600 ;
        RECT 517.950 475.500 520.050 477.600 ;
        RECT 520.950 475.500 523.050 477.600 ;
        RECT 502.950 472.950 505.050 475.050 ;
        RECT 502.950 469.950 505.050 472.050 ;
        RECT 503.400 457.050 504.450 469.950 ;
        RECT 520.950 466.950 523.050 469.050 ;
        RECT 517.950 457.950 520.050 460.050 ;
        RECT 496.950 454.950 499.050 457.050 ;
        RECT 499.950 454.950 502.050 457.050 ;
        RECT 502.950 454.950 505.050 457.050 ;
        RECT 490.950 451.950 493.050 454.050 ;
        RECT 494.250 452.250 496.050 453.150 ;
        RECT 484.950 449.850 486.750 450.750 ;
        RECT 487.950 448.950 490.050 451.050 ;
        RECT 491.250 449.850 492.750 450.750 ;
        RECT 493.950 448.950 496.050 451.050 ;
        RECT 487.950 446.850 490.050 447.750 ;
        RECT 484.950 442.950 487.050 445.050 ;
        RECT 485.400 427.050 486.450 442.950 ;
        RECT 484.950 424.950 487.050 427.050 ;
        RECT 481.950 421.950 484.050 424.050 ;
        RECT 481.950 418.950 484.050 421.050 ;
        RECT 487.950 418.950 490.050 421.050 ;
        RECT 475.950 409.950 478.050 412.050 ;
        RECT 472.950 406.950 475.050 409.050 ;
        RECT 482.400 397.050 483.450 418.950 ;
        RECT 488.400 415.050 489.450 418.950 ;
        RECT 493.950 416.250 496.050 417.150 ;
        RECT 484.950 413.250 486.750 414.150 ;
        RECT 487.950 412.950 490.050 415.050 ;
        RECT 491.250 413.250 492.750 414.150 ;
        RECT 493.950 412.950 496.050 415.050 ;
        RECT 484.950 409.950 487.050 412.050 ;
        RECT 488.250 410.850 489.750 411.750 ;
        RECT 490.950 409.950 493.050 412.050 ;
        RECT 491.400 409.050 492.450 409.950 ;
        RECT 490.950 406.950 493.050 409.050 ;
        RECT 484.950 403.950 487.050 406.050 ;
        RECT 481.950 394.950 484.050 397.050 ;
        RECT 469.950 388.950 472.050 391.050 ;
        RECT 481.950 388.950 484.050 391.050 ;
        RECT 482.400 388.050 483.450 388.950 ;
        RECT 475.950 385.950 478.050 388.050 ;
        RECT 481.950 385.950 484.050 388.050 ;
        RECT 457.950 382.950 460.050 385.050 ;
        RECT 460.950 382.950 463.050 385.050 ;
        RECT 469.950 382.950 472.050 385.050 ;
        RECT 458.400 381.450 459.450 382.950 ;
        RECT 460.950 381.450 463.050 382.050 ;
        RECT 458.400 380.400 463.050 381.450 ;
        RECT 460.950 379.950 463.050 380.400 ;
        RECT 466.950 380.250 469.050 381.150 ;
        RECT 460.950 377.850 463.050 378.750 ;
        RECT 463.950 376.950 466.050 379.050 ;
        RECT 457.950 373.950 460.050 376.050 ;
        RECT 424.800 367.800 426.900 369.900 ;
        RECT 448.950 367.950 451.050 370.050 ;
        RECT 451.950 367.950 454.050 370.050 ;
        RECT 454.950 367.950 457.050 370.050 ;
        RECT 436.950 358.950 439.050 361.050 ;
        RECT 445.950 358.950 448.050 361.050 ;
        RECT 433.950 355.950 436.050 358.050 ;
        RECT 409.950 343.950 412.050 346.050 ;
        RECT 418.950 343.950 421.050 346.050 ;
        RECT 409.950 341.250 412.050 342.150 ;
        RECT 415.950 341.250 418.050 342.150 ;
        RECT 409.950 339.450 412.050 340.050 ;
        RECT 407.400 338.400 412.050 339.450 ;
        RECT 397.950 334.950 400.050 337.050 ;
        RECT 400.950 334.950 403.050 337.050 ;
        RECT 394.950 319.950 397.050 322.050 ;
        RECT 394.950 316.950 397.050 319.050 ;
        RECT 391.950 310.950 394.050 313.050 ;
        RECT 395.400 310.050 396.450 316.950 ;
        RECT 398.400 313.050 399.450 334.950 ;
        RECT 401.400 331.050 402.450 334.950 ;
        RECT 404.400 331.050 405.450 337.950 ;
        RECT 400.950 328.950 403.050 331.050 ;
        RECT 403.950 328.950 406.050 331.050 ;
        RECT 407.400 328.050 408.450 338.400 ;
        RECT 409.950 337.950 412.050 338.400 ;
        RECT 413.250 338.250 414.750 339.150 ;
        RECT 415.950 337.950 418.050 340.050 ;
        RECT 412.950 334.950 415.050 337.050 ;
        RECT 409.950 331.950 412.050 334.050 ;
        RECT 406.950 325.950 409.050 328.050 ;
        RECT 397.950 310.950 400.050 313.050 ;
        RECT 403.950 312.450 406.050 313.050 ;
        RECT 401.250 311.250 402.750 312.150 ;
        RECT 403.950 311.400 408.450 312.450 ;
        RECT 403.950 310.950 406.050 311.400 ;
        RECT 379.950 308.250 381.750 309.150 ;
        RECT 382.950 307.950 385.050 310.050 ;
        RECT 386.250 308.250 388.050 309.150 ;
        RECT 394.950 307.950 397.050 310.050 ;
        RECT 398.250 308.850 399.750 309.750 ;
        RECT 400.950 307.950 403.050 310.050 ;
        RECT 404.250 308.850 406.050 309.750 ;
        RECT 379.950 304.950 382.050 307.050 ;
        RECT 383.250 305.850 384.750 306.750 ;
        RECT 385.950 304.950 388.050 307.050 ;
        RECT 394.950 305.850 397.050 306.750 ;
        RECT 380.400 304.050 381.450 304.950 ;
        RECT 379.950 301.950 382.050 304.050 ;
        RECT 385.950 301.950 388.050 304.050 ;
        RECT 394.950 301.950 397.050 304.050 ;
        RECT 386.400 280.050 387.450 301.950 ;
        RECT 388.950 295.950 391.050 298.050 ;
        RECT 379.950 277.950 382.050 280.050 ;
        RECT 385.950 277.950 388.050 280.050 ;
        RECT 376.950 273.450 379.050 274.050 ;
        RECT 374.400 272.400 379.050 273.450 ;
        RECT 374.400 271.050 375.450 272.400 ;
        RECT 376.950 271.950 379.050 272.400 ;
        RECT 367.950 268.950 370.050 271.050 ;
        RECT 370.950 269.250 372.750 270.150 ;
        RECT 373.950 268.950 376.050 271.050 ;
        RECT 376.950 268.950 379.050 271.050 ;
        RECT 367.950 265.950 370.050 268.050 ;
        RECT 370.950 265.950 373.050 268.050 ;
        RECT 374.250 266.850 376.050 267.750 ;
        RECT 364.950 262.950 367.050 265.050 ;
        RECT 368.400 261.450 369.450 265.950 ;
        RECT 371.400 264.450 372.450 265.950 ;
        RECT 371.400 263.400 375.450 264.450 ;
        RECT 365.400 260.400 369.450 261.450 ;
        RECT 365.400 241.050 366.450 260.400 ;
        RECT 370.950 259.950 373.050 262.050 ;
        RECT 367.950 253.950 370.050 256.050 ;
        RECT 364.950 238.950 367.050 241.050 ;
        RECT 364.950 235.950 367.050 238.050 ;
        RECT 364.950 233.850 367.050 234.750 ;
        RECT 368.400 232.050 369.450 253.950 ;
        RECT 362.400 230.400 366.450 231.450 ;
        RECT 359.400 227.400 363.450 228.450 ;
        RECT 335.400 212.400 339.450 213.450 ;
        RECT 335.400 175.050 336.450 212.400 ;
        RECT 340.950 203.250 343.050 204.150 ;
        RECT 346.950 202.950 349.050 205.050 ;
        RECT 347.400 202.050 348.450 202.950 ;
        RECT 337.950 200.250 339.750 201.150 ;
        RECT 340.950 199.950 343.050 202.050 ;
        RECT 344.250 200.250 345.750 201.150 ;
        RECT 346.950 199.950 349.050 202.050 ;
        RECT 337.950 196.950 340.050 199.050 ;
        RECT 341.400 196.050 342.450 199.950 ;
        RECT 343.950 196.950 346.050 199.050 ;
        RECT 347.250 197.850 349.050 198.750 ;
        RECT 340.950 193.950 343.050 196.050 ;
        RECT 334.950 172.950 337.050 175.050 ;
        RECT 341.400 172.050 342.450 193.950 ;
        RECT 344.400 193.050 345.450 196.950 ;
        RECT 343.950 190.950 346.050 193.050 ;
        RECT 346.950 187.950 349.050 190.050 ;
        RECT 334.950 169.950 337.050 172.050 ;
        RECT 340.950 169.950 343.050 172.050 ;
        RECT 328.950 163.950 331.050 166.050 ;
        RECT 331.950 163.950 334.050 166.050 ;
        RECT 325.950 160.950 328.050 163.050 ;
        RECT 326.400 160.050 327.450 160.950 ;
        RECT 329.400 160.050 330.450 163.950 ;
        RECT 335.400 163.050 336.450 169.950 ;
        RECT 347.400 169.050 348.450 187.950 ;
        RECT 350.400 169.050 351.450 223.950 ;
        RECT 356.100 223.800 358.200 225.900 ;
        RECT 358.950 214.950 361.050 217.050 ;
        RECT 352.950 205.950 355.050 208.050 ;
        RECT 353.400 199.050 354.450 205.950 ;
        RECT 359.400 199.050 360.450 214.950 ;
        RECT 362.400 214.050 363.450 227.400 ;
        RECT 361.950 211.950 364.050 214.050 ;
        RECT 365.400 202.050 366.450 230.400 ;
        RECT 367.950 229.950 370.050 232.050 ;
        RECT 371.400 228.450 372.450 259.950 ;
        RECT 368.400 227.400 372.450 228.450 ;
        RECT 364.950 199.950 367.050 202.050 ;
        RECT 352.950 196.950 355.050 199.050 ;
        RECT 358.950 196.950 361.050 199.050 ;
        RECT 362.250 197.250 364.050 198.150 ;
        RECT 364.950 196.950 367.050 199.050 ;
        RECT 352.950 194.850 355.050 195.750 ;
        RECT 355.950 194.250 358.050 195.150 ;
        RECT 358.950 194.850 360.750 195.750 ;
        RECT 361.950 193.950 364.050 196.050 ;
        RECT 352.950 190.950 355.050 193.050 ;
        RECT 355.950 190.950 358.050 193.050 ;
        RECT 337.950 167.250 340.050 168.150 ;
        RECT 340.950 167.850 343.050 168.750 ;
        RECT 343.950 167.250 345.750 168.150 ;
        RECT 346.950 166.950 349.050 169.050 ;
        RECT 349.950 166.950 352.050 169.050 ;
        RECT 337.950 163.950 340.050 166.050 ;
        RECT 343.950 163.950 346.050 166.050 ;
        RECT 347.250 164.850 349.050 165.750 ;
        RECT 349.950 163.950 352.050 166.050 ;
        RECT 331.950 160.950 334.050 163.050 ;
        RECT 334.950 160.950 337.050 163.050 ;
        RECT 325.950 157.950 328.050 160.050 ;
        RECT 328.950 157.950 331.050 160.050 ;
        RECT 325.950 154.950 328.050 157.050 ;
        RECT 316.950 120.450 319.050 121.050 ;
        RECT 311.400 119.400 319.050 120.450 ;
        RECT 295.950 112.950 298.050 115.050 ;
        RECT 292.950 97.950 295.050 100.050 ;
        RECT 296.400 97.050 297.450 112.950 ;
        RECT 301.950 103.950 304.050 106.050 ;
        RECT 289.950 94.950 292.050 97.050 ;
        RECT 293.250 95.250 294.750 96.150 ;
        RECT 295.950 94.950 298.050 97.050 ;
        RECT 289.950 92.850 291.750 93.750 ;
        RECT 292.950 91.950 295.050 94.050 ;
        RECT 296.250 92.850 297.750 93.750 ;
        RECT 298.950 91.950 301.050 94.050 ;
        RECT 298.950 89.850 301.050 90.750 ;
        RECT 298.950 85.950 301.050 88.050 ;
        RECT 286.950 58.950 289.050 61.050 ;
        RECT 289.950 59.250 292.050 60.150 ;
        RECT 295.950 58.950 298.050 61.050 ;
        RECT 265.950 55.950 268.050 58.050 ;
        RECT 268.950 55.950 271.050 58.050 ;
        RECT 274.950 57.450 277.050 58.050 ;
        RECT 272.250 56.250 273.750 57.150 ;
        RECT 274.950 56.400 279.450 57.450 ;
        RECT 274.950 55.950 277.050 56.400 ;
        RECT 259.950 52.950 262.050 55.050 ;
        RECT 259.950 50.850 262.050 51.750 ;
        RECT 262.950 50.250 265.050 51.150 ;
        RECT 256.950 46.950 259.050 49.050 ;
        RECT 262.950 48.450 265.050 49.050 ;
        RECT 266.400 48.450 267.450 55.950 ;
        RECT 268.950 53.850 270.750 54.750 ;
        RECT 271.950 52.950 274.050 55.050 ;
        RECT 275.250 53.850 277.050 54.750 ;
        RECT 278.400 52.050 279.450 56.400 ;
        RECT 283.950 55.950 286.050 58.050 ;
        RECT 287.250 56.250 288.750 57.150 ;
        RECT 289.950 55.950 292.050 58.050 ;
        RECT 293.250 56.250 295.050 57.150 ;
        RECT 283.950 53.850 285.750 54.750 ;
        RECT 286.950 52.950 289.050 55.050 ;
        RECT 287.400 52.050 288.450 52.950 ;
        RECT 277.950 49.950 280.050 52.050 ;
        RECT 286.950 49.950 289.050 52.050 ;
        RECT 262.950 47.400 267.450 48.450 ;
        RECT 262.950 46.950 265.050 47.400 ;
        RECT 286.950 46.950 289.050 49.050 ;
        RECT 257.400 25.050 258.450 46.950 ;
        RECT 274.950 40.950 277.050 43.050 ;
        RECT 262.950 31.950 265.050 34.050 ;
        RECT 263.400 25.050 264.450 31.950 ;
        RECT 256.950 22.950 259.050 25.050 ;
        RECT 260.250 23.250 261.750 24.150 ;
        RECT 262.950 22.950 265.050 25.050 ;
        RECT 247.950 20.400 252.450 21.450 ;
        RECT 247.950 19.950 250.050 20.400 ;
        RECT 253.950 19.950 256.050 22.050 ;
        RECT 256.950 20.850 258.750 21.750 ;
        RECT 259.950 19.950 262.050 22.050 ;
        RECT 263.250 20.850 264.750 21.750 ;
        RECT 265.950 19.950 268.050 22.050 ;
        RECT 235.950 17.850 238.050 18.750 ;
        RECT 265.950 17.850 268.050 18.750 ;
        RECT 275.400 18.450 276.450 40.950 ;
        RECT 287.400 40.050 288.450 46.950 ;
        RECT 290.400 40.050 291.450 55.950 ;
        RECT 292.950 54.450 295.050 55.050 ;
        RECT 296.400 54.450 297.450 58.950 ;
        RECT 299.400 55.050 300.450 85.950 ;
        RECT 302.400 57.450 303.450 103.950 ;
        RECT 304.950 100.950 307.050 103.050 ;
        RECT 305.400 70.050 306.450 100.950 ;
        RECT 314.400 97.050 315.450 119.400 ;
        RECT 316.950 118.950 319.050 119.400 ;
        RECT 322.950 118.950 325.050 121.050 ;
        RECT 319.950 106.950 322.050 109.050 ;
        RECT 316.950 97.950 319.050 100.050 ;
        RECT 307.950 94.950 310.050 97.050 ;
        RECT 311.250 95.250 312.750 96.150 ;
        RECT 313.950 94.950 316.050 97.050 ;
        RECT 317.400 94.050 318.450 97.950 ;
        RECT 307.950 92.850 309.750 93.750 ;
        RECT 310.950 91.950 313.050 94.050 ;
        RECT 314.250 92.850 315.750 93.750 ;
        RECT 316.950 91.950 319.050 94.050 ;
        RECT 311.400 90.450 312.450 91.950 ;
        RECT 308.400 89.400 312.450 90.450 ;
        RECT 316.950 89.850 319.050 90.750 ;
        RECT 304.950 67.950 307.050 70.050 ;
        RECT 302.400 56.400 306.450 57.450 ;
        RECT 292.950 53.400 297.450 54.450 ;
        RECT 292.950 52.950 295.050 53.400 ;
        RECT 296.400 52.050 297.450 53.400 ;
        RECT 298.950 52.950 301.050 55.050 ;
        RECT 301.950 52.950 304.050 55.050 ;
        RECT 295.950 49.950 298.050 52.050 ;
        RECT 298.950 50.250 301.050 51.150 ;
        RECT 301.950 50.850 304.050 51.750 ;
        RECT 298.950 46.950 301.050 49.050 ;
        RECT 299.400 40.050 300.450 46.950 ;
        RECT 286.950 37.950 289.050 40.050 ;
        RECT 289.950 37.950 292.050 40.050 ;
        RECT 298.950 37.950 301.050 40.050 ;
        RECT 287.400 22.050 288.450 37.950 ;
        RECT 290.400 31.050 291.450 37.950 ;
        RECT 299.400 34.050 300.450 37.950 ;
        RECT 298.950 31.950 301.050 34.050 ;
        RECT 289.950 28.950 292.050 31.050 ;
        RECT 298.950 28.950 301.050 31.050 ;
        RECT 292.950 25.950 295.050 28.050 ;
        RECT 295.950 25.950 298.050 28.050 ;
        RECT 293.400 25.050 294.450 25.950 ;
        RECT 299.400 25.050 300.450 28.950 ;
        RECT 301.950 25.950 304.050 28.050 ;
        RECT 292.950 22.950 295.050 25.050 ;
        RECT 296.250 23.850 297.750 24.750 ;
        RECT 298.950 22.950 301.050 25.050 ;
        RECT 277.950 20.250 279.750 21.150 ;
        RECT 280.950 19.950 283.050 22.050 ;
        RECT 284.250 20.250 286.050 21.150 ;
        RECT 286.950 19.950 289.050 22.050 ;
        RECT 292.950 20.850 295.050 21.750 ;
        RECT 298.950 20.850 301.050 21.750 ;
        RECT 277.950 18.450 280.050 19.050 ;
        RECT 275.400 17.400 280.050 18.450 ;
        RECT 281.250 17.850 282.750 18.750 ;
        RECT 277.950 16.950 280.050 17.400 ;
        RECT 283.950 16.950 286.050 19.050 ;
        RECT 226.950 13.650 229.050 15.750 ;
        RECT 223.950 10.050 226.050 12.150 ;
        RECT 47.100 7.800 49.200 9.900 ;
        RECT 184.950 7.950 187.050 10.050 ;
        RECT 196.950 7.950 199.050 10.050 ;
        RECT 199.950 7.950 202.050 10.050 ;
        RECT 202.950 7.950 205.050 10.050 ;
        RECT 227.250 9.900 228.450 13.650 ;
        RECT 284.400 13.050 285.450 16.950 ;
        RECT 302.400 16.050 303.450 25.950 ;
        RECT 305.400 25.050 306.450 56.400 ;
        RECT 308.400 55.050 309.450 89.400 ;
        RECT 310.950 79.950 313.050 82.050 ;
        RECT 311.400 58.050 312.450 79.950 ;
        RECT 320.400 61.050 321.450 106.950 ;
        RECT 326.400 103.050 327.450 154.950 ;
        RECT 328.950 133.950 331.050 136.050 ;
        RECT 329.400 124.050 330.450 133.950 ;
        RECT 332.400 133.050 333.450 160.950 ;
        RECT 338.400 157.050 339.450 163.950 ;
        RECT 344.400 160.050 345.450 163.950 ;
        RECT 343.950 157.950 346.050 160.050 ;
        RECT 337.950 154.950 340.050 157.050 ;
        RECT 350.400 154.050 351.450 163.950 ;
        RECT 349.950 151.950 352.050 154.050 ;
        RECT 346.950 136.950 349.050 139.050 ;
        RECT 347.400 133.050 348.450 136.950 ;
        RECT 331.950 130.950 334.050 133.050 ;
        RECT 346.950 130.950 349.050 133.050 ;
        RECT 349.950 130.950 352.050 133.050 ;
        RECT 331.950 127.950 334.050 130.050 ;
        RECT 334.950 128.250 337.050 129.150 ;
        RECT 340.950 127.950 343.050 130.050 ;
        RECT 328.950 121.950 331.050 124.050 ;
        RECT 332.400 120.450 333.450 127.950 ;
        RECT 341.400 127.050 342.450 127.950 ;
        RECT 350.400 127.050 351.450 130.950 ;
        RECT 353.400 130.050 354.450 190.950 ;
        RECT 356.400 190.050 357.450 190.950 ;
        RECT 365.400 190.050 366.450 196.950 ;
        RECT 368.400 193.050 369.450 227.400 ;
        RECT 374.400 226.050 375.450 263.400 ;
        RECT 377.400 256.050 378.450 268.950 ;
        RECT 380.400 267.450 381.450 277.950 ;
        RECT 389.400 271.050 390.450 295.950 ;
        RECT 391.950 280.950 394.050 283.050 ;
        RECT 392.400 271.050 393.450 280.950 ;
        RECT 395.400 274.050 396.450 301.950 ;
        RECT 401.400 301.050 402.450 307.950 ;
        RECT 400.950 298.950 403.050 301.050 ;
        RECT 407.400 292.050 408.450 311.400 ;
        RECT 406.950 289.950 409.050 292.050 ;
        RECT 394.950 271.950 397.050 274.050 ;
        RECT 400.950 271.950 403.050 274.050 ;
        RECT 406.950 272.250 409.050 273.150 ;
        RECT 401.400 271.050 402.450 271.950 ;
        RECT 382.950 269.250 384.750 270.150 ;
        RECT 385.950 268.950 388.050 271.050 ;
        RECT 388.950 268.950 391.050 271.050 ;
        RECT 391.950 270.450 394.050 271.050 ;
        RECT 391.950 269.400 396.450 270.450 ;
        RECT 391.950 268.950 394.050 269.400 ;
        RECT 382.950 267.450 385.050 268.050 ;
        RECT 380.400 266.400 385.050 267.450 ;
        RECT 386.250 266.850 388.050 267.750 ;
        RECT 382.950 265.950 385.050 266.400 ;
        RECT 388.950 266.250 391.050 267.150 ;
        RECT 391.950 266.850 394.050 267.750 ;
        RECT 395.400 267.450 396.450 269.400 ;
        RECT 397.950 269.250 399.750 270.150 ;
        RECT 400.950 268.950 403.050 271.050 ;
        RECT 404.250 269.250 405.750 270.150 ;
        RECT 406.950 268.950 409.050 271.050 ;
        RECT 397.950 267.450 400.050 268.050 ;
        RECT 395.400 266.400 400.050 267.450 ;
        RECT 401.250 266.850 402.750 267.750 ;
        RECT 403.950 267.450 406.050 268.050 ;
        RECT 397.950 265.950 400.050 266.400 ;
        RECT 403.950 266.400 408.450 267.450 ;
        RECT 403.950 265.950 406.050 266.400 ;
        RECT 379.950 264.450 382.050 265.050 ;
        RECT 385.950 264.450 388.050 265.050 ;
        RECT 388.950 264.450 391.050 265.050 ;
        RECT 379.950 263.400 384.450 264.450 ;
        RECT 379.950 262.950 382.050 263.400 ;
        RECT 379.950 259.950 382.050 262.050 ;
        RECT 376.950 253.950 379.050 256.050 ;
        RECT 376.950 239.250 379.050 240.150 ;
        RECT 376.950 237.450 379.050 238.050 ;
        RECT 380.400 237.450 381.450 259.950 ;
        RECT 383.400 247.050 384.450 263.400 ;
        RECT 385.950 263.400 391.050 264.450 ;
        RECT 385.950 262.950 388.050 263.400 ;
        RECT 388.950 262.950 391.050 263.400 ;
        RECT 394.950 262.950 397.050 265.050 ;
        RECT 397.950 262.950 400.050 265.050 ;
        RECT 403.950 262.950 406.050 265.050 ;
        RECT 382.950 244.950 385.050 247.050 ;
        RECT 382.950 238.950 385.050 241.050 ;
        RECT 376.950 236.400 381.450 237.450 ;
        RECT 376.950 235.950 379.050 236.400 ;
        RECT 376.950 232.950 379.050 235.050 ;
        RECT 373.950 223.950 376.050 226.050 ;
        RECT 377.400 222.450 378.450 232.950 ;
        RECT 379.950 223.950 382.050 226.050 ;
        RECT 374.400 221.400 378.450 222.450 ;
        RECT 370.950 202.950 373.050 205.050 ;
        RECT 371.400 193.050 372.450 202.950 ;
        RECT 374.400 196.050 375.450 221.400 ;
        RECT 380.400 205.050 381.450 223.950 ;
        RECT 383.400 217.050 384.450 238.950 ;
        RECT 385.950 235.950 388.050 238.050 ;
        RECT 382.950 214.950 385.050 217.050 ;
        RECT 386.400 208.050 387.450 235.950 ;
        RECT 389.400 234.450 390.450 262.950 ;
        RECT 395.400 259.050 396.450 262.950 ;
        RECT 391.950 256.950 394.050 259.050 ;
        RECT 394.950 256.950 397.050 259.050 ;
        RECT 392.400 241.050 393.450 256.950 ;
        RECT 398.400 244.050 399.450 262.950 ;
        RECT 397.950 241.950 400.050 244.050 ;
        RECT 404.400 241.050 405.450 262.950 ;
        RECT 407.400 256.050 408.450 266.400 ;
        RECT 410.400 262.050 411.450 331.950 ;
        RECT 412.950 319.950 415.050 322.050 ;
        RECT 413.400 316.050 414.450 319.950 ;
        RECT 419.400 319.050 420.450 343.950 ;
        RECT 421.950 340.950 424.050 343.050 ;
        RECT 424.950 341.250 427.050 342.150 ;
        RECT 430.950 341.250 433.050 342.150 ;
        RECT 422.400 334.050 423.450 340.950 ;
        RECT 424.950 337.950 427.050 340.050 ;
        RECT 428.250 338.250 429.750 339.150 ;
        RECT 430.950 337.950 433.050 340.050 ;
        RECT 421.950 331.950 424.050 334.050 ;
        RECT 425.400 331.050 426.450 337.950 ;
        RECT 427.950 334.950 430.050 337.050 ;
        RECT 424.950 328.950 427.050 331.050 ;
        RECT 428.400 325.050 429.450 334.950 ;
        RECT 431.400 325.050 432.450 337.950 ;
        RECT 434.400 328.050 435.450 355.950 ;
        RECT 437.400 340.050 438.450 358.950 ;
        RECT 446.400 355.050 447.450 358.950 ;
        RECT 445.950 352.950 448.050 355.050 ;
        RECT 451.950 346.950 454.050 349.050 ;
        RECT 452.400 346.050 453.450 346.950 ;
        RECT 451.950 343.950 454.050 346.050 ;
        RECT 458.400 343.050 459.450 373.950 ;
        RECT 464.400 367.050 465.450 376.950 ;
        RECT 463.950 364.950 466.050 367.050 ;
        RECT 442.950 341.250 445.050 342.150 ;
        RECT 448.950 341.250 451.050 342.150 ;
        RECT 451.950 340.950 454.050 343.050 ;
        RECT 454.950 341.250 457.050 342.150 ;
        RECT 457.950 340.950 460.050 343.050 ;
        RECT 460.950 341.250 463.050 342.150 ;
        RECT 436.950 337.950 439.050 340.050 ;
        RECT 442.950 337.950 445.050 340.050 ;
        RECT 446.250 338.250 447.750 339.150 ;
        RECT 448.950 337.950 451.050 340.050 ;
        RECT 443.400 337.050 444.450 337.950 ;
        RECT 449.400 337.050 450.450 337.950 ;
        RECT 442.950 334.950 445.050 337.050 ;
        RECT 445.950 334.950 448.050 337.050 ;
        RECT 448.950 334.950 451.050 337.050 ;
        RECT 433.950 325.950 436.050 328.050 ;
        RECT 427.950 322.950 430.050 325.050 ;
        RECT 430.950 322.950 433.050 325.050 ;
        RECT 418.950 316.950 421.050 319.050 ;
        RECT 427.950 316.950 430.050 319.050 ;
        RECT 412.950 313.950 415.050 316.050 ;
        RECT 418.950 313.950 421.050 316.050 ;
        RECT 419.400 313.050 420.450 313.950 ;
        RECT 412.950 310.950 415.050 313.050 ;
        RECT 416.250 311.250 417.750 312.150 ;
        RECT 418.950 310.950 421.050 313.050 ;
        RECT 422.250 311.250 423.750 312.150 ;
        RECT 424.950 310.950 427.050 313.050 ;
        RECT 428.400 310.050 429.450 316.950 ;
        RECT 434.400 315.450 435.450 325.950 ;
        RECT 431.400 314.400 435.450 315.450 ;
        RECT 431.400 313.050 432.450 314.400 ;
        RECT 436.950 313.950 439.050 316.050 ;
        RECT 437.400 313.050 438.450 313.950 ;
        RECT 443.400 313.050 444.450 334.950 ;
        RECT 446.400 325.050 447.450 334.950 ;
        RECT 445.950 322.950 448.050 325.050 ;
        RECT 448.950 313.950 451.050 316.050 ;
        RECT 430.950 310.950 433.050 313.050 ;
        RECT 434.250 311.250 435.750 312.150 ;
        RECT 436.950 310.950 439.050 313.050 ;
        RECT 440.250 311.250 441.750 312.150 ;
        RECT 442.950 310.950 445.050 313.050 ;
        RECT 412.950 308.850 414.750 309.750 ;
        RECT 415.950 307.950 418.050 310.050 ;
        RECT 419.250 308.850 420.750 309.750 ;
        RECT 421.950 307.950 424.050 310.050 ;
        RECT 425.250 308.850 427.050 309.750 ;
        RECT 427.950 307.950 430.050 310.050 ;
        RECT 430.950 308.850 432.750 309.750 ;
        RECT 433.950 307.950 436.050 310.050 ;
        RECT 437.250 308.850 438.750 309.750 ;
        RECT 439.950 307.950 442.050 310.050 ;
        RECT 443.250 308.850 445.050 309.750 ;
        RECT 415.950 304.950 418.050 307.050 ;
        RECT 416.400 295.050 417.450 304.950 ;
        RECT 422.400 304.050 423.450 307.950 ;
        RECT 434.400 307.050 435.450 307.950 ;
        RECT 427.950 304.950 430.050 307.050 ;
        RECT 433.950 304.950 436.050 307.050 ;
        RECT 421.950 301.950 424.050 304.050 ;
        RECT 418.950 298.950 421.050 301.050 ;
        RECT 412.950 292.950 415.050 295.050 ;
        RECT 415.950 292.950 418.050 295.050 ;
        RECT 413.400 262.050 414.450 292.950 ;
        RECT 415.950 283.950 418.050 286.050 ;
        RECT 416.400 274.050 417.450 283.950 ;
        RECT 419.400 277.050 420.450 298.950 ;
        RECT 422.400 298.050 423.450 301.950 ;
        RECT 421.950 295.950 424.050 298.050 ;
        RECT 424.950 277.950 427.050 280.050 ;
        RECT 418.950 274.950 421.050 277.050 ;
        RECT 415.950 271.950 418.050 274.050 ;
        RECT 419.400 273.450 420.450 274.950 ;
        RECT 425.400 274.050 426.450 277.950 ;
        RECT 428.400 277.050 429.450 304.950 ;
        RECT 440.400 298.050 441.450 307.950 ;
        RECT 445.950 298.950 448.050 301.050 ;
        RECT 439.950 295.950 442.050 298.050 ;
        RECT 446.400 277.050 447.450 298.950 ;
        RECT 449.400 286.050 450.450 313.950 ;
        RECT 448.950 283.950 451.050 286.050 ;
        RECT 452.400 283.050 453.450 340.950 ;
        RECT 454.950 337.950 457.050 340.050 ;
        RECT 458.250 338.250 459.750 339.150 ;
        RECT 460.950 337.950 463.050 340.050 ;
        RECT 455.400 316.050 456.450 337.950 ;
        RECT 457.950 334.950 460.050 337.050 ;
        RECT 458.400 331.050 459.450 334.950 ;
        RECT 457.950 328.950 460.050 331.050 ;
        RECT 461.400 328.050 462.450 337.950 ;
        RECT 466.950 331.950 469.050 334.050 ;
        RECT 460.950 325.950 463.050 328.050 ;
        RECT 463.950 325.950 466.050 328.050 ;
        RECT 454.950 315.450 457.050 316.050 ;
        RECT 457.950 315.450 460.050 316.050 ;
        RECT 454.950 314.400 460.050 315.450 ;
        RECT 454.950 313.950 457.050 314.400 ;
        RECT 457.950 313.950 460.050 314.400 ;
        RECT 460.950 313.950 463.050 316.050 ;
        RECT 454.950 311.250 457.050 312.150 ;
        RECT 457.950 311.850 460.050 312.750 ;
        RECT 454.950 307.950 457.050 310.050 ;
        RECT 457.950 307.950 460.050 310.050 ;
        RECT 448.950 280.950 451.050 283.050 ;
        RECT 451.950 280.950 454.050 283.050 ;
        RECT 427.950 274.950 430.050 277.050 ;
        RECT 430.950 276.450 433.050 277.050 ;
        RECT 430.950 275.400 438.450 276.450 ;
        RECT 430.950 274.950 433.050 275.400 ;
        RECT 437.400 274.050 438.450 275.400 ;
        RECT 442.950 275.250 445.050 276.150 ;
        RECT 445.950 274.950 448.050 277.050 ;
        RECT 419.400 272.400 423.450 273.450 ;
        RECT 422.400 271.050 423.450 272.400 ;
        RECT 424.950 271.950 427.050 274.050 ;
        RECT 427.950 272.250 430.050 273.150 ;
        RECT 430.950 271.950 433.050 274.050 ;
        RECT 436.950 271.950 439.050 274.050 ;
        RECT 440.250 272.250 441.750 273.150 ;
        RECT 442.950 271.950 445.050 274.050 ;
        RECT 446.250 272.250 448.050 273.150 ;
        RECT 415.950 268.950 418.050 271.050 ;
        RECT 418.950 269.250 420.750 270.150 ;
        RECT 421.950 268.950 424.050 271.050 ;
        RECT 425.250 269.250 426.750 270.150 ;
        RECT 427.950 268.950 430.050 271.050 ;
        RECT 409.950 259.950 412.050 262.050 ;
        RECT 412.950 259.950 415.050 262.050 ;
        RECT 406.950 253.950 409.050 256.050 ;
        RECT 410.400 250.050 411.450 259.950 ;
        RECT 416.400 253.050 417.450 268.950 ;
        RECT 428.400 268.050 429.450 268.950 ;
        RECT 418.950 265.950 421.050 268.050 ;
        RECT 422.250 266.850 423.750 267.750 ;
        RECT 424.950 265.950 427.050 268.050 ;
        RECT 427.950 265.950 430.050 268.050 ;
        RECT 425.400 259.050 426.450 265.950 ;
        RECT 431.400 259.050 432.450 271.950 ;
        RECT 436.950 269.850 438.750 270.750 ;
        RECT 439.950 268.950 442.050 271.050 ;
        RECT 424.950 256.950 427.050 259.050 ;
        RECT 430.950 256.950 433.050 259.050 ;
        RECT 436.950 256.950 439.050 259.050 ;
        RECT 412.950 250.950 415.050 253.050 ;
        RECT 415.950 250.950 418.050 253.050 ;
        RECT 409.950 247.950 412.050 250.050 ;
        RECT 406.950 244.950 409.050 247.050 ;
        RECT 391.950 238.950 394.050 241.050 ;
        RECT 395.250 239.250 396.750 240.150 ;
        RECT 397.950 238.950 400.050 241.050 ;
        RECT 401.250 239.250 402.750 240.150 ;
        RECT 403.950 238.950 406.050 241.050 ;
        RECT 391.950 236.850 393.750 237.750 ;
        RECT 394.950 235.950 397.050 238.050 ;
        RECT 398.250 236.850 399.750 237.750 ;
        RECT 400.950 235.950 403.050 238.050 ;
        RECT 404.250 236.850 406.050 237.750 ;
        RECT 389.400 233.400 393.450 234.450 ;
        RECT 392.400 232.050 393.450 233.400 ;
        RECT 397.950 232.950 400.050 235.050 ;
        RECT 388.950 229.950 391.050 232.050 ;
        RECT 391.950 229.950 394.050 232.050 ;
        RECT 389.400 217.050 390.450 229.950 ;
        RECT 394.950 226.950 397.050 229.050 ;
        RECT 388.950 214.950 391.050 217.050 ;
        RECT 385.950 205.950 388.050 208.050 ;
        RECT 391.950 205.950 394.050 208.050 ;
        RECT 379.950 202.950 382.050 205.050 ;
        RECT 376.950 197.250 378.750 198.150 ;
        RECT 379.950 196.950 382.050 199.050 ;
        RECT 383.250 197.250 384.750 198.150 ;
        RECT 385.950 196.950 388.050 199.050 ;
        RECT 389.250 197.250 391.050 198.150 ;
        RECT 373.950 193.950 376.050 196.050 ;
        RECT 376.950 193.950 379.050 196.050 ;
        RECT 380.250 194.850 381.750 195.750 ;
        RECT 382.950 193.950 385.050 196.050 ;
        RECT 386.250 194.850 387.750 195.750 ;
        RECT 388.950 193.950 391.050 196.050 ;
        RECT 367.950 190.950 370.050 193.050 ;
        RECT 370.950 190.950 373.050 193.050 ;
        RECT 355.950 187.950 358.050 190.050 ;
        RECT 364.950 187.950 367.050 190.050 ;
        RECT 370.950 187.950 373.050 190.050 ;
        RECT 355.950 175.950 358.050 178.050 ;
        RECT 356.400 157.050 357.450 175.950 ;
        RECT 367.950 166.950 370.050 169.050 ;
        RECT 371.400 168.450 372.450 187.950 ;
        RECT 377.400 187.050 378.450 193.950 ;
        RECT 383.400 193.050 384.450 193.950 ;
        RECT 382.950 190.950 385.050 193.050 ;
        RECT 392.400 187.050 393.450 205.950 ;
        RECT 376.950 184.950 379.050 187.050 ;
        RECT 391.950 184.950 394.050 187.050 ;
        RECT 379.950 169.950 382.050 172.050 ;
        RECT 380.400 169.050 381.450 169.950 ;
        RECT 373.950 168.450 376.050 169.050 ;
        RECT 371.400 167.400 376.050 168.450 ;
        RECT 368.400 166.050 369.450 166.950 ;
        RECT 358.950 164.250 360.750 165.150 ;
        RECT 361.950 163.950 364.050 166.050 ;
        RECT 367.950 163.950 370.050 166.050 ;
        RECT 358.950 160.950 361.050 163.050 ;
        RECT 362.250 161.850 363.750 162.750 ;
        RECT 364.950 160.950 367.050 163.050 ;
        RECT 368.250 161.850 370.050 162.750 ;
        RECT 371.400 162.450 372.450 167.400 ;
        RECT 373.950 166.950 376.050 167.400 ;
        RECT 377.250 167.250 378.750 168.150 ;
        RECT 379.950 166.950 382.050 169.050 ;
        RECT 385.950 168.450 388.050 169.050 ;
        RECT 383.250 167.250 384.750 168.150 ;
        RECT 385.950 167.400 390.450 168.450 ;
        RECT 385.950 166.950 388.050 167.400 ;
        RECT 373.950 164.850 375.750 165.750 ;
        RECT 376.950 163.950 379.050 166.050 ;
        RECT 380.250 164.850 381.750 165.750 ;
        RECT 382.950 163.950 385.050 166.050 ;
        RECT 386.250 164.850 388.050 165.750 ;
        RECT 371.400 161.400 375.450 162.450 ;
        RECT 361.950 157.950 364.050 160.050 ;
        RECT 364.950 158.850 367.050 159.750 ;
        RECT 367.950 157.950 370.050 160.050 ;
        RECT 355.950 154.950 358.050 157.050 ;
        RECT 358.950 133.950 361.050 136.050 ;
        RECT 359.400 133.050 360.450 133.950 ;
        RECT 358.950 130.950 361.050 133.050 ;
        RECT 352.950 127.950 355.050 130.050 ;
        RECT 355.950 128.250 358.050 129.150 ;
        RECT 358.950 127.950 361.050 130.050 ;
        RECT 334.950 124.950 337.050 127.050 ;
        RECT 338.250 125.250 339.750 126.150 ;
        RECT 340.950 124.950 343.050 127.050 ;
        RECT 344.250 125.250 346.050 126.150 ;
        RECT 346.950 125.250 348.750 126.150 ;
        RECT 349.950 124.950 352.050 127.050 ;
        RECT 353.250 125.250 354.750 126.150 ;
        RECT 355.950 124.950 358.050 127.050 ;
        RECT 334.950 121.950 337.050 124.050 ;
        RECT 337.950 121.950 340.050 124.050 ;
        RECT 341.250 122.850 342.750 123.750 ;
        RECT 343.950 121.950 346.050 124.050 ;
        RECT 346.950 121.950 349.050 124.050 ;
        RECT 350.250 122.850 351.750 123.750 ;
        RECT 352.950 121.950 355.050 124.050 ;
        RECT 355.950 121.950 358.050 124.050 ;
        RECT 329.400 119.400 333.450 120.450 ;
        RECT 325.950 100.950 328.050 103.050 ;
        RECT 329.400 100.050 330.450 119.400 ;
        RECT 332.400 118.050 333.450 119.400 ;
        RECT 331.950 115.950 334.050 118.050 ;
        RECT 335.400 117.450 336.450 121.950 ;
        RECT 338.400 121.050 339.450 121.950 ;
        RECT 337.950 118.950 340.050 121.050 ;
        RECT 335.400 116.400 339.450 117.450 ;
        RECT 334.950 106.950 337.050 109.050 ;
        RECT 331.950 100.950 334.050 103.050 ;
        RECT 328.950 97.950 331.050 100.050 ;
        RECT 332.400 97.050 333.450 100.950 ;
        RECT 335.400 97.050 336.450 106.950 ;
        RECT 338.400 97.050 339.450 116.400 ;
        RECT 344.400 112.050 345.450 121.950 ;
        RECT 343.950 109.950 346.050 112.050 ;
        RECT 344.400 97.050 345.450 109.950 ;
        RECT 322.950 96.450 325.050 97.050 ;
        RECT 325.950 96.450 328.050 97.050 ;
        RECT 322.950 95.400 328.050 96.450 ;
        RECT 329.250 95.850 330.750 96.750 ;
        RECT 322.950 94.950 325.050 95.400 ;
        RECT 325.950 94.950 328.050 95.400 ;
        RECT 331.950 94.950 334.050 97.050 ;
        RECT 334.950 94.950 337.050 97.050 ;
        RECT 337.950 94.950 340.050 97.050 ;
        RECT 343.950 94.950 346.050 97.050 ;
        RECT 323.400 82.050 324.450 94.950 ;
        RECT 325.950 92.850 328.050 93.750 ;
        RECT 331.950 92.850 334.050 93.750 ;
        RECT 334.950 92.850 337.050 93.750 ;
        RECT 340.950 92.250 343.050 93.150 ;
        RECT 343.950 92.850 346.050 93.750 ;
        RECT 340.950 88.950 343.050 91.050 ;
        RECT 343.950 88.950 346.050 91.050 ;
        RECT 322.950 79.950 325.050 82.050 ;
        RECT 325.950 79.950 328.050 82.050 ;
        RECT 319.950 58.950 322.050 61.050 ;
        RECT 310.950 55.950 313.050 58.050 ;
        RECT 322.950 56.250 325.050 57.150 ;
        RECT 307.950 52.950 310.050 55.050 ;
        RECT 307.950 49.950 310.050 52.050 ;
        RECT 311.400 51.450 312.450 55.950 ;
        RECT 313.950 53.250 315.750 54.150 ;
        RECT 316.950 52.950 319.050 55.050 ;
        RECT 320.250 53.250 321.750 54.150 ;
        RECT 322.950 52.950 325.050 55.050 ;
        RECT 326.400 52.050 327.450 79.950 ;
        RECT 328.950 58.950 331.050 61.050 ;
        RECT 313.950 51.450 316.050 52.050 ;
        RECT 311.400 50.400 316.050 51.450 ;
        RECT 317.250 50.850 318.750 51.750 ;
        RECT 313.950 49.950 316.050 50.400 ;
        RECT 319.950 49.950 322.050 52.050 ;
        RECT 325.950 49.950 328.050 52.050 ;
        RECT 329.400 51.450 330.450 58.950 ;
        RECT 331.950 53.250 334.050 54.150 ;
        RECT 337.950 53.250 340.050 54.150 ;
        RECT 331.950 51.450 334.050 52.050 ;
        RECT 329.400 50.400 334.050 51.450 ;
        RECT 331.950 49.950 334.050 50.400 ;
        RECT 335.250 50.250 336.750 51.150 ;
        RECT 337.950 49.950 340.050 52.050 ;
        RECT 308.400 40.050 309.450 49.950 ;
        RECT 334.950 48.450 337.050 49.050 ;
        RECT 337.950 48.450 340.050 49.050 ;
        RECT 334.950 47.400 340.050 48.450 ;
        RECT 334.950 46.950 337.050 47.400 ;
        RECT 337.950 46.950 340.050 47.400 ;
        RECT 334.950 43.950 337.050 46.050 ;
        RECT 307.950 37.950 310.050 40.050 ;
        RECT 322.950 34.950 325.050 37.050 ;
        RECT 313.950 25.950 316.050 28.050 ;
        RECT 304.950 22.950 307.050 25.050 ;
        RECT 308.250 23.250 309.750 24.150 ;
        RECT 310.950 22.950 313.050 25.050 ;
        RECT 314.400 22.050 315.450 25.950 ;
        RECT 316.950 22.950 319.050 25.050 ;
        RECT 319.950 22.950 322.050 25.050 ;
        RECT 304.950 20.850 306.750 21.750 ;
        RECT 307.950 19.950 310.050 22.050 ;
        RECT 311.250 20.850 312.750 21.750 ;
        RECT 313.950 19.950 316.050 22.050 ;
        RECT 313.950 17.850 316.050 18.750 ;
        RECT 301.950 13.950 304.050 16.050 ;
        RECT 317.400 13.050 318.450 22.950 ;
        RECT 320.400 16.050 321.450 22.950 ;
        RECT 323.400 22.050 324.450 34.950 ;
        RECT 328.950 25.950 331.050 28.050 ;
        RECT 329.400 25.050 330.450 25.950 ;
        RECT 335.400 25.050 336.450 43.950 ;
        RECT 337.950 37.950 340.050 40.050 ;
        RECT 325.950 22.950 328.050 25.050 ;
        RECT 328.950 22.950 331.050 25.050 ;
        RECT 332.250 23.250 333.750 24.150 ;
        RECT 334.950 22.950 337.050 25.050 ;
        RECT 326.400 22.050 327.450 22.950 ;
        RECT 322.950 19.950 325.050 22.050 ;
        RECT 325.950 19.950 328.050 22.050 ;
        RECT 329.250 20.850 330.750 21.750 ;
        RECT 331.950 19.950 334.050 22.050 ;
        RECT 335.250 20.850 337.050 21.750 ;
        RECT 325.950 17.850 328.050 18.750 ;
        RECT 319.950 13.950 322.050 16.050 ;
        RECT 283.950 10.950 286.050 13.050 ;
        RECT 316.950 10.950 319.050 13.050 ;
        RECT 227.100 7.800 229.200 9.900 ;
        RECT 338.400 7.050 339.450 37.950 ;
        RECT 341.400 28.050 342.450 88.950 ;
        RECT 344.400 43.050 345.450 88.950 ;
        RECT 347.400 58.050 348.450 121.950 ;
        RECT 356.400 106.050 357.450 121.950 ;
        RECT 359.400 106.050 360.450 127.950 ;
        RECT 362.400 115.050 363.450 157.950 ;
        RECT 364.950 151.950 367.050 154.050 ;
        RECT 365.400 130.050 366.450 151.950 ;
        RECT 364.950 127.950 367.050 130.050 ;
        RECT 364.950 124.950 367.050 127.050 ;
        RECT 365.400 118.050 366.450 124.950 ;
        RECT 364.950 115.950 367.050 118.050 ;
        RECT 361.950 112.950 364.050 115.050 ;
        RECT 355.950 103.950 358.050 106.050 ;
        RECT 358.950 103.950 361.050 106.050 ;
        RECT 364.950 103.950 367.050 106.050 ;
        RECT 352.950 97.950 355.050 100.050 ;
        RECT 361.950 97.950 364.050 100.050 ;
        RECT 349.950 95.250 352.050 96.150 ;
        RECT 352.950 95.850 355.050 96.750 ;
        RECT 355.950 95.250 357.750 96.150 ;
        RECT 358.950 94.950 361.050 97.050 ;
        RECT 349.950 91.950 352.050 94.050 ;
        RECT 355.950 91.950 358.050 94.050 ;
        RECT 359.250 92.850 361.050 93.750 ;
        RECT 350.400 91.050 351.450 91.950 ;
        RECT 349.950 88.950 352.050 91.050 ;
        RECT 356.400 70.050 357.450 91.950 ;
        RECT 358.950 82.950 361.050 85.050 ;
        RECT 355.950 67.950 358.050 70.050 ;
        RECT 355.950 58.950 358.050 61.050 ;
        RECT 346.950 55.950 349.050 58.050 ;
        RECT 346.950 53.250 349.050 54.150 ;
        RECT 352.950 53.250 355.050 54.150 ;
        RECT 356.400 52.050 357.450 58.950 ;
        RECT 346.950 49.950 349.050 52.050 ;
        RECT 350.250 50.250 351.750 51.150 ;
        RECT 352.950 49.950 355.050 52.050 ;
        RECT 355.950 49.950 358.050 52.050 ;
        RECT 347.400 49.050 348.450 49.950 ;
        RECT 353.400 49.050 354.450 49.950 ;
        RECT 346.950 46.950 349.050 49.050 ;
        RECT 349.950 46.950 352.050 49.050 ;
        RECT 352.950 46.950 355.050 49.050 ;
        RECT 343.950 40.950 346.050 43.050 ;
        RECT 350.400 40.050 351.450 46.950 ;
        RECT 349.950 37.950 352.050 40.050 ;
        RECT 340.950 25.950 343.050 28.050 ;
        RECT 352.950 25.950 355.050 28.050 ;
        RECT 340.950 19.950 343.050 22.050 ;
        RECT 343.950 20.250 345.750 21.150 ;
        RECT 346.950 19.950 349.050 22.050 ;
        RECT 350.250 20.250 352.050 21.150 ;
        RECT 341.400 18.450 342.450 19.950 ;
        RECT 343.950 18.450 346.050 19.050 ;
        RECT 341.400 17.400 346.050 18.450 ;
        RECT 347.250 17.850 348.750 18.750 ;
        RECT 349.950 18.450 352.050 19.050 ;
        RECT 353.400 18.450 354.450 25.950 ;
        RECT 359.400 25.050 360.450 82.950 ;
        RECT 362.400 58.050 363.450 97.950 ;
        RECT 365.400 70.050 366.450 103.950 ;
        RECT 368.400 76.050 369.450 157.950 ;
        RECT 374.400 130.050 375.450 161.400 ;
        RECT 377.400 145.050 378.450 163.950 ;
        RECT 383.400 154.050 384.450 163.950 ;
        RECT 389.400 163.050 390.450 167.400 ;
        RECT 391.950 163.950 394.050 166.050 ;
        RECT 388.950 160.950 391.050 163.050 ;
        RECT 382.950 151.950 385.050 154.050 ;
        RECT 376.950 142.950 379.050 145.050 ;
        RECT 379.950 142.950 382.050 145.050 ;
        RECT 380.400 139.050 381.450 142.950 ;
        RECT 379.950 136.950 382.050 139.050 ;
        RECT 383.400 133.050 384.450 151.950 ;
        RECT 392.400 133.050 393.450 163.950 ;
        RECT 395.400 160.050 396.450 226.950 ;
        RECT 398.400 199.050 399.450 232.950 ;
        RECT 401.400 232.050 402.450 235.950 ;
        RECT 407.400 234.450 408.450 244.950 ;
        RECT 413.400 238.050 414.450 250.950 ;
        RECT 427.950 247.950 430.050 250.050 ;
        RECT 418.950 241.950 421.050 244.050 ;
        RECT 421.950 241.950 424.050 244.050 ;
        RECT 409.950 236.250 411.750 237.150 ;
        RECT 412.950 235.950 415.050 238.050 ;
        RECT 416.250 236.250 418.050 237.150 ;
        RECT 409.950 234.450 412.050 235.050 ;
        RECT 407.400 233.400 412.050 234.450 ;
        RECT 413.250 233.850 414.750 234.750 ;
        RECT 400.950 229.950 403.050 232.050 ;
        RECT 407.400 220.050 408.450 233.400 ;
        RECT 409.950 232.950 412.050 233.400 ;
        RECT 415.950 232.950 418.050 235.050 ;
        RECT 412.950 229.950 415.050 232.050 ;
        RECT 409.950 226.950 412.050 229.050 ;
        RECT 406.950 217.950 409.050 220.050 ;
        RECT 397.950 196.950 400.050 199.050 ;
        RECT 400.950 197.250 403.050 198.150 ;
        RECT 406.950 197.250 409.050 198.150 ;
        RECT 398.400 193.050 399.450 196.950 ;
        RECT 400.950 193.950 403.050 196.050 ;
        RECT 404.250 194.250 405.750 195.150 ;
        RECT 406.950 193.950 409.050 196.050 ;
        RECT 397.950 190.950 400.050 193.050 ;
        RECT 401.400 189.450 402.450 193.950 ;
        RECT 403.950 190.950 406.050 193.050 ;
        RECT 401.400 188.400 405.450 189.450 ;
        RECT 404.400 184.050 405.450 188.400 ;
        RECT 407.400 187.050 408.450 193.950 ;
        RECT 410.400 190.050 411.450 226.950 ;
        RECT 413.400 202.050 414.450 229.950 ;
        RECT 416.400 229.050 417.450 232.950 ;
        RECT 415.950 226.950 418.050 229.050 ;
        RECT 419.400 220.050 420.450 241.950 ;
        RECT 418.950 217.950 421.050 220.050 ;
        RECT 422.400 208.050 423.450 241.950 ;
        RECT 424.950 238.950 427.050 241.050 ;
        RECT 425.400 238.050 426.450 238.950 ;
        RECT 424.950 235.950 427.050 238.050 ;
        RECT 428.400 235.050 429.450 247.950 ;
        RECT 430.950 241.950 433.050 244.050 ;
        RECT 431.400 238.050 432.450 241.950 ;
        RECT 430.950 235.950 433.050 238.050 ;
        RECT 434.250 236.250 436.050 237.150 ;
        RECT 424.950 233.850 426.750 234.750 ;
        RECT 427.950 232.950 430.050 235.050 ;
        RECT 431.250 233.850 432.750 234.750 ;
        RECT 433.950 232.950 436.050 235.050 ;
        RECT 434.400 232.050 435.450 232.950 ;
        RECT 427.950 230.850 430.050 231.750 ;
        RECT 433.950 229.950 436.050 232.050 ;
        RECT 427.950 226.950 430.050 229.050 ;
        RECT 433.950 226.950 436.050 229.050 ;
        RECT 424.950 214.950 427.050 217.050 ;
        RECT 421.950 205.950 424.050 208.050 ;
        RECT 425.400 205.050 426.450 214.950 ;
        RECT 428.400 208.050 429.450 226.950 ;
        RECT 430.950 223.950 433.050 226.050 ;
        RECT 431.400 217.050 432.450 223.950 ;
        RECT 430.950 214.950 433.050 217.050 ;
        RECT 427.950 205.950 430.050 208.050 ;
        RECT 415.950 202.950 418.050 205.050 ;
        RECT 424.950 202.950 427.050 205.050 ;
        RECT 412.950 199.950 415.050 202.050 ;
        RECT 413.400 199.050 414.450 199.950 ;
        RECT 412.950 196.950 415.050 199.050 ;
        RECT 416.400 196.050 417.450 202.950 ;
        RECT 418.950 197.250 421.050 198.150 ;
        RECT 424.950 197.250 427.050 198.150 ;
        RECT 430.950 197.250 433.050 198.150 ;
        RECT 412.950 194.850 415.050 195.750 ;
        RECT 415.950 193.950 418.050 196.050 ;
        RECT 418.950 193.950 421.050 196.050 ;
        RECT 422.250 194.250 424.050 195.150 ;
        RECT 424.950 193.950 427.050 196.050 ;
        RECT 428.250 194.250 429.750 195.150 ;
        RECT 430.950 193.950 433.050 196.050 ;
        RECT 409.950 187.950 412.050 190.050 ;
        RECT 419.400 187.050 420.450 193.950 ;
        RECT 421.950 190.950 424.050 193.050 ;
        RECT 406.950 184.950 409.050 187.050 ;
        RECT 418.950 184.950 421.050 187.050 ;
        RECT 422.400 184.050 423.450 190.950 ;
        RECT 425.400 190.050 426.450 193.950 ;
        RECT 427.950 190.950 430.050 193.050 ;
        RECT 424.950 187.950 427.050 190.050 ;
        RECT 403.950 181.950 406.050 184.050 ;
        RECT 421.950 181.950 424.050 184.050 ;
        RECT 425.400 183.450 426.450 187.950 ;
        RECT 428.400 187.050 429.450 190.950 ;
        RECT 427.950 184.950 430.050 187.050 ;
        RECT 425.400 182.400 429.450 183.450 ;
        RECT 400.950 175.950 403.050 178.050 ;
        RECT 401.400 166.050 402.450 175.950 ;
        RECT 404.400 172.050 405.450 181.950 ;
        RECT 415.950 175.950 418.050 178.050 ;
        RECT 418.950 175.950 421.050 178.050 ;
        RECT 409.950 172.950 412.050 175.050 ;
        RECT 403.950 169.950 406.050 172.050 ;
        RECT 406.950 169.950 409.050 172.050 ;
        RECT 407.400 166.050 408.450 169.950 ;
        RECT 397.950 164.250 399.750 165.150 ;
        RECT 400.950 163.950 403.050 166.050 ;
        RECT 404.250 164.250 406.050 165.150 ;
        RECT 406.950 163.950 409.050 166.050 ;
        RECT 397.950 160.950 400.050 163.050 ;
        RECT 401.250 161.850 402.750 162.750 ;
        RECT 403.950 160.950 406.050 163.050 ;
        RECT 406.950 160.950 409.050 163.050 ;
        RECT 394.950 157.950 397.050 160.050 ;
        RECT 398.400 154.050 399.450 160.950 ;
        RECT 404.400 159.450 405.450 160.950 ;
        RECT 401.400 158.400 405.450 159.450 ;
        RECT 397.950 151.950 400.050 154.050 ;
        RECT 394.950 136.950 397.050 139.050 ;
        RECT 382.950 130.950 385.050 133.050 ;
        RECT 385.950 131.250 388.050 132.150 ;
        RECT 391.950 130.950 394.050 133.050 ;
        RECT 370.950 128.250 373.050 129.150 ;
        RECT 373.950 127.950 376.050 130.050 ;
        RECT 382.950 128.250 384.750 129.150 ;
        RECT 385.950 127.950 388.050 130.050 ;
        RECT 391.950 129.450 394.050 130.050 ;
        RECT 395.400 129.450 396.450 136.950 ;
        RECT 397.950 130.950 400.050 133.050 ;
        RECT 389.250 128.250 390.750 129.150 ;
        RECT 391.950 128.400 396.450 129.450 ;
        RECT 391.950 127.950 394.050 128.400 ;
        RECT 370.950 124.950 373.050 127.050 ;
        RECT 374.250 125.250 375.750 126.150 ;
        RECT 376.950 124.950 379.050 127.050 ;
        RECT 380.250 125.250 382.050 126.150 ;
        RECT 382.950 124.950 385.050 127.050 ;
        RECT 388.950 124.950 391.050 127.050 ;
        RECT 392.250 125.850 394.050 126.750 ;
        RECT 394.950 124.950 397.050 127.050 ;
        RECT 371.400 124.050 372.450 124.950 ;
        RECT 383.400 124.050 384.450 124.950 ;
        RECT 370.950 121.950 373.050 124.050 ;
        RECT 373.950 121.950 376.050 124.050 ;
        RECT 377.250 122.850 378.750 123.750 ;
        RECT 379.950 121.950 382.050 124.050 ;
        RECT 382.950 121.950 385.050 124.050 ;
        RECT 371.400 91.050 372.450 121.950 ;
        RECT 374.400 121.050 375.450 121.950 ;
        RECT 373.950 118.950 376.050 121.050 ;
        RECT 376.950 118.950 379.050 121.050 ;
        RECT 377.400 94.050 378.450 118.950 ;
        RECT 380.400 112.050 381.450 121.950 ;
        RECT 389.400 121.050 390.450 124.950 ;
        RECT 388.950 118.950 391.050 121.050 ;
        RECT 379.950 109.950 382.050 112.050 ;
        RECT 382.950 97.950 385.050 100.050 ;
        RECT 383.400 94.050 384.450 97.950 ;
        RECT 395.400 97.050 396.450 124.950 ;
        RECT 398.400 123.450 399.450 130.950 ;
        RECT 401.400 130.050 402.450 158.400 ;
        RECT 407.400 154.050 408.450 160.950 ;
        RECT 410.400 160.050 411.450 172.950 ;
        RECT 412.950 166.950 415.050 169.050 ;
        RECT 413.400 163.050 414.450 166.950 ;
        RECT 416.400 166.050 417.450 175.950 ;
        RECT 419.400 169.050 420.450 175.950 ;
        RECT 424.950 172.950 427.050 175.050 ;
        RECT 425.400 172.050 426.450 172.950 ;
        RECT 424.950 169.950 427.050 172.050 ;
        RECT 418.950 166.950 421.050 169.050 ;
        RECT 422.250 167.250 423.750 168.150 ;
        RECT 424.950 166.950 427.050 169.050 ;
        RECT 415.950 163.950 418.050 166.050 ;
        RECT 419.250 164.850 420.750 165.750 ;
        RECT 421.950 163.950 424.050 166.050 ;
        RECT 425.250 164.850 427.050 165.750 ;
        RECT 412.950 160.950 415.050 163.050 ;
        RECT 415.950 161.850 418.050 162.750 ;
        RECT 409.950 157.950 412.050 160.050 ;
        RECT 406.950 151.950 409.050 154.050 ;
        RECT 413.400 139.050 414.450 160.950 ;
        RECT 422.400 142.050 423.450 163.950 ;
        RECT 428.400 162.450 429.450 182.400 ;
        RECT 425.400 161.400 429.450 162.450 ;
        RECT 431.400 162.450 432.450 193.950 ;
        RECT 434.400 178.050 435.450 226.950 ;
        RECT 437.400 199.050 438.450 256.950 ;
        RECT 440.400 253.050 441.450 268.950 ;
        RECT 443.400 264.450 444.450 271.950 ;
        RECT 445.950 268.950 448.050 271.050 ;
        RECT 446.400 268.050 447.450 268.950 ;
        RECT 445.950 265.950 448.050 268.050 ;
        RECT 443.400 263.400 447.450 264.450 ;
        RECT 446.400 256.050 447.450 263.400 ;
        RECT 445.950 253.950 448.050 256.050 ;
        RECT 449.400 253.050 450.450 280.950 ;
        RECT 455.400 279.450 456.450 307.950 ;
        RECT 458.400 292.050 459.450 307.950 ;
        RECT 457.950 289.950 460.050 292.050 ;
        RECT 461.400 280.050 462.450 313.950 ;
        RECT 455.400 278.400 459.450 279.450 ;
        RECT 454.950 274.950 457.050 277.050 ;
        RECT 458.400 276.450 459.450 278.400 ;
        RECT 460.950 277.950 463.050 280.050 ;
        RECT 458.400 275.400 462.450 276.450 ;
        RECT 455.400 274.050 456.450 274.950 ;
        RECT 461.400 274.050 462.450 275.400 ;
        RECT 451.950 271.950 454.050 274.050 ;
        RECT 454.950 271.950 457.050 274.050 ;
        RECT 458.250 272.250 459.750 273.150 ;
        RECT 460.950 271.950 463.050 274.050 ;
        RECT 452.400 268.050 453.450 271.950 ;
        RECT 454.950 269.850 456.750 270.750 ;
        RECT 457.950 268.950 460.050 271.050 ;
        RECT 461.250 269.850 463.050 270.750 ;
        RECT 458.400 268.050 459.450 268.950 ;
        RECT 464.400 268.050 465.450 325.950 ;
        RECT 467.400 316.050 468.450 331.950 ;
        RECT 470.400 316.050 471.450 382.950 ;
        RECT 476.400 379.050 477.450 385.950 ;
        RECT 485.400 385.050 486.450 403.950 ;
        RECT 494.400 403.050 495.450 412.950 ;
        RECT 487.950 400.950 490.050 403.050 ;
        RECT 493.950 400.950 496.050 403.050 ;
        RECT 478.950 382.950 481.050 385.050 ;
        RECT 482.250 383.850 483.750 384.750 ;
        RECT 484.950 382.950 487.050 385.050 ;
        RECT 478.950 380.850 481.050 381.750 ;
        RECT 484.950 380.850 487.050 381.750 ;
        RECT 475.950 376.950 478.050 379.050 ;
        RECT 481.950 376.950 484.050 379.050 ;
        RECT 475.950 370.950 478.050 373.050 ;
        RECT 476.400 343.050 477.450 370.950 ;
        RECT 472.950 341.250 474.750 342.150 ;
        RECT 475.950 340.950 478.050 343.050 ;
        RECT 472.950 337.950 475.050 340.050 ;
        RECT 476.250 338.850 478.050 339.750 ;
        RECT 473.400 325.050 474.450 337.950 ;
        RECT 475.950 328.950 478.050 331.050 ;
        RECT 472.950 322.950 475.050 325.050 ;
        RECT 476.400 322.050 477.450 328.950 ;
        RECT 475.950 319.950 478.050 322.050 ;
        RECT 466.950 313.950 469.050 316.050 ;
        RECT 469.950 313.950 472.050 316.050 ;
        RECT 466.950 310.950 469.050 313.050 ;
        RECT 470.250 311.250 471.750 312.150 ;
        RECT 472.950 310.950 475.050 313.050 ;
        RECT 466.950 308.850 468.750 309.750 ;
        RECT 469.950 307.950 472.050 310.050 ;
        RECT 473.250 308.850 474.750 309.750 ;
        RECT 475.950 309.450 478.050 310.050 ;
        RECT 475.950 308.400 480.450 309.450 ;
        RECT 475.950 307.950 478.050 308.400 ;
        RECT 466.950 304.950 469.050 307.050 ;
        RECT 467.400 285.450 468.450 304.950 ;
        RECT 470.400 289.050 471.450 307.950 ;
        RECT 475.950 305.850 478.050 306.750 ;
        RECT 479.400 304.050 480.450 308.400 ;
        RECT 478.950 301.950 481.050 304.050 ;
        RECT 482.400 300.450 483.450 376.950 ;
        RECT 488.400 373.050 489.450 400.950 ;
        RECT 490.950 394.950 493.050 397.050 ;
        RECT 491.400 385.050 492.450 394.950 ;
        RECT 493.950 388.950 496.050 391.050 ;
        RECT 490.950 382.950 493.050 385.050 ;
        RECT 490.950 380.850 493.050 381.750 ;
        RECT 494.400 378.450 495.450 388.950 ;
        RECT 497.400 385.050 498.450 454.950 ;
        RECT 499.950 451.950 502.050 454.050 ;
        RECT 505.950 453.450 508.050 454.050 ;
        RECT 503.400 452.400 508.050 453.450 ;
        RECT 500.400 448.050 501.450 451.950 ;
        RECT 503.400 451.050 504.450 452.400 ;
        RECT 505.950 451.950 508.050 452.400 ;
        RECT 508.950 451.950 511.050 454.050 ;
        RECT 511.950 451.950 514.050 454.050 ;
        RECT 515.250 452.250 517.050 453.150 ;
        RECT 509.400 451.050 510.450 451.950 ;
        RECT 502.950 448.950 505.050 451.050 ;
        RECT 505.950 449.850 507.750 450.750 ;
        RECT 508.950 448.950 511.050 451.050 ;
        RECT 512.250 449.850 513.750 450.750 ;
        RECT 514.950 448.950 517.050 451.050 ;
        RECT 499.950 445.950 502.050 448.050 ;
        RECT 502.950 445.950 505.050 448.050 ;
        RECT 505.950 445.950 508.050 448.050 ;
        RECT 508.950 446.850 511.050 447.750 ;
        RECT 503.400 445.050 504.450 445.950 ;
        RECT 502.950 442.950 505.050 445.050 ;
        RECT 499.950 421.950 502.050 424.050 ;
        RECT 500.400 415.050 501.450 421.950 ;
        RECT 499.950 412.950 502.050 415.050 ;
        RECT 502.950 413.250 505.050 414.150 ;
        RECT 499.950 410.250 501.750 411.150 ;
        RECT 502.950 409.950 505.050 412.050 ;
        RECT 499.950 406.950 502.050 409.050 ;
        RECT 506.400 408.450 507.450 445.950 ;
        RECT 511.950 442.950 514.050 445.050 ;
        RECT 508.950 412.950 511.050 415.050 ;
        RECT 508.950 410.850 511.050 411.750 ;
        RECT 512.400 408.450 513.450 442.950 ;
        RECT 518.400 417.450 519.450 457.950 ;
        RECT 521.400 451.050 522.450 466.950 ;
        RECT 524.400 457.050 525.450 493.950 ;
        RECT 527.400 460.050 528.450 500.400 ;
        RECT 536.400 495.450 537.450 520.950 ;
        RECT 538.950 511.950 541.050 514.050 ;
        RECT 533.400 494.400 537.450 495.450 ;
        RECT 529.950 488.250 532.050 489.150 ;
        RECT 529.950 484.950 532.050 487.050 ;
        RECT 530.400 484.050 531.450 484.950 ;
        RECT 529.950 481.950 532.050 484.050 ;
        RECT 526.950 457.950 529.050 460.050 ;
        RECT 533.400 457.050 534.450 494.400 ;
        RECT 535.950 490.950 538.050 493.050 ;
        RECT 536.400 487.050 537.450 490.950 ;
        RECT 535.950 484.950 538.050 487.050 ;
        RECT 539.400 484.050 540.450 511.950 ;
        RECT 542.400 493.050 543.450 529.950 ;
        RECT 560.400 529.050 561.450 538.950 ;
        RECT 562.950 529.950 565.050 532.050 ;
        RECT 547.950 528.450 550.050 529.050 ;
        RECT 545.400 527.400 550.050 528.450 ;
        RECT 545.400 523.050 546.450 527.400 ;
        RECT 547.950 526.950 550.050 527.400 ;
        RECT 551.250 527.250 552.750 528.150 ;
        RECT 553.950 526.950 556.050 529.050 ;
        RECT 557.250 527.250 558.750 528.150 ;
        RECT 559.950 526.950 562.050 529.050 ;
        RECT 563.400 526.050 564.450 529.950 ;
        RECT 566.400 526.050 567.450 550.950 ;
        RECT 568.950 541.950 571.050 544.050 ;
        RECT 547.950 524.850 549.750 525.750 ;
        RECT 550.950 523.950 553.050 526.050 ;
        RECT 554.250 524.850 555.750 525.750 ;
        RECT 556.950 523.950 559.050 526.050 ;
        RECT 560.250 524.850 562.050 525.750 ;
        RECT 562.950 523.950 565.050 526.050 ;
        RECT 565.950 523.950 568.050 526.050 ;
        RECT 544.950 520.950 547.050 523.050 ;
        RECT 551.400 520.050 552.450 523.950 ;
        RECT 553.950 520.950 556.050 523.050 ;
        RECT 544.950 517.950 547.050 520.050 ;
        RECT 550.950 517.950 553.050 520.050 ;
        RECT 541.950 490.950 544.050 493.050 ;
        RECT 541.950 487.950 544.050 490.050 ;
        RECT 542.400 487.050 543.450 487.950 ;
        RECT 541.950 484.950 544.050 487.050 ;
        RECT 538.950 481.950 541.050 484.050 ;
        RECT 541.950 482.850 544.050 483.750 ;
        RECT 523.950 454.950 526.050 457.050 ;
        RECT 526.950 454.950 529.050 457.050 ;
        RECT 529.950 454.950 532.050 457.050 ;
        RECT 532.950 454.950 535.050 457.050 ;
        RECT 520.950 448.950 523.050 451.050 ;
        RECT 524.400 421.050 525.450 454.950 ;
        RECT 527.400 454.050 528.450 454.950 ;
        RECT 526.950 451.950 529.050 454.050 ;
        RECT 530.400 453.450 531.450 454.950 ;
        RECT 532.950 453.450 535.050 454.050 ;
        RECT 530.400 452.400 535.050 453.450 ;
        RECT 532.950 451.950 535.050 452.400 ;
        RECT 536.250 452.250 538.050 453.150 ;
        RECT 526.950 449.850 528.750 450.750 ;
        RECT 529.950 448.950 532.050 451.050 ;
        RECT 533.250 449.850 534.750 450.750 ;
        RECT 535.950 448.950 538.050 451.050 ;
        RECT 526.950 445.950 529.050 448.050 ;
        RECT 529.950 446.850 532.050 447.750 ;
        RECT 532.950 445.950 535.050 448.050 ;
        RECT 523.950 418.950 526.050 421.050 ;
        RECT 527.400 418.050 528.450 445.950 ;
        RECT 503.400 407.400 507.450 408.450 ;
        RECT 509.400 407.400 513.450 408.450 ;
        RECT 515.400 416.400 519.450 417.450 ;
        RECT 500.400 406.050 501.450 406.950 ;
        RECT 499.950 403.950 502.050 406.050 ;
        RECT 496.950 382.950 499.050 385.050 ;
        RECT 499.950 382.950 502.050 385.050 ;
        RECT 496.950 380.250 499.050 381.150 ;
        RECT 499.950 380.850 502.050 381.750 ;
        RECT 496.950 378.450 499.050 379.050 ;
        RECT 494.400 377.400 499.050 378.450 ;
        RECT 496.950 376.950 499.050 377.400 ;
        RECT 487.950 370.950 490.050 373.050 ;
        RECT 487.950 352.950 490.050 355.050 ;
        RECT 488.400 343.050 489.450 352.950 ;
        RECT 499.950 346.950 502.050 349.050 ;
        RECT 493.950 343.950 496.050 346.050 ;
        RECT 494.400 343.050 495.450 343.950 ;
        RECT 484.950 341.250 486.750 342.150 ;
        RECT 487.950 340.950 490.050 343.050 ;
        RECT 491.250 341.250 492.750 342.150 ;
        RECT 493.950 340.950 496.050 343.050 ;
        RECT 497.250 341.250 499.050 342.150 ;
        RECT 484.950 337.950 487.050 340.050 ;
        RECT 488.250 338.850 489.750 339.750 ;
        RECT 490.950 337.950 493.050 340.050 ;
        RECT 494.250 338.850 495.750 339.750 ;
        RECT 496.950 337.950 499.050 340.050 ;
        RECT 485.400 337.050 486.450 337.950 ;
        RECT 484.950 334.950 487.050 337.050 ;
        RECT 487.950 334.950 490.050 337.050 ;
        RECT 488.400 310.050 489.450 334.950 ;
        RECT 493.950 322.950 496.050 325.050 ;
        RECT 484.950 308.250 486.750 309.150 ;
        RECT 487.950 307.950 490.050 310.050 ;
        RECT 491.250 308.250 493.050 309.150 ;
        RECT 484.950 304.950 487.050 307.050 ;
        RECT 488.250 305.850 489.750 306.750 ;
        RECT 490.950 304.950 493.050 307.050 ;
        RECT 491.400 301.050 492.450 304.950 ;
        RECT 479.400 299.400 483.450 300.450 ;
        RECT 472.950 295.950 475.050 298.050 ;
        RECT 473.400 289.050 474.450 295.950 ;
        RECT 475.950 289.950 478.050 292.050 ;
        RECT 469.950 286.950 472.050 289.050 ;
        RECT 472.950 286.950 475.050 289.050 ;
        RECT 467.400 284.400 471.450 285.450 ;
        RECT 470.400 277.050 471.450 284.400 ;
        RECT 466.950 274.950 469.050 277.050 ;
        RECT 469.950 274.950 472.050 277.050 ;
        RECT 467.400 274.050 468.450 274.950 ;
        RECT 466.950 271.950 469.050 274.050 ;
        RECT 470.250 272.250 471.750 273.150 ;
        RECT 472.950 271.950 475.050 274.050 ;
        RECT 466.950 269.850 468.750 270.750 ;
        RECT 469.950 268.950 472.050 271.050 ;
        RECT 473.250 269.850 475.050 270.750 ;
        RECT 451.950 265.950 454.050 268.050 ;
        RECT 457.950 265.950 460.050 268.050 ;
        RECT 463.950 265.950 466.050 268.050 ;
        RECT 472.950 265.950 475.050 268.050 ;
        RECT 457.950 262.950 460.050 265.050 ;
        RECT 463.950 264.450 466.050 265.050 ;
        RECT 466.950 264.450 469.050 265.050 ;
        RECT 463.950 263.400 469.050 264.450 ;
        RECT 463.950 262.950 466.050 263.400 ;
        RECT 466.950 262.950 469.050 263.400 ;
        RECT 439.950 250.950 442.050 253.050 ;
        RECT 448.950 250.950 451.050 253.050 ;
        RECT 454.950 247.950 457.050 250.050 ;
        RECT 439.950 241.950 442.050 244.050 ;
        RECT 442.950 243.450 445.050 244.050 ;
        RECT 448.950 243.450 451.050 244.050 ;
        RECT 442.950 242.400 451.050 243.450 ;
        RECT 442.950 241.950 445.050 242.400 ;
        RECT 448.950 241.950 451.050 242.400 ;
        RECT 440.400 226.050 441.450 241.950 ;
        RECT 455.400 241.050 456.450 247.950 ;
        RECT 442.950 238.950 445.050 241.050 ;
        RECT 445.950 239.250 448.050 240.150 ;
        RECT 448.950 239.850 451.050 240.750 ;
        RECT 451.950 239.250 453.750 240.150 ;
        RECT 454.950 238.950 457.050 241.050 ;
        RECT 439.950 223.950 442.050 226.050 ;
        RECT 443.400 225.450 444.450 238.950 ;
        RECT 458.400 238.050 459.450 262.950 ;
        RECT 460.950 256.950 463.050 259.050 ;
        RECT 469.950 256.950 472.050 259.050 ;
        RECT 461.400 241.050 462.450 256.950 ;
        RECT 470.400 244.050 471.450 256.950 ;
        RECT 466.950 241.950 469.050 244.050 ;
        RECT 469.950 241.950 472.050 244.050 ;
        RECT 467.400 241.050 468.450 241.950 ;
        RECT 473.400 241.050 474.450 265.950 ;
        RECT 460.950 238.950 463.050 241.050 ;
        RECT 464.250 239.250 465.750 240.150 ;
        RECT 466.950 238.950 469.050 241.050 ;
        RECT 470.250 239.250 471.750 240.150 ;
        RECT 472.950 238.950 475.050 241.050 ;
        RECT 445.950 235.950 448.050 238.050 ;
        RECT 451.950 235.950 454.050 238.050 ;
        RECT 455.250 236.850 457.050 237.750 ;
        RECT 457.950 235.950 460.050 238.050 ;
        RECT 460.950 236.850 462.750 237.750 ;
        RECT 463.950 235.950 466.050 238.050 ;
        RECT 467.250 236.850 468.750 237.750 ;
        RECT 469.950 235.950 472.050 238.050 ;
        RECT 473.250 236.850 475.050 237.750 ;
        RECT 446.400 229.050 447.450 235.950 ;
        RECT 448.950 232.950 451.050 235.050 ;
        RECT 445.950 226.950 448.050 229.050 ;
        RECT 443.400 224.400 447.450 225.450 ;
        RECT 439.950 220.950 442.050 223.050 ;
        RECT 440.400 217.050 441.450 220.950 ;
        RECT 442.950 217.950 445.050 220.050 ;
        RECT 439.950 214.950 442.050 217.050 ;
        RECT 443.400 199.050 444.450 217.950 ;
        RECT 446.400 217.050 447.450 224.400 ;
        RECT 445.950 214.950 448.050 217.050 ;
        RECT 445.950 199.950 448.050 202.050 ;
        RECT 436.950 196.950 439.050 199.050 ;
        RECT 442.950 196.950 445.050 199.050 ;
        RECT 446.400 196.050 447.450 199.950 ;
        RECT 439.950 194.250 442.050 195.150 ;
        RECT 442.950 194.850 445.050 195.750 ;
        RECT 445.950 193.950 448.050 196.050 ;
        RECT 439.950 190.950 442.050 193.050 ;
        RECT 445.950 190.950 448.050 193.050 ;
        RECT 440.400 187.050 441.450 190.950 ;
        RECT 439.950 184.950 442.050 187.050 ;
        RECT 433.950 175.950 436.050 178.050 ;
        RECT 440.400 175.050 441.450 184.950 ;
        RECT 439.950 172.950 442.050 175.050 ;
        RECT 433.950 169.950 436.050 172.050 ;
        RECT 434.400 169.050 435.450 169.950 ;
        RECT 446.400 169.050 447.450 190.950 ;
        RECT 433.950 166.950 436.050 169.050 ;
        RECT 437.250 167.250 438.750 168.150 ;
        RECT 439.950 166.950 442.050 169.050 ;
        RECT 443.250 167.250 444.750 168.150 ;
        RECT 445.950 166.950 448.050 169.050 ;
        RECT 433.950 164.850 435.750 165.750 ;
        RECT 436.950 163.950 439.050 166.050 ;
        RECT 440.250 164.850 441.750 165.750 ;
        RECT 442.950 163.950 445.050 166.050 ;
        RECT 446.250 164.850 448.050 165.750 ;
        RECT 437.400 163.050 438.450 163.950 ;
        RECT 443.400 163.050 444.450 163.950 ;
        RECT 431.400 161.400 435.450 162.450 ;
        RECT 425.400 142.050 426.450 161.400 ;
        RECT 427.950 159.450 430.050 160.050 ;
        RECT 430.950 159.450 433.050 160.050 ;
        RECT 427.950 158.400 433.050 159.450 ;
        RECT 427.950 157.950 430.050 158.400 ;
        RECT 430.950 157.950 433.050 158.400 ;
        RECT 430.950 154.950 433.050 157.050 ;
        RECT 421.950 139.950 424.050 142.050 ;
        RECT 424.950 139.950 427.050 142.050 ;
        RECT 412.950 136.950 415.050 139.050 ;
        RECT 406.950 131.250 409.050 132.150 ;
        RECT 412.950 130.950 415.050 133.050 ;
        RECT 400.950 127.950 403.050 130.050 ;
        RECT 404.250 128.250 405.750 129.150 ;
        RECT 406.950 127.950 409.050 130.050 ;
        RECT 410.250 128.250 412.050 129.150 ;
        RECT 400.950 125.850 402.750 126.750 ;
        RECT 403.950 124.950 406.050 127.050 ;
        RECT 404.400 123.450 405.450 124.950 ;
        RECT 398.400 122.400 405.450 123.450 ;
        RECT 401.400 109.050 402.450 122.400 ;
        RECT 403.950 115.950 406.050 118.050 ;
        RECT 400.950 106.950 403.050 109.050 ;
        RECT 400.950 103.950 403.050 106.050 ;
        RECT 401.400 97.050 402.450 103.950 ;
        RECT 388.950 96.450 391.050 97.050 ;
        RECT 386.400 95.400 391.050 96.450 ;
        RECT 373.950 92.250 375.750 93.150 ;
        RECT 376.950 91.950 379.050 94.050 ;
        RECT 380.250 92.250 382.050 93.150 ;
        RECT 382.950 91.950 385.050 94.050 ;
        RECT 370.950 88.950 373.050 91.050 ;
        RECT 373.950 88.950 376.050 91.050 ;
        RECT 377.250 89.850 378.750 90.750 ;
        RECT 379.950 88.950 382.050 91.050 ;
        RECT 374.400 82.050 375.450 88.950 ;
        RECT 373.950 79.950 376.050 82.050 ;
        RECT 380.400 79.050 381.450 88.950 ;
        RECT 386.400 82.050 387.450 95.400 ;
        RECT 388.950 94.950 391.050 95.400 ;
        RECT 392.250 95.250 393.750 96.150 ;
        RECT 394.950 94.950 397.050 97.050 ;
        RECT 398.250 95.250 399.750 96.150 ;
        RECT 400.950 94.950 403.050 97.050 ;
        RECT 404.400 94.050 405.450 115.950 ;
        RECT 407.400 115.050 408.450 127.950 ;
        RECT 409.950 124.950 412.050 127.050 ;
        RECT 410.400 118.050 411.450 124.950 ;
        RECT 409.950 115.950 412.050 118.050 ;
        RECT 406.950 112.950 409.050 115.050 ;
        RECT 406.950 109.950 409.050 112.050 ;
        RECT 407.400 97.050 408.450 109.950 ;
        RECT 413.400 100.050 414.450 130.950 ;
        RECT 427.950 127.950 430.050 130.050 ;
        RECT 418.950 125.250 421.050 126.150 ;
        RECT 424.950 125.250 427.050 126.150 ;
        RECT 418.950 121.950 421.050 124.050 ;
        RECT 422.250 122.250 423.750 123.150 ;
        RECT 424.950 121.950 427.050 124.050 ;
        RECT 425.400 121.050 426.450 121.950 ;
        RECT 418.950 118.950 421.050 121.050 ;
        RECT 421.950 118.950 424.050 121.050 ;
        RECT 424.950 118.950 427.050 121.050 ;
        RECT 415.950 115.950 418.050 118.050 ;
        RECT 412.950 97.950 415.050 100.050 ;
        RECT 406.950 94.950 409.050 97.050 ;
        RECT 410.250 95.250 411.750 96.150 ;
        RECT 412.950 94.950 415.050 97.050 ;
        RECT 416.400 94.050 417.450 115.950 ;
        RECT 419.400 112.050 420.450 118.950 ;
        RECT 422.400 112.050 423.450 118.950 ;
        RECT 418.950 109.950 421.050 112.050 ;
        RECT 421.950 109.950 424.050 112.050 ;
        RECT 418.950 100.950 421.050 103.050 ;
        RECT 388.950 92.850 390.750 93.750 ;
        RECT 391.950 91.950 394.050 94.050 ;
        RECT 395.250 92.850 396.750 93.750 ;
        RECT 397.950 91.950 400.050 94.050 ;
        RECT 401.250 92.850 403.050 93.750 ;
        RECT 403.950 91.950 406.050 94.050 ;
        RECT 406.950 92.850 408.750 93.750 ;
        RECT 409.950 91.950 412.050 94.050 ;
        RECT 413.250 92.850 414.750 93.750 ;
        RECT 415.950 91.950 418.050 94.050 ;
        RECT 385.950 79.950 388.050 82.050 ;
        RECT 388.950 79.950 391.050 82.050 ;
        RECT 379.950 76.950 382.050 79.050 ;
        RECT 389.400 76.050 390.450 79.950 ;
        RECT 392.400 79.050 393.450 91.950 ;
        RECT 415.950 89.850 418.050 90.750 ;
        RECT 419.400 79.050 420.450 100.950 ;
        RECT 421.950 97.950 424.050 100.050 ;
        RECT 391.950 76.950 394.050 79.050 ;
        RECT 418.950 76.950 421.050 79.050 ;
        RECT 367.950 73.950 370.050 76.050 ;
        RECT 388.950 73.950 391.050 76.050 ;
        RECT 394.950 73.950 397.050 76.050 ;
        RECT 364.950 67.950 367.050 70.050 ;
        RECT 364.950 64.950 367.050 67.050 ;
        RECT 361.950 55.950 364.050 58.050 ;
        RECT 361.950 52.950 364.050 55.050 ;
        RECT 362.400 40.050 363.450 52.950 ;
        RECT 361.950 37.950 364.050 40.050 ;
        RECT 362.400 37.050 363.450 37.950 ;
        RECT 361.950 34.950 364.050 37.050 ;
        RECT 361.950 25.950 364.050 28.050 ;
        RECT 365.400 25.050 366.450 64.950 ;
        RECT 379.950 55.950 382.050 58.050 ;
        RECT 367.950 53.250 369.750 54.150 ;
        RECT 370.950 52.950 373.050 55.050 ;
        RECT 376.950 52.950 379.050 55.050 ;
        RECT 367.950 49.950 370.050 52.050 ;
        RECT 371.250 50.850 373.050 51.750 ;
        RECT 373.950 50.250 376.050 51.150 ;
        RECT 376.950 50.850 379.050 51.750 ;
        RECT 380.400 49.050 381.450 55.950 ;
        RECT 382.950 52.950 385.050 55.050 ;
        RECT 388.950 53.250 391.050 54.150 ;
        RECT 395.400 52.050 396.450 73.950 ;
        RECT 412.950 67.950 415.050 70.050 ;
        RECT 406.950 56.250 409.050 57.150 ;
        RECT 413.400 55.050 414.450 67.950 ;
        RECT 422.400 58.050 423.450 97.950 ;
        RECT 424.950 94.950 427.050 97.050 ;
        RECT 425.400 58.050 426.450 94.950 ;
        RECT 428.400 94.050 429.450 127.950 ;
        RECT 431.400 121.050 432.450 154.950 ;
        RECT 430.950 118.950 433.050 121.050 ;
        RECT 434.400 115.050 435.450 161.400 ;
        RECT 436.950 160.950 439.050 163.050 ;
        RECT 442.950 160.950 445.050 163.050 ;
        RECT 439.950 154.950 442.050 157.050 ;
        RECT 436.950 151.950 439.050 154.050 ;
        RECT 430.950 112.950 433.050 115.050 ;
        RECT 433.950 112.950 436.050 115.050 ;
        RECT 427.950 91.950 430.050 94.050 ;
        RECT 431.400 91.050 432.450 112.950 ;
        RECT 437.400 112.050 438.450 151.950 ;
        RECT 440.400 145.050 441.450 154.950 ;
        RECT 442.950 151.950 445.050 154.050 ;
        RECT 439.950 142.950 442.050 145.050 ;
        RECT 443.400 127.050 444.450 151.950 ;
        RECT 445.950 139.950 448.050 142.050 ;
        RECT 449.400 141.450 450.450 232.950 ;
        RECT 452.400 226.050 453.450 235.950 ;
        RECT 451.950 223.950 454.050 226.050 ;
        RECT 457.950 220.950 460.050 223.050 ;
        RECT 451.950 214.950 454.050 217.050 ;
        RECT 452.400 193.050 453.450 214.950 ;
        RECT 458.400 199.050 459.450 220.950 ;
        RECT 470.400 220.050 471.450 235.950 ;
        RECT 469.950 217.950 472.050 220.050 ;
        RECT 472.950 211.950 475.050 214.050 ;
        RECT 473.400 199.050 474.450 211.950 ;
        RECT 476.400 199.050 477.450 289.950 ;
        RECT 479.400 241.050 480.450 299.400 ;
        RECT 490.950 298.950 493.050 301.050 ;
        RECT 484.950 283.950 487.050 286.050 ;
        RECT 485.400 277.050 486.450 283.950 ;
        RECT 490.950 280.950 493.050 283.050 ;
        RECT 491.400 277.050 492.450 280.950 ;
        RECT 484.950 274.950 487.050 277.050 ;
        RECT 490.950 274.950 493.050 277.050 ;
        RECT 494.400 274.050 495.450 322.950 ;
        RECT 497.400 322.050 498.450 337.950 ;
        RECT 496.950 319.950 499.050 322.050 ;
        RECT 500.400 312.450 501.450 346.950 ;
        RECT 503.400 337.050 504.450 407.400 ;
        RECT 505.950 352.950 508.050 355.050 ;
        RECT 506.400 343.050 507.450 352.950 ;
        RECT 509.400 343.050 510.450 407.400 ;
        RECT 511.950 403.950 514.050 406.050 ;
        RECT 512.400 385.050 513.450 403.950 ;
        RECT 511.950 382.950 514.050 385.050 ;
        RECT 511.950 380.850 514.050 381.750 ;
        RECT 505.950 340.950 508.050 343.050 ;
        RECT 508.950 340.950 511.050 343.050 ;
        RECT 505.950 338.850 508.050 339.750 ;
        RECT 508.950 338.250 511.050 339.150 ;
        RECT 502.950 334.950 505.050 337.050 ;
        RECT 508.950 334.950 511.050 337.050 ;
        RECT 502.950 313.950 505.050 316.050 ;
        RECT 497.400 311.400 501.450 312.450 ;
        RECT 497.400 292.050 498.450 311.400 ;
        RECT 503.400 310.050 504.450 313.950 ;
        RECT 509.400 313.050 510.450 334.950 ;
        RECT 515.400 319.050 516.450 416.400 ;
        RECT 526.950 415.950 529.050 418.050 ;
        RECT 533.400 415.050 534.450 445.950 ;
        RECT 536.400 415.050 537.450 448.950 ;
        RECT 538.950 415.950 541.050 418.050 ;
        RECT 539.400 415.050 540.450 415.950 ;
        RECT 517.950 412.950 520.050 415.050 ;
        RECT 520.950 413.250 523.050 414.150 ;
        RECT 526.950 413.250 529.050 414.150 ;
        RECT 529.950 412.950 532.050 415.050 ;
        RECT 532.950 412.950 535.050 415.050 ;
        RECT 535.950 412.950 538.050 415.050 ;
        RECT 538.950 412.950 541.050 415.050 ;
        RECT 542.250 413.250 544.050 414.150 ;
        RECT 518.400 411.450 519.450 412.950 ;
        RECT 520.950 411.450 523.050 412.050 ;
        RECT 518.400 410.400 523.050 411.450 ;
        RECT 526.950 411.450 529.050 412.050 ;
        RECT 530.400 411.450 531.450 412.950 ;
        RECT 520.950 409.950 523.050 410.400 ;
        RECT 524.250 410.250 525.750 411.150 ;
        RECT 526.950 410.400 531.450 411.450 ;
        RECT 532.950 410.850 535.050 411.750 ;
        RECT 526.950 409.950 529.050 410.400 ;
        RECT 530.400 409.050 531.450 410.400 ;
        RECT 535.950 410.250 538.050 411.150 ;
        RECT 538.950 410.850 540.750 411.750 ;
        RECT 541.950 409.950 544.050 412.050 ;
        RECT 523.950 406.950 526.050 409.050 ;
        RECT 529.950 406.950 532.050 409.050 ;
        RECT 535.950 406.950 538.050 409.050 ;
        RECT 524.400 403.050 525.450 406.950 ;
        RECT 523.950 400.950 526.050 403.050 ;
        RECT 536.400 400.050 537.450 406.950 ;
        RECT 535.950 397.950 538.050 400.050 ;
        RECT 542.400 385.050 543.450 409.950 ;
        RECT 520.950 382.950 523.050 385.050 ;
        RECT 523.950 382.950 526.050 385.050 ;
        RECT 541.950 382.950 544.050 385.050 ;
        RECT 517.950 380.850 520.050 381.750 ;
        RECT 521.400 355.050 522.450 382.950 ;
        RECT 520.950 352.950 523.050 355.050 ;
        RECT 524.400 343.050 525.450 382.950 ;
        RECT 529.950 379.950 532.050 382.050 ;
        RECT 535.950 379.950 538.050 382.050 ;
        RECT 539.250 380.250 541.050 381.150 ;
        RECT 541.950 379.950 544.050 382.050 ;
        RECT 545.400 381.450 546.450 517.950 ;
        RECT 554.400 493.050 555.450 520.950 ;
        RECT 550.950 491.250 553.050 492.150 ;
        RECT 553.950 490.950 556.050 493.050 ;
        RECT 563.400 492.450 564.450 523.950 ;
        RECT 563.400 491.400 567.450 492.450 ;
        RECT 547.950 488.250 549.750 489.150 ;
        RECT 550.950 487.950 553.050 490.050 ;
        RECT 556.950 489.450 559.050 490.050 ;
        RECT 554.250 488.250 555.750 489.150 ;
        RECT 556.950 488.400 561.450 489.450 ;
        RECT 556.950 487.950 559.050 488.400 ;
        RECT 547.950 484.950 550.050 487.050 ;
        RECT 553.950 484.950 556.050 487.050 ;
        RECT 557.250 485.850 559.050 486.750 ;
        RECT 554.400 483.450 555.450 484.950 ;
        RECT 554.400 482.400 558.450 483.450 ;
        RECT 553.950 457.950 556.050 460.050 ;
        RECT 550.950 455.250 553.050 456.150 ;
        RECT 553.950 455.850 556.050 456.750 ;
        RECT 550.950 451.950 553.050 454.050 ;
        RECT 551.400 436.050 552.450 451.950 ;
        RECT 550.950 433.950 553.050 436.050 ;
        RECT 557.400 415.050 558.450 482.400 ;
        RECT 560.400 460.050 561.450 488.400 ;
        RECT 566.400 487.050 567.450 491.400 ;
        RECT 565.950 484.950 568.050 487.050 ;
        RECT 565.950 482.850 568.050 483.750 ;
        RECT 565.950 475.950 568.050 478.050 ;
        RECT 559.950 457.950 562.050 460.050 ;
        RECT 562.950 457.950 565.050 460.050 ;
        RECT 559.950 455.250 562.050 456.150 ;
        RECT 559.950 453.450 562.050 454.050 ;
        RECT 563.400 453.450 564.450 457.950 ;
        RECT 559.950 452.400 564.450 453.450 ;
        RECT 559.950 451.950 562.050 452.400 ;
        RECT 562.950 433.950 565.050 436.050 ;
        RECT 559.950 415.950 562.050 418.050 ;
        RECT 560.400 415.050 561.450 415.950 ;
        RECT 550.950 414.450 553.050 415.050 ;
        RECT 550.950 413.400 555.450 414.450 ;
        RECT 550.950 412.950 553.050 413.400 ;
        RECT 547.950 410.250 550.050 411.150 ;
        RECT 550.950 410.850 553.050 411.750 ;
        RECT 547.950 406.950 550.050 409.050 ;
        RECT 554.400 408.450 555.450 413.400 ;
        RECT 556.950 412.950 559.050 415.050 ;
        RECT 559.950 412.950 562.050 415.050 ;
        RECT 556.950 410.250 559.050 411.150 ;
        RECT 559.950 410.850 562.050 411.750 ;
        RECT 556.950 408.450 559.050 409.050 ;
        RECT 554.400 407.400 559.050 408.450 ;
        RECT 556.950 406.950 559.050 407.400 ;
        RECT 556.950 403.950 559.050 406.050 ;
        RECT 547.950 383.250 550.050 384.150 ;
        RECT 547.950 381.450 550.050 382.050 ;
        RECT 545.400 380.400 550.050 381.450 ;
        RECT 547.950 379.950 550.050 380.400 ;
        RECT 526.950 376.950 529.050 379.050 ;
        RECT 529.950 377.850 531.750 378.750 ;
        RECT 532.950 376.950 535.050 379.050 ;
        RECT 536.250 377.850 537.750 378.750 ;
        RECT 538.950 376.950 541.050 379.050 ;
        RECT 527.400 358.050 528.450 376.950 ;
        RECT 532.950 374.850 535.050 375.750 ;
        RECT 532.950 361.950 535.050 364.050 ;
        RECT 526.950 355.950 529.050 358.050 ;
        RECT 520.950 341.250 523.050 342.150 ;
        RECT 523.950 340.950 526.050 343.050 ;
        RECT 526.950 341.250 529.050 342.150 ;
        RECT 529.950 341.250 532.050 342.150 ;
        RECT 520.950 339.450 523.050 340.050 ;
        RECT 518.400 338.400 523.050 339.450 ;
        RECT 518.400 322.050 519.450 338.400 ;
        RECT 520.950 337.950 523.050 338.400 ;
        RECT 524.250 338.250 525.750 339.150 ;
        RECT 526.950 337.950 529.050 340.050 ;
        RECT 529.950 337.950 532.050 340.050 ;
        RECT 523.950 336.450 526.050 337.050 ;
        RECT 521.400 335.400 526.050 336.450 ;
        RECT 517.950 319.950 520.050 322.050 ;
        RECT 514.950 316.950 517.050 319.050 ;
        RECT 521.400 316.050 522.450 335.400 ;
        RECT 523.950 334.950 526.050 335.400 ;
        RECT 527.400 333.450 528.450 337.950 ;
        RECT 533.400 337.050 534.450 361.950 ;
        RECT 538.950 352.950 541.050 355.050 ;
        RECT 535.950 341.250 538.050 342.150 ;
        RECT 539.400 339.450 540.450 352.950 ;
        RECT 542.400 346.050 543.450 379.950 ;
        RECT 548.400 355.050 549.450 379.950 ;
        RECT 557.400 379.050 558.450 403.950 ;
        RECT 563.400 394.050 564.450 433.950 ;
        RECT 562.950 391.950 565.050 394.050 ;
        RECT 559.950 381.450 562.050 382.050 ;
        RECT 563.400 381.450 564.450 391.950 ;
        RECT 559.950 380.400 564.450 381.450 ;
        RECT 559.950 379.950 562.050 380.400 ;
        RECT 556.950 376.950 559.050 379.050 ;
        RECT 559.950 377.850 562.050 378.750 ;
        RECT 566.400 373.050 567.450 475.950 ;
        RECT 569.400 400.050 570.450 541.950 ;
        RECT 571.950 529.950 574.050 532.050 ;
        RECT 571.950 527.850 574.050 528.750 ;
        RECT 574.950 527.250 577.050 528.150 ;
        RECT 574.950 523.950 577.050 526.050 ;
        RECT 571.950 508.950 574.050 511.050 ;
        RECT 572.400 460.050 573.450 508.950 ;
        RECT 578.400 492.450 579.450 571.950 ;
        RECT 580.950 556.950 583.050 559.050 ;
        RECT 587.400 556.050 588.450 634.950 ;
        RECT 592.950 629.250 595.050 630.150 ;
        RECT 595.950 628.950 598.050 631.050 ;
        RECT 598.950 628.950 601.050 631.050 ;
        RECT 589.950 626.250 591.750 627.150 ;
        RECT 592.950 625.950 595.050 628.050 ;
        RECT 593.400 625.050 594.450 625.950 ;
        RECT 589.950 622.950 592.050 625.050 ;
        RECT 592.950 622.950 595.050 625.050 ;
        RECT 590.400 622.050 591.450 622.950 ;
        RECT 589.950 619.950 592.050 622.050 ;
        RECT 596.400 621.450 597.450 628.950 ;
        RECT 605.400 628.050 606.450 635.400 ;
        RECT 610.950 635.250 613.050 636.150 ;
        RECT 613.950 634.950 616.050 637.050 ;
        RECT 617.400 634.050 618.450 661.950 ;
        RECT 623.400 640.050 624.450 667.950 ;
        RECT 629.400 666.450 630.450 671.400 ;
        RECT 626.400 665.400 630.450 666.450 ;
        RECT 622.950 637.950 625.050 640.050 ;
        RECT 607.950 632.250 609.750 633.150 ;
        RECT 610.950 631.950 613.050 634.050 ;
        RECT 614.250 632.250 615.750 633.150 ;
        RECT 616.950 631.950 619.050 634.050 ;
        RECT 607.950 628.950 610.050 631.050 ;
        RECT 598.950 626.850 601.050 627.750 ;
        RECT 604.950 625.950 607.050 628.050 ;
        RECT 593.400 620.400 597.450 621.450 ;
        RECT 593.400 598.050 594.450 620.400 ;
        RECT 605.400 607.050 606.450 625.950 ;
        RECT 604.950 604.950 607.050 607.050 ;
        RECT 608.400 604.050 609.450 628.950 ;
        RECT 611.400 616.050 612.450 631.950 ;
        RECT 613.950 628.950 616.050 631.050 ;
        RECT 617.250 629.850 619.050 630.750 ;
        RECT 614.400 625.050 615.450 628.950 ;
        RECT 616.950 625.950 619.050 628.050 ;
        RECT 613.950 622.950 616.050 625.050 ;
        RECT 610.950 613.950 613.050 616.050 ;
        RECT 598.950 601.950 601.050 604.050 ;
        RECT 604.950 601.950 607.050 604.050 ;
        RECT 607.950 601.950 610.050 604.050 ;
        RECT 595.950 599.250 598.050 600.150 ;
        RECT 598.950 599.850 601.050 600.750 ;
        RECT 601.950 598.950 604.050 601.050 ;
        RECT 592.950 595.950 595.050 598.050 ;
        RECT 595.950 595.950 598.050 598.050 ;
        RECT 602.400 592.050 603.450 598.950 ;
        RECT 605.400 594.450 606.450 601.950 ;
        RECT 607.950 596.250 609.750 597.150 ;
        RECT 610.950 595.950 613.050 598.050 ;
        RECT 614.250 596.250 616.050 597.150 ;
        RECT 607.950 594.450 610.050 595.050 ;
        RECT 605.400 593.400 610.050 594.450 ;
        RECT 611.250 593.850 612.750 594.750 ;
        RECT 601.950 589.950 604.050 592.050 ;
        RECT 592.950 560.250 595.050 561.150 ;
        RECT 592.950 558.450 595.050 559.050 ;
        RECT 590.400 557.400 595.050 558.450 ;
        RECT 580.950 554.850 583.050 555.750 ;
        RECT 583.950 554.250 586.050 555.150 ;
        RECT 586.950 553.950 589.050 556.050 ;
        RECT 583.950 550.950 586.050 553.050 ;
        RECT 580.950 544.950 583.050 547.050 ;
        RECT 581.400 520.050 582.450 544.950 ;
        RECT 584.400 541.050 585.450 550.950 ;
        RECT 583.950 538.950 586.050 541.050 ;
        RECT 590.400 535.050 591.450 557.400 ;
        RECT 592.950 556.950 595.050 557.400 ;
        RECT 596.250 557.250 597.750 558.150 ;
        RECT 598.950 556.950 601.050 559.050 ;
        RECT 602.250 557.250 604.050 558.150 ;
        RECT 605.400 556.050 606.450 593.400 ;
        RECT 607.950 592.950 610.050 593.400 ;
        RECT 613.950 592.950 616.050 595.050 ;
        RECT 617.400 589.050 618.450 625.950 ;
        RECT 623.400 616.050 624.450 637.950 ;
        RECT 619.950 613.950 622.050 616.050 ;
        RECT 622.950 613.950 625.050 616.050 ;
        RECT 620.400 595.050 621.450 613.950 ;
        RECT 626.400 610.050 627.450 665.400 ;
        RECT 632.400 664.050 633.450 694.950 ;
        RECT 646.950 679.950 649.050 682.050 ;
        RECT 637.950 673.950 640.050 676.050 ;
        RECT 638.400 673.050 639.450 673.950 ;
        RECT 634.950 670.950 637.050 673.050 ;
        RECT 637.950 670.950 640.050 673.050 ;
        RECT 641.250 671.250 642.750 672.150 ;
        RECT 643.950 670.950 646.050 673.050 ;
        RECT 635.400 670.050 636.450 670.950 ;
        RECT 634.950 667.950 637.050 670.050 ;
        RECT 638.250 668.850 639.750 669.750 ;
        RECT 640.950 667.950 643.050 670.050 ;
        RECT 644.250 668.850 646.050 669.750 ;
        RECT 647.400 669.450 648.450 679.950 ;
        RECT 649.950 671.250 652.050 672.150 ;
        RECT 652.950 670.950 655.050 673.050 ;
        RECT 649.950 669.450 652.050 670.050 ;
        RECT 647.400 668.400 652.050 669.450 ;
        RECT 649.950 667.950 652.050 668.400 ;
        RECT 653.400 667.050 654.450 670.950 ;
        RECT 659.400 670.050 660.450 704.400 ;
        RECT 661.950 703.950 664.050 704.400 ;
        RECT 665.250 704.250 666.750 705.150 ;
        RECT 667.950 703.950 670.050 706.050 ;
        RECT 671.250 704.250 673.050 705.150 ;
        RECT 674.400 703.050 675.450 706.950 ;
        RECT 677.400 706.050 678.450 710.400 ;
        RECT 685.950 706.950 688.050 709.050 ;
        RECT 686.400 706.050 687.450 706.950 ;
        RECT 676.950 703.950 679.050 706.050 ;
        RECT 679.950 703.950 682.050 706.050 ;
        RECT 683.250 704.250 684.750 705.150 ;
        RECT 685.950 703.950 688.050 706.050 ;
        RECT 661.950 701.850 663.750 702.750 ;
        RECT 664.950 700.950 667.050 703.050 ;
        RECT 670.950 702.450 673.050 703.050 ;
        RECT 673.950 702.450 676.050 703.050 ;
        RECT 670.950 701.400 676.050 702.450 ;
        RECT 679.950 701.850 681.750 702.750 ;
        RECT 670.950 700.950 673.050 701.400 ;
        RECT 673.950 700.950 676.050 701.400 ;
        RECT 682.950 700.950 685.050 703.050 ;
        RECT 686.250 701.850 688.050 702.750 ;
        RECT 665.400 700.050 666.450 700.950 ;
        RECT 664.950 697.950 667.050 700.050 ;
        RECT 664.950 691.950 667.050 694.050 ;
        RECT 658.950 667.950 661.050 670.050 ;
        RECT 661.950 667.950 664.050 670.050 ;
        RECT 634.950 665.850 637.050 666.750 ;
        RECT 640.950 664.950 643.050 667.050 ;
        RECT 652.950 664.950 655.050 667.050 ;
        RECT 661.950 665.850 664.050 666.750 ;
        RECT 631.950 661.950 634.050 664.050 ;
        RECT 634.950 635.250 637.050 636.150 ;
        RECT 628.950 631.950 631.050 634.050 ;
        RECT 632.250 632.250 633.750 633.150 ;
        RECT 634.950 631.950 637.050 634.050 ;
        RECT 638.250 632.250 640.050 633.150 ;
        RECT 628.950 629.850 630.750 630.750 ;
        RECT 631.950 628.950 634.050 631.050 ;
        RECT 635.400 625.050 636.450 631.950 ;
        RECT 637.950 628.950 640.050 631.050 ;
        RECT 638.400 628.050 639.450 628.950 ;
        RECT 637.950 625.950 640.050 628.050 ;
        RECT 634.950 622.950 637.050 625.050 ;
        RECT 635.400 619.050 636.450 622.950 ;
        RECT 638.400 622.050 639.450 625.950 ;
        RECT 637.950 619.950 640.050 622.050 ;
        RECT 634.950 616.950 637.050 619.050 ;
        RECT 634.950 613.950 637.050 616.050 ;
        RECT 625.950 607.950 628.050 610.050 ;
        RECT 622.950 601.950 625.050 604.050 ;
        RECT 619.950 592.950 622.050 595.050 ;
        RECT 616.950 586.950 619.050 589.050 ;
        RECT 617.400 565.050 618.450 586.950 ;
        RECT 619.950 565.950 622.050 568.050 ;
        RECT 616.950 562.950 619.050 565.050 ;
        RECT 620.400 559.050 621.450 565.950 ;
        RECT 613.950 557.250 616.050 558.150 ;
        RECT 616.950 556.950 619.050 559.050 ;
        RECT 619.950 556.950 622.050 559.050 ;
        RECT 595.950 553.950 598.050 556.050 ;
        RECT 599.250 554.850 600.750 555.750 ;
        RECT 601.950 553.950 604.050 556.050 ;
        RECT 604.950 553.950 607.050 556.050 ;
        RECT 610.950 554.250 612.750 555.150 ;
        RECT 613.950 553.950 616.050 556.050 ;
        RECT 602.400 541.050 603.450 553.950 ;
        RECT 610.950 550.950 613.050 553.050 ;
        RECT 613.950 550.950 616.050 553.050 ;
        RECT 614.400 547.050 615.450 550.950 ;
        RECT 613.950 544.950 616.050 547.050 ;
        RECT 601.950 538.950 604.050 541.050 ;
        RECT 589.950 532.950 592.050 535.050 ;
        RECT 590.400 526.050 591.450 532.950 ;
        RECT 595.950 529.950 598.050 532.050 ;
        RECT 601.950 531.450 604.050 532.050 ;
        RECT 604.950 531.450 607.050 532.050 ;
        RECT 601.950 530.400 607.050 531.450 ;
        RECT 601.950 529.950 604.050 530.400 ;
        RECT 604.950 529.950 607.050 530.400 ;
        RECT 586.950 524.250 588.750 525.150 ;
        RECT 589.950 523.950 592.050 526.050 ;
        RECT 593.250 524.250 595.050 525.150 ;
        RECT 586.950 520.950 589.050 523.050 ;
        RECT 590.250 521.850 591.750 522.750 ;
        RECT 592.950 520.950 595.050 523.050 ;
        RECT 580.950 517.950 583.050 520.050 ;
        RECT 587.400 511.050 588.450 520.950 ;
        RECT 593.400 520.050 594.450 520.950 ;
        RECT 592.950 517.950 595.050 520.050 ;
        RECT 596.400 511.050 597.450 529.950 ;
        RECT 614.400 529.050 615.450 544.950 ;
        RECT 617.400 538.050 618.450 556.950 ;
        RECT 619.950 554.850 622.050 555.750 ;
        RECT 616.950 535.950 619.050 538.050 ;
        RECT 617.400 532.050 618.450 535.950 ;
        RECT 616.950 529.950 619.050 532.050 ;
        RECT 619.950 529.950 622.050 532.050 ;
        RECT 620.400 529.050 621.450 529.950 ;
        RECT 598.950 526.950 601.050 529.050 ;
        RECT 602.250 527.850 603.750 528.750 ;
        RECT 604.950 526.950 607.050 529.050 ;
        RECT 607.950 526.950 610.050 529.050 ;
        RECT 613.950 526.950 616.050 529.050 ;
        RECT 617.250 527.850 618.750 528.750 ;
        RECT 619.950 526.950 622.050 529.050 ;
        RECT 598.950 524.850 601.050 525.750 ;
        RECT 604.950 524.850 607.050 525.750 ;
        RECT 586.950 508.950 589.050 511.050 ;
        RECT 595.950 508.950 598.050 511.050 ;
        RECT 586.800 497.100 588.900 499.200 ;
        RECT 587.550 493.350 588.750 497.100 ;
        RECT 589.950 494.850 592.050 496.950 ;
        RECT 578.400 491.400 582.450 492.450 ;
        RECT 577.950 488.250 580.050 489.150 ;
        RECT 577.950 486.450 580.050 487.050 ;
        RECT 575.400 485.400 580.050 486.450 ;
        RECT 575.400 484.050 576.450 485.400 ;
        RECT 577.950 484.950 580.050 485.400 ;
        RECT 574.950 481.950 577.050 484.050 ;
        RECT 571.950 457.950 574.050 460.050 ;
        RECT 571.950 453.450 574.050 454.050 ;
        RECT 575.400 453.450 576.450 481.950 ;
        RECT 581.400 469.050 582.450 491.400 ;
        RECT 586.950 491.250 589.050 493.350 ;
        RECT 587.550 477.600 588.750 491.250 ;
        RECT 590.250 477.600 591.450 494.850 ;
        RECT 597.900 494.400 600.000 496.500 ;
        RECT 601.950 494.400 604.050 496.500 ;
        RECT 592.950 491.250 595.050 493.350 ;
        RECT 593.400 477.600 594.600 491.250 ;
        RECT 598.350 485.550 599.550 494.400 ;
        RECT 602.550 488.250 603.750 494.400 ;
        RECT 601.950 486.150 604.050 488.250 ;
        RECT 597.750 483.450 599.850 485.550 ;
        RECT 598.350 477.600 599.550 483.450 ;
        RECT 602.550 477.600 603.750 486.150 ;
        RECT 604.950 482.250 607.050 483.150 ;
        RECT 604.950 480.450 607.050 481.050 ;
        RECT 608.400 480.450 609.450 526.950 ;
        RECT 613.950 524.850 616.050 525.750 ;
        RECT 619.950 524.850 622.050 525.750 ;
        RECT 623.400 517.050 624.450 601.950 ;
        RECT 628.950 598.950 631.050 601.050 ;
        RECT 629.400 598.050 630.450 598.950 ;
        RECT 625.950 596.250 627.750 597.150 ;
        RECT 628.950 595.950 631.050 598.050 ;
        RECT 632.250 596.250 634.050 597.150 ;
        RECT 625.950 592.950 628.050 595.050 ;
        RECT 629.250 593.850 630.750 594.750 ;
        RECT 631.950 592.950 634.050 595.050 ;
        RECT 632.400 592.050 633.450 592.950 ;
        RECT 631.950 589.950 634.050 592.050 ;
        RECT 635.400 577.050 636.450 613.950 ;
        RECT 641.400 604.050 642.450 664.950 ;
        RECT 643.950 631.950 646.050 634.050 ;
        RECT 665.400 633.450 666.450 691.950 ;
        RECT 683.400 685.050 684.450 700.950 ;
        RECT 689.400 697.050 690.450 733.950 ;
        RECT 701.400 706.050 702.450 743.400 ;
        RECT 707.400 736.050 708.450 746.400 ;
        RECT 709.950 745.950 712.050 746.400 ;
        RECT 715.950 745.950 718.050 748.050 ;
        RECT 709.950 743.850 712.050 744.750 ;
        RECT 712.950 743.250 715.050 744.150 ;
        RECT 712.950 741.450 715.050 742.050 ;
        RECT 716.400 741.450 717.450 745.950 ;
        RECT 712.950 740.400 717.450 741.450 ;
        RECT 725.400 741.450 726.450 763.950 ;
        RECT 733.950 748.950 736.050 751.050 ;
        RECT 734.400 745.050 735.450 748.950 ;
        RECT 736.950 745.950 739.050 748.050 ;
        RECT 727.950 743.250 730.050 744.150 ;
        RECT 733.950 742.950 736.050 745.050 ;
        RECT 737.250 743.850 739.050 744.750 ;
        RECT 727.950 741.450 730.050 742.050 ;
        RECT 725.400 740.400 730.050 741.450 ;
        RECT 733.950 740.850 736.050 741.750 ;
        RECT 712.950 739.950 715.050 740.400 ;
        RECT 727.950 739.950 730.050 740.400 ;
        RECT 706.950 733.950 709.050 736.050 ;
        RECT 740.400 706.050 741.450 772.950 ;
        RECT 746.400 771.450 747.450 776.400 ;
        RECT 749.400 774.450 750.450 808.950 ;
        RECT 767.400 802.050 768.450 808.950 ;
        RECT 773.400 808.050 774.450 808.950 ;
        RECT 772.950 805.950 775.050 808.050 ;
        RECT 778.950 806.850 781.050 807.750 ;
        RECT 763.950 799.950 766.050 802.050 ;
        RECT 766.950 799.950 769.050 802.050 ;
        RECT 757.950 781.950 760.050 784.050 ;
        RECT 751.950 776.250 754.050 777.150 ;
        RECT 758.400 775.050 759.450 781.950 ;
        RECT 751.950 774.450 754.050 775.050 ;
        RECT 749.400 773.400 754.050 774.450 ;
        RECT 751.950 772.950 754.050 773.400 ;
        RECT 755.250 773.250 756.750 774.150 ;
        RECT 757.950 772.950 760.050 775.050 ;
        RECT 761.250 773.250 763.050 774.150 ;
        RECT 746.400 770.400 750.450 771.450 ;
        RECT 742.950 748.950 745.050 751.050 ;
        RECT 743.400 742.050 744.450 748.950 ;
        RECT 749.400 748.050 750.450 770.400 ;
        RECT 752.400 748.050 753.450 772.950 ;
        RECT 754.950 769.950 757.050 772.050 ;
        RECT 758.250 770.850 759.750 771.750 ;
        RECT 760.950 769.950 763.050 772.050 ;
        RECT 754.950 766.950 757.050 769.050 ;
        RECT 745.950 745.950 748.050 748.050 ;
        RECT 748.950 745.950 751.050 748.050 ;
        RECT 751.950 745.950 754.050 748.050 ;
        RECT 746.400 745.050 747.450 745.950 ;
        RECT 745.950 742.950 748.050 745.050 ;
        RECT 749.250 743.250 750.750 744.150 ;
        RECT 751.950 742.950 754.050 745.050 ;
        RECT 755.400 742.050 756.450 766.950 ;
        RECT 761.400 760.050 762.450 769.950 ;
        RECT 764.400 768.450 765.450 799.950 ;
        RECT 769.950 773.250 772.050 774.150 ;
        RECT 766.950 770.250 768.750 771.150 ;
        RECT 769.950 769.950 772.050 772.050 ;
        RECT 770.400 769.050 771.450 769.950 ;
        RECT 773.400 769.050 774.450 805.950 ;
        RECT 778.950 781.950 781.050 784.050 ;
        RECT 775.950 775.950 778.050 778.050 ;
        RECT 776.400 775.050 777.450 775.950 ;
        RECT 775.950 772.950 778.050 775.050 ;
        RECT 775.950 770.850 778.050 771.750 ;
        RECT 766.950 768.450 769.050 769.050 ;
        RECT 764.400 767.400 769.050 768.450 ;
        RECT 766.950 766.950 769.050 767.400 ;
        RECT 769.950 766.950 772.050 769.050 ;
        RECT 772.950 766.950 775.050 769.050 ;
        RECT 779.400 760.050 780.450 781.950 ;
        RECT 785.400 780.450 786.450 808.950 ;
        RECT 788.400 808.050 789.450 815.400 ;
        RECT 791.400 814.050 792.450 817.950 ;
        RECT 797.400 817.050 798.450 820.950 ;
        RECT 811.950 817.950 814.050 820.050 ;
        RECT 820.950 817.950 823.050 820.050 ;
        RECT 829.950 817.950 832.050 820.050 ;
        RECT 838.950 817.950 841.050 820.050 ;
        RECT 793.950 814.950 796.050 817.050 ;
        RECT 796.950 814.950 799.050 817.050 ;
        RECT 800.250 815.250 801.750 816.150 ;
        RECT 802.950 814.950 805.050 817.050 ;
        RECT 805.950 814.950 808.050 817.050 ;
        RECT 811.950 815.850 814.050 816.750 ;
        RECT 814.950 815.250 817.050 816.150 ;
        RECT 817.950 814.950 820.050 817.050 ;
        RECT 794.400 814.050 795.450 814.950 ;
        RECT 790.950 811.950 793.050 814.050 ;
        RECT 793.950 811.950 796.050 814.050 ;
        RECT 797.250 812.850 798.750 813.750 ;
        RECT 799.950 811.950 802.050 814.050 ;
        RECT 803.250 812.850 805.050 813.750 ;
        RECT 787.950 805.950 790.050 808.050 ;
        RECT 791.400 781.050 792.450 811.950 ;
        RECT 793.950 809.850 796.050 810.750 ;
        RECT 800.400 810.450 801.450 811.950 ;
        RECT 806.400 810.450 807.450 814.950 ;
        RECT 811.950 811.950 814.050 814.050 ;
        RECT 814.950 813.450 817.050 814.050 ;
        RECT 818.400 813.450 819.450 814.950 ;
        RECT 814.950 812.400 819.450 813.450 ;
        RECT 814.950 811.950 817.050 812.400 ;
        RECT 800.400 809.400 807.450 810.450 ;
        RECT 793.950 802.950 796.050 805.050 ;
        RECT 785.400 779.400 789.450 780.450 ;
        RECT 788.400 778.050 789.450 779.400 ;
        RECT 790.950 778.950 793.050 781.050 ;
        RECT 794.400 778.050 795.450 802.950 ;
        RECT 802.950 778.950 805.050 781.050 ;
        RECT 803.400 778.050 804.450 778.950 ;
        RECT 787.950 775.950 790.050 778.050 ;
        RECT 791.250 776.250 792.750 777.150 ;
        RECT 793.950 775.950 796.050 778.050 ;
        RECT 802.950 775.950 805.050 778.050 ;
        RECT 806.250 776.250 807.750 777.150 ;
        RECT 808.950 775.950 811.050 778.050 ;
        RECT 787.950 773.850 789.750 774.750 ;
        RECT 790.950 772.950 793.050 775.050 ;
        RECT 794.250 773.850 796.050 774.750 ;
        RECT 802.950 773.850 804.750 774.750 ;
        RECT 805.950 772.950 808.050 775.050 ;
        RECT 809.250 773.850 811.050 774.750 ;
        RECT 760.950 757.950 763.050 760.050 ;
        RECT 772.950 757.950 775.050 760.050 ;
        RECT 778.950 757.950 781.050 760.050 ;
        RECT 761.400 757.050 762.450 757.950 ;
        RECT 760.950 754.950 763.050 757.050 ;
        RECT 763.950 748.950 766.050 751.050 ;
        RECT 764.400 748.050 765.450 748.950 ;
        RECT 763.950 745.950 766.050 748.050 ;
        RECT 766.950 745.950 769.050 748.050 ;
        RECT 769.950 745.950 772.050 748.050 ;
        RECT 767.400 745.050 768.450 745.950 ;
        RECT 760.950 744.450 763.050 745.050 ;
        RECT 758.400 743.400 763.050 744.450 ;
        RECT 764.250 743.850 765.750 744.750 ;
        RECT 742.950 739.950 745.050 742.050 ;
        RECT 745.950 740.850 747.750 741.750 ;
        RECT 748.950 739.950 751.050 742.050 ;
        RECT 752.250 740.850 753.750 741.750 ;
        RECT 754.950 739.950 757.050 742.050 ;
        RECT 754.950 737.850 757.050 738.750 ;
        RECT 758.400 727.050 759.450 743.400 ;
        RECT 760.950 742.950 763.050 743.400 ;
        RECT 766.950 742.950 769.050 745.050 ;
        RECT 760.950 740.850 763.050 741.750 ;
        RECT 766.950 740.850 769.050 741.750 ;
        RECT 757.950 724.950 760.050 727.050 ;
        RECT 766.950 724.950 769.050 727.050 ;
        RECT 751.950 715.950 754.050 718.050 ;
        RECT 748.950 706.950 751.050 709.050 ;
        RECT 749.400 706.050 750.450 706.950 ;
        RECT 752.400 706.050 753.450 715.950 ;
        RECT 694.950 704.250 697.050 705.150 ;
        RECT 700.950 703.950 703.050 706.050 ;
        RECT 724.950 703.950 727.050 706.050 ;
        RECT 736.950 703.950 739.050 706.050 ;
        RECT 739.950 703.950 742.050 706.050 ;
        RECT 742.950 703.950 745.050 706.050 ;
        RECT 746.250 704.250 747.750 705.150 ;
        RECT 748.950 703.950 751.050 706.050 ;
        RECT 751.950 703.950 754.050 706.050 ;
        RECT 763.950 704.250 766.050 705.150 ;
        RECT 701.400 703.050 702.450 703.950 ;
        RECT 725.400 703.050 726.450 703.950 ;
        RECT 694.950 700.950 697.050 703.050 ;
        RECT 698.250 701.250 699.750 702.150 ;
        RECT 700.950 700.950 703.050 703.050 ;
        RECT 704.250 701.250 706.050 702.150 ;
        RECT 715.950 700.950 718.050 703.050 ;
        RECT 721.950 701.250 723.750 702.150 ;
        RECT 724.950 700.950 727.050 703.050 ;
        RECT 730.950 701.250 733.050 702.150 ;
        RECT 697.950 697.950 700.050 700.050 ;
        RECT 701.250 698.850 702.750 699.750 ;
        RECT 703.950 697.950 706.050 700.050 ;
        RECT 715.950 698.850 718.050 699.750 ;
        RECT 721.950 697.950 724.050 700.050 ;
        RECT 725.250 698.850 727.050 699.750 ;
        RECT 730.950 697.950 733.050 700.050 ;
        RECT 688.950 694.950 691.050 697.050 ;
        RECT 698.400 694.050 699.450 697.950 ;
        RECT 731.400 697.050 732.450 697.950 ;
        RECT 724.950 694.950 727.050 697.050 ;
        RECT 730.950 694.950 733.050 697.050 ;
        RECT 697.950 691.950 700.050 694.050 ;
        RECT 682.950 682.950 685.050 685.050 ;
        RECT 691.950 682.950 694.050 685.050 ;
        RECT 670.950 677.400 673.050 679.500 ;
        RECT 673.950 677.400 676.050 679.500 ;
        RECT 676.950 677.400 679.050 679.500 ;
        RECT 681.750 677.400 683.850 679.500 ;
        RECT 685.950 677.400 688.050 679.500 ;
        RECT 671.550 663.750 672.750 677.400 ;
        RECT 670.950 661.650 673.050 663.750 ;
        RECT 671.550 657.900 672.750 661.650 ;
        RECT 674.250 660.150 675.450 677.400 ;
        RECT 677.400 663.750 678.600 677.400 ;
        RECT 682.350 671.550 683.550 677.400 ;
        RECT 681.750 669.450 683.850 671.550 ;
        RECT 676.950 661.650 679.050 663.750 ;
        RECT 682.350 660.600 683.550 669.450 ;
        RECT 686.550 668.850 687.750 677.400 ;
        RECT 688.950 673.950 691.050 676.050 ;
        RECT 688.950 671.850 691.050 672.750 ;
        RECT 685.950 666.750 688.050 668.850 ;
        RECT 686.550 660.600 687.750 666.750 ;
        RECT 673.950 658.050 676.050 660.150 ;
        RECT 681.900 658.500 684.000 660.600 ;
        RECT 685.950 658.500 688.050 660.600 ;
        RECT 670.800 655.800 672.900 657.900 ;
        RECT 676.950 655.950 679.050 658.050 ;
        RECT 662.400 632.400 669.450 633.450 ;
        RECT 644.400 619.050 645.450 631.950 ;
        RECT 646.950 628.950 649.050 631.050 ;
        RECT 652.950 628.950 655.050 631.050 ;
        RECT 656.250 629.250 658.050 630.150 ;
        RECT 658.950 628.950 661.050 631.050 ;
        RECT 646.950 626.850 649.050 627.750 ;
        RECT 649.950 626.250 652.050 627.150 ;
        RECT 652.950 626.850 654.750 627.750 ;
        RECT 655.950 625.950 658.050 628.050 ;
        RECT 659.400 625.050 660.450 628.950 ;
        RECT 649.950 622.950 652.050 625.050 ;
        RECT 658.950 622.950 661.050 625.050 ;
        RECT 643.950 616.950 646.050 619.050 ;
        RECT 643.950 610.950 646.050 613.050 ;
        RECT 640.950 601.950 643.050 604.050 ;
        RECT 644.400 601.050 645.450 610.950 ;
        RECT 649.950 607.950 652.050 610.050 ;
        RECT 643.950 598.950 646.050 601.050 ;
        RECT 644.400 598.050 645.450 598.950 ;
        RECT 637.950 595.950 640.050 598.050 ;
        RECT 640.950 595.950 643.050 598.050 ;
        RECT 643.950 595.950 646.050 598.050 ;
        RECT 647.250 596.250 649.050 597.150 ;
        RECT 641.400 595.050 642.450 595.950 ;
        RECT 637.950 593.850 639.750 594.750 ;
        RECT 640.950 592.950 643.050 595.050 ;
        RECT 644.250 593.850 645.750 594.750 ;
        RECT 646.950 592.950 649.050 595.050 ;
        RECT 647.400 592.050 648.450 592.950 ;
        RECT 640.950 590.850 643.050 591.750 ;
        RECT 646.950 589.950 649.050 592.050 ;
        RECT 650.400 583.050 651.450 607.950 ;
        RECT 655.950 601.950 658.050 604.050 ;
        RECT 652.950 598.950 655.050 601.050 ;
        RECT 655.950 599.850 657.750 600.750 ;
        RECT 658.950 598.950 661.050 601.050 ;
        RECT 653.400 598.050 654.450 598.950 ;
        RECT 652.950 595.950 655.050 598.050 ;
        RECT 658.950 596.850 661.050 597.750 ;
        RECT 649.950 580.950 652.050 583.050 ;
        RECT 649.950 577.950 652.050 580.050 ;
        RECT 634.950 574.950 637.050 577.050 ;
        RECT 640.950 574.950 643.050 577.050 ;
        RECT 628.950 559.950 631.050 562.050 ;
        RECT 632.250 560.250 633.750 561.150 ;
        RECT 634.950 559.950 637.050 562.050 ;
        RECT 641.400 559.050 642.450 574.950 ;
        RECT 646.950 560.250 649.050 561.150 ;
        RECT 628.950 557.850 630.750 558.750 ;
        RECT 631.950 556.950 634.050 559.050 ;
        RECT 635.250 557.850 637.050 558.750 ;
        RECT 637.950 557.250 639.750 558.150 ;
        RECT 640.950 556.950 643.050 559.050 ;
        RECT 646.950 558.450 649.050 559.050 ;
        RECT 650.400 558.450 651.450 577.950 ;
        RECT 644.250 557.250 645.750 558.150 ;
        RECT 646.950 557.400 651.450 558.450 ;
        RECT 646.950 556.950 649.050 557.400 ;
        RECT 625.950 553.950 628.050 556.050 ;
        RECT 626.400 544.050 627.450 553.950 ;
        RECT 632.400 550.050 633.450 556.950 ;
        RECT 634.950 553.950 637.050 556.050 ;
        RECT 637.950 553.950 640.050 556.050 ;
        RECT 641.250 554.850 642.750 555.750 ;
        RECT 643.950 553.950 646.050 556.050 ;
        RECT 631.950 547.950 634.050 550.050 ;
        RECT 635.400 547.050 636.450 553.950 ;
        RECT 650.400 547.050 651.450 557.400 ;
        RECT 653.400 550.050 654.450 595.950 ;
        RECT 658.950 592.950 661.050 595.050 ;
        RECT 655.950 580.950 658.050 583.050 ;
        RECT 656.400 559.050 657.450 580.950 ;
        RECT 659.400 568.050 660.450 592.950 ;
        RECT 658.950 565.950 661.050 568.050 ;
        RECT 662.400 561.450 663.450 632.400 ;
        RECT 668.400 631.050 669.450 632.400 ;
        RECT 673.950 632.250 676.050 633.150 ;
        RECT 677.400 631.050 678.450 655.950 ;
        RECT 692.400 643.050 693.450 682.950 ;
        RECT 694.950 676.950 697.050 679.050 ;
        RECT 697.950 676.950 700.050 679.050 ;
        RECT 700.950 676.950 703.050 679.050 ;
        RECT 695.250 658.050 696.450 676.950 ;
        RECT 698.250 664.350 699.450 676.950 ;
        RECT 697.950 662.250 700.050 664.350 ;
        RECT 698.250 658.050 699.450 662.250 ;
        RECT 701.250 658.050 702.450 676.950 ;
        RECT 725.400 670.050 726.450 694.950 ;
        RECT 737.400 675.450 738.450 703.950 ;
        RECT 742.950 701.850 744.750 702.750 ;
        RECT 745.950 700.950 748.050 703.050 ;
        RECT 749.250 701.850 751.050 702.750 ;
        RECT 751.950 700.950 754.050 703.050 ;
        RECT 754.950 701.250 756.750 702.150 ;
        RECT 757.950 700.950 760.050 703.050 ;
        RECT 761.250 701.250 762.750 702.150 ;
        RECT 763.950 700.950 766.050 703.050 ;
        RECT 746.400 700.050 747.450 700.950 ;
        RECT 745.950 697.950 748.050 700.050 ;
        RECT 752.400 694.050 753.450 700.950 ;
        RECT 754.950 697.950 757.050 700.050 ;
        RECT 758.250 698.850 759.750 699.750 ;
        RECT 760.950 697.950 763.050 700.050 ;
        RECT 764.400 697.050 765.450 700.950 ;
        RECT 763.950 694.950 766.050 697.050 ;
        RECT 767.400 694.050 768.450 724.950 ;
        RECT 770.400 718.050 771.450 745.950 ;
        RECT 769.950 715.950 772.050 718.050 ;
        RECT 769.950 706.950 772.050 709.050 ;
        RECT 751.950 691.950 754.050 694.050 ;
        RECT 760.950 691.950 763.050 694.050 ;
        RECT 766.950 691.950 769.050 694.050 ;
        RECT 737.400 674.400 741.450 675.450 ;
        RECT 736.950 671.250 739.050 672.150 ;
        RECT 712.950 668.250 715.050 669.150 ;
        RECT 715.950 667.950 718.050 670.050 ;
        RECT 721.950 668.250 723.750 669.150 ;
        RECT 724.950 667.950 727.050 670.050 ;
        RECT 728.250 668.250 730.050 669.150 ;
        RECT 706.950 665.850 709.050 666.750 ;
        RECT 712.950 664.950 715.050 667.050 ;
        RECT 694.950 655.950 697.050 658.050 ;
        RECT 697.950 655.950 700.050 658.050 ;
        RECT 700.950 655.950 703.050 658.050 ;
        RECT 691.950 640.950 694.050 643.050 ;
        RECT 697.950 640.950 700.050 643.050 ;
        RECT 691.950 637.950 694.050 640.050 ;
        RECT 685.950 632.250 688.050 633.150 ;
        RECT 692.400 631.050 693.450 637.950 ;
        RECT 664.950 629.250 666.750 630.150 ;
        RECT 667.950 628.950 670.050 631.050 ;
        RECT 671.250 629.250 672.750 630.150 ;
        RECT 673.950 628.950 676.050 631.050 ;
        RECT 676.950 628.950 679.050 631.050 ;
        RECT 685.950 628.950 688.050 631.050 ;
        RECT 689.250 629.250 690.750 630.150 ;
        RECT 691.950 628.950 694.050 631.050 ;
        RECT 695.250 629.250 697.050 630.150 ;
        RECT 674.400 628.050 675.450 628.950 ;
        RECT 664.950 625.950 667.050 628.050 ;
        RECT 668.250 626.850 669.750 627.750 ;
        RECT 670.950 625.950 673.050 628.050 ;
        RECT 673.950 625.950 676.050 628.050 ;
        RECT 688.950 625.950 691.050 628.050 ;
        RECT 692.250 626.850 693.750 627.750 ;
        RECT 694.950 625.950 697.050 628.050 ;
        RECT 665.400 619.050 666.450 625.950 ;
        RECT 671.400 625.050 672.450 625.950 ;
        RECT 667.950 622.950 670.050 625.050 ;
        RECT 670.950 622.950 673.050 625.050 ;
        RECT 664.950 616.950 667.050 619.050 ;
        RECT 664.950 599.250 667.050 600.150 ;
        RECT 664.950 595.950 667.050 598.050 ;
        RECT 668.400 592.050 669.450 622.950 ;
        RECT 679.950 613.950 682.050 616.050 ;
        RECT 680.400 601.050 681.450 613.950 ;
        RECT 695.400 610.050 696.450 625.950 ;
        RECT 694.950 607.950 697.050 610.050 ;
        RECT 695.400 607.050 696.450 607.950 ;
        RECT 691.950 604.950 694.050 607.050 ;
        RECT 694.950 604.950 697.050 607.050 ;
        RECT 673.950 600.450 676.050 601.050 ;
        RECT 671.400 599.400 676.050 600.450 ;
        RECT 667.950 589.950 670.050 592.050 ;
        RECT 671.400 586.050 672.450 599.400 ;
        RECT 673.950 598.950 676.050 599.400 ;
        RECT 677.250 599.250 678.750 600.150 ;
        RECT 679.950 598.950 682.050 601.050 ;
        RECT 683.250 599.250 684.750 600.150 ;
        RECT 685.950 598.950 688.050 601.050 ;
        RECT 673.950 596.850 675.750 597.750 ;
        RECT 676.950 595.950 679.050 598.050 ;
        RECT 680.250 596.850 681.750 597.750 ;
        RECT 682.950 595.950 685.050 598.050 ;
        RECT 686.250 596.850 688.050 597.750 ;
        RECT 677.400 592.050 678.450 595.950 ;
        RECT 673.950 589.950 676.050 592.050 ;
        RECT 676.950 589.950 679.050 592.050 ;
        RECT 670.950 583.950 673.050 586.050 ;
        RECT 664.950 561.450 667.050 562.050 ;
        RECT 658.950 560.250 661.050 561.150 ;
        RECT 662.400 560.400 667.050 561.450 ;
        RECT 664.950 559.950 667.050 560.400 ;
        RECT 665.400 559.050 666.450 559.950 ;
        RECT 655.950 556.950 658.050 559.050 ;
        RECT 658.950 556.950 661.050 559.050 ;
        RECT 662.250 557.250 663.750 558.150 ;
        RECT 664.950 556.950 667.050 559.050 ;
        RECT 668.250 557.250 670.050 558.150 ;
        RECT 659.400 556.050 660.450 556.950 ;
        RECT 658.950 553.950 661.050 556.050 ;
        RECT 661.950 553.950 664.050 556.050 ;
        RECT 665.250 554.850 666.750 555.750 ;
        RECT 667.950 553.950 670.050 556.050 ;
        RECT 652.950 547.950 655.050 550.050 ;
        RECT 634.950 544.950 637.050 547.050 ;
        RECT 646.950 544.950 649.050 547.050 ;
        RECT 649.950 544.950 652.050 547.050 ;
        RECT 655.950 544.950 658.050 547.050 ;
        RECT 625.950 541.950 628.050 544.050 ;
        RECT 640.950 535.950 643.050 538.050 ;
        RECT 625.950 532.950 628.050 535.050 ;
        RECT 626.400 532.050 627.450 532.950 ;
        RECT 625.950 529.950 628.050 532.050 ;
        RECT 641.400 529.050 642.450 535.950 ;
        RECT 647.400 529.050 648.450 544.950 ;
        RECT 649.950 538.950 652.050 541.050 ;
        RECT 625.950 527.850 628.050 528.750 ;
        RECT 628.950 527.250 631.050 528.150 ;
        RECT 640.950 526.950 643.050 529.050 ;
        RECT 644.250 527.250 645.750 528.150 ;
        RECT 646.950 526.950 649.050 529.050 ;
        RECT 650.400 526.050 651.450 538.950 ;
        RECT 656.400 529.050 657.450 544.950 ;
        RECT 658.950 541.950 661.050 544.050 ;
        RECT 659.400 532.050 660.450 541.950 ;
        RECT 662.400 532.050 663.450 553.950 ;
        RECT 658.950 529.950 661.050 532.050 ;
        RECT 661.950 529.950 664.050 532.050 ;
        RECT 674.400 529.050 675.450 589.950 ;
        RECT 688.950 586.950 691.050 589.050 ;
        RECT 679.950 565.950 682.050 568.050 ;
        RECT 676.950 556.950 679.050 559.050 ;
        RECT 676.950 554.850 679.050 555.750 ;
        RECT 680.400 555.450 681.450 565.950 ;
        RECT 682.950 557.250 685.050 558.150 ;
        RECT 682.950 555.450 685.050 556.050 ;
        RECT 680.400 554.400 685.050 555.450 ;
        RECT 682.950 553.950 685.050 554.400 ;
        RECT 686.250 554.250 688.050 555.150 ;
        RECT 689.400 553.050 690.450 586.950 ;
        RECT 685.950 550.950 688.050 553.050 ;
        RECT 688.950 550.950 691.050 553.050 ;
        RECT 686.400 550.050 687.450 550.950 ;
        RECT 685.950 547.950 688.050 550.050 ;
        RECT 682.950 544.950 685.050 547.050 ;
        RECT 655.950 526.950 658.050 529.050 ;
        RECT 659.250 527.850 660.750 528.750 ;
        RECT 661.950 528.450 664.050 529.050 ;
        RECT 661.950 527.400 666.450 528.450 ;
        RECT 661.950 526.950 664.050 527.400 ;
        RECT 628.950 523.950 631.050 526.050 ;
        RECT 640.950 524.850 642.750 525.750 ;
        RECT 643.950 523.950 646.050 526.050 ;
        RECT 647.250 524.850 648.750 525.750 ;
        RECT 649.950 523.950 652.050 526.050 ;
        RECT 655.950 524.850 658.050 525.750 ;
        RECT 661.950 524.850 664.050 525.750 ;
        RECT 665.400 523.050 666.450 527.400 ;
        RECT 673.950 526.950 676.050 529.050 ;
        RECT 673.950 524.250 675.750 525.150 ;
        RECT 676.950 523.950 679.050 526.050 ;
        RECT 683.400 525.450 684.450 544.950 ;
        RECT 685.950 527.250 688.050 528.150 ;
        RECT 688.950 526.950 691.050 529.050 ;
        RECT 685.950 525.450 688.050 526.050 ;
        RECT 680.250 524.250 682.050 525.150 ;
        RECT 683.400 524.400 688.050 525.450 ;
        RECT 649.950 521.850 652.050 522.750 ;
        RECT 652.950 520.950 655.050 523.050 ;
        RECT 664.950 520.950 667.050 523.050 ;
        RECT 673.950 520.950 676.050 523.050 ;
        RECT 677.250 521.850 678.750 522.750 ;
        RECT 679.950 522.450 682.050 523.050 ;
        RECT 683.400 522.450 684.450 524.400 ;
        RECT 685.950 523.950 688.050 524.400 ;
        RECT 679.950 521.400 684.450 522.450 ;
        RECT 679.950 520.950 682.050 521.400 ;
        RECT 622.950 514.950 625.050 517.050 ;
        RECT 640.950 514.950 643.050 517.050 ;
        RECT 610.950 496.950 613.050 499.050 ;
        RECT 613.950 496.950 616.050 499.050 ;
        RECT 616.950 496.950 619.050 499.050 ;
        RECT 604.950 479.400 609.450 480.450 ;
        RECT 604.950 478.950 607.050 479.400 ;
        RECT 611.250 478.050 612.450 496.950 ;
        RECT 614.250 492.750 615.450 496.950 ;
        RECT 613.950 490.650 616.050 492.750 ;
        RECT 614.250 478.050 615.450 490.650 ;
        RECT 617.250 478.050 618.450 496.950 ;
        RECT 622.950 488.250 625.050 489.150 ;
        RECT 628.950 487.950 631.050 490.050 ;
        RECT 634.950 487.950 637.050 490.050 ;
        RECT 628.950 485.850 631.050 486.750 ;
        RECT 619.950 481.950 622.050 484.050 ;
        RECT 586.950 475.500 589.050 477.600 ;
        RECT 589.950 475.500 592.050 477.600 ;
        RECT 592.950 475.500 595.050 477.600 ;
        RECT 597.750 475.500 599.850 477.600 ;
        RECT 601.950 475.500 604.050 477.600 ;
        RECT 610.950 475.950 613.050 478.050 ;
        RECT 613.950 475.950 616.050 478.050 ;
        RECT 616.950 475.950 619.050 478.050 ;
        RECT 616.950 472.950 619.050 475.050 ;
        RECT 580.950 466.950 583.050 469.050 ;
        RECT 580.950 461.400 583.050 463.500 ;
        RECT 583.950 461.400 586.050 463.500 ;
        RECT 586.950 461.400 589.050 463.500 ;
        RECT 591.750 461.400 593.850 463.500 ;
        RECT 595.950 461.400 598.050 463.500 ;
        RECT 571.950 452.400 576.450 453.450 ;
        RECT 571.950 451.950 574.050 452.400 ;
        RECT 571.950 449.850 574.050 450.750 ;
        RECT 575.400 436.050 576.450 452.400 ;
        RECT 581.550 447.750 582.750 461.400 ;
        RECT 580.950 445.650 583.050 447.750 ;
        RECT 581.550 441.900 582.750 445.650 ;
        RECT 584.250 444.150 585.450 461.400 ;
        RECT 587.400 447.750 588.600 461.400 ;
        RECT 592.350 455.550 593.550 461.400 ;
        RECT 591.750 453.450 593.850 455.550 ;
        RECT 586.950 445.650 589.050 447.750 ;
        RECT 592.350 444.600 593.550 453.450 ;
        RECT 596.550 452.850 597.750 461.400 ;
        RECT 598.950 460.950 601.050 463.050 ;
        RECT 604.950 460.950 607.050 463.050 ;
        RECT 607.950 460.950 610.050 463.050 ;
        RECT 610.950 460.950 613.050 463.050 ;
        RECT 599.400 460.050 600.450 460.950 ;
        RECT 598.950 457.950 601.050 460.050 ;
        RECT 598.950 455.850 601.050 456.750 ;
        RECT 595.950 450.750 598.050 452.850 ;
        RECT 596.550 444.600 597.750 450.750 ;
        RECT 583.950 442.050 586.050 444.150 ;
        RECT 591.900 442.500 594.000 444.600 ;
        RECT 595.950 442.500 598.050 444.600 ;
        RECT 605.250 442.050 606.450 460.950 ;
        RECT 608.250 448.350 609.450 460.950 ;
        RECT 607.950 446.250 610.050 448.350 ;
        RECT 608.250 442.050 609.450 446.250 ;
        RECT 611.250 442.050 612.450 460.950 ;
        RECT 617.400 454.050 618.450 472.950 ;
        RECT 616.950 451.950 619.050 454.050 ;
        RECT 616.950 449.850 619.050 450.750 ;
        RECT 616.950 445.950 619.050 448.050 ;
        RECT 580.800 439.800 582.900 441.900 ;
        RECT 604.950 439.950 607.050 442.050 ;
        RECT 607.950 439.950 610.050 442.050 ;
        RECT 610.950 439.950 613.050 442.050 ;
        RECT 574.950 433.950 577.050 436.050 ;
        RECT 586.950 433.950 589.050 436.050 ;
        RECT 587.400 415.050 588.450 433.950 ;
        RECT 617.400 424.050 618.450 445.950 ;
        RECT 616.950 421.950 619.050 424.050 ;
        RECT 610.950 418.950 613.050 421.050 ;
        RECT 620.400 420.450 621.450 481.950 ;
        RECT 635.400 475.050 636.450 487.950 ;
        RECT 634.950 472.950 637.050 475.050 ;
        RECT 631.950 457.950 634.050 460.050 ;
        RECT 637.950 457.950 640.050 460.050 ;
        RECT 631.950 455.850 634.050 456.750 ;
        RECT 634.950 455.250 637.050 456.150 ;
        RECT 622.950 452.250 625.050 453.150 ;
        RECT 631.950 451.950 634.050 454.050 ;
        RECT 634.950 453.450 637.050 454.050 ;
        RECT 638.400 453.450 639.450 457.950 ;
        RECT 634.950 452.400 639.450 453.450 ;
        RECT 634.950 451.950 637.050 452.400 ;
        RECT 617.400 419.400 621.450 420.450 ;
        RECT 571.950 413.250 574.050 414.150 ;
        RECT 577.950 413.250 580.050 414.150 ;
        RECT 586.950 412.950 589.050 415.050 ;
        RECT 571.950 409.950 574.050 412.050 ;
        RECT 586.950 410.850 589.050 411.750 ;
        RECT 607.950 410.850 610.050 411.750 ;
        RECT 572.400 403.050 573.450 409.950 ;
        RECT 571.950 400.950 574.050 403.050 ;
        RECT 568.950 397.950 571.050 400.050 ;
        RECT 607.950 397.950 610.050 400.050 ;
        RECT 568.950 389.400 571.050 391.500 ;
        RECT 571.950 389.400 574.050 391.500 ;
        RECT 574.950 389.400 577.050 391.500 ;
        RECT 579.750 389.400 581.850 391.500 ;
        RECT 583.950 389.400 586.050 391.500 ;
        RECT 569.550 375.750 570.750 389.400 ;
        RECT 568.950 373.650 571.050 375.750 ;
        RECT 565.950 370.950 568.050 373.050 ;
        RECT 553.950 367.950 556.050 370.050 ;
        RECT 556.950 367.950 559.050 370.050 ;
        RECT 569.550 369.900 570.750 373.650 ;
        RECT 572.250 372.150 573.450 389.400 ;
        RECT 575.400 375.750 576.600 389.400 ;
        RECT 580.350 383.550 581.550 389.400 ;
        RECT 579.750 381.450 581.850 383.550 ;
        RECT 574.950 373.650 577.050 375.750 ;
        RECT 580.350 372.600 581.550 381.450 ;
        RECT 584.550 380.850 585.750 389.400 ;
        RECT 592.950 388.950 595.050 391.050 ;
        RECT 595.950 388.950 598.050 391.050 ;
        RECT 598.950 388.950 601.050 391.050 ;
        RECT 586.950 387.450 589.050 388.050 ;
        RECT 586.950 386.400 591.450 387.450 ;
        RECT 586.950 385.950 589.050 386.400 ;
        RECT 586.950 383.850 589.050 384.750 ;
        RECT 583.950 378.750 586.050 380.850 ;
        RECT 584.550 372.600 585.750 378.750 ;
        RECT 571.950 370.050 574.050 372.150 ;
        RECT 579.900 370.500 582.000 372.600 ;
        RECT 583.950 370.500 586.050 372.600 ;
        RECT 547.950 352.950 550.050 355.050 ;
        RECT 541.950 343.950 544.050 346.050 ;
        RECT 541.950 341.250 544.050 342.150 ;
        RECT 547.950 341.250 550.050 342.150 ;
        RECT 541.950 339.450 544.050 340.050 ;
        RECT 539.400 338.400 544.050 339.450 ;
        RECT 541.950 337.950 544.050 338.400 ;
        RECT 529.950 334.950 532.050 337.050 ;
        RECT 532.950 334.950 535.050 337.050 ;
        RECT 524.400 332.400 528.450 333.450 ;
        RECT 524.400 331.050 525.450 332.400 ;
        RECT 523.950 328.950 526.050 331.050 ;
        RECT 514.950 313.950 517.050 316.050 ;
        RECT 520.950 313.950 523.050 316.050 ;
        RECT 524.400 313.050 525.450 328.950 ;
        RECT 508.950 310.950 511.050 313.050 ;
        RECT 514.950 311.850 517.050 312.750 ;
        RECT 517.950 311.250 520.050 312.150 ;
        RECT 523.950 310.950 526.050 313.050 ;
        RECT 499.950 308.250 501.750 309.150 ;
        RECT 502.950 307.950 505.050 310.050 ;
        RECT 508.950 307.950 511.050 310.050 ;
        RECT 517.950 307.950 520.050 310.050 ;
        RECT 520.950 307.950 523.050 310.050 ;
        RECT 499.950 304.950 502.050 307.050 ;
        RECT 503.250 305.850 504.750 306.750 ;
        RECT 505.950 304.950 508.050 307.050 ;
        RECT 509.250 305.850 511.050 306.750 ;
        RECT 496.950 289.950 499.050 292.050 ;
        RECT 500.400 283.050 501.450 304.950 ;
        RECT 505.950 302.850 508.050 303.750 ;
        RECT 508.950 301.950 511.050 304.050 ;
        RECT 499.950 280.950 502.050 283.050 ;
        RECT 496.950 274.950 499.050 277.050 ;
        RECT 481.950 271.950 484.050 274.050 ;
        RECT 487.950 273.450 490.050 274.050 ;
        RECT 485.250 272.250 486.750 273.150 ;
        RECT 487.950 272.400 492.450 273.450 ;
        RECT 487.950 271.950 490.050 272.400 ;
        RECT 481.950 269.850 483.750 270.750 ;
        RECT 484.950 268.950 487.050 271.050 ;
        RECT 488.250 269.850 490.050 270.750 ;
        RECT 481.950 265.950 484.050 268.050 ;
        RECT 478.950 238.950 481.050 241.050 ;
        RECT 482.400 229.050 483.450 265.950 ;
        RECT 485.400 265.050 486.450 268.950 ;
        RECT 491.400 267.450 492.450 272.400 ;
        RECT 493.950 271.950 496.050 274.050 ;
        RECT 497.400 271.050 498.450 274.950 ;
        RECT 502.950 271.950 505.050 274.050 ;
        RECT 503.400 271.050 504.450 271.950 ;
        RECT 493.950 269.250 495.750 270.150 ;
        RECT 496.950 268.950 499.050 271.050 ;
        RECT 500.250 269.250 501.750 270.150 ;
        RECT 502.950 268.950 505.050 271.050 ;
        RECT 506.250 269.250 508.050 270.150 ;
        RECT 488.400 266.400 492.450 267.450 ;
        RECT 484.950 262.950 487.050 265.050 ;
        RECT 488.400 259.050 489.450 266.400 ;
        RECT 493.950 265.950 496.050 268.050 ;
        RECT 497.250 266.850 498.750 267.750 ;
        RECT 499.950 265.950 502.050 268.050 ;
        RECT 503.250 266.850 504.750 267.750 ;
        RECT 505.950 265.950 508.050 268.050 ;
        RECT 490.950 262.950 493.050 265.050 ;
        RECT 494.400 264.450 495.450 265.950 ;
        RECT 500.400 265.050 501.450 265.950 ;
        RECT 509.400 265.050 510.450 301.950 ;
        RECT 511.950 295.950 514.050 298.050 ;
        RECT 512.400 268.050 513.450 295.950 ;
        RECT 521.400 295.050 522.450 307.950 ;
        RECT 520.950 292.950 523.050 295.050 ;
        RECT 514.950 271.950 517.050 274.050 ;
        RECT 511.950 265.950 514.050 268.050 ;
        RECT 494.400 263.400 498.450 264.450 ;
        RECT 487.950 256.950 490.050 259.050 ;
        RECT 487.950 241.950 490.050 244.050 ;
        RECT 488.400 238.050 489.450 241.950 ;
        RECT 484.950 236.250 486.750 237.150 ;
        RECT 487.950 235.950 490.050 238.050 ;
        RECT 491.400 235.050 492.450 262.950 ;
        RECT 493.950 253.950 496.050 256.050 ;
        RECT 494.400 244.050 495.450 253.950 ;
        RECT 493.950 241.950 496.050 244.050 ;
        RECT 493.950 238.950 496.050 241.050 ;
        RECT 494.400 238.050 495.450 238.950 ;
        RECT 493.950 235.950 496.050 238.050 ;
        RECT 484.950 232.950 487.050 235.050 ;
        RECT 488.250 233.850 489.750 234.750 ;
        RECT 490.950 232.950 493.050 235.050 ;
        RECT 494.250 233.850 496.050 234.750 ;
        RECT 481.950 226.950 484.050 229.050 ;
        RECT 485.400 214.050 486.450 232.950 ;
        RECT 490.950 230.850 493.050 231.750 ;
        RECT 487.950 226.950 490.050 229.050 ;
        RECT 484.950 211.950 487.050 214.050 ;
        RECT 484.950 199.950 487.050 202.050 ;
        RECT 454.950 197.250 456.750 198.150 ;
        RECT 457.950 196.950 460.050 199.050 ;
        RECT 461.250 197.250 462.750 198.150 ;
        RECT 463.950 196.950 466.050 199.050 ;
        RECT 467.250 197.250 469.050 198.150 ;
        RECT 469.950 196.950 472.050 199.050 ;
        RECT 472.950 196.950 475.050 199.050 ;
        RECT 475.950 196.950 478.050 199.050 ;
        RECT 478.950 196.950 481.050 199.050 ;
        RECT 482.250 197.250 484.050 198.150 ;
        RECT 454.950 193.950 457.050 196.050 ;
        RECT 458.250 194.850 459.750 195.750 ;
        RECT 460.950 193.950 463.050 196.050 ;
        RECT 464.250 194.850 465.750 195.750 ;
        RECT 466.950 193.950 469.050 196.050 ;
        RECT 451.950 190.950 454.050 193.050 ;
        RECT 451.950 187.950 454.050 190.050 ;
        RECT 452.400 172.050 453.450 187.950 ;
        RECT 455.400 172.050 456.450 193.950 ;
        RECT 457.950 172.950 460.050 175.050 ;
        RECT 451.950 169.950 454.050 172.050 ;
        RECT 454.950 169.950 457.050 172.050 ;
        RECT 458.400 169.050 459.450 172.950 ;
        RECT 451.950 166.950 454.050 169.050 ;
        RECT 455.250 167.250 456.750 168.150 ;
        RECT 457.950 166.950 460.050 169.050 ;
        RECT 461.400 166.050 462.450 193.950 ;
        RECT 463.950 190.950 466.050 193.050 ;
        RECT 451.950 164.850 453.750 165.750 ;
        RECT 454.950 163.950 457.050 166.050 ;
        RECT 458.250 164.850 459.750 165.750 ;
        RECT 460.950 163.950 463.050 166.050 ;
        RECT 460.950 161.850 463.050 162.750 ;
        RECT 460.950 142.950 463.050 145.050 ;
        RECT 449.400 140.400 453.450 141.450 ;
        RECT 439.950 125.250 441.750 126.150 ;
        RECT 442.950 124.950 445.050 127.050 ;
        RECT 446.400 124.050 447.450 139.950 ;
        RECT 448.950 136.950 451.050 139.050 ;
        RECT 439.950 121.950 442.050 124.050 ;
        RECT 443.250 122.850 445.050 123.750 ;
        RECT 445.950 121.950 448.050 124.050 ;
        RECT 436.950 109.950 439.050 112.050 ;
        RECT 440.400 109.050 441.450 121.950 ;
        RECT 433.950 106.950 436.050 109.050 ;
        RECT 439.950 106.950 442.050 109.050 ;
        RECT 449.400 108.450 450.450 136.950 ;
        RECT 452.400 124.050 453.450 140.400 ;
        RECT 457.950 139.950 460.050 142.050 ;
        RECT 458.400 130.050 459.450 139.950 ;
        RECT 454.950 128.250 457.050 129.150 ;
        RECT 457.950 127.950 460.050 130.050 ;
        RECT 461.400 127.050 462.450 142.950 ;
        RECT 464.400 139.050 465.450 190.950 ;
        RECT 470.400 187.050 471.450 196.950 ;
        RECT 485.400 196.050 486.450 199.950 ;
        RECT 472.950 194.850 475.050 195.750 ;
        RECT 475.950 194.250 478.050 195.150 ;
        RECT 478.950 194.850 480.750 195.750 ;
        RECT 481.950 193.950 484.050 196.050 ;
        RECT 484.950 193.950 487.050 196.050 ;
        RECT 482.400 193.050 483.450 193.950 ;
        RECT 475.950 190.950 478.050 193.050 ;
        RECT 481.950 190.950 484.050 193.050 ;
        RECT 469.950 184.950 472.050 187.050 ;
        RECT 472.950 184.950 475.050 187.050 ;
        RECT 469.950 172.950 472.050 175.050 ;
        RECT 473.400 174.450 474.450 184.950 ;
        RECT 476.400 178.050 477.450 190.950 ;
        RECT 481.950 187.950 484.050 190.050 ;
        RECT 475.950 175.950 478.050 178.050 ;
        RECT 473.400 173.400 477.450 174.450 ;
        RECT 470.400 166.050 471.450 172.950 ;
        RECT 472.950 169.950 475.050 172.050 ;
        RECT 473.400 166.050 474.450 169.950 ;
        RECT 476.400 169.050 477.450 173.400 ;
        RECT 478.950 172.950 481.050 175.050 ;
        RECT 475.950 166.950 478.050 169.050 ;
        RECT 469.950 163.950 472.050 166.050 ;
        RECT 472.950 163.950 475.050 166.050 ;
        RECT 476.250 164.250 478.050 165.150 ;
        RECT 466.950 161.850 468.750 162.750 ;
        RECT 469.950 160.950 472.050 163.050 ;
        RECT 473.250 161.850 474.750 162.750 ;
        RECT 475.950 160.950 478.050 163.050 ;
        RECT 469.950 158.850 472.050 159.750 ;
        RECT 476.400 145.050 477.450 160.950 ;
        RECT 479.400 145.050 480.450 172.950 ;
        RECT 482.400 154.050 483.450 187.950 ;
        RECT 488.400 187.050 489.450 226.950 ;
        RECT 493.950 214.950 496.050 217.050 ;
        RECT 494.400 199.050 495.450 214.950 ;
        RECT 497.400 202.050 498.450 263.400 ;
        RECT 499.950 262.950 502.050 265.050 ;
        RECT 508.950 262.950 511.050 265.050 ;
        RECT 508.950 259.950 511.050 262.050 ;
        RECT 499.950 256.950 502.050 259.050 ;
        RECT 500.400 208.050 501.450 256.950 ;
        RECT 509.400 253.050 510.450 259.950 ;
        RECT 508.950 250.950 511.050 253.050 ;
        RECT 512.400 247.050 513.450 265.950 ;
        RECT 515.400 256.050 516.450 271.950 ;
        RECT 521.400 271.050 522.450 292.950 ;
        RECT 530.400 274.050 531.450 334.950 ;
        RECT 554.400 325.050 555.450 367.950 ;
        RECT 557.400 337.050 558.450 367.950 ;
        RECT 568.800 367.800 570.900 369.900 ;
        RECT 590.400 367.050 591.450 386.400 ;
        RECT 593.250 370.050 594.450 388.950 ;
        RECT 596.250 376.350 597.450 388.950 ;
        RECT 595.950 374.250 598.050 376.350 ;
        RECT 596.250 370.050 597.450 374.250 ;
        RECT 599.250 370.050 600.450 388.950 ;
        RECT 604.950 377.850 607.050 378.750 ;
        RECT 592.950 367.950 595.050 370.050 ;
        RECT 595.950 367.950 598.050 370.050 ;
        RECT 598.950 367.950 601.050 370.050 ;
        RECT 589.950 364.950 592.050 367.050 ;
        RECT 595.950 364.950 598.050 367.050 ;
        RECT 559.950 355.950 562.050 358.050 ;
        RECT 560.400 349.050 561.450 355.950 ;
        RECT 577.950 352.950 580.050 355.050 ;
        RECT 559.950 346.950 562.050 349.050 ;
        RECT 568.950 346.950 571.050 349.050 ;
        RECT 571.950 346.950 574.050 349.050 ;
        RECT 560.400 340.050 561.450 346.950 ;
        RECT 569.400 346.050 570.450 346.950 ;
        RECT 562.950 343.950 565.050 346.050 ;
        RECT 566.250 344.250 567.750 345.150 ;
        RECT 568.950 343.950 571.050 346.050 ;
        RECT 562.950 341.850 564.750 342.750 ;
        RECT 565.950 340.950 568.050 343.050 ;
        RECT 569.250 341.850 571.050 342.750 ;
        RECT 559.950 337.950 562.050 340.050 ;
        RECT 556.950 334.950 559.050 337.050 ;
        RECT 556.950 325.950 559.050 328.050 ;
        RECT 553.950 322.950 556.050 325.050 ;
        RECT 541.950 316.950 544.050 319.050 ;
        RECT 532.950 313.950 535.050 316.050 ;
        RECT 535.950 313.950 538.050 316.050 ;
        RECT 533.400 313.050 534.450 313.950 ;
        RECT 532.950 310.950 535.050 313.050 ;
        RECT 536.400 310.050 537.450 313.950 ;
        RECT 542.400 313.050 543.450 316.950 ;
        RECT 538.950 311.250 540.750 312.150 ;
        RECT 541.950 310.950 544.050 313.050 ;
        RECT 547.950 311.250 550.050 312.150 ;
        RECT 532.950 308.850 535.050 309.750 ;
        RECT 535.950 307.950 538.050 310.050 ;
        RECT 538.950 307.950 541.050 310.050 ;
        RECT 542.250 308.850 544.050 309.750 ;
        RECT 547.950 307.950 550.050 310.050 ;
        RECT 535.950 298.950 538.050 301.050 ;
        RECT 532.950 289.950 535.050 292.050 ;
        RECT 529.950 271.950 532.050 274.050 ;
        RECT 517.950 269.250 519.750 270.150 ;
        RECT 520.950 268.950 523.050 271.050 ;
        RECT 524.250 269.250 525.750 270.150 ;
        RECT 526.950 268.950 529.050 271.050 ;
        RECT 530.250 269.250 532.050 270.150 ;
        RECT 517.950 265.950 520.050 268.050 ;
        RECT 521.250 266.850 522.750 267.750 ;
        RECT 523.950 265.950 526.050 268.050 ;
        RECT 527.250 266.850 528.750 267.750 ;
        RECT 529.950 265.950 532.050 268.050 ;
        RECT 517.950 264.450 520.050 265.050 ;
        RECT 520.950 264.450 523.050 265.050 ;
        RECT 517.950 263.400 523.050 264.450 ;
        RECT 517.950 262.950 520.050 263.400 ;
        RECT 520.950 262.950 523.050 263.400 ;
        RECT 524.400 261.450 525.450 265.950 ;
        RECT 529.950 262.950 532.050 265.050 ;
        RECT 524.400 260.400 528.450 261.450 ;
        RECT 523.950 256.950 526.050 259.050 ;
        RECT 514.950 253.950 517.050 256.050 ;
        RECT 514.950 250.950 517.050 253.050 ;
        RECT 511.950 244.950 514.050 247.050 ;
        RECT 505.950 241.950 508.050 244.050 ;
        RECT 511.950 243.450 514.050 244.050 ;
        RECT 515.400 243.450 516.450 250.950 ;
        RECT 511.950 242.400 516.450 243.450 ;
        RECT 511.950 241.950 514.050 242.400 ;
        RECT 502.950 239.250 505.050 240.150 ;
        RECT 505.950 239.850 508.050 240.750 ;
        RECT 508.950 238.950 511.050 241.050 ;
        RECT 514.950 238.950 517.050 241.050 ;
        RECT 502.950 235.950 505.050 238.050 ;
        RECT 503.400 235.050 504.450 235.950 ;
        RECT 502.950 232.950 505.050 235.050 ;
        RECT 505.950 232.950 508.050 235.050 ;
        RECT 503.400 229.050 504.450 232.950 ;
        RECT 502.950 226.950 505.050 229.050 ;
        RECT 506.400 217.050 507.450 232.950 ;
        RECT 509.400 220.050 510.450 238.950 ;
        RECT 515.400 238.050 516.450 238.950 ;
        RECT 511.950 236.250 513.750 237.150 ;
        RECT 514.950 235.950 517.050 238.050 ;
        RECT 518.250 236.250 520.050 237.150 ;
        RECT 520.950 235.950 523.050 238.050 ;
        RECT 511.950 232.950 514.050 235.050 ;
        RECT 515.250 233.850 516.750 234.750 ;
        RECT 517.950 232.950 520.050 235.050 ;
        RECT 512.400 232.050 513.450 232.950 ;
        RECT 511.950 229.950 514.050 232.050 ;
        RECT 508.950 217.950 511.050 220.050 ;
        RECT 505.950 214.950 508.050 217.050 ;
        RECT 505.950 211.950 508.050 214.050 ;
        RECT 499.950 205.950 502.050 208.050 ;
        RECT 502.950 205.950 505.050 208.050 ;
        RECT 496.950 199.950 499.050 202.050 ;
        RECT 499.950 200.250 502.050 201.150 ;
        RECT 490.950 197.250 492.750 198.150 ;
        RECT 493.950 196.950 496.050 199.050 ;
        RECT 497.250 197.250 498.750 198.150 ;
        RECT 499.950 196.950 502.050 199.050 ;
        RECT 490.950 193.950 493.050 196.050 ;
        RECT 494.250 194.850 495.750 195.750 ;
        RECT 496.950 193.950 499.050 196.050 ;
        RECT 490.950 190.950 493.050 193.050 ;
        RECT 487.950 184.950 490.050 187.050 ;
        RECT 484.950 181.950 487.050 184.050 ;
        RECT 481.950 151.950 484.050 154.050 ;
        RECT 475.950 142.950 478.050 145.050 ;
        RECT 478.950 142.950 481.050 145.050 ;
        RECT 478.950 139.950 481.050 142.050 ;
        RECT 463.950 136.950 466.050 139.050 ;
        RECT 479.400 133.050 480.450 139.950 ;
        RECT 481.950 136.950 484.050 139.050 ;
        RECT 478.950 130.950 481.050 133.050 ;
        RECT 478.950 128.250 481.050 129.150 ;
        RECT 454.950 124.950 457.050 127.050 ;
        RECT 458.250 125.250 459.750 126.150 ;
        RECT 460.950 124.950 463.050 127.050 ;
        RECT 464.250 125.250 466.050 126.150 ;
        RECT 466.950 124.950 469.050 127.050 ;
        RECT 469.950 125.250 471.750 126.150 ;
        RECT 472.950 124.950 475.050 127.050 ;
        RECT 476.250 125.250 477.750 126.150 ;
        RECT 478.950 124.950 481.050 127.050 ;
        RECT 451.950 121.950 454.050 124.050 ;
        RECT 446.400 107.400 450.450 108.450 ;
        RECT 434.400 94.050 435.450 106.950 ;
        RECT 440.400 97.050 441.450 106.950 ;
        RECT 442.950 103.950 445.050 106.050 ;
        RECT 439.950 94.950 442.050 97.050 ;
        RECT 433.950 91.950 436.050 94.050 ;
        RECT 437.250 92.250 439.050 93.150 ;
        RECT 439.950 91.950 442.050 94.050 ;
        RECT 427.950 89.850 429.750 90.750 ;
        RECT 430.950 88.950 433.050 91.050 ;
        RECT 434.250 89.850 435.750 90.750 ;
        RECT 436.950 88.950 439.050 91.050 ;
        RECT 440.400 88.050 441.450 91.950 ;
        RECT 443.400 91.050 444.450 103.950 ;
        RECT 442.950 88.950 445.050 91.050 ;
        RECT 430.950 86.850 433.050 87.750 ;
        RECT 439.950 85.950 442.050 88.050 ;
        RECT 442.950 76.950 445.050 79.050 ;
        RECT 433.950 73.950 436.050 76.050 ;
        RECT 430.950 67.950 433.050 70.050 ;
        RECT 431.400 58.050 432.450 67.950 ;
        RECT 434.400 61.050 435.450 73.950 ;
        RECT 439.950 64.950 442.050 67.050 ;
        RECT 433.950 58.950 436.050 61.050 ;
        RECT 418.950 56.250 421.050 57.150 ;
        RECT 421.950 55.950 424.050 58.050 ;
        RECT 424.950 55.950 427.050 58.050 ;
        RECT 430.950 55.950 433.050 58.050 ;
        RECT 434.250 56.250 435.750 57.150 ;
        RECT 436.950 55.950 439.050 58.050 ;
        RECT 440.400 55.050 441.450 64.950 ;
        RECT 443.400 61.050 444.450 76.950 ;
        RECT 446.400 70.050 447.450 107.400 ;
        RECT 455.400 100.050 456.450 124.950 ;
        RECT 457.950 121.950 460.050 124.050 ;
        RECT 461.250 122.850 462.750 123.750 ;
        RECT 463.950 121.950 466.050 124.050 ;
        RECT 458.400 106.050 459.450 121.950 ;
        RECT 463.950 118.950 466.050 121.050 ;
        RECT 457.950 103.950 460.050 106.050 ;
        RECT 454.950 97.950 457.050 100.050 ;
        RECT 455.400 97.050 456.450 97.950 ;
        RECT 448.950 94.950 451.050 97.050 ;
        RECT 452.250 95.250 453.750 96.150 ;
        RECT 454.950 94.950 457.050 97.050 ;
        RECT 464.400 94.050 465.450 118.950 ;
        RECT 467.400 115.050 468.450 124.950 ;
        RECT 482.400 124.050 483.450 136.950 ;
        RECT 485.400 133.050 486.450 181.950 ;
        RECT 491.400 169.050 492.450 190.950 ;
        RECT 497.400 187.050 498.450 193.950 ;
        RECT 500.400 193.050 501.450 196.950 ;
        RECT 499.950 190.950 502.050 193.050 ;
        RECT 496.950 184.950 499.050 187.050 ;
        RECT 503.400 175.050 504.450 205.950 ;
        RECT 506.400 196.050 507.450 211.950 ;
        RECT 508.950 207.450 511.050 208.050 ;
        RECT 511.950 207.450 514.050 208.050 ;
        RECT 508.950 206.400 514.050 207.450 ;
        RECT 508.950 205.950 511.050 206.400 ;
        RECT 511.950 205.950 514.050 206.400 ;
        RECT 517.950 205.950 520.050 208.050 ;
        RECT 511.950 203.250 514.050 204.150 ;
        RECT 518.400 202.050 519.450 205.950 ;
        RECT 521.400 205.050 522.450 235.950 ;
        RECT 524.400 217.050 525.450 256.950 ;
        RECT 527.400 256.050 528.450 260.400 ;
        RECT 526.950 253.950 529.050 256.050 ;
        RECT 530.400 253.050 531.450 262.950 ;
        RECT 533.400 253.050 534.450 289.950 ;
        RECT 536.400 256.050 537.450 298.950 ;
        RECT 548.400 289.050 549.450 307.950 ;
        RECT 547.950 286.950 550.050 289.050 ;
        RECT 541.950 274.950 544.050 277.050 ;
        RECT 542.400 271.050 543.450 274.950 ;
        RECT 554.400 274.050 555.450 322.950 ;
        RECT 557.400 274.050 558.450 325.950 ;
        RECT 566.400 322.050 567.450 340.950 ;
        RECT 572.400 325.050 573.450 346.950 ;
        RECT 574.950 343.950 577.050 346.050 ;
        RECT 575.400 339.450 576.450 343.950 ;
        RECT 578.400 342.450 579.450 352.950 ;
        RECT 580.950 344.250 583.050 345.150 ;
        RECT 580.950 342.450 583.050 343.050 ;
        RECT 578.400 341.400 583.050 342.450 ;
        RECT 580.950 340.950 583.050 341.400 ;
        RECT 584.250 341.250 585.750 342.150 ;
        RECT 586.950 340.950 589.050 343.050 ;
        RECT 590.250 341.250 592.050 342.150 ;
        RECT 592.950 340.950 595.050 343.050 ;
        RECT 575.400 338.400 579.450 339.450 ;
        RECT 574.950 331.950 577.050 334.050 ;
        RECT 571.950 322.950 574.050 325.050 ;
        RECT 565.950 319.950 568.050 322.050 ;
        RECT 566.400 316.050 567.450 319.950 ;
        RECT 565.950 313.950 568.050 316.050 ;
        RECT 571.950 313.950 574.050 316.050 ;
        RECT 562.950 311.250 565.050 312.150 ;
        RECT 568.950 310.950 571.050 313.050 ;
        RECT 572.250 311.850 574.050 312.750 ;
        RECT 562.950 307.950 565.050 310.050 ;
        RECT 565.950 307.950 568.050 310.050 ;
        RECT 568.950 308.850 571.050 309.750 ;
        RECT 563.400 307.050 564.450 307.950 ;
        RECT 562.950 304.950 565.050 307.050 ;
        RECT 559.950 283.950 562.050 286.050 ;
        RECT 547.950 271.950 550.050 274.050 ;
        RECT 553.950 271.950 556.050 274.050 ;
        RECT 556.950 271.950 559.050 274.050 ;
        RECT 538.950 268.950 541.050 271.050 ;
        RECT 541.950 268.950 544.050 271.050 ;
        RECT 538.950 266.850 541.050 267.750 ;
        RECT 541.950 266.250 544.050 267.150 ;
        RECT 541.950 264.450 544.050 265.050 ;
        RECT 539.400 263.400 544.050 264.450 ;
        RECT 535.950 253.950 538.050 256.050 ;
        RECT 529.950 250.950 532.050 253.050 ;
        RECT 532.950 250.950 535.050 253.050 ;
        RECT 539.400 247.050 540.450 263.400 ;
        RECT 541.950 262.950 544.050 263.400 ;
        RECT 541.950 259.950 544.050 262.050 ;
        RECT 542.400 256.050 543.450 259.950 ;
        RECT 548.400 259.050 549.450 271.950 ;
        RECT 560.400 271.050 561.450 283.950 ;
        RECT 550.950 269.250 552.750 270.150 ;
        RECT 553.950 268.950 556.050 271.050 ;
        RECT 557.250 269.250 558.750 270.150 ;
        RECT 559.950 268.950 562.050 271.050 ;
        RECT 563.250 269.250 565.050 270.150 ;
        RECT 566.400 268.050 567.450 307.950 ;
        RECT 575.400 286.050 576.450 331.950 ;
        RECT 574.950 283.950 577.050 286.050 ;
        RECT 578.400 283.050 579.450 338.400 ;
        RECT 583.950 337.950 586.050 340.050 ;
        RECT 587.250 338.850 588.750 339.750 ;
        RECT 589.950 337.950 592.050 340.050 ;
        RECT 580.950 334.950 583.050 337.050 ;
        RECT 581.400 292.050 582.450 334.950 ;
        RECT 586.950 331.950 589.050 334.050 ;
        RECT 587.400 310.050 588.450 331.950 ;
        RECT 590.400 328.050 591.450 337.950 ;
        RECT 593.400 337.050 594.450 340.950 ;
        RECT 592.950 334.950 595.050 337.050 ;
        RECT 596.400 334.050 597.450 364.950 ;
        RECT 604.950 352.950 607.050 355.050 ;
        RECT 601.950 349.950 604.050 352.050 ;
        RECT 602.400 343.050 603.450 349.950 ;
        RECT 598.950 341.250 600.750 342.150 ;
        RECT 601.950 340.950 604.050 343.050 ;
        RECT 598.950 337.950 601.050 340.050 ;
        RECT 602.250 338.850 604.050 339.750 ;
        RECT 595.950 331.950 598.050 334.050 ;
        RECT 589.950 325.950 592.050 328.050 ;
        RECT 598.950 322.950 601.050 325.050 ;
        RECT 595.950 319.950 598.050 322.050 ;
        RECT 596.400 316.050 597.450 319.950 ;
        RECT 595.950 313.950 598.050 316.050 ;
        RECT 595.950 310.950 598.050 313.050 ;
        RECT 583.950 308.250 585.750 309.150 ;
        RECT 586.950 307.950 589.050 310.050 ;
        RECT 590.250 308.250 592.050 309.150 ;
        RECT 583.950 304.950 586.050 307.050 ;
        RECT 587.250 305.850 588.750 306.750 ;
        RECT 589.950 304.950 592.050 307.050 ;
        RECT 590.400 304.050 591.450 304.950 ;
        RECT 583.950 301.950 586.050 304.050 ;
        RECT 589.950 301.950 592.050 304.050 ;
        RECT 580.950 289.950 583.050 292.050 ;
        RECT 574.950 280.950 577.050 283.050 ;
        RECT 577.950 280.950 580.050 283.050 ;
        RECT 568.950 274.950 571.050 277.050 ;
        RECT 569.400 271.050 570.450 274.950 ;
        RECT 575.400 271.050 576.450 280.950 ;
        RECT 568.950 268.950 571.050 271.050 ;
        RECT 574.950 268.950 577.050 271.050 ;
        RECT 578.250 269.250 580.050 270.150 ;
        RECT 584.400 268.050 585.450 301.950 ;
        RECT 596.400 280.050 597.450 310.950 ;
        RECT 599.400 304.050 600.450 322.950 ;
        RECT 605.400 312.450 606.450 352.950 ;
        RECT 608.400 346.050 609.450 397.950 ;
        RECT 611.400 388.050 612.450 418.950 ;
        RECT 617.400 414.450 618.450 419.400 ;
        RECT 619.950 416.250 622.050 417.150 ;
        RECT 619.950 414.450 622.050 415.050 ;
        RECT 617.400 413.400 622.050 414.450 ;
        RECT 619.950 412.950 622.050 413.400 ;
        RECT 623.250 413.250 624.750 414.150 ;
        RECT 625.950 412.950 628.050 415.050 ;
        RECT 629.250 413.250 631.050 414.150 ;
        RECT 616.950 409.950 619.050 412.050 ;
        RECT 619.950 411.450 622.050 412.050 ;
        RECT 622.950 411.450 625.050 412.050 ;
        RECT 619.950 410.400 625.050 411.450 ;
        RECT 626.250 410.850 627.750 411.750 ;
        RECT 619.950 409.950 622.050 410.400 ;
        RECT 622.950 409.950 625.050 410.400 ;
        RECT 628.950 409.950 631.050 412.050 ;
        RECT 610.950 385.950 613.050 388.050 ;
        RECT 610.950 380.250 613.050 381.150 ;
        RECT 610.950 376.950 613.050 379.050 ;
        RECT 607.950 343.950 610.050 346.050 ;
        RECT 607.950 340.950 610.050 343.050 ;
        RECT 607.950 338.850 610.050 339.750 ;
        RECT 617.400 328.050 618.450 409.950 ;
        RECT 619.950 397.950 622.050 400.050 ;
        RECT 620.400 388.050 621.450 397.950 ;
        RECT 629.400 397.050 630.450 409.950 ;
        RECT 632.400 403.050 633.450 451.950 ;
        RECT 637.950 436.950 640.050 439.050 ;
        RECT 634.950 418.950 637.050 421.050 ;
        RECT 635.400 418.050 636.450 418.950 ;
        RECT 634.950 415.950 637.050 418.050 ;
        RECT 635.400 415.050 636.450 415.950 ;
        RECT 634.950 412.950 637.050 415.050 ;
        RECT 634.950 410.850 637.050 411.750 ;
        RECT 634.950 406.950 637.050 409.050 ;
        RECT 631.950 400.950 634.050 403.050 ;
        RECT 628.950 394.950 631.050 397.050 ;
        RECT 628.950 388.950 631.050 391.050 ;
        RECT 619.950 385.950 622.050 388.050 ;
        RECT 625.950 385.950 628.050 388.050 ;
        RECT 619.950 383.850 622.050 384.750 ;
        RECT 622.950 383.250 625.050 384.150 ;
        RECT 622.950 381.450 625.050 382.050 ;
        RECT 626.400 381.450 627.450 385.950 ;
        RECT 622.950 380.400 627.450 381.450 ;
        RECT 622.950 379.950 625.050 380.400 ;
        RECT 629.400 361.050 630.450 388.950 ;
        RECT 635.400 385.050 636.450 406.950 ;
        RECT 638.400 394.050 639.450 436.950 ;
        RECT 637.950 391.950 640.050 394.050 ;
        RECT 641.400 391.050 642.450 514.950 ;
        RECT 653.400 487.050 654.450 520.950 ;
        RECT 689.400 505.050 690.450 526.950 ;
        RECT 688.950 502.950 691.050 505.050 ;
        RECT 673.800 497.100 675.900 499.200 ;
        RECT 674.550 493.350 675.750 497.100 ;
        RECT 676.950 494.850 679.050 496.950 ;
        RECT 673.950 491.250 676.050 493.350 ;
        RECT 664.950 488.250 667.050 489.150 ;
        RECT 643.950 484.950 646.050 487.050 ;
        RECT 652.950 486.450 655.050 487.050 ;
        RECT 650.400 485.400 655.050 486.450 ;
        RECT 643.950 482.850 646.050 483.750 ;
        RECT 646.950 482.250 649.050 483.150 ;
        RECT 646.950 480.450 649.050 481.050 ;
        RECT 650.400 480.450 651.450 485.400 ;
        RECT 652.950 484.950 655.050 485.400 ;
        RECT 664.950 484.950 667.050 487.050 ;
        RECT 652.950 482.850 655.050 483.750 ;
        RECT 646.950 479.400 651.450 480.450 ;
        RECT 646.950 478.950 649.050 479.400 ;
        RECT 661.950 478.950 664.050 481.050 ;
        RECT 652.950 460.950 655.050 463.050 ;
        RECT 646.950 457.950 649.050 460.050 ;
        RECT 647.400 457.050 648.450 457.950 ;
        RECT 653.400 457.050 654.450 460.950 ;
        RECT 643.950 454.950 646.050 457.050 ;
        RECT 646.950 454.950 649.050 457.050 ;
        RECT 650.250 455.250 651.750 456.150 ;
        RECT 652.950 454.950 655.050 457.050 ;
        RECT 655.950 454.950 658.050 457.050 ;
        RECT 644.400 400.050 645.450 454.950 ;
        RECT 656.400 454.050 657.450 454.950 ;
        RECT 646.950 452.850 648.750 453.750 ;
        RECT 649.950 451.950 652.050 454.050 ;
        RECT 653.250 452.850 654.750 453.750 ;
        RECT 655.950 451.950 658.050 454.050 ;
        RECT 646.950 416.250 649.050 417.150 ;
        RECT 646.950 412.950 649.050 415.050 ;
        RECT 643.950 397.950 646.050 400.050 ;
        RECT 647.400 391.050 648.450 412.950 ;
        RECT 650.400 409.050 651.450 451.950 ;
        RECT 655.950 449.850 658.050 450.750 ;
        RECT 662.400 448.050 663.450 478.950 ;
        RECT 674.550 477.600 675.750 491.250 ;
        RECT 677.250 477.600 678.450 494.850 ;
        RECT 684.900 494.400 687.000 496.500 ;
        RECT 688.950 494.400 691.050 496.500 ;
        RECT 679.950 491.250 682.050 493.350 ;
        RECT 680.400 477.600 681.600 491.250 ;
        RECT 685.350 485.550 686.550 494.400 ;
        RECT 689.550 488.250 690.750 494.400 ;
        RECT 692.400 493.050 693.450 604.950 ;
        RECT 694.950 599.250 697.050 600.150 ;
        RECT 698.400 598.050 699.450 640.950 ;
        RECT 700.950 634.950 703.050 637.050 ;
        RECT 701.400 631.050 702.450 634.950 ;
        RECT 712.950 632.250 715.050 633.150 ;
        RECT 700.950 628.950 703.050 631.050 ;
        RECT 712.950 630.450 715.050 631.050 ;
        RECT 716.400 630.450 717.450 667.950 ;
        RECT 721.950 664.950 724.050 667.050 ;
        RECT 725.250 665.850 726.750 666.750 ;
        RECT 727.950 664.950 730.050 667.050 ;
        RECT 722.400 658.050 723.450 664.950 ;
        RECT 728.400 661.050 729.450 664.950 ;
        RECT 727.950 658.950 730.050 661.050 ;
        RECT 721.950 655.950 724.050 658.050 ;
        RECT 721.800 641.100 723.900 643.200 ;
        RECT 722.550 637.350 723.750 641.100 ;
        RECT 724.950 638.850 727.050 640.950 ;
        RECT 721.950 635.250 724.050 637.350 ;
        RECT 712.950 629.400 717.450 630.450 ;
        RECT 712.950 628.950 715.050 629.400 ;
        RECT 700.950 626.850 703.050 627.750 ;
        RECT 703.950 610.950 706.050 613.050 ;
        RECT 694.950 595.950 697.050 598.050 ;
        RECT 697.950 595.950 700.050 598.050 ;
        RECT 695.400 589.050 696.450 595.950 ;
        RECT 704.400 589.050 705.450 610.950 ;
        RECT 713.400 610.050 714.450 628.950 ;
        RECT 716.400 628.050 717.450 629.400 ;
        RECT 718.950 628.950 721.050 631.050 ;
        RECT 715.950 625.950 718.050 628.050 ;
        RECT 719.400 613.050 720.450 628.950 ;
        RECT 722.550 621.600 723.750 635.250 ;
        RECT 725.250 621.600 726.450 638.850 ;
        RECT 732.900 638.400 735.000 640.500 ;
        RECT 736.950 638.400 739.050 640.500 ;
        RECT 727.950 635.250 730.050 637.350 ;
        RECT 728.400 621.600 729.600 635.250 ;
        RECT 733.350 629.550 734.550 638.400 ;
        RECT 737.550 632.250 738.750 638.400 ;
        RECT 736.950 630.150 739.050 632.250 ;
        RECT 740.400 631.050 741.450 674.400 ;
        RECT 752.400 664.050 753.450 691.950 ;
        RECT 754.950 676.950 757.050 679.050 ;
        RECT 751.950 661.950 754.050 664.050 ;
        RECT 745.950 640.950 748.050 643.050 ;
        RECT 748.950 640.950 751.050 643.050 ;
        RECT 751.950 640.950 754.050 643.050 ;
        RECT 732.750 627.450 734.850 629.550 ;
        RECT 733.350 621.600 734.550 627.450 ;
        RECT 737.550 621.600 738.750 630.150 ;
        RECT 739.950 628.950 742.050 631.050 ;
        RECT 739.950 626.250 742.050 627.150 ;
        RECT 739.950 622.950 742.050 625.050 ;
        RECT 746.250 622.050 747.450 640.950 ;
        RECT 749.250 636.750 750.450 640.950 ;
        RECT 748.950 634.650 751.050 636.750 ;
        RECT 749.250 622.050 750.450 634.650 ;
        RECT 752.250 622.050 753.450 640.950 ;
        RECT 755.400 622.050 756.450 676.950 ;
        RECT 757.950 671.250 760.050 672.150 ;
        RECT 757.950 667.950 760.050 670.050 ;
        RECT 757.950 632.250 760.050 633.150 ;
        RECT 721.950 619.500 724.050 621.600 ;
        RECT 724.950 619.500 727.050 621.600 ;
        RECT 727.950 619.500 730.050 621.600 ;
        RECT 732.750 619.500 734.850 621.600 ;
        RECT 736.950 619.500 739.050 621.600 ;
        RECT 745.950 619.950 748.050 622.050 ;
        RECT 748.950 619.950 751.050 622.050 ;
        RECT 751.950 619.950 754.050 622.050 ;
        RECT 754.950 619.950 757.050 622.050 ;
        RECT 733.950 613.950 736.050 616.050 ;
        RECT 718.950 610.950 721.050 613.050 ;
        RECT 706.950 607.950 709.050 610.050 ;
        RECT 712.950 607.950 715.050 610.050 ;
        RECT 707.400 598.050 708.450 607.950 ;
        RECT 715.950 605.400 718.050 607.500 ;
        RECT 718.950 605.400 721.050 607.500 ;
        RECT 721.950 605.400 724.050 607.500 ;
        RECT 726.750 605.400 728.850 607.500 ;
        RECT 730.950 605.400 733.050 607.500 ;
        RECT 712.950 601.950 715.050 604.050 ;
        RECT 706.950 595.950 709.050 598.050 ;
        RECT 706.950 593.850 709.050 594.750 ;
        RECT 713.400 592.050 714.450 601.950 ;
        RECT 712.950 589.950 715.050 592.050 ;
        RECT 716.550 591.750 717.750 605.400 ;
        RECT 715.950 589.650 718.050 591.750 ;
        RECT 694.950 586.950 697.050 589.050 ;
        RECT 703.950 586.950 706.050 589.050 ;
        RECT 716.550 585.900 717.750 589.650 ;
        RECT 719.250 588.150 720.450 605.400 ;
        RECT 722.400 591.750 723.600 605.400 ;
        RECT 727.350 599.550 728.550 605.400 ;
        RECT 726.750 597.450 728.850 599.550 ;
        RECT 721.950 589.650 724.050 591.750 ;
        RECT 727.350 588.600 728.550 597.450 ;
        RECT 731.550 596.850 732.750 605.400 ;
        RECT 734.400 604.050 735.450 613.950 ;
        RECT 736.950 610.950 739.050 613.050 ;
        RECT 733.950 601.950 736.050 604.050 ;
        RECT 733.950 599.850 736.050 600.750 ;
        RECT 730.950 594.750 733.050 596.850 ;
        RECT 731.550 588.600 732.750 594.750 ;
        RECT 718.950 586.050 721.050 588.150 ;
        RECT 726.900 586.500 729.000 588.600 ;
        RECT 730.950 586.500 733.050 588.600 ;
        RECT 715.800 583.800 717.900 585.900 ;
        RECT 737.400 568.050 738.450 610.950 ;
        RECT 748.950 607.950 751.050 610.050 ;
        RECT 739.950 604.950 742.050 607.050 ;
        RECT 742.950 604.950 745.050 607.050 ;
        RECT 745.950 604.950 748.050 607.050 ;
        RECT 740.250 586.050 741.450 604.950 ;
        RECT 743.250 592.350 744.450 604.950 ;
        RECT 742.950 590.250 745.050 592.350 ;
        RECT 743.250 586.050 744.450 590.250 ;
        RECT 746.250 586.050 747.450 604.950 ;
        RECT 739.950 583.950 742.050 586.050 ;
        RECT 742.950 583.950 745.050 586.050 ;
        RECT 745.950 583.950 748.050 586.050 ;
        RECT 730.950 565.950 733.050 568.050 ;
        RECT 736.950 565.950 739.050 568.050 ;
        RECT 731.400 562.050 732.450 565.950 ;
        RECT 749.400 565.050 750.450 607.950 ;
        RECT 761.400 600.450 762.450 691.950 ;
        RECT 766.950 688.950 769.050 691.050 ;
        RECT 763.950 685.950 766.050 688.050 ;
        RECT 764.400 667.050 765.450 685.950 ;
        RECT 767.400 670.050 768.450 688.950 ;
        RECT 770.400 679.050 771.450 706.950 ;
        RECT 773.400 703.050 774.450 757.950 ;
        RECT 778.950 754.950 781.050 757.050 ;
        RECT 784.950 754.950 787.050 757.050 ;
        RECT 775.950 743.250 778.050 744.150 ;
        RECT 775.950 741.450 778.050 742.050 ;
        RECT 779.400 741.450 780.450 754.950 ;
        RECT 781.950 742.950 784.050 745.050 ;
        RECT 775.950 740.400 780.450 741.450 ;
        RECT 775.950 739.950 778.050 740.400 ;
        RECT 772.950 700.950 775.050 703.050 ;
        RECT 772.950 698.850 775.050 699.750 ;
        RECT 772.950 694.950 775.050 697.050 ;
        RECT 769.950 676.950 772.050 679.050 ;
        RECT 769.950 673.950 772.050 676.050 ;
        RECT 770.400 670.050 771.450 673.950 ;
        RECT 773.400 673.050 774.450 694.950 ;
        RECT 776.400 676.050 777.450 739.950 ;
        RECT 778.950 736.950 781.050 739.050 ;
        RECT 779.400 700.050 780.450 736.950 ;
        RECT 778.950 697.950 781.050 700.050 ;
        RECT 775.950 673.950 778.050 676.050 ;
        RECT 772.950 670.950 775.050 673.050 ;
        RECT 776.250 671.250 777.750 672.150 ;
        RECT 778.950 670.950 781.050 673.050 ;
        RECT 766.950 667.950 769.050 670.050 ;
        RECT 769.950 667.950 772.050 670.050 ;
        RECT 773.250 668.850 774.750 669.750 ;
        RECT 775.950 667.950 778.050 670.050 ;
        RECT 779.250 668.850 781.050 669.750 ;
        RECT 776.400 667.050 777.450 667.950 ;
        RECT 763.950 664.950 766.050 667.050 ;
        RECT 769.950 665.850 772.050 666.750 ;
        RECT 775.950 664.950 778.050 667.050 ;
        RECT 764.400 634.050 765.450 664.950 ;
        RECT 769.950 655.950 772.050 658.050 ;
        RECT 763.950 631.950 766.050 634.050 ;
        RECT 763.950 629.850 766.050 630.750 ;
        RECT 770.400 613.050 771.450 655.950 ;
        RECT 772.950 646.950 775.050 649.050 ;
        RECT 773.400 637.050 774.450 646.950 ;
        RECT 776.400 640.050 777.450 664.950 ;
        RECT 775.950 637.950 778.050 640.050 ;
        RECT 772.950 634.950 775.050 637.050 ;
        RECT 773.400 631.050 774.450 634.950 ;
        RECT 772.950 628.950 775.050 631.050 ;
        RECT 772.950 626.850 775.050 627.750 ;
        RECT 772.950 613.950 775.050 616.050 ;
        RECT 769.950 610.950 772.050 613.050 ;
        RECT 766.950 607.950 769.050 610.050 ;
        RECT 761.400 599.400 765.450 600.450 ;
        RECT 757.950 596.250 760.050 597.150 ;
        RECT 760.950 595.950 763.050 598.050 ;
        RECT 751.950 593.850 754.050 594.750 ;
        RECT 757.950 594.450 760.050 595.050 ;
        RECT 761.400 594.450 762.450 595.950 ;
        RECT 757.950 593.400 762.450 594.450 ;
        RECT 757.950 592.950 760.050 593.400 ;
        RECT 757.950 589.950 760.050 592.050 ;
        RECT 754.950 571.950 757.050 574.050 ;
        RECT 736.950 562.950 739.050 565.050 ;
        RECT 739.950 562.950 742.050 565.050 ;
        RECT 748.950 562.950 751.050 565.050 ;
        RECT 737.400 562.050 738.450 562.950 ;
        RECT 730.950 559.950 733.050 562.050 ;
        RECT 734.250 560.250 735.750 561.150 ;
        RECT 736.950 559.950 739.050 562.050 ;
        RECT 697.950 558.450 700.050 559.050 ;
        RECT 695.400 557.400 700.050 558.450 ;
        RECT 730.950 557.850 732.750 558.750 ;
        RECT 695.400 525.450 696.450 557.400 ;
        RECT 697.950 556.950 700.050 557.400 ;
        RECT 733.950 556.950 736.050 559.050 ;
        RECT 737.250 557.850 739.050 558.750 ;
        RECT 734.400 556.050 735.450 556.950 ;
        RECT 697.950 554.850 700.050 555.750 ;
        RECT 718.950 554.850 721.050 555.750 ;
        RECT 733.950 553.950 736.050 556.050 ;
        RECT 706.950 533.400 709.050 535.500 ;
        RECT 709.950 533.400 712.050 535.500 ;
        RECT 712.950 533.400 715.050 535.500 ;
        RECT 717.750 533.400 719.850 535.500 ;
        RECT 721.950 533.400 724.050 535.500 ;
        RECT 697.950 525.450 700.050 526.050 ;
        RECT 695.400 524.400 700.050 525.450 ;
        RECT 691.950 490.950 694.050 493.050 ;
        RECT 688.950 486.150 691.050 488.250 ;
        RECT 695.400 487.050 696.450 524.400 ;
        RECT 697.950 523.950 700.050 524.400 ;
        RECT 697.950 521.850 700.050 522.750 ;
        RECT 707.550 519.750 708.750 533.400 ;
        RECT 706.950 517.650 709.050 519.750 ;
        RECT 707.550 513.900 708.750 517.650 ;
        RECT 710.250 516.150 711.450 533.400 ;
        RECT 713.400 519.750 714.600 533.400 ;
        RECT 718.350 527.550 719.550 533.400 ;
        RECT 717.750 525.450 719.850 527.550 ;
        RECT 712.950 517.650 715.050 519.750 ;
        RECT 718.350 516.600 719.550 525.450 ;
        RECT 722.550 524.850 723.750 533.400 ;
        RECT 730.950 532.950 733.050 535.050 ;
        RECT 733.950 532.950 736.050 535.050 ;
        RECT 736.950 532.950 739.050 535.050 ;
        RECT 724.950 529.950 727.050 532.050 ;
        RECT 724.950 527.850 727.050 528.750 ;
        RECT 721.950 522.750 724.050 524.850 ;
        RECT 722.550 516.600 723.750 522.750 ;
        RECT 709.950 514.050 712.050 516.150 ;
        RECT 717.900 514.500 720.000 516.600 ;
        RECT 721.950 514.500 724.050 516.600 ;
        RECT 731.250 514.050 732.450 532.950 ;
        RECT 734.250 520.350 735.450 532.950 ;
        RECT 733.950 518.250 736.050 520.350 ;
        RECT 734.250 514.050 735.450 518.250 ;
        RECT 737.250 514.050 738.450 532.950 ;
        RECT 706.800 511.800 708.900 513.900 ;
        RECT 730.950 511.950 733.050 514.050 ;
        RECT 733.950 511.950 736.050 514.050 ;
        RECT 736.950 511.950 739.050 514.050 ;
        RECT 730.950 508.950 733.050 511.050 ;
        RECT 706.950 502.950 709.050 505.050 ;
        RECT 697.950 496.950 700.050 499.050 ;
        RECT 700.950 496.950 703.050 499.050 ;
        RECT 703.950 496.950 706.050 499.050 ;
        RECT 684.750 483.450 686.850 485.550 ;
        RECT 685.350 477.600 686.550 483.450 ;
        RECT 689.550 477.600 690.750 486.150 ;
        RECT 694.950 484.950 697.050 487.050 ;
        RECT 691.950 482.250 694.050 483.150 ;
        RECT 691.950 478.950 694.050 481.050 ;
        RECT 698.250 478.050 699.450 496.950 ;
        RECT 701.250 492.750 702.450 496.950 ;
        RECT 700.950 490.650 703.050 492.750 ;
        RECT 701.250 478.050 702.450 490.650 ;
        RECT 704.250 478.050 705.450 496.950 ;
        RECT 673.950 475.500 676.050 477.600 ;
        RECT 676.950 475.500 679.050 477.600 ;
        RECT 679.950 475.500 682.050 477.600 ;
        RECT 684.750 475.500 686.850 477.600 ;
        RECT 688.950 475.500 691.050 477.600 ;
        RECT 697.950 475.950 700.050 478.050 ;
        RECT 700.950 475.950 703.050 478.050 ;
        RECT 703.950 475.950 706.050 478.050 ;
        RECT 697.950 469.950 700.050 472.050 ;
        RECT 667.950 466.950 670.050 469.050 ;
        RECT 673.950 466.950 676.050 469.050 ;
        RECT 668.400 457.050 669.450 466.950 ;
        RECT 674.400 457.050 675.450 466.950 ;
        RECT 667.950 454.950 670.050 457.050 ;
        RECT 671.250 455.250 672.750 456.150 ;
        RECT 673.950 454.950 676.050 457.050 ;
        RECT 676.950 454.950 679.050 457.050 ;
        RECT 679.950 454.950 682.050 457.050 ;
        RECT 685.950 456.450 688.050 457.050 ;
        RECT 683.400 455.400 688.050 456.450 ;
        RECT 677.400 454.050 678.450 454.950 ;
        RECT 667.950 452.850 669.750 453.750 ;
        RECT 670.950 451.950 673.050 454.050 ;
        RECT 674.250 452.850 675.750 453.750 ;
        RECT 676.950 451.950 679.050 454.050 ;
        RECT 676.950 449.850 679.050 450.750 ;
        RECT 661.950 445.950 664.050 448.050 ;
        RECT 680.400 429.450 681.450 454.950 ;
        RECT 683.400 430.050 684.450 455.400 ;
        RECT 685.950 454.950 688.050 455.400 ;
        RECT 689.250 455.250 690.750 456.150 ;
        RECT 691.950 454.950 694.050 457.050 ;
        RECT 694.950 454.950 697.050 457.050 ;
        RECT 695.400 454.050 696.450 454.950 ;
        RECT 685.950 452.850 687.750 453.750 ;
        RECT 688.950 451.950 691.050 454.050 ;
        RECT 692.250 452.850 693.750 453.750 ;
        RECT 694.950 451.950 697.050 454.050 ;
        RECT 694.950 449.850 697.050 450.750 ;
        RECT 677.400 428.400 681.450 429.450 ;
        RECT 655.800 425.100 657.900 427.200 ;
        RECT 656.550 421.350 657.750 425.100 ;
        RECT 658.950 422.850 661.050 424.950 ;
        RECT 655.950 419.250 658.050 421.350 ;
        RECT 649.950 406.950 652.050 409.050 ;
        RECT 656.550 405.600 657.750 419.250 ;
        RECT 659.250 405.600 660.450 422.850 ;
        RECT 666.900 422.400 669.000 424.500 ;
        RECT 670.950 422.400 673.050 424.500 ;
        RECT 661.950 419.250 664.050 421.350 ;
        RECT 662.400 405.600 663.600 419.250 ;
        RECT 667.350 413.550 668.550 422.400 ;
        RECT 671.550 416.250 672.750 422.400 ;
        RECT 670.950 414.150 673.050 416.250 ;
        RECT 666.750 411.450 668.850 413.550 ;
        RECT 667.350 405.600 668.550 411.450 ;
        RECT 671.550 405.600 672.750 414.150 ;
        RECT 673.950 410.250 676.050 411.150 ;
        RECT 673.950 408.450 676.050 409.050 ;
        RECT 677.400 408.450 678.450 428.400 ;
        RECT 682.950 427.950 685.050 430.050 ;
        RECT 679.950 424.950 682.050 427.050 ;
        RECT 682.950 424.950 685.050 427.050 ;
        RECT 685.950 424.950 688.050 427.050 ;
        RECT 673.950 407.400 678.450 408.450 ;
        RECT 673.950 406.950 676.050 407.400 ;
        RECT 680.250 406.050 681.450 424.950 ;
        RECT 683.250 420.750 684.450 424.950 ;
        RECT 682.950 418.650 685.050 420.750 ;
        RECT 683.250 406.050 684.450 418.650 ;
        RECT 686.250 406.050 687.450 424.950 ;
        RECT 698.400 418.050 699.450 469.950 ;
        RECT 700.950 457.950 703.050 460.050 ;
        RECT 691.950 416.250 694.050 417.150 ;
        RECT 697.950 415.950 700.050 418.050 ;
        RECT 697.950 413.850 700.050 414.750 ;
        RECT 655.950 403.500 658.050 405.600 ;
        RECT 658.950 403.500 661.050 405.600 ;
        RECT 661.950 403.500 664.050 405.600 ;
        RECT 666.750 403.500 668.850 405.600 ;
        RECT 670.950 403.500 673.050 405.600 ;
        RECT 679.950 403.950 682.050 406.050 ;
        RECT 682.950 403.950 685.050 406.050 ;
        RECT 685.950 403.950 688.050 406.050 ;
        RECT 694.950 403.950 697.050 406.050 ;
        RECT 676.950 400.950 679.050 403.050 ;
        RECT 661.950 397.950 664.050 400.050 ;
        RECT 664.950 397.950 667.050 400.050 ;
        RECT 640.950 388.950 643.050 391.050 ;
        RECT 646.950 388.950 649.050 391.050 ;
        RECT 640.950 385.950 643.050 388.050 ;
        RECT 655.950 385.950 658.050 388.050 ;
        RECT 634.950 382.950 637.050 385.050 ;
        RECT 638.250 383.250 640.050 384.150 ;
        RECT 640.950 383.850 643.050 384.750 ;
        RECT 643.950 383.250 646.050 384.150 ;
        RECT 646.950 382.950 649.050 385.050 ;
        RECT 652.950 382.950 655.050 385.050 ;
        RECT 634.950 380.850 636.750 381.750 ;
        RECT 637.950 379.950 640.050 382.050 ;
        RECT 643.950 379.950 646.050 382.050 ;
        RECT 644.400 367.050 645.450 379.950 ;
        RECT 647.400 369.450 648.450 382.950 ;
        RECT 653.400 382.050 654.450 382.950 ;
        RECT 649.950 380.250 651.750 381.150 ;
        RECT 652.950 379.950 655.050 382.050 ;
        RECT 656.400 379.050 657.450 385.950 ;
        RECT 658.950 382.950 661.050 385.050 ;
        RECT 659.400 382.050 660.450 382.950 ;
        RECT 658.950 379.950 661.050 382.050 ;
        RECT 649.950 376.950 652.050 379.050 ;
        RECT 653.250 377.850 654.750 378.750 ;
        RECT 655.950 376.950 658.050 379.050 ;
        RECT 659.250 377.850 661.050 378.750 ;
        RECT 650.400 373.050 651.450 376.950 ;
        RECT 655.950 374.850 658.050 375.750 ;
        RECT 662.400 373.050 663.450 397.950 ;
        RECT 665.400 385.050 666.450 397.950 ;
        RECT 670.950 394.950 673.050 397.050 ;
        RECT 671.400 388.050 672.450 394.950 ;
        RECT 670.950 387.450 673.050 388.050 ;
        RECT 670.950 386.400 675.450 387.450 ;
        RECT 670.950 385.950 673.050 386.400 ;
        RECT 664.950 382.950 667.050 385.050 ;
        RECT 667.950 383.250 670.050 384.150 ;
        RECT 670.950 383.850 673.050 384.750 ;
        RECT 665.400 381.450 666.450 382.950 ;
        RECT 674.400 382.050 675.450 386.400 ;
        RECT 677.400 385.050 678.450 400.950 ;
        RECT 682.950 391.950 685.050 394.050 ;
        RECT 683.400 385.050 684.450 391.950 ;
        RECT 695.400 385.050 696.450 403.950 ;
        RECT 701.400 399.450 702.450 457.950 ;
        RECT 703.950 454.950 706.050 457.050 ;
        RECT 707.400 456.450 708.450 502.950 ;
        RECT 715.950 489.450 718.050 490.050 ;
        RECT 709.950 488.250 712.050 489.150 ;
        RECT 715.950 488.400 720.450 489.450 ;
        RECT 715.950 487.950 718.050 488.400 ;
        RECT 715.950 485.850 718.050 486.750 ;
        RECT 719.400 484.050 720.450 488.400 ;
        RECT 731.400 487.050 732.450 508.950 ;
        RECT 736.950 505.950 739.050 508.050 ;
        RECT 724.950 484.950 727.050 487.050 ;
        RECT 727.950 485.250 729.750 486.150 ;
        RECT 730.950 484.950 733.050 487.050 ;
        RECT 733.950 485.250 736.050 486.150 ;
        RECT 718.950 481.950 721.050 484.050 ;
        RECT 719.400 472.050 720.450 481.950 ;
        RECT 718.950 469.950 721.050 472.050 ;
        RECT 725.400 460.050 726.450 484.950 ;
        RECT 727.950 481.950 730.050 484.050 ;
        RECT 731.250 482.850 733.050 483.750 ;
        RECT 733.950 483.450 736.050 484.050 ;
        RECT 737.400 483.450 738.450 505.950 ;
        RECT 740.400 490.050 741.450 562.950 ;
        RECT 745.950 559.950 748.050 562.050 ;
        RECT 751.950 560.250 754.050 561.150 ;
        RECT 746.400 559.050 747.450 559.950 ;
        RECT 742.950 557.250 744.750 558.150 ;
        RECT 745.950 556.950 748.050 559.050 ;
        RECT 749.250 557.250 750.750 558.150 ;
        RECT 751.950 556.950 754.050 559.050 ;
        RECT 752.400 556.050 753.450 556.950 ;
        RECT 742.950 553.950 745.050 556.050 ;
        RECT 746.250 554.850 747.750 555.750 ;
        RECT 748.950 553.950 751.050 556.050 ;
        RECT 751.950 553.950 754.050 556.050 ;
        RECT 749.400 547.050 750.450 553.950 ;
        RECT 751.950 550.950 754.050 553.050 ;
        RECT 748.950 544.950 751.050 547.050 ;
        RECT 748.950 524.250 751.050 525.150 ;
        RECT 742.950 521.850 745.050 522.750 ;
        RECT 748.950 520.950 751.050 523.050 ;
        RECT 749.400 501.450 750.450 520.950 ;
        RECT 752.400 508.050 753.450 550.950 ;
        RECT 755.400 550.050 756.450 571.950 ;
        RECT 758.400 553.050 759.450 589.950 ;
        RECT 764.400 568.050 765.450 599.400 ;
        RECT 767.400 592.050 768.450 607.950 ;
        RECT 769.950 598.950 772.050 601.050 ;
        RECT 769.950 596.850 772.050 597.750 ;
        RECT 766.950 589.950 769.050 592.050 ;
        RECT 767.400 582.450 768.450 589.950 ;
        RECT 767.400 581.400 771.450 582.450 ;
        RECT 763.950 565.950 766.050 568.050 ;
        RECT 764.400 564.450 765.450 565.950 ;
        RECT 761.400 563.400 765.450 564.450 ;
        RECT 761.400 558.450 762.450 563.400 ;
        RECT 763.950 560.250 766.050 561.150 ;
        RECT 770.400 559.050 771.450 581.400 ;
        RECT 773.400 561.450 774.450 613.950 ;
        RECT 776.400 610.050 777.450 637.950 ;
        RECT 778.950 628.950 781.050 631.050 ;
        RECT 779.400 616.050 780.450 628.950 ;
        RECT 778.950 613.950 781.050 616.050 ;
        RECT 775.950 607.950 778.050 610.050 ;
        RECT 778.950 604.950 781.050 607.050 ;
        RECT 775.950 598.950 778.050 601.050 ;
        RECT 775.950 596.850 778.050 597.750 ;
        RECT 779.400 562.050 780.450 604.950 ;
        RECT 773.400 560.400 777.450 561.450 ;
        RECT 763.950 558.450 766.050 559.050 ;
        RECT 761.400 557.400 766.050 558.450 ;
        RECT 763.950 556.950 766.050 557.400 ;
        RECT 767.250 557.250 768.750 558.150 ;
        RECT 769.950 556.950 772.050 559.050 ;
        RECT 773.250 557.250 775.050 558.150 ;
        RECT 766.950 553.950 769.050 556.050 ;
        RECT 770.250 554.850 771.750 555.750 ;
        RECT 772.950 553.950 775.050 556.050 ;
        RECT 757.950 550.950 760.050 553.050 ;
        RECT 754.950 547.950 757.050 550.050 ;
        RECT 755.400 523.050 756.450 547.950 ;
        RECT 757.950 529.950 760.050 532.050 ;
        RECT 758.400 529.050 759.450 529.950 ;
        RECT 757.950 526.950 760.050 529.050 ;
        RECT 761.250 527.250 762.750 528.150 ;
        RECT 763.950 526.950 766.050 529.050 ;
        RECT 776.400 528.450 777.450 560.400 ;
        RECT 778.950 559.950 781.050 562.050 ;
        RECT 778.950 556.950 781.050 559.050 ;
        RECT 778.950 554.850 781.050 555.750 ;
        RECT 782.400 546.450 783.450 742.950 ;
        RECT 785.400 709.050 786.450 754.950 ;
        RECT 791.400 748.050 792.450 772.950 ;
        RECT 806.400 757.050 807.450 772.950 ;
        RECT 812.400 772.050 813.450 811.950 ;
        RECT 821.400 808.050 822.450 817.950 ;
        RECT 826.950 815.250 829.050 816.150 ;
        RECT 829.950 815.850 832.050 816.750 ;
        RECT 839.400 814.050 840.450 817.950 ;
        RECT 826.950 811.950 829.050 814.050 ;
        RECT 835.950 812.250 837.750 813.150 ;
        RECT 838.950 811.950 841.050 814.050 ;
        RECT 842.250 812.250 844.050 813.150 ;
        RECT 835.950 808.950 838.050 811.050 ;
        RECT 839.250 809.850 840.750 810.750 ;
        RECT 841.950 808.950 844.050 811.050 ;
        RECT 820.950 805.950 823.050 808.050 ;
        RECT 836.400 784.050 837.450 808.950 ;
        RECT 829.950 781.950 832.050 784.050 ;
        RECT 835.950 781.950 838.050 784.050 ;
        RECT 820.950 773.250 823.050 774.150 ;
        RECT 826.950 773.250 829.050 774.150 ;
        RECT 811.950 769.950 814.050 772.050 ;
        RECT 820.950 769.950 823.050 772.050 ;
        RECT 824.250 770.250 825.750 771.150 ;
        RECT 826.950 769.950 829.050 772.050 ;
        RECT 830.400 771.450 831.450 781.950 ;
        RECT 832.950 773.250 835.050 774.150 ;
        RECT 838.950 773.250 841.050 774.150 ;
        RECT 832.950 771.450 835.050 772.050 ;
        RECT 830.400 770.400 835.050 771.450 ;
        RECT 838.950 771.450 841.050 772.050 ;
        RECT 842.400 771.450 843.450 808.950 ;
        RECT 847.950 772.950 850.050 775.050 ;
        RECT 851.250 773.250 853.050 774.150 ;
        RECT 853.950 772.950 856.050 775.050 ;
        RECT 832.950 769.950 835.050 770.400 ;
        RECT 836.250 770.250 837.750 771.150 ;
        RECT 838.950 770.400 843.450 771.450 ;
        RECT 847.950 770.850 849.750 771.750 ;
        RECT 838.950 769.950 841.050 770.400 ;
        RECT 850.950 769.950 853.050 772.050 ;
        RECT 827.400 769.050 828.450 769.950 ;
        RECT 823.950 766.950 826.050 769.050 ;
        RECT 826.950 766.950 829.050 769.050 ;
        RECT 835.950 766.950 838.050 769.050 ;
        RECT 805.950 754.950 808.050 757.050 ;
        RECT 796.950 749.400 799.050 751.500 ;
        RECT 799.950 749.400 802.050 751.500 ;
        RECT 802.950 749.400 805.050 751.500 ;
        RECT 807.750 749.400 809.850 751.500 ;
        RECT 811.950 749.400 814.050 751.500 ;
        RECT 851.400 751.050 852.450 769.950 ;
        RECT 790.950 745.950 793.050 748.050 ;
        RECT 787.950 741.450 790.050 742.050 ;
        RECT 787.950 740.400 792.450 741.450 ;
        RECT 787.950 739.950 790.050 740.400 ;
        RECT 787.950 737.850 790.050 738.750 ;
        RECT 791.400 735.450 792.450 740.400 ;
        RECT 797.550 735.750 798.750 749.400 ;
        RECT 788.400 734.400 792.450 735.450 ;
        RECT 784.950 706.950 787.050 709.050 ;
        RECT 784.950 704.250 787.050 705.150 ;
        RECT 784.950 702.450 787.050 703.050 ;
        RECT 788.400 702.450 789.450 734.400 ;
        RECT 796.950 733.650 799.050 735.750 ;
        RECT 797.550 729.900 798.750 733.650 ;
        RECT 800.250 732.150 801.450 749.400 ;
        RECT 803.400 735.750 804.600 749.400 ;
        RECT 808.350 743.550 809.550 749.400 ;
        RECT 807.750 741.450 809.850 743.550 ;
        RECT 802.950 733.650 805.050 735.750 ;
        RECT 808.350 732.600 809.550 741.450 ;
        RECT 812.550 740.850 813.750 749.400 ;
        RECT 820.950 748.950 823.050 751.050 ;
        RECT 823.950 748.950 826.050 751.050 ;
        RECT 826.950 748.950 829.050 751.050 ;
        RECT 829.950 748.950 832.050 751.050 ;
        RECT 850.950 748.950 853.050 751.050 ;
        RECT 814.950 747.450 817.050 748.050 ;
        RECT 814.950 746.400 819.450 747.450 ;
        RECT 814.950 745.950 817.050 746.400 ;
        RECT 814.950 743.850 817.050 744.750 ;
        RECT 811.950 738.750 814.050 740.850 ;
        RECT 818.400 739.050 819.450 746.400 ;
        RECT 812.550 732.600 813.750 738.750 ;
        RECT 817.950 736.950 820.050 739.050 ;
        RECT 799.950 730.050 802.050 732.150 ;
        RECT 807.900 730.500 810.000 732.600 ;
        RECT 811.950 730.500 814.050 732.600 ;
        RECT 821.250 730.050 822.450 748.950 ;
        RECT 824.250 736.350 825.450 748.950 ;
        RECT 823.950 734.250 826.050 736.350 ;
        RECT 824.250 730.050 825.450 734.250 ;
        RECT 827.250 730.050 828.450 748.950 ;
        RECT 796.800 727.800 798.900 729.900 ;
        RECT 820.950 727.950 823.050 730.050 ;
        RECT 823.950 727.950 826.050 730.050 ;
        RECT 826.950 727.950 829.050 730.050 ;
        RECT 826.950 724.950 829.050 727.050 ;
        RECT 793.800 713.100 795.900 715.200 ;
        RECT 794.550 709.350 795.750 713.100 ;
        RECT 817.950 712.950 820.050 715.050 ;
        RECT 820.950 712.950 823.050 715.050 ;
        RECT 823.950 712.950 826.050 715.050 ;
        RECT 796.950 710.850 799.050 712.950 ;
        RECT 790.950 706.950 793.050 709.050 ;
        RECT 793.950 707.250 796.050 709.350 ;
        RECT 784.950 701.400 789.450 702.450 ;
        RECT 784.950 700.950 787.050 701.400 ;
        RECT 785.400 691.050 786.450 700.950 ;
        RECT 784.950 688.950 787.050 691.050 ;
        RECT 784.950 676.950 787.050 679.050 ;
        RECT 785.400 676.050 786.450 676.950 ;
        RECT 791.400 676.050 792.450 706.950 ;
        RECT 794.550 693.600 795.750 707.250 ;
        RECT 797.250 693.600 798.450 710.850 ;
        RECT 804.900 710.400 807.000 712.500 ;
        RECT 808.950 710.400 811.050 712.500 ;
        RECT 799.950 707.250 802.050 709.350 ;
        RECT 800.400 693.600 801.600 707.250 ;
        RECT 805.350 701.550 806.550 710.400 ;
        RECT 809.550 704.250 810.750 710.400 ;
        RECT 814.950 706.950 817.050 709.050 ;
        RECT 808.950 702.150 811.050 704.250 ;
        RECT 804.750 699.450 806.850 701.550 ;
        RECT 805.350 693.600 806.550 699.450 ;
        RECT 809.550 693.600 810.750 702.150 ;
        RECT 811.950 698.250 814.050 699.150 ;
        RECT 811.950 694.950 814.050 697.050 ;
        RECT 793.950 691.500 796.050 693.600 ;
        RECT 796.950 691.500 799.050 693.600 ;
        RECT 799.950 691.500 802.050 693.600 ;
        RECT 804.750 691.500 806.850 693.600 ;
        RECT 808.950 691.500 811.050 693.600 ;
        RECT 812.400 691.050 813.450 694.950 ;
        RECT 811.950 688.950 814.050 691.050 ;
        RECT 815.400 678.450 816.450 706.950 ;
        RECT 818.250 694.050 819.450 712.950 ;
        RECT 821.250 708.750 822.450 712.950 ;
        RECT 820.950 706.650 823.050 708.750 ;
        RECT 821.250 694.050 822.450 706.650 ;
        RECT 824.250 694.050 825.450 712.950 ;
        RECT 817.950 691.950 820.050 694.050 ;
        RECT 820.950 691.950 823.050 694.050 ;
        RECT 823.950 691.950 826.050 694.050 ;
        RECT 820.950 688.950 823.050 691.050 ;
        RECT 812.400 677.400 816.450 678.450 ;
        RECT 784.950 673.950 787.050 676.050 ;
        RECT 790.950 673.950 793.050 676.050 ;
        RECT 796.950 673.950 799.050 676.050 ;
        RECT 808.950 673.950 811.050 676.050 ;
        RECT 784.950 671.850 787.050 672.750 ;
        RECT 787.950 671.250 790.050 672.150 ;
        RECT 787.950 667.950 790.050 670.050 ;
        RECT 788.400 658.050 789.450 667.950 ;
        RECT 791.400 661.050 792.450 673.950 ;
        RECT 796.950 671.850 798.750 672.750 ;
        RECT 799.950 672.450 802.050 673.050 ;
        RECT 799.950 671.400 804.450 672.450 ;
        RECT 799.950 670.950 802.050 671.400 ;
        RECT 803.400 670.050 804.450 671.400 ;
        RECT 805.950 671.250 808.050 672.150 ;
        RECT 799.950 668.850 802.050 669.750 ;
        RECT 802.950 667.950 805.050 670.050 ;
        RECT 805.950 669.450 808.050 670.050 ;
        RECT 809.400 669.450 810.450 673.950 ;
        RECT 805.950 668.400 810.450 669.450 ;
        RECT 805.950 667.950 808.050 668.400 ;
        RECT 790.950 658.950 793.050 661.050 ;
        RECT 787.950 655.950 790.050 658.050 ;
        RECT 787.950 652.950 790.050 655.050 ;
        RECT 784.950 632.250 787.050 633.150 ;
        RECT 784.950 628.950 787.050 631.050 ;
        RECT 785.400 628.050 786.450 628.950 ;
        RECT 784.950 625.950 787.050 628.050 ;
        RECT 788.400 619.050 789.450 652.950 ;
        RECT 793.800 641.100 795.900 643.200 ;
        RECT 794.550 637.350 795.750 641.100 ;
        RECT 796.950 638.850 799.050 640.950 ;
        RECT 793.950 635.250 796.050 637.350 ;
        RECT 790.950 631.950 793.050 634.050 ;
        RECT 787.950 616.950 790.050 619.050 ;
        RECT 787.950 613.950 790.050 616.050 ;
        RECT 784.950 610.950 787.050 613.050 ;
        RECT 785.400 604.050 786.450 610.950 ;
        RECT 784.950 601.950 787.050 604.050 ;
        RECT 788.400 601.050 789.450 613.950 ;
        RECT 791.400 601.050 792.450 631.950 ;
        RECT 794.550 621.600 795.750 635.250 ;
        RECT 797.250 621.600 798.450 638.850 ;
        RECT 804.900 638.400 807.000 640.500 ;
        RECT 808.950 638.400 811.050 640.500 ;
        RECT 799.950 635.250 802.050 637.350 ;
        RECT 800.400 621.600 801.600 635.250 ;
        RECT 805.350 629.550 806.550 638.400 ;
        RECT 809.550 632.250 810.750 638.400 ;
        RECT 808.950 630.150 811.050 632.250 ;
        RECT 812.400 631.050 813.450 677.400 ;
        RECT 814.950 673.950 817.050 676.050 ;
        RECT 815.400 673.050 816.450 673.950 ;
        RECT 821.400 673.050 822.450 688.950 ;
        RECT 823.950 673.950 826.050 676.050 ;
        RECT 814.950 670.950 817.050 673.050 ;
        RECT 818.250 671.250 819.750 672.150 ;
        RECT 820.950 670.950 823.050 673.050 ;
        RECT 824.400 670.050 825.450 673.950 ;
        RECT 814.950 668.850 816.750 669.750 ;
        RECT 817.950 667.950 820.050 670.050 ;
        RECT 821.250 668.850 822.750 669.750 ;
        RECT 823.950 667.950 826.050 670.050 ;
        RECT 818.400 664.050 819.450 667.950 ;
        RECT 823.950 665.850 826.050 666.750 ;
        RECT 814.950 661.950 817.050 664.050 ;
        RECT 817.950 661.950 820.050 664.050 ;
        RECT 804.750 627.450 806.850 629.550 ;
        RECT 805.350 621.600 806.550 627.450 ;
        RECT 809.550 621.600 810.750 630.150 ;
        RECT 811.950 628.950 814.050 631.050 ;
        RECT 811.950 626.250 814.050 627.150 ;
        RECT 811.950 622.950 814.050 625.050 ;
        RECT 793.950 619.500 796.050 621.600 ;
        RECT 796.950 619.500 799.050 621.600 ;
        RECT 799.950 619.500 802.050 621.600 ;
        RECT 804.750 619.500 806.850 621.600 ;
        RECT 808.950 619.500 811.050 621.600 ;
        RECT 812.400 619.050 813.450 622.950 ;
        RECT 811.950 616.950 814.050 619.050 ;
        RECT 799.950 613.950 802.050 616.050 ;
        RECT 811.950 613.950 814.050 616.050 ;
        RECT 796.950 610.950 799.050 613.050 ;
        RECT 784.950 599.850 786.750 600.750 ;
        RECT 787.950 598.950 790.050 601.050 ;
        RECT 790.950 598.950 793.050 601.050 ;
        RECT 793.950 599.250 796.050 600.150 ;
        RECT 787.950 596.850 790.050 597.750 ;
        RECT 784.950 565.950 787.050 568.050 ;
        RECT 785.400 559.050 786.450 565.950 ;
        RECT 791.400 565.050 792.450 598.950 ;
        RECT 793.950 595.950 796.050 598.050 ;
        RECT 793.950 592.950 796.050 595.050 ;
        RECT 787.950 562.950 790.050 565.050 ;
        RECT 790.950 562.950 793.050 565.050 ;
        RECT 784.950 556.950 787.050 559.050 ;
        RECT 788.400 558.450 789.450 562.950 ;
        RECT 790.950 560.250 793.050 561.150 ;
        RECT 790.950 558.450 793.050 559.050 ;
        RECT 788.400 557.400 793.050 558.450 ;
        RECT 790.950 556.950 793.050 557.400 ;
        RECT 782.400 545.400 786.450 546.450 ;
        RECT 778.950 529.950 781.050 532.050 ;
        RECT 773.400 527.400 777.450 528.450 ;
        RECT 757.950 524.850 759.750 525.750 ;
        RECT 760.950 523.950 763.050 526.050 ;
        RECT 764.250 524.850 765.750 525.750 ;
        RECT 766.950 525.450 769.050 526.050 ;
        RECT 766.950 524.400 771.450 525.450 ;
        RECT 766.950 523.950 769.050 524.400 ;
        RECT 761.400 523.050 762.450 523.950 ;
        RECT 754.950 520.950 757.050 523.050 ;
        RECT 760.950 520.950 763.050 523.050 ;
        RECT 766.950 521.850 769.050 522.750 ;
        RECT 754.950 517.950 757.050 520.050 ;
        RECT 755.400 513.450 756.450 517.950 ;
        RECT 755.400 512.400 759.450 513.450 ;
        RECT 751.950 505.950 754.050 508.050 ;
        RECT 746.400 500.400 750.450 501.450 ;
        RECT 746.400 496.050 747.450 500.400 ;
        RECT 745.950 493.950 748.050 496.050 ;
        RECT 739.950 487.950 742.050 490.050 ;
        RECT 739.950 485.250 742.050 486.150 ;
        RECT 746.400 484.050 747.450 493.950 ;
        RECT 748.950 485.250 751.050 486.150 ;
        RECT 754.950 485.250 757.050 486.150 ;
        RECT 733.950 482.400 738.450 483.450 ;
        RECT 733.950 481.950 736.050 482.400 ;
        RECT 728.400 481.050 729.450 481.950 ;
        RECT 727.950 478.950 730.050 481.050 ;
        RECT 728.400 478.050 729.450 478.950 ;
        RECT 727.950 475.950 730.050 478.050 ;
        RECT 724.950 457.950 727.050 460.050 ;
        RECT 733.950 457.950 736.050 460.050 ;
        RECT 707.400 455.400 711.450 456.450 ;
        RECT 704.400 450.450 705.450 454.950 ;
        RECT 710.400 454.050 711.450 455.400 ;
        RECT 724.950 455.250 727.050 456.150 ;
        RECT 730.950 454.950 733.050 457.050 ;
        RECT 734.250 455.850 736.050 456.750 ;
        RECT 706.950 452.250 708.750 453.150 ;
        RECT 709.950 451.950 712.050 454.050 ;
        RECT 715.950 453.450 718.050 454.050 ;
        RECT 715.950 452.400 720.450 453.450 ;
        RECT 715.950 451.950 718.050 452.400 ;
        RECT 706.950 450.450 709.050 451.050 ;
        RECT 704.400 449.400 709.050 450.450 ;
        RECT 710.250 449.850 711.750 450.750 ;
        RECT 706.950 448.950 709.050 449.400 ;
        RECT 712.950 448.950 715.050 451.050 ;
        RECT 716.250 449.850 718.050 450.750 ;
        RECT 719.400 448.050 720.450 452.400 ;
        RECT 724.950 451.950 727.050 454.050 ;
        RECT 727.950 451.950 730.050 454.050 ;
        RECT 730.950 452.850 733.050 453.750 ;
        RECT 733.950 451.950 736.050 454.050 ;
        RECT 725.400 451.050 726.450 451.950 ;
        RECT 724.950 448.950 727.050 451.050 ;
        RECT 712.950 446.850 715.050 447.750 ;
        RECT 718.950 445.950 721.050 448.050 ;
        RECT 718.950 442.950 721.050 445.050 ;
        RECT 703.950 418.950 706.050 421.050 ;
        RECT 704.400 415.050 705.450 418.950 ;
        RECT 706.950 415.950 709.050 418.050 ;
        RECT 710.250 416.250 711.750 417.150 ;
        RECT 712.950 415.950 715.050 418.050 ;
        RECT 715.950 415.950 718.050 418.050 ;
        RECT 703.950 412.950 706.050 415.050 ;
        RECT 706.950 413.850 708.750 414.750 ;
        RECT 709.950 412.950 712.050 415.050 ;
        RECT 713.250 413.850 715.050 414.750 ;
        RECT 710.400 412.050 711.450 412.950 ;
        RECT 709.950 409.950 712.050 412.050 ;
        RECT 701.400 398.400 705.450 399.450 ;
        RECT 700.950 394.950 703.050 397.050 ;
        RECT 701.400 385.050 702.450 394.950 ;
        RECT 676.950 384.450 679.050 385.050 ;
        RECT 676.950 383.400 681.450 384.450 ;
        RECT 676.950 382.950 679.050 383.400 ;
        RECT 667.950 381.450 670.050 382.050 ;
        RECT 665.400 380.400 670.050 381.450 ;
        RECT 667.950 379.950 670.050 380.400 ;
        RECT 673.950 379.950 676.050 382.050 ;
        RECT 676.950 380.850 679.050 381.750 ;
        RECT 674.400 373.050 675.450 379.950 ;
        RECT 680.400 379.050 681.450 383.400 ;
        RECT 682.950 382.950 685.050 385.050 ;
        RECT 685.950 382.950 688.050 385.050 ;
        RECT 691.950 382.950 694.050 385.050 ;
        RECT 694.950 382.950 697.050 385.050 ;
        RECT 698.250 383.250 699.750 384.150 ;
        RECT 700.950 382.950 703.050 385.050 ;
        RECT 682.950 380.850 685.050 381.750 ;
        RECT 679.950 376.950 682.050 379.050 ;
        RECT 649.950 370.950 652.050 373.050 ;
        RECT 661.950 370.950 664.050 373.050 ;
        RECT 673.950 370.950 676.050 373.050 ;
        RECT 647.400 368.400 651.450 369.450 ;
        RECT 643.950 364.950 646.050 367.050 ;
        RECT 628.950 358.950 631.050 361.050 ;
        RECT 628.800 353.100 630.900 355.200 ;
        RECT 629.550 349.350 630.750 353.100 ;
        RECT 631.950 350.850 634.050 352.950 ;
        RECT 628.950 347.250 631.050 349.350 ;
        RECT 619.950 344.250 622.050 345.150 ;
        RECT 625.950 343.950 628.050 346.050 ;
        RECT 619.950 340.950 622.050 343.050 ;
        RECT 619.950 337.950 622.050 340.050 ;
        RECT 616.950 325.950 619.050 328.050 ;
        RECT 616.950 319.950 619.050 322.050 ;
        RECT 610.950 316.950 613.050 319.050 ;
        RECT 611.400 316.050 612.450 316.950 ;
        RECT 610.950 313.950 613.050 316.050 ;
        RECT 607.950 312.450 610.050 313.050 ;
        RECT 601.950 311.250 604.050 312.150 ;
        RECT 605.400 311.400 610.050 312.450 ;
        RECT 611.250 311.850 613.050 312.750 ;
        RECT 601.950 307.950 604.050 310.050 ;
        RECT 602.400 307.050 603.450 307.950 ;
        RECT 605.400 307.050 606.450 311.400 ;
        RECT 607.950 310.950 610.050 311.400 ;
        RECT 617.400 310.050 618.450 319.950 ;
        RECT 620.400 313.050 621.450 337.950 ;
        RECT 626.400 321.450 627.450 343.950 ;
        RECT 629.550 333.600 630.750 347.250 ;
        RECT 632.250 333.600 633.450 350.850 ;
        RECT 639.900 350.400 642.000 352.500 ;
        RECT 643.950 350.400 646.050 352.500 ;
        RECT 634.950 347.250 637.050 349.350 ;
        RECT 635.400 333.600 636.600 347.250 ;
        RECT 640.350 341.550 641.550 350.400 ;
        RECT 644.550 344.250 645.750 350.400 ;
        RECT 643.950 342.150 646.050 344.250 ;
        RECT 639.750 339.450 641.850 341.550 ;
        RECT 640.350 333.600 641.550 339.450 ;
        RECT 644.550 333.600 645.750 342.150 ;
        RECT 646.950 338.250 649.050 339.150 ;
        RECT 646.950 334.950 649.050 337.050 ;
        RECT 628.950 331.500 631.050 333.600 ;
        RECT 631.950 331.500 634.050 333.600 ;
        RECT 634.950 331.500 637.050 333.600 ;
        RECT 639.750 331.500 641.850 333.600 ;
        RECT 643.950 331.500 646.050 333.600 ;
        RECT 647.400 331.050 648.450 334.950 ;
        RECT 646.950 328.950 649.050 331.050 ;
        RECT 650.400 328.050 651.450 368.400 ;
        RECT 673.950 367.950 676.050 370.050 ;
        RECT 661.950 364.950 664.050 367.050 ;
        RECT 652.950 352.950 655.050 355.050 ;
        RECT 655.950 352.950 658.050 355.050 ;
        RECT 658.950 352.950 661.050 355.050 ;
        RECT 653.250 334.050 654.450 352.950 ;
        RECT 656.250 348.750 657.450 352.950 ;
        RECT 655.950 346.650 658.050 348.750 ;
        RECT 656.250 334.050 657.450 346.650 ;
        RECT 659.250 334.050 660.450 352.950 ;
        RECT 652.950 331.950 655.050 334.050 ;
        RECT 655.950 331.950 658.050 334.050 ;
        RECT 658.950 331.950 661.050 334.050 ;
        RECT 652.950 328.950 655.050 331.050 ;
        RECT 631.950 325.950 634.050 328.050 ;
        RECT 649.950 325.950 652.050 328.050 ;
        RECT 626.400 320.400 630.450 321.450 ;
        RECT 625.950 316.950 628.050 319.050 ;
        RECT 622.950 313.950 625.050 316.050 ;
        RECT 619.950 310.950 622.050 313.050 ;
        RECT 607.950 308.850 610.050 309.750 ;
        RECT 613.950 308.250 615.750 309.150 ;
        RECT 616.950 307.950 619.050 310.050 ;
        RECT 620.250 308.250 622.050 309.150 ;
        RECT 601.950 304.950 604.050 307.050 ;
        RECT 604.950 304.950 607.050 307.050 ;
        RECT 613.950 304.950 616.050 307.050 ;
        RECT 617.250 305.850 618.750 306.750 ;
        RECT 619.950 304.950 622.050 307.050 ;
        RECT 598.950 301.950 601.050 304.050 ;
        RECT 601.950 295.950 604.050 298.050 ;
        RECT 602.400 289.050 603.450 295.950 ;
        RECT 598.950 286.950 601.050 289.050 ;
        RECT 601.950 286.950 604.050 289.050 ;
        RECT 595.950 277.950 598.050 280.050 ;
        RECT 599.400 274.050 600.450 286.950 ;
        RECT 598.950 271.950 601.050 274.050 ;
        RECT 601.950 272.250 604.050 273.150 ;
        RECT 586.950 268.950 589.050 271.050 ;
        RECT 592.950 269.250 594.750 270.150 ;
        RECT 595.950 268.950 598.050 271.050 ;
        RECT 599.250 269.250 600.750 270.150 ;
        RECT 601.950 268.950 604.050 271.050 ;
        RECT 550.950 265.950 553.050 268.050 ;
        RECT 554.250 266.850 555.750 267.750 ;
        RECT 556.950 265.950 559.050 268.050 ;
        RECT 560.250 266.850 561.750 267.750 ;
        RECT 562.950 265.950 565.050 268.050 ;
        RECT 565.950 265.950 568.050 268.050 ;
        RECT 568.950 266.850 571.050 267.750 ;
        RECT 571.950 266.250 574.050 267.150 ;
        RECT 574.950 266.850 576.750 267.750 ;
        RECT 577.950 265.950 580.050 268.050 ;
        RECT 583.950 265.950 586.050 268.050 ;
        RECT 586.950 266.850 589.050 267.750 ;
        RECT 589.950 266.250 592.050 267.150 ;
        RECT 592.950 265.950 595.050 268.050 ;
        RECT 596.250 266.850 597.750 267.750 ;
        RECT 598.950 265.950 601.050 268.050 ;
        RECT 601.950 265.950 604.050 268.050 ;
        RECT 551.400 265.050 552.450 265.950 ;
        RECT 550.950 262.950 553.050 265.050 ;
        RECT 553.950 262.950 556.050 265.050 ;
        RECT 550.950 259.950 553.050 262.050 ;
        RECT 547.950 256.950 550.050 259.050 ;
        RECT 541.950 253.950 544.050 256.050 ;
        RECT 547.950 253.950 550.050 256.050 ;
        RECT 542.400 253.050 543.450 253.950 ;
        RECT 541.950 250.950 544.050 253.050 ;
        RECT 538.950 244.950 541.050 247.050 ;
        RECT 541.950 244.950 544.050 247.050 ;
        RECT 529.950 241.950 532.050 244.050 ;
        RECT 542.400 243.450 543.450 244.950 ;
        RECT 536.400 242.400 543.450 243.450 ;
        RECT 536.400 241.050 537.450 242.400 ;
        RECT 548.400 241.050 549.450 253.950 ;
        RECT 526.950 239.250 529.050 240.150 ;
        RECT 529.950 239.850 532.050 240.750 ;
        RECT 532.950 239.250 534.750 240.150 ;
        RECT 535.950 238.950 538.050 241.050 ;
        RECT 541.950 238.950 544.050 241.050 ;
        RECT 547.950 238.950 550.050 241.050 ;
        RECT 526.950 235.950 529.050 238.050 ;
        RECT 529.950 235.950 532.050 238.050 ;
        RECT 532.950 235.950 535.050 238.050 ;
        RECT 536.250 236.850 538.050 237.750 ;
        RECT 527.400 235.050 528.450 235.950 ;
        RECT 526.950 232.950 529.050 235.050 ;
        RECT 530.400 232.050 531.450 235.950 ;
        RECT 542.400 232.050 543.450 238.950 ;
        RECT 551.400 238.050 552.450 259.950 ;
        RECT 554.400 252.450 555.450 262.950 ;
        RECT 557.400 262.050 558.450 265.950 ;
        RECT 593.400 265.050 594.450 265.950 ;
        RECT 559.950 262.950 562.050 265.050 ;
        RECT 562.950 262.950 565.050 265.050 ;
        RECT 565.950 262.950 568.050 265.050 ;
        RECT 571.950 262.950 574.050 265.050 ;
        RECT 589.950 262.950 592.050 265.050 ;
        RECT 592.950 262.950 595.050 265.050 ;
        RECT 598.950 262.950 601.050 265.050 ;
        RECT 556.950 259.950 559.050 262.050 ;
        RECT 560.400 259.050 561.450 262.950 ;
        RECT 559.950 256.950 562.050 259.050 ;
        RECT 554.400 251.400 558.450 252.450 ;
        RECT 547.950 236.250 549.750 237.150 ;
        RECT 550.950 235.950 553.050 238.050 ;
        RECT 554.250 236.250 556.050 237.150 ;
        RECT 547.950 232.950 550.050 235.050 ;
        RECT 551.250 233.850 552.750 234.750 ;
        RECT 553.950 232.950 556.050 235.050 ;
        RECT 526.950 229.950 529.050 232.050 ;
        RECT 529.950 229.950 532.050 232.050 ;
        RECT 541.950 229.950 544.050 232.050 ;
        RECT 523.950 214.950 526.050 217.050 ;
        RECT 523.950 205.950 526.050 208.050 ;
        RECT 520.950 202.950 523.050 205.050 ;
        RECT 508.950 200.250 510.750 201.150 ;
        RECT 511.950 199.950 514.050 202.050 ;
        RECT 515.250 200.250 516.750 201.150 ;
        RECT 517.950 199.950 520.050 202.050 ;
        RECT 520.950 199.950 523.050 202.050 ;
        RECT 508.950 196.950 511.050 199.050 ;
        RECT 505.950 193.950 508.050 196.050 ;
        RECT 505.950 190.950 508.050 193.050 ;
        RECT 506.400 178.050 507.450 190.950 ;
        RECT 509.400 184.050 510.450 196.950 ;
        RECT 512.400 196.050 513.450 199.950 ;
        RECT 514.950 196.950 517.050 199.050 ;
        RECT 518.250 197.850 520.050 198.750 ;
        RECT 515.400 196.050 516.450 196.950 ;
        RECT 511.950 193.950 514.050 196.050 ;
        RECT 514.950 193.950 517.050 196.050 ;
        RECT 511.950 190.950 514.050 193.050 ;
        RECT 514.950 190.950 517.050 193.050 ;
        RECT 508.950 181.950 511.050 184.050 ;
        RECT 505.950 175.950 508.050 178.050 ;
        RECT 506.400 175.050 507.450 175.950 ;
        RECT 502.950 172.950 505.050 175.050 ;
        RECT 505.950 172.950 508.050 175.050 ;
        RECT 496.950 169.950 499.050 172.050 ;
        RECT 497.400 169.050 498.450 169.950 ;
        RECT 512.400 169.050 513.450 190.950 ;
        RECT 515.400 169.050 516.450 190.950 ;
        RECT 521.400 190.050 522.450 199.950 ;
        RECT 520.950 187.950 523.050 190.050 ;
        RECT 520.950 175.950 523.050 178.050 ;
        RECT 487.950 166.950 490.050 169.050 ;
        RECT 490.950 166.950 493.050 169.050 ;
        RECT 496.950 166.950 499.050 169.050 ;
        RECT 499.950 166.950 502.050 169.050 ;
        RECT 505.950 166.950 508.050 169.050 ;
        RECT 509.250 167.250 510.750 168.150 ;
        RECT 511.950 166.950 514.050 169.050 ;
        RECT 514.950 166.950 517.050 169.050 ;
        RECT 487.950 164.850 490.050 165.750 ;
        RECT 493.950 164.250 496.050 165.150 ;
        RECT 496.950 164.850 499.050 165.750 ;
        RECT 487.950 160.950 490.050 163.050 ;
        RECT 493.950 162.450 496.050 163.050 ;
        RECT 491.400 161.400 496.050 162.450 ;
        RECT 488.400 157.050 489.450 160.950 ;
        RECT 487.950 154.950 490.050 157.050 ;
        RECT 491.400 151.050 492.450 161.400 ;
        RECT 493.950 160.950 496.050 161.400 ;
        RECT 493.950 154.950 496.050 157.050 ;
        RECT 490.950 148.950 493.050 151.050 ;
        RECT 484.950 130.950 487.050 133.050 ;
        RECT 484.950 127.950 487.050 130.050 ;
        RECT 487.950 128.250 490.050 129.150 ;
        RECT 469.950 121.950 472.050 124.050 ;
        RECT 473.250 122.850 474.750 123.750 ;
        RECT 475.950 121.950 478.050 124.050 ;
        RECT 478.950 121.950 481.050 124.050 ;
        RECT 481.950 121.950 484.050 124.050 ;
        RECT 470.400 121.050 471.450 121.950 ;
        RECT 476.400 121.050 477.450 121.950 ;
        RECT 469.950 118.950 472.050 121.050 ;
        RECT 472.950 118.950 475.050 121.050 ;
        RECT 475.950 118.950 478.050 121.050 ;
        RECT 466.950 112.950 469.050 115.050 ;
        RECT 467.400 97.050 468.450 112.950 ;
        RECT 473.400 97.050 474.450 118.950 ;
        RECT 466.950 94.950 469.050 97.050 ;
        RECT 470.250 95.250 471.750 96.150 ;
        RECT 472.950 94.950 475.050 97.050 ;
        RECT 475.950 94.950 478.050 97.050 ;
        RECT 476.400 94.050 477.450 94.950 ;
        RECT 448.950 92.850 450.750 93.750 ;
        RECT 451.950 91.950 454.050 94.050 ;
        RECT 455.250 92.850 456.750 93.750 ;
        RECT 460.950 91.950 463.050 94.050 ;
        RECT 463.950 91.950 466.050 94.050 ;
        RECT 466.950 92.850 468.750 93.750 ;
        RECT 469.950 91.950 472.050 94.050 ;
        RECT 473.250 92.850 474.750 93.750 ;
        RECT 475.950 91.950 478.050 94.050 ;
        RECT 451.950 88.950 454.050 91.050 ;
        RECT 457.950 89.850 460.050 90.750 ;
        RECT 445.950 67.950 448.050 70.050 ;
        RECT 442.950 58.950 445.050 61.050 ;
        RECT 397.950 53.250 399.750 54.150 ;
        RECT 400.950 52.950 403.050 55.050 ;
        RECT 404.250 53.250 405.750 54.150 ;
        RECT 406.950 52.950 409.050 55.050 ;
        RECT 409.950 52.950 412.050 55.050 ;
        RECT 412.950 52.950 415.050 55.050 ;
        RECT 418.950 52.950 421.050 55.050 ;
        RECT 422.250 53.250 423.750 54.150 ;
        RECT 424.950 52.950 427.050 55.050 ;
        RECT 428.250 53.250 430.050 54.150 ;
        RECT 430.950 53.850 432.750 54.750 ;
        RECT 433.950 52.950 436.050 55.050 ;
        RECT 437.250 53.850 439.050 54.750 ;
        RECT 439.950 52.950 442.050 55.050 ;
        RECT 407.400 52.050 408.450 52.950 ;
        RECT 382.950 50.850 385.050 51.750 ;
        RECT 388.950 49.950 391.050 52.050 ;
        RECT 394.950 51.450 397.050 52.050 ;
        RECT 397.950 51.450 400.050 52.050 ;
        RECT 392.250 50.250 394.050 51.150 ;
        RECT 394.950 50.400 400.050 51.450 ;
        RECT 401.250 50.850 402.750 51.750 ;
        RECT 394.950 49.950 397.050 50.400 ;
        RECT 397.950 49.950 400.050 50.400 ;
        RECT 403.950 49.950 406.050 52.050 ;
        RECT 406.950 49.950 409.050 52.050 ;
        RECT 373.950 46.950 376.050 49.050 ;
        RECT 379.950 46.950 382.050 49.050 ;
        RECT 391.950 46.950 394.050 49.050 ;
        RECT 385.950 43.950 388.050 46.050 ;
        RECT 370.950 31.950 373.050 34.050 ;
        RECT 382.950 31.950 385.050 34.050 ;
        RECT 371.400 28.050 372.450 31.950 ;
        RECT 376.950 28.950 379.050 31.050 ;
        RECT 377.400 28.050 378.450 28.950 ;
        RECT 370.950 25.950 373.050 28.050 ;
        RECT 376.950 25.950 379.050 28.050 ;
        RECT 358.950 22.950 361.050 25.050 ;
        RECT 362.250 23.850 363.750 24.750 ;
        RECT 364.950 22.950 367.050 25.050 ;
        RECT 358.950 20.850 361.050 21.750 ;
        RECT 364.950 20.850 367.050 21.750 ;
        RECT 371.400 21.450 372.450 25.950 ;
        RECT 383.400 25.050 384.450 31.950 ;
        RECT 373.950 23.250 376.050 24.150 ;
        RECT 376.950 23.850 379.050 24.750 ;
        RECT 379.950 23.250 381.750 24.150 ;
        RECT 382.950 22.950 385.050 25.050 ;
        RECT 373.950 21.450 376.050 22.050 ;
        RECT 371.400 20.400 376.050 21.450 ;
        RECT 373.950 19.950 376.050 20.400 ;
        RECT 379.950 19.950 382.050 22.050 ;
        RECT 383.250 20.850 385.050 21.750 ;
        RECT 386.400 21.450 387.450 43.950 ;
        RECT 392.400 40.050 393.450 46.950 ;
        RECT 391.950 37.950 394.050 40.050 ;
        RECT 397.950 37.950 400.050 40.050 ;
        RECT 394.950 31.950 397.050 34.050 ;
        RECT 388.950 23.250 390.750 24.150 ;
        RECT 391.950 22.950 394.050 25.050 ;
        RECT 388.950 21.450 391.050 22.050 ;
        RECT 386.400 20.400 391.050 21.450 ;
        RECT 392.250 20.850 394.050 21.750 ;
        RECT 388.950 19.950 391.050 20.400 ;
        RECT 343.950 16.950 346.050 17.400 ;
        RECT 349.950 17.400 354.450 18.450 ;
        RECT 349.950 16.950 352.050 17.400 ;
        RECT 380.400 16.050 381.450 19.950 ;
        RECT 395.400 16.050 396.450 31.950 ;
        RECT 398.400 22.050 399.450 37.950 ;
        RECT 404.400 36.450 405.450 49.950 ;
        RECT 410.400 40.050 411.450 52.950 ;
        RECT 409.950 37.950 412.050 40.050 ;
        RECT 404.400 35.400 411.450 36.450 ;
        RECT 406.950 31.950 409.050 34.050 ;
        RECT 400.950 28.950 403.050 31.050 ;
        RECT 401.400 25.050 402.450 28.950 ;
        RECT 407.400 25.050 408.450 31.950 ;
        RECT 410.400 25.050 411.450 35.400 ;
        RECT 400.950 22.950 403.050 25.050 ;
        RECT 404.250 23.250 405.750 24.150 ;
        RECT 406.950 22.950 409.050 25.050 ;
        RECT 409.950 22.950 412.050 25.050 ;
        RECT 397.950 19.950 400.050 22.050 ;
        RECT 400.950 20.850 402.750 21.750 ;
        RECT 403.950 19.950 406.050 22.050 ;
        RECT 407.250 20.850 408.750 21.750 ;
        RECT 409.950 19.950 412.050 22.050 ;
        RECT 409.950 17.850 412.050 18.750 ;
        RECT 379.950 13.950 382.050 16.050 ;
        RECT 394.950 13.950 397.050 16.050 ;
        RECT 413.400 10.050 414.450 52.950 ;
        RECT 415.950 49.950 418.050 52.050 ;
        RECT 418.950 49.950 421.050 52.050 ;
        RECT 421.950 49.950 424.050 52.050 ;
        RECT 425.250 50.850 426.750 51.750 ;
        RECT 427.950 49.950 430.050 52.050 ;
        RECT 416.400 36.450 417.450 49.950 ;
        RECT 419.400 40.050 420.450 49.950 ;
        RECT 418.950 37.950 421.050 40.050 ;
        RECT 422.400 36.450 423.450 49.950 ;
        RECT 416.400 35.400 423.450 36.450 ;
        RECT 418.950 28.950 421.050 31.050 ;
        RECT 430.950 28.950 433.050 31.050 ;
        RECT 439.950 28.950 442.050 31.050 ;
        RECT 419.400 18.450 420.450 28.950 ;
        RECT 421.950 20.250 423.750 21.150 ;
        RECT 424.950 19.950 427.050 22.050 ;
        RECT 428.250 20.250 430.050 21.150 ;
        RECT 421.950 18.450 424.050 19.050 ;
        RECT 419.400 17.400 424.050 18.450 ;
        RECT 425.250 17.850 426.750 18.750 ;
        RECT 427.950 18.450 430.050 19.050 ;
        RECT 431.400 18.450 432.450 28.950 ;
        RECT 440.400 28.050 441.450 28.950 ;
        RECT 436.950 25.950 439.050 28.050 ;
        RECT 439.950 25.950 442.050 28.050 ;
        RECT 437.400 25.050 438.450 25.950 ;
        RECT 443.400 25.050 444.450 58.950 ;
        RECT 452.400 58.050 453.450 88.950 ;
        RECT 461.400 73.050 462.450 91.950 ;
        RECT 463.950 82.950 466.050 85.050 ;
        RECT 460.950 70.950 463.050 73.050 ;
        RECT 457.950 59.250 460.050 60.150 ;
        RECT 445.950 55.950 448.050 58.050 ;
        RECT 451.950 57.450 454.050 58.050 ;
        RECT 449.400 56.400 454.050 57.450 ;
        RECT 446.400 40.050 447.450 55.950 ;
        RECT 449.400 52.050 450.450 56.400 ;
        RECT 451.950 55.950 454.050 56.400 ;
        RECT 455.250 56.250 456.750 57.150 ;
        RECT 457.950 55.950 460.050 58.050 ;
        RECT 461.250 56.250 463.050 57.150 ;
        RECT 458.400 55.050 459.450 55.950 ;
        RECT 464.400 55.050 465.450 82.950 ;
        RECT 470.400 76.050 471.450 91.950 ;
        RECT 475.950 89.850 478.050 90.750 ;
        RECT 479.400 88.050 480.450 121.950 ;
        RECT 481.950 112.950 484.050 115.050 ;
        RECT 482.400 94.050 483.450 112.950 ;
        RECT 485.400 112.050 486.450 127.950 ;
        RECT 494.400 127.050 495.450 154.950 ;
        RECT 500.400 139.050 501.450 166.950 ;
        RECT 505.950 164.850 507.750 165.750 ;
        RECT 508.950 163.950 511.050 166.050 ;
        RECT 512.250 164.850 513.750 165.750 ;
        RECT 514.950 163.950 517.050 166.050 ;
        RECT 509.400 157.050 510.450 163.950 ;
        RECT 514.950 161.850 517.050 162.750 ;
        RECT 514.950 157.950 517.050 160.050 ;
        RECT 515.400 157.050 516.450 157.950 ;
        RECT 521.400 157.050 522.450 175.950 ;
        RECT 524.400 169.050 525.450 205.950 ;
        RECT 527.400 184.050 528.450 229.950 ;
        RECT 535.950 226.950 538.050 229.050 ;
        RECT 529.950 214.950 532.050 217.050 ;
        RECT 530.400 202.050 531.450 214.950 ;
        RECT 536.400 205.050 537.450 226.950 ;
        RECT 541.950 220.950 544.050 223.050 ;
        RECT 538.950 214.950 541.050 217.050 ;
        RECT 535.950 202.950 538.050 205.050 ;
        RECT 529.950 199.950 532.050 202.050 ;
        RECT 536.400 199.050 537.450 202.950 ;
        RECT 539.400 202.050 540.450 214.950 ;
        RECT 538.950 199.950 541.050 202.050 ;
        RECT 529.950 197.250 532.050 198.150 ;
        RECT 535.950 196.950 538.050 199.050 ;
        RECT 539.250 197.250 541.050 198.150 ;
        RECT 529.950 193.950 532.050 196.050 ;
        RECT 535.950 194.850 537.750 195.750 ;
        RECT 538.950 193.950 541.050 196.050 ;
        RECT 539.400 187.050 540.450 193.950 ;
        RECT 538.950 184.950 541.050 187.050 ;
        RECT 526.950 181.950 529.050 184.050 ;
        RECT 532.950 181.950 535.050 184.050 ;
        RECT 538.950 181.950 541.050 184.050 ;
        RECT 526.950 175.950 529.050 178.050 ;
        RECT 523.950 166.950 526.050 169.050 ;
        RECT 527.400 166.050 528.450 175.950 ;
        RECT 523.950 164.250 525.750 165.150 ;
        RECT 526.950 163.950 529.050 166.050 ;
        RECT 530.250 164.250 532.050 165.150 ;
        RECT 523.950 160.950 526.050 163.050 ;
        RECT 527.250 161.850 528.750 162.750 ;
        RECT 529.950 160.950 532.050 163.050 ;
        RECT 508.950 154.950 511.050 157.050 ;
        RECT 514.950 154.950 517.050 157.050 ;
        RECT 520.950 154.950 523.050 157.050 ;
        RECT 502.950 142.950 505.050 145.050 ;
        RECT 499.950 136.950 502.050 139.050 ;
        RECT 503.400 130.050 504.450 142.950 ;
        RECT 511.950 139.950 514.050 142.050 ;
        RECT 508.950 136.950 511.050 139.050 ;
        RECT 509.400 130.050 510.450 136.950 ;
        RECT 502.950 129.450 505.050 130.050 ;
        RECT 500.400 128.400 505.050 129.450 ;
        RECT 487.950 124.950 490.050 127.050 ;
        RECT 491.250 125.250 492.750 126.150 ;
        RECT 493.950 124.950 496.050 127.050 ;
        RECT 497.250 125.250 499.050 126.150 ;
        RECT 488.400 115.050 489.450 124.950 ;
        RECT 490.950 121.950 493.050 124.050 ;
        RECT 494.250 122.850 495.750 123.750 ;
        RECT 496.950 121.950 499.050 124.050 ;
        RECT 487.950 112.950 490.050 115.050 ;
        RECT 484.950 109.950 487.050 112.050 ;
        RECT 484.950 106.950 487.050 109.050 ;
        RECT 485.400 100.050 486.450 106.950 ;
        RECT 491.400 103.050 492.450 121.950 ;
        RECT 500.400 118.050 501.450 128.400 ;
        RECT 502.950 127.950 505.050 128.400 ;
        RECT 506.250 128.250 507.750 129.150 ;
        RECT 508.950 127.950 511.050 130.050 ;
        RECT 512.400 127.050 513.450 139.950 ;
        RECT 524.400 139.050 525.450 160.950 ;
        RECT 523.950 136.950 526.050 139.050 ;
        RECT 517.950 127.950 520.050 130.050 ;
        RECT 523.950 129.450 526.050 130.050 ;
        RECT 521.250 128.250 522.750 129.150 ;
        RECT 523.950 128.400 528.450 129.450 ;
        RECT 523.950 127.950 526.050 128.400 ;
        RECT 502.950 125.850 504.750 126.750 ;
        RECT 505.950 124.950 508.050 127.050 ;
        RECT 509.250 125.850 511.050 126.750 ;
        RECT 511.950 124.950 514.050 127.050 ;
        RECT 517.950 125.850 519.750 126.750 ;
        RECT 520.950 124.950 523.050 127.050 ;
        RECT 524.250 125.850 526.050 126.750 ;
        RECT 505.950 121.950 508.050 124.050 ;
        RECT 499.950 115.950 502.050 118.050 ;
        RECT 496.950 112.950 499.050 115.050 ;
        RECT 490.950 100.950 493.050 103.050 ;
        RECT 484.950 97.950 487.050 100.050 ;
        RECT 485.400 97.050 486.450 97.950 ;
        RECT 484.950 94.950 487.050 97.050 ;
        RECT 488.250 95.250 489.750 96.150 ;
        RECT 490.950 94.950 493.050 97.050 ;
        RECT 481.950 91.950 484.050 94.050 ;
        RECT 484.950 92.850 486.750 93.750 ;
        RECT 487.950 91.950 490.050 94.050 ;
        RECT 491.250 92.850 492.750 93.750 ;
        RECT 493.950 91.950 496.050 94.050 ;
        RECT 497.400 91.050 498.450 112.950 ;
        RECT 502.950 109.950 505.050 112.050 ;
        RECT 499.950 91.950 502.050 94.050 ;
        RECT 484.950 88.950 487.050 91.050 ;
        RECT 493.950 89.850 496.050 90.750 ;
        RECT 496.950 88.950 499.050 91.050 ;
        RECT 478.950 85.950 481.050 88.050 ;
        RECT 469.950 73.950 472.050 76.050 ;
        RECT 469.950 67.950 472.050 70.050 ;
        RECT 466.950 61.950 469.050 64.050 ;
        RECT 451.950 53.850 453.750 54.750 ;
        RECT 454.950 52.950 457.050 55.050 ;
        RECT 457.950 52.950 460.050 55.050 ;
        RECT 460.950 52.950 463.050 55.050 ;
        RECT 463.950 52.950 466.050 55.050 ;
        RECT 448.950 49.950 451.050 52.050 ;
        RECT 448.950 46.950 451.050 49.050 ;
        RECT 445.950 37.950 448.050 40.050 ;
        RECT 436.950 22.950 439.050 25.050 ;
        RECT 440.250 23.850 441.750 24.750 ;
        RECT 442.950 22.950 445.050 25.050 ;
        RECT 449.400 22.050 450.450 46.950 ;
        RECT 455.400 28.050 456.450 52.950 ;
        RECT 463.950 34.950 466.050 37.050 ;
        RECT 454.950 25.950 457.050 28.050 ;
        RECT 464.400 25.050 465.450 34.950 ;
        RECT 467.400 25.050 468.450 61.950 ;
        RECT 470.400 58.050 471.450 67.950 ;
        RECT 478.950 61.950 481.050 64.050 ;
        RECT 469.950 55.950 472.050 58.050 ;
        RECT 472.950 56.250 475.050 57.150 ;
        RECT 479.400 55.050 480.450 61.950 ;
        RECT 469.950 52.950 472.050 55.050 ;
        RECT 472.950 52.950 475.050 55.050 ;
        RECT 476.250 53.250 477.750 54.150 ;
        RECT 478.950 52.950 481.050 55.050 ;
        RECT 482.250 53.250 484.050 54.150 ;
        RECT 470.400 37.050 471.450 52.950 ;
        RECT 469.950 34.950 472.050 37.050 ;
        RECT 451.950 22.950 454.050 25.050 ;
        RECT 455.250 23.250 456.750 24.150 ;
        RECT 457.950 22.950 460.050 25.050 ;
        RECT 461.250 23.250 462.750 24.150 ;
        RECT 463.950 22.950 466.050 25.050 ;
        RECT 466.950 22.950 469.050 25.050 ;
        RECT 473.400 22.050 474.450 52.950 ;
        RECT 475.950 49.950 478.050 52.050 ;
        RECT 479.250 50.850 480.750 51.750 ;
        RECT 481.950 49.950 484.050 52.050 ;
        RECT 482.400 49.050 483.450 49.950 ;
        RECT 481.950 46.950 484.050 49.050 ;
        RECT 485.400 46.050 486.450 88.950 ;
        RECT 490.950 58.950 493.050 61.050 ;
        RECT 491.400 55.050 492.450 58.950 ;
        RECT 490.950 52.950 493.050 55.050 ;
        RECT 494.250 53.250 496.050 54.150 ;
        RECT 490.950 50.850 492.750 51.750 ;
        RECT 493.950 49.950 496.050 52.050 ;
        RECT 484.950 43.950 487.050 46.050 ;
        RECT 490.950 43.950 493.050 46.050 ;
        RECT 484.950 28.950 487.050 31.050 ;
        RECT 485.400 28.050 486.450 28.950 ;
        RECT 484.950 25.950 487.050 28.050 ;
        RECT 478.950 22.950 481.050 25.050 ;
        RECT 481.950 22.950 484.050 25.050 ;
        RECT 484.950 23.850 487.050 24.750 ;
        RECT 487.950 23.250 490.050 24.150 ;
        RECT 436.950 20.850 439.050 21.750 ;
        RECT 442.950 20.850 445.050 21.750 ;
        RECT 448.950 19.950 451.050 22.050 ;
        RECT 451.950 20.850 453.750 21.750 ;
        RECT 454.950 19.950 457.050 22.050 ;
        RECT 458.250 20.850 459.750 21.750 ;
        RECT 460.950 19.950 463.050 22.050 ;
        RECT 464.250 20.850 466.050 21.750 ;
        RECT 466.950 19.950 469.050 22.050 ;
        RECT 469.950 20.250 471.750 21.150 ;
        RECT 472.950 19.950 475.050 22.050 ;
        RECT 476.250 20.250 478.050 21.150 ;
        RECT 421.950 16.950 424.050 17.400 ;
        RECT 427.950 17.400 432.450 18.450 ;
        RECT 427.950 16.950 430.050 17.400 ;
        RECT 461.400 13.050 462.450 19.950 ;
        RECT 467.400 18.450 468.450 19.950 ;
        RECT 469.950 18.450 472.050 19.050 ;
        RECT 467.400 17.400 472.050 18.450 ;
        RECT 473.250 17.850 474.750 18.750 ;
        RECT 475.950 18.450 478.050 19.050 ;
        RECT 479.400 18.450 480.450 22.950 ;
        RECT 469.950 16.950 472.050 17.400 ;
        RECT 475.950 17.400 480.450 18.450 ;
        RECT 475.950 16.950 478.050 17.400 ;
        RECT 482.400 13.050 483.450 22.950 ;
        RECT 487.950 19.950 490.050 22.050 ;
        RECT 460.950 10.950 463.050 13.050 ;
        RECT 481.950 10.950 484.050 13.050 ;
        RECT 491.400 10.050 492.450 43.950 ;
        RECT 494.400 37.050 495.450 49.950 ;
        RECT 500.400 46.050 501.450 91.950 ;
        RECT 503.400 91.050 504.450 109.950 ;
        RECT 506.400 97.050 507.450 121.950 ;
        RECT 508.950 112.950 511.050 115.050 ;
        RECT 509.400 100.050 510.450 112.950 ;
        RECT 527.400 112.050 528.450 128.400 ;
        RECT 511.950 109.950 514.050 112.050 ;
        RECT 526.950 109.950 529.050 112.050 ;
        RECT 512.400 100.050 513.450 109.950 ;
        RECT 508.950 97.950 511.050 100.050 ;
        RECT 511.950 97.950 514.050 100.050 ;
        RECT 505.950 94.950 508.050 97.050 ;
        RECT 509.250 95.250 511.050 96.150 ;
        RECT 511.950 95.850 514.050 96.750 ;
        RECT 526.950 96.450 529.050 97.050 ;
        RECT 530.400 96.450 531.450 160.950 ;
        RECT 533.400 121.050 534.450 181.950 ;
        RECT 535.950 166.950 538.050 169.050 ;
        RECT 536.400 163.050 537.450 166.950 ;
        RECT 535.950 160.950 538.050 163.050 ;
        RECT 539.400 154.050 540.450 181.950 ;
        RECT 542.400 178.050 543.450 220.950 ;
        RECT 548.400 211.050 549.450 232.950 ;
        RECT 557.400 232.050 558.450 251.400 ;
        RECT 559.950 250.950 562.050 253.050 ;
        RECT 560.400 235.050 561.450 250.950 ;
        RECT 563.400 247.050 564.450 262.950 ;
        RECT 566.400 250.050 567.450 262.950 ;
        RECT 572.400 262.050 573.450 262.950 ;
        RECT 590.400 262.050 591.450 262.950 ;
        RECT 571.950 259.950 574.050 262.050 ;
        RECT 589.950 259.950 592.050 262.050 ;
        RECT 574.950 256.950 577.050 259.050 ;
        RECT 571.950 253.950 574.050 256.050 ;
        RECT 565.950 247.950 568.050 250.050 ;
        RECT 568.950 247.950 571.050 250.050 ;
        RECT 562.950 244.950 565.050 247.050 ;
        RECT 565.950 244.950 568.050 247.050 ;
        RECT 566.400 238.050 567.450 244.950 ;
        RECT 569.400 244.050 570.450 247.950 ;
        RECT 568.950 241.950 571.050 244.050 ;
        RECT 572.400 240.450 573.450 253.950 ;
        RECT 575.400 250.050 576.450 256.950 ;
        RECT 574.950 247.950 577.050 250.050 ;
        RECT 580.950 244.950 583.050 247.050 ;
        RECT 583.950 244.950 586.050 247.050 ;
        RECT 589.950 244.950 592.050 247.050 ;
        RECT 595.950 244.950 598.050 247.050 ;
        RECT 581.400 244.050 582.450 244.950 ;
        RECT 584.400 244.050 585.450 244.950 ;
        RECT 580.950 241.950 583.050 244.050 ;
        RECT 583.950 241.950 586.050 244.050 ;
        RECT 577.950 240.450 580.050 241.050 ;
        RECT 572.400 239.400 580.050 240.450 ;
        RECT 581.250 239.850 582.750 240.750 ;
        RECT 577.950 238.950 580.050 239.400 ;
        RECT 583.950 238.950 586.050 241.050 ;
        RECT 562.950 236.250 564.750 237.150 ;
        RECT 565.950 235.950 568.050 238.050 ;
        RECT 571.950 237.450 574.050 238.050 ;
        RECT 571.950 236.400 576.450 237.450 ;
        RECT 577.950 236.850 580.050 237.750 ;
        RECT 571.950 235.950 574.050 236.400 ;
        RECT 559.950 232.950 562.050 235.050 ;
        RECT 562.950 232.950 565.050 235.050 ;
        RECT 566.250 233.850 567.750 234.750 ;
        RECT 568.950 232.950 571.050 235.050 ;
        RECT 572.250 233.850 574.050 234.750 ;
        RECT 550.950 229.950 553.050 232.050 ;
        RECT 556.950 229.950 559.050 232.050 ;
        RECT 568.950 230.850 571.050 231.750 ;
        RECT 571.950 229.950 574.050 232.050 ;
        RECT 547.950 208.950 550.050 211.050 ;
        RECT 551.400 207.450 552.450 229.950 ;
        RECT 572.400 223.050 573.450 229.950 ;
        RECT 575.400 226.050 576.450 236.400 ;
        RECT 580.950 235.950 583.050 238.050 ;
        RECT 583.950 236.850 586.050 237.750 ;
        RECT 581.400 229.050 582.450 235.950 ;
        RECT 580.950 226.950 583.050 229.050 ;
        RECT 574.950 223.950 577.050 226.050 ;
        RECT 577.950 223.950 580.050 226.050 ;
        RECT 571.950 220.950 574.050 223.050 ;
        RECT 572.400 220.050 573.450 220.950 ;
        RECT 575.400 220.050 576.450 223.950 ;
        RECT 571.950 217.950 574.050 220.050 ;
        RECT 574.950 217.950 577.050 220.050 ;
        RECT 556.950 211.950 559.050 214.050 ;
        RECT 571.950 211.950 574.050 214.050 ;
        RECT 548.400 206.400 552.450 207.450 ;
        RECT 544.950 196.950 547.050 199.050 ;
        RECT 544.950 194.850 547.050 195.750 ;
        RECT 544.950 190.950 547.050 193.050 ;
        RECT 545.400 184.050 546.450 190.950 ;
        RECT 548.400 190.050 549.450 206.400 ;
        RECT 557.400 199.050 558.450 211.950 ;
        RECT 565.950 203.250 568.050 204.150 ;
        RECT 559.950 199.950 562.050 202.050 ;
        RECT 563.250 200.250 564.750 201.150 ;
        RECT 565.950 199.950 568.050 202.050 ;
        RECT 569.250 200.250 571.050 201.150 ;
        RECT 556.950 196.950 559.050 199.050 ;
        RECT 559.950 197.850 561.750 198.750 ;
        RECT 562.950 196.950 565.050 199.050 ;
        RECT 568.950 196.950 571.050 199.050 ;
        RECT 562.950 193.950 565.050 196.050 ;
        RECT 547.950 187.950 550.050 190.050 ;
        RECT 559.950 187.950 562.050 190.050 ;
        RECT 544.950 181.950 547.050 184.050 ;
        RECT 541.950 175.950 544.050 178.050 ;
        RECT 544.950 166.950 547.050 169.050 ;
        RECT 548.250 167.250 549.750 168.150 ;
        RECT 550.950 166.950 553.050 169.050 ;
        RECT 541.950 163.950 544.050 166.050 ;
        RECT 545.250 164.850 546.750 165.750 ;
        RECT 547.950 163.950 550.050 166.050 ;
        RECT 551.250 164.850 553.050 165.750 ;
        RECT 541.950 161.850 544.050 162.750 ;
        RECT 548.400 154.050 549.450 163.950 ;
        RECT 538.950 151.950 541.050 154.050 ;
        RECT 547.950 151.950 550.050 154.050 ;
        RECT 560.400 139.050 561.450 187.950 ;
        RECT 563.400 171.450 564.450 193.950 ;
        RECT 569.400 192.450 570.450 196.950 ;
        RECT 566.400 191.400 570.450 192.450 ;
        RECT 566.400 175.050 567.450 191.400 ;
        RECT 572.400 187.050 573.450 211.950 ;
        RECT 571.950 184.950 574.050 187.050 ;
        RECT 568.950 181.950 571.050 184.050 ;
        RECT 571.950 181.950 574.050 184.050 ;
        RECT 565.950 172.950 568.050 175.050 ;
        RECT 563.400 170.400 567.450 171.450 ;
        RECT 562.950 167.250 565.050 168.150 ;
        RECT 562.950 163.950 565.050 166.050 ;
        RECT 563.400 157.050 564.450 163.950 ;
        RECT 566.400 160.050 567.450 170.400 ;
        RECT 569.400 169.050 570.450 181.950 ;
        RECT 572.400 178.050 573.450 181.950 ;
        RECT 571.950 175.950 574.050 178.050 ;
        RECT 578.400 171.450 579.450 223.950 ;
        RECT 590.400 223.050 591.450 244.950 ;
        RECT 596.400 244.050 597.450 244.950 ;
        RECT 595.950 243.450 598.050 244.050 ;
        RECT 599.400 243.450 600.450 262.950 ;
        RECT 602.400 261.450 603.450 265.950 ;
        RECT 605.400 264.450 606.450 304.950 ;
        RECT 607.950 289.950 610.050 292.050 ;
        RECT 608.400 274.050 609.450 289.950 ;
        RECT 616.950 277.950 619.050 280.050 ;
        RECT 613.950 274.950 616.050 277.050 ;
        RECT 607.950 271.950 610.050 274.050 ;
        RECT 610.950 271.950 613.050 274.050 ;
        RECT 611.400 271.050 612.450 271.950 ;
        RECT 610.950 268.950 613.050 271.050 ;
        RECT 607.950 266.250 610.050 267.150 ;
        RECT 610.950 266.850 613.050 267.750 ;
        RECT 607.950 264.450 610.050 265.050 ;
        RECT 614.400 264.450 615.450 274.950 ;
        RECT 617.400 274.050 618.450 277.950 ;
        RECT 623.400 274.050 624.450 313.950 ;
        RECT 626.400 307.050 627.450 316.950 ;
        RECT 629.400 310.050 630.450 320.400 ;
        RECT 632.400 313.050 633.450 325.950 ;
        RECT 637.950 322.950 640.050 325.050 ;
        RECT 638.400 316.050 639.450 322.950 ;
        RECT 637.950 313.950 640.050 316.050 ;
        RECT 653.400 313.050 654.450 328.950 ;
        RECT 658.950 325.950 661.050 328.050 ;
        RECT 631.950 310.950 634.050 313.050 ;
        RECT 635.250 311.250 637.050 312.150 ;
        RECT 637.950 311.850 640.050 312.750 ;
        RECT 640.950 311.250 643.050 312.150 ;
        RECT 646.950 310.950 649.050 313.050 ;
        RECT 650.250 311.250 651.750 312.150 ;
        RECT 652.950 310.950 655.050 313.050 ;
        RECT 628.950 307.950 631.050 310.050 ;
        RECT 631.950 308.850 633.750 309.750 ;
        RECT 634.950 307.950 637.050 310.050 ;
        RECT 640.950 307.950 643.050 310.050 ;
        RECT 646.950 308.850 648.750 309.750 ;
        RECT 649.950 307.950 652.050 310.050 ;
        RECT 653.250 308.850 654.750 309.750 ;
        RECT 655.950 307.950 658.050 310.050 ;
        RECT 625.950 304.950 628.050 307.050 ;
        RECT 641.400 304.050 642.450 307.950 ;
        RECT 640.950 301.950 643.050 304.050 ;
        RECT 650.400 301.050 651.450 307.950 ;
        RECT 655.950 305.850 658.050 306.750 ;
        RECT 649.950 298.950 652.050 301.050 ;
        RECT 637.950 295.950 640.050 298.050 ;
        RECT 638.400 280.050 639.450 295.950 ;
        RECT 659.400 294.450 660.450 325.950 ;
        RECT 662.400 298.050 663.450 364.950 ;
        RECT 664.950 344.250 667.050 345.150 ;
        RECT 670.950 343.950 673.050 346.050 ;
        RECT 670.950 341.850 673.050 342.750 ;
        RECT 674.400 316.050 675.450 367.950 ;
        RECT 676.950 349.950 679.050 352.050 ;
        RECT 677.400 322.050 678.450 349.950 ;
        RECT 680.400 346.050 681.450 376.950 ;
        RECT 686.400 370.050 687.450 382.950 ;
        RECT 692.400 382.050 693.450 382.950 ;
        RECT 691.950 379.950 694.050 382.050 ;
        RECT 695.250 380.850 696.750 381.750 ;
        RECT 697.950 379.950 700.050 382.050 ;
        RECT 701.250 380.850 703.050 381.750 ;
        RECT 691.950 377.850 694.050 378.750 ;
        RECT 698.400 378.450 699.450 379.950 ;
        RECT 698.400 377.400 702.450 378.450 ;
        RECT 701.400 373.050 702.450 377.400 ;
        RECT 700.950 370.950 703.050 373.050 ;
        RECT 685.950 367.950 688.050 370.050 ;
        RECT 682.950 361.950 685.050 364.050 ;
        RECT 683.400 346.050 684.450 361.950 ;
        RECT 691.950 352.950 694.050 355.050 ;
        RECT 694.950 352.950 697.050 355.050 ;
        RECT 697.950 352.950 700.050 355.050 ;
        RECT 679.950 343.950 682.050 346.050 ;
        RECT 682.950 343.950 685.050 346.050 ;
        RECT 685.950 344.250 688.050 345.150 ;
        RECT 679.950 341.850 682.050 342.750 ;
        RECT 676.950 319.950 679.050 322.050 ;
        RECT 683.400 319.050 684.450 343.950 ;
        RECT 692.550 334.050 693.750 352.950 ;
        RECT 695.550 348.750 696.750 352.950 ;
        RECT 694.950 346.650 697.050 348.750 ;
        RECT 695.550 334.050 696.750 346.650 ;
        RECT 698.550 334.050 699.750 352.950 ;
        RECT 691.950 331.950 694.050 334.050 ;
        RECT 694.950 331.950 697.050 334.050 ;
        RECT 697.950 331.950 700.050 334.050 ;
        RECT 701.400 330.450 702.450 370.950 ;
        RECT 704.400 346.050 705.450 398.400 ;
        RECT 716.400 397.050 717.450 415.950 ;
        RECT 719.400 400.050 720.450 442.950 ;
        RECT 728.400 423.450 729.450 451.950 ;
        RECT 734.400 448.050 735.450 451.950 ;
        RECT 733.950 445.950 736.050 448.050 ;
        RECT 737.400 439.050 738.450 482.400 ;
        RECT 739.950 481.950 742.050 484.050 ;
        RECT 745.950 481.950 748.050 484.050 ;
        RECT 748.950 481.950 751.050 484.050 ;
        RECT 754.950 483.450 757.050 484.050 ;
        RECT 758.400 483.450 759.450 512.400 ;
        RECT 770.400 511.050 771.450 524.400 ;
        RECT 769.950 508.950 772.050 511.050 ;
        RECT 769.950 502.950 772.050 505.050 ;
        RECT 770.400 492.450 771.450 502.950 ;
        RECT 773.400 495.450 774.450 527.400 ;
        RECT 779.400 526.050 780.450 529.950 ;
        RECT 775.950 524.250 777.750 525.150 ;
        RECT 778.950 523.950 781.050 526.050 ;
        RECT 782.250 524.250 784.050 525.150 ;
        RECT 775.950 520.950 778.050 523.050 ;
        RECT 779.250 521.850 780.750 522.750 ;
        RECT 781.950 520.950 784.050 523.050 ;
        RECT 776.400 505.050 777.450 520.950 ;
        RECT 775.950 502.950 778.050 505.050 ;
        RECT 773.400 494.400 777.450 495.450 ;
        RECT 766.950 491.250 769.050 492.150 ;
        RECT 770.400 491.400 774.450 492.450 ;
        RECT 773.400 490.050 774.450 491.400 ;
        RECT 763.950 488.250 765.750 489.150 ;
        RECT 766.950 487.950 769.050 490.050 ;
        RECT 770.250 488.250 771.750 489.150 ;
        RECT 772.950 487.950 775.050 490.050 ;
        RECT 763.950 484.950 766.050 487.050 ;
        RECT 752.250 482.250 753.750 483.150 ;
        RECT 754.950 482.400 759.450 483.450 ;
        RECT 754.950 481.950 757.050 482.400 ;
        RECT 749.400 481.050 750.450 481.950 ;
        RECT 748.950 478.950 751.050 481.050 ;
        RECT 751.950 478.950 754.050 481.050 ;
        RECT 739.950 457.950 742.050 460.050 ;
        RECT 740.400 450.450 741.450 457.950 ;
        RECT 752.400 457.050 753.450 478.950 ;
        RECT 751.950 454.950 754.050 457.050 ;
        RECT 742.950 452.250 744.750 453.150 ;
        RECT 745.950 451.950 748.050 454.050 ;
        RECT 749.250 452.250 751.050 453.150 ;
        RECT 742.950 450.450 745.050 451.050 ;
        RECT 740.400 449.400 745.050 450.450 ;
        RECT 746.250 449.850 747.750 450.750 ;
        RECT 748.950 450.450 751.050 451.050 ;
        RECT 752.400 450.450 753.450 454.950 ;
        RECT 755.400 451.050 756.450 481.950 ;
        RECT 764.400 481.050 765.450 484.950 ;
        RECT 763.950 478.950 766.050 481.050 ;
        RECT 767.400 472.050 768.450 487.950 ;
        RECT 769.950 484.950 772.050 487.050 ;
        RECT 773.250 485.850 775.050 486.750 ;
        RECT 766.950 469.950 769.050 472.050 ;
        RECT 772.950 469.950 775.050 472.050 ;
        RECT 760.950 457.950 763.050 460.050 ;
        RECT 761.400 454.050 762.450 457.950 ;
        RECT 767.400 454.050 768.450 469.950 ;
        RECT 773.400 460.050 774.450 469.950 ;
        RECT 772.950 457.950 775.050 460.050 ;
        RECT 769.950 455.250 772.050 456.150 ;
        RECT 772.950 455.850 775.050 456.750 ;
        RECT 757.950 452.250 759.750 453.150 ;
        RECT 760.950 451.950 763.050 454.050 ;
        RECT 764.250 452.250 766.050 453.150 ;
        RECT 766.950 451.950 769.050 454.050 ;
        RECT 769.950 451.950 772.050 454.050 ;
        RECT 770.400 451.050 771.450 451.950 ;
        RECT 742.950 448.950 745.050 449.400 ;
        RECT 748.950 449.400 753.450 450.450 ;
        RECT 748.950 448.950 751.050 449.400 ;
        RECT 754.950 448.950 757.050 451.050 ;
        RECT 757.950 448.950 760.050 451.050 ;
        RECT 761.250 449.850 762.750 450.750 ;
        RECT 763.950 448.950 766.050 451.050 ;
        RECT 769.950 448.950 772.050 451.050 ;
        RECT 736.950 436.950 739.050 439.050 ;
        RECT 736.950 427.950 739.050 430.050 ;
        RECT 733.950 424.950 736.050 427.050 ;
        RECT 728.400 422.400 732.450 423.450 ;
        RECT 721.950 418.950 724.050 421.050 ;
        RECT 727.950 418.950 730.050 421.050 ;
        RECT 722.400 418.050 723.450 418.950 ;
        RECT 728.400 418.050 729.450 418.950 ;
        RECT 721.950 415.950 724.050 418.050 ;
        RECT 725.250 416.250 726.750 417.150 ;
        RECT 727.950 415.950 730.050 418.050 ;
        RECT 721.950 413.850 723.750 414.750 ;
        RECT 724.950 412.950 727.050 415.050 ;
        RECT 728.250 413.850 730.050 414.750 ;
        RECT 725.400 412.050 726.450 412.950 ;
        RECT 721.950 409.950 724.050 412.050 ;
        RECT 724.950 409.950 727.050 412.050 ;
        RECT 722.400 409.050 723.450 409.950 ;
        RECT 721.950 406.950 724.050 409.050 ;
        RECT 718.950 397.950 721.050 400.050 ;
        RECT 715.950 394.950 718.050 397.050 ;
        RECT 731.400 394.050 732.450 422.400 ;
        RECT 734.400 412.050 735.450 424.950 ;
        RECT 737.400 417.450 738.450 427.950 ;
        RECT 743.400 427.050 744.450 448.950 ;
        RECT 758.400 445.050 759.450 448.950 ;
        RECT 763.950 445.950 766.050 448.050 ;
        RECT 757.950 442.950 760.050 445.050 ;
        RECT 742.950 424.950 745.050 427.050 ;
        RECT 739.950 417.450 742.050 418.050 ;
        RECT 737.400 416.400 742.050 417.450 ;
        RECT 745.950 417.450 748.050 418.050 ;
        RECT 737.400 412.050 738.450 416.400 ;
        RECT 739.950 415.950 742.050 416.400 ;
        RECT 743.250 416.250 744.750 417.150 ;
        RECT 745.950 416.400 750.450 417.450 ;
        RECT 745.950 415.950 748.050 416.400 ;
        RECT 739.950 413.850 741.750 414.750 ;
        RECT 742.950 412.950 745.050 415.050 ;
        RECT 746.250 413.850 748.050 414.750 ;
        RECT 733.950 409.950 736.050 412.050 ;
        RECT 736.950 409.950 739.050 412.050 ;
        RECT 749.400 409.050 750.450 416.400 ;
        RECT 754.950 415.950 757.050 418.050 ;
        RECT 760.950 416.250 763.050 417.150 ;
        RECT 755.400 415.050 756.450 415.950 ;
        RECT 751.950 413.250 753.750 414.150 ;
        RECT 754.950 412.950 757.050 415.050 ;
        RECT 760.950 414.450 763.050 415.050 ;
        RECT 764.400 414.450 765.450 445.950 ;
        RECT 772.950 415.950 775.050 418.050 ;
        RECT 773.400 415.050 774.450 415.950 ;
        RECT 776.400 415.050 777.450 494.400 ;
        RECT 781.950 490.950 784.050 493.050 ;
        RECT 782.400 487.050 783.450 490.950 ;
        RECT 781.950 484.950 784.050 487.050 ;
        RECT 781.950 482.850 784.050 483.750 ;
        RECT 778.950 455.250 781.050 456.150 ;
        RECT 778.950 451.950 781.050 454.050 ;
        RECT 758.250 413.250 759.750 414.150 ;
        RECT 760.950 413.400 765.450 414.450 ;
        RECT 760.950 412.950 763.050 413.400 ;
        RECT 766.950 412.950 769.050 415.050 ;
        RECT 772.950 412.950 775.050 415.050 ;
        RECT 775.950 412.950 778.050 415.050 ;
        RECT 781.950 414.450 784.050 415.050 ;
        RECT 779.400 413.400 784.050 414.450 ;
        RECT 751.950 409.950 754.050 412.050 ;
        RECT 755.250 410.850 756.750 411.750 ;
        RECT 757.950 409.950 760.050 412.050 ;
        RECT 763.950 409.950 766.050 412.050 ;
        RECT 748.950 406.950 751.050 409.050 ;
        RECT 715.950 391.950 718.050 394.050 ;
        RECT 730.950 391.950 733.050 394.050 ;
        RECT 706.950 380.250 709.050 381.150 ;
        RECT 706.950 376.950 709.050 379.050 ;
        RECT 712.950 377.850 715.050 378.750 ;
        RECT 716.400 355.050 717.450 391.950 ;
        RECT 718.950 388.950 721.050 391.050 ;
        RECT 721.950 388.950 724.050 391.050 ;
        RECT 724.950 388.950 727.050 391.050 ;
        RECT 733.950 389.400 736.050 391.500 ;
        RECT 738.150 389.400 740.250 391.500 ;
        RECT 742.950 389.400 745.050 391.500 ;
        RECT 745.950 389.400 748.050 391.500 ;
        RECT 748.950 389.400 751.050 391.500 ;
        RECT 719.550 370.050 720.750 388.950 ;
        RECT 722.550 376.350 723.750 388.950 ;
        RECT 721.950 374.250 724.050 376.350 ;
        RECT 722.550 370.050 723.750 374.250 ;
        RECT 725.550 370.050 726.750 388.950 ;
        RECT 730.950 385.950 733.050 388.050 ;
        RECT 730.950 383.850 733.050 384.750 ;
        RECT 734.250 380.850 735.450 389.400 ;
        RECT 738.450 383.550 739.650 389.400 ;
        RECT 738.150 381.450 740.250 383.550 ;
        RECT 727.950 376.950 730.050 379.050 ;
        RECT 733.950 378.750 736.050 380.850 ;
        RECT 718.950 367.950 721.050 370.050 ;
        RECT 721.950 367.950 724.050 370.050 ;
        RECT 724.950 367.950 727.050 370.050 ;
        RECT 715.950 352.950 718.050 355.050 ;
        RECT 722.100 353.100 724.200 355.200 ;
        RECT 706.950 350.400 709.050 352.500 ;
        RECT 711.000 350.400 713.100 352.500 ;
        RECT 718.950 350.850 721.050 352.950 ;
        RECT 703.950 343.950 706.050 346.050 ;
        RECT 707.250 344.250 708.450 350.400 ;
        RECT 706.950 342.150 709.050 344.250 ;
        RECT 703.950 338.250 706.050 339.150 ;
        RECT 703.950 334.950 706.050 337.050 ;
        RECT 698.400 329.400 702.450 330.450 ;
        RECT 691.950 319.950 694.050 322.050 ;
        RECT 682.950 316.950 685.050 319.050 ;
        RECT 670.950 313.950 673.050 316.050 ;
        RECT 673.950 313.950 676.050 316.050 ;
        RECT 676.950 313.950 679.050 316.050 ;
        RECT 679.950 313.950 682.050 316.050 ;
        RECT 671.400 313.050 672.450 313.950 ;
        RECT 677.400 313.050 678.450 313.950 ;
        RECT 667.950 310.950 670.050 313.050 ;
        RECT 670.950 310.950 673.050 313.050 ;
        RECT 674.250 311.850 675.750 312.750 ;
        RECT 676.950 310.950 679.050 313.050 ;
        RECT 661.950 295.950 664.050 298.050 ;
        RECT 659.400 293.400 663.450 294.450 ;
        RECT 640.950 280.950 643.050 283.050 ;
        RECT 637.950 277.950 640.050 280.050 ;
        RECT 634.950 274.950 637.050 277.050 ;
        RECT 641.400 276.450 642.450 280.950 ;
        RECT 643.950 277.950 646.050 280.050 ;
        RECT 652.950 277.950 655.050 280.050 ;
        RECT 638.400 275.400 642.450 276.450 ;
        RECT 635.400 274.050 636.450 274.950 ;
        RECT 616.950 271.950 619.050 274.050 ;
        RECT 620.250 272.250 621.750 273.150 ;
        RECT 622.950 271.950 625.050 274.050 ;
        RECT 628.950 271.950 631.050 274.050 ;
        RECT 632.250 272.250 633.750 273.150 ;
        RECT 634.950 271.950 637.050 274.050 ;
        RECT 616.950 269.850 618.750 270.750 ;
        RECT 619.950 268.950 622.050 271.050 ;
        RECT 623.250 269.850 625.050 270.750 ;
        RECT 628.950 269.850 630.750 270.750 ;
        RECT 631.950 268.950 634.050 271.050 ;
        RECT 635.250 269.850 637.050 270.750 ;
        RECT 605.400 263.400 610.050 264.450 ;
        RECT 607.950 262.950 610.050 263.400 ;
        RECT 611.400 263.400 615.450 264.450 ;
        RECT 602.400 260.400 606.450 261.450 ;
        RECT 595.950 242.400 600.450 243.450 ;
        RECT 595.950 241.950 598.050 242.400 ;
        RECT 592.950 239.250 595.050 240.150 ;
        RECT 595.950 239.850 598.050 240.750 ;
        RECT 598.950 239.250 600.750 240.150 ;
        RECT 601.950 238.950 604.050 241.050 ;
        RECT 592.950 235.950 595.050 238.050 ;
        RECT 598.950 237.450 601.050 238.050 ;
        RECT 596.400 236.400 601.050 237.450 ;
        RECT 602.250 236.850 604.050 237.750 ;
        RECT 593.400 235.050 594.450 235.950 ;
        RECT 592.950 232.950 595.050 235.050 ;
        RECT 589.950 220.950 592.050 223.050 ;
        RECT 596.400 220.050 597.450 236.400 ;
        RECT 598.950 235.950 601.050 236.400 ;
        RECT 601.950 232.950 604.050 235.050 ;
        RECT 598.950 226.950 601.050 229.050 ;
        RECT 595.950 217.950 598.050 220.050 ;
        RECT 580.950 202.950 583.050 205.050 ;
        RECT 581.400 202.050 582.450 202.950 ;
        RECT 596.400 202.050 597.450 217.950 ;
        RECT 580.950 199.950 583.050 202.050 ;
        RECT 595.950 199.950 598.050 202.050 ;
        RECT 581.400 199.050 582.450 199.950 ;
        RECT 599.400 199.050 600.450 226.950 ;
        RECT 602.400 217.050 603.450 232.950 ;
        RECT 605.400 226.050 606.450 260.400 ;
        RECT 607.950 241.950 610.050 244.050 ;
        RECT 608.400 238.050 609.450 241.950 ;
        RECT 611.400 238.050 612.450 263.400 ;
        RECT 620.400 262.050 621.450 268.950 ;
        RECT 632.400 267.450 633.450 268.950 ;
        RECT 638.400 267.450 639.450 275.400 ;
        RECT 640.950 271.950 643.050 274.050 ;
        RECT 632.400 266.400 639.450 267.450 ;
        RECT 628.950 262.950 631.050 265.050 ;
        RECT 616.950 259.950 619.050 262.050 ;
        RECT 619.950 259.950 622.050 262.050 ;
        RECT 617.400 247.050 618.450 259.950 ;
        RECT 629.400 259.050 630.450 262.950 ;
        RECT 641.400 262.050 642.450 271.950 ;
        RECT 644.400 268.050 645.450 277.950 ;
        RECT 646.950 274.950 649.050 277.050 ;
        RECT 643.950 265.950 646.050 268.050 ;
        RECT 647.400 265.050 648.450 274.950 ;
        RECT 653.400 271.050 654.450 277.950 ;
        RECT 658.950 274.950 661.050 277.050 ;
        RECT 659.400 271.050 660.450 274.950 ;
        RECT 649.950 269.250 651.750 270.150 ;
        RECT 652.950 268.950 655.050 271.050 ;
        RECT 658.950 268.950 661.050 271.050 ;
        RECT 662.400 268.050 663.450 293.400 ;
        RECT 668.400 277.050 669.450 310.950 ;
        RECT 670.950 308.850 673.050 309.750 ;
        RECT 676.950 308.850 679.050 309.750 ;
        RECT 673.950 304.950 676.050 307.050 ;
        RECT 680.400 306.450 681.450 313.950 ;
        RECT 685.950 310.950 688.050 313.050 ;
        RECT 686.400 310.050 687.450 310.950 ;
        RECT 682.950 308.250 684.750 309.150 ;
        RECT 685.950 307.950 688.050 310.050 ;
        RECT 689.250 308.250 691.050 309.150 ;
        RECT 682.950 306.450 685.050 307.050 ;
        RECT 680.400 305.400 685.050 306.450 ;
        RECT 686.250 305.850 687.750 306.750 ;
        RECT 682.950 304.950 685.050 305.400 ;
        RECT 688.950 304.950 691.050 307.050 ;
        RECT 664.950 274.950 667.050 277.050 ;
        RECT 667.950 274.950 670.050 277.050 ;
        RECT 649.950 265.950 652.050 268.050 ;
        RECT 653.250 266.850 655.050 267.750 ;
        RECT 655.950 266.250 658.050 267.150 ;
        RECT 658.950 266.850 661.050 267.750 ;
        RECT 661.950 265.950 664.050 268.050 ;
        RECT 665.400 267.450 666.450 274.950 ;
        RECT 670.950 271.950 673.050 274.050 ;
        RECT 667.950 269.250 670.050 270.150 ;
        RECT 670.950 269.850 673.050 270.750 ;
        RECT 667.950 267.450 670.050 268.050 ;
        RECT 665.400 266.400 670.050 267.450 ;
        RECT 667.950 265.950 670.050 266.400 ;
        RECT 670.950 265.950 673.050 268.050 ;
        RECT 646.950 262.950 649.050 265.050 ;
        RECT 655.950 262.950 658.050 265.050 ;
        RECT 661.950 262.950 664.050 265.050 ;
        RECT 640.950 259.950 643.050 262.050 ;
        RECT 646.950 259.950 649.050 262.050 ;
        RECT 652.950 259.950 655.050 262.050 ;
        RECT 628.950 256.950 631.050 259.050 ;
        RECT 634.950 253.950 637.050 256.050 ;
        RECT 616.950 244.950 619.050 247.050 ;
        RECT 635.400 244.050 636.450 253.950 ;
        RECT 643.950 244.950 646.050 247.050 ;
        RECT 619.950 241.950 622.050 244.050 ;
        RECT 625.950 241.950 628.050 244.050 ;
        RECT 634.950 241.950 637.050 244.050 ;
        RECT 613.950 238.950 616.050 241.050 ;
        RECT 614.400 238.050 615.450 238.950 ;
        RECT 607.950 235.950 610.050 238.050 ;
        RECT 610.950 235.950 613.050 238.050 ;
        RECT 613.950 235.950 616.050 238.050 ;
        RECT 617.250 236.250 619.050 237.150 ;
        RECT 620.400 235.050 621.450 241.950 ;
        RECT 622.950 239.250 625.050 240.150 ;
        RECT 625.950 239.850 628.050 240.750 ;
        RECT 631.950 240.450 634.050 241.050 ;
        RECT 628.950 239.250 630.750 240.150 ;
        RECT 631.950 239.400 636.450 240.450 ;
        RECT 631.950 238.950 634.050 239.400 ;
        RECT 622.950 235.950 625.050 238.050 ;
        RECT 625.950 235.950 628.050 238.050 ;
        RECT 628.950 235.950 631.050 238.050 ;
        RECT 632.250 236.850 634.050 237.750 ;
        RECT 607.950 233.850 609.750 234.750 ;
        RECT 610.950 232.950 613.050 235.050 ;
        RECT 614.250 233.850 615.750 234.750 ;
        RECT 616.950 232.950 619.050 235.050 ;
        RECT 619.950 232.950 622.050 235.050 ;
        RECT 610.950 230.850 613.050 231.750 ;
        RECT 617.400 226.050 618.450 232.950 ;
        RECT 604.950 223.950 607.050 226.050 ;
        RECT 616.950 223.950 619.050 226.050 ;
        RECT 616.950 220.950 619.050 223.050 ;
        RECT 601.950 214.950 604.050 217.050 ;
        RECT 604.950 208.950 607.050 211.050 ;
        RECT 613.950 208.950 616.050 211.050 ;
        RECT 580.950 196.950 583.050 199.050 ;
        RECT 592.950 198.450 595.050 199.050 ;
        RECT 590.400 197.400 595.050 198.450 ;
        RECT 580.950 194.850 583.050 195.750 ;
        RECT 583.950 194.250 586.050 195.150 ;
        RECT 583.950 190.950 586.050 193.050 ;
        RECT 575.400 170.400 579.450 171.450 ;
        RECT 568.950 166.950 571.050 169.050 ;
        RECT 572.250 167.250 574.050 168.150 ;
        RECT 568.950 164.850 570.750 165.750 ;
        RECT 571.950 163.950 574.050 166.050 ;
        RECT 565.950 157.950 568.050 160.050 ;
        RECT 568.950 157.950 571.050 160.050 ;
        RECT 562.950 154.950 565.050 157.050 ;
        RECT 562.950 151.950 565.050 154.050 ;
        RECT 563.400 142.050 564.450 151.950 ;
        RECT 562.950 139.950 565.050 142.050 ;
        RECT 541.950 136.950 544.050 139.050 ;
        RECT 559.950 136.950 562.050 139.050 ;
        RECT 535.950 128.250 538.050 129.150 ;
        RECT 542.400 127.050 543.450 136.950 ;
        RECT 550.950 131.250 553.050 132.150 ;
        RECT 556.950 130.950 559.050 133.050 ;
        RECT 559.950 130.950 562.050 133.050 ;
        RECT 557.400 130.050 558.450 130.950 ;
        RECT 547.950 128.250 549.750 129.150 ;
        RECT 550.950 127.950 553.050 130.050 ;
        RECT 554.250 128.250 555.750 129.150 ;
        RECT 556.950 127.950 559.050 130.050 ;
        RECT 551.400 127.050 552.450 127.950 ;
        RECT 560.400 127.050 561.450 130.950 ;
        RECT 535.950 124.950 538.050 127.050 ;
        RECT 539.250 125.250 540.750 126.150 ;
        RECT 541.950 124.950 544.050 127.050 ;
        RECT 545.250 125.250 547.050 126.150 ;
        RECT 547.950 124.950 550.050 127.050 ;
        RECT 550.950 124.950 553.050 127.050 ;
        RECT 553.950 124.950 556.050 127.050 ;
        RECT 557.250 125.850 559.050 126.750 ;
        RECT 559.950 124.950 562.050 127.050 ;
        RECT 538.950 121.950 541.050 124.050 ;
        RECT 542.250 122.850 543.750 123.750 ;
        RECT 544.950 123.450 547.050 124.050 ;
        RECT 548.400 123.450 549.450 124.950 ;
        RECT 554.400 124.050 555.450 124.950 ;
        RECT 563.400 124.050 564.450 139.950 ;
        RECT 569.400 133.050 570.450 157.950 ;
        RECT 575.400 147.450 576.450 170.400 ;
        RECT 584.400 169.050 585.450 190.950 ;
        RECT 590.400 187.050 591.450 197.400 ;
        RECT 592.950 196.950 595.050 197.400 ;
        RECT 598.950 196.950 601.050 199.050 ;
        RECT 592.950 194.850 595.050 195.750 ;
        RECT 595.950 194.250 598.050 195.150 ;
        RECT 598.950 193.950 601.050 196.050 ;
        RECT 595.950 190.950 598.050 193.050 ;
        RECT 589.950 184.950 592.050 187.050 ;
        RECT 596.400 181.050 597.450 190.950 ;
        RECT 595.950 178.950 598.050 181.050 ;
        RECT 589.950 175.950 592.050 178.050 ;
        RECT 590.400 171.450 591.450 175.950 ;
        RECT 599.400 175.050 600.450 193.950 ;
        RECT 601.950 187.950 604.050 190.050 ;
        RECT 598.950 172.950 601.050 175.050 ;
        RECT 587.400 170.400 591.450 171.450 ;
        RECT 577.950 168.450 580.050 169.050 ;
        RECT 577.950 167.400 582.450 168.450 ;
        RECT 577.950 166.950 580.050 167.400 ;
        RECT 577.950 164.850 580.050 165.750 ;
        RECT 581.400 163.050 582.450 167.400 ;
        RECT 583.950 166.950 586.050 169.050 ;
        RECT 580.950 160.950 583.050 163.050 ;
        RECT 572.400 146.400 576.450 147.450 ;
        RECT 568.950 130.950 571.050 133.050 ;
        RECT 572.400 127.050 573.450 146.400 ;
        RECT 574.950 142.950 577.050 145.050 ;
        RECT 575.400 130.050 576.450 142.950 ;
        RECT 581.400 136.050 582.450 160.950 ;
        RECT 580.950 133.950 583.050 136.050 ;
        RECT 580.950 130.950 583.050 133.050 ;
        RECT 574.950 127.950 577.050 130.050 ;
        RECT 568.950 125.250 571.050 126.150 ;
        RECT 571.950 124.950 574.050 127.050 ;
        RECT 574.950 125.850 577.050 126.750 ;
        RECT 577.950 125.250 580.050 126.150 ;
        RECT 544.950 122.400 552.450 123.450 ;
        RECT 544.950 121.950 547.050 122.400 ;
        RECT 539.400 121.050 540.450 121.950 ;
        RECT 532.950 118.950 535.050 121.050 ;
        RECT 538.950 118.950 541.050 121.050 ;
        RECT 547.950 103.950 550.050 106.050 ;
        RECT 535.950 97.950 538.050 100.050 ;
        RECT 514.950 95.250 517.050 96.150 ;
        RECT 526.950 95.400 531.450 96.450 ;
        RECT 526.950 94.950 529.050 95.400 ;
        RECT 530.400 94.050 531.450 95.400 ;
        RECT 505.950 92.850 507.750 93.750 ;
        RECT 508.950 91.950 511.050 94.050 ;
        RECT 514.950 91.950 517.050 94.050 ;
        RECT 523.950 91.950 526.050 94.050 ;
        RECT 529.950 91.950 532.050 94.050 ;
        RECT 533.250 92.250 535.050 93.150 ;
        RECT 502.950 88.950 505.050 91.050 ;
        RECT 509.400 67.050 510.450 91.950 ;
        RECT 515.400 91.050 516.450 91.950 ;
        RECT 514.950 88.950 517.050 91.050 ;
        RECT 523.950 89.850 525.750 90.750 ;
        RECT 526.950 88.950 529.050 91.050 ;
        RECT 530.250 89.850 531.750 90.750 ;
        RECT 532.950 88.950 535.050 91.050 ;
        RECT 523.950 85.950 526.050 88.050 ;
        RECT 526.950 86.850 529.050 87.750 ;
        RECT 508.950 64.950 511.050 67.050 ;
        RECT 505.950 55.950 508.050 58.050 ;
        RECT 511.950 55.950 514.050 58.050 ;
        RECT 502.950 52.950 505.050 55.050 ;
        RECT 503.400 49.050 504.450 52.950 ;
        RECT 502.950 46.950 505.050 49.050 ;
        RECT 499.950 43.950 502.050 46.050 ;
        RECT 496.950 37.950 499.050 40.050 ;
        RECT 493.950 34.950 496.050 37.050 ;
        RECT 493.950 25.950 496.050 28.050 ;
        RECT 494.400 19.050 495.450 25.950 ;
        RECT 497.400 25.050 498.450 37.950 ;
        RECT 506.400 25.050 507.450 55.950 ;
        RECT 512.400 55.050 513.450 55.950 ;
        RECT 508.950 53.250 510.750 54.150 ;
        RECT 511.950 52.950 514.050 55.050 ;
        RECT 508.950 49.950 511.050 52.050 ;
        RECT 512.250 50.850 514.050 51.750 ;
        RECT 517.950 50.850 520.050 51.750 ;
        RECT 509.400 46.050 510.450 49.950 ;
        RECT 508.950 43.950 511.050 46.050 ;
        RECT 517.950 37.950 520.050 40.050 ;
        RECT 514.950 28.950 517.050 31.050 ;
        RECT 515.400 28.050 516.450 28.950 ;
        RECT 514.950 25.950 517.050 28.050 ;
        RECT 518.400 25.050 519.450 37.950 ;
        RECT 496.950 22.950 499.050 25.050 ;
        RECT 500.250 23.250 501.750 24.150 ;
        RECT 502.950 22.950 505.050 25.050 ;
        RECT 505.950 22.950 508.050 25.050 ;
        RECT 511.950 22.950 514.050 25.050 ;
        RECT 515.250 23.850 516.750 24.750 ;
        RECT 517.950 22.950 520.050 25.050 ;
        RECT 506.400 22.050 507.450 22.950 ;
        RECT 496.950 20.850 498.750 21.750 ;
        RECT 499.950 19.950 502.050 22.050 ;
        RECT 503.250 20.850 504.750 21.750 ;
        RECT 505.950 19.950 508.050 22.050 ;
        RECT 511.950 20.850 514.050 21.750 ;
        RECT 517.950 20.850 520.050 21.750 ;
        RECT 493.950 16.950 496.050 19.050 ;
        RECT 505.950 17.850 508.050 18.750 ;
        RECT 412.950 7.950 415.050 10.050 ;
        RECT 490.950 7.950 493.050 10.050 ;
        RECT 524.400 7.050 525.450 85.950 ;
        RECT 526.950 82.950 529.050 85.050 ;
        RECT 527.400 28.050 528.450 82.950 ;
        RECT 533.400 79.050 534.450 88.950 ;
        RECT 532.950 76.950 535.050 79.050 ;
        RECT 529.950 64.950 532.050 67.050 ;
        RECT 530.400 40.050 531.450 64.950 ;
        RECT 536.400 43.050 537.450 97.950 ;
        RECT 548.400 97.050 549.450 103.950 ;
        RECT 547.950 94.950 550.050 97.050 ;
        RECT 538.950 91.950 541.050 94.050 ;
        RECT 541.950 92.250 543.750 93.150 ;
        RECT 544.950 91.950 547.050 94.050 ;
        RECT 548.250 92.250 550.050 93.150 ;
        RECT 539.400 85.050 540.450 91.950 ;
        RECT 541.950 88.950 544.050 91.050 ;
        RECT 545.250 89.850 546.750 90.750 ;
        RECT 547.950 88.950 550.050 91.050 ;
        RECT 548.400 88.050 549.450 88.950 ;
        RECT 547.950 85.950 550.050 88.050 ;
        RECT 538.950 82.950 541.050 85.050 ;
        RECT 538.950 79.950 541.050 82.050 ;
        RECT 547.950 79.950 550.050 82.050 ;
        RECT 539.400 58.050 540.450 79.950 ;
        RECT 538.950 55.950 541.050 58.050 ;
        RECT 539.400 55.050 540.450 55.950 ;
        RECT 548.400 55.050 549.450 79.950 ;
        RECT 538.950 52.950 541.050 55.050 ;
        RECT 547.950 52.950 550.050 55.050 ;
        RECT 551.400 52.050 552.450 122.400 ;
        RECT 553.950 121.950 556.050 124.050 ;
        RECT 562.950 121.950 565.050 124.050 ;
        RECT 568.950 121.950 571.050 124.050 ;
        RECT 577.950 121.950 580.050 124.050 ;
        RECT 569.400 106.050 570.450 121.950 ;
        RECT 568.950 103.950 571.050 106.050 ;
        RECT 553.950 100.950 556.050 103.050 ;
        RECT 554.400 97.050 555.450 100.950 ;
        RECT 578.400 100.050 579.450 121.950 ;
        RECT 581.400 112.050 582.450 130.950 ;
        RECT 587.400 124.050 588.450 170.400 ;
        RECT 598.950 169.950 601.050 172.050 ;
        RECT 599.400 169.050 600.450 169.950 ;
        RECT 589.950 168.450 592.050 169.050 ;
        RECT 589.950 167.400 597.450 168.450 ;
        RECT 589.950 166.950 592.050 167.400 ;
        RECT 589.950 164.850 592.050 165.750 ;
        RECT 592.950 164.250 595.050 165.150 ;
        RECT 592.950 160.950 595.050 163.050 ;
        RECT 593.400 160.050 594.450 160.950 ;
        RECT 592.950 157.950 595.050 160.050 ;
        RECT 593.400 157.050 594.450 157.950 ;
        RECT 592.950 154.950 595.050 157.050 ;
        RECT 596.400 142.050 597.450 167.400 ;
        RECT 598.950 166.950 601.050 169.050 ;
        RECT 598.950 164.850 601.050 165.750 ;
        RECT 602.400 142.050 603.450 187.950 ;
        RECT 605.400 175.050 606.450 208.950 ;
        RECT 607.950 200.250 610.050 201.150 ;
        RECT 614.400 199.050 615.450 208.950 ;
        RECT 617.400 202.050 618.450 220.950 ;
        RECT 623.400 208.050 624.450 235.950 ;
        RECT 626.400 235.050 627.450 235.950 ;
        RECT 629.400 235.050 630.450 235.950 ;
        RECT 625.950 232.950 628.050 235.050 ;
        RECT 628.950 234.450 631.050 235.050 ;
        RECT 628.950 233.400 633.450 234.450 ;
        RECT 628.950 232.950 631.050 233.400 ;
        RECT 622.950 205.950 625.050 208.050 ;
        RECT 626.400 205.050 627.450 232.950 ;
        RECT 628.950 223.950 631.050 226.050 ;
        RECT 622.950 203.250 625.050 204.150 ;
        RECT 625.950 202.950 628.050 205.050 ;
        RECT 629.400 202.050 630.450 223.950 ;
        RECT 632.400 219.450 633.450 233.400 ;
        RECT 635.400 229.050 636.450 239.400 ;
        RECT 637.950 238.950 640.050 241.050 ;
        RECT 640.950 238.950 643.050 241.050 ;
        RECT 634.950 226.950 637.050 229.050 ;
        RECT 635.400 223.050 636.450 226.950 ;
        RECT 634.950 220.950 637.050 223.050 ;
        RECT 632.400 218.400 636.450 219.450 ;
        RECT 635.400 208.050 636.450 218.400 ;
        RECT 638.400 214.050 639.450 238.950 ;
        RECT 637.950 211.950 640.050 214.050 ;
        RECT 631.950 205.950 634.050 208.050 ;
        RECT 634.950 205.950 637.050 208.050 ;
        RECT 616.950 199.950 619.050 202.050 ;
        RECT 619.950 200.250 621.750 201.150 ;
        RECT 622.950 199.950 625.050 202.050 ;
        RECT 626.250 200.250 627.750 201.150 ;
        RECT 628.950 199.950 631.050 202.050 ;
        RECT 607.950 196.950 610.050 199.050 ;
        RECT 611.250 197.250 612.750 198.150 ;
        RECT 613.950 196.950 616.050 199.050 ;
        RECT 617.250 197.250 619.050 198.150 ;
        RECT 619.950 196.950 622.050 199.050 ;
        RECT 608.400 190.050 609.450 196.950 ;
        RECT 610.950 193.950 613.050 196.050 ;
        RECT 614.250 194.850 615.750 195.750 ;
        RECT 616.950 193.950 619.050 196.050 ;
        RECT 619.950 193.950 622.050 196.050 ;
        RECT 607.950 187.950 610.050 190.050 ;
        RECT 604.950 172.950 607.050 175.050 ;
        RECT 607.950 172.950 610.050 175.050 ;
        RECT 608.400 172.050 609.450 172.950 ;
        RECT 604.950 169.950 607.050 172.050 ;
        RECT 607.950 169.950 610.050 172.050 ;
        RECT 605.400 168.450 606.450 169.950 ;
        RECT 611.400 169.050 612.450 193.950 ;
        RECT 620.400 184.050 621.450 193.950 ;
        RECT 623.400 190.050 624.450 199.950 ;
        RECT 632.400 199.050 633.450 205.950 ;
        RECT 635.400 202.050 636.450 205.950 ;
        RECT 641.400 202.050 642.450 238.950 ;
        RECT 644.400 238.050 645.450 244.950 ;
        RECT 647.400 241.050 648.450 259.950 ;
        RECT 653.400 243.450 654.450 259.950 ;
        RECT 656.400 247.050 657.450 262.950 ;
        RECT 655.950 244.950 658.050 247.050 ;
        RECT 653.400 242.400 657.450 243.450 ;
        RECT 646.950 238.950 649.050 241.050 ;
        RECT 650.250 239.250 651.750 240.150 ;
        RECT 652.950 238.950 655.050 241.050 ;
        RECT 656.400 238.050 657.450 242.400 ;
        RECT 658.950 241.950 661.050 244.050 ;
        RECT 643.950 235.950 646.050 238.050 ;
        RECT 647.250 236.850 648.750 237.750 ;
        RECT 649.950 235.950 652.050 238.050 ;
        RECT 653.250 236.850 655.050 237.750 ;
        RECT 655.950 235.950 658.050 238.050 ;
        RECT 643.950 233.850 646.050 234.750 ;
        RECT 634.950 199.950 637.050 202.050 ;
        RECT 640.950 199.950 643.050 202.050 ;
        RECT 646.950 200.250 649.050 201.150 ;
        RECT 625.950 196.950 628.050 199.050 ;
        RECT 629.250 197.850 631.050 198.750 ;
        RECT 631.950 196.950 634.050 199.050 ;
        RECT 634.950 196.950 637.050 199.050 ;
        RECT 637.950 197.250 639.750 198.150 ;
        RECT 640.950 196.950 643.050 199.050 ;
        RECT 644.250 197.250 645.750 198.150 ;
        RECT 646.950 196.950 649.050 199.050 ;
        RECT 622.950 187.950 625.050 190.050 ;
        RECT 635.400 187.050 636.450 196.950 ;
        RECT 637.950 193.950 640.050 196.050 ;
        RECT 641.250 194.850 642.750 195.750 ;
        RECT 643.950 193.950 646.050 196.050 ;
        RECT 634.950 184.950 637.050 187.050 ;
        RECT 619.950 181.950 622.050 184.050 ;
        RECT 613.950 175.950 616.050 178.050 ;
        RECT 614.400 169.050 615.450 175.950 ;
        RECT 619.950 172.950 622.050 175.050 ;
        RECT 631.950 172.950 634.050 175.050 ;
        RECT 620.400 169.050 621.450 172.950 ;
        RECT 628.950 169.950 631.050 172.050 ;
        RECT 629.400 169.050 630.450 169.950 ;
        RECT 605.400 167.400 609.450 168.450 ;
        RECT 604.950 163.950 607.050 166.050 ;
        RECT 608.400 165.450 609.450 167.400 ;
        RECT 610.950 166.950 613.050 169.050 ;
        RECT 613.950 166.950 616.050 169.050 ;
        RECT 617.250 167.250 618.750 168.150 ;
        RECT 619.950 166.950 622.050 169.050 ;
        RECT 622.950 166.950 625.050 169.050 ;
        RECT 626.250 167.250 627.750 168.150 ;
        RECT 628.950 166.950 631.050 169.050 ;
        RECT 632.400 166.050 633.450 172.950 ;
        RECT 638.400 172.050 639.450 193.950 ;
        RECT 634.950 169.950 637.050 172.050 ;
        RECT 637.950 169.950 640.050 172.050 ;
        RECT 610.950 165.450 613.050 166.050 ;
        RECT 608.400 164.400 613.050 165.450 ;
        RECT 614.250 164.850 615.750 165.750 ;
        RECT 605.400 163.050 606.450 163.950 ;
        RECT 604.950 160.950 607.050 163.050 ;
        RECT 604.950 157.950 607.050 160.050 ;
        RECT 595.950 139.950 598.050 142.050 ;
        RECT 601.950 139.950 604.050 142.050 ;
        RECT 592.950 131.250 595.050 132.150 ;
        RECT 598.950 130.950 601.050 133.050 ;
        RECT 599.400 130.050 600.450 130.950 ;
        RECT 589.950 128.250 591.750 129.150 ;
        RECT 592.950 127.950 595.050 130.050 ;
        RECT 596.250 128.250 597.750 129.150 ;
        RECT 598.950 127.950 601.050 130.050 ;
        RECT 605.400 129.450 606.450 157.950 ;
        RECT 608.400 154.050 609.450 164.400 ;
        RECT 610.950 163.950 613.050 164.400 ;
        RECT 616.950 163.950 619.050 166.050 ;
        RECT 620.250 164.850 622.050 165.750 ;
        RECT 622.950 164.850 624.750 165.750 ;
        RECT 625.950 163.950 628.050 166.050 ;
        RECT 629.250 164.850 630.750 165.750 ;
        RECT 631.950 163.950 634.050 166.050 ;
        RECT 626.400 163.050 627.450 163.950 ;
        RECT 610.950 161.850 613.050 162.750 ;
        RECT 625.950 160.950 628.050 163.050 ;
        RECT 628.950 160.950 631.050 163.050 ;
        RECT 631.950 161.850 634.050 162.750 ;
        RECT 607.950 151.950 610.050 154.050 ;
        RECT 610.950 151.950 613.050 154.050 ;
        RECT 611.400 145.050 612.450 151.950 ;
        RECT 610.950 142.950 613.050 145.050 ;
        RECT 616.950 139.950 619.050 142.050 ;
        RECT 613.950 130.950 616.050 133.050 ;
        RECT 614.400 130.050 615.450 130.950 ;
        RECT 607.950 129.450 610.050 130.050 ;
        RECT 605.400 128.400 610.050 129.450 ;
        RECT 593.400 127.050 594.450 127.950 ;
        RECT 589.950 124.950 592.050 127.050 ;
        RECT 592.950 124.950 595.050 127.050 ;
        RECT 595.950 124.950 598.050 127.050 ;
        RECT 599.250 125.850 601.050 126.750 ;
        RECT 586.950 121.950 589.050 124.050 ;
        RECT 590.400 115.050 591.450 124.950 ;
        RECT 596.400 121.050 597.450 124.950 ;
        RECT 605.400 124.050 606.450 128.400 ;
        RECT 607.950 127.950 610.050 128.400 ;
        RECT 611.250 128.250 612.750 129.150 ;
        RECT 613.950 127.950 616.050 130.050 ;
        RECT 607.950 125.850 609.750 126.750 ;
        RECT 610.950 124.950 613.050 127.050 ;
        RECT 614.250 125.850 616.050 126.750 ;
        RECT 598.950 121.950 601.050 124.050 ;
        RECT 604.950 121.950 607.050 124.050 ;
        RECT 592.950 118.950 595.050 121.050 ;
        RECT 595.950 118.950 598.050 121.050 ;
        RECT 593.400 115.050 594.450 118.950 ;
        RECT 586.950 112.950 589.050 115.050 ;
        RECT 589.950 112.950 592.050 115.050 ;
        RECT 592.950 112.950 595.050 115.050 ;
        RECT 580.950 109.950 583.050 112.050 ;
        RECT 577.950 97.950 580.050 100.050 ;
        RECT 581.400 97.050 582.450 109.950 ;
        RECT 553.950 94.950 556.050 97.050 ;
        RECT 562.950 96.450 565.050 97.050 ;
        RECT 562.950 95.400 567.450 96.450 ;
        RECT 562.950 94.950 565.050 95.400 ;
        RECT 553.950 92.850 556.050 93.750 ;
        RECT 559.950 92.250 562.050 93.150 ;
        RECT 562.950 92.850 565.050 93.750 ;
        RECT 559.950 88.950 562.050 91.050 ;
        RECT 560.400 79.050 561.450 88.950 ;
        RECT 562.950 85.950 565.050 88.050 ;
        RECT 563.400 79.050 564.450 85.950 ;
        RECT 566.400 85.050 567.450 95.400 ;
        RECT 577.950 94.950 580.050 97.050 ;
        RECT 580.950 94.950 583.050 97.050 ;
        RECT 574.950 91.950 577.050 94.050 ;
        RECT 578.400 91.050 579.450 94.950 ;
        RECT 581.400 94.050 582.450 94.950 ;
        RECT 580.950 91.950 583.050 94.050 ;
        RECT 584.250 92.250 586.050 93.150 ;
        RECT 574.950 89.850 576.750 90.750 ;
        RECT 577.950 88.950 580.050 91.050 ;
        RECT 581.250 89.850 582.750 90.750 ;
        RECT 583.950 88.950 586.050 91.050 ;
        RECT 584.400 88.050 585.450 88.950 ;
        RECT 577.950 86.850 580.050 87.750 ;
        RECT 583.950 85.950 586.050 88.050 ;
        RECT 565.950 82.950 568.050 85.050 ;
        RECT 559.950 76.950 562.050 79.050 ;
        RECT 562.950 76.950 565.050 79.050 ;
        RECT 587.400 76.050 588.450 112.950 ;
        RECT 592.950 100.950 595.050 103.050 ;
        RECT 589.950 97.950 592.050 100.050 ;
        RECT 590.400 91.050 591.450 97.950 ;
        RECT 593.400 97.050 594.450 100.950 ;
        RECT 599.400 100.050 600.450 121.950 ;
        RECT 604.950 109.950 607.050 112.050 ;
        RECT 598.950 97.950 601.050 100.050 ;
        RECT 592.950 94.950 595.050 97.050 ;
        RECT 596.250 95.250 598.050 96.150 ;
        RECT 598.950 95.850 601.050 96.750 ;
        RECT 601.950 95.250 604.050 96.150 ;
        RECT 592.950 92.850 594.750 93.750 ;
        RECT 595.950 91.950 598.050 94.050 ;
        RECT 601.950 91.950 604.050 94.050 ;
        RECT 589.950 88.950 592.050 91.050 ;
        RECT 596.400 88.050 597.450 91.950 ;
        RECT 602.400 88.050 603.450 91.950 ;
        RECT 595.950 85.950 598.050 88.050 ;
        RECT 601.950 85.950 604.050 88.050 ;
        RECT 586.950 73.950 589.050 76.050 ;
        RECT 568.800 65.100 570.900 67.200 ;
        RECT 569.550 61.350 570.750 65.100 ;
        RECT 592.950 64.950 595.050 67.050 ;
        RECT 595.950 64.950 598.050 67.050 ;
        RECT 598.950 64.950 601.050 67.050 ;
        RECT 571.950 62.850 574.050 64.950 ;
        RECT 553.950 58.950 556.050 61.050 ;
        RECT 568.950 59.250 571.050 61.350 ;
        RECT 538.950 50.850 541.050 51.750 ;
        RECT 541.950 49.950 544.050 52.050 ;
        RECT 547.950 50.850 550.050 51.750 ;
        RECT 550.950 49.950 553.050 52.050 ;
        RECT 535.950 40.950 538.050 43.050 ;
        RECT 529.950 37.950 532.050 40.050 ;
        RECT 526.950 25.950 529.050 28.050 ;
        RECT 532.950 25.950 535.050 28.050 ;
        RECT 526.950 22.950 529.050 25.050 ;
        RECT 527.400 18.450 528.450 22.950 ;
        RECT 533.400 22.050 534.450 25.950 ;
        RECT 536.400 25.050 537.450 40.950 ;
        RECT 535.950 22.950 538.050 25.050 ;
        RECT 542.400 22.050 543.450 49.950 ;
        RECT 547.950 22.950 550.050 25.050 ;
        RECT 548.400 22.050 549.450 22.950 ;
        RECT 529.950 20.250 531.750 21.150 ;
        RECT 532.950 19.950 535.050 22.050 ;
        RECT 536.250 20.250 538.050 21.150 ;
        RECT 541.950 19.950 544.050 22.050 ;
        RECT 547.950 19.950 550.050 22.050 ;
        RECT 551.250 20.250 553.050 21.150 ;
        RECT 554.400 19.050 555.450 58.950 ;
        RECT 559.950 56.250 562.050 57.150 ;
        RECT 559.950 52.950 562.050 55.050 ;
        RECT 569.550 45.600 570.750 59.250 ;
        RECT 572.250 45.600 573.450 62.850 ;
        RECT 579.900 62.400 582.000 64.500 ;
        RECT 583.950 62.400 586.050 64.500 ;
        RECT 574.950 59.250 577.050 61.350 ;
        RECT 575.400 45.600 576.600 59.250 ;
        RECT 580.350 53.550 581.550 62.400 ;
        RECT 584.550 56.250 585.750 62.400 ;
        RECT 583.950 54.150 586.050 56.250 ;
        RECT 579.750 51.450 581.850 53.550 ;
        RECT 580.350 45.600 581.550 51.450 ;
        RECT 584.550 45.600 585.750 54.150 ;
        RECT 586.950 50.250 589.050 51.150 ;
        RECT 586.950 46.950 589.050 49.050 ;
        RECT 593.250 46.050 594.450 64.950 ;
        RECT 596.250 60.750 597.450 64.950 ;
        RECT 595.950 58.650 598.050 60.750 ;
        RECT 596.250 46.050 597.450 58.650 ;
        RECT 599.250 46.050 600.450 64.950 ;
        RECT 602.400 61.050 603.450 85.950 ;
        RECT 605.400 67.050 606.450 109.950 ;
        RECT 611.400 106.050 612.450 124.950 ;
        RECT 617.400 112.050 618.450 139.950 ;
        RECT 629.400 139.050 630.450 160.950 ;
        RECT 628.950 136.950 631.050 139.050 ;
        RECT 625.950 130.950 628.050 133.050 ;
        RECT 626.400 130.050 627.450 130.950 ;
        RECT 629.400 130.050 630.450 136.950 ;
        RECT 625.950 127.950 628.050 130.050 ;
        RECT 628.950 127.950 631.050 130.050 ;
        RECT 619.950 125.250 622.050 126.150 ;
        RECT 625.950 125.850 628.050 126.750 ;
        RECT 628.950 125.250 631.050 126.150 ;
        RECT 631.950 124.950 634.050 127.050 ;
        RECT 619.950 121.950 622.050 124.050 ;
        RECT 628.950 121.950 631.050 124.050 ;
        RECT 625.950 118.950 628.050 121.050 ;
        RECT 616.950 109.950 619.050 112.050 ;
        RECT 610.950 103.950 613.050 106.050 ;
        RECT 626.400 94.050 627.450 118.950 ;
        RECT 632.400 100.050 633.450 124.950 ;
        RECT 635.400 121.050 636.450 169.950 ;
        RECT 640.950 166.950 643.050 169.050 ;
        RECT 641.400 166.050 642.450 166.950 ;
        RECT 637.950 164.250 639.750 165.150 ;
        RECT 640.950 163.950 643.050 166.050 ;
        RECT 644.250 164.250 646.050 165.150 ;
        RECT 637.950 160.950 640.050 163.050 ;
        RECT 641.250 161.850 642.750 162.750 ;
        RECT 643.950 160.950 646.050 163.050 ;
        RECT 640.950 157.950 643.050 160.050 ;
        RECT 641.400 130.050 642.450 157.950 ;
        RECT 644.400 145.050 645.450 160.950 ;
        RECT 643.950 142.950 646.050 145.050 ;
        RECT 650.400 133.050 651.450 235.950 ;
        RECT 652.950 232.950 655.050 235.050 ;
        RECT 655.950 232.950 658.050 235.050 ;
        RECT 659.400 234.450 660.450 241.950 ;
        RECT 662.400 237.450 663.450 262.950 ;
        RECT 671.400 250.050 672.450 265.950 ;
        RECT 674.400 265.050 675.450 304.950 ;
        RECT 679.950 301.950 682.050 304.050 ;
        RECT 676.950 269.250 679.050 270.150 ;
        RECT 676.950 265.950 679.050 268.050 ;
        RECT 673.950 262.950 676.050 265.050 ;
        RECT 677.400 262.050 678.450 265.950 ;
        RECT 676.950 259.950 679.050 262.050 ;
        RECT 680.400 258.450 681.450 301.950 ;
        RECT 689.400 295.050 690.450 304.950 ;
        RECT 682.950 292.950 685.050 295.050 ;
        RECT 688.950 292.950 691.050 295.050 ;
        RECT 683.400 274.050 684.450 292.950 ;
        RECT 692.400 283.050 693.450 319.950 ;
        RECT 698.400 313.050 699.450 329.400 ;
        RECT 700.950 313.950 703.050 316.050 ;
        RECT 697.950 310.950 700.050 313.050 ;
        RECT 698.400 307.050 699.450 310.950 ;
        RECT 701.400 310.050 702.450 313.950 ;
        RECT 704.400 313.050 705.450 334.950 ;
        RECT 707.250 333.600 708.450 342.150 ;
        RECT 711.450 341.550 712.650 350.400 ;
        RECT 715.950 347.250 718.050 349.350 ;
        RECT 711.150 339.450 713.250 341.550 ;
        RECT 711.450 333.600 712.650 339.450 ;
        RECT 716.400 333.600 717.600 347.250 ;
        RECT 719.550 333.600 720.750 350.850 ;
        RECT 722.250 349.350 723.450 353.100 ;
        RECT 721.950 347.250 724.050 349.350 ;
        RECT 728.400 349.050 729.450 376.950 ;
        RECT 734.250 372.600 735.450 378.750 ;
        RECT 738.450 372.600 739.650 381.450 ;
        RECT 743.400 375.750 744.600 389.400 ;
        RECT 742.950 373.650 745.050 375.750 ;
        RECT 733.950 370.500 736.050 372.600 ;
        RECT 738.000 370.500 740.100 372.600 ;
        RECT 746.550 372.150 747.750 389.400 ;
        RECT 749.250 375.750 750.450 389.400 ;
        RECT 752.400 376.050 753.450 409.950 ;
        RECT 758.400 391.050 759.450 409.950 ;
        RECT 757.950 388.950 760.050 391.050 ;
        RECT 755.400 386.400 762.450 387.450 ;
        RECT 755.400 385.050 756.450 386.400 ;
        RECT 761.400 385.050 762.450 386.400 ;
        RECT 754.950 382.950 757.050 385.050 ;
        RECT 757.950 382.950 760.050 385.050 ;
        RECT 760.950 382.950 763.050 385.050 ;
        RECT 758.400 382.050 759.450 382.950 ;
        RECT 754.950 379.950 757.050 382.050 ;
        RECT 757.950 379.950 760.050 382.050 ;
        RECT 748.950 373.650 751.050 375.750 ;
        RECT 751.950 373.950 754.050 376.050 ;
        RECT 745.950 370.050 748.050 372.150 ;
        RECT 749.250 369.900 750.450 373.650 ;
        RECT 749.100 367.800 751.200 369.900 ;
        RECT 751.950 364.950 754.050 367.050 ;
        RECT 739.950 358.950 742.050 361.050 ;
        RECT 736.950 352.950 739.050 355.050 ;
        RECT 722.250 333.600 723.450 347.250 ;
        RECT 727.950 346.950 730.050 349.050 ;
        RECT 706.950 331.500 709.050 333.600 ;
        RECT 711.150 331.500 713.250 333.600 ;
        RECT 715.950 331.500 718.050 333.600 ;
        RECT 718.950 331.500 721.050 333.600 ;
        RECT 721.950 331.500 724.050 333.600 ;
        RECT 718.950 319.950 721.050 322.050 ;
        RECT 715.950 316.950 718.050 319.050 ;
        RECT 709.950 313.950 712.050 316.050 ;
        RECT 710.400 313.050 711.450 313.950 ;
        RECT 703.950 310.950 706.050 313.050 ;
        RECT 707.250 311.250 708.750 312.150 ;
        RECT 709.950 310.950 712.050 313.050 ;
        RECT 700.950 307.950 703.050 310.050 ;
        RECT 704.250 308.850 705.750 309.750 ;
        RECT 706.950 307.950 709.050 310.050 ;
        RECT 710.250 308.850 712.050 309.750 ;
        RECT 712.950 307.950 715.050 310.050 ;
        RECT 707.400 307.050 708.450 307.950 ;
        RECT 697.950 304.950 700.050 307.050 ;
        RECT 700.950 305.850 703.050 306.750 ;
        RECT 706.950 304.950 709.050 307.050 ;
        RECT 694.950 301.950 697.050 304.050 ;
        RECT 691.950 280.950 694.050 283.050 ;
        RECT 688.950 275.250 691.050 276.150 ;
        RECT 695.400 274.050 696.450 301.950 ;
        RECT 713.400 301.050 714.450 307.950 ;
        RECT 712.950 298.950 715.050 301.050 ;
        RECT 709.950 289.950 712.050 292.050 ;
        RECT 700.950 286.950 703.050 289.050 ;
        RECT 697.950 283.950 700.050 286.050 ;
        RECT 682.950 271.950 685.050 274.050 ;
        RECT 685.950 272.250 687.750 273.150 ;
        RECT 688.950 271.950 691.050 274.050 ;
        RECT 692.250 272.250 693.750 273.150 ;
        RECT 694.950 271.950 697.050 274.050 ;
        RECT 685.950 270.450 688.050 271.050 ;
        RECT 683.400 269.400 688.050 270.450 ;
        RECT 683.400 262.050 684.450 269.400 ;
        RECT 685.950 268.950 688.050 269.400 ;
        RECT 688.950 268.950 691.050 271.050 ;
        RECT 691.950 268.950 694.050 271.050 ;
        RECT 695.250 269.850 697.050 270.750 ;
        RECT 685.950 265.950 688.050 268.050 ;
        RECT 682.950 259.950 685.050 262.050 ;
        RECT 677.400 257.400 681.450 258.450 ;
        RECT 670.950 247.950 673.050 250.050 ;
        RECT 667.950 241.950 670.050 244.050 ;
        RECT 677.400 241.050 678.450 257.400 ;
        RECT 664.950 239.250 667.050 240.150 ;
        RECT 667.950 239.850 670.050 240.750 ;
        RECT 670.950 238.950 673.050 241.050 ;
        RECT 674.250 239.250 675.750 240.150 ;
        RECT 676.950 238.950 679.050 241.050 ;
        RECT 664.950 237.450 667.050 238.050 ;
        RECT 662.400 236.400 667.050 237.450 ;
        RECT 664.950 235.950 667.050 236.400 ;
        RECT 667.950 235.950 670.050 238.050 ;
        RECT 670.950 236.850 672.750 237.750 ;
        RECT 673.950 235.950 676.050 238.050 ;
        RECT 677.250 236.850 678.750 237.750 ;
        RECT 679.950 235.950 682.050 238.050 ;
        RECT 659.400 233.400 663.450 234.450 ;
        RECT 653.400 199.050 654.450 232.950 ;
        RECT 652.950 196.950 655.050 199.050 ;
        RECT 652.950 193.950 655.050 196.050 ;
        RECT 653.400 157.050 654.450 193.950 ;
        RECT 656.400 169.050 657.450 232.950 ;
        RECT 662.400 226.050 663.450 233.400 ;
        RECT 661.950 223.950 664.050 226.050 ;
        RECT 662.400 202.050 663.450 223.950 ;
        RECT 668.400 211.050 669.450 235.950 ;
        RECT 674.400 229.050 675.450 235.950 ;
        RECT 679.950 233.850 682.050 234.750 ;
        RECT 673.950 226.950 676.050 229.050 ;
        RECT 683.400 226.050 684.450 259.950 ;
        RECT 686.400 238.050 687.450 265.950 ;
        RECT 689.400 262.050 690.450 268.950 ;
        RECT 688.950 259.950 691.050 262.050 ;
        RECT 692.400 250.050 693.450 268.950 ;
        RECT 698.400 262.050 699.450 283.950 ;
        RECT 701.400 271.050 702.450 286.950 ;
        RECT 706.950 274.950 709.050 277.050 ;
        RECT 703.950 271.950 706.050 274.050 ;
        RECT 704.400 271.050 705.450 271.950 ;
        RECT 700.950 268.950 703.050 271.050 ;
        RECT 703.950 268.950 706.050 271.050 ;
        RECT 700.950 266.250 703.050 267.150 ;
        RECT 703.950 266.850 706.050 267.750 ;
        RECT 700.950 262.950 703.050 265.050 ;
        RECT 694.950 259.950 697.050 262.050 ;
        RECT 697.950 259.950 700.050 262.050 ;
        RECT 691.950 247.950 694.050 250.050 ;
        RECT 692.400 247.050 693.450 247.950 ;
        RECT 691.950 244.950 694.050 247.050 ;
        RECT 695.400 244.050 696.450 259.950 ;
        RECT 701.400 253.050 702.450 262.950 ;
        RECT 700.950 250.950 703.050 253.050 ;
        RECT 700.950 247.950 703.050 250.050 ;
        RECT 694.950 241.950 697.050 244.050 ;
        RECT 691.950 240.450 694.050 241.050 ;
        RECT 689.400 239.400 694.050 240.450 ;
        RECT 695.250 239.850 696.750 240.750 ;
        RECT 685.950 235.950 688.050 238.050 ;
        RECT 670.950 223.950 673.050 226.050 ;
        RECT 682.950 223.950 685.050 226.050 ;
        RECT 664.950 208.950 667.050 211.050 ;
        RECT 667.950 208.950 670.050 211.050 ;
        RECT 661.950 199.950 664.050 202.050 ;
        RECT 665.400 199.050 666.450 208.950 ;
        RECT 661.950 197.250 664.050 198.150 ;
        RECT 664.950 196.950 667.050 199.050 ;
        RECT 667.950 197.250 670.050 198.150 ;
        RECT 661.950 193.950 664.050 196.050 ;
        RECT 665.250 194.250 666.750 195.150 ;
        RECT 667.950 193.950 670.050 196.050 ;
        RECT 664.950 190.950 667.050 193.050 ;
        RECT 658.950 187.950 661.050 190.050 ;
        RECT 659.400 172.050 660.450 187.950 ;
        RECT 664.950 184.950 667.050 187.050 ;
        RECT 661.950 172.950 664.050 175.050 ;
        RECT 658.950 169.950 661.050 172.050 ;
        RECT 662.400 169.050 663.450 172.950 ;
        RECT 655.950 166.950 658.050 169.050 ;
        RECT 659.250 167.850 660.750 168.750 ;
        RECT 661.950 166.950 664.050 169.050 ;
        RECT 655.950 164.850 658.050 165.750 ;
        RECT 661.950 164.850 664.050 165.750 ;
        RECT 652.950 154.950 655.050 157.050 ;
        RECT 665.400 151.050 666.450 184.950 ;
        RECT 671.400 169.050 672.450 223.950 ;
        RECT 673.950 208.950 676.050 211.050 ;
        RECT 674.400 208.050 675.450 208.950 ;
        RECT 673.950 205.950 676.050 208.050 ;
        RECT 674.400 199.050 675.450 205.950 ;
        RECT 676.950 199.950 679.050 202.050 ;
        RECT 673.950 196.950 676.050 199.050 ;
        RECT 673.950 194.850 676.050 195.750 ;
        RECT 677.400 184.050 678.450 199.950 ;
        RECT 679.950 196.950 682.050 199.050 ;
        RECT 679.950 194.850 682.050 195.750 ;
        RECT 686.400 187.050 687.450 235.950 ;
        RECT 689.400 229.050 690.450 239.400 ;
        RECT 691.950 238.950 694.050 239.400 ;
        RECT 697.950 238.950 700.050 241.050 ;
        RECT 691.950 236.850 694.050 237.750 ;
        RECT 697.950 236.850 700.050 237.750 ;
        RECT 688.950 226.950 691.050 229.050 ;
        RECT 691.950 197.250 694.050 198.150 ;
        RECT 697.950 197.250 700.050 198.150 ;
        RECT 691.950 193.950 694.050 196.050 ;
        RECT 695.250 194.250 696.750 195.150 ;
        RECT 697.950 193.950 700.050 196.050 ;
        RECT 692.400 187.050 693.450 193.950 ;
        RECT 694.950 190.950 697.050 193.050 ;
        RECT 698.400 190.050 699.450 193.950 ;
        RECT 697.950 187.950 700.050 190.050 ;
        RECT 685.950 184.950 688.050 187.050 ;
        RECT 691.950 184.950 694.050 187.050 ;
        RECT 676.950 181.950 679.050 184.050 ;
        RECT 676.950 178.950 679.050 181.050 ;
        RECT 670.950 166.950 673.050 169.050 ;
        RECT 673.950 165.450 676.050 166.050 ;
        RECT 671.400 164.400 676.050 165.450 ;
        RECT 652.950 148.950 655.050 151.050 ;
        RECT 664.950 148.950 667.050 151.050 ;
        RECT 646.950 131.250 649.050 132.150 ;
        RECT 649.950 130.950 652.050 133.050 ;
        RECT 640.950 127.950 643.050 130.050 ;
        RECT 644.250 128.250 645.750 129.150 ;
        RECT 646.950 127.950 649.050 130.050 ;
        RECT 650.250 128.250 652.050 129.150 ;
        RECT 640.950 125.850 642.750 126.750 ;
        RECT 643.950 124.950 646.050 127.050 ;
        RECT 634.950 118.950 637.050 121.050 ;
        RECT 644.400 103.050 645.450 124.950 ;
        RECT 647.400 121.050 648.450 127.950 ;
        RECT 649.950 124.950 652.050 127.050 ;
        RECT 650.400 124.050 651.450 124.950 ;
        RECT 649.950 121.950 652.050 124.050 ;
        RECT 646.950 118.950 649.050 121.050 ;
        RECT 643.950 100.950 646.050 103.050 ;
        RECT 631.950 97.950 634.050 100.050 ;
        RECT 643.950 97.950 646.050 100.050 ;
        RECT 628.950 94.950 631.050 97.050 ;
        RECT 634.950 94.950 637.050 97.050 ;
        RECT 640.950 95.250 643.050 96.150 ;
        RECT 643.950 95.850 646.050 96.750 ;
        RECT 646.950 95.250 648.750 96.150 ;
        RECT 649.950 94.950 652.050 97.050 ;
        RECT 629.400 94.050 630.450 94.950 ;
        RECT 607.950 92.250 609.750 93.150 ;
        RECT 610.950 91.950 613.050 94.050 ;
        RECT 619.950 93.450 622.050 94.050 ;
        RECT 622.950 93.450 625.050 94.050 ;
        RECT 614.250 92.250 616.050 93.150 ;
        RECT 619.950 92.400 625.050 93.450 ;
        RECT 619.950 91.950 622.050 92.400 ;
        RECT 622.950 91.950 625.050 92.400 ;
        RECT 625.950 91.950 628.050 94.050 ;
        RECT 628.950 91.950 631.050 94.050 ;
        RECT 632.250 92.250 634.050 93.150 ;
        RECT 607.950 88.950 610.050 91.050 ;
        RECT 611.250 89.850 612.750 90.750 ;
        RECT 613.950 88.950 616.050 91.050 ;
        RECT 622.950 89.850 624.750 90.750 ;
        RECT 625.950 88.950 628.050 91.050 ;
        RECT 629.250 89.850 630.750 90.750 ;
        RECT 631.950 88.950 634.050 91.050 ;
        RECT 608.400 88.050 609.450 88.950 ;
        RECT 632.400 88.050 633.450 88.950 ;
        RECT 607.950 85.950 610.050 88.050 ;
        RECT 625.950 86.850 628.050 87.750 ;
        RECT 631.950 85.950 634.050 88.050 ;
        RECT 635.400 85.050 636.450 94.950 ;
        RECT 640.950 91.950 643.050 94.050 ;
        RECT 646.950 91.950 649.050 94.050 ;
        RECT 650.250 92.850 652.050 93.750 ;
        RECT 634.950 82.950 637.050 85.050 ;
        RECT 647.400 76.050 648.450 91.950 ;
        RECT 653.400 91.050 654.450 148.950 ;
        RECT 664.950 139.950 667.050 142.050 ;
        RECT 658.950 131.250 661.050 132.150 ;
        RECT 665.400 130.050 666.450 139.950 ;
        RECT 655.950 128.250 657.750 129.150 ;
        RECT 658.950 127.950 661.050 130.050 ;
        RECT 662.250 128.250 663.750 129.150 ;
        RECT 664.950 127.950 667.050 130.050 ;
        RECT 655.950 124.950 658.050 127.050 ;
        RECT 656.400 115.050 657.450 124.950 ;
        RECT 659.400 124.050 660.450 127.950 ;
        RECT 671.400 127.050 672.450 164.400 ;
        RECT 673.950 163.950 676.050 164.400 ;
        RECT 677.400 163.050 678.450 178.950 ;
        RECT 701.400 178.050 702.450 247.950 ;
        RECT 707.400 244.050 708.450 274.950 ;
        RECT 710.400 259.050 711.450 289.950 ;
        RECT 709.950 256.950 712.050 259.050 ;
        RECT 713.400 247.050 714.450 298.950 ;
        RECT 716.400 280.050 717.450 316.950 ;
        RECT 719.400 313.050 720.450 319.950 ;
        RECT 718.950 310.950 721.050 313.050 ;
        RECT 724.950 310.950 727.050 313.050 ;
        RECT 718.950 308.850 721.050 309.750 ;
        RECT 724.950 308.850 727.050 309.750 ;
        RECT 728.400 298.050 729.450 346.950 ;
        RECT 730.950 344.250 733.050 345.150 ;
        RECT 730.950 340.950 733.050 343.050 ;
        RECT 731.400 337.050 732.450 340.950 ;
        RECT 730.950 334.950 733.050 337.050 ;
        RECT 727.950 295.950 730.050 298.050 ;
        RECT 724.950 292.950 727.050 295.050 ;
        RECT 715.950 277.950 718.050 280.050 ;
        RECT 718.950 275.250 721.050 276.150 ;
        RECT 725.400 274.050 726.450 292.950 ;
        RECT 715.950 272.250 717.750 273.150 ;
        RECT 718.950 271.950 721.050 274.050 ;
        RECT 722.250 272.250 723.750 273.150 ;
        RECT 724.950 271.950 727.050 274.050 ;
        RECT 727.950 271.950 730.050 274.050 ;
        RECT 715.950 268.950 718.050 271.050 ;
        RECT 721.950 268.950 724.050 271.050 ;
        RECT 725.250 269.850 727.050 270.750 ;
        RECT 716.400 268.050 717.450 268.950 ;
        RECT 715.950 265.950 718.050 268.050 ;
        RECT 722.400 267.450 723.450 268.950 ;
        RECT 728.400 267.450 729.450 271.950 ;
        RECT 722.400 266.400 729.450 267.450 ;
        RECT 712.950 244.950 715.050 247.050 ;
        RECT 718.950 244.950 721.050 247.050 ;
        RECT 706.950 241.950 709.050 244.050 ;
        RECT 707.400 235.050 708.450 241.950 ;
        RECT 712.950 238.950 715.050 241.050 ;
        RECT 713.400 238.050 714.450 238.950 ;
        RECT 709.950 236.250 711.750 237.150 ;
        RECT 712.950 235.950 715.050 238.050 ;
        RECT 716.250 236.250 718.050 237.150 ;
        RECT 706.950 232.950 709.050 235.050 ;
        RECT 709.950 232.950 712.050 235.050 ;
        RECT 713.250 233.850 714.750 234.750 ;
        RECT 715.950 232.950 718.050 235.050 ;
        RECT 710.400 232.050 711.450 232.950 ;
        RECT 706.950 229.950 709.050 232.050 ;
        RECT 709.950 229.950 712.050 232.050 ;
        RECT 707.400 226.050 708.450 229.950 ;
        RECT 706.950 223.950 709.050 226.050 ;
        RECT 706.950 220.950 709.050 223.050 ;
        RECT 707.400 199.050 708.450 220.950 ;
        RECT 706.950 196.950 709.050 199.050 ;
        RECT 710.400 196.050 711.450 229.950 ;
        RECT 712.950 199.950 715.050 202.050 ;
        RECT 703.950 194.250 706.050 195.150 ;
        RECT 706.950 194.850 709.050 195.750 ;
        RECT 709.950 193.950 712.050 196.050 ;
        RECT 713.400 193.050 714.450 199.950 ;
        RECT 719.400 199.050 720.450 244.950 ;
        RECT 725.400 244.050 726.450 266.400 ;
        RECT 727.950 262.950 730.050 265.050 ;
        RECT 728.400 253.050 729.450 262.950 ;
        RECT 727.950 250.950 730.050 253.050 ;
        RECT 731.400 247.050 732.450 334.950 ;
        RECT 737.400 322.050 738.450 352.950 ;
        RECT 736.950 319.950 739.050 322.050 ;
        RECT 736.950 316.950 739.050 319.050 ;
        RECT 733.950 313.950 736.050 316.050 ;
        RECT 734.400 286.050 735.450 313.950 ;
        RECT 733.950 283.950 736.050 286.050 ;
        RECT 733.950 277.950 736.050 280.050 ;
        RECT 734.400 256.050 735.450 277.950 ;
        RECT 737.400 277.050 738.450 316.950 ;
        RECT 740.400 315.450 741.450 358.950 ;
        RECT 742.950 340.950 745.050 343.050 ;
        RECT 742.950 338.850 745.050 339.750 ;
        RECT 752.400 337.050 753.450 364.950 ;
        RECT 751.950 334.950 754.050 337.050 ;
        RECT 755.400 322.050 756.450 379.950 ;
        RECT 757.950 377.850 760.050 378.750 ;
        RECT 764.400 372.450 765.450 409.950 ;
        RECT 761.400 371.400 765.450 372.450 ;
        RECT 761.400 343.050 762.450 371.400 ;
        RECT 767.400 343.050 768.450 412.950 ;
        RECT 772.950 410.850 775.050 411.750 ;
        RECT 775.950 410.250 778.050 411.150 ;
        RECT 775.950 408.450 778.050 409.050 ;
        RECT 779.400 408.450 780.450 413.400 ;
        RECT 781.950 412.950 784.050 413.400 ;
        RECT 785.400 412.050 786.450 545.400 ;
        RECT 787.950 526.950 790.050 529.050 ;
        RECT 790.950 527.250 793.050 528.150 ;
        RECT 788.400 523.050 789.450 526.950 ;
        RECT 790.950 523.950 793.050 526.050 ;
        RECT 787.950 520.950 790.050 523.050 ;
        RECT 787.950 514.950 790.050 517.050 ;
        RECT 788.400 412.050 789.450 514.950 ;
        RECT 791.400 511.050 792.450 523.950 ;
        RECT 794.400 517.050 795.450 592.950 ;
        RECT 797.400 574.050 798.450 610.950 ;
        RECT 800.400 589.050 801.450 613.950 ;
        RECT 808.950 607.950 811.050 610.050 ;
        RECT 802.950 604.950 805.050 607.050 ;
        RECT 803.400 601.050 804.450 604.950 ;
        RECT 805.950 601.950 808.050 604.050 ;
        RECT 809.400 601.050 810.450 607.950 ;
        RECT 802.950 598.950 805.050 601.050 ;
        RECT 806.250 599.850 807.750 600.750 ;
        RECT 808.950 598.950 811.050 601.050 ;
        RECT 802.950 596.850 805.050 597.750 ;
        RECT 808.950 596.850 811.050 597.750 ;
        RECT 812.400 595.050 813.450 613.950 ;
        RECT 815.400 598.050 816.450 661.950 ;
        RECT 827.400 655.050 828.450 724.950 ;
        RECT 830.400 709.050 831.450 748.950 ;
        RECT 850.950 745.950 853.050 748.050 ;
        RECT 851.400 745.050 852.450 745.950 ;
        RECT 854.400 745.050 855.450 772.950 ;
        RECT 856.950 745.950 859.050 748.050 ;
        RECT 844.950 744.450 847.050 745.050 ;
        RECT 842.400 743.400 847.050 744.450 ;
        RECT 838.950 740.250 841.050 741.150 ;
        RECT 832.950 737.850 835.050 738.750 ;
        RECT 838.950 738.450 841.050 739.050 ;
        RECT 836.400 737.400 841.050 738.450 ;
        RECT 829.950 706.950 832.050 709.050 ;
        RECT 836.400 706.050 837.450 737.400 ;
        RECT 838.950 736.950 841.050 737.400 ;
        RECT 842.400 736.050 843.450 743.400 ;
        RECT 844.950 742.950 847.050 743.400 ;
        RECT 848.250 743.250 849.750 744.150 ;
        RECT 850.950 742.950 853.050 745.050 ;
        RECT 853.950 742.950 856.050 745.050 ;
        RECT 854.400 742.050 855.450 742.950 ;
        RECT 844.950 740.850 846.750 741.750 ;
        RECT 847.950 739.950 850.050 742.050 ;
        RECT 851.250 740.850 852.750 741.750 ;
        RECT 853.950 739.950 856.050 742.050 ;
        RECT 841.950 733.950 844.050 736.050 ;
        RECT 848.400 727.050 849.450 739.950 ;
        RECT 853.950 737.850 856.050 738.750 ;
        RECT 853.950 733.950 856.050 736.050 ;
        RECT 847.950 724.950 850.050 727.050 ;
        RECT 835.950 705.450 838.050 706.050 ;
        RECT 829.950 704.250 832.050 705.150 ;
        RECT 833.400 704.400 838.050 705.450 ;
        RECT 833.400 688.050 834.450 704.400 ;
        RECT 835.950 703.950 838.050 704.400 ;
        RECT 835.950 701.850 838.050 702.750 ;
        RECT 841.950 700.950 844.050 703.050 ;
        RECT 847.950 700.950 850.050 703.050 ;
        RECT 832.950 685.950 835.050 688.050 ;
        RECT 838.950 673.950 841.050 676.050 ;
        RECT 839.400 673.050 840.450 673.950 ;
        RECT 829.950 672.450 832.050 673.050 ;
        RECT 832.950 672.450 835.050 673.050 ;
        RECT 829.950 671.400 835.050 672.450 ;
        RECT 829.950 670.950 832.050 671.400 ;
        RECT 832.950 670.950 835.050 671.400 ;
        RECT 836.250 671.250 837.750 672.150 ;
        RECT 838.950 670.950 841.050 673.050 ;
        RECT 826.950 652.950 829.050 655.050 ;
        RECT 817.950 640.950 820.050 643.050 ;
        RECT 820.950 640.950 823.050 643.050 ;
        RECT 823.950 640.950 826.050 643.050 ;
        RECT 830.400 642.450 831.450 670.950 ;
        RECT 842.400 670.050 843.450 700.950 ;
        RECT 847.950 698.850 850.050 699.750 ;
        RECT 850.950 698.250 853.050 699.150 ;
        RECT 844.950 694.950 847.050 697.050 ;
        RECT 850.950 694.950 853.050 697.050 ;
        RECT 832.950 668.850 834.750 669.750 ;
        RECT 835.950 667.950 838.050 670.050 ;
        RECT 839.250 668.850 840.750 669.750 ;
        RECT 841.950 667.950 844.050 670.050 ;
        RECT 836.400 667.050 837.450 667.950 ;
        RECT 835.950 664.950 838.050 667.050 ;
        RECT 841.950 665.850 844.050 666.750 ;
        RECT 841.950 661.950 844.050 664.050 ;
        RECT 830.400 641.400 834.450 642.450 ;
        RECT 818.250 622.050 819.450 640.950 ;
        RECT 821.250 636.750 822.450 640.950 ;
        RECT 820.950 634.650 823.050 636.750 ;
        RECT 821.250 622.050 822.450 634.650 ;
        RECT 824.250 622.050 825.450 640.950 ;
        RECT 829.950 632.250 832.050 633.150 ;
        RECT 817.950 619.950 820.050 622.050 ;
        RECT 820.950 619.950 823.050 622.050 ;
        RECT 823.950 619.950 826.050 622.050 ;
        RECT 823.950 616.950 826.050 619.050 ;
        RECT 824.400 601.050 825.450 616.950 ;
        RECT 829.950 607.950 832.050 610.050 ;
        RECT 817.950 598.950 820.050 601.050 ;
        RECT 821.250 599.250 822.750 600.150 ;
        RECT 823.950 598.950 826.050 601.050 ;
        RECT 826.950 598.950 829.050 601.050 ;
        RECT 827.400 598.050 828.450 598.950 ;
        RECT 814.950 595.950 817.050 598.050 ;
        RECT 817.950 596.850 819.750 597.750 ;
        RECT 820.950 595.950 823.050 598.050 ;
        RECT 824.250 596.850 825.750 597.750 ;
        RECT 826.950 595.950 829.050 598.050 ;
        RECT 811.950 592.950 814.050 595.050 ;
        RECT 826.950 593.850 829.050 594.750 ;
        RECT 799.950 586.950 802.050 589.050 ;
        RECT 796.950 571.950 799.050 574.050 ;
        RECT 830.400 573.450 831.450 607.950 ;
        RECT 833.400 607.050 834.450 641.400 ;
        RECT 838.950 634.950 841.050 637.050 ;
        RECT 835.950 631.950 838.050 634.050 ;
        RECT 835.950 629.850 838.050 630.750 ;
        RECT 832.950 604.950 835.050 607.050 ;
        RECT 835.950 604.950 838.050 607.050 ;
        RECT 836.400 601.050 837.450 604.950 ;
        RECT 839.400 604.050 840.450 634.950 ;
        RECT 842.400 607.050 843.450 661.950 ;
        RECT 845.400 627.450 846.450 694.950 ;
        RECT 854.400 664.050 855.450 733.950 ;
        RECT 853.950 661.950 856.050 664.050 ;
        RECT 857.400 636.450 858.450 745.950 ;
        RECT 862.950 700.950 865.050 703.050 ;
        RECT 857.400 635.400 861.450 636.450 ;
        RECT 847.950 631.950 850.050 634.050 ;
        RECT 853.950 633.450 856.050 634.050 ;
        RECT 851.250 632.250 852.750 633.150 ;
        RECT 853.950 632.400 858.450 633.450 ;
        RECT 853.950 631.950 856.050 632.400 ;
        RECT 847.950 629.850 849.750 630.750 ;
        RECT 850.950 628.950 853.050 631.050 ;
        RECT 854.250 629.850 856.050 630.750 ;
        RECT 845.400 626.400 849.450 627.450 ;
        RECT 841.950 604.950 844.050 607.050 ;
        RECT 838.950 601.950 841.050 604.050 ;
        RECT 844.950 601.950 847.050 604.050 ;
        RECT 835.950 598.950 838.050 601.050 ;
        RECT 839.250 599.250 840.750 600.150 ;
        RECT 841.950 598.950 844.050 601.050 ;
        RECT 845.400 598.050 846.450 601.950 ;
        RECT 835.950 596.850 837.750 597.750 ;
        RECT 838.950 595.950 841.050 598.050 ;
        RECT 842.250 596.850 843.750 597.750 ;
        RECT 844.950 595.950 847.050 598.050 ;
        RECT 839.400 592.050 840.450 595.950 ;
        RECT 844.950 593.850 847.050 594.750 ;
        RECT 838.950 589.950 841.050 592.050 ;
        RECT 848.400 591.450 849.450 626.400 ;
        RECT 851.400 610.050 852.450 628.950 ;
        RECT 857.400 627.450 858.450 632.400 ;
        RECT 854.400 626.400 858.450 627.450 ;
        RECT 850.950 607.950 853.050 610.050 ;
        RECT 850.950 604.950 853.050 607.050 ;
        RECT 845.400 590.400 849.450 591.450 ;
        RECT 830.400 572.400 834.450 573.450 ;
        RECT 799.800 569.100 801.900 571.200 ;
        RECT 800.550 565.350 801.750 569.100 ;
        RECT 823.950 568.950 826.050 571.050 ;
        RECT 826.950 568.950 829.050 571.050 ;
        RECT 829.950 568.950 832.050 571.050 ;
        RECT 802.950 566.850 805.050 568.950 ;
        RECT 799.950 563.250 802.050 565.350 ;
        RECT 800.550 549.600 801.750 563.250 ;
        RECT 803.250 549.600 804.450 566.850 ;
        RECT 810.900 566.400 813.000 568.500 ;
        RECT 814.950 566.400 817.050 568.500 ;
        RECT 805.950 563.250 808.050 565.350 ;
        RECT 806.400 549.600 807.600 563.250 ;
        RECT 811.350 557.550 812.550 566.400 ;
        RECT 815.550 560.250 816.750 566.400 ;
        RECT 814.950 558.150 817.050 560.250 ;
        RECT 810.750 555.450 812.850 557.550 ;
        RECT 811.350 549.600 812.550 555.450 ;
        RECT 815.550 549.600 816.750 558.150 ;
        RECT 817.950 554.250 820.050 555.150 ;
        RECT 817.950 550.950 820.050 553.050 ;
        RECT 799.950 547.500 802.050 549.600 ;
        RECT 802.950 547.500 805.050 549.600 ;
        RECT 805.950 547.500 808.050 549.600 ;
        RECT 810.750 547.500 812.850 549.600 ;
        RECT 814.950 547.500 817.050 549.600 ;
        RECT 818.400 547.050 819.450 550.950 ;
        RECT 824.250 550.050 825.450 568.950 ;
        RECT 827.250 564.750 828.450 568.950 ;
        RECT 826.950 562.650 829.050 564.750 ;
        RECT 827.250 550.050 828.450 562.650 ;
        RECT 830.250 550.050 831.450 568.950 ;
        RECT 823.950 547.950 826.050 550.050 ;
        RECT 826.950 547.950 829.050 550.050 ;
        RECT 829.950 547.950 832.050 550.050 ;
        RECT 817.950 544.950 820.050 547.050 ;
        RECT 811.950 533.400 814.050 535.500 ;
        RECT 814.950 533.400 817.050 535.500 ;
        RECT 817.950 533.400 820.050 535.500 ;
        RECT 822.750 533.400 824.850 535.500 ;
        RECT 826.950 533.400 829.050 535.500 ;
        RECT 796.950 523.950 799.050 526.050 ;
        RECT 802.950 523.950 805.050 526.050 ;
        RECT 793.950 514.950 796.050 517.050 ;
        RECT 790.950 508.950 793.050 511.050 ;
        RECT 793.950 488.250 796.050 489.150 ;
        RECT 793.950 486.450 796.050 487.050 ;
        RECT 797.400 486.450 798.450 523.950 ;
        RECT 802.950 521.850 805.050 522.750 ;
        RECT 812.550 519.750 813.750 533.400 ;
        RECT 811.950 517.650 814.050 519.750 ;
        RECT 812.550 513.900 813.750 517.650 ;
        RECT 815.250 516.150 816.450 533.400 ;
        RECT 818.400 519.750 819.600 533.400 ;
        RECT 823.350 527.550 824.550 533.400 ;
        RECT 822.750 525.450 824.850 527.550 ;
        RECT 817.950 517.650 820.050 519.750 ;
        RECT 823.350 516.600 824.550 525.450 ;
        RECT 827.550 524.850 828.750 533.400 ;
        RECT 829.950 529.950 832.050 532.050 ;
        RECT 829.950 527.850 832.050 528.750 ;
        RECT 826.950 522.750 829.050 524.850 ;
        RECT 827.550 516.600 828.750 522.750 ;
        RECT 814.950 514.050 817.050 516.150 ;
        RECT 822.900 514.500 825.000 516.600 ;
        RECT 826.950 514.500 829.050 516.600 ;
        RECT 811.800 511.800 813.900 513.900 ;
        RECT 833.400 502.050 834.450 572.400 ;
        RECT 841.950 562.950 844.050 565.050 ;
        RECT 842.400 562.050 843.450 562.950 ;
        RECT 835.950 560.250 838.050 561.150 ;
        RECT 841.950 559.950 844.050 562.050 ;
        RECT 841.950 557.850 844.050 558.750 ;
        RECT 835.950 532.950 838.050 535.050 ;
        RECT 838.950 532.950 841.050 535.050 ;
        RECT 841.950 532.950 844.050 535.050 ;
        RECT 836.250 514.050 837.450 532.950 ;
        RECT 839.250 520.350 840.450 532.950 ;
        RECT 838.950 518.250 841.050 520.350 ;
        RECT 839.250 514.050 840.450 518.250 ;
        RECT 842.250 514.050 843.450 532.950 ;
        RECT 835.950 511.950 838.050 514.050 ;
        RECT 838.950 511.950 841.050 514.050 ;
        RECT 841.950 511.950 844.050 514.050 ;
        RECT 841.950 508.950 844.050 511.050 ;
        RECT 823.950 499.950 826.050 502.050 ;
        RECT 832.950 499.950 835.050 502.050 ;
        RECT 802.800 497.100 804.900 499.200 ;
        RECT 803.550 493.350 804.750 497.100 ;
        RECT 805.950 494.850 808.050 496.950 ;
        RECT 802.950 491.250 805.050 493.350 ;
        RECT 793.950 485.400 798.450 486.450 ;
        RECT 793.950 484.950 796.050 485.400 ;
        RECT 790.950 453.450 793.050 454.050 ;
        RECT 794.400 453.450 795.450 484.950 ;
        RECT 803.550 477.600 804.750 491.250 ;
        RECT 806.250 477.600 807.450 494.850 ;
        RECT 813.900 494.400 816.000 496.500 ;
        RECT 817.950 494.400 820.050 496.500 ;
        RECT 808.950 491.250 811.050 493.350 ;
        RECT 809.400 477.600 810.600 491.250 ;
        RECT 814.350 485.550 815.550 494.400 ;
        RECT 818.550 488.250 819.750 494.400 ;
        RECT 817.950 486.150 820.050 488.250 ;
        RECT 813.750 483.450 815.850 485.550 ;
        RECT 814.350 477.600 815.550 483.450 ;
        RECT 818.550 477.600 819.750 486.150 ;
        RECT 820.950 482.250 823.050 483.150 ;
        RECT 820.950 478.950 823.050 481.050 ;
        RECT 802.950 475.500 805.050 477.600 ;
        RECT 805.950 475.500 808.050 477.600 ;
        RECT 808.950 475.500 811.050 477.600 ;
        RECT 813.750 475.500 815.850 477.600 ;
        RECT 817.950 475.500 820.050 477.600 ;
        RECT 821.400 469.050 822.450 478.950 ;
        RECT 820.950 466.950 823.050 469.050 ;
        RECT 824.400 465.450 825.450 499.950 ;
        RECT 826.950 496.950 829.050 499.050 ;
        RECT 829.950 496.950 832.050 499.050 ;
        RECT 832.950 496.950 835.050 499.050 ;
        RECT 827.250 478.050 828.450 496.950 ;
        RECT 830.250 492.750 831.450 496.950 ;
        RECT 829.950 490.650 832.050 492.750 ;
        RECT 830.250 478.050 831.450 490.650 ;
        RECT 833.250 478.050 834.450 496.950 ;
        RECT 842.400 493.050 843.450 508.950 ;
        RECT 845.400 507.450 846.450 590.400 ;
        RECT 847.950 577.950 850.050 580.050 ;
        RECT 848.400 532.050 849.450 577.950 ;
        RECT 847.950 529.950 850.050 532.050 ;
        RECT 847.950 521.850 850.050 522.750 ;
        RECT 847.950 517.950 850.050 520.050 ;
        RECT 848.400 511.050 849.450 517.950 ;
        RECT 847.950 508.950 850.050 511.050 ;
        RECT 845.400 506.400 849.450 507.450 ;
        RECT 844.950 493.950 847.050 496.050 ;
        RECT 841.950 490.950 844.050 493.050 ;
        RECT 845.400 490.050 846.450 493.950 ;
        RECT 844.950 489.450 847.050 490.050 ;
        RECT 838.950 488.250 841.050 489.150 ;
        RECT 842.400 488.400 847.050 489.450 ;
        RECT 826.950 475.950 829.050 478.050 ;
        RECT 829.950 475.950 832.050 478.050 ;
        RECT 832.950 475.950 835.050 478.050 ;
        RECT 821.400 464.400 825.450 465.450 ;
        RECT 799.950 461.400 802.050 463.500 ;
        RECT 802.950 461.400 805.050 463.500 ;
        RECT 805.950 461.400 808.050 463.500 ;
        RECT 810.750 461.400 812.850 463.500 ;
        RECT 814.950 461.400 817.050 463.500 ;
        RECT 790.950 452.400 795.450 453.450 ;
        RECT 790.950 451.950 793.050 452.400 ;
        RECT 790.950 449.850 793.050 450.750 ;
        RECT 794.400 420.450 795.450 452.400 ;
        RECT 800.550 447.750 801.750 461.400 ;
        RECT 799.950 445.650 802.050 447.750 ;
        RECT 800.550 441.900 801.750 445.650 ;
        RECT 803.250 444.150 804.450 461.400 ;
        RECT 806.400 447.750 807.600 461.400 ;
        RECT 811.350 455.550 812.550 461.400 ;
        RECT 810.750 453.450 812.850 455.550 ;
        RECT 805.950 445.650 808.050 447.750 ;
        RECT 811.350 444.600 812.550 453.450 ;
        RECT 815.550 452.850 816.750 461.400 ;
        RECT 817.950 457.950 820.050 460.050 ;
        RECT 817.950 455.850 820.050 456.750 ;
        RECT 814.950 450.750 817.050 452.850 ;
        RECT 815.550 444.600 816.750 450.750 ;
        RECT 802.950 442.050 805.050 444.150 ;
        RECT 810.900 442.500 813.000 444.600 ;
        RECT 814.950 442.500 817.050 444.600 ;
        RECT 799.800 439.800 801.900 441.900 ;
        RECT 802.800 425.100 804.900 427.200 ;
        RECT 803.550 421.350 804.750 425.100 ;
        RECT 805.950 422.850 808.050 424.950 ;
        RECT 791.400 419.400 795.450 420.450 ;
        RECT 791.400 414.450 792.450 419.400 ;
        RECT 802.950 419.250 805.050 421.350 ;
        RECT 793.950 416.250 796.050 417.150 ;
        RECT 793.950 414.450 796.050 415.050 ;
        RECT 791.400 413.400 796.050 414.450 ;
        RECT 781.950 410.850 784.050 411.750 ;
        RECT 784.950 409.950 787.050 412.050 ;
        RECT 787.950 409.950 790.050 412.050 ;
        RECT 775.950 407.400 780.450 408.450 ;
        RECT 775.950 406.950 778.050 407.400 ;
        RECT 791.400 388.050 792.450 413.400 ;
        RECT 793.950 412.950 796.050 413.400 ;
        RECT 793.950 409.950 796.050 412.050 ;
        RECT 790.950 385.950 793.050 388.050 ;
        RECT 781.950 384.450 784.050 385.050 ;
        RECT 769.950 383.250 772.050 384.150 ;
        RECT 779.400 383.400 784.050 384.450 ;
        RECT 769.950 379.950 772.050 382.050 ;
        RECT 770.400 379.050 771.450 379.950 ;
        RECT 769.950 376.950 772.050 379.050 ;
        RECT 779.400 373.050 780.450 383.400 ;
        RECT 781.950 382.950 784.050 383.400 ;
        RECT 785.250 383.250 786.750 384.150 ;
        RECT 787.950 382.950 790.050 385.050 ;
        RECT 790.950 382.950 793.050 385.050 ;
        RECT 791.400 382.050 792.450 382.950 ;
        RECT 781.950 380.850 783.750 381.750 ;
        RECT 784.950 379.950 787.050 382.050 ;
        RECT 788.250 380.850 789.750 381.750 ;
        RECT 790.950 379.950 793.050 382.050 ;
        RECT 794.400 379.050 795.450 409.950 ;
        RECT 803.550 405.600 804.750 419.250 ;
        RECT 806.250 405.600 807.450 422.850 ;
        RECT 813.900 422.400 816.000 424.500 ;
        RECT 817.950 422.400 820.050 424.500 ;
        RECT 808.950 419.250 811.050 421.350 ;
        RECT 809.400 405.600 810.600 419.250 ;
        RECT 814.350 413.550 815.550 422.400 ;
        RECT 818.550 416.250 819.750 422.400 ;
        RECT 817.950 414.150 820.050 416.250 ;
        RECT 821.400 414.450 822.450 464.400 ;
        RECT 823.950 460.950 826.050 463.050 ;
        RECT 826.950 460.950 829.050 463.050 ;
        RECT 829.950 460.950 832.050 463.050 ;
        RECT 824.250 442.050 825.450 460.950 ;
        RECT 827.250 448.350 828.450 460.950 ;
        RECT 826.950 446.250 829.050 448.350 ;
        RECT 827.250 442.050 828.450 446.250 ;
        RECT 830.250 442.050 831.450 460.950 ;
        RECT 842.400 456.450 843.450 488.400 ;
        RECT 844.950 487.950 847.050 488.400 ;
        RECT 844.950 485.850 847.050 486.750 ;
        RECT 842.400 455.400 846.450 456.450 ;
        RECT 841.950 452.250 844.050 453.150 ;
        RECT 835.950 449.850 838.050 450.750 ;
        RECT 841.950 450.450 844.050 451.050 ;
        RECT 845.400 450.450 846.450 455.400 ;
        RECT 841.950 449.400 846.450 450.450 ;
        RECT 841.950 448.950 844.050 449.400 ;
        RECT 835.950 445.950 838.050 448.050 ;
        RECT 823.950 439.950 826.050 442.050 ;
        RECT 826.950 439.950 829.050 442.050 ;
        RECT 829.950 439.950 832.050 442.050 ;
        RECT 826.950 424.950 829.050 427.050 ;
        RECT 829.950 424.950 832.050 427.050 ;
        RECT 832.950 424.950 835.050 427.050 ;
        RECT 813.750 411.450 815.850 413.550 ;
        RECT 814.350 405.600 815.550 411.450 ;
        RECT 818.550 405.600 819.750 414.150 ;
        RECT 821.400 413.400 825.450 414.450 ;
        RECT 820.950 410.250 823.050 411.150 ;
        RECT 820.950 406.950 823.050 409.050 ;
        RECT 821.400 406.050 822.450 406.950 ;
        RECT 802.950 403.500 805.050 405.600 ;
        RECT 805.950 403.500 808.050 405.600 ;
        RECT 808.950 403.500 811.050 405.600 ;
        RECT 813.750 403.500 815.850 405.600 ;
        RECT 817.950 403.500 820.050 405.600 ;
        RECT 820.950 403.950 823.050 406.050 ;
        RECT 808.950 391.950 811.050 394.050 ;
        RECT 796.950 382.950 799.050 385.050 ;
        RECT 802.950 382.950 805.050 385.050 ;
        RECT 787.950 376.950 790.050 379.050 ;
        RECT 790.950 377.850 793.050 378.750 ;
        RECT 793.950 376.950 796.050 379.050 ;
        RECT 797.400 378.450 798.450 382.950 ;
        RECT 803.400 382.050 804.450 382.950 ;
        RECT 809.400 382.050 810.450 391.950 ;
        RECT 820.950 388.950 823.050 391.050 ;
        RECT 814.950 385.950 817.050 388.050 ;
        RECT 814.950 383.850 817.050 384.750 ;
        RECT 817.950 383.250 820.050 384.150 ;
        RECT 799.950 380.250 801.750 381.150 ;
        RECT 802.950 379.950 805.050 382.050 ;
        RECT 808.950 379.950 811.050 382.050 ;
        RECT 817.950 379.950 820.050 382.050 ;
        RECT 799.950 378.450 802.050 379.050 ;
        RECT 797.400 377.400 802.050 378.450 ;
        RECT 803.250 377.850 804.750 378.750 ;
        RECT 799.950 376.950 802.050 377.400 ;
        RECT 805.950 376.950 808.050 379.050 ;
        RECT 809.250 377.850 811.050 378.750 ;
        RECT 811.950 376.950 814.050 379.050 ;
        RECT 769.950 370.950 772.050 373.050 ;
        RECT 778.950 370.950 781.050 373.050 ;
        RECT 770.400 358.050 771.450 370.950 ;
        RECT 769.950 355.950 772.050 358.050 ;
        RECT 757.950 341.250 760.050 342.150 ;
        RECT 760.950 340.950 763.050 343.050 ;
        RECT 763.950 341.250 766.050 342.150 ;
        RECT 766.950 340.950 769.050 343.050 ;
        RECT 757.950 337.950 760.050 340.050 ;
        RECT 761.250 338.250 762.750 339.150 ;
        RECT 763.950 337.950 766.050 340.050 ;
        RECT 754.950 319.950 757.050 322.050 ;
        RECT 758.400 319.050 759.450 337.950 ;
        RECT 764.400 337.050 765.450 337.950 ;
        RECT 760.950 334.950 763.050 337.050 ;
        RECT 763.950 334.950 766.050 337.050 ;
        RECT 761.400 334.050 762.450 334.950 ;
        RECT 760.950 331.950 763.050 334.050 ;
        RECT 760.950 319.950 763.050 322.050 ;
        RECT 754.950 316.950 757.050 319.050 ;
        RECT 757.950 316.950 760.050 319.050 ;
        RECT 742.950 315.450 745.050 316.050 ;
        RECT 740.400 314.400 747.450 315.450 ;
        RECT 742.950 313.950 745.050 314.400 ;
        RECT 739.950 311.250 742.050 312.150 ;
        RECT 742.950 311.850 745.050 312.750 ;
        RECT 739.950 307.950 742.050 310.050 ;
        RECT 740.400 301.050 741.450 307.950 ;
        RECT 739.950 298.950 742.050 301.050 ;
        RECT 739.950 280.950 742.050 283.050 ;
        RECT 742.950 280.950 745.050 283.050 ;
        RECT 740.400 277.050 741.450 280.950 ;
        RECT 736.950 274.950 739.050 277.050 ;
        RECT 739.950 274.950 742.050 277.050 ;
        RECT 743.400 274.050 744.450 280.950 ;
        RECT 746.400 277.050 747.450 314.400 ;
        RECT 748.950 310.950 751.050 313.050 ;
        RECT 745.950 274.950 748.050 277.050 ;
        RECT 749.400 274.050 750.450 310.950 ;
        RECT 755.400 310.050 756.450 316.950 ;
        RECT 761.400 310.050 762.450 319.950 ;
        RECT 751.950 308.250 753.750 309.150 ;
        RECT 754.950 307.950 757.050 310.050 ;
        RECT 760.950 307.950 763.050 310.050 ;
        RECT 751.950 304.950 754.050 307.050 ;
        RECT 755.250 305.850 756.750 306.750 ;
        RECT 757.950 304.950 760.050 307.050 ;
        RECT 761.250 305.850 763.050 306.750 ;
        RECT 757.950 302.850 760.050 303.750 ;
        RECT 764.400 295.050 765.450 334.950 ;
        RECT 767.400 325.050 768.450 340.950 ;
        RECT 770.400 331.050 771.450 355.950 ;
        RECT 784.950 352.950 787.050 355.050 ;
        RECT 781.950 343.950 784.050 346.050 ;
        RECT 772.950 341.250 775.050 342.150 ;
        RECT 778.950 341.250 781.050 342.150 ;
        RECT 772.950 337.950 775.050 340.050 ;
        RECT 776.250 338.250 777.750 339.150 ;
        RECT 778.950 337.950 781.050 340.050 ;
        RECT 773.400 334.050 774.450 337.950 ;
        RECT 775.950 334.950 778.050 337.050 ;
        RECT 772.950 331.950 775.050 334.050 ;
        RECT 769.950 328.950 772.050 331.050 ;
        RECT 779.400 328.050 780.450 337.950 ;
        RECT 782.400 337.050 783.450 343.950 ;
        RECT 785.400 340.050 786.450 352.950 ;
        RECT 784.950 337.950 787.050 340.050 ;
        RECT 781.950 334.950 784.050 337.050 ;
        RECT 769.950 325.950 772.050 328.050 ;
        RECT 778.950 325.950 781.050 328.050 ;
        RECT 766.950 322.950 769.050 325.050 ;
        RECT 767.400 316.050 768.450 322.950 ;
        RECT 770.400 316.050 771.450 325.950 ;
        RECT 775.950 316.950 778.050 319.050 ;
        RECT 766.950 313.950 769.050 316.050 ;
        RECT 769.950 313.950 772.050 316.050 ;
        RECT 767.400 313.050 768.450 313.950 ;
        RECT 766.950 310.950 769.050 313.050 ;
        RECT 770.250 311.850 771.750 312.750 ;
        RECT 772.950 310.950 775.050 313.050 ;
        RECT 766.950 308.850 769.050 309.750 ;
        RECT 772.950 308.850 775.050 309.750 ;
        RECT 766.950 304.950 769.050 307.050 ;
        RECT 763.950 292.950 766.050 295.050 ;
        RECT 760.950 283.950 763.050 286.050 ;
        RECT 757.950 277.950 760.050 280.050 ;
        RECT 754.950 274.950 757.050 277.050 ;
        RECT 736.950 271.950 739.050 274.050 ;
        RECT 742.950 273.450 745.050 274.050 ;
        RECT 740.250 272.250 741.750 273.150 ;
        RECT 742.950 272.400 747.450 273.450 ;
        RECT 742.950 271.950 745.050 272.400 ;
        RECT 736.950 269.850 738.750 270.750 ;
        RECT 739.950 268.950 742.050 271.050 ;
        RECT 743.250 269.850 745.050 270.750 ;
        RECT 736.950 259.950 739.050 262.050 ;
        RECT 733.950 253.950 736.050 256.050 ;
        RECT 733.950 250.950 736.050 253.050 ;
        RECT 730.950 244.950 733.050 247.050 ;
        RECT 724.950 241.950 727.050 244.050 ;
        RECT 721.950 238.950 724.050 241.050 ;
        RECT 725.250 239.850 726.750 240.750 ;
        RECT 727.950 238.950 730.050 241.050 ;
        RECT 721.950 236.850 724.050 237.750 ;
        RECT 724.950 235.950 727.050 238.050 ;
        RECT 727.950 236.850 730.050 237.750 ;
        RECT 725.400 223.050 726.450 235.950 ;
        RECT 724.950 220.950 727.050 223.050 ;
        RECT 724.950 200.250 727.050 201.150 ;
        RECT 715.950 197.250 717.750 198.150 ;
        RECT 718.950 196.950 721.050 199.050 ;
        RECT 722.250 197.250 723.750 198.150 ;
        RECT 724.950 196.950 727.050 199.050 ;
        RECT 727.950 196.950 730.050 199.050 ;
        RECT 715.950 193.950 718.050 196.050 ;
        RECT 719.250 194.850 720.750 195.750 ;
        RECT 721.950 193.950 724.050 196.050 ;
        RECT 703.950 190.950 706.050 193.050 ;
        RECT 712.950 190.950 715.050 193.050 ;
        RECT 703.950 181.950 706.050 184.050 ;
        RECT 700.950 175.950 703.050 178.050 ;
        RECT 679.950 169.950 682.050 172.050 ;
        RECT 685.950 169.950 688.050 172.050 ;
        RECT 697.950 169.950 700.050 172.050 ;
        RECT 680.400 166.050 681.450 169.950 ;
        RECT 679.950 163.950 682.050 166.050 ;
        RECT 683.250 164.250 685.050 165.150 ;
        RECT 673.950 161.850 675.750 162.750 ;
        RECT 676.950 160.950 679.050 163.050 ;
        RECT 680.250 161.850 681.750 162.750 ;
        RECT 682.950 160.950 685.050 163.050 ;
        RECT 683.400 160.050 684.450 160.950 ;
        RECT 673.950 157.950 676.050 160.050 ;
        RECT 676.950 158.850 679.050 159.750 ;
        RECT 682.950 157.950 685.050 160.050 ;
        RECT 674.400 157.050 675.450 157.950 ;
        RECT 673.950 154.950 676.050 157.050 ;
        RECT 673.950 145.950 676.050 148.050 ;
        RECT 661.950 124.950 664.050 127.050 ;
        RECT 665.250 125.850 667.050 126.750 ;
        RECT 670.950 124.950 673.050 127.050 ;
        RECT 658.950 121.950 661.050 124.050 ;
        RECT 658.950 120.450 661.050 121.050 ;
        RECT 662.400 120.450 663.450 124.950 ;
        RECT 674.400 121.050 675.450 145.950 ;
        RECT 686.400 144.450 687.450 169.950 ;
        RECT 698.400 166.050 699.450 169.950 ;
        RECT 691.950 163.950 694.050 166.050 ;
        RECT 697.950 163.950 700.050 166.050 ;
        RECT 701.250 164.250 703.050 165.150 ;
        RECT 688.950 160.950 691.050 163.050 ;
        RECT 691.950 161.850 693.750 162.750 ;
        RECT 694.950 160.950 697.050 163.050 ;
        RECT 698.250 161.850 699.750 162.750 ;
        RECT 700.950 160.950 703.050 163.050 ;
        RECT 689.400 148.050 690.450 160.950 ;
        RECT 694.950 158.850 697.050 159.750 ;
        RECT 700.950 157.950 703.050 160.050 ;
        RECT 688.950 145.950 691.050 148.050 ;
        RECT 686.400 143.400 690.450 144.450 ;
        RECT 679.950 127.950 682.050 130.050 ;
        RECT 680.400 127.050 681.450 127.950 ;
        RECT 676.950 125.250 678.750 126.150 ;
        RECT 679.950 124.950 682.050 127.050 ;
        RECT 685.950 124.950 688.050 127.050 ;
        RECT 689.400 124.050 690.450 143.400 ;
        RECT 697.950 139.950 700.050 142.050 ;
        RECT 698.400 130.050 699.450 139.950 ;
        RECT 701.400 130.050 702.450 157.950 ;
        RECT 691.950 127.950 694.050 130.050 ;
        RECT 695.250 128.250 696.750 129.150 ;
        RECT 697.950 127.950 700.050 130.050 ;
        RECT 700.950 127.950 703.050 130.050 ;
        RECT 691.950 125.850 693.750 126.750 ;
        RECT 694.950 124.950 697.050 127.050 ;
        RECT 698.250 125.850 700.050 126.750 ;
        RECT 676.950 121.950 679.050 124.050 ;
        RECT 680.250 122.850 682.050 123.750 ;
        RECT 682.950 122.250 685.050 123.150 ;
        RECT 685.950 122.850 688.050 123.750 ;
        RECT 688.950 121.950 691.050 124.050 ;
        RECT 694.950 121.950 697.050 124.050 ;
        RECT 658.950 119.400 663.450 120.450 ;
        RECT 658.950 118.950 661.050 119.400 ;
        RECT 673.950 118.950 676.050 121.050 ;
        RECT 682.950 118.950 685.050 121.050 ;
        RECT 655.950 112.950 658.050 115.050 ;
        RECT 652.950 88.950 655.050 91.050 ;
        RECT 646.950 73.950 649.050 76.050 ;
        RECT 604.950 64.950 607.050 67.050 ;
        RECT 619.950 64.950 622.050 67.050 ;
        RECT 640.800 65.100 642.900 67.200 ;
        RECT 659.400 67.050 660.450 118.950 ;
        RECT 685.950 112.950 688.050 115.050 ;
        RECT 673.950 100.950 676.050 103.050 ;
        RECT 670.950 97.950 673.050 100.050 ;
        RECT 671.400 97.050 672.450 97.950 ;
        RECT 661.950 94.950 664.050 97.050 ;
        RECT 664.950 94.950 667.050 97.050 ;
        RECT 668.250 95.250 669.750 96.150 ;
        RECT 670.950 94.950 673.050 97.050 ;
        RECT 662.400 94.050 663.450 94.950 ;
        RECT 661.950 91.950 664.050 94.050 ;
        RECT 665.250 92.850 666.750 93.750 ;
        RECT 667.950 91.950 670.050 94.050 ;
        RECT 671.250 92.850 673.050 93.750 ;
        RECT 668.400 91.050 669.450 91.950 ;
        RECT 661.950 89.850 664.050 90.750 ;
        RECT 667.950 88.950 670.050 91.050 ;
        RECT 674.400 88.050 675.450 100.950 ;
        RECT 679.950 97.950 682.050 100.050 ;
        RECT 676.950 94.950 679.050 97.050 ;
        RECT 676.950 92.850 679.050 93.750 ;
        RECT 673.950 85.950 676.050 88.050 ;
        RECT 680.400 82.050 681.450 97.950 ;
        RECT 686.400 97.050 687.450 112.950 ;
        RECT 691.950 103.950 694.050 106.050 ;
        RECT 692.400 97.050 693.450 103.950 ;
        RECT 695.400 100.050 696.450 121.950 ;
        RECT 701.400 115.050 702.450 127.950 ;
        RECT 700.950 112.950 703.050 115.050 ;
        RECT 694.950 97.950 697.050 100.050 ;
        RECT 685.950 94.950 688.050 97.050 ;
        RECT 688.950 94.950 691.050 97.050 ;
        RECT 691.950 94.950 694.050 97.050 ;
        RECT 695.250 95.850 696.750 96.750 ;
        RECT 697.950 96.450 700.050 97.050 ;
        RECT 697.950 95.400 702.450 96.450 ;
        RECT 697.950 94.950 700.050 95.400 ;
        RECT 682.950 92.250 685.050 93.150 ;
        RECT 685.950 92.850 688.050 93.750 ;
        RECT 682.950 88.950 685.050 91.050 ;
        RECT 683.400 88.050 684.450 88.950 ;
        RECT 689.400 88.050 690.450 94.950 ;
        RECT 691.950 92.850 694.050 93.750 ;
        RECT 697.950 92.850 700.050 93.750 ;
        RECT 682.950 85.950 685.050 88.050 ;
        RECT 688.950 85.950 691.050 88.050 ;
        RECT 697.950 85.950 700.050 88.050 ;
        RECT 679.950 79.950 682.050 82.050 ;
        RECT 694.950 73.950 697.050 76.050 ;
        RECT 601.950 58.950 604.050 61.050 ;
        RECT 610.950 58.950 613.050 61.050 ;
        RECT 611.400 58.050 612.450 58.950 ;
        RECT 604.950 56.250 607.050 57.150 ;
        RECT 610.950 55.950 613.050 58.050 ;
        RECT 620.400 55.050 621.450 64.950 ;
        RECT 641.550 61.350 642.750 65.100 ;
        RECT 658.950 64.950 661.050 67.050 ;
        RECT 664.950 64.950 667.050 67.050 ;
        RECT 667.950 64.950 670.050 67.050 ;
        RECT 670.950 64.950 673.050 67.050 ;
        RECT 643.950 62.850 646.050 64.950 ;
        RECT 640.950 59.250 643.050 61.350 ;
        RECT 631.950 56.250 634.050 57.150 ;
        RECT 601.950 52.950 604.050 55.050 ;
        RECT 610.950 53.850 613.050 54.750 ;
        RECT 619.950 52.950 622.050 55.050 ;
        RECT 631.950 52.950 634.050 55.050 ;
        RECT 568.950 43.500 571.050 45.600 ;
        RECT 571.950 43.500 574.050 45.600 ;
        RECT 574.950 43.500 577.050 45.600 ;
        RECT 579.750 43.500 581.850 45.600 ;
        RECT 583.950 43.500 586.050 45.600 ;
        RECT 592.950 43.950 595.050 46.050 ;
        RECT 595.950 43.950 598.050 46.050 ;
        RECT 598.950 43.950 601.050 46.050 ;
        RECT 559.950 25.950 562.050 28.050 ;
        RECT 577.950 25.950 580.050 28.050 ;
        RECT 529.950 18.450 532.050 19.050 ;
        RECT 527.400 17.400 532.050 18.450 ;
        RECT 533.250 17.850 534.750 18.750 ;
        RECT 529.950 16.950 532.050 17.400 ;
        RECT 535.950 16.950 538.050 19.050 ;
        RECT 541.950 17.850 543.750 18.750 ;
        RECT 544.950 16.950 547.050 19.050 ;
        RECT 548.250 17.850 549.750 18.750 ;
        RECT 550.950 16.950 553.050 19.050 ;
        RECT 553.950 16.950 556.050 19.050 ;
        RECT 560.400 18.450 561.450 25.950 ;
        RECT 565.950 22.950 568.050 25.050 ;
        RECT 566.400 22.050 567.450 22.950 ;
        RECT 578.400 22.050 579.450 25.950 ;
        RECT 583.950 22.950 586.050 25.050 ;
        RECT 589.950 23.250 592.050 24.150 ;
        RECT 562.950 20.250 564.750 21.150 ;
        RECT 565.950 19.950 568.050 22.050 ;
        RECT 569.250 20.250 571.050 21.150 ;
        RECT 574.950 20.250 576.750 21.150 ;
        RECT 577.950 19.950 580.050 22.050 ;
        RECT 581.250 20.250 583.050 21.150 ;
        RECT 562.950 18.450 565.050 19.050 ;
        RECT 560.400 17.400 565.050 18.450 ;
        RECT 566.250 17.850 567.750 18.750 ;
        RECT 562.950 16.950 565.050 17.400 ;
        RECT 568.950 16.950 571.050 19.050 ;
        RECT 574.950 16.950 577.050 19.050 ;
        RECT 578.250 17.850 579.750 18.750 ;
        RECT 580.950 18.450 583.050 19.050 ;
        RECT 584.400 18.450 585.450 22.950 ;
        RECT 602.400 22.050 603.450 52.950 ;
        RECT 619.950 50.850 622.050 51.750 ;
        RECT 632.400 49.050 633.450 52.950 ;
        RECT 631.950 46.950 634.050 49.050 ;
        RECT 641.550 45.600 642.750 59.250 ;
        RECT 644.250 45.600 645.450 62.850 ;
        RECT 651.900 62.400 654.000 64.500 ;
        RECT 655.950 62.400 658.050 64.500 ;
        RECT 646.950 59.250 649.050 61.350 ;
        RECT 647.400 45.600 648.600 59.250 ;
        RECT 652.350 53.550 653.550 62.400 ;
        RECT 656.550 56.250 657.750 62.400 ;
        RECT 661.950 58.950 664.050 61.050 ;
        RECT 655.950 54.150 658.050 56.250 ;
        RECT 651.750 51.450 653.850 53.550 ;
        RECT 652.350 45.600 653.550 51.450 ;
        RECT 656.550 45.600 657.750 54.150 ;
        RECT 658.950 50.250 661.050 51.150 ;
        RECT 658.950 46.950 661.050 49.050 ;
        RECT 640.950 43.500 643.050 45.600 ;
        RECT 643.950 43.500 646.050 45.600 ;
        RECT 646.950 43.500 649.050 45.600 ;
        RECT 651.750 43.500 653.850 45.600 ;
        RECT 655.950 43.500 658.050 45.600 ;
        RECT 659.400 37.050 660.450 46.950 ;
        RECT 658.950 34.950 661.050 37.050 ;
        RECT 610.950 29.400 613.050 31.500 ;
        RECT 613.950 29.400 616.050 31.500 ;
        RECT 616.950 29.400 619.050 31.500 ;
        RECT 621.750 29.400 623.850 31.500 ;
        RECT 625.950 29.400 628.050 31.500 ;
        RECT 589.950 19.950 592.050 22.050 ;
        RECT 601.950 19.950 604.050 22.050 ;
        RECT 590.400 19.050 591.450 19.950 ;
        RECT 580.950 17.400 585.450 18.450 ;
        RECT 580.950 16.950 583.050 17.400 ;
        RECT 589.950 16.950 592.050 19.050 ;
        RECT 601.950 17.850 604.050 18.750 ;
        RECT 536.400 16.050 537.450 16.950 ;
        RECT 551.400 16.050 552.450 16.950 ;
        RECT 575.400 16.050 576.450 16.950 ;
        RECT 535.950 13.950 538.050 16.050 ;
        RECT 544.950 14.850 547.050 15.750 ;
        RECT 550.950 13.950 553.050 16.050 ;
        RECT 574.950 13.950 577.050 16.050 ;
        RECT 611.550 15.750 612.750 29.400 ;
        RECT 610.950 13.650 613.050 15.750 ;
        RECT 611.550 9.900 612.750 13.650 ;
        RECT 614.250 12.150 615.450 29.400 ;
        RECT 617.400 15.750 618.600 29.400 ;
        RECT 622.350 23.550 623.550 29.400 ;
        RECT 621.750 21.450 623.850 23.550 ;
        RECT 616.950 13.650 619.050 15.750 ;
        RECT 622.350 12.600 623.550 21.450 ;
        RECT 626.550 20.850 627.750 29.400 ;
        RECT 634.950 28.950 637.050 31.050 ;
        RECT 637.950 28.950 640.050 31.050 ;
        RECT 640.950 28.950 643.050 31.050 ;
        RECT 628.950 25.950 631.050 28.050 ;
        RECT 628.950 23.850 631.050 24.750 ;
        RECT 625.950 18.750 628.050 20.850 ;
        RECT 626.550 12.600 627.750 18.750 ;
        RECT 613.950 10.050 616.050 12.150 ;
        RECT 621.900 10.500 624.000 12.600 ;
        RECT 625.950 10.500 628.050 12.600 ;
        RECT 635.250 10.050 636.450 28.950 ;
        RECT 638.250 16.350 639.450 28.950 ;
        RECT 637.950 14.250 640.050 16.350 ;
        RECT 638.250 10.050 639.450 14.250 ;
        RECT 641.250 10.050 642.450 28.950 ;
        RECT 662.400 28.050 663.450 58.950 ;
        RECT 665.250 46.050 666.450 64.950 ;
        RECT 668.250 60.750 669.450 64.950 ;
        RECT 667.950 58.650 670.050 60.750 ;
        RECT 668.250 46.050 669.450 58.650 ;
        RECT 671.250 46.050 672.450 64.950 ;
        RECT 682.950 58.950 685.050 61.050 ;
        RECT 683.400 58.050 684.450 58.950 ;
        RECT 676.950 56.250 679.050 57.150 ;
        RECT 682.950 55.950 685.050 58.050 ;
        RECT 673.950 52.950 676.050 55.050 ;
        RECT 682.950 53.850 685.050 54.750 ;
        RECT 664.950 43.950 667.050 46.050 ;
        RECT 667.950 43.950 670.050 46.050 ;
        RECT 670.950 43.950 673.050 46.050 ;
        RECT 664.950 31.950 667.050 34.050 ;
        RECT 665.400 28.050 666.450 31.950 ;
        RECT 655.950 25.950 658.050 28.050 ;
        RECT 661.950 25.950 664.050 28.050 ;
        RECT 664.950 25.950 667.050 28.050 ;
        RECT 670.950 25.950 673.050 28.050 ;
        RECT 652.950 20.250 655.050 21.150 ;
        RECT 646.950 17.850 649.050 18.750 ;
        RECT 652.950 18.450 655.050 19.050 ;
        RECT 656.400 18.450 657.450 25.950 ;
        RECT 671.400 25.050 672.450 25.950 ;
        RECT 661.950 23.250 664.050 24.150 ;
        RECT 664.950 23.850 667.050 24.750 ;
        RECT 667.950 23.250 669.750 24.150 ;
        RECT 670.950 22.950 673.050 25.050 ;
        RECT 674.400 22.050 675.450 52.950 ;
        RECT 682.950 34.950 685.050 37.050 ;
        RECT 683.400 28.050 684.450 34.950 ;
        RECT 679.950 25.950 682.050 28.050 ;
        RECT 682.950 25.950 685.050 28.050 ;
        RECT 685.950 25.950 688.050 28.050 ;
        RECT 680.400 25.050 681.450 25.950 ;
        RECT 686.400 25.050 687.450 25.950 ;
        RECT 695.400 25.050 696.450 73.950 ;
        RECT 698.400 58.050 699.450 85.950 ;
        RECT 701.400 70.050 702.450 95.400 ;
        RECT 700.950 67.950 703.050 70.050 ;
        RECT 704.400 63.450 705.450 181.950 ;
        RECT 716.400 172.050 717.450 193.950 ;
        RECT 722.400 181.050 723.450 193.950 ;
        RECT 725.400 193.050 726.450 196.950 ;
        RECT 724.950 190.950 727.050 193.050 ;
        RECT 724.950 187.950 727.050 190.050 ;
        RECT 721.950 178.950 724.050 181.050 ;
        RECT 721.950 175.950 724.050 178.050 ;
        RECT 715.950 169.950 718.050 172.050 ;
        RECT 709.950 165.450 712.050 166.050 ;
        RECT 707.400 164.400 712.050 165.450 ;
        RECT 707.400 142.050 708.450 164.400 ;
        RECT 709.950 163.950 712.050 164.400 ;
        RECT 715.950 163.950 718.050 166.050 ;
        RECT 719.250 164.250 721.050 165.150 ;
        RECT 709.950 161.850 711.750 162.750 ;
        RECT 712.950 160.950 715.050 163.050 ;
        RECT 716.250 161.850 717.750 162.750 ;
        RECT 718.950 162.450 721.050 163.050 ;
        RECT 722.400 162.450 723.450 175.950 ;
        RECT 718.950 161.400 723.450 162.450 ;
        RECT 718.950 160.950 721.050 161.400 ;
        RECT 712.950 158.850 715.050 159.750 ;
        RECT 706.950 139.950 709.050 142.050 ;
        RECT 725.400 139.050 726.450 187.950 ;
        RECT 724.950 136.950 727.050 139.050 ;
        RECT 718.950 132.450 721.050 133.050 ;
        RECT 721.950 132.450 724.050 133.050 ;
        RECT 718.950 131.400 724.050 132.450 ;
        RECT 728.400 132.450 729.450 196.950 ;
        RECT 731.400 193.050 732.450 244.950 ;
        RECT 734.400 229.050 735.450 250.950 ;
        RECT 737.400 232.050 738.450 259.950 ;
        RECT 740.400 259.050 741.450 268.950 ;
        RECT 742.950 265.950 745.050 268.050 ;
        RECT 739.950 256.950 742.050 259.050 ;
        RECT 743.400 250.050 744.450 265.950 ;
        RECT 746.400 253.050 747.450 272.400 ;
        RECT 748.950 271.950 751.050 274.050 ;
        RECT 745.950 250.950 748.050 253.050 ;
        RECT 742.950 247.950 745.050 250.050 ;
        RECT 739.950 241.950 742.050 244.050 ;
        RECT 742.950 241.950 745.050 244.050 ;
        RECT 740.400 241.050 741.450 241.950 ;
        RECT 746.400 241.050 747.450 250.950 ;
        RECT 739.950 238.950 742.050 241.050 ;
        RECT 743.250 239.850 744.750 240.750 ;
        RECT 745.950 238.950 748.050 241.050 ;
        RECT 739.950 236.850 742.050 237.750 ;
        RECT 745.950 236.850 748.050 237.750 ;
        RECT 736.950 229.950 739.050 232.050 ;
        RECT 733.950 226.950 736.050 229.050 ;
        RECT 749.400 214.050 750.450 271.950 ;
        RECT 755.400 271.050 756.450 274.950 ;
        RECT 758.400 271.050 759.450 277.950 ;
        RECT 761.400 273.450 762.450 283.950 ;
        RECT 761.400 272.400 765.450 273.450 ;
        RECT 751.950 269.250 753.750 270.150 ;
        RECT 754.950 268.950 757.050 271.050 ;
        RECT 757.950 268.950 760.050 271.050 ;
        RECT 760.950 268.950 763.050 271.050 ;
        RECT 751.950 265.950 754.050 268.050 ;
        RECT 755.250 266.850 757.050 267.750 ;
        RECT 757.950 266.250 760.050 267.150 ;
        RECT 760.950 266.850 763.050 267.750 ;
        RECT 752.400 262.050 753.450 265.950 ;
        RECT 757.950 262.950 760.050 265.050 ;
        RECT 751.950 259.950 754.050 262.050 ;
        RECT 758.400 259.050 759.450 262.950 ;
        RECT 757.950 256.950 760.050 259.050 ;
        RECT 751.950 247.950 754.050 250.050 ;
        RECT 754.950 247.950 757.050 250.050 ;
        RECT 752.400 241.050 753.450 247.950 ;
        RECT 755.400 244.050 756.450 247.950 ;
        RECT 764.400 244.050 765.450 272.400 ;
        RECT 767.400 271.050 768.450 304.950 ;
        RECT 776.400 283.050 777.450 316.950 ;
        RECT 782.400 316.050 783.450 334.950 ;
        RECT 788.400 328.050 789.450 376.950 ;
        RECT 805.950 374.850 808.050 375.750 ;
        RECT 802.950 349.950 805.050 352.050 ;
        RECT 793.950 347.250 796.050 348.150 ;
        RECT 799.950 346.950 802.050 349.050 ;
        RECT 800.400 346.050 801.450 346.950 ;
        RECT 790.950 344.250 792.750 345.150 ;
        RECT 793.950 343.950 796.050 346.050 ;
        RECT 797.250 344.250 798.750 345.150 ;
        RECT 799.950 343.950 802.050 346.050 ;
        RECT 790.950 340.950 793.050 343.050 ;
        RECT 796.950 340.950 799.050 343.050 ;
        RECT 800.250 341.850 802.050 342.750 ;
        RECT 791.400 340.050 792.450 340.950 ;
        RECT 790.950 337.950 793.050 340.050 ;
        RECT 797.400 339.450 798.450 340.950 ;
        RECT 803.400 339.450 804.450 349.950 ;
        RECT 812.400 346.050 813.450 376.950 ;
        RECT 818.400 346.050 819.450 379.950 ;
        RECT 821.400 379.050 822.450 388.950 ;
        RECT 820.950 376.950 823.050 379.050 ;
        RECT 821.400 352.050 822.450 376.950 ;
        RECT 820.950 349.950 823.050 352.050 ;
        RECT 824.400 348.450 825.450 413.400 ;
        RECT 827.250 406.050 828.450 424.950 ;
        RECT 830.250 420.750 831.450 424.950 ;
        RECT 829.950 418.650 832.050 420.750 ;
        RECT 830.250 406.050 831.450 418.650 ;
        RECT 833.250 406.050 834.450 424.950 ;
        RECT 836.400 411.450 837.450 445.950 ;
        RECT 838.950 416.250 841.050 417.150 ;
        RECT 838.950 414.450 841.050 415.050 ;
        RECT 842.400 414.450 843.450 448.950 ;
        RECT 838.950 413.400 843.450 414.450 ;
        RECT 844.950 413.850 847.050 414.750 ;
        RECT 838.950 412.950 841.050 413.400 ;
        RECT 836.400 410.400 840.450 411.450 ;
        RECT 835.950 406.950 838.050 409.050 ;
        RECT 826.950 403.950 829.050 406.050 ;
        RECT 829.950 403.950 832.050 406.050 ;
        RECT 832.950 403.950 835.050 406.050 ;
        RECT 826.950 380.250 828.750 381.150 ;
        RECT 829.950 379.950 832.050 382.050 ;
        RECT 833.250 380.250 835.050 381.150 ;
        RECT 826.950 376.950 829.050 379.050 ;
        RECT 830.250 377.850 831.750 378.750 ;
        RECT 832.950 376.950 835.050 379.050 ;
        RECT 827.400 373.050 828.450 376.950 ;
        RECT 836.400 376.050 837.450 406.950 ;
        RECT 835.950 373.950 838.050 376.050 ;
        RECT 826.950 370.950 829.050 373.050 ;
        RECT 827.400 355.050 828.450 370.950 ;
        RECT 839.400 370.050 840.450 410.400 ;
        RECT 841.950 409.950 844.050 412.050 ;
        RECT 842.400 379.050 843.450 409.950 ;
        RECT 848.400 409.050 849.450 506.400 ;
        RECT 847.950 406.950 850.050 409.050 ;
        RECT 844.950 385.950 847.050 388.050 ;
        RECT 841.950 376.950 844.050 379.050 ;
        RECT 838.950 367.950 841.050 370.050 ;
        RECT 845.400 366.450 846.450 385.950 ;
        RECT 847.950 383.250 850.050 384.150 ;
        RECT 847.950 379.950 850.050 382.050 ;
        RECT 847.950 373.950 850.050 376.050 ;
        RECT 842.400 365.400 846.450 366.450 ;
        RECT 826.950 352.950 829.050 355.050 ;
        RECT 821.400 347.400 825.450 348.450 ;
        RECT 805.950 343.950 808.050 346.050 ;
        RECT 808.950 344.250 811.050 345.150 ;
        RECT 811.950 343.950 814.050 346.050 ;
        RECT 817.950 343.950 820.050 346.050 ;
        RECT 806.400 342.450 807.450 343.950 ;
        RECT 808.950 342.450 811.050 343.050 ;
        RECT 806.400 341.400 811.050 342.450 ;
        RECT 808.950 340.950 811.050 341.400 ;
        RECT 812.250 341.250 813.750 342.150 ;
        RECT 814.950 340.950 817.050 343.050 ;
        RECT 818.250 341.250 820.050 342.150 ;
        RECT 797.400 338.400 804.450 339.450 ;
        RECT 811.950 337.950 814.050 340.050 ;
        RECT 815.250 338.850 816.750 339.750 ;
        RECT 817.950 337.950 820.050 340.050 ;
        RECT 793.950 334.950 796.050 337.050 ;
        RECT 787.950 325.950 790.050 328.050 ;
        RECT 781.950 313.950 784.050 316.050 ;
        RECT 778.950 312.450 781.050 313.050 ;
        RECT 781.950 312.450 784.050 313.050 ;
        RECT 778.950 311.400 784.050 312.450 ;
        RECT 778.950 310.950 781.050 311.400 ;
        RECT 781.950 310.950 784.050 311.400 ;
        RECT 785.250 311.250 786.750 312.150 ;
        RECT 787.950 310.950 790.050 313.050 ;
        RECT 779.400 304.050 780.450 310.950 ;
        RECT 781.950 308.850 783.750 309.750 ;
        RECT 784.950 307.950 787.050 310.050 ;
        RECT 788.250 308.850 789.750 309.750 ;
        RECT 790.950 307.950 793.050 310.050 ;
        RECT 790.950 305.850 793.050 306.750 ;
        RECT 778.950 301.950 781.050 304.050 ;
        RECT 787.950 295.950 790.050 298.050 ;
        RECT 781.950 286.950 784.050 289.050 ;
        RECT 775.950 280.950 778.050 283.050 ;
        RECT 775.950 277.950 778.050 280.050 ;
        RECT 769.950 272.250 772.050 273.150 ;
        RECT 776.400 271.050 777.450 277.950 ;
        RECT 766.950 268.950 769.050 271.050 ;
        RECT 769.950 268.950 772.050 271.050 ;
        RECT 773.250 269.250 774.750 270.150 ;
        RECT 775.950 268.950 778.050 271.050 ;
        RECT 779.250 269.250 781.050 270.150 ;
        RECT 766.950 265.950 769.050 268.050 ;
        RECT 767.400 256.050 768.450 265.950 ;
        RECT 770.400 262.050 771.450 268.950 ;
        RECT 772.950 265.950 775.050 268.050 ;
        RECT 776.250 266.850 777.750 267.750 ;
        RECT 778.950 265.950 781.050 268.050 ;
        RECT 773.400 265.050 774.450 265.950 ;
        RECT 772.950 262.950 775.050 265.050 ;
        RECT 769.950 259.950 772.050 262.050 ;
        RECT 766.950 253.950 769.050 256.050 ;
        RECT 779.400 244.050 780.450 265.950 ;
        RECT 754.950 241.950 757.050 244.050 ;
        RECT 757.950 241.950 760.050 244.050 ;
        RECT 763.950 241.950 766.050 244.050 ;
        RECT 778.950 241.950 781.050 244.050 ;
        RECT 758.400 241.050 759.450 241.950 ;
        RECT 751.950 238.950 754.050 241.050 ;
        RECT 755.250 239.850 756.750 240.750 ;
        RECT 757.950 238.950 760.050 241.050 ;
        RECT 760.950 238.950 763.050 241.050 ;
        RECT 751.950 236.850 754.050 237.750 ;
        RECT 757.950 236.850 760.050 237.750 ;
        RECT 761.400 232.050 762.450 238.950 ;
        RECT 764.400 238.050 765.450 241.950 ;
        RECT 779.400 241.050 780.450 241.950 ;
        RECT 766.950 238.950 769.050 241.050 ;
        RECT 772.950 240.450 775.050 241.050 ;
        RECT 775.950 240.450 778.050 241.050 ;
        RECT 770.250 239.250 771.750 240.150 ;
        RECT 772.950 239.400 778.050 240.450 ;
        RECT 772.950 238.950 775.050 239.400 ;
        RECT 775.950 238.950 778.050 239.400 ;
        RECT 778.950 238.950 781.050 241.050 ;
        RECT 763.950 235.950 766.050 238.050 ;
        RECT 766.950 236.850 768.750 237.750 ;
        RECT 769.950 235.950 772.050 238.050 ;
        RECT 773.250 236.850 774.750 237.750 ;
        RECT 775.950 235.950 778.050 238.050 ;
        RECT 760.950 229.950 763.050 232.050 ;
        RECT 748.950 211.950 751.050 214.050 ;
        RECT 748.950 208.950 751.050 211.050 ;
        RECT 733.950 202.950 736.050 205.050 ;
        RECT 742.950 203.250 745.050 204.150 ;
        RECT 734.400 196.050 735.450 202.950 ;
        RECT 736.950 199.950 739.050 202.050 ;
        RECT 740.250 200.250 741.750 201.150 ;
        RECT 742.950 199.950 745.050 202.050 ;
        RECT 746.250 200.250 748.050 201.150 ;
        RECT 736.950 197.850 738.750 198.750 ;
        RECT 739.950 196.950 742.050 199.050 ;
        RECT 740.400 196.050 741.450 196.950 ;
        RECT 743.400 196.050 744.450 199.950 ;
        RECT 745.950 196.950 748.050 199.050 ;
        RECT 733.950 193.950 736.050 196.050 ;
        RECT 739.950 193.950 742.050 196.050 ;
        RECT 742.950 193.950 745.050 196.050 ;
        RECT 730.950 190.950 733.050 193.050 ;
        RECT 745.950 190.950 748.050 193.050 ;
        RECT 730.950 172.950 733.050 175.050 ;
        RECT 731.400 172.050 732.450 172.950 ;
        RECT 730.950 169.950 733.050 172.050 ;
        RECT 736.950 169.950 739.050 172.050 ;
        RECT 742.950 169.950 745.050 172.050 ;
        RECT 731.400 169.050 732.450 169.950 ;
        RECT 737.400 169.050 738.450 169.950 ;
        RECT 730.950 166.950 733.050 169.050 ;
        RECT 734.250 167.250 735.750 168.150 ;
        RECT 736.950 166.950 739.050 169.050 ;
        RECT 739.950 166.950 742.050 169.050 ;
        RECT 740.400 166.050 741.450 166.950 ;
        RECT 730.950 164.850 732.750 165.750 ;
        RECT 733.950 163.950 736.050 166.050 ;
        RECT 737.250 164.850 738.750 165.750 ;
        RECT 739.950 163.950 742.050 166.050 ;
        RECT 734.400 157.050 735.450 163.950 ;
        RECT 739.950 161.850 742.050 162.750 ;
        RECT 733.950 154.950 736.050 157.050 ;
        RECT 736.950 136.950 739.050 139.050 ;
        RECT 728.400 131.400 732.450 132.450 ;
        RECT 718.950 130.950 721.050 131.400 ;
        RECT 721.950 130.950 724.050 131.400 ;
        RECT 706.950 127.950 709.050 130.050 ;
        RECT 712.950 129.450 715.050 130.050 ;
        RECT 721.950 129.450 724.050 130.050 ;
        RECT 710.250 128.250 711.750 129.150 ;
        RECT 712.950 128.400 717.450 129.450 ;
        RECT 712.950 127.950 715.050 128.400 ;
        RECT 706.950 125.850 708.750 126.750 ;
        RECT 709.950 124.950 712.050 127.050 ;
        RECT 713.250 125.850 715.050 126.750 ;
        RECT 710.400 124.050 711.450 124.950 ;
        RECT 709.950 121.950 712.050 124.050 ;
        RECT 716.400 121.050 717.450 128.400 ;
        RECT 719.400 128.400 724.050 129.450 ;
        RECT 719.400 124.050 720.450 128.400 ;
        RECT 721.950 127.950 724.050 128.400 ;
        RECT 725.250 128.250 726.750 129.150 ;
        RECT 727.950 127.950 730.050 130.050 ;
        RECT 721.950 125.850 723.750 126.750 ;
        RECT 724.950 124.950 727.050 127.050 ;
        RECT 728.250 125.850 730.050 126.750 ;
        RECT 718.950 121.950 721.050 124.050 ;
        RECT 706.950 118.950 709.050 121.050 ;
        RECT 715.950 118.950 718.050 121.050 ;
        RECT 718.950 118.950 721.050 121.050 ;
        RECT 707.400 94.050 708.450 118.950 ;
        RECT 716.400 118.050 717.450 118.950 ;
        RECT 719.400 118.050 720.450 118.950 ;
        RECT 715.950 115.950 718.050 118.050 ;
        RECT 718.950 115.950 721.050 118.050 ;
        RECT 725.400 106.050 726.450 124.950 ;
        RECT 727.950 112.950 730.050 115.050 ;
        RECT 709.950 103.950 712.050 106.050 ;
        RECT 724.950 103.950 727.050 106.050 ;
        RECT 710.400 97.050 711.450 103.950 ;
        RECT 718.950 100.950 721.050 103.050 ;
        RECT 719.400 97.050 720.450 100.950 ;
        RECT 709.950 94.950 712.050 97.050 ;
        RECT 715.950 95.250 717.750 96.150 ;
        RECT 718.950 94.950 721.050 97.050 ;
        RECT 724.950 95.250 727.050 96.150 ;
        RECT 706.950 91.950 709.050 94.050 ;
        RECT 709.950 92.850 712.050 93.750 ;
        RECT 715.950 91.950 718.050 94.050 ;
        RECT 719.250 92.850 721.050 93.750 ;
        RECT 724.950 91.950 727.050 94.050 ;
        RECT 716.400 70.050 717.450 91.950 ;
        RECT 709.950 67.950 712.050 70.050 ;
        RECT 715.950 67.950 718.050 70.050 ;
        RECT 704.400 62.400 708.450 63.450 ;
        RECT 703.950 58.950 706.050 61.050 ;
        RECT 704.400 58.050 705.450 58.950 ;
        RECT 707.400 58.050 708.450 62.400 ;
        RECT 697.950 55.950 700.050 58.050 ;
        RECT 701.250 56.250 702.750 57.150 ;
        RECT 703.950 55.950 706.050 58.050 ;
        RECT 706.950 55.950 709.050 58.050 ;
        RECT 710.400 55.050 711.450 67.950 ;
        RECT 712.950 60.450 715.050 61.050 ;
        RECT 712.950 59.400 717.450 60.450 ;
        RECT 712.950 58.950 715.050 59.400 ;
        RECT 716.400 58.050 717.450 59.400 ;
        RECT 721.950 59.250 724.050 60.150 ;
        RECT 715.950 55.950 718.050 58.050 ;
        RECT 719.250 56.250 720.750 57.150 ;
        RECT 721.950 55.950 724.050 58.050 ;
        RECT 725.250 56.250 727.050 57.150 ;
        RECT 697.950 53.850 699.750 54.750 ;
        RECT 700.950 52.950 703.050 55.050 ;
        RECT 704.250 53.850 706.050 54.750 ;
        RECT 709.950 52.950 712.050 55.050 ;
        RECT 715.950 53.850 717.750 54.750 ;
        RECT 718.950 52.950 721.050 55.050 ;
        RECT 719.400 46.050 720.450 52.950 ;
        RECT 718.950 43.950 721.050 46.050 ;
        RECT 706.950 40.950 709.050 43.050 ;
        RECT 703.950 31.950 706.050 34.050 ;
        RECT 697.950 25.950 700.050 28.050 ;
        RECT 679.950 22.950 682.050 25.050 ;
        RECT 683.250 23.850 684.750 24.750 ;
        RECT 685.950 22.950 688.050 25.050 ;
        RECT 694.950 22.950 697.050 25.050 ;
        RECT 698.250 23.850 699.750 24.750 ;
        RECT 700.950 22.950 703.050 25.050 ;
        RECT 661.950 19.950 664.050 22.050 ;
        RECT 667.950 19.950 670.050 22.050 ;
        RECT 671.250 20.850 673.050 21.750 ;
        RECT 673.950 19.950 676.050 22.050 ;
        RECT 679.950 20.850 682.050 21.750 ;
        RECT 685.950 20.850 688.050 21.750 ;
        RECT 694.950 20.850 697.050 21.750 ;
        RECT 700.950 20.850 703.050 21.750 ;
        RECT 662.400 19.050 663.450 19.950 ;
        RECT 652.950 17.400 657.450 18.450 ;
        RECT 652.950 16.950 655.050 17.400 ;
        RECT 661.950 16.950 664.050 19.050 ;
        RECT 704.400 16.050 705.450 31.950 ;
        RECT 707.400 19.050 708.450 40.950 ;
        RECT 712.950 22.950 715.050 25.050 ;
        RECT 713.400 22.050 714.450 22.950 ;
        RECT 709.950 20.250 711.750 21.150 ;
        RECT 712.950 19.950 715.050 22.050 ;
        RECT 716.250 20.250 718.050 21.150 ;
        RECT 718.950 19.950 721.050 22.050 ;
        RECT 706.950 16.950 709.050 19.050 ;
        RECT 709.950 16.950 712.050 19.050 ;
        RECT 713.250 17.850 714.750 18.750 ;
        RECT 715.950 18.450 718.050 19.050 ;
        RECT 719.400 18.450 720.450 19.950 ;
        RECT 715.950 17.400 720.450 18.450 ;
        RECT 715.950 16.950 718.050 17.400 ;
        RECT 710.400 16.050 711.450 16.950 ;
        RECT 722.400 16.050 723.450 55.950 ;
        RECT 724.950 52.950 727.050 55.050 ;
        RECT 725.400 43.050 726.450 52.950 ;
        RECT 728.400 52.050 729.450 112.950 ;
        RECT 731.400 94.050 732.450 131.400 ;
        RECT 733.950 130.950 736.050 133.050 ;
        RECT 730.950 91.950 733.050 94.050 ;
        RECT 731.400 79.050 732.450 91.950 ;
        RECT 730.950 76.950 733.050 79.050 ;
        RECT 730.950 52.950 733.050 55.050 ;
        RECT 727.950 49.950 730.050 52.050 ;
        RECT 731.400 49.050 732.450 52.950 ;
        RECT 730.950 46.950 733.050 49.050 ;
        RECT 734.400 46.050 735.450 130.950 ;
        RECT 737.400 130.050 738.450 136.950 ;
        RECT 743.400 133.050 744.450 169.950 ;
        RECT 746.400 166.050 747.450 190.950 ;
        RECT 745.950 163.950 748.050 166.050 ;
        RECT 742.950 130.950 745.050 133.050 ;
        RECT 736.950 127.950 739.050 130.050 ;
        RECT 740.250 128.250 741.750 129.150 ;
        RECT 742.950 127.950 745.050 130.050 ;
        RECT 736.950 125.850 738.750 126.750 ;
        RECT 739.950 124.950 742.050 127.050 ;
        RECT 743.250 125.850 745.050 126.750 ;
        RECT 740.400 118.050 741.450 124.950 ;
        RECT 739.950 115.950 742.050 118.050 ;
        RECT 739.950 94.950 742.050 97.050 ;
        RECT 740.400 94.050 741.450 94.950 ;
        RECT 736.950 92.250 738.750 93.150 ;
        RECT 739.950 91.950 742.050 94.050 ;
        RECT 743.250 92.250 745.050 93.150 ;
        RECT 736.950 88.950 739.050 91.050 ;
        RECT 740.250 89.850 741.750 90.750 ;
        RECT 742.950 88.950 745.050 91.050 ;
        RECT 737.400 87.450 738.450 88.950 ;
        RECT 737.400 86.400 741.450 87.450 ;
        RECT 736.950 50.850 739.050 51.750 ;
        RECT 733.950 43.950 736.050 46.050 ;
        RECT 724.950 40.950 727.050 43.050 ;
        RECT 727.950 22.950 730.050 25.050 ;
        RECT 728.400 22.050 729.450 22.950 ;
        RECT 740.400 22.050 741.450 86.400 ;
        RECT 743.400 82.050 744.450 88.950 ;
        RECT 742.950 79.950 745.050 82.050 ;
        RECT 746.400 55.050 747.450 163.950 ;
        RECT 749.400 163.050 750.450 208.950 ;
        RECT 770.400 201.450 771.450 235.950 ;
        RECT 775.950 233.850 778.050 234.750 ;
        RECT 754.950 200.250 757.050 201.150 ;
        RECT 767.400 200.400 771.450 201.450 ;
        RECT 751.950 196.950 754.050 199.050 ;
        RECT 754.950 196.950 757.050 199.050 ;
        RECT 758.250 197.250 759.750 198.150 ;
        RECT 760.950 196.950 763.050 199.050 ;
        RECT 764.250 197.250 766.050 198.150 ;
        RECT 752.400 184.050 753.450 196.950 ;
        RECT 755.400 193.050 756.450 196.950 ;
        RECT 757.950 193.950 760.050 196.050 ;
        RECT 761.250 194.850 762.750 195.750 ;
        RECT 763.950 193.950 766.050 196.050 ;
        RECT 754.950 190.950 757.050 193.050 ;
        RECT 760.950 184.950 763.050 187.050 ;
        RECT 751.950 181.950 754.050 184.050 ;
        RECT 754.950 181.950 757.050 184.050 ;
        RECT 755.400 172.050 756.450 181.950 ;
        RECT 757.950 172.950 760.050 175.050 ;
        RECT 751.950 169.950 754.050 172.050 ;
        RECT 754.950 169.950 757.050 172.050 ;
        RECT 752.400 169.050 753.450 169.950 ;
        RECT 758.400 169.050 759.450 172.950 ;
        RECT 751.950 166.950 754.050 169.050 ;
        RECT 755.250 167.850 756.750 168.750 ;
        RECT 757.950 166.950 760.050 169.050 ;
        RECT 751.950 164.850 754.050 165.750 ;
        RECT 757.950 164.850 760.050 165.750 ;
        RECT 748.950 160.950 751.050 163.050 ;
        RECT 761.400 145.050 762.450 184.950 ;
        RECT 763.950 172.950 766.050 175.050 ;
        RECT 764.400 163.050 765.450 172.950 ;
        RECT 767.400 172.050 768.450 200.400 ;
        RECT 778.950 199.950 781.050 202.050 ;
        RECT 769.950 197.250 772.050 198.150 ;
        RECT 775.950 197.250 778.050 198.150 ;
        RECT 769.950 193.950 772.050 196.050 ;
        RECT 773.250 194.250 774.750 195.150 ;
        RECT 775.950 193.950 778.050 196.050 ;
        RECT 770.400 172.050 771.450 193.950 ;
        RECT 772.950 190.950 775.050 193.050 ;
        RECT 773.400 181.050 774.450 190.950 ;
        RECT 776.400 184.050 777.450 193.950 ;
        RECT 775.950 181.950 778.050 184.050 ;
        RECT 772.950 178.950 775.050 181.050 ;
        RECT 772.950 172.950 775.050 175.050 ;
        RECT 766.950 169.950 769.050 172.050 ;
        RECT 769.950 169.950 772.050 172.050 ;
        RECT 773.400 169.050 774.450 172.950 ;
        RECT 775.950 169.950 778.050 172.050 ;
        RECT 779.400 171.450 780.450 199.950 ;
        RECT 782.400 175.050 783.450 286.950 ;
        RECT 784.950 271.950 787.050 274.050 ;
        RECT 784.950 269.850 787.050 270.750 ;
        RECT 788.400 259.050 789.450 295.950 ;
        RECT 790.950 272.250 793.050 273.150 ;
        RECT 790.950 265.950 793.050 268.050 ;
        RECT 787.950 256.950 790.050 259.050 ;
        RECT 784.950 250.950 787.050 253.050 ;
        RECT 785.400 196.050 786.450 250.950 ;
        RECT 791.400 241.050 792.450 265.950 ;
        RECT 794.400 244.050 795.450 334.950 ;
        RECT 812.400 334.050 813.450 337.950 ;
        RECT 811.950 331.950 814.050 334.050 ;
        RECT 818.400 331.050 819.450 337.950 ;
        RECT 811.950 328.950 814.050 331.050 ;
        RECT 817.950 328.950 820.050 331.050 ;
        RECT 805.950 316.950 808.050 319.050 ;
        RECT 796.950 310.950 799.050 313.050 ;
        RECT 797.400 286.050 798.450 310.950 ;
        RECT 799.950 308.250 801.750 309.150 ;
        RECT 802.950 307.950 805.050 310.050 ;
        RECT 806.400 307.050 807.450 316.950 ;
        RECT 812.400 313.050 813.450 328.950 ;
        RECT 821.400 324.450 822.450 347.400 ;
        RECT 827.400 346.050 828.450 352.950 ;
        RECT 829.950 346.950 832.050 349.050 ;
        RECT 823.950 343.950 826.050 346.050 ;
        RECT 826.950 343.950 829.050 346.050 ;
        RECT 824.400 337.050 825.450 343.950 ;
        RECT 830.400 343.050 831.450 346.950 ;
        RECT 835.950 343.950 838.050 346.050 ;
        RECT 826.950 341.250 829.050 342.150 ;
        RECT 829.950 340.950 832.050 343.050 ;
        RECT 832.950 341.250 835.050 342.150 ;
        RECT 826.950 337.950 829.050 340.050 ;
        RECT 830.250 338.250 831.750 339.150 ;
        RECT 832.950 337.950 835.050 340.050 ;
        RECT 823.950 334.950 826.050 337.050 ;
        RECT 826.950 334.950 829.050 337.050 ;
        RECT 829.950 334.950 832.050 337.050 ;
        RECT 823.950 331.950 826.050 334.050 ;
        RECT 818.400 323.400 822.450 324.450 ;
        RECT 811.950 310.950 814.050 313.050 ;
        RECT 814.950 311.250 817.050 312.150 ;
        RECT 808.950 309.450 811.050 310.050 ;
        RECT 808.950 308.400 813.450 309.450 ;
        RECT 808.950 307.950 811.050 308.400 ;
        RECT 799.950 304.950 802.050 307.050 ;
        RECT 803.250 305.850 804.750 306.750 ;
        RECT 805.950 304.950 808.050 307.050 ;
        RECT 809.250 305.850 811.050 306.750 ;
        RECT 805.950 302.850 808.050 303.750 ;
        RECT 812.400 301.050 813.450 308.400 ;
        RECT 814.950 307.950 817.050 310.050 ;
        RECT 808.950 298.950 811.050 301.050 ;
        RECT 811.950 298.950 814.050 301.050 ;
        RECT 796.950 283.950 799.050 286.050 ;
        RECT 805.950 283.950 808.050 286.050 ;
        RECT 796.950 280.950 799.050 283.050 ;
        RECT 799.950 280.950 802.050 283.050 ;
        RECT 802.950 280.950 805.050 283.050 ;
        RECT 797.550 262.050 798.750 280.950 ;
        RECT 800.550 276.750 801.750 280.950 ;
        RECT 799.950 274.650 802.050 276.750 ;
        RECT 800.550 262.050 801.750 274.650 ;
        RECT 803.550 262.050 804.750 280.950 ;
        RECT 806.400 264.450 807.450 283.950 ;
        RECT 809.400 271.050 810.450 298.950 ;
        RECT 818.400 289.050 819.450 323.400 ;
        RECT 820.950 319.950 823.050 322.050 ;
        RECT 821.400 316.050 822.450 319.950 ;
        RECT 824.400 316.050 825.450 331.950 ;
        RECT 827.400 318.450 828.450 334.950 ;
        RECT 830.400 331.050 831.450 334.950 ;
        RECT 829.950 328.950 832.050 331.050 ;
        RECT 833.400 328.050 834.450 337.950 ;
        RECT 836.400 334.050 837.450 343.950 ;
        RECT 842.400 343.050 843.450 365.400 ;
        RECT 838.950 341.250 841.050 342.150 ;
        RECT 841.950 340.950 844.050 343.050 ;
        RECT 844.950 341.250 847.050 342.150 ;
        RECT 838.950 337.950 841.050 340.050 ;
        RECT 842.250 338.250 843.750 339.150 ;
        RECT 844.950 337.950 847.050 340.050 ;
        RECT 835.950 331.950 838.050 334.050 ;
        RECT 839.400 331.050 840.450 337.950 ;
        RECT 841.950 334.950 844.050 337.050 ;
        RECT 844.950 334.950 847.050 337.050 ;
        RECT 842.400 334.050 843.450 334.950 ;
        RECT 841.950 331.950 844.050 334.050 ;
        RECT 838.950 328.950 841.050 331.050 ;
        RECT 841.950 328.950 844.050 331.050 ;
        RECT 832.950 325.950 835.050 328.050 ;
        RECT 832.950 319.950 835.050 322.050 ;
        RECT 827.400 317.400 831.450 318.450 ;
        RECT 820.950 313.950 823.050 316.050 ;
        RECT 823.950 315.450 826.050 316.050 ;
        RECT 823.950 314.400 828.450 315.450 ;
        RECT 823.950 313.950 826.050 314.400 ;
        RECT 821.400 313.050 822.450 313.950 ;
        RECT 820.950 310.950 823.050 313.050 ;
        RECT 824.250 311.850 826.050 312.750 ;
        RECT 820.950 308.850 823.050 309.750 ;
        RECT 823.950 307.950 826.050 310.050 ;
        RECT 820.950 304.950 823.050 307.050 ;
        RECT 821.400 292.050 822.450 304.950 ;
        RECT 824.400 298.050 825.450 307.950 ;
        RECT 827.400 301.050 828.450 314.400 ;
        RECT 826.950 298.950 829.050 301.050 ;
        RECT 823.950 295.950 826.050 298.050 ;
        RECT 820.950 289.950 823.050 292.050 ;
        RECT 817.950 286.950 820.050 289.050 ;
        RECT 830.400 286.050 831.450 317.400 ;
        RECT 833.400 313.050 834.450 319.950 ;
        RECT 835.950 316.950 838.050 319.050 ;
        RECT 832.950 310.950 835.050 313.050 ;
        RECT 836.400 310.050 837.450 316.950 ;
        RECT 832.950 308.250 834.750 309.150 ;
        RECT 835.950 307.950 838.050 310.050 ;
        RECT 839.250 308.250 841.050 309.150 ;
        RECT 832.950 304.950 835.050 307.050 ;
        RECT 836.250 305.850 837.750 306.750 ;
        RECT 838.950 304.950 841.050 307.050 ;
        RECT 839.400 301.050 840.450 304.950 ;
        RECT 838.950 298.950 841.050 301.050 ;
        RECT 832.950 295.950 835.050 298.050 ;
        RECT 829.950 283.950 832.050 286.050 ;
        RECT 827.100 281.100 829.200 283.200 ;
        RECT 811.950 278.400 814.050 280.500 ;
        RECT 816.000 278.400 818.100 280.500 ;
        RECT 823.950 278.850 826.050 280.950 ;
        RECT 812.250 272.250 813.450 278.400 ;
        RECT 808.950 268.950 811.050 271.050 ;
        RECT 811.950 270.150 814.050 272.250 ;
        RECT 808.950 266.250 811.050 267.150 ;
        RECT 808.950 264.450 811.050 265.050 ;
        RECT 806.400 263.400 811.050 264.450 ;
        RECT 808.950 262.950 811.050 263.400 ;
        RECT 796.950 259.950 799.050 262.050 ;
        RECT 799.950 259.950 802.050 262.050 ;
        RECT 802.950 259.950 805.050 262.050 ;
        RECT 808.950 259.950 811.050 262.050 ;
        RECT 812.250 261.600 813.450 270.150 ;
        RECT 816.450 269.550 817.650 278.400 ;
        RECT 820.950 275.250 823.050 277.350 ;
        RECT 816.150 267.450 818.250 269.550 ;
        RECT 816.450 261.600 817.650 267.450 ;
        RECT 821.400 261.600 822.600 275.250 ;
        RECT 824.550 261.600 825.750 278.850 ;
        RECT 827.250 277.350 828.450 281.100 ;
        RECT 826.950 275.250 829.050 277.350 ;
        RECT 827.250 261.600 828.450 275.250 ;
        RECT 829.950 274.950 832.050 277.050 ;
        RECT 802.950 256.950 805.050 259.050 ;
        RECT 805.950 256.950 808.050 259.050 ;
        RECT 803.400 244.050 804.450 256.950 ;
        RECT 806.400 244.050 807.450 256.950 ;
        RECT 809.400 252.450 810.450 259.950 ;
        RECT 811.950 259.500 814.050 261.600 ;
        RECT 816.150 259.500 818.250 261.600 ;
        RECT 820.950 259.500 823.050 261.600 ;
        RECT 823.950 259.500 826.050 261.600 ;
        RECT 826.950 259.500 829.050 261.600 ;
        RECT 814.950 253.950 817.050 256.050 ;
        RECT 817.950 253.950 820.050 256.050 ;
        RECT 809.400 251.400 813.450 252.450 ;
        RECT 808.950 247.950 811.050 250.050 ;
        RECT 793.950 241.950 796.050 244.050 ;
        RECT 799.950 241.950 802.050 244.050 ;
        RECT 802.950 241.950 805.050 244.050 ;
        RECT 805.950 241.950 808.050 244.050 ;
        RECT 787.950 238.950 790.050 241.050 ;
        RECT 790.950 238.950 793.050 241.050 ;
        RECT 794.250 239.250 795.750 240.150 ;
        RECT 796.950 238.950 799.050 241.050 ;
        RECT 788.400 238.050 789.450 238.950 ;
        RECT 787.950 235.950 790.050 238.050 ;
        RECT 791.250 236.850 792.750 237.750 ;
        RECT 793.950 235.950 796.050 238.050 ;
        RECT 797.250 236.850 799.050 237.750 ;
        RECT 787.950 233.850 790.050 234.750 ;
        RECT 787.950 229.950 790.050 232.050 ;
        RECT 788.400 205.050 789.450 229.950 ;
        RECT 787.950 202.950 790.050 205.050 ;
        RECT 788.400 199.050 789.450 202.950 ;
        RECT 787.950 196.950 790.050 199.050 ;
        RECT 793.950 197.250 796.050 198.150 ;
        RECT 784.950 193.950 787.050 196.050 ;
        RECT 787.950 194.850 790.050 195.750 ;
        RECT 793.950 193.950 796.050 196.050 ;
        RECT 797.250 194.250 799.050 195.150 ;
        RECT 781.950 172.950 784.050 175.050 ;
        RECT 779.400 170.400 783.450 171.450 ;
        RECT 766.950 166.950 769.050 169.050 ;
        RECT 770.250 167.850 771.750 168.750 ;
        RECT 772.950 166.950 775.050 169.050 ;
        RECT 766.950 164.850 769.050 165.750 ;
        RECT 772.950 164.850 775.050 165.750 ;
        RECT 763.950 160.950 766.050 163.050 ;
        RECT 748.950 142.950 751.050 145.050 ;
        RECT 760.950 142.950 763.050 145.050 ;
        RECT 749.400 91.050 750.450 142.950 ;
        RECT 754.950 136.950 757.050 139.050 ;
        RECT 751.950 133.950 754.050 136.050 ;
        RECT 752.400 115.050 753.450 133.950 ;
        RECT 751.950 112.950 754.050 115.050 ;
        RECT 755.400 100.050 756.450 136.950 ;
        RECT 776.400 127.050 777.450 169.950 ;
        RECT 778.950 167.250 781.050 168.150 ;
        RECT 778.950 163.950 781.050 166.050 ;
        RECT 779.400 163.050 780.450 163.950 ;
        RECT 778.950 160.950 781.050 163.050 ;
        RECT 782.400 154.050 783.450 170.400 ;
        RECT 785.400 169.050 786.450 193.950 ;
        RECT 794.400 184.050 795.450 193.950 ;
        RECT 796.950 190.950 799.050 193.050 ;
        RECT 797.400 190.050 798.450 190.950 ;
        RECT 796.950 187.950 799.050 190.050 ;
        RECT 800.400 187.050 801.450 241.950 ;
        RECT 809.400 241.050 810.450 247.950 ;
        RECT 802.950 238.950 805.050 241.050 ;
        RECT 806.250 239.850 807.750 240.750 ;
        RECT 808.950 238.950 811.050 241.050 ;
        RECT 802.950 236.850 805.050 237.750 ;
        RECT 808.950 236.850 811.050 237.750 ;
        RECT 808.950 232.950 811.050 235.050 ;
        RECT 805.950 226.950 808.050 229.050 ;
        RECT 806.400 199.050 807.450 226.950 ;
        RECT 805.950 196.950 808.050 199.050 ;
        RECT 805.950 194.850 808.050 195.750 ;
        RECT 809.400 193.050 810.450 232.950 ;
        RECT 812.400 202.050 813.450 251.400 ;
        RECT 815.400 235.050 816.450 253.950 ;
        RECT 814.950 232.950 817.050 235.050 ;
        RECT 811.950 199.950 814.050 202.050 ;
        RECT 811.950 197.250 814.050 198.150 ;
        RECT 811.950 193.950 814.050 196.050 ;
        RECT 815.250 194.250 817.050 195.150 ;
        RECT 808.950 190.950 811.050 193.050 ;
        RECT 812.400 187.050 813.450 193.950 ;
        RECT 814.950 190.950 817.050 193.050 ;
        RECT 799.950 184.950 802.050 187.050 ;
        RECT 811.950 184.950 814.050 187.050 ;
        RECT 793.950 181.950 796.050 184.050 ;
        RECT 818.400 181.050 819.450 253.950 ;
        RECT 823.950 250.950 826.050 253.050 ;
        RECT 824.400 241.050 825.450 250.950 ;
        RECT 823.950 240.450 826.050 241.050 ;
        RECT 821.400 239.400 826.050 240.450 ;
        RECT 821.400 220.050 822.450 239.400 ;
        RECT 823.950 238.950 826.050 239.400 ;
        RECT 827.250 239.250 829.050 240.150 ;
        RECT 823.950 236.850 825.750 237.750 ;
        RECT 826.950 235.950 829.050 238.050 ;
        RECT 823.950 232.950 826.050 235.050 ;
        RECT 820.950 217.950 823.050 220.050 ;
        RECT 820.950 211.950 823.050 214.050 ;
        RECT 817.950 178.950 820.050 181.050 ;
        RECT 817.950 175.950 820.050 178.050 ;
        RECT 787.950 172.950 790.050 175.050 ;
        RECT 799.950 173.400 802.050 175.500 ;
        RECT 802.950 173.400 805.050 175.500 ;
        RECT 805.950 173.400 808.050 175.500 ;
        RECT 810.750 173.400 812.850 175.500 ;
        RECT 814.950 173.400 817.050 175.500 ;
        RECT 784.950 166.950 787.050 169.050 ;
        RECT 781.950 151.950 784.050 154.050 ;
        RECT 785.400 130.050 786.450 166.950 ;
        RECT 781.950 128.250 784.050 129.150 ;
        RECT 784.950 127.950 787.050 130.050 ;
        RECT 757.950 125.250 760.050 126.150 ;
        RECT 763.950 125.250 766.050 126.150 ;
        RECT 772.950 125.250 774.750 126.150 ;
        RECT 775.950 124.950 778.050 127.050 ;
        RECT 779.250 125.250 780.750 126.150 ;
        RECT 781.950 124.950 784.050 127.050 ;
        RECT 757.950 121.950 760.050 124.050 ;
        RECT 761.250 122.250 762.750 123.150 ;
        RECT 763.950 121.950 766.050 124.050 ;
        RECT 772.950 121.950 775.050 124.050 ;
        RECT 776.250 122.850 777.750 123.750 ;
        RECT 778.950 121.950 781.050 124.050 ;
        RECT 757.950 118.950 760.050 121.050 ;
        RECT 760.950 118.950 763.050 121.050 ;
        RECT 754.950 97.950 757.050 100.050 ;
        RECT 751.950 95.250 754.050 96.150 ;
        RECT 754.950 95.850 757.050 96.750 ;
        RECT 758.400 96.450 759.450 118.950 ;
        RECT 761.400 118.050 762.450 118.950 ;
        RECT 760.950 115.950 763.050 118.050 ;
        RECT 764.400 115.050 765.450 121.950 ;
        RECT 773.400 115.050 774.450 121.950 ;
        RECT 763.950 112.950 766.050 115.050 ;
        RECT 772.950 112.950 775.050 115.050 ;
        RECT 775.950 112.950 778.050 115.050 ;
        RECT 760.950 100.950 763.050 103.050 ;
        RECT 766.950 100.950 769.050 103.050 ;
        RECT 769.950 100.950 772.050 103.050 ;
        RECT 761.400 100.050 762.450 100.950 ;
        RECT 760.950 97.950 763.050 100.050 ;
        RECT 767.400 97.050 768.450 100.950 ;
        RECT 760.950 96.450 763.050 97.050 ;
        RECT 758.400 95.400 763.050 96.450 ;
        RECT 751.950 93.450 754.050 94.050 ;
        RECT 758.400 93.450 759.450 95.400 ;
        RECT 760.950 94.950 763.050 95.400 ;
        RECT 764.250 95.250 765.750 96.150 ;
        RECT 766.950 94.950 769.050 97.050 ;
        RECT 770.400 94.050 771.450 100.950 ;
        RECT 772.950 97.950 775.050 100.050 ;
        RECT 751.950 92.400 759.450 93.450 ;
        RECT 760.950 92.850 762.750 93.750 ;
        RECT 751.950 91.950 754.050 92.400 ;
        RECT 763.950 91.950 766.050 94.050 ;
        RECT 767.250 92.850 768.750 93.750 ;
        RECT 769.950 91.950 772.050 94.050 ;
        RECT 748.950 88.950 751.050 91.050 ;
        RECT 757.950 88.950 760.050 91.050 ;
        RECT 766.950 88.950 769.050 91.050 ;
        RECT 769.950 89.850 772.050 90.750 ;
        RECT 751.950 79.950 754.050 82.050 ;
        RECT 745.950 52.950 748.050 55.050 ;
        RECT 745.950 43.950 748.050 46.050 ;
        RECT 724.950 20.250 726.750 21.150 ;
        RECT 727.950 19.950 730.050 22.050 ;
        RECT 731.250 20.250 733.050 21.150 ;
        RECT 733.950 19.950 736.050 22.050 ;
        RECT 736.950 20.250 738.750 21.150 ;
        RECT 739.950 19.950 742.050 22.050 ;
        RECT 743.250 20.250 745.050 21.150 ;
        RECT 724.950 16.950 727.050 19.050 ;
        RECT 728.250 17.850 729.750 18.750 ;
        RECT 730.950 18.450 733.050 19.050 ;
        RECT 734.400 18.450 735.450 19.950 ;
        RECT 730.950 17.400 735.450 18.450 ;
        RECT 730.950 16.950 733.050 17.400 ;
        RECT 736.950 16.950 739.050 19.050 ;
        RECT 740.250 17.850 741.750 18.750 ;
        RECT 742.950 18.450 745.050 19.050 ;
        RECT 746.400 18.450 747.450 43.950 ;
        RECT 752.400 22.050 753.450 79.950 ;
        RECT 758.400 60.450 759.450 88.950 ;
        RECT 758.400 59.400 762.450 60.450 ;
        RECT 757.950 52.950 760.050 55.050 ;
        RECT 757.950 50.850 760.050 51.750 ;
        RECT 761.400 49.050 762.450 59.400 ;
        RECT 767.400 55.050 768.450 88.950 ;
        RECT 773.400 73.050 774.450 97.950 ;
        RECT 776.400 97.050 777.450 112.950 ;
        RECT 779.400 100.050 780.450 121.950 ;
        RECT 785.400 121.050 786.450 127.950 ;
        RECT 788.400 127.050 789.450 172.950 ;
        RECT 790.950 163.950 793.050 166.050 ;
        RECT 790.950 161.850 793.050 162.750 ;
        RECT 800.550 159.750 801.750 173.400 ;
        RECT 799.950 157.650 802.050 159.750 ;
        RECT 800.550 153.900 801.750 157.650 ;
        RECT 803.250 156.150 804.450 173.400 ;
        RECT 806.400 159.750 807.600 173.400 ;
        RECT 811.350 167.550 812.550 173.400 ;
        RECT 810.750 165.450 812.850 167.550 ;
        RECT 805.950 157.650 808.050 159.750 ;
        RECT 811.350 156.600 812.550 165.450 ;
        RECT 815.550 164.850 816.750 173.400 ;
        RECT 818.400 172.050 819.450 175.950 ;
        RECT 817.950 169.950 820.050 172.050 ;
        RECT 817.950 167.850 820.050 168.750 ;
        RECT 814.950 162.750 817.050 164.850 ;
        RECT 821.400 163.050 822.450 211.950 ;
        RECT 824.400 202.050 825.450 232.950 ;
        RECT 827.400 226.050 828.450 235.950 ;
        RECT 830.400 235.050 831.450 274.950 ;
        RECT 833.400 256.050 834.450 295.950 ;
        RECT 838.950 292.950 841.050 295.050 ;
        RECT 835.950 283.950 838.050 286.050 ;
        RECT 836.400 277.050 837.450 283.950 ;
        RECT 835.950 274.950 838.050 277.050 ;
        RECT 835.950 272.250 838.050 273.150 ;
        RECT 839.400 271.050 840.450 292.950 ;
        RECT 835.950 268.950 838.050 271.050 ;
        RECT 838.950 268.950 841.050 271.050 ;
        RECT 832.950 253.950 835.050 256.050 ;
        RECT 836.400 247.050 837.450 268.950 ;
        RECT 835.950 244.950 838.050 247.050 ;
        RECT 835.950 241.950 838.050 244.050 ;
        RECT 836.400 241.050 837.450 241.950 ;
        RECT 832.950 239.250 834.750 240.150 ;
        RECT 835.950 238.950 838.050 241.050 ;
        RECT 832.950 235.950 835.050 238.050 ;
        RECT 836.250 236.850 838.050 237.750 ;
        RECT 829.950 232.950 832.050 235.050 ;
        RECT 839.400 226.050 840.450 268.950 ;
        RECT 842.400 238.050 843.450 328.950 ;
        RECT 845.400 259.050 846.450 334.950 ;
        RECT 848.400 316.050 849.450 373.950 ;
        RECT 851.400 367.050 852.450 604.950 ;
        RECT 854.400 529.050 855.450 626.400 ;
        RECT 856.950 622.950 859.050 625.050 ;
        RECT 853.950 526.950 856.050 529.050 ;
        RECT 853.950 524.250 856.050 525.150 ;
        RECT 853.950 520.950 856.050 523.050 ;
        RECT 854.400 496.050 855.450 520.950 ;
        RECT 853.950 493.950 856.050 496.050 ;
        RECT 853.950 490.950 856.050 493.050 ;
        RECT 854.400 412.050 855.450 490.950 ;
        RECT 857.400 448.050 858.450 622.950 ;
        RECT 860.400 580.050 861.450 635.400 ;
        RECT 859.950 577.950 862.050 580.050 ;
        RECT 859.950 502.950 862.050 505.050 ;
        RECT 856.950 445.950 859.050 448.050 ;
        RECT 853.950 409.950 856.050 412.050 ;
        RECT 856.950 388.950 859.050 391.050 ;
        RECT 857.400 388.050 858.450 388.950 ;
        RECT 856.950 385.950 859.050 388.050 ;
        RECT 853.950 382.950 856.050 385.050 ;
        RECT 857.250 383.850 859.050 384.750 ;
        RECT 853.950 380.850 856.050 381.750 ;
        RECT 856.950 379.950 859.050 382.050 ;
        RECT 853.950 376.950 856.050 379.050 ;
        RECT 850.950 364.950 853.050 367.050 ;
        RECT 850.950 337.950 853.050 340.050 ;
        RECT 851.400 316.050 852.450 337.950 ;
        RECT 854.400 331.050 855.450 376.950 ;
        RECT 857.400 373.050 858.450 379.950 ;
        RECT 856.950 370.950 859.050 373.050 ;
        RECT 856.950 367.950 859.050 370.050 ;
        RECT 853.950 328.950 856.050 331.050 ;
        RECT 853.950 322.950 856.050 325.050 ;
        RECT 847.950 313.950 850.050 316.050 ;
        RECT 850.950 313.950 853.050 316.050 ;
        RECT 854.400 313.050 855.450 322.950 ;
        RECT 847.950 310.950 850.050 313.050 ;
        RECT 851.250 311.850 852.750 312.750 ;
        RECT 853.950 310.950 856.050 313.050 ;
        RECT 847.950 308.850 850.050 309.750 ;
        RECT 853.950 308.850 856.050 309.750 ;
        RECT 853.950 304.950 856.050 307.050 ;
        RECT 850.950 301.950 853.050 304.050 ;
        RECT 847.950 268.950 850.050 271.050 ;
        RECT 847.950 266.850 850.050 267.750 ;
        RECT 844.950 256.950 847.050 259.050 ;
        RECT 851.400 253.050 852.450 301.950 ;
        RECT 854.400 292.050 855.450 304.950 ;
        RECT 853.950 289.950 856.050 292.050 ;
        RECT 850.950 250.950 853.050 253.050 ;
        RECT 854.400 244.050 855.450 289.950 ;
        RECT 853.950 241.950 856.050 244.050 ;
        RECT 841.950 235.950 844.050 238.050 ;
        RECT 844.950 236.250 846.750 237.150 ;
        RECT 847.950 235.950 850.050 238.050 ;
        RECT 851.250 236.250 853.050 237.150 ;
        RECT 853.950 235.950 856.050 238.050 ;
        RECT 844.950 232.950 847.050 235.050 ;
        RECT 848.250 233.850 849.750 234.750 ;
        RECT 850.950 232.950 853.050 235.050 ;
        RECT 826.950 223.950 829.050 226.050 ;
        RECT 838.950 223.950 841.050 226.050 ;
        RECT 841.950 220.950 844.050 223.050 ;
        RECT 829.950 203.250 832.050 204.150 ;
        RECT 823.950 199.950 826.050 202.050 ;
        RECT 827.250 200.250 828.750 201.150 ;
        RECT 829.950 199.950 832.050 202.050 ;
        RECT 833.250 200.250 835.050 201.150 ;
        RECT 823.950 197.850 825.750 198.750 ;
        RECT 826.950 196.950 829.050 199.050 ;
        RECT 830.400 181.050 831.450 199.950 ;
        RECT 842.400 199.050 843.450 220.950 ;
        RECT 854.400 205.050 855.450 235.950 ;
        RECT 853.950 202.950 856.050 205.050 ;
        RECT 847.950 199.950 850.050 202.050 ;
        RECT 853.950 199.950 856.050 202.050 ;
        RECT 848.400 199.050 849.450 199.950 ;
        RECT 832.950 196.950 835.050 199.050 ;
        RECT 838.950 197.250 840.750 198.150 ;
        RECT 841.950 196.950 844.050 199.050 ;
        RECT 845.250 197.250 846.750 198.150 ;
        RECT 847.950 196.950 850.050 199.050 ;
        RECT 851.250 197.250 853.050 198.150 ;
        RECT 829.950 178.950 832.050 181.050 ;
        RECT 823.950 172.950 826.050 175.050 ;
        RECT 826.950 172.950 829.050 175.050 ;
        RECT 829.950 172.950 832.050 175.050 ;
        RECT 815.550 156.600 816.750 162.750 ;
        RECT 820.950 160.950 823.050 163.050 ;
        RECT 802.950 154.050 805.050 156.150 ;
        RECT 810.900 154.500 813.000 156.600 ;
        RECT 814.950 154.500 817.050 156.600 ;
        RECT 824.250 154.050 825.450 172.950 ;
        RECT 827.250 160.350 828.450 172.950 ;
        RECT 826.950 158.250 829.050 160.350 ;
        RECT 827.250 154.050 828.450 158.250 ;
        RECT 830.250 154.050 831.450 172.950 ;
        RECT 833.400 166.050 834.450 196.950 ;
        RECT 838.950 193.950 841.050 196.050 ;
        RECT 842.250 194.850 843.750 195.750 ;
        RECT 844.950 193.950 847.050 196.050 ;
        RECT 848.250 194.850 849.750 195.750 ;
        RECT 850.950 193.950 853.050 196.050 ;
        RECT 845.400 190.050 846.450 193.950 ;
        RECT 844.950 187.950 847.050 190.050 ;
        RECT 844.950 166.950 847.050 169.050 ;
        RECT 850.950 167.250 853.050 168.150 ;
        RECT 832.950 163.950 835.050 166.050 ;
        RECT 841.950 164.250 844.050 165.150 ;
        RECT 835.950 161.850 838.050 162.750 ;
        RECT 841.950 160.950 844.050 163.050 ;
        RECT 799.800 151.800 801.900 153.900 ;
        RECT 823.950 151.950 826.050 154.050 ;
        RECT 826.950 151.950 829.050 154.050 ;
        RECT 829.950 151.950 832.050 154.050 ;
        RECT 802.950 131.250 805.050 132.150 ;
        RECT 796.950 129.450 799.050 130.050 ;
        RECT 794.400 128.400 799.050 129.450 ;
        RECT 787.950 124.950 790.050 127.050 ;
        RECT 784.950 118.950 787.050 121.050 ;
        RECT 788.400 115.050 789.450 124.950 ;
        RECT 787.950 112.950 790.050 115.050 ;
        RECT 778.950 97.950 781.050 100.050 ;
        RECT 794.400 97.050 795.450 128.400 ;
        RECT 796.950 127.950 799.050 128.400 ;
        RECT 800.250 128.250 801.750 129.150 ;
        RECT 802.950 127.950 805.050 130.050 ;
        RECT 806.250 128.250 808.050 129.150 ;
        RECT 796.950 125.850 798.750 126.750 ;
        RECT 799.950 124.950 802.050 127.050 ;
        RECT 796.950 121.950 799.050 124.050 ;
        RECT 775.950 94.950 778.050 97.050 ;
        RECT 779.250 95.250 780.750 96.150 ;
        RECT 781.950 94.950 784.050 97.050 ;
        RECT 784.950 94.950 787.050 97.050 ;
        RECT 787.950 94.950 790.050 97.050 ;
        RECT 793.950 94.950 796.050 97.050 ;
        RECT 785.400 94.050 786.450 94.950 ;
        RECT 775.950 92.850 777.750 93.750 ;
        RECT 778.950 91.950 781.050 94.050 ;
        RECT 782.250 92.850 783.750 93.750 ;
        RECT 784.950 91.950 787.050 94.050 ;
        RECT 784.950 89.850 787.050 90.750 ;
        RECT 772.950 70.950 775.050 73.050 ;
        RECT 778.950 70.950 781.050 73.050 ;
        RECT 772.950 64.950 775.050 67.050 ;
        RECT 766.950 54.450 769.050 55.050 ;
        RECT 764.400 53.400 769.050 54.450 ;
        RECT 760.950 46.950 763.050 49.050 ;
        RECT 757.950 43.950 760.050 46.050 ;
        RECT 758.400 22.050 759.450 43.950 ;
        RECT 751.950 19.950 754.050 22.050 ;
        RECT 757.950 19.950 760.050 22.050 ;
        RECT 761.250 20.250 763.050 21.150 ;
        RECT 742.950 17.400 747.450 18.450 ;
        RECT 751.950 17.850 753.750 18.750 ;
        RECT 742.950 16.950 745.050 17.400 ;
        RECT 754.950 16.950 757.050 19.050 ;
        RECT 758.250 17.850 759.750 18.750 ;
        RECT 760.950 16.950 763.050 19.050 ;
        RECT 737.400 16.050 738.450 16.950 ;
        RECT 703.950 13.950 706.050 16.050 ;
        RECT 709.950 13.950 712.050 16.050 ;
        RECT 721.950 13.950 724.050 16.050 ;
        RECT 736.950 13.950 739.050 16.050 ;
        RECT 754.950 14.850 757.050 15.750 ;
        RECT 764.400 10.050 765.450 53.400 ;
        RECT 766.950 52.950 769.050 53.400 ;
        RECT 770.250 53.250 772.050 54.150 ;
        RECT 766.950 50.850 768.750 51.750 ;
        RECT 769.950 49.950 772.050 52.050 ;
        RECT 766.950 22.950 769.050 25.050 ;
        RECT 767.400 16.050 768.450 22.950 ;
        RECT 773.400 22.050 774.450 64.950 ;
        RECT 779.400 55.050 780.450 70.950 ;
        RECT 778.950 52.950 781.050 55.050 ;
        RECT 778.950 50.850 781.050 51.750 ;
        RECT 788.400 28.050 789.450 94.950 ;
        RECT 797.400 94.050 798.450 121.950 ;
        RECT 803.400 115.050 804.450 127.950 ;
        RECT 845.400 127.050 846.450 166.950 ;
        RECT 854.400 166.050 855.450 199.950 ;
        RECT 857.400 169.050 858.450 367.950 ;
        RECT 860.400 235.050 861.450 502.950 ;
        RECT 859.950 232.950 862.050 235.050 ;
        RECT 859.950 202.950 862.050 205.050 ;
        RECT 860.400 199.050 861.450 202.950 ;
        RECT 859.950 196.950 862.050 199.050 ;
        RECT 860.400 196.050 861.450 196.950 ;
        RECT 859.950 193.950 862.050 196.050 ;
        RECT 860.400 172.050 861.450 193.950 ;
        RECT 863.400 184.050 864.450 700.950 ;
        RECT 862.950 181.950 865.050 184.050 ;
        RECT 859.950 169.950 862.050 172.050 ;
        RECT 856.950 166.950 859.050 169.050 ;
        RECT 860.250 167.850 862.050 168.750 ;
        RECT 847.950 163.950 850.050 166.050 ;
        RECT 850.950 163.950 853.050 166.050 ;
        RECT 853.950 163.950 856.050 166.050 ;
        RECT 856.950 164.850 859.050 165.750 ;
        RECT 805.950 124.950 808.050 127.050 ;
        RECT 808.950 125.250 811.050 126.150 ;
        RECT 814.950 125.250 817.050 126.150 ;
        RECT 823.950 125.250 826.050 126.150 ;
        RECT 829.950 124.950 832.050 127.050 ;
        RECT 838.950 124.950 841.050 127.050 ;
        RECT 844.950 124.950 847.050 127.050 ;
        RECT 806.400 124.050 807.450 124.950 ;
        RECT 805.950 121.950 808.050 124.050 ;
        RECT 808.950 121.950 811.050 124.050 ;
        RECT 812.250 122.250 813.750 123.150 ;
        RECT 814.950 121.950 817.050 124.050 ;
        RECT 817.950 121.950 820.050 124.050 ;
        RECT 820.950 122.250 822.750 123.150 ;
        RECT 823.950 121.950 826.050 124.050 ;
        RECT 829.950 122.850 832.050 123.750 ;
        RECT 802.950 112.950 805.050 115.050 ;
        RECT 799.950 100.950 802.050 103.050 ;
        RECT 805.950 100.950 808.050 103.050 ;
        RECT 800.400 97.050 801.450 100.950 ;
        RECT 806.400 97.050 807.450 100.950 ;
        RECT 799.950 94.950 802.050 97.050 ;
        RECT 803.250 95.250 804.750 96.150 ;
        RECT 805.950 94.950 808.050 97.050 ;
        RECT 796.950 91.950 799.050 94.050 ;
        RECT 800.250 92.850 801.750 93.750 ;
        RECT 802.950 91.950 805.050 94.050 ;
        RECT 806.250 92.850 808.050 93.750 ;
        RECT 809.400 91.050 810.450 121.950 ;
        RECT 815.400 121.050 816.450 121.950 ;
        RECT 811.950 118.950 814.050 121.050 ;
        RECT 814.950 118.950 817.050 121.050 ;
        RECT 812.400 117.450 813.450 118.950 ;
        RECT 818.400 117.450 819.450 121.950 ;
        RECT 820.950 118.950 823.050 121.050 ;
        RECT 839.400 120.450 840.450 124.950 ;
        RECT 841.950 122.250 844.050 123.150 ;
        RECT 844.950 122.850 847.050 123.750 ;
        RECT 841.950 120.450 844.050 121.050 ;
        RECT 839.400 119.400 844.050 120.450 ;
        RECT 841.950 118.950 844.050 119.400 ;
        RECT 821.400 118.050 822.450 118.950 ;
        RECT 812.400 116.400 819.450 117.450 ;
        RECT 820.950 115.950 823.050 118.050 ;
        RECT 811.950 103.950 814.050 106.050 ;
        RECT 829.950 103.950 832.050 106.050 ;
        RECT 844.950 103.950 847.050 106.050 ;
        RECT 812.400 97.050 813.450 103.950 ;
        RECT 814.950 100.950 817.050 103.050 ;
        RECT 815.400 100.050 816.450 100.950 ;
        RECT 814.950 97.950 817.050 100.050 ;
        RECT 817.950 97.950 820.050 100.050 ;
        RECT 826.950 97.950 829.050 100.050 ;
        RECT 818.400 97.050 819.450 97.950 ;
        RECT 827.400 97.050 828.450 97.950 ;
        RECT 811.950 94.950 814.050 97.050 ;
        RECT 815.250 95.850 816.750 96.750 ;
        RECT 817.950 94.950 820.050 97.050 ;
        RECT 826.950 94.950 829.050 97.050 ;
        RECT 811.950 92.850 814.050 93.750 ;
        RECT 817.950 92.850 820.050 93.750 ;
        RECT 826.950 92.850 829.050 93.750 ;
        RECT 796.950 89.850 799.050 90.750 ;
        RECT 808.950 88.950 811.050 91.050 ;
        RECT 830.400 90.450 831.450 103.950 ;
        RECT 845.400 97.050 846.450 103.950 ;
        RECT 848.400 100.050 849.450 163.950 ;
        RECT 851.400 130.050 852.450 163.950 ;
        RECT 853.950 160.950 856.050 163.050 ;
        RECT 850.950 127.950 853.050 130.050 ;
        RECT 850.950 124.950 853.050 127.050 ;
        RECT 847.950 97.950 850.050 100.050 ;
        RECT 851.400 97.050 852.450 124.950 ;
        RECT 835.950 94.950 838.050 97.050 ;
        RECT 844.950 94.950 847.050 97.050 ;
        RECT 848.250 95.850 849.750 96.750 ;
        RECT 850.950 94.950 853.050 97.050 ;
        RECT 832.950 92.250 835.050 93.150 ;
        RECT 835.950 92.850 838.050 93.750 ;
        RECT 844.950 92.850 847.050 93.750 ;
        RECT 850.950 92.850 853.050 93.750 ;
        RECT 832.950 90.450 835.050 91.050 ;
        RECT 830.400 89.400 835.050 90.450 ;
        RECT 832.950 88.950 835.050 89.400 ;
        RECT 799.800 65.100 801.900 67.200 ;
        RECT 800.550 61.350 801.750 65.100 ;
        RECT 823.950 64.950 826.050 67.050 ;
        RECT 826.950 64.950 829.050 67.050 ;
        RECT 829.950 64.950 832.050 67.050 ;
        RECT 802.950 62.850 805.050 64.950 ;
        RECT 799.950 59.250 802.050 61.350 ;
        RECT 790.950 56.250 793.050 57.150 ;
        RECT 790.950 52.950 793.050 55.050 ;
        RECT 796.950 52.950 799.050 55.050 ;
        RECT 787.950 25.950 790.050 28.050 ;
        RECT 784.950 23.250 787.050 24.150 ;
        RECT 797.400 22.050 798.450 52.950 ;
        RECT 800.550 45.600 801.750 59.250 ;
        RECT 803.250 45.600 804.450 62.850 ;
        RECT 810.900 62.400 813.000 64.500 ;
        RECT 814.950 62.400 817.050 64.500 ;
        RECT 805.950 59.250 808.050 61.350 ;
        RECT 806.400 45.600 807.600 59.250 ;
        RECT 811.350 53.550 812.550 62.400 ;
        RECT 815.550 56.250 816.750 62.400 ;
        RECT 814.950 54.150 817.050 56.250 ;
        RECT 810.750 51.450 812.850 53.550 ;
        RECT 811.350 45.600 812.550 51.450 ;
        RECT 815.550 45.600 816.750 54.150 ;
        RECT 817.950 50.250 820.050 51.150 ;
        RECT 817.950 46.950 820.050 49.050 ;
        RECT 824.250 46.050 825.450 64.950 ;
        RECT 827.250 60.750 828.450 64.950 ;
        RECT 826.950 58.650 829.050 60.750 ;
        RECT 827.250 46.050 828.450 58.650 ;
        RECT 830.250 46.050 831.450 64.950 ;
        RECT 841.950 58.950 844.050 61.050 ;
        RECT 842.400 58.050 843.450 58.950 ;
        RECT 854.400 58.050 855.450 160.950 ;
        RECT 835.950 56.250 838.050 57.150 ;
        RECT 841.950 55.950 844.050 58.050 ;
        RECT 853.950 55.950 856.050 58.050 ;
        RECT 841.950 53.850 844.050 54.750 ;
        RECT 799.950 43.500 802.050 45.600 ;
        RECT 802.950 43.500 805.050 45.600 ;
        RECT 805.950 43.500 808.050 45.600 ;
        RECT 810.750 43.500 812.850 45.600 ;
        RECT 814.950 43.500 817.050 45.600 ;
        RECT 823.950 43.950 826.050 46.050 ;
        RECT 826.950 43.950 829.050 46.050 ;
        RECT 829.950 43.950 832.050 46.050 ;
        RECT 805.950 29.400 808.050 31.500 ;
        RECT 808.950 29.400 811.050 31.500 ;
        RECT 811.950 29.400 814.050 31.500 ;
        RECT 816.750 29.400 818.850 31.500 ;
        RECT 820.950 29.400 823.050 31.500 ;
        RECT 769.950 20.250 771.750 21.150 ;
        RECT 772.950 19.950 775.050 22.050 ;
        RECT 776.250 20.250 778.050 21.150 ;
        RECT 784.950 19.950 787.050 22.050 ;
        RECT 796.950 19.950 799.050 22.050 ;
        RECT 769.950 16.950 772.050 19.050 ;
        RECT 773.250 17.850 774.750 18.750 ;
        RECT 775.950 16.950 778.050 19.050 ;
        RECT 776.400 16.050 777.450 16.950 ;
        RECT 766.950 13.950 769.050 16.050 ;
        RECT 775.950 13.950 778.050 16.050 ;
        RECT 785.400 10.050 786.450 19.950 ;
        RECT 796.950 17.850 799.050 18.750 ;
        RECT 806.550 15.750 807.750 29.400 ;
        RECT 805.950 13.650 808.050 15.750 ;
        RECT 610.800 7.800 612.900 9.900 ;
        RECT 634.950 7.950 637.050 10.050 ;
        RECT 637.950 7.950 640.050 10.050 ;
        RECT 640.950 7.950 643.050 10.050 ;
        RECT 763.950 7.950 766.050 10.050 ;
        RECT 784.950 7.950 787.050 10.050 ;
        RECT 806.550 9.900 807.750 13.650 ;
        RECT 809.250 12.150 810.450 29.400 ;
        RECT 812.400 15.750 813.600 29.400 ;
        RECT 817.350 23.550 818.550 29.400 ;
        RECT 816.750 21.450 818.850 23.550 ;
        RECT 811.950 13.650 814.050 15.750 ;
        RECT 817.350 12.600 818.550 21.450 ;
        RECT 821.550 20.850 822.750 29.400 ;
        RECT 829.950 28.950 832.050 31.050 ;
        RECT 832.950 28.950 835.050 31.050 ;
        RECT 835.950 28.950 838.050 31.050 ;
        RECT 823.950 25.950 826.050 28.050 ;
        RECT 823.950 23.850 826.050 24.750 ;
        RECT 820.950 18.750 823.050 20.850 ;
        RECT 821.550 12.600 822.750 18.750 ;
        RECT 808.950 10.050 811.050 12.150 ;
        RECT 816.900 10.500 819.000 12.600 ;
        RECT 820.950 10.500 823.050 12.600 ;
        RECT 830.250 10.050 831.450 28.950 ;
        RECT 833.250 16.350 834.450 28.950 ;
        RECT 832.950 14.250 835.050 16.350 ;
        RECT 833.250 10.050 834.450 14.250 ;
        RECT 836.250 10.050 837.450 28.950 ;
        RECT 847.950 20.250 850.050 21.150 ;
        RECT 854.400 19.050 855.450 55.950 ;
        RECT 841.950 17.850 844.050 18.750 ;
        RECT 847.950 16.950 850.050 19.050 ;
        RECT 853.950 16.950 856.050 19.050 ;
        RECT 805.800 7.800 807.900 9.900 ;
        RECT 829.950 7.950 832.050 10.050 ;
        RECT 832.950 7.950 835.050 10.050 ;
        RECT 835.950 7.950 838.050 10.050 ;
        RECT 337.950 4.950 340.050 7.050 ;
        RECT 523.950 4.950 526.050 7.050 ;
      LAYER metal3 ;
        RECT 181.950 822.600 184.050 823.050 ;
        RECT 241.950 822.600 244.050 823.050 ;
        RECT 274.950 822.600 277.050 823.050 ;
        RECT 181.950 821.400 277.050 822.600 ;
        RECT 181.950 820.950 184.050 821.400 ;
        RECT 241.950 820.950 244.050 821.400 ;
        RECT 274.950 820.950 277.050 821.400 ;
        RECT 442.950 822.600 445.050 823.050 ;
        RECT 451.950 822.600 454.050 823.050 ;
        RECT 502.950 822.600 505.050 823.050 ;
        RECT 442.950 821.400 505.050 822.600 ;
        RECT 442.950 820.950 445.050 821.400 ;
        RECT 451.950 820.950 454.050 821.400 ;
        RECT 502.950 820.950 505.050 821.400 ;
        RECT 508.950 822.600 511.050 823.050 ;
        RECT 523.950 822.600 526.050 823.050 ;
        RECT 508.950 821.400 526.050 822.600 ;
        RECT 508.950 820.950 511.050 821.400 ;
        RECT 523.950 820.950 526.050 821.400 ;
        RECT 787.950 822.600 790.050 823.050 ;
        RECT 796.950 822.600 799.050 823.050 ;
        RECT 787.950 821.400 799.050 822.600 ;
        RECT 787.950 820.950 790.050 821.400 ;
        RECT 796.950 820.950 799.050 821.400 ;
        RECT 10.950 819.600 13.050 820.050 ;
        RECT 22.950 819.600 25.050 820.050 ;
        RECT 10.950 818.400 25.050 819.600 ;
        RECT 10.950 817.950 13.050 818.400 ;
        RECT 22.950 817.950 25.050 818.400 ;
        RECT 28.950 819.600 31.050 820.050 ;
        RECT 37.950 819.600 40.050 820.050 ;
        RECT 28.950 818.400 40.050 819.600 ;
        RECT 28.950 817.950 31.050 818.400 ;
        RECT 37.950 817.950 40.050 818.400 ;
        RECT 40.950 819.600 43.050 820.050 ;
        RECT 76.950 819.600 79.050 820.050 ;
        RECT 40.950 818.400 79.050 819.600 ;
        RECT 40.950 817.950 43.050 818.400 ;
        RECT 76.950 817.950 79.050 818.400 ;
        RECT 118.950 819.600 121.050 820.050 ;
        RECT 130.950 819.600 133.050 820.050 ;
        RECT 136.950 819.600 139.050 820.050 ;
        RECT 118.950 818.400 139.050 819.600 ;
        RECT 118.950 817.950 121.050 818.400 ;
        RECT 130.950 817.950 133.050 818.400 ;
        RECT 136.950 817.950 139.050 818.400 ;
        RECT 187.950 819.600 190.050 820.050 ;
        RECT 256.950 819.600 259.050 820.050 ;
        RECT 187.950 818.400 259.050 819.600 ;
        RECT 187.950 817.950 190.050 818.400 ;
        RECT 256.950 817.950 259.050 818.400 ;
        RECT 259.950 819.600 262.050 820.050 ;
        RECT 295.950 819.600 298.050 820.050 ;
        RECT 259.950 818.400 298.050 819.600 ;
        RECT 259.950 817.950 262.050 818.400 ;
        RECT 295.950 817.950 298.050 818.400 ;
        RECT 340.950 819.600 343.050 820.050 ;
        RECT 421.950 819.600 424.050 820.050 ;
        RECT 445.950 819.600 448.050 820.050 ;
        RECT 340.950 818.400 448.050 819.600 ;
        RECT 340.950 817.950 343.050 818.400 ;
        RECT 421.950 817.950 424.050 818.400 ;
        RECT 445.950 817.950 448.050 818.400 ;
        RECT 475.950 819.600 478.050 820.050 ;
        RECT 484.950 819.600 487.050 820.050 ;
        RECT 475.950 818.400 487.050 819.600 ;
        RECT 475.950 817.950 478.050 818.400 ;
        RECT 484.950 817.950 487.050 818.400 ;
        RECT 511.950 819.600 514.050 820.050 ;
        RECT 538.950 819.600 541.050 820.050 ;
        RECT 559.950 819.600 562.050 820.050 ;
        RECT 511.950 818.400 562.050 819.600 ;
        RECT 511.950 817.950 514.050 818.400 ;
        RECT 538.950 817.950 541.050 818.400 ;
        RECT 559.950 817.950 562.050 818.400 ;
        RECT 691.950 819.600 694.050 820.050 ;
        RECT 754.950 819.600 757.050 820.050 ;
        RECT 790.950 819.600 793.050 820.050 ;
        RECT 811.950 819.600 814.050 820.050 ;
        RECT 691.950 818.400 789.600 819.600 ;
        RECT 691.950 817.950 694.050 818.400 ;
        RECT 754.950 817.950 757.050 818.400 ;
        RECT 7.950 816.600 10.050 817.050 ;
        RECT 139.950 816.600 142.050 817.050 ;
        RECT 7.950 815.400 142.050 816.600 ;
        RECT 7.950 814.950 10.050 815.400 ;
        RECT 139.950 814.950 142.050 815.400 ;
        RECT 193.950 816.600 196.050 817.050 ;
        RECT 199.950 816.600 202.050 817.050 ;
        RECT 193.950 815.400 202.050 816.600 ;
        RECT 193.950 814.950 196.050 815.400 ;
        RECT 199.950 814.950 202.050 815.400 ;
        RECT 214.950 814.950 217.050 817.050 ;
        RECT 223.950 816.600 226.050 817.050 ;
        RECT 235.950 816.600 238.050 817.050 ;
        RECT 223.950 815.400 238.050 816.600 ;
        RECT 223.950 814.950 226.050 815.400 ;
        RECT 235.950 814.950 238.050 815.400 ;
        RECT 328.950 816.600 331.050 817.050 ;
        RECT 346.950 816.600 349.050 817.050 ;
        RECT 370.950 816.600 373.050 817.050 ;
        RECT 328.950 815.400 373.050 816.600 ;
        RECT 328.950 814.950 331.050 815.400 ;
        RECT 346.950 814.950 349.050 815.400 ;
        RECT 370.950 814.950 373.050 815.400 ;
        RECT 484.950 816.600 487.050 817.050 ;
        RECT 541.950 816.600 544.050 817.050 ;
        RECT 484.950 815.400 544.050 816.600 ;
        RECT 484.950 814.950 487.050 815.400 ;
        RECT 541.950 814.950 544.050 815.400 ;
        RECT 553.950 814.950 556.050 817.050 ;
        RECT 601.950 816.600 604.050 817.050 ;
        RECT 613.950 816.600 616.050 817.050 ;
        RECT 601.950 815.400 616.050 816.600 ;
        RECT 601.950 814.950 604.050 815.400 ;
        RECT 613.950 814.950 616.050 815.400 ;
        RECT 619.950 816.600 622.050 817.050 ;
        RECT 637.950 816.600 640.050 817.050 ;
        RECT 619.950 815.400 640.050 816.600 ;
        RECT 619.950 814.950 622.050 815.400 ;
        RECT 637.950 814.950 640.050 815.400 ;
        RECT 643.950 816.600 646.050 817.050 ;
        RECT 652.950 816.600 655.050 817.050 ;
        RECT 643.950 815.400 655.050 816.600 ;
        RECT 643.950 814.950 646.050 815.400 ;
        RECT 652.950 814.950 655.050 815.400 ;
        RECT 676.950 816.600 679.050 817.050 ;
        RECT 712.950 816.600 715.050 817.050 ;
        RECT 733.950 816.600 736.050 817.050 ;
        RECT 676.950 815.400 736.050 816.600 ;
        RECT 676.950 814.950 679.050 815.400 ;
        RECT 712.950 814.950 715.050 815.400 ;
        RECT 733.950 814.950 736.050 815.400 ;
        RECT 742.950 816.600 745.050 817.050 ;
        RECT 775.950 816.600 778.050 817.050 ;
        RECT 742.950 815.400 778.050 816.600 ;
        RECT 742.950 814.950 745.050 815.400 ;
        RECT 775.950 814.950 778.050 815.400 ;
        RECT 778.950 816.600 781.050 817.050 ;
        RECT 784.950 816.600 787.050 817.050 ;
        RECT 778.950 815.400 787.050 816.600 ;
        RECT 788.400 816.600 789.600 818.400 ;
        RECT 790.950 818.400 814.050 819.600 ;
        RECT 790.950 817.950 793.050 818.400 ;
        RECT 811.950 817.950 814.050 818.400 ;
        RECT 820.950 819.600 823.050 820.050 ;
        RECT 829.950 819.600 832.050 820.050 ;
        RECT 838.950 819.600 841.050 820.050 ;
        RECT 820.950 818.400 841.050 819.600 ;
        RECT 820.950 817.950 823.050 818.400 ;
        RECT 829.950 817.950 832.050 818.400 ;
        RECT 838.950 817.950 841.050 818.400 ;
        RECT 793.950 816.600 796.050 817.050 ;
        RECT 788.400 815.400 796.050 816.600 ;
        RECT 778.950 814.950 781.050 815.400 ;
        RECT 784.950 814.950 787.050 815.400 ;
        RECT 793.950 814.950 796.050 815.400 ;
        RECT 802.950 814.950 805.050 817.050 ;
        RECT 805.950 816.600 808.050 817.050 ;
        RECT 817.950 816.600 820.050 817.050 ;
        RECT 805.950 815.400 820.050 816.600 ;
        RECT 805.950 814.950 808.050 815.400 ;
        RECT 817.950 814.950 820.050 815.400 ;
        RECT 103.950 813.600 106.050 814.050 ;
        RECT 121.950 813.600 124.050 814.050 ;
        RECT 103.950 812.400 124.050 813.600 ;
        RECT 103.950 811.950 106.050 812.400 ;
        RECT 121.950 811.950 124.050 812.400 ;
        RECT 127.950 813.600 130.050 814.050 ;
        RECT 140.400 813.600 141.600 814.950 ;
        RECT 127.950 812.400 141.600 813.600 ;
        RECT 175.950 813.600 178.050 814.050 ;
        RECT 215.400 813.600 216.600 814.950 ;
        RECT 244.950 813.600 247.050 814.050 ;
        RECT 175.950 812.400 186.600 813.600 ;
        RECT 127.950 811.950 130.050 812.400 ;
        RECT 175.950 811.950 178.050 812.400 ;
        RECT 185.400 811.050 186.600 812.400 ;
        RECT 197.400 812.400 247.050 813.600 ;
        RECT 197.400 811.050 198.600 812.400 ;
        RECT 244.950 811.950 247.050 812.400 ;
        RECT 274.950 813.600 277.050 814.050 ;
        RECT 334.950 813.600 337.050 814.050 ;
        RECT 274.950 812.400 337.050 813.600 ;
        RECT 274.950 811.950 277.050 812.400 ;
        RECT 334.950 811.950 337.050 812.400 ;
        RECT 415.950 813.600 418.050 814.050 ;
        RECT 436.950 813.600 439.050 814.050 ;
        RECT 415.950 812.400 439.050 813.600 ;
        RECT 415.950 811.950 418.050 812.400 ;
        RECT 436.950 811.950 439.050 812.400 ;
        RECT 451.950 813.600 454.050 814.050 ;
        RECT 490.950 813.600 493.050 814.050 ;
        RECT 451.950 812.400 493.050 813.600 ;
        RECT 451.950 811.950 454.050 812.400 ;
        RECT 490.950 811.950 493.050 812.400 ;
        RECT 520.950 813.600 523.050 814.050 ;
        RECT 554.400 813.600 555.600 814.950 ;
        RECT 574.950 813.600 577.050 814.050 ;
        RECT 586.950 813.600 589.050 814.050 ;
        RECT 520.950 812.400 577.050 813.600 ;
        RECT 520.950 811.950 523.050 812.400 ;
        RECT 574.950 811.950 577.050 812.400 ;
        RECT 578.400 812.400 589.050 813.600 ;
        RECT 578.400 811.050 579.600 812.400 ;
        RECT 586.950 811.950 589.050 812.400 ;
        RECT 610.950 811.950 613.050 814.050 ;
        RECT 616.950 813.600 619.050 814.050 ;
        RECT 631.950 813.600 634.050 814.050 ;
        RECT 646.950 813.600 649.050 814.050 ;
        RECT 616.950 812.400 649.050 813.600 ;
        RECT 616.950 811.950 619.050 812.400 ;
        RECT 631.950 811.950 634.050 812.400 ;
        RECT 646.950 811.950 649.050 812.400 ;
        RECT 658.950 813.600 661.050 814.050 ;
        RECT 664.950 813.600 667.050 814.050 ;
        RECT 658.950 812.400 667.050 813.600 ;
        RECT 658.950 811.950 661.050 812.400 ;
        RECT 664.950 811.950 667.050 812.400 ;
        RECT 667.950 813.600 670.050 814.050 ;
        RECT 673.950 813.600 676.050 814.050 ;
        RECT 667.950 812.400 676.050 813.600 ;
        RECT 667.950 811.950 670.050 812.400 ;
        RECT 673.950 811.950 676.050 812.400 ;
        RECT 697.950 813.600 700.050 814.050 ;
        RECT 703.950 813.600 706.050 814.050 ;
        RECT 697.950 812.400 706.050 813.600 ;
        RECT 697.950 811.950 700.050 812.400 ;
        RECT 703.950 811.950 706.050 812.400 ;
        RECT 718.950 813.600 721.050 814.050 ;
        RECT 730.950 813.600 733.050 814.050 ;
        RECT 718.950 812.400 733.050 813.600 ;
        RECT 743.400 813.600 744.600 814.950 ;
        RECT 751.950 813.600 754.050 814.050 ;
        RECT 743.400 812.400 754.050 813.600 ;
        RECT 718.950 811.950 721.050 812.400 ;
        RECT 730.950 811.950 733.050 812.400 ;
        RECT 751.950 811.950 754.050 812.400 ;
        RECT 769.950 813.600 772.050 814.050 ;
        RECT 781.950 813.600 784.050 814.050 ;
        RECT 790.950 813.600 793.050 814.050 ;
        RECT 769.950 812.400 793.050 813.600 ;
        RECT 803.400 813.600 804.600 814.950 ;
        RECT 811.950 813.600 814.050 814.050 ;
        RECT 826.950 813.600 829.050 814.050 ;
        RECT 803.400 812.400 829.050 813.600 ;
        RECT 769.950 811.950 772.050 812.400 ;
        RECT 781.950 811.950 784.050 812.400 ;
        RECT 790.950 811.950 793.050 812.400 ;
        RECT 811.950 811.950 814.050 812.400 ;
        RECT 826.950 811.950 829.050 812.400 ;
        RECT 22.950 810.600 25.050 811.050 ;
        RECT 31.950 810.600 34.050 811.050 ;
        RECT 22.950 809.400 34.050 810.600 ;
        RECT 22.950 808.950 25.050 809.400 ;
        RECT 31.950 808.950 34.050 809.400 ;
        RECT 124.950 810.600 127.050 811.050 ;
        RECT 145.950 810.600 148.050 811.050 ;
        RECT 124.950 809.400 148.050 810.600 ;
        RECT 124.950 808.950 127.050 809.400 ;
        RECT 145.950 808.950 148.050 809.400 ;
        RECT 154.950 810.600 157.050 811.050 ;
        RECT 163.950 810.600 166.050 811.050 ;
        RECT 172.950 810.600 175.050 811.050 ;
        RECT 154.950 809.400 175.050 810.600 ;
        RECT 154.950 808.950 157.050 809.400 ;
        RECT 163.950 808.950 166.050 809.400 ;
        RECT 172.950 808.950 175.050 809.400 ;
        RECT 184.950 808.950 187.050 811.050 ;
        RECT 196.950 808.950 199.050 811.050 ;
        RECT 202.950 810.600 205.050 811.050 ;
        RECT 217.950 810.600 220.050 811.050 ;
        RECT 202.950 809.400 220.050 810.600 ;
        RECT 202.950 808.950 205.050 809.400 ;
        RECT 217.950 808.950 220.050 809.400 ;
        RECT 295.950 810.600 298.050 811.050 ;
        RECT 325.950 810.600 328.050 811.050 ;
        RECT 391.950 810.600 394.050 811.050 ;
        RECT 295.950 809.400 394.050 810.600 ;
        RECT 295.950 808.950 298.050 809.400 ;
        RECT 325.950 808.950 328.050 809.400 ;
        RECT 391.950 808.950 394.050 809.400 ;
        RECT 424.950 810.600 427.050 811.050 ;
        RECT 433.950 810.600 436.050 811.050 ;
        RECT 448.950 810.600 451.050 811.050 ;
        RECT 424.950 809.400 451.050 810.600 ;
        RECT 424.950 808.950 427.050 809.400 ;
        RECT 433.950 808.950 436.050 809.400 ;
        RECT 448.950 808.950 451.050 809.400 ;
        RECT 460.950 810.600 463.050 811.050 ;
        RECT 472.950 810.600 475.050 811.050 ;
        RECT 460.950 809.400 475.050 810.600 ;
        RECT 460.950 808.950 463.050 809.400 ;
        RECT 472.950 808.950 475.050 809.400 ;
        RECT 505.950 810.600 508.050 811.050 ;
        RECT 517.950 810.600 520.050 811.050 ;
        RECT 505.950 809.400 520.050 810.600 ;
        RECT 505.950 808.950 508.050 809.400 ;
        RECT 517.950 808.950 520.050 809.400 ;
        RECT 544.950 810.600 547.050 811.050 ;
        RECT 577.950 810.600 580.050 811.050 ;
        RECT 544.950 809.400 580.050 810.600 ;
        RECT 611.400 810.600 612.600 811.950 ;
        RECT 628.950 810.600 631.050 811.050 ;
        RECT 611.400 809.400 631.050 810.600 ;
        RECT 544.950 808.950 547.050 809.400 ;
        RECT 577.950 808.950 580.050 809.400 ;
        RECT 628.950 808.950 631.050 809.400 ;
        RECT 634.950 808.950 637.050 811.050 ;
        RECT 640.950 810.600 643.050 811.050 ;
        RECT 706.950 810.600 709.050 811.050 ;
        RECT 748.950 810.600 751.050 811.050 ;
        RECT 841.950 810.600 844.050 811.050 ;
        RECT 640.950 809.400 844.050 810.600 ;
        RECT 640.950 808.950 643.050 809.400 ;
        RECT 706.950 808.950 709.050 809.400 ;
        RECT 748.950 808.950 751.050 809.400 ;
        RECT 841.950 808.950 844.050 809.400 ;
        RECT 7.950 807.600 10.050 808.050 ;
        RECT 13.950 807.600 16.050 808.050 ;
        RECT 151.950 807.600 154.050 808.050 ;
        RECT 7.950 806.400 154.050 807.600 ;
        RECT 7.950 805.950 10.050 806.400 ;
        RECT 13.950 805.950 16.050 806.400 ;
        RECT 151.950 805.950 154.050 806.400 ;
        RECT 208.950 807.600 211.050 808.050 ;
        RECT 265.950 807.600 268.050 808.050 ;
        RECT 208.950 806.400 268.050 807.600 ;
        RECT 208.950 805.950 211.050 806.400 ;
        RECT 265.950 805.950 268.050 806.400 ;
        RECT 271.950 807.600 274.050 808.050 ;
        RECT 349.950 807.600 352.050 808.050 ;
        RECT 271.950 806.400 352.050 807.600 ;
        RECT 271.950 805.950 274.050 806.400 ;
        RECT 349.950 805.950 352.050 806.400 ;
        RECT 445.950 807.600 448.050 808.050 ;
        RECT 478.950 807.600 481.050 808.050 ;
        RECT 493.950 807.600 496.050 808.050 ;
        RECT 445.950 806.400 496.050 807.600 ;
        RECT 445.950 805.950 448.050 806.400 ;
        RECT 478.950 805.950 481.050 806.400 ;
        RECT 493.950 805.950 496.050 806.400 ;
        RECT 526.950 807.600 529.050 808.050 ;
        RECT 541.950 807.600 544.050 808.050 ;
        RECT 565.950 807.600 568.050 808.050 ;
        RECT 598.950 807.600 601.050 808.050 ;
        RECT 526.950 806.400 601.050 807.600 ;
        RECT 526.950 805.950 529.050 806.400 ;
        RECT 541.950 805.950 544.050 806.400 ;
        RECT 565.950 805.950 568.050 806.400 ;
        RECT 598.950 805.950 601.050 806.400 ;
        RECT 631.950 807.600 634.050 808.050 ;
        RECT 635.400 807.600 636.600 808.950 ;
        RECT 631.950 806.400 636.600 807.600 ;
        RECT 646.950 807.600 649.050 808.050 ;
        RECT 670.950 807.600 673.050 808.050 ;
        RECT 646.950 806.400 673.050 807.600 ;
        RECT 631.950 805.950 634.050 806.400 ;
        RECT 646.950 805.950 649.050 806.400 ;
        RECT 670.950 805.950 673.050 806.400 ;
        RECT 736.950 807.600 739.050 808.050 ;
        RECT 772.950 807.600 775.050 808.050 ;
        RECT 736.950 806.400 775.050 807.600 ;
        RECT 736.950 805.950 739.050 806.400 ;
        RECT 772.950 805.950 775.050 806.400 ;
        RECT 787.950 807.600 790.050 808.050 ;
        RECT 820.950 807.600 823.050 808.050 ;
        RECT 787.950 806.400 823.050 807.600 ;
        RECT 787.950 805.950 790.050 806.400 ;
        RECT 820.950 805.950 823.050 806.400 ;
        RECT 25.950 804.600 28.050 805.050 ;
        RECT 202.950 804.600 205.050 805.050 ;
        RECT 25.950 803.400 205.050 804.600 ;
        RECT 25.950 802.950 28.050 803.400 ;
        RECT 202.950 802.950 205.050 803.400 ;
        RECT 454.950 804.600 457.050 805.050 ;
        RECT 463.950 804.600 466.050 805.050 ;
        RECT 454.950 803.400 466.050 804.600 ;
        RECT 454.950 802.950 457.050 803.400 ;
        RECT 463.950 802.950 466.050 803.400 ;
        RECT 493.950 804.600 496.050 805.050 ;
        RECT 532.950 804.600 535.050 805.050 ;
        RECT 493.950 803.400 535.050 804.600 ;
        RECT 493.950 802.950 496.050 803.400 ;
        RECT 532.950 802.950 535.050 803.400 ;
        RECT 550.950 804.600 553.050 805.050 ;
        RECT 556.950 804.600 559.050 805.050 ;
        RECT 550.950 803.400 559.050 804.600 ;
        RECT 550.950 802.950 553.050 803.400 ;
        RECT 556.950 802.950 559.050 803.400 ;
        RECT 598.950 804.600 601.050 805.050 ;
        RECT 661.950 804.600 664.050 805.050 ;
        RECT 598.950 803.400 664.050 804.600 ;
        RECT 598.950 802.950 601.050 803.400 ;
        RECT 661.950 802.950 664.050 803.400 ;
        RECT 664.950 804.600 667.050 805.050 ;
        RECT 688.950 804.600 691.050 805.050 ;
        RECT 664.950 803.400 691.050 804.600 ;
        RECT 664.950 802.950 667.050 803.400 ;
        RECT 688.950 802.950 691.050 803.400 ;
        RECT 628.950 801.600 631.050 802.050 ;
        RECT 667.950 801.600 670.050 802.050 ;
        RECT 721.950 801.600 724.050 802.050 ;
        RECT 763.950 801.600 766.050 802.050 ;
        RECT 766.950 801.600 769.050 802.050 ;
        RECT 628.950 800.400 769.050 801.600 ;
        RECT 628.950 799.950 631.050 800.400 ;
        RECT 667.950 799.950 670.050 800.400 ;
        RECT 721.950 799.950 724.050 800.400 ;
        RECT 763.950 799.950 766.050 800.400 ;
        RECT 766.950 799.950 769.050 800.400 ;
        RECT 52.950 798.600 55.050 799.050 ;
        RECT 67.950 798.600 70.050 799.050 ;
        RECT 52.950 797.400 70.050 798.600 ;
        RECT 52.950 796.950 55.050 797.400 ;
        RECT 67.950 796.950 70.050 797.400 ;
        RECT 169.950 789.600 172.050 790.050 ;
        RECT 226.950 789.600 229.050 790.050 ;
        RECT 235.950 789.600 238.050 790.050 ;
        RECT 277.950 789.600 280.050 790.050 ;
        RECT 340.950 789.600 343.050 790.050 ;
        RECT 169.950 788.400 343.050 789.600 ;
        RECT 169.950 787.950 172.050 788.400 ;
        RECT 226.950 787.950 229.050 788.400 ;
        RECT 235.950 787.950 238.050 788.400 ;
        RECT 277.950 787.950 280.050 788.400 ;
        RECT 340.950 787.950 343.050 788.400 ;
        RECT 346.950 783.600 349.050 784.050 ;
        RECT 460.950 783.600 463.050 784.050 ;
        RECT 514.950 783.600 517.050 784.050 ;
        RECT 346.950 782.400 517.050 783.600 ;
        RECT 346.950 781.950 349.050 782.400 ;
        RECT 460.950 781.950 463.050 782.400 ;
        RECT 514.950 781.950 517.050 782.400 ;
        RECT 643.950 783.600 646.050 784.050 ;
        RECT 757.950 783.600 760.050 784.050 ;
        RECT 778.950 783.600 781.050 784.050 ;
        RECT 829.950 783.600 832.050 784.050 ;
        RECT 835.950 783.600 838.050 784.050 ;
        RECT 643.950 782.400 838.050 783.600 ;
        RECT 643.950 781.950 646.050 782.400 ;
        RECT 757.950 781.950 760.050 782.400 ;
        RECT 778.950 781.950 781.050 782.400 ;
        RECT 829.950 781.950 832.050 782.400 ;
        RECT 835.950 781.950 838.050 782.400 ;
        RECT 412.950 780.600 415.050 781.050 ;
        RECT 424.950 780.600 427.050 781.050 ;
        RECT 451.950 780.600 454.050 781.050 ;
        RECT 412.950 779.400 454.050 780.600 ;
        RECT 412.950 778.950 415.050 779.400 ;
        RECT 424.950 778.950 427.050 779.400 ;
        RECT 451.950 778.950 454.050 779.400 ;
        RECT 508.950 780.600 511.050 781.050 ;
        RECT 574.950 780.600 577.050 781.050 ;
        RECT 601.950 780.600 604.050 781.050 ;
        RECT 508.950 779.400 528.600 780.600 ;
        RECT 508.950 778.950 511.050 779.400 ;
        RECT 28.950 777.600 31.050 778.050 ;
        RECT 40.950 777.600 43.050 778.050 ;
        RECT 28.950 776.400 43.050 777.600 ;
        RECT 28.950 775.950 31.050 776.400 ;
        RECT 40.950 775.950 43.050 776.400 ;
        RECT 46.950 775.950 49.050 778.050 ;
        RECT 139.950 777.600 142.050 778.050 ;
        RECT 145.950 777.600 148.050 778.050 ;
        RECT 139.950 776.400 148.050 777.600 ;
        RECT 139.950 775.950 142.050 776.400 ;
        RECT 145.950 775.950 148.050 776.400 ;
        RECT 148.950 777.600 151.050 778.050 ;
        RECT 160.950 777.600 163.050 778.050 ;
        RECT 148.950 776.400 163.050 777.600 ;
        RECT 148.950 775.950 151.050 776.400 ;
        RECT 160.950 775.950 163.050 776.400 ;
        RECT 214.950 777.600 217.050 778.050 ;
        RECT 223.950 777.600 226.050 778.050 ;
        RECT 271.950 777.600 274.050 778.050 ;
        RECT 214.950 776.400 274.050 777.600 ;
        RECT 214.950 775.950 217.050 776.400 ;
        RECT 223.950 775.950 226.050 776.400 ;
        RECT 271.950 775.950 274.050 776.400 ;
        RECT 388.950 777.600 391.050 778.050 ;
        RECT 403.950 777.600 406.050 778.050 ;
        RECT 388.950 776.400 406.050 777.600 ;
        RECT 388.950 775.950 391.050 776.400 ;
        RECT 403.950 775.950 406.050 776.400 ;
        RECT 451.950 777.600 454.050 778.050 ;
        RECT 508.950 777.600 511.050 778.050 ;
        RECT 520.950 777.600 523.050 778.050 ;
        RECT 451.950 776.400 523.050 777.600 ;
        RECT 451.950 775.950 454.050 776.400 ;
        RECT 508.950 775.950 511.050 776.400 ;
        RECT 520.950 775.950 523.050 776.400 ;
        RECT 10.950 774.600 13.050 775.050 ;
        RECT 47.400 774.600 48.600 775.950 ;
        RECT 10.950 773.400 48.600 774.600 ;
        RECT 130.950 774.600 133.050 775.050 ;
        RECT 133.950 774.600 136.050 775.050 ;
        RECT 151.950 774.600 154.050 775.050 ;
        RECT 130.950 773.400 154.050 774.600 ;
        RECT 10.950 772.950 13.050 773.400 ;
        RECT 130.950 772.950 133.050 773.400 ;
        RECT 133.950 772.950 136.050 773.400 ;
        RECT 151.950 772.950 154.050 773.400 ;
        RECT 157.950 774.600 160.050 775.050 ;
        RECT 163.950 774.600 166.050 775.050 ;
        RECT 157.950 773.400 166.050 774.600 ;
        RECT 157.950 772.950 160.050 773.400 ;
        RECT 163.950 772.950 166.050 773.400 ;
        RECT 172.950 774.600 175.050 775.050 ;
        RECT 187.950 774.600 190.050 775.050 ;
        RECT 172.950 773.400 190.050 774.600 ;
        RECT 172.950 772.950 175.050 773.400 ;
        RECT 187.950 772.950 190.050 773.400 ;
        RECT 193.950 774.600 196.050 775.050 ;
        RECT 211.950 774.600 214.050 775.050 ;
        RECT 193.950 773.400 214.050 774.600 ;
        RECT 193.950 772.950 196.050 773.400 ;
        RECT 211.950 772.950 214.050 773.400 ;
        RECT 406.950 774.600 409.050 775.050 ;
        RECT 415.950 774.600 418.050 775.050 ;
        RECT 406.950 773.400 418.050 774.600 ;
        RECT 406.950 772.950 409.050 773.400 ;
        RECT 415.950 772.950 418.050 773.400 ;
        RECT 484.950 774.600 487.050 775.050 ;
        RECT 502.950 774.600 505.050 775.050 ;
        RECT 523.950 774.600 526.050 775.050 ;
        RECT 484.950 773.400 505.050 774.600 ;
        RECT 484.950 772.950 487.050 773.400 ;
        RECT 502.950 772.950 505.050 773.400 ;
        RECT 518.400 773.400 526.050 774.600 ;
        RECT 49.950 771.600 52.050 772.050 ;
        RECT 58.950 771.600 61.050 772.050 ;
        RECT 49.950 770.400 61.050 771.600 ;
        RECT 49.950 769.950 52.050 770.400 ;
        RECT 58.950 769.950 61.050 770.400 ;
        RECT 139.950 771.600 142.050 772.050 ;
        RECT 154.950 771.600 157.050 772.050 ;
        RECT 139.950 770.400 157.050 771.600 ;
        RECT 139.950 769.950 142.050 770.400 ;
        RECT 154.950 769.950 157.050 770.400 ;
        RECT 190.950 771.600 193.050 772.050 ;
        RECT 199.950 771.600 202.050 772.050 ;
        RECT 190.950 770.400 202.050 771.600 ;
        RECT 190.950 769.950 193.050 770.400 ;
        RECT 199.950 769.950 202.050 770.400 ;
        RECT 265.950 771.600 268.050 772.050 ;
        RECT 295.950 771.600 298.050 772.050 ;
        RECT 265.950 770.400 298.050 771.600 ;
        RECT 265.950 769.950 268.050 770.400 ;
        RECT 295.950 769.950 298.050 770.400 ;
        RECT 409.950 771.600 412.050 772.050 ;
        RECT 430.950 771.600 433.050 772.050 ;
        RECT 457.950 771.600 460.050 772.050 ;
        RECT 463.950 771.600 466.050 772.050 ;
        RECT 409.950 770.400 466.050 771.600 ;
        RECT 409.950 769.950 412.050 770.400 ;
        RECT 430.950 769.950 433.050 770.400 ;
        RECT 457.950 769.950 460.050 770.400 ;
        RECT 463.950 769.950 466.050 770.400 ;
        RECT 505.950 771.600 508.050 772.050 ;
        RECT 518.400 771.600 519.600 773.400 ;
        RECT 523.950 772.950 526.050 773.400 ;
        RECT 505.950 770.400 519.600 771.600 ;
        RECT 520.950 771.600 523.050 772.050 ;
        RECT 527.400 771.600 528.600 779.400 ;
        RECT 574.950 779.400 604.050 780.600 ;
        RECT 574.950 778.950 577.050 779.400 ;
        RECT 601.950 778.950 604.050 779.400 ;
        RECT 676.950 780.600 679.050 781.050 ;
        RECT 730.950 780.600 733.050 781.050 ;
        RECT 676.950 779.400 733.050 780.600 ;
        RECT 676.950 778.950 679.050 779.400 ;
        RECT 730.950 778.950 733.050 779.400 ;
        RECT 790.950 780.600 793.050 781.050 ;
        RECT 802.950 780.600 805.050 781.050 ;
        RECT 790.950 779.400 805.050 780.600 ;
        RECT 790.950 778.950 793.050 779.400 ;
        RECT 802.950 778.950 805.050 779.400 ;
        RECT 571.950 777.600 574.050 778.050 ;
        RECT 583.950 777.600 586.050 778.050 ;
        RECT 571.950 776.400 586.050 777.600 ;
        RECT 571.950 775.950 574.050 776.400 ;
        RECT 583.950 775.950 586.050 776.400 ;
        RECT 589.950 777.600 592.050 778.050 ;
        RECT 607.950 777.600 610.050 778.050 ;
        RECT 589.950 776.400 610.050 777.600 ;
        RECT 589.950 775.950 592.050 776.400 ;
        RECT 607.950 775.950 610.050 776.400 ;
        RECT 625.950 775.950 628.050 778.050 ;
        RECT 655.950 777.600 658.050 778.050 ;
        RECT 661.950 777.600 664.050 778.050 ;
        RECT 655.950 776.400 664.050 777.600 ;
        RECT 655.950 775.950 658.050 776.400 ;
        RECT 661.950 775.950 664.050 776.400 ;
        RECT 691.950 777.600 694.050 778.050 ;
        RECT 709.950 777.600 712.050 778.050 ;
        RECT 691.950 776.400 712.050 777.600 ;
        RECT 691.950 775.950 694.050 776.400 ;
        RECT 709.950 775.950 712.050 776.400 ;
        RECT 730.950 777.600 733.050 778.050 ;
        RECT 736.950 777.600 739.050 778.050 ;
        RECT 730.950 776.400 739.050 777.600 ;
        RECT 730.950 775.950 733.050 776.400 ;
        RECT 736.950 775.950 739.050 776.400 ;
        RECT 775.950 777.600 778.050 778.050 ;
        RECT 808.950 777.600 811.050 778.050 ;
        RECT 775.950 776.400 811.050 777.600 ;
        RECT 775.950 775.950 778.050 776.400 ;
        RECT 808.950 775.950 811.050 776.400 ;
        RECT 535.950 774.600 538.050 775.050 ;
        RECT 547.950 774.600 550.050 775.050 ;
        RECT 535.950 773.400 550.050 774.600 ;
        RECT 535.950 772.950 538.050 773.400 ;
        RECT 547.950 772.950 550.050 773.400 ;
        RECT 553.950 774.600 556.050 775.050 ;
        RECT 598.950 774.600 601.050 775.050 ;
        RECT 553.950 773.400 601.050 774.600 ;
        RECT 626.400 774.600 627.600 775.950 ;
        RECT 658.950 774.600 661.050 775.050 ;
        RECT 667.950 774.600 670.050 775.050 ;
        RECT 626.400 773.400 670.050 774.600 ;
        RECT 553.950 772.950 556.050 773.400 ;
        RECT 598.950 772.950 601.050 773.400 ;
        RECT 658.950 772.950 661.050 773.400 ;
        RECT 667.950 772.950 670.050 773.400 ;
        RECT 682.950 772.950 685.050 775.050 ;
        RECT 709.950 774.600 712.050 775.050 ;
        RECT 721.950 774.600 724.050 775.050 ;
        RECT 709.950 773.400 724.050 774.600 ;
        RECT 709.950 772.950 712.050 773.400 ;
        RECT 721.950 772.950 724.050 773.400 ;
        RECT 727.950 774.600 730.050 775.050 ;
        RECT 733.950 774.600 736.050 775.050 ;
        RECT 727.950 773.400 736.050 774.600 ;
        RECT 727.950 772.950 730.050 773.400 ;
        RECT 733.950 772.950 736.050 773.400 ;
        RECT 847.950 774.600 850.050 775.050 ;
        RECT 853.950 774.600 856.050 775.050 ;
        RECT 847.950 773.400 856.050 774.600 ;
        RECT 847.950 772.950 850.050 773.400 ;
        RECT 853.950 772.950 856.050 773.400 ;
        RECT 520.950 770.400 528.600 771.600 ;
        RECT 529.950 771.600 532.050 772.050 ;
        RECT 544.950 771.600 547.050 772.050 ;
        RECT 529.950 770.400 547.050 771.600 ;
        RECT 505.950 769.950 508.050 770.400 ;
        RECT 520.950 769.950 523.050 770.400 ;
        RECT 529.950 769.950 532.050 770.400 ;
        RECT 544.950 769.950 547.050 770.400 ;
        RECT 550.950 771.600 553.050 772.050 ;
        RECT 562.950 771.600 565.050 772.050 ;
        RECT 550.950 770.400 565.050 771.600 ;
        RECT 550.950 769.950 553.050 770.400 ;
        RECT 562.950 769.950 565.050 770.400 ;
        RECT 577.950 771.600 580.050 772.050 ;
        RECT 595.950 771.600 598.050 772.050 ;
        RECT 577.950 770.400 598.050 771.600 ;
        RECT 577.950 769.950 580.050 770.400 ;
        RECT 595.950 769.950 598.050 770.400 ;
        RECT 601.950 771.600 604.050 772.050 ;
        RECT 607.950 771.600 610.050 772.050 ;
        RECT 601.950 770.400 610.050 771.600 ;
        RECT 601.950 769.950 604.050 770.400 ;
        RECT 607.950 769.950 610.050 770.400 ;
        RECT 676.950 771.600 679.050 772.050 ;
        RECT 683.400 771.600 684.600 772.950 ;
        RECT 676.950 770.400 684.600 771.600 ;
        RECT 724.950 771.600 727.050 772.050 ;
        RECT 754.950 771.600 757.050 772.050 ;
        RECT 724.950 770.400 757.050 771.600 ;
        RECT 676.950 769.950 679.050 770.400 ;
        RECT 724.950 769.950 727.050 770.400 ;
        RECT 754.950 769.950 757.050 770.400 ;
        RECT 811.950 771.600 814.050 772.050 ;
        RECT 820.950 771.600 823.050 772.050 ;
        RECT 811.950 770.400 823.050 771.600 ;
        RECT 811.950 769.950 814.050 770.400 ;
        RECT 820.950 769.950 823.050 770.400 ;
        RECT 4.950 768.600 7.050 769.050 ;
        RECT 19.950 768.600 22.050 769.050 ;
        RECT 25.950 768.600 28.050 769.050 ;
        RECT 4.950 767.400 28.050 768.600 ;
        RECT 4.950 766.950 7.050 767.400 ;
        RECT 19.950 766.950 22.050 767.400 ;
        RECT 25.950 766.950 28.050 767.400 ;
        RECT 43.950 768.600 46.050 769.050 ;
        RECT 52.950 768.600 55.050 769.050 ;
        RECT 43.950 767.400 55.050 768.600 ;
        RECT 43.950 766.950 46.050 767.400 ;
        RECT 52.950 766.950 55.050 767.400 ;
        RECT 115.950 768.600 118.050 769.050 ;
        RECT 142.950 768.600 145.050 769.050 ;
        RECT 172.950 768.600 175.050 769.050 ;
        RECT 115.950 767.400 175.050 768.600 ;
        RECT 115.950 766.950 118.050 767.400 ;
        RECT 142.950 766.950 145.050 767.400 ;
        RECT 172.950 766.950 175.050 767.400 ;
        RECT 202.950 768.600 205.050 769.050 ;
        RECT 238.950 768.600 241.050 769.050 ;
        RECT 202.950 767.400 241.050 768.600 ;
        RECT 202.950 766.950 205.050 767.400 ;
        RECT 238.950 766.950 241.050 767.400 ;
        RECT 325.950 768.600 328.050 769.050 ;
        RECT 358.950 768.600 361.050 769.050 ;
        RECT 325.950 767.400 361.050 768.600 ;
        RECT 325.950 766.950 328.050 767.400 ;
        RECT 358.950 766.950 361.050 767.400 ;
        RECT 364.950 768.600 367.050 769.050 ;
        RECT 448.950 768.600 451.050 769.050 ;
        RECT 457.950 768.600 460.050 769.050 ;
        RECT 364.950 767.400 460.050 768.600 ;
        RECT 364.950 766.950 367.050 767.400 ;
        RECT 448.950 766.950 451.050 767.400 ;
        RECT 457.950 766.950 460.050 767.400 ;
        RECT 472.950 768.600 475.050 769.050 ;
        RECT 481.950 768.600 484.050 769.050 ;
        RECT 472.950 767.400 484.050 768.600 ;
        RECT 472.950 766.950 475.050 767.400 ;
        RECT 481.950 766.950 484.050 767.400 ;
        RECT 532.950 768.600 535.050 769.050 ;
        RECT 538.950 768.600 541.050 769.050 ;
        RECT 532.950 767.400 541.050 768.600 ;
        RECT 532.950 766.950 535.050 767.400 ;
        RECT 538.950 766.950 541.050 767.400 ;
        RECT 550.950 768.600 553.050 769.050 ;
        RECT 556.950 768.600 559.050 769.050 ;
        RECT 550.950 767.400 559.050 768.600 ;
        RECT 550.950 766.950 553.050 767.400 ;
        RECT 556.950 766.950 559.050 767.400 ;
        RECT 559.950 768.600 562.050 769.050 ;
        RECT 568.950 768.600 571.050 769.050 ;
        RECT 559.950 767.400 571.050 768.600 ;
        RECT 559.950 766.950 562.050 767.400 ;
        RECT 568.950 766.950 571.050 767.400 ;
        RECT 601.950 768.600 604.050 769.050 ;
        RECT 616.950 768.600 619.050 769.050 ;
        RECT 601.950 767.400 619.050 768.600 ;
        RECT 601.950 766.950 604.050 767.400 ;
        RECT 616.950 766.950 619.050 767.400 ;
        RECT 622.950 768.600 625.050 769.050 ;
        RECT 625.950 768.600 628.050 769.050 ;
        RECT 631.950 768.600 634.050 769.050 ;
        RECT 622.950 767.400 634.050 768.600 ;
        RECT 622.950 766.950 625.050 767.400 ;
        RECT 625.950 766.950 628.050 767.400 ;
        RECT 631.950 766.950 634.050 767.400 ;
        RECT 652.950 768.600 655.050 769.050 ;
        RECT 658.950 768.600 661.050 769.050 ;
        RECT 652.950 767.400 661.050 768.600 ;
        RECT 652.950 766.950 655.050 767.400 ;
        RECT 658.950 766.950 661.050 767.400 ;
        RECT 670.950 768.600 673.050 769.050 ;
        RECT 700.950 768.600 703.050 769.050 ;
        RECT 754.950 768.600 757.050 769.050 ;
        RECT 670.950 767.400 757.050 768.600 ;
        RECT 670.950 766.950 673.050 767.400 ;
        RECT 700.950 766.950 703.050 767.400 ;
        RECT 754.950 766.950 757.050 767.400 ;
        RECT 769.950 768.600 772.050 769.050 ;
        RECT 772.950 768.600 775.050 769.050 ;
        RECT 823.950 768.600 826.050 769.050 ;
        RECT 769.950 767.400 826.050 768.600 ;
        RECT 769.950 766.950 772.050 767.400 ;
        RECT 772.950 766.950 775.050 767.400 ;
        RECT 823.950 766.950 826.050 767.400 ;
        RECT 826.950 768.600 829.050 769.050 ;
        RECT 835.950 768.600 838.050 769.050 ;
        RECT 826.950 767.400 838.050 768.600 ;
        RECT 826.950 766.950 829.050 767.400 ;
        RECT 835.950 766.950 838.050 767.400 ;
        RECT 184.950 765.600 187.050 766.050 ;
        RECT 217.950 765.600 220.050 766.050 ;
        RECT 184.950 764.400 220.050 765.600 ;
        RECT 184.950 763.950 187.050 764.400 ;
        RECT 217.950 763.950 220.050 764.400 ;
        RECT 355.950 765.600 358.050 766.050 ;
        RECT 499.950 765.600 502.050 766.050 ;
        RECT 355.950 764.400 502.050 765.600 ;
        RECT 355.950 763.950 358.050 764.400 ;
        RECT 499.950 763.950 502.050 764.400 ;
        RECT 517.950 765.600 520.050 766.050 ;
        RECT 550.950 765.600 553.050 766.050 ;
        RECT 517.950 764.400 553.050 765.600 ;
        RECT 517.950 763.950 520.050 764.400 ;
        RECT 550.950 763.950 553.050 764.400 ;
        RECT 580.950 765.600 583.050 766.050 ;
        RECT 643.950 765.600 646.050 766.050 ;
        RECT 649.950 765.600 652.050 766.050 ;
        RECT 580.950 764.400 652.050 765.600 ;
        RECT 580.950 763.950 583.050 764.400 ;
        RECT 643.950 763.950 646.050 764.400 ;
        RECT 649.950 763.950 652.050 764.400 ;
        RECT 676.950 765.600 679.050 766.050 ;
        RECT 682.950 765.600 685.050 766.050 ;
        RECT 676.950 764.400 685.050 765.600 ;
        RECT 676.950 763.950 679.050 764.400 ;
        RECT 682.950 763.950 685.050 764.400 ;
        RECT 685.950 765.600 688.050 766.050 ;
        RECT 712.950 765.600 715.050 766.050 ;
        RECT 724.950 765.600 727.050 766.050 ;
        RECT 685.950 764.400 727.050 765.600 ;
        RECT 685.950 763.950 688.050 764.400 ;
        RECT 712.950 763.950 715.050 764.400 ;
        RECT 724.950 763.950 727.050 764.400 ;
        RECT 16.950 762.600 19.050 763.050 ;
        RECT 22.950 762.600 25.050 763.050 ;
        RECT 124.950 762.600 127.050 763.050 ;
        RECT 16.950 761.400 127.050 762.600 ;
        RECT 16.950 760.950 19.050 761.400 ;
        RECT 22.950 760.950 25.050 761.400 ;
        RECT 124.950 760.950 127.050 761.400 ;
        RECT 301.950 762.600 304.050 763.050 ;
        RECT 367.950 762.600 370.050 763.050 ;
        RECT 301.950 761.400 370.050 762.600 ;
        RECT 301.950 760.950 304.050 761.400 ;
        RECT 367.950 760.950 370.050 761.400 ;
        RECT 433.950 762.600 436.050 763.050 ;
        RECT 466.950 762.600 469.050 763.050 ;
        RECT 433.950 761.400 469.050 762.600 ;
        RECT 433.950 760.950 436.050 761.400 ;
        RECT 466.950 760.950 469.050 761.400 ;
        RECT 76.950 759.600 79.050 760.050 ;
        RECT 91.950 759.600 94.050 760.050 ;
        RECT 76.950 758.400 94.050 759.600 ;
        RECT 76.950 757.950 79.050 758.400 ;
        RECT 91.950 757.950 94.050 758.400 ;
        RECT 283.950 759.600 286.050 760.050 ;
        RECT 304.950 759.600 307.050 760.050 ;
        RECT 283.950 758.400 307.050 759.600 ;
        RECT 283.950 757.950 286.050 758.400 ;
        RECT 304.950 757.950 307.050 758.400 ;
        RECT 466.950 759.600 469.050 760.050 ;
        RECT 535.950 759.600 538.050 760.050 ;
        RECT 466.950 758.400 538.050 759.600 ;
        RECT 466.950 757.950 469.050 758.400 ;
        RECT 535.950 757.950 538.050 758.400 ;
        RECT 592.950 759.600 595.050 760.050 ;
        RECT 655.950 759.600 658.050 760.050 ;
        RECT 706.950 759.600 709.050 760.050 ;
        RECT 760.950 759.600 763.050 760.050 ;
        RECT 592.950 758.400 763.050 759.600 ;
        RECT 592.950 757.950 595.050 758.400 ;
        RECT 655.950 757.950 658.050 758.400 ;
        RECT 706.950 757.950 709.050 758.400 ;
        RECT 760.950 757.950 763.050 758.400 ;
        RECT 772.950 759.600 775.050 760.050 ;
        RECT 778.950 759.600 781.050 760.050 ;
        RECT 772.950 758.400 781.050 759.600 ;
        RECT 772.950 757.950 775.050 758.400 ;
        RECT 778.950 757.950 781.050 758.400 ;
        RECT 28.950 756.600 31.050 757.050 ;
        RECT 55.950 756.600 58.050 757.050 ;
        RECT 28.950 755.400 58.050 756.600 ;
        RECT 28.950 754.950 31.050 755.400 ;
        RECT 55.950 754.950 58.050 755.400 ;
        RECT 118.950 756.600 121.050 757.050 ;
        RECT 178.950 756.600 181.050 757.050 ;
        RECT 265.950 756.600 268.050 757.050 ;
        RECT 118.950 755.400 268.050 756.600 ;
        RECT 118.950 754.950 121.050 755.400 ;
        RECT 178.950 754.950 181.050 755.400 ;
        RECT 265.950 754.950 268.050 755.400 ;
        RECT 277.950 756.600 280.050 757.050 ;
        RECT 295.950 756.600 298.050 757.050 ;
        RECT 277.950 755.400 298.050 756.600 ;
        RECT 277.950 754.950 280.050 755.400 ;
        RECT 295.950 754.950 298.050 755.400 ;
        RECT 379.950 756.600 382.050 757.050 ;
        RECT 406.950 756.600 409.050 757.050 ;
        RECT 379.950 755.400 409.050 756.600 ;
        RECT 379.950 754.950 382.050 755.400 ;
        RECT 406.950 754.950 409.050 755.400 ;
        RECT 409.950 756.600 412.050 757.050 ;
        RECT 421.950 756.600 424.050 757.050 ;
        RECT 409.950 755.400 424.050 756.600 ;
        RECT 409.950 754.950 412.050 755.400 ;
        RECT 421.950 754.950 424.050 755.400 ;
        RECT 640.950 756.600 643.050 757.050 ;
        RECT 652.950 756.600 655.050 757.050 ;
        RECT 640.950 755.400 655.050 756.600 ;
        RECT 640.950 754.950 643.050 755.400 ;
        RECT 652.950 754.950 655.050 755.400 ;
        RECT 760.950 756.600 763.050 757.050 ;
        RECT 778.950 756.600 781.050 757.050 ;
        RECT 760.950 755.400 781.050 756.600 ;
        RECT 760.950 754.950 763.050 755.400 ;
        RECT 778.950 754.950 781.050 755.400 ;
        RECT 784.950 756.600 787.050 757.050 ;
        RECT 805.950 756.600 808.050 757.050 ;
        RECT 784.950 755.400 808.050 756.600 ;
        RECT 784.950 754.950 787.050 755.400 ;
        RECT 805.950 754.950 808.050 755.400 ;
        RECT 55.950 753.600 58.050 754.050 ;
        RECT 118.950 753.600 121.050 754.050 ;
        RECT 55.950 752.400 121.050 753.600 ;
        RECT 55.950 751.950 58.050 752.400 ;
        RECT 118.950 751.950 121.050 752.400 ;
        RECT 238.950 753.600 241.050 754.050 ;
        RECT 244.950 753.600 247.050 754.050 ;
        RECT 292.950 753.600 295.050 754.050 ;
        RECT 238.950 752.400 295.050 753.600 ;
        RECT 238.950 751.950 241.050 752.400 ;
        RECT 244.950 751.950 247.050 752.400 ;
        RECT 292.950 751.950 295.050 752.400 ;
        RECT 322.950 753.600 325.050 754.050 ;
        RECT 397.950 753.600 400.050 754.050 ;
        RECT 322.950 752.400 400.050 753.600 ;
        RECT 322.950 751.950 325.050 752.400 ;
        RECT 397.950 751.950 400.050 752.400 ;
        RECT 400.950 753.600 403.050 754.050 ;
        RECT 418.950 753.600 421.050 754.050 ;
        RECT 400.950 752.400 421.050 753.600 ;
        RECT 400.950 751.950 403.050 752.400 ;
        RECT 418.950 751.950 421.050 752.400 ;
        RECT 478.950 753.600 481.050 754.050 ;
        RECT 526.950 753.600 529.050 754.050 ;
        RECT 478.950 752.400 529.050 753.600 ;
        RECT 478.950 751.950 481.050 752.400 ;
        RECT 526.950 751.950 529.050 752.400 ;
        RECT 565.950 753.600 568.050 754.050 ;
        RECT 640.950 753.600 643.050 754.050 ;
        RECT 643.950 753.600 646.050 754.050 ;
        RECT 679.950 753.600 682.050 754.050 ;
        RECT 565.950 752.400 682.050 753.600 ;
        RECT 565.950 751.950 568.050 752.400 ;
        RECT 640.950 751.950 643.050 752.400 ;
        RECT 643.950 751.950 646.050 752.400 ;
        RECT 679.950 751.950 682.050 752.400 ;
        RECT 91.950 750.600 94.050 751.050 ;
        RECT 148.950 750.600 151.050 751.050 ;
        RECT 91.950 749.400 151.050 750.600 ;
        RECT 91.950 748.950 94.050 749.400 ;
        RECT 148.950 748.950 151.050 749.400 ;
        RECT 151.950 750.600 154.050 751.050 ;
        RECT 247.950 750.600 250.050 751.050 ;
        RECT 322.950 750.600 325.050 751.050 ;
        RECT 151.950 749.400 325.050 750.600 ;
        RECT 151.950 748.950 154.050 749.400 ;
        RECT 247.950 748.950 250.050 749.400 ;
        RECT 322.950 748.950 325.050 749.400 ;
        RECT 331.950 750.600 334.050 751.050 ;
        RECT 346.950 750.600 349.050 751.050 ;
        RECT 331.950 749.400 349.050 750.600 ;
        RECT 331.950 748.950 334.050 749.400 ;
        RECT 346.950 748.950 349.050 749.400 ;
        RECT 367.950 750.600 370.050 751.050 ;
        RECT 439.950 750.600 442.050 751.050 ;
        RECT 367.950 749.400 442.050 750.600 ;
        RECT 367.950 748.950 370.050 749.400 ;
        RECT 439.950 748.950 442.050 749.400 ;
        RECT 451.950 750.600 454.050 751.050 ;
        RECT 463.950 750.600 466.050 751.050 ;
        RECT 475.950 750.600 478.050 751.050 ;
        RECT 451.950 749.400 478.050 750.600 ;
        RECT 451.950 748.950 454.050 749.400 ;
        RECT 463.950 748.950 466.050 749.400 ;
        RECT 475.950 748.950 478.050 749.400 ;
        RECT 508.950 750.600 511.050 751.050 ;
        RECT 514.950 750.600 517.050 751.050 ;
        RECT 508.950 749.400 517.050 750.600 ;
        RECT 508.950 748.950 511.050 749.400 ;
        RECT 514.950 748.950 517.050 749.400 ;
        RECT 562.950 750.600 565.050 751.050 ;
        RECT 586.950 750.600 589.050 751.050 ;
        RECT 562.950 749.400 589.050 750.600 ;
        RECT 562.950 748.950 565.050 749.400 ;
        RECT 586.950 748.950 589.050 749.400 ;
        RECT 733.950 750.600 736.050 751.050 ;
        RECT 742.950 750.600 745.050 751.050 ;
        RECT 763.950 750.600 766.050 751.050 ;
        RECT 733.950 749.400 766.050 750.600 ;
        RECT 733.950 748.950 736.050 749.400 ;
        RECT 742.950 748.950 745.050 749.400 ;
        RECT 763.950 748.950 766.050 749.400 ;
        RECT 829.950 750.600 832.050 751.050 ;
        RECT 850.950 750.600 853.050 751.050 ;
        RECT 829.950 749.400 853.050 750.600 ;
        RECT 829.950 748.950 832.050 749.400 ;
        RECT 850.950 748.950 853.050 749.400 ;
        RECT 58.950 747.600 61.050 748.050 ;
        RECT 73.950 747.600 76.050 748.050 ;
        RECT 118.950 747.600 121.050 748.050 ;
        RECT 58.950 746.400 121.050 747.600 ;
        RECT 58.950 745.950 61.050 746.400 ;
        RECT 73.950 745.950 76.050 746.400 ;
        RECT 118.950 745.950 121.050 746.400 ;
        RECT 145.950 747.600 148.050 748.050 ;
        RECT 157.950 747.600 160.050 748.050 ;
        RECT 205.950 747.600 208.050 748.050 ;
        RECT 145.950 746.400 150.600 747.600 ;
        RECT 145.950 745.950 148.050 746.400 ;
        RECT 79.950 744.600 82.050 745.050 ;
        RECT 97.950 744.600 100.050 745.050 ;
        RECT 79.950 743.400 100.050 744.600 ;
        RECT 79.950 742.950 82.050 743.400 ;
        RECT 97.950 742.950 100.050 743.400 ;
        RECT 103.950 744.600 106.050 745.050 ;
        RECT 109.950 744.600 112.050 745.050 ;
        RECT 103.950 743.400 112.050 744.600 ;
        RECT 149.400 744.600 150.600 746.400 ;
        RECT 157.950 746.400 208.050 747.600 ;
        RECT 157.950 745.950 160.050 746.400 ;
        RECT 205.950 745.950 208.050 746.400 ;
        RECT 289.950 747.600 292.050 748.050 ;
        RECT 307.950 747.600 310.050 748.050 ;
        RECT 289.950 746.400 310.050 747.600 ;
        RECT 289.950 745.950 292.050 746.400 ;
        RECT 307.950 745.950 310.050 746.400 ;
        RECT 319.950 747.600 322.050 748.050 ;
        RECT 343.950 747.600 346.050 748.050 ;
        RECT 373.950 747.600 376.050 748.050 ;
        RECT 319.950 746.400 376.050 747.600 ;
        RECT 319.950 745.950 322.050 746.400 ;
        RECT 343.950 745.950 346.050 746.400 ;
        RECT 373.950 745.950 376.050 746.400 ;
        RECT 397.950 747.600 400.050 748.050 ;
        RECT 466.950 747.600 469.050 748.050 ;
        RECT 397.950 746.400 469.050 747.600 ;
        RECT 397.950 745.950 400.050 746.400 ;
        RECT 466.950 745.950 469.050 746.400 ;
        RECT 502.950 747.600 505.050 748.050 ;
        RECT 535.950 747.600 538.050 748.050 ;
        RECT 577.950 747.600 580.050 748.050 ;
        RECT 502.950 746.400 516.600 747.600 ;
        RECT 502.950 745.950 505.050 746.400 ;
        RECT 163.950 744.600 166.050 745.050 ;
        RECT 149.400 743.400 166.050 744.600 ;
        RECT 103.950 742.950 106.050 743.400 ;
        RECT 109.950 742.950 112.050 743.400 ;
        RECT 163.950 742.950 166.050 743.400 ;
        RECT 235.950 744.600 238.050 745.050 ;
        RECT 241.950 744.600 244.050 745.050 ;
        RECT 235.950 743.400 244.050 744.600 ;
        RECT 235.950 742.950 238.050 743.400 ;
        RECT 241.950 742.950 244.050 743.400 ;
        RECT 274.950 744.600 277.050 745.050 ;
        RECT 331.950 744.600 334.050 745.050 ;
        RECT 337.950 744.600 340.050 745.050 ;
        RECT 274.950 743.400 340.050 744.600 ;
        RECT 274.950 742.950 277.050 743.400 ;
        RECT 331.950 742.950 334.050 743.400 ;
        RECT 337.950 742.950 340.050 743.400 ;
        RECT 391.950 744.600 394.050 745.050 ;
        RECT 442.950 744.600 445.050 745.050 ;
        RECT 454.950 744.600 457.050 745.050 ;
        RECT 391.950 743.400 408.600 744.600 ;
        RECT 391.950 742.950 394.050 743.400 ;
        RECT 106.950 741.600 109.050 742.050 ;
        RECT 127.950 741.600 130.050 742.050 ;
        RECT 106.950 740.400 130.050 741.600 ;
        RECT 106.950 739.950 109.050 740.400 ;
        RECT 127.950 739.950 130.050 740.400 ;
        RECT 142.950 741.600 145.050 742.050 ;
        RECT 148.950 741.600 151.050 742.050 ;
        RECT 142.950 740.400 151.050 741.600 ;
        RECT 142.950 739.950 145.050 740.400 ;
        RECT 148.950 739.950 151.050 740.400 ;
        RECT 268.950 741.600 271.050 742.050 ;
        RECT 286.950 741.600 289.050 742.050 ;
        RECT 268.950 740.400 289.050 741.600 ;
        RECT 268.950 739.950 271.050 740.400 ;
        RECT 286.950 739.950 289.050 740.400 ;
        RECT 349.950 741.600 352.050 742.050 ;
        RECT 361.950 741.600 364.050 742.050 ;
        RECT 349.950 740.400 364.050 741.600 ;
        RECT 349.950 739.950 352.050 740.400 ;
        RECT 361.950 739.950 364.050 740.400 ;
        RECT 67.950 738.600 70.050 739.050 ;
        RECT 115.950 738.600 118.050 739.050 ;
        RECT 67.950 737.400 118.050 738.600 ;
        RECT 67.950 736.950 70.050 737.400 ;
        RECT 115.950 736.950 118.050 737.400 ;
        RECT 157.950 738.600 160.050 739.050 ;
        RECT 184.950 738.600 187.050 739.050 ;
        RECT 157.950 737.400 187.050 738.600 ;
        RECT 157.950 736.950 160.050 737.400 ;
        RECT 184.950 736.950 187.050 737.400 ;
        RECT 382.950 738.600 385.050 739.050 ;
        RECT 397.950 738.600 400.050 739.050 ;
        RECT 382.950 737.400 400.050 738.600 ;
        RECT 407.400 738.600 408.600 743.400 ;
        RECT 442.950 743.400 457.050 744.600 ;
        RECT 442.950 742.950 445.050 743.400 ;
        RECT 454.950 742.950 457.050 743.400 ;
        RECT 511.950 742.950 514.050 745.050 ;
        RECT 515.400 744.600 516.600 746.400 ;
        RECT 535.950 746.400 580.050 747.600 ;
        RECT 535.950 745.950 538.050 746.400 ;
        RECT 577.950 745.950 580.050 746.400 ;
        RECT 586.950 747.600 589.050 748.050 ;
        RECT 604.950 747.600 607.050 748.050 ;
        RECT 607.950 747.600 610.050 748.050 ;
        RECT 586.950 746.400 610.050 747.600 ;
        RECT 586.950 745.950 589.050 746.400 ;
        RECT 604.950 745.950 607.050 746.400 ;
        RECT 607.950 745.950 610.050 746.400 ;
        RECT 619.950 747.600 622.050 748.050 ;
        RECT 661.950 747.600 664.050 748.050 ;
        RECT 619.950 746.400 664.050 747.600 ;
        RECT 619.950 745.950 622.050 746.400 ;
        RECT 661.950 745.950 664.050 746.400 ;
        RECT 673.950 747.600 676.050 748.050 ;
        RECT 679.950 747.600 682.050 748.050 ;
        RECT 673.950 746.400 682.050 747.600 ;
        RECT 673.950 745.950 676.050 746.400 ;
        RECT 679.950 745.950 682.050 746.400 ;
        RECT 715.950 747.600 718.050 748.050 ;
        RECT 736.950 747.600 739.050 748.050 ;
        RECT 745.950 747.600 748.050 748.050 ;
        RECT 715.950 746.400 748.050 747.600 ;
        RECT 715.950 745.950 718.050 746.400 ;
        RECT 736.950 745.950 739.050 746.400 ;
        RECT 745.950 745.950 748.050 746.400 ;
        RECT 748.950 745.950 751.050 748.050 ;
        RECT 751.950 747.600 754.050 748.050 ;
        RECT 766.950 747.600 769.050 748.050 ;
        RECT 751.950 746.400 769.050 747.600 ;
        RECT 751.950 745.950 754.050 746.400 ;
        RECT 766.950 745.950 769.050 746.400 ;
        RECT 769.950 747.600 772.050 748.050 ;
        RECT 790.950 747.600 793.050 748.050 ;
        RECT 769.950 746.400 793.050 747.600 ;
        RECT 769.950 745.950 772.050 746.400 ;
        RECT 790.950 745.950 793.050 746.400 ;
        RECT 850.950 747.600 853.050 748.050 ;
        RECT 856.950 747.600 859.050 748.050 ;
        RECT 850.950 746.400 859.050 747.600 ;
        RECT 850.950 745.950 853.050 746.400 ;
        RECT 856.950 745.950 859.050 746.400 ;
        RECT 595.950 744.600 598.050 745.050 ;
        RECT 604.950 744.600 607.050 745.050 ;
        RECT 515.400 743.400 598.050 744.600 ;
        RECT 595.950 742.950 598.050 743.400 ;
        RECT 599.400 743.400 607.050 744.600 ;
        RECT 415.950 741.600 418.050 742.050 ;
        RECT 433.950 741.600 436.050 742.050 ;
        RECT 415.950 740.400 436.050 741.600 ;
        RECT 415.950 739.950 418.050 740.400 ;
        RECT 433.950 739.950 436.050 740.400 ;
        RECT 475.950 741.600 478.050 742.050 ;
        RECT 484.950 741.600 487.050 742.050 ;
        RECT 475.950 740.400 487.050 741.600 ;
        RECT 475.950 739.950 478.050 740.400 ;
        RECT 484.950 739.950 487.050 740.400 ;
        RECT 499.950 741.600 502.050 742.050 ;
        RECT 508.950 741.600 511.050 742.050 ;
        RECT 499.950 740.400 511.050 741.600 ;
        RECT 512.400 741.600 513.600 742.950 ;
        RECT 514.950 741.600 517.050 742.050 ;
        RECT 512.400 740.400 517.050 741.600 ;
        RECT 499.950 739.950 502.050 740.400 ;
        RECT 508.950 739.950 511.050 740.400 ;
        RECT 514.950 739.950 517.050 740.400 ;
        RECT 541.950 741.600 544.050 742.050 ;
        RECT 568.950 741.600 571.050 742.050 ;
        RECT 577.950 741.600 580.050 742.050 ;
        RECT 541.950 740.400 561.600 741.600 ;
        RECT 541.950 739.950 544.050 740.400 ;
        RECT 560.400 739.050 561.600 740.400 ;
        RECT 568.950 740.400 580.050 741.600 ;
        RECT 568.950 739.950 571.050 740.400 ;
        RECT 577.950 739.950 580.050 740.400 ;
        RECT 421.950 738.600 424.050 739.050 ;
        RECT 407.400 737.400 424.050 738.600 ;
        RECT 382.950 736.950 385.050 737.400 ;
        RECT 397.950 736.950 400.050 737.400 ;
        RECT 421.950 736.950 424.050 737.400 ;
        RECT 487.950 738.600 490.050 739.050 ;
        RECT 493.950 738.600 496.050 739.050 ;
        RECT 487.950 737.400 496.050 738.600 ;
        RECT 487.950 736.950 490.050 737.400 ;
        RECT 493.950 736.950 496.050 737.400 ;
        RECT 520.950 738.600 523.050 739.050 ;
        RECT 538.950 738.600 541.050 739.050 ;
        RECT 520.950 737.400 541.050 738.600 ;
        RECT 520.950 736.950 523.050 737.400 ;
        RECT 538.950 736.950 541.050 737.400 ;
        RECT 559.950 736.950 562.050 739.050 ;
        RECT 574.950 738.600 577.050 739.050 ;
        RECT 599.400 738.600 600.600 743.400 ;
        RECT 604.950 742.950 607.050 743.400 ;
        RECT 613.950 742.950 616.050 745.050 ;
        RECT 616.950 744.600 619.050 745.050 ;
        RECT 664.950 744.600 667.050 745.050 ;
        RECT 694.950 744.600 697.050 745.050 ;
        RECT 616.950 743.400 697.050 744.600 ;
        RECT 749.400 744.600 750.600 745.950 ;
        RECT 751.950 744.600 754.050 745.050 ;
        RECT 749.400 743.400 754.050 744.600 ;
        RECT 616.950 742.950 619.050 743.400 ;
        RECT 664.950 742.950 667.050 743.400 ;
        RECT 694.950 742.950 697.050 743.400 ;
        RECT 751.950 742.950 754.050 743.400 ;
        RECT 781.950 744.600 784.050 745.050 ;
        RECT 853.950 744.600 856.050 745.050 ;
        RECT 781.950 743.400 856.050 744.600 ;
        RECT 781.950 742.950 784.050 743.400 ;
        RECT 853.950 742.950 856.050 743.400 ;
        RECT 614.400 741.600 615.600 742.950 ;
        RECT 634.950 741.600 637.050 742.050 ;
        RECT 685.950 741.600 688.050 742.050 ;
        RECT 614.400 740.400 633.600 741.600 ;
        RECT 632.400 739.050 633.600 740.400 ;
        RECT 634.950 740.400 688.050 741.600 ;
        RECT 634.950 739.950 637.050 740.400 ;
        RECT 685.950 739.950 688.050 740.400 ;
        RECT 742.950 741.600 745.050 742.050 ;
        RECT 748.950 741.600 751.050 742.050 ;
        RECT 742.950 740.400 751.050 741.600 ;
        RECT 742.950 739.950 745.050 740.400 ;
        RECT 748.950 739.950 751.050 740.400 ;
        RECT 574.950 737.400 600.600 738.600 ;
        RECT 610.950 738.600 613.050 739.050 ;
        RECT 619.950 738.600 622.050 739.050 ;
        RECT 610.950 737.400 622.050 738.600 ;
        RECT 574.950 736.950 577.050 737.400 ;
        RECT 610.950 736.950 613.050 737.400 ;
        RECT 619.950 736.950 622.050 737.400 ;
        RECT 631.950 736.950 634.050 739.050 ;
        RECT 661.950 736.950 664.050 739.050 ;
        RECT 667.950 738.600 670.050 739.050 ;
        RECT 676.950 738.600 679.050 739.050 ;
        RECT 694.950 738.600 697.050 739.050 ;
        RECT 667.950 737.400 697.050 738.600 ;
        RECT 667.950 736.950 670.050 737.400 ;
        RECT 676.950 736.950 679.050 737.400 ;
        RECT 694.950 736.950 697.050 737.400 ;
        RECT 778.950 738.600 781.050 739.050 ;
        RECT 817.950 738.600 820.050 739.050 ;
        RECT 778.950 737.400 820.050 738.600 ;
        RECT 778.950 736.950 781.050 737.400 ;
        RECT 817.950 736.950 820.050 737.400 ;
        RECT 109.950 735.600 112.050 736.050 ;
        RECT 124.950 735.600 127.050 736.050 ;
        RECT 109.950 734.400 127.050 735.600 ;
        RECT 109.950 733.950 112.050 734.400 ;
        RECT 124.950 733.950 127.050 734.400 ;
        RECT 148.950 735.600 151.050 736.050 ;
        RECT 262.950 735.600 265.050 736.050 ;
        RECT 295.950 735.600 298.050 736.050 ;
        RECT 301.950 735.600 304.050 736.050 ;
        RECT 148.950 734.400 304.050 735.600 ;
        RECT 148.950 733.950 151.050 734.400 ;
        RECT 262.950 733.950 265.050 734.400 ;
        RECT 295.950 733.950 298.050 734.400 ;
        RECT 301.950 733.950 304.050 734.400 ;
        RECT 469.950 735.600 472.050 736.050 ;
        RECT 499.950 735.600 502.050 736.050 ;
        RECT 505.950 735.600 508.050 736.050 ;
        RECT 469.950 734.400 508.050 735.600 ;
        RECT 469.950 733.950 472.050 734.400 ;
        RECT 499.950 733.950 502.050 734.400 ;
        RECT 505.950 733.950 508.050 734.400 ;
        RECT 544.950 735.600 547.050 736.050 ;
        RECT 610.950 735.600 613.050 736.050 ;
        RECT 544.950 734.400 613.050 735.600 ;
        RECT 544.950 733.950 547.050 734.400 ;
        RECT 610.950 733.950 613.050 734.400 ;
        RECT 646.950 735.600 649.050 736.050 ;
        RECT 652.950 735.600 655.050 736.050 ;
        RECT 646.950 734.400 655.050 735.600 ;
        RECT 662.400 735.600 663.600 736.950 ;
        RECT 688.950 735.600 691.050 736.050 ;
        RECT 706.950 735.600 709.050 736.050 ;
        RECT 662.400 734.400 709.050 735.600 ;
        RECT 646.950 733.950 649.050 734.400 ;
        RECT 652.950 733.950 655.050 734.400 ;
        RECT 688.950 733.950 691.050 734.400 ;
        RECT 706.950 733.950 709.050 734.400 ;
        RECT 841.950 735.600 844.050 736.050 ;
        RECT 853.950 735.600 856.050 736.050 ;
        RECT 841.950 734.400 856.050 735.600 ;
        RECT 841.950 733.950 844.050 734.400 ;
        RECT 853.950 733.950 856.050 734.400 ;
        RECT 118.950 732.600 121.050 733.050 ;
        RECT 154.950 732.600 157.050 733.050 ;
        RECT 208.950 732.600 211.050 733.050 ;
        RECT 289.950 732.600 292.050 733.050 ;
        RECT 118.950 731.400 292.050 732.600 ;
        RECT 118.950 730.950 121.050 731.400 ;
        RECT 154.950 730.950 157.050 731.400 ;
        RECT 208.950 730.950 211.050 731.400 ;
        RECT 289.950 730.950 292.050 731.400 ;
        RECT 394.950 732.600 397.050 733.050 ;
        RECT 583.950 732.600 586.050 733.050 ;
        RECT 394.950 731.400 586.050 732.600 ;
        RECT 394.950 730.950 397.050 731.400 ;
        RECT 533.400 730.050 534.600 731.400 ;
        RECT 583.950 730.950 586.050 731.400 ;
        RECT 532.950 727.950 535.050 730.050 ;
        RECT 502.950 726.600 505.050 727.050 ;
        RECT 550.950 726.600 553.050 727.050 ;
        RECT 502.950 725.400 553.050 726.600 ;
        RECT 502.950 724.950 505.050 725.400 ;
        RECT 550.950 724.950 553.050 725.400 ;
        RECT 580.950 726.600 583.050 727.050 ;
        RECT 646.950 726.600 649.050 727.050 ;
        RECT 580.950 725.400 649.050 726.600 ;
        RECT 580.950 724.950 583.050 725.400 ;
        RECT 646.950 724.950 649.050 725.400 ;
        RECT 655.950 726.600 658.050 727.050 ;
        RECT 757.950 726.600 760.050 727.050 ;
        RECT 766.950 726.600 769.050 727.050 ;
        RECT 655.950 725.400 769.050 726.600 ;
        RECT 655.950 724.950 658.050 725.400 ;
        RECT 757.950 724.950 760.050 725.400 ;
        RECT 766.950 724.950 769.050 725.400 ;
        RECT 826.950 726.600 829.050 727.050 ;
        RECT 847.950 726.600 850.050 727.050 ;
        RECT 826.950 725.400 850.050 726.600 ;
        RECT 826.950 724.950 829.050 725.400 ;
        RECT 847.950 724.950 850.050 725.400 ;
        RECT 166.950 720.600 169.050 721.050 ;
        RECT 220.950 720.600 223.050 721.050 ;
        RECT 166.950 719.400 223.050 720.600 ;
        RECT 166.950 718.950 169.050 719.400 ;
        RECT 220.950 718.950 223.050 719.400 ;
        RECT 28.950 717.600 31.050 718.050 ;
        RECT 58.950 717.600 61.050 718.050 ;
        RECT 28.950 716.400 61.050 717.600 ;
        RECT 28.950 715.950 31.050 716.400 ;
        RECT 58.950 715.950 61.050 716.400 ;
        RECT 112.950 717.600 115.050 718.050 ;
        RECT 157.950 717.600 160.050 718.050 ;
        RECT 112.950 716.400 160.050 717.600 ;
        RECT 112.950 715.950 115.050 716.400 ;
        RECT 157.950 715.950 160.050 716.400 ;
        RECT 187.950 717.600 190.050 718.050 ;
        RECT 313.950 717.600 316.050 718.050 ;
        RECT 379.950 717.600 382.050 718.050 ;
        RECT 187.950 716.400 382.050 717.600 ;
        RECT 187.950 715.950 190.050 716.400 ;
        RECT 313.950 715.950 316.050 716.400 ;
        RECT 379.950 715.950 382.050 716.400 ;
        RECT 751.950 717.600 754.050 718.050 ;
        RECT 769.950 717.600 772.050 718.050 ;
        RECT 751.950 716.400 772.050 717.600 ;
        RECT 751.950 715.950 754.050 716.400 ;
        RECT 769.950 715.950 772.050 716.400 ;
        RECT 4.950 714.600 7.050 715.050 ;
        RECT 34.950 714.600 37.050 715.050 ;
        RECT 70.950 714.600 73.050 715.050 ;
        RECT 208.950 714.600 211.050 715.050 ;
        RECT 4.950 713.400 211.050 714.600 ;
        RECT 4.950 712.950 7.050 713.400 ;
        RECT 34.950 712.950 37.050 713.400 ;
        RECT 70.950 712.950 73.050 713.400 ;
        RECT 208.950 712.950 211.050 713.400 ;
        RECT 214.950 714.600 217.050 715.050 ;
        RECT 325.950 714.600 328.050 715.050 ;
        RECT 214.950 713.400 328.050 714.600 ;
        RECT 214.950 712.950 217.050 713.400 ;
        RECT 325.950 712.950 328.050 713.400 ;
        RECT 451.950 714.600 454.050 715.050 ;
        RECT 496.950 714.600 499.050 715.050 ;
        RECT 451.950 713.400 499.050 714.600 ;
        RECT 451.950 712.950 454.050 713.400 ;
        RECT 496.950 712.950 499.050 713.400 ;
        RECT 169.950 711.600 172.050 712.050 ;
        RECT 178.950 711.600 181.050 712.050 ;
        RECT 286.950 711.600 289.050 712.050 ;
        RECT 316.950 711.600 319.050 712.050 ;
        RECT 169.950 710.400 319.050 711.600 ;
        RECT 169.950 709.950 172.050 710.400 ;
        RECT 178.950 709.950 181.050 710.400 ;
        RECT 286.950 709.950 289.050 710.400 ;
        RECT 316.950 709.950 319.050 710.400 ;
        RECT 433.950 711.600 436.050 712.050 ;
        RECT 451.950 711.600 454.050 712.050 ;
        RECT 433.950 710.400 454.050 711.600 ;
        RECT 433.950 709.950 436.050 710.400 ;
        RECT 451.950 709.950 454.050 710.400 ;
        RECT 478.950 711.600 481.050 712.050 ;
        RECT 553.950 711.600 556.050 712.050 ;
        RECT 559.950 711.600 562.050 712.050 ;
        RECT 634.950 711.600 637.050 712.050 ;
        RECT 637.950 711.600 640.050 712.050 ;
        RECT 478.950 710.400 562.050 711.600 ;
        RECT 632.400 710.400 640.050 711.600 ;
        RECT 478.950 709.950 481.050 710.400 ;
        RECT 553.950 709.950 556.050 710.400 ;
        RECT 559.950 709.950 562.050 710.400 ;
        RECT 634.950 709.950 637.050 710.400 ;
        RECT 637.950 709.950 640.050 710.400 ;
        RECT 13.950 708.600 16.050 709.050 ;
        RECT 25.950 708.600 28.050 709.050 ;
        RECT 121.950 708.600 124.050 709.050 ;
        RECT 13.950 707.400 124.050 708.600 ;
        RECT 13.950 706.950 16.050 707.400 ;
        RECT 25.950 706.950 28.050 707.400 ;
        RECT 121.950 706.950 124.050 707.400 ;
        RECT 142.950 708.600 145.050 709.050 ;
        RECT 187.950 708.600 190.050 709.050 ;
        RECT 142.950 707.400 190.050 708.600 ;
        RECT 142.950 706.950 145.050 707.400 ;
        RECT 187.950 706.950 190.050 707.400 ;
        RECT 262.950 708.600 265.050 709.050 ;
        RECT 268.950 708.600 271.050 709.050 ;
        RECT 262.950 707.400 271.050 708.600 ;
        RECT 262.950 706.950 265.050 707.400 ;
        RECT 268.950 706.950 271.050 707.400 ;
        RECT 298.950 708.600 301.050 709.050 ;
        RECT 313.950 708.600 316.050 709.050 ;
        RECT 337.950 708.600 340.050 709.050 ;
        RECT 298.950 707.400 340.050 708.600 ;
        RECT 298.950 706.950 301.050 707.400 ;
        RECT 313.950 706.950 316.050 707.400 ;
        RECT 337.950 706.950 340.050 707.400 ;
        RECT 370.950 708.600 373.050 709.050 ;
        RECT 436.950 708.600 439.050 709.050 ;
        RECT 445.950 708.600 448.050 709.050 ;
        RECT 448.950 708.600 451.050 709.050 ;
        RECT 370.950 707.400 393.600 708.600 ;
        RECT 370.950 706.950 373.050 707.400 ;
        RECT 392.400 706.050 393.600 707.400 ;
        RECT 436.950 707.400 451.050 708.600 ;
        RECT 436.950 706.950 439.050 707.400 ;
        RECT 445.950 706.950 448.050 707.400 ;
        RECT 448.950 706.950 451.050 707.400 ;
        RECT 463.950 708.600 466.050 709.050 ;
        RECT 481.950 708.600 484.050 709.050 ;
        RECT 463.950 707.400 513.600 708.600 ;
        RECT 463.950 706.950 466.050 707.400 ;
        RECT 481.950 706.950 484.050 707.400 ;
        RECT 7.950 705.600 10.050 706.050 ;
        RECT 82.950 705.600 85.050 706.050 ;
        RECT 97.950 705.600 100.050 706.050 ;
        RECT 127.950 705.600 130.050 706.050 ;
        RECT 7.950 704.400 15.600 705.600 ;
        RECT 7.950 703.950 10.050 704.400 ;
        RECT 10.950 702.600 13.050 703.050 ;
        RECT 8.400 701.400 13.050 702.600 ;
        RECT 14.400 702.600 15.600 704.400 ;
        RECT 82.950 704.400 130.050 705.600 ;
        RECT 82.950 703.950 85.050 704.400 ;
        RECT 97.950 703.950 100.050 704.400 ;
        RECT 127.950 703.950 130.050 704.400 ;
        RECT 136.950 705.600 139.050 706.050 ;
        RECT 142.950 705.600 145.050 706.050 ;
        RECT 136.950 704.400 145.050 705.600 ;
        RECT 136.950 703.950 139.050 704.400 ;
        RECT 142.950 703.950 145.050 704.400 ;
        RECT 208.950 705.600 211.050 706.050 ;
        RECT 217.950 705.600 220.050 706.050 ;
        RECT 208.950 704.400 220.050 705.600 ;
        RECT 208.950 703.950 211.050 704.400 ;
        RECT 217.950 703.950 220.050 704.400 ;
        RECT 307.950 705.600 310.050 706.050 ;
        RECT 319.950 705.600 322.050 706.050 ;
        RECT 307.950 704.400 322.050 705.600 ;
        RECT 307.950 703.950 310.050 704.400 ;
        RECT 319.950 703.950 322.050 704.400 ;
        RECT 334.950 705.600 337.050 706.050 ;
        RECT 370.950 705.600 373.050 706.050 ;
        RECT 334.950 704.400 373.050 705.600 ;
        RECT 334.950 703.950 337.050 704.400 ;
        RECT 370.950 703.950 373.050 704.400 ;
        RECT 379.950 705.600 382.050 706.050 ;
        RECT 391.950 705.600 394.050 706.050 ;
        RECT 418.950 705.600 421.050 706.050 ;
        RECT 427.950 705.600 430.050 706.050 ;
        RECT 379.950 704.400 390.600 705.600 ;
        RECT 379.950 703.950 382.050 704.400 ;
        RECT 94.950 702.600 97.050 703.050 ;
        RECT 14.400 701.400 97.050 702.600 ;
        RECT 8.400 696.600 9.600 701.400 ;
        RECT 10.950 700.950 13.050 701.400 ;
        RECT 94.950 700.950 97.050 701.400 ;
        RECT 118.950 702.600 121.050 703.050 ;
        RECT 124.950 702.600 127.050 703.050 ;
        RECT 166.950 702.600 169.050 703.050 ;
        RECT 118.950 701.400 169.050 702.600 ;
        RECT 118.950 700.950 121.050 701.400 ;
        RECT 124.950 700.950 127.050 701.400 ;
        RECT 166.950 700.950 169.050 701.400 ;
        RECT 226.950 702.600 229.050 703.050 ;
        RECT 268.950 702.600 271.050 703.050 ;
        RECT 226.950 701.400 271.050 702.600 ;
        RECT 226.950 700.950 229.050 701.400 ;
        RECT 268.950 700.950 271.050 701.400 ;
        RECT 271.950 702.600 274.050 703.050 ;
        RECT 280.950 702.600 283.050 703.050 ;
        RECT 322.950 702.600 325.050 703.050 ;
        RECT 328.950 702.600 331.050 703.050 ;
        RECT 343.950 702.600 346.050 703.050 ;
        RECT 271.950 701.400 346.050 702.600 ;
        RECT 389.400 702.600 390.600 704.400 ;
        RECT 391.950 704.400 421.050 705.600 ;
        RECT 391.950 703.950 394.050 704.400 ;
        RECT 418.950 703.950 421.050 704.400 ;
        RECT 425.400 704.400 430.050 705.600 ;
        RECT 391.950 702.600 394.050 703.050 ;
        RECT 389.400 701.400 394.050 702.600 ;
        RECT 271.950 700.950 274.050 701.400 ;
        RECT 280.950 700.950 283.050 701.400 ;
        RECT 322.950 700.950 325.050 701.400 ;
        RECT 328.950 700.950 331.050 701.400 ;
        RECT 343.950 700.950 346.050 701.400 ;
        RECT 391.950 700.950 394.050 701.400 ;
        RECT 394.950 702.600 397.050 703.050 ;
        RECT 400.950 702.600 403.050 703.050 ;
        RECT 394.950 701.400 403.050 702.600 ;
        RECT 394.950 700.950 397.050 701.400 ;
        RECT 400.950 700.950 403.050 701.400 ;
        RECT 409.950 702.600 412.050 703.050 ;
        RECT 415.950 702.600 418.050 703.050 ;
        RECT 409.950 701.400 418.050 702.600 ;
        RECT 409.950 700.950 412.050 701.400 ;
        RECT 415.950 700.950 418.050 701.400 ;
        RECT 127.950 699.600 130.050 700.050 ;
        RECT 136.950 699.600 139.050 700.050 ;
        RECT 127.950 698.400 139.050 699.600 ;
        RECT 127.950 697.950 130.050 698.400 ;
        RECT 136.950 697.950 139.050 698.400 ;
        RECT 145.950 699.600 148.050 700.050 ;
        RECT 160.950 699.600 163.050 700.050 ;
        RECT 145.950 698.400 163.050 699.600 ;
        RECT 145.950 697.950 148.050 698.400 ;
        RECT 160.950 697.950 163.050 698.400 ;
        RECT 163.950 699.600 166.050 700.050 ;
        RECT 175.950 699.600 178.050 700.050 ;
        RECT 163.950 698.400 178.050 699.600 ;
        RECT 163.950 697.950 166.050 698.400 ;
        RECT 175.950 697.950 178.050 698.400 ;
        RECT 181.950 699.600 184.050 700.050 ;
        RECT 196.950 699.600 199.050 700.050 ;
        RECT 181.950 698.400 199.050 699.600 ;
        RECT 181.950 697.950 184.050 698.400 ;
        RECT 196.950 697.950 199.050 698.400 ;
        RECT 217.950 699.600 220.050 700.050 ;
        RECT 238.950 699.600 241.050 700.050 ;
        RECT 217.950 698.400 241.050 699.600 ;
        RECT 217.950 697.950 220.050 698.400 ;
        RECT 238.950 697.950 241.050 698.400 ;
        RECT 304.950 699.600 307.050 700.050 ;
        RECT 310.950 699.600 313.050 700.050 ;
        RECT 304.950 698.400 313.050 699.600 ;
        RECT 304.950 697.950 307.050 698.400 ;
        RECT 310.950 697.950 313.050 698.400 ;
        RECT 349.950 699.600 352.050 700.050 ;
        RECT 364.950 699.600 367.050 700.050 ;
        RECT 349.950 698.400 367.050 699.600 ;
        RECT 349.950 697.950 352.050 698.400 ;
        RECT 364.950 697.950 367.050 698.400 ;
        RECT 382.950 699.600 385.050 700.050 ;
        RECT 412.950 699.600 415.050 700.050 ;
        RECT 382.950 698.400 415.050 699.600 ;
        RECT 425.400 699.600 426.600 704.400 ;
        RECT 427.950 703.950 430.050 704.400 ;
        RECT 442.950 703.950 445.050 706.050 ;
        RECT 457.950 705.600 460.050 706.050 ;
        RECT 460.950 705.600 463.050 706.050 ;
        RECT 469.950 705.600 472.050 706.050 ;
        RECT 457.950 704.400 472.050 705.600 ;
        RECT 457.950 703.950 460.050 704.400 ;
        RECT 460.950 703.950 463.050 704.400 ;
        RECT 469.950 703.950 472.050 704.400 ;
        RECT 487.950 705.600 490.050 706.050 ;
        RECT 493.950 705.600 496.050 706.050 ;
        RECT 487.950 704.400 496.050 705.600 ;
        RECT 487.950 703.950 490.050 704.400 ;
        RECT 493.950 703.950 496.050 704.400 ;
        RECT 427.950 702.600 430.050 703.050 ;
        RECT 439.950 702.600 442.050 703.050 ;
        RECT 427.950 701.400 442.050 702.600 ;
        RECT 427.950 700.950 430.050 701.400 ;
        RECT 439.950 700.950 442.050 701.400 ;
        RECT 443.400 702.600 444.600 703.950 ;
        RECT 512.400 703.050 513.600 707.400 ;
        RECT 541.950 706.950 544.050 709.050 ;
        RECT 544.950 708.600 547.050 709.050 ;
        RECT 574.950 708.600 577.050 709.050 ;
        RECT 583.950 708.600 586.050 709.050 ;
        RECT 544.950 707.400 586.050 708.600 ;
        RECT 544.950 706.950 547.050 707.400 ;
        RECT 542.400 705.600 543.600 706.950 ;
        RECT 547.950 705.600 550.050 706.050 ;
        RECT 542.400 704.400 550.050 705.600 ;
        RECT 547.950 703.950 550.050 704.400 ;
        RECT 454.950 702.600 457.050 703.050 ;
        RECT 443.400 701.400 457.050 702.600 ;
        RECT 443.400 700.050 444.600 701.400 ;
        RECT 454.950 700.950 457.050 701.400 ;
        RECT 511.950 700.950 514.050 703.050 ;
        RECT 535.950 702.600 538.050 703.050 ;
        RECT 550.950 702.600 553.050 703.050 ;
        RECT 515.400 701.400 553.050 702.600 ;
        RECT 436.950 699.600 439.050 700.050 ;
        RECT 425.400 698.400 439.050 699.600 ;
        RECT 382.950 697.950 385.050 698.400 ;
        RECT 412.950 697.950 415.050 698.400 ;
        RECT 436.950 697.950 439.050 698.400 ;
        RECT 442.950 697.950 445.050 700.050 ;
        RECT 445.950 699.600 448.050 700.050 ;
        RECT 478.950 699.600 481.050 700.050 ;
        RECT 484.950 699.600 487.050 700.050 ;
        RECT 445.950 698.400 487.050 699.600 ;
        RECT 445.950 697.950 448.050 698.400 ;
        RECT 478.950 697.950 481.050 698.400 ;
        RECT 484.950 697.950 487.050 698.400 ;
        RECT 508.950 699.600 511.050 700.050 ;
        RECT 515.400 699.600 516.600 701.400 ;
        RECT 535.950 700.950 538.050 701.400 ;
        RECT 550.950 700.950 553.050 701.400 ;
        RECT 556.950 702.600 559.050 703.050 ;
        RECT 560.400 702.600 561.600 707.400 ;
        RECT 574.950 706.950 577.050 707.400 ;
        RECT 583.950 706.950 586.050 707.400 ;
        RECT 589.950 708.600 592.050 709.050 ;
        RECT 595.950 708.600 598.050 709.050 ;
        RECT 589.950 707.400 598.050 708.600 ;
        RECT 589.950 706.950 592.050 707.400 ;
        RECT 595.950 706.950 598.050 707.400 ;
        RECT 607.950 708.600 610.050 709.050 ;
        RECT 673.950 708.600 676.050 709.050 ;
        RECT 685.950 708.600 688.050 709.050 ;
        RECT 607.950 707.400 688.050 708.600 ;
        RECT 607.950 706.950 610.050 707.400 ;
        RECT 673.950 706.950 676.050 707.400 ;
        RECT 685.950 706.950 688.050 707.400 ;
        RECT 748.950 708.600 751.050 709.050 ;
        RECT 769.950 708.600 772.050 709.050 ;
        RECT 748.950 707.400 772.050 708.600 ;
        RECT 748.950 706.950 751.050 707.400 ;
        RECT 769.950 706.950 772.050 707.400 ;
        RECT 784.950 708.600 787.050 709.050 ;
        RECT 790.950 708.600 793.050 709.050 ;
        RECT 784.950 707.400 793.050 708.600 ;
        RECT 784.950 706.950 787.050 707.400 ;
        RECT 790.950 706.950 793.050 707.400 ;
        RECT 814.950 708.600 817.050 709.050 ;
        RECT 829.950 708.600 832.050 709.050 ;
        RECT 814.950 707.400 832.050 708.600 ;
        RECT 814.950 706.950 817.050 707.400 ;
        RECT 829.950 706.950 832.050 707.400 ;
        RECT 562.950 703.950 565.050 706.050 ;
        RECT 586.950 705.600 589.050 706.050 ;
        RECT 601.950 705.600 604.050 706.050 ;
        RECT 586.950 704.400 604.050 705.600 ;
        RECT 586.950 703.950 589.050 704.400 ;
        RECT 601.950 703.950 604.050 704.400 ;
        RECT 604.950 705.600 607.050 706.050 ;
        RECT 616.950 705.600 619.050 706.050 ;
        RECT 646.950 705.600 649.050 706.050 ;
        RECT 604.950 704.400 619.050 705.600 ;
        RECT 604.950 703.950 607.050 704.400 ;
        RECT 616.950 703.950 619.050 704.400 ;
        RECT 623.400 704.400 649.050 705.600 ;
        RECT 556.950 701.400 561.600 702.600 ;
        RECT 563.400 702.600 564.600 703.950 ;
        RECT 623.400 703.050 624.600 704.400 ;
        RECT 646.950 703.950 649.050 704.400 ;
        RECT 667.950 705.600 670.050 706.050 ;
        RECT 676.950 705.600 679.050 706.050 ;
        RECT 667.950 704.400 679.050 705.600 ;
        RECT 667.950 703.950 670.050 704.400 ;
        RECT 676.950 703.950 679.050 704.400 ;
        RECT 679.950 705.600 682.050 706.050 ;
        RECT 700.950 705.600 703.050 706.050 ;
        RECT 679.950 704.400 703.050 705.600 ;
        RECT 679.950 703.950 682.050 704.400 ;
        RECT 700.950 703.950 703.050 704.400 ;
        RECT 724.950 705.600 727.050 706.050 ;
        RECT 736.950 705.600 739.050 706.050 ;
        RECT 739.950 705.600 742.050 706.050 ;
        RECT 724.950 704.400 742.050 705.600 ;
        RECT 724.950 703.950 727.050 704.400 ;
        RECT 736.950 703.950 739.050 704.400 ;
        RECT 739.950 703.950 742.050 704.400 ;
        RECT 742.950 705.600 745.050 706.050 ;
        RECT 751.950 705.600 754.050 706.050 ;
        RECT 742.950 704.400 754.050 705.600 ;
        RECT 742.950 703.950 745.050 704.400 ;
        RECT 751.950 703.950 754.050 704.400 ;
        RECT 571.950 702.600 574.050 703.050 ;
        RECT 563.400 701.400 574.050 702.600 ;
        RECT 556.950 700.950 559.050 701.400 ;
        RECT 571.950 700.950 574.050 701.400 ;
        RECT 598.950 702.600 601.050 703.050 ;
        RECT 607.950 702.600 610.050 703.050 ;
        RECT 598.950 701.400 610.050 702.600 ;
        RECT 598.950 700.950 601.050 701.400 ;
        RECT 607.950 700.950 610.050 701.400 ;
        RECT 622.950 700.950 625.050 703.050 ;
        RECT 628.950 702.600 631.050 703.050 ;
        RECT 634.950 702.600 637.050 703.050 ;
        RECT 628.950 701.400 637.050 702.600 ;
        RECT 628.950 700.950 631.050 701.400 ;
        RECT 634.950 700.950 637.050 701.400 ;
        RECT 673.950 702.600 676.050 703.050 ;
        RECT 694.950 702.600 697.050 703.050 ;
        RECT 715.950 702.600 718.050 703.050 ;
        RECT 743.400 702.600 744.600 703.950 ;
        RECT 673.950 701.400 697.050 702.600 ;
        RECT 673.950 700.950 676.050 701.400 ;
        RECT 694.950 700.950 697.050 701.400 ;
        RECT 704.400 701.400 718.050 702.600 ;
        RECT 704.400 700.050 705.600 701.400 ;
        RECT 715.950 700.950 718.050 701.400 ;
        RECT 722.400 701.400 744.600 702.600 ;
        RECT 751.950 702.600 754.050 703.050 ;
        RECT 757.950 702.600 760.050 703.050 ;
        RECT 751.950 701.400 760.050 702.600 ;
        RECT 722.400 700.050 723.600 701.400 ;
        RECT 751.950 700.950 754.050 701.400 ;
        RECT 757.950 700.950 760.050 701.400 ;
        RECT 772.950 702.600 775.050 703.050 ;
        RECT 841.950 702.600 844.050 703.050 ;
        RECT 772.950 701.400 844.050 702.600 ;
        RECT 772.950 700.950 775.050 701.400 ;
        RECT 841.950 700.950 844.050 701.400 ;
        RECT 847.950 702.600 850.050 703.050 ;
        RECT 862.950 702.600 865.050 703.050 ;
        RECT 847.950 701.400 865.050 702.600 ;
        RECT 847.950 700.950 850.050 701.400 ;
        RECT 862.950 700.950 865.050 701.400 ;
        RECT 517.950 699.600 520.050 700.050 ;
        RECT 508.950 698.400 520.050 699.600 ;
        RECT 508.950 697.950 511.050 698.400 ;
        RECT 517.950 697.950 520.050 698.400 ;
        RECT 529.950 699.600 532.050 700.050 ;
        RECT 544.950 699.600 547.050 700.050 ;
        RECT 529.950 698.400 547.050 699.600 ;
        RECT 529.950 697.950 532.050 698.400 ;
        RECT 544.950 697.950 547.050 698.400 ;
        RECT 553.950 699.600 556.050 700.050 ;
        RECT 592.950 699.600 595.050 700.050 ;
        RECT 655.950 699.600 658.050 700.050 ;
        RECT 553.950 698.400 658.050 699.600 ;
        RECT 553.950 697.950 556.050 698.400 ;
        RECT 592.950 697.950 595.050 698.400 ;
        RECT 655.950 697.950 658.050 698.400 ;
        RECT 664.950 699.600 667.050 700.050 ;
        RECT 703.950 699.600 706.050 700.050 ;
        RECT 664.950 698.400 706.050 699.600 ;
        RECT 664.950 697.950 667.050 698.400 ;
        RECT 703.950 697.950 706.050 698.400 ;
        RECT 721.950 697.950 724.050 700.050 ;
        RECT 745.950 699.600 748.050 700.050 ;
        RECT 754.950 699.600 757.050 700.050 ;
        RECT 745.950 698.400 757.050 699.600 ;
        RECT 745.950 697.950 748.050 698.400 ;
        RECT 754.950 697.950 757.050 698.400 ;
        RECT 760.950 699.600 763.050 700.050 ;
        RECT 778.950 699.600 781.050 700.050 ;
        RECT 760.950 698.400 781.050 699.600 ;
        RECT 760.950 697.950 763.050 698.400 ;
        RECT 778.950 697.950 781.050 698.400 ;
        RECT 19.950 696.600 22.050 697.050 ;
        RECT 8.400 695.400 22.050 696.600 ;
        RECT 19.950 694.950 22.050 695.400 ;
        RECT 22.950 696.600 25.050 697.050 ;
        RECT 58.950 696.600 61.050 697.050 ;
        RECT 22.950 695.400 61.050 696.600 ;
        RECT 22.950 694.950 25.050 695.400 ;
        RECT 58.950 694.950 61.050 695.400 ;
        RECT 133.950 696.600 136.050 697.050 ;
        RECT 184.950 696.600 187.050 697.050 ;
        RECT 133.950 695.400 187.050 696.600 ;
        RECT 133.950 694.950 136.050 695.400 ;
        RECT 184.950 694.950 187.050 695.400 ;
        RECT 220.950 696.600 223.050 697.050 ;
        RECT 319.950 696.600 322.050 697.050 ;
        RECT 331.950 696.600 334.050 697.050 ;
        RECT 340.950 696.600 343.050 697.050 ;
        RECT 358.950 696.600 361.050 697.050 ;
        RECT 382.950 696.600 385.050 697.050 ;
        RECT 220.950 695.400 385.050 696.600 ;
        RECT 220.950 694.950 223.050 695.400 ;
        RECT 319.950 694.950 322.050 695.400 ;
        RECT 331.950 694.950 334.050 695.400 ;
        RECT 340.950 694.950 343.050 695.400 ;
        RECT 358.950 694.950 361.050 695.400 ;
        RECT 382.950 694.950 385.050 695.400 ;
        RECT 385.950 696.600 388.050 697.050 ;
        RECT 499.950 696.600 502.050 697.050 ;
        RECT 385.950 695.400 502.050 696.600 ;
        RECT 385.950 694.950 388.050 695.400 ;
        RECT 499.950 694.950 502.050 695.400 ;
        RECT 535.950 696.600 538.050 697.050 ;
        RECT 571.950 696.600 574.050 697.050 ;
        RECT 580.950 696.600 583.050 697.050 ;
        RECT 535.950 695.400 583.050 696.600 ;
        RECT 535.950 694.950 538.050 695.400 ;
        RECT 571.950 694.950 574.050 695.400 ;
        RECT 580.950 694.950 583.050 695.400 ;
        RECT 595.950 696.600 598.050 697.050 ;
        RECT 604.950 696.600 607.050 697.050 ;
        RECT 595.950 695.400 607.050 696.600 ;
        RECT 595.950 694.950 598.050 695.400 ;
        RECT 604.950 694.950 607.050 695.400 ;
        RECT 619.950 696.600 622.050 697.050 ;
        RECT 628.950 696.600 631.050 697.050 ;
        RECT 619.950 695.400 631.050 696.600 ;
        RECT 619.950 694.950 622.050 695.400 ;
        RECT 628.950 694.950 631.050 695.400 ;
        RECT 649.950 696.600 652.050 697.050 ;
        RECT 688.950 696.600 691.050 697.050 ;
        RECT 649.950 695.400 691.050 696.600 ;
        RECT 649.950 694.950 652.050 695.400 ;
        RECT 688.950 694.950 691.050 695.400 ;
        RECT 724.950 696.600 727.050 697.050 ;
        RECT 730.950 696.600 733.050 697.050 ;
        RECT 724.950 695.400 733.050 696.600 ;
        RECT 724.950 694.950 727.050 695.400 ;
        RECT 730.950 694.950 733.050 695.400 ;
        RECT 763.950 696.600 766.050 697.050 ;
        RECT 772.950 696.600 775.050 697.050 ;
        RECT 763.950 695.400 775.050 696.600 ;
        RECT 763.950 694.950 766.050 695.400 ;
        RECT 772.950 694.950 775.050 695.400 ;
        RECT 844.950 696.600 847.050 697.050 ;
        RECT 850.950 696.600 853.050 697.050 ;
        RECT 844.950 695.400 853.050 696.600 ;
        RECT 844.950 694.950 847.050 695.400 ;
        RECT 850.950 694.950 853.050 695.400 ;
        RECT 238.950 693.600 241.050 694.050 ;
        RECT 262.950 693.600 265.050 694.050 ;
        RECT 238.950 692.400 265.050 693.600 ;
        RECT 238.950 691.950 241.050 692.400 ;
        RECT 262.950 691.950 265.050 692.400 ;
        RECT 334.950 693.600 337.050 694.050 ;
        RECT 349.950 693.600 352.050 694.050 ;
        RECT 334.950 692.400 352.050 693.600 ;
        RECT 334.950 691.950 337.050 692.400 ;
        RECT 349.950 691.950 352.050 692.400 ;
        RECT 352.950 693.600 355.050 694.050 ;
        RECT 388.950 693.600 391.050 694.050 ;
        RECT 352.950 692.400 391.050 693.600 ;
        RECT 352.950 691.950 355.050 692.400 ;
        RECT 388.950 691.950 391.050 692.400 ;
        RECT 415.950 693.600 418.050 694.050 ;
        RECT 424.950 693.600 427.050 694.050 ;
        RECT 415.950 692.400 427.050 693.600 ;
        RECT 415.950 691.950 418.050 692.400 ;
        RECT 424.950 691.950 427.050 692.400 ;
        RECT 448.950 693.600 451.050 694.050 ;
        RECT 466.950 693.600 469.050 694.050 ;
        RECT 493.950 693.600 496.050 694.050 ;
        RECT 505.950 693.600 508.050 694.050 ;
        RECT 448.950 692.400 508.050 693.600 ;
        RECT 448.950 691.950 451.050 692.400 ;
        RECT 466.950 691.950 469.050 692.400 ;
        RECT 493.950 691.950 496.050 692.400 ;
        RECT 505.950 691.950 508.050 692.400 ;
        RECT 523.950 693.600 526.050 694.050 ;
        RECT 556.950 693.600 559.050 694.050 ;
        RECT 523.950 692.400 559.050 693.600 ;
        RECT 523.950 691.950 526.050 692.400 ;
        RECT 556.950 691.950 559.050 692.400 ;
        RECT 565.950 693.600 568.050 694.050 ;
        RECT 589.950 693.600 592.050 694.050 ;
        RECT 565.950 692.400 592.050 693.600 ;
        RECT 565.950 691.950 568.050 692.400 ;
        RECT 589.950 691.950 592.050 692.400 ;
        RECT 664.950 693.600 667.050 694.050 ;
        RECT 697.950 693.600 700.050 694.050 ;
        RECT 751.950 693.600 754.050 694.050 ;
        RECT 664.950 692.400 754.050 693.600 ;
        RECT 664.950 691.950 667.050 692.400 ;
        RECT 697.950 691.950 700.050 692.400 ;
        RECT 751.950 691.950 754.050 692.400 ;
        RECT 760.950 693.600 763.050 694.050 ;
        RECT 766.950 693.600 769.050 694.050 ;
        RECT 760.950 692.400 769.050 693.600 ;
        RECT 760.950 691.950 763.050 692.400 ;
        RECT 766.950 691.950 769.050 692.400 ;
        RECT 85.950 690.600 88.050 691.050 ;
        RECT 226.950 690.600 229.050 691.050 ;
        RECT 85.950 689.400 229.050 690.600 ;
        RECT 85.950 688.950 88.050 689.400 ;
        RECT 226.950 688.950 229.050 689.400 ;
        RECT 235.950 690.600 238.050 691.050 ;
        RECT 241.950 690.600 244.050 691.050 ;
        RECT 235.950 689.400 244.050 690.600 ;
        RECT 235.950 688.950 238.050 689.400 ;
        RECT 241.950 688.950 244.050 689.400 ;
        RECT 289.950 690.600 292.050 691.050 ;
        RECT 406.950 690.600 409.050 691.050 ;
        RECT 289.950 689.400 409.050 690.600 ;
        RECT 289.950 688.950 292.050 689.400 ;
        RECT 406.950 688.950 409.050 689.400 ;
        RECT 430.950 690.600 433.050 691.050 ;
        RECT 472.950 690.600 475.050 691.050 ;
        RECT 430.950 689.400 475.050 690.600 ;
        RECT 430.950 688.950 433.050 689.400 ;
        RECT 472.950 688.950 475.050 689.400 ;
        RECT 508.950 690.600 511.050 691.050 ;
        RECT 532.950 690.600 535.050 691.050 ;
        RECT 508.950 689.400 535.050 690.600 ;
        RECT 508.950 688.950 511.050 689.400 ;
        RECT 532.950 688.950 535.050 689.400 ;
        RECT 766.950 690.600 769.050 691.050 ;
        RECT 784.950 690.600 787.050 691.050 ;
        RECT 766.950 689.400 787.050 690.600 ;
        RECT 766.950 688.950 769.050 689.400 ;
        RECT 784.950 688.950 787.050 689.400 ;
        RECT 811.950 690.600 814.050 691.050 ;
        RECT 820.950 690.600 823.050 691.050 ;
        RECT 811.950 689.400 823.050 690.600 ;
        RECT 811.950 688.950 814.050 689.400 ;
        RECT 820.950 688.950 823.050 689.400 ;
        RECT 190.950 687.600 193.050 688.050 ;
        RECT 325.950 687.600 328.050 688.050 ;
        RECT 190.950 686.400 328.050 687.600 ;
        RECT 190.950 685.950 193.050 686.400 ;
        RECT 325.950 685.950 328.050 686.400 ;
        RECT 346.950 687.600 349.050 688.050 ;
        RECT 367.950 687.600 370.050 688.050 ;
        RECT 346.950 686.400 370.050 687.600 ;
        RECT 346.950 685.950 349.050 686.400 ;
        RECT 367.950 685.950 370.050 686.400 ;
        RECT 415.950 687.600 418.050 688.050 ;
        RECT 433.950 687.600 436.050 688.050 ;
        RECT 415.950 686.400 436.050 687.600 ;
        RECT 415.950 685.950 418.050 686.400 ;
        RECT 433.950 685.950 436.050 686.400 ;
        RECT 475.950 687.600 478.050 688.050 ;
        RECT 505.950 687.600 508.050 688.050 ;
        RECT 475.950 686.400 508.050 687.600 ;
        RECT 475.950 685.950 478.050 686.400 ;
        RECT 505.950 685.950 508.050 686.400 ;
        RECT 511.950 687.600 514.050 688.050 ;
        RECT 598.950 687.600 601.050 688.050 ;
        RECT 613.950 687.600 616.050 688.050 ;
        RECT 511.950 686.400 616.050 687.600 ;
        RECT 511.950 685.950 514.050 686.400 ;
        RECT 598.950 685.950 601.050 686.400 ;
        RECT 613.950 685.950 616.050 686.400 ;
        RECT 763.950 687.600 766.050 688.050 ;
        RECT 832.950 687.600 835.050 688.050 ;
        RECT 763.950 686.400 835.050 687.600 ;
        RECT 763.950 685.950 766.050 686.400 ;
        RECT 832.950 685.950 835.050 686.400 ;
        RECT 166.950 684.600 169.050 685.050 ;
        RECT 238.950 684.600 241.050 685.050 ;
        RECT 166.950 683.400 241.050 684.600 ;
        RECT 166.950 682.950 169.050 683.400 ;
        RECT 238.950 682.950 241.050 683.400 ;
        RECT 331.950 684.600 334.050 685.050 ;
        RECT 361.950 684.600 364.050 685.050 ;
        RECT 331.950 683.400 364.050 684.600 ;
        RECT 331.950 682.950 334.050 683.400 ;
        RECT 361.950 682.950 364.050 683.400 ;
        RECT 412.950 684.600 415.050 685.050 ;
        RECT 439.950 684.600 442.050 685.050 ;
        RECT 412.950 683.400 442.050 684.600 ;
        RECT 412.950 682.950 415.050 683.400 ;
        RECT 439.950 682.950 442.050 683.400 ;
        RECT 460.950 684.600 463.050 685.050 ;
        RECT 493.950 684.600 496.050 685.050 ;
        RECT 460.950 683.400 496.050 684.600 ;
        RECT 460.950 682.950 463.050 683.400 ;
        RECT 493.950 682.950 496.050 683.400 ;
        RECT 502.950 684.600 505.050 685.050 ;
        RECT 538.950 684.600 541.050 685.050 ;
        RECT 502.950 683.400 541.050 684.600 ;
        RECT 502.950 682.950 505.050 683.400 ;
        RECT 538.950 682.950 541.050 683.400 ;
        RECT 580.950 684.600 583.050 685.050 ;
        RECT 625.950 684.600 628.050 685.050 ;
        RECT 580.950 683.400 628.050 684.600 ;
        RECT 580.950 682.950 583.050 683.400 ;
        RECT 625.950 682.950 628.050 683.400 ;
        RECT 682.950 684.600 685.050 685.050 ;
        RECT 691.950 684.600 694.050 685.050 ;
        RECT 682.950 683.400 694.050 684.600 ;
        RECT 682.950 682.950 685.050 683.400 ;
        RECT 691.950 682.950 694.050 683.400 ;
        RECT 256.950 681.600 259.050 682.050 ;
        RECT 355.950 681.600 358.050 682.050 ;
        RECT 256.950 680.400 358.050 681.600 ;
        RECT 256.950 679.950 259.050 680.400 ;
        RECT 355.950 679.950 358.050 680.400 ;
        RECT 409.950 681.600 412.050 682.050 ;
        RECT 466.950 681.600 469.050 682.050 ;
        RECT 409.950 680.400 469.050 681.600 ;
        RECT 409.950 679.950 412.050 680.400 ;
        RECT 466.950 679.950 469.050 680.400 ;
        RECT 478.950 681.600 481.050 682.050 ;
        RECT 523.950 681.600 526.050 682.050 ;
        RECT 478.950 680.400 526.050 681.600 ;
        RECT 478.950 679.950 481.050 680.400 ;
        RECT 523.950 679.950 526.050 680.400 ;
        RECT 583.950 681.600 586.050 682.050 ;
        RECT 616.950 681.600 619.050 682.050 ;
        RECT 646.950 681.600 649.050 682.050 ;
        RECT 583.950 680.400 649.050 681.600 ;
        RECT 583.950 679.950 586.050 680.400 ;
        RECT 616.950 679.950 619.050 680.400 ;
        RECT 646.950 679.950 649.050 680.400 ;
        RECT 112.950 678.600 115.050 679.050 ;
        RECT 157.950 678.600 160.050 679.050 ;
        RECT 169.950 678.600 172.050 679.050 ;
        RECT 112.950 677.400 172.050 678.600 ;
        RECT 112.950 676.950 115.050 677.400 ;
        RECT 157.950 676.950 160.050 677.400 ;
        RECT 169.950 676.950 172.050 677.400 ;
        RECT 247.950 678.600 250.050 679.050 ;
        RECT 271.950 678.600 274.050 679.050 ;
        RECT 247.950 677.400 274.050 678.600 ;
        RECT 247.950 676.950 250.050 677.400 ;
        RECT 271.950 676.950 274.050 677.400 ;
        RECT 304.950 678.600 307.050 679.050 ;
        RECT 313.950 678.600 316.050 679.050 ;
        RECT 304.950 677.400 316.050 678.600 ;
        RECT 304.950 676.950 307.050 677.400 ;
        RECT 313.950 676.950 316.050 677.400 ;
        RECT 346.950 678.600 349.050 679.050 ;
        RECT 388.950 678.600 391.050 679.050 ;
        RECT 346.950 677.400 391.050 678.600 ;
        RECT 346.950 676.950 349.050 677.400 ;
        RECT 388.950 676.950 391.050 677.400 ;
        RECT 391.950 678.600 394.050 679.050 ;
        RECT 403.950 678.600 406.050 679.050 ;
        RECT 430.950 678.600 433.050 679.050 ;
        RECT 391.950 677.400 433.050 678.600 ;
        RECT 391.950 676.950 394.050 677.400 ;
        RECT 403.950 676.950 406.050 677.400 ;
        RECT 430.950 676.950 433.050 677.400 ;
        RECT 439.950 678.600 442.050 679.050 ;
        RECT 445.950 678.600 448.050 679.050 ;
        RECT 439.950 677.400 448.050 678.600 ;
        RECT 439.950 676.950 442.050 677.400 ;
        RECT 445.950 676.950 448.050 677.400 ;
        RECT 451.950 678.600 454.050 679.050 ;
        RECT 472.950 678.600 475.050 679.050 ;
        RECT 451.950 677.400 475.050 678.600 ;
        RECT 451.950 676.950 454.050 677.400 ;
        RECT 472.950 676.950 475.050 677.400 ;
        RECT 481.950 678.600 484.050 679.050 ;
        RECT 514.950 678.600 517.050 679.050 ;
        RECT 481.950 677.400 517.050 678.600 ;
        RECT 481.950 676.950 484.050 677.400 ;
        RECT 514.950 676.950 517.050 677.400 ;
        RECT 535.950 678.600 538.050 679.050 ;
        RECT 556.950 678.600 559.050 679.050 ;
        RECT 535.950 677.400 559.050 678.600 ;
        RECT 535.950 676.950 538.050 677.400 ;
        RECT 556.950 676.950 559.050 677.400 ;
        RECT 562.950 678.600 565.050 679.050 ;
        RECT 574.950 678.600 577.050 679.050 ;
        RECT 610.950 678.600 613.050 679.050 ;
        RECT 562.950 677.400 613.050 678.600 ;
        RECT 562.950 676.950 565.050 677.400 ;
        RECT 574.950 676.950 577.050 677.400 ;
        RECT 610.950 676.950 613.050 677.400 ;
        RECT 754.950 678.600 757.050 679.050 ;
        RECT 769.950 678.600 772.050 679.050 ;
        RECT 784.950 678.600 787.050 679.050 ;
        RECT 754.950 677.400 787.050 678.600 ;
        RECT 754.950 676.950 757.050 677.400 ;
        RECT 769.950 676.950 772.050 677.400 ;
        RECT 784.950 676.950 787.050 677.400 ;
        RECT 28.950 675.600 31.050 676.050 ;
        RECT 127.950 675.600 130.050 676.050 ;
        RECT 28.950 674.400 130.050 675.600 ;
        RECT 28.950 673.950 31.050 674.400 ;
        RECT 127.950 673.950 130.050 674.400 ;
        RECT 160.950 675.600 163.050 676.050 ;
        RECT 169.950 675.600 172.050 676.050 ;
        RECT 160.950 674.400 172.050 675.600 ;
        RECT 160.950 673.950 163.050 674.400 ;
        RECT 169.950 673.950 172.050 674.400 ;
        RECT 181.950 675.600 184.050 676.050 ;
        RECT 193.950 675.600 196.050 676.050 ;
        RECT 181.950 674.400 196.050 675.600 ;
        RECT 181.950 673.950 184.050 674.400 ;
        RECT 193.950 673.950 196.050 674.400 ;
        RECT 217.950 675.600 220.050 676.050 ;
        RECT 232.950 675.600 235.050 676.050 ;
        RECT 241.950 675.600 244.050 676.050 ;
        RECT 298.950 675.600 301.050 676.050 ;
        RECT 217.950 674.400 301.050 675.600 ;
        RECT 217.950 673.950 220.050 674.400 ;
        RECT 232.950 673.950 235.050 674.400 ;
        RECT 241.950 673.950 244.050 674.400 ;
        RECT 298.950 673.950 301.050 674.400 ;
        RECT 307.950 673.950 310.050 676.050 ;
        RECT 322.950 675.600 325.050 676.050 ;
        RECT 358.950 675.600 361.050 676.050 ;
        RECT 373.950 675.600 376.050 676.050 ;
        RECT 322.950 674.400 376.050 675.600 ;
        RECT 322.950 673.950 325.050 674.400 ;
        RECT 358.950 673.950 361.050 674.400 ;
        RECT 373.950 673.950 376.050 674.400 ;
        RECT 382.950 675.600 385.050 676.050 ;
        RECT 421.950 675.600 424.050 676.050 ;
        RECT 481.950 675.600 484.050 676.050 ;
        RECT 382.950 674.400 484.050 675.600 ;
        RECT 382.950 673.950 385.050 674.400 ;
        RECT 421.950 673.950 424.050 674.400 ;
        RECT 481.950 673.950 484.050 674.400 ;
        RECT 496.950 675.600 499.050 676.050 ;
        RECT 547.950 675.600 550.050 676.050 ;
        RECT 568.950 675.600 571.050 676.050 ;
        RECT 496.950 674.400 571.050 675.600 ;
        RECT 496.950 673.950 499.050 674.400 ;
        RECT 547.950 673.950 550.050 674.400 ;
        RECT 568.950 673.950 571.050 674.400 ;
        RECT 571.950 675.600 574.050 676.050 ;
        RECT 583.950 675.600 586.050 676.050 ;
        RECT 589.950 675.600 592.050 676.050 ;
        RECT 571.950 674.400 582.600 675.600 ;
        RECT 571.950 673.950 574.050 674.400 ;
        RECT 100.950 672.600 103.050 673.050 ;
        RECT 106.950 672.600 109.050 673.050 ;
        RECT 100.950 671.400 109.050 672.600 ;
        RECT 100.950 670.950 103.050 671.400 ;
        RECT 106.950 670.950 109.050 671.400 ;
        RECT 112.950 672.600 115.050 673.050 ;
        RECT 121.950 672.600 124.050 673.050 ;
        RECT 112.950 671.400 124.050 672.600 ;
        RECT 112.950 670.950 115.050 671.400 ;
        RECT 121.950 670.950 124.050 671.400 ;
        RECT 136.950 672.600 139.050 673.050 ;
        RECT 163.950 672.600 166.050 673.050 ;
        RECT 166.950 672.600 169.050 673.050 ;
        RECT 136.950 671.400 169.050 672.600 ;
        RECT 136.950 670.950 139.050 671.400 ;
        RECT 163.950 670.950 166.050 671.400 ;
        RECT 166.950 670.950 169.050 671.400 ;
        RECT 172.950 672.600 175.050 673.050 ;
        RECT 178.950 672.600 181.050 673.050 ;
        RECT 193.950 672.600 196.050 673.050 ;
        RECT 172.950 671.400 177.600 672.600 ;
        RECT 172.950 670.950 175.050 671.400 ;
        RECT 55.950 669.600 58.050 670.050 ;
        RECT 85.950 669.600 88.050 670.050 ;
        RECT 55.950 668.400 88.050 669.600 ;
        RECT 55.950 667.950 58.050 668.400 ;
        RECT 85.950 667.950 88.050 668.400 ;
        RECT 130.950 669.600 133.050 670.050 ;
        RECT 142.950 669.600 145.050 670.050 ;
        RECT 130.950 668.400 145.050 669.600 ;
        RECT 176.400 669.600 177.600 671.400 ;
        RECT 178.950 671.400 196.050 672.600 ;
        RECT 178.950 670.950 181.050 671.400 ;
        RECT 193.950 670.950 196.050 671.400 ;
        RECT 250.950 672.600 253.050 673.050 ;
        RECT 268.950 672.600 271.050 673.050 ;
        RECT 295.950 672.600 298.050 673.050 ;
        RECT 250.950 671.400 298.050 672.600 ;
        RECT 250.950 670.950 253.050 671.400 ;
        RECT 268.950 670.950 271.050 671.400 ;
        RECT 295.950 670.950 298.050 671.400 ;
        RECT 301.950 670.950 304.050 673.050 ;
        RECT 196.950 669.600 199.050 670.050 ;
        RECT 176.400 668.400 199.050 669.600 ;
        RECT 130.950 667.950 133.050 668.400 ;
        RECT 142.950 667.950 145.050 668.400 ;
        RECT 196.950 667.950 199.050 668.400 ;
        RECT 235.950 669.600 238.050 670.050 ;
        RECT 292.950 669.600 295.050 670.050 ;
        RECT 235.950 668.400 295.050 669.600 ;
        RECT 235.950 667.950 238.050 668.400 ;
        RECT 292.950 667.950 295.050 668.400 ;
        RECT 79.950 666.600 82.050 667.050 ;
        RECT 88.950 666.600 91.050 667.050 ;
        RECT 79.950 665.400 91.050 666.600 ;
        RECT 79.950 664.950 82.050 665.400 ;
        RECT 88.950 664.950 91.050 665.400 ;
        RECT 133.950 666.600 136.050 667.050 ;
        RECT 139.950 666.600 142.050 667.050 ;
        RECT 133.950 665.400 142.050 666.600 ;
        RECT 133.950 664.950 136.050 665.400 ;
        RECT 139.950 664.950 142.050 665.400 ;
        RECT 169.950 666.600 172.050 667.050 ;
        RECT 175.950 666.600 178.050 667.050 ;
        RECT 169.950 665.400 178.050 666.600 ;
        RECT 169.950 664.950 172.050 665.400 ;
        RECT 175.950 664.950 178.050 665.400 ;
        RECT 202.950 666.600 205.050 667.050 ;
        RECT 211.950 666.600 214.050 667.050 ;
        RECT 202.950 665.400 214.050 666.600 ;
        RECT 302.400 666.600 303.600 670.950 ;
        RECT 308.400 670.050 309.600 673.950 ;
        RECT 310.950 672.600 313.050 673.050 ;
        RECT 364.950 672.600 367.050 673.050 ;
        RECT 385.950 672.600 388.050 673.050 ;
        RECT 310.950 671.400 342.600 672.600 ;
        RECT 310.950 670.950 313.050 671.400 ;
        RECT 307.950 667.950 310.050 670.050 ;
        RECT 322.950 669.600 325.050 670.050 ;
        RECT 328.950 669.600 331.050 670.050 ;
        RECT 322.950 668.400 331.050 669.600 ;
        RECT 341.400 669.600 342.600 671.400 ;
        RECT 364.950 671.400 388.050 672.600 ;
        RECT 364.950 670.950 367.050 671.400 ;
        RECT 385.950 670.950 388.050 671.400 ;
        RECT 388.950 672.600 391.050 673.050 ;
        RECT 427.950 672.600 430.050 673.050 ;
        RECT 433.950 672.600 436.050 673.050 ;
        RECT 388.950 671.400 436.050 672.600 ;
        RECT 388.950 670.950 391.050 671.400 ;
        RECT 427.950 670.950 430.050 671.400 ;
        RECT 433.950 670.950 436.050 671.400 ;
        RECT 436.950 672.600 439.050 673.050 ;
        RECT 445.950 672.600 448.050 673.050 ;
        RECT 454.950 672.600 457.050 673.050 ;
        RECT 436.950 671.400 444.600 672.600 ;
        RECT 436.950 670.950 439.050 671.400 ;
        RECT 343.950 669.600 346.050 670.050 ;
        RECT 341.400 668.400 346.050 669.600 ;
        RECT 322.950 667.950 325.050 668.400 ;
        RECT 328.950 667.950 331.050 668.400 ;
        RECT 343.950 667.950 346.050 668.400 ;
        RECT 370.950 669.600 373.050 670.050 ;
        RECT 382.950 669.600 385.050 670.050 ;
        RECT 370.950 668.400 385.050 669.600 ;
        RECT 370.950 667.950 373.050 668.400 ;
        RECT 382.950 667.950 385.050 668.400 ;
        RECT 388.950 667.950 391.050 670.050 ;
        RECT 406.950 669.600 409.050 670.050 ;
        RECT 412.950 669.600 415.050 670.050 ;
        RECT 406.950 668.400 415.050 669.600 ;
        RECT 443.400 669.600 444.600 671.400 ;
        RECT 445.950 671.400 457.050 672.600 ;
        RECT 445.950 670.950 448.050 671.400 ;
        RECT 454.950 670.950 457.050 671.400 ;
        RECT 523.950 670.950 526.050 673.050 ;
        RECT 529.950 672.600 532.050 673.050 ;
        RECT 535.950 672.600 538.050 673.050 ;
        RECT 559.950 672.600 562.050 673.050 ;
        RECT 529.950 671.400 538.050 672.600 ;
        RECT 529.950 670.950 532.050 671.400 ;
        RECT 535.950 670.950 538.050 671.400 ;
        RECT 542.400 671.400 562.050 672.600 ;
        RECT 581.400 672.600 582.600 674.400 ;
        RECT 583.950 674.400 592.050 675.600 ;
        RECT 583.950 673.950 586.050 674.400 ;
        RECT 589.950 673.950 592.050 674.400 ;
        RECT 592.950 675.600 595.050 676.050 ;
        RECT 601.950 675.600 604.050 676.050 ;
        RECT 592.950 674.400 604.050 675.600 ;
        RECT 592.950 673.950 595.050 674.400 ;
        RECT 601.950 673.950 604.050 674.400 ;
        RECT 604.950 675.600 607.050 676.050 ;
        RECT 607.950 675.600 610.050 676.050 ;
        RECT 622.950 675.600 625.050 676.050 ;
        RECT 604.950 674.400 625.050 675.600 ;
        RECT 604.950 673.950 607.050 674.400 ;
        RECT 607.950 673.950 610.050 674.400 ;
        RECT 622.950 673.950 625.050 674.400 ;
        RECT 637.950 675.600 640.050 676.050 ;
        RECT 688.950 675.600 691.050 676.050 ;
        RECT 637.950 674.400 691.050 675.600 ;
        RECT 637.950 673.950 640.050 674.400 ;
        RECT 688.950 673.950 691.050 674.400 ;
        RECT 769.950 675.600 772.050 676.050 ;
        RECT 775.950 675.600 778.050 676.050 ;
        RECT 769.950 674.400 778.050 675.600 ;
        RECT 769.950 673.950 772.050 674.400 ;
        RECT 775.950 673.950 778.050 674.400 ;
        RECT 790.950 675.600 793.050 676.050 ;
        RECT 796.950 675.600 799.050 676.050 ;
        RECT 790.950 674.400 799.050 675.600 ;
        RECT 790.950 673.950 793.050 674.400 ;
        RECT 796.950 673.950 799.050 674.400 ;
        RECT 823.950 675.600 826.050 676.050 ;
        RECT 838.950 675.600 841.050 676.050 ;
        RECT 823.950 674.400 841.050 675.600 ;
        RECT 823.950 673.950 826.050 674.400 ;
        RECT 838.950 673.950 841.050 674.400 ;
        RECT 586.950 672.600 589.050 673.050 ;
        RECT 581.400 671.400 589.050 672.600 ;
        RECT 457.950 669.600 460.050 670.050 ;
        RECT 443.400 668.400 460.050 669.600 ;
        RECT 406.950 667.950 409.050 668.400 ;
        RECT 412.950 667.950 415.050 668.400 ;
        RECT 457.950 667.950 460.050 668.400 ;
        RECT 490.950 669.600 493.050 670.050 ;
        RECT 514.950 669.600 517.050 670.050 ;
        RECT 490.950 668.400 517.050 669.600 ;
        RECT 524.400 669.600 525.600 670.950 ;
        RECT 526.950 669.600 529.050 670.050 ;
        RECT 524.400 668.400 529.050 669.600 ;
        RECT 490.950 667.950 493.050 668.400 ;
        RECT 514.950 667.950 517.050 668.400 ;
        RECT 526.950 667.950 529.050 668.400 ;
        RECT 343.950 666.600 346.050 667.050 ;
        RECT 302.400 665.400 346.050 666.600 ;
        RECT 389.400 666.600 390.600 667.950 ;
        RECT 530.400 667.050 531.600 670.950 ;
        RECT 542.400 670.050 543.600 671.400 ;
        RECT 559.950 670.950 562.050 671.400 ;
        RECT 586.950 670.950 589.050 671.400 ;
        RECT 619.950 672.600 622.050 673.050 ;
        RECT 634.950 672.600 637.050 673.050 ;
        RECT 619.950 671.400 637.050 672.600 ;
        RECT 619.950 670.950 622.050 671.400 ;
        RECT 634.950 670.950 637.050 671.400 ;
        RECT 643.950 672.600 646.050 673.050 ;
        RECT 652.950 672.600 655.050 673.050 ;
        RECT 643.950 671.400 655.050 672.600 ;
        RECT 643.950 670.950 646.050 671.400 ;
        RECT 652.950 670.950 655.050 671.400 ;
        RECT 778.950 672.600 781.050 673.050 ;
        RECT 829.950 672.600 832.050 673.050 ;
        RECT 778.950 671.400 832.050 672.600 ;
        RECT 778.950 670.950 781.050 671.400 ;
        RECT 829.950 670.950 832.050 671.400 ;
        RECT 541.950 667.950 544.050 670.050 ;
        RECT 556.950 669.600 559.050 670.050 ;
        RECT 595.950 669.600 598.050 670.050 ;
        RECT 556.950 668.400 598.050 669.600 ;
        RECT 556.950 667.950 559.050 668.400 ;
        RECT 595.950 667.950 598.050 668.400 ;
        RECT 640.950 669.600 643.050 670.050 ;
        RECT 658.950 669.600 661.050 670.050 ;
        RECT 640.950 668.400 661.050 669.600 ;
        RECT 640.950 667.950 643.050 668.400 ;
        RECT 658.950 667.950 661.050 668.400 ;
        RECT 661.950 669.600 664.050 670.050 ;
        RECT 715.950 669.600 718.050 670.050 ;
        RECT 757.950 669.600 760.050 670.050 ;
        RECT 766.950 669.600 769.050 670.050 ;
        RECT 661.950 668.400 769.050 669.600 ;
        RECT 661.950 667.950 664.050 668.400 ;
        RECT 715.950 667.950 718.050 668.400 ;
        RECT 757.950 667.950 760.050 668.400 ;
        RECT 766.950 667.950 769.050 668.400 ;
        RECT 787.950 669.600 790.050 670.050 ;
        RECT 802.950 669.600 805.050 670.050 ;
        RECT 787.950 668.400 805.050 669.600 ;
        RECT 787.950 667.950 790.050 668.400 ;
        RECT 802.950 667.950 805.050 668.400 ;
        RECT 418.950 666.600 421.050 667.050 ;
        RECT 475.950 666.600 478.050 667.050 ;
        RECT 484.950 666.600 487.050 667.050 ;
        RECT 389.400 665.400 487.050 666.600 ;
        RECT 202.950 664.950 205.050 665.400 ;
        RECT 211.950 664.950 214.050 665.400 ;
        RECT 343.950 664.950 346.050 665.400 ;
        RECT 418.950 664.950 421.050 665.400 ;
        RECT 475.950 664.950 478.050 665.400 ;
        RECT 484.950 664.950 487.050 665.400 ;
        RECT 496.950 666.600 499.050 667.050 ;
        RECT 499.950 666.600 502.050 667.050 ;
        RECT 511.950 666.600 514.050 667.050 ;
        RECT 496.950 665.400 514.050 666.600 ;
        RECT 496.950 664.950 499.050 665.400 ;
        RECT 499.950 664.950 502.050 665.400 ;
        RECT 511.950 664.950 514.050 665.400 ;
        RECT 529.950 664.950 532.050 667.050 ;
        RECT 532.950 666.600 535.050 667.050 ;
        RECT 568.950 666.600 571.050 667.050 ;
        RECT 532.950 665.400 571.050 666.600 ;
        RECT 532.950 664.950 535.050 665.400 ;
        RECT 568.950 664.950 571.050 665.400 ;
        RECT 640.950 666.600 643.050 667.050 ;
        RECT 652.950 666.600 655.050 667.050 ;
        RECT 640.950 665.400 655.050 666.600 ;
        RECT 640.950 664.950 643.050 665.400 ;
        RECT 652.950 664.950 655.050 665.400 ;
        RECT 712.950 666.600 715.050 667.050 ;
        RECT 763.950 666.600 766.050 667.050 ;
        RECT 712.950 665.400 766.050 666.600 ;
        RECT 712.950 664.950 715.050 665.400 ;
        RECT 763.950 664.950 766.050 665.400 ;
        RECT 775.950 666.600 778.050 667.050 ;
        RECT 835.950 666.600 838.050 667.050 ;
        RECT 775.950 665.400 838.050 666.600 ;
        RECT 775.950 664.950 778.050 665.400 ;
        RECT 835.950 664.950 838.050 665.400 ;
        RECT 67.950 663.600 70.050 664.050 ;
        RECT 118.950 663.600 121.050 664.050 ;
        RECT 133.950 663.600 136.050 664.050 ;
        RECT 67.950 662.400 136.050 663.600 ;
        RECT 67.950 661.950 70.050 662.400 ;
        RECT 118.950 661.950 121.050 662.400 ;
        RECT 133.950 661.950 136.050 662.400 ;
        RECT 175.950 663.600 178.050 664.050 ;
        RECT 253.950 663.600 256.050 664.050 ;
        RECT 175.950 662.400 256.050 663.600 ;
        RECT 175.950 661.950 178.050 662.400 ;
        RECT 253.950 661.950 256.050 662.400 ;
        RECT 277.950 663.600 280.050 664.050 ;
        RECT 307.950 663.600 310.050 664.050 ;
        RECT 277.950 662.400 310.050 663.600 ;
        RECT 277.950 661.950 280.050 662.400 ;
        RECT 307.950 661.950 310.050 662.400 ;
        RECT 526.950 663.600 529.050 664.050 ;
        RECT 532.950 663.600 535.050 664.050 ;
        RECT 526.950 662.400 535.050 663.600 ;
        RECT 526.950 661.950 529.050 662.400 ;
        RECT 532.950 661.950 535.050 662.400 ;
        RECT 616.950 663.600 619.050 664.050 ;
        RECT 631.950 663.600 634.050 664.050 ;
        RECT 616.950 662.400 634.050 663.600 ;
        RECT 616.950 661.950 619.050 662.400 ;
        RECT 631.950 661.950 634.050 662.400 ;
        RECT 751.950 663.600 754.050 664.050 ;
        RECT 814.950 663.600 817.050 664.050 ;
        RECT 817.950 663.600 820.050 664.050 ;
        RECT 751.950 662.400 820.050 663.600 ;
        RECT 751.950 661.950 754.050 662.400 ;
        RECT 814.950 661.950 817.050 662.400 ;
        RECT 817.950 661.950 820.050 662.400 ;
        RECT 841.950 663.600 844.050 664.050 ;
        RECT 853.950 663.600 856.050 664.050 ;
        RECT 841.950 662.400 856.050 663.600 ;
        RECT 841.950 661.950 844.050 662.400 ;
        RECT 853.950 661.950 856.050 662.400 ;
        RECT 97.950 660.600 100.050 661.050 ;
        RECT 142.950 660.600 145.050 661.050 ;
        RECT 97.950 659.400 145.050 660.600 ;
        RECT 97.950 658.950 100.050 659.400 ;
        RECT 142.950 658.950 145.050 659.400 ;
        RECT 247.950 660.600 250.050 661.050 ;
        RECT 349.950 660.600 352.050 661.050 ;
        RECT 247.950 659.400 352.050 660.600 ;
        RECT 247.950 658.950 250.050 659.400 ;
        RECT 349.950 658.950 352.050 659.400 ;
        RECT 727.950 660.600 730.050 661.050 ;
        RECT 790.950 660.600 793.050 661.050 ;
        RECT 727.950 659.400 793.050 660.600 ;
        RECT 727.950 658.950 730.050 659.400 ;
        RECT 790.950 658.950 793.050 659.400 ;
        RECT 253.950 657.600 256.050 658.050 ;
        RECT 271.950 657.600 274.050 658.050 ;
        RECT 253.950 656.400 274.050 657.600 ;
        RECT 253.950 655.950 256.050 656.400 ;
        RECT 271.950 655.950 274.050 656.400 ;
        RECT 322.950 657.600 325.050 658.050 ;
        RECT 337.950 657.600 340.050 658.050 ;
        RECT 322.950 656.400 340.050 657.600 ;
        RECT 322.950 655.950 325.050 656.400 ;
        RECT 337.950 655.950 340.050 656.400 ;
        RECT 676.950 657.600 679.050 658.050 ;
        RECT 721.950 657.600 724.050 658.050 ;
        RECT 676.950 656.400 724.050 657.600 ;
        RECT 676.950 655.950 679.050 656.400 ;
        RECT 721.950 655.950 724.050 656.400 ;
        RECT 769.950 657.600 772.050 658.050 ;
        RECT 787.950 657.600 790.050 658.050 ;
        RECT 769.950 656.400 790.050 657.600 ;
        RECT 769.950 655.950 772.050 656.400 ;
        RECT 787.950 655.950 790.050 656.400 ;
        RECT 124.950 654.600 127.050 655.050 ;
        RECT 160.950 654.600 163.050 655.050 ;
        RECT 178.950 654.600 181.050 655.050 ;
        RECT 124.950 653.400 181.050 654.600 ;
        RECT 124.950 652.950 127.050 653.400 ;
        RECT 160.950 652.950 163.050 653.400 ;
        RECT 178.950 652.950 181.050 653.400 ;
        RECT 271.950 654.600 274.050 655.050 ;
        RECT 283.950 654.600 286.050 655.050 ;
        RECT 271.950 653.400 286.050 654.600 ;
        RECT 271.950 652.950 274.050 653.400 ;
        RECT 283.950 652.950 286.050 653.400 ;
        RECT 346.950 654.600 349.050 655.050 ;
        RECT 391.950 654.600 394.050 655.050 ;
        RECT 346.950 653.400 394.050 654.600 ;
        RECT 346.950 652.950 349.050 653.400 ;
        RECT 391.950 652.950 394.050 653.400 ;
        RECT 472.950 654.600 475.050 655.050 ;
        RECT 505.950 654.600 508.050 655.050 ;
        RECT 472.950 653.400 508.050 654.600 ;
        RECT 472.950 652.950 475.050 653.400 ;
        RECT 505.950 652.950 508.050 653.400 ;
        RECT 787.950 654.600 790.050 655.050 ;
        RECT 826.950 654.600 829.050 655.050 ;
        RECT 787.950 653.400 829.050 654.600 ;
        RECT 787.950 652.950 790.050 653.400 ;
        RECT 826.950 652.950 829.050 653.400 ;
        RECT 124.950 651.600 127.050 652.050 ;
        RECT 208.950 651.600 211.050 652.050 ;
        RECT 250.950 651.600 253.050 652.050 ;
        RECT 124.950 650.400 253.050 651.600 ;
        RECT 124.950 649.950 127.050 650.400 ;
        RECT 208.950 649.950 211.050 650.400 ;
        RECT 250.950 649.950 253.050 650.400 ;
        RECT 373.950 651.600 376.050 652.050 ;
        RECT 505.950 651.600 508.050 652.050 ;
        RECT 373.950 650.400 508.050 651.600 ;
        RECT 373.950 649.950 376.050 650.400 ;
        RECT 505.950 649.950 508.050 650.400 ;
        RECT 361.950 648.600 364.050 649.050 ;
        RECT 379.950 648.600 382.050 649.050 ;
        RECT 361.950 647.400 382.050 648.600 ;
        RECT 361.950 646.950 364.050 647.400 ;
        RECT 379.950 646.950 382.050 647.400 ;
        RECT 469.950 648.600 472.050 649.050 ;
        RECT 478.950 648.600 481.050 649.050 ;
        RECT 469.950 647.400 481.050 648.600 ;
        RECT 469.950 646.950 472.050 647.400 ;
        RECT 478.950 646.950 481.050 647.400 ;
        RECT 595.950 648.600 598.050 649.050 ;
        RECT 772.950 648.600 775.050 649.050 ;
        RECT 595.950 647.400 775.050 648.600 ;
        RECT 595.950 646.950 598.050 647.400 ;
        RECT 772.950 646.950 775.050 647.400 ;
        RECT 268.950 645.600 271.050 646.050 ;
        RECT 286.950 645.600 289.050 646.050 ;
        RECT 379.950 645.600 382.050 646.050 ;
        RECT 268.950 644.400 382.050 645.600 ;
        RECT 268.950 643.950 271.050 644.400 ;
        RECT 286.950 643.950 289.050 644.400 ;
        RECT 379.950 643.950 382.050 644.400 ;
        RECT 274.950 642.600 277.050 643.050 ;
        RECT 325.950 642.600 328.050 643.050 ;
        RECT 274.950 641.400 328.050 642.600 ;
        RECT 274.950 640.950 277.050 641.400 ;
        RECT 325.950 640.950 328.050 641.400 ;
        RECT 376.950 642.600 379.050 643.050 ;
        RECT 391.950 642.600 394.050 643.050 ;
        RECT 376.950 641.400 394.050 642.600 ;
        RECT 376.950 640.950 379.050 641.400 ;
        RECT 391.950 640.950 394.050 641.400 ;
        RECT 490.950 642.600 493.050 643.050 ;
        RECT 502.950 642.600 505.050 643.050 ;
        RECT 490.950 641.400 505.050 642.600 ;
        RECT 490.950 640.950 493.050 641.400 ;
        RECT 502.950 640.950 505.050 641.400 ;
        RECT 691.950 642.600 694.050 643.050 ;
        RECT 697.950 642.600 700.050 643.050 ;
        RECT 691.950 641.400 700.050 642.600 ;
        RECT 691.950 640.950 694.050 641.400 ;
        RECT 697.950 640.950 700.050 641.400 ;
        RECT 298.950 639.600 301.050 640.050 ;
        RECT 313.950 639.600 316.050 640.050 ;
        RECT 421.950 639.600 424.050 640.050 ;
        RECT 463.950 639.600 466.050 640.050 ;
        RECT 298.950 638.400 466.050 639.600 ;
        RECT 298.950 637.950 301.050 638.400 ;
        RECT 313.950 637.950 316.050 638.400 ;
        RECT 421.950 637.950 424.050 638.400 ;
        RECT 463.950 637.950 466.050 638.400 ;
        RECT 622.950 639.600 625.050 640.050 ;
        RECT 691.950 639.600 694.050 640.050 ;
        RECT 775.950 639.600 778.050 640.050 ;
        RECT 622.950 638.400 778.050 639.600 ;
        RECT 622.950 637.950 625.050 638.400 ;
        RECT 691.950 637.950 694.050 638.400 ;
        RECT 775.950 637.950 778.050 638.400 ;
        RECT 115.950 636.600 118.050 637.050 ;
        RECT 172.950 636.600 175.050 637.050 ;
        RECT 115.950 635.400 175.050 636.600 ;
        RECT 115.950 634.950 118.050 635.400 ;
        RECT 172.950 634.950 175.050 635.400 ;
        RECT 190.950 636.600 193.050 637.050 ;
        RECT 262.950 636.600 265.050 637.050 ;
        RECT 295.950 636.600 298.050 637.050 ;
        RECT 190.950 635.400 243.600 636.600 ;
        RECT 190.950 634.950 193.050 635.400 ;
        RECT 242.400 634.050 243.600 635.400 ;
        RECT 262.950 635.400 298.050 636.600 ;
        RECT 262.950 634.950 265.050 635.400 ;
        RECT 295.950 634.950 298.050 635.400 ;
        RECT 304.950 636.600 307.050 637.050 ;
        RECT 316.950 636.600 319.050 637.050 ;
        RECT 304.950 635.400 319.050 636.600 ;
        RECT 304.950 634.950 307.050 635.400 ;
        RECT 316.950 634.950 319.050 635.400 ;
        RECT 331.950 636.600 334.050 637.050 ;
        RECT 343.950 636.600 346.050 637.050 ;
        RECT 331.950 635.400 346.050 636.600 ;
        RECT 331.950 634.950 334.050 635.400 ;
        RECT 343.950 634.950 346.050 635.400 ;
        RECT 376.950 636.600 379.050 637.050 ;
        RECT 424.950 636.600 427.050 637.050 ;
        RECT 376.950 635.400 427.050 636.600 ;
        RECT 376.950 634.950 379.050 635.400 ;
        RECT 424.950 634.950 427.050 635.400 ;
        RECT 439.950 636.600 442.050 637.050 ;
        RECT 445.950 636.600 448.050 637.050 ;
        RECT 439.950 635.400 448.050 636.600 ;
        RECT 439.950 634.950 442.050 635.400 ;
        RECT 445.950 634.950 448.050 635.400 ;
        RECT 466.950 636.600 469.050 637.050 ;
        RECT 508.950 636.600 511.050 637.050 ;
        RECT 466.950 635.400 511.050 636.600 ;
        RECT 466.950 634.950 469.050 635.400 ;
        RECT 508.950 634.950 511.050 635.400 ;
        RECT 511.950 636.600 514.050 637.050 ;
        RECT 517.950 636.600 520.050 637.050 ;
        RECT 511.950 635.400 520.050 636.600 ;
        RECT 511.950 634.950 514.050 635.400 ;
        RECT 517.950 634.950 520.050 635.400 ;
        RECT 541.950 636.600 544.050 637.050 ;
        RECT 547.950 636.600 550.050 637.050 ;
        RECT 541.950 635.400 550.050 636.600 ;
        RECT 541.950 634.950 544.050 635.400 ;
        RECT 547.950 634.950 550.050 635.400 ;
        RECT 580.950 636.600 583.050 637.050 ;
        RECT 586.950 636.600 589.050 637.050 ;
        RECT 580.950 635.400 589.050 636.600 ;
        RECT 580.950 634.950 583.050 635.400 ;
        RECT 586.950 634.950 589.050 635.400 ;
        RECT 613.950 636.600 616.050 637.050 ;
        RECT 700.950 636.600 703.050 637.050 ;
        RECT 613.950 635.400 703.050 636.600 ;
        RECT 613.950 634.950 616.050 635.400 ;
        RECT 700.950 634.950 703.050 635.400 ;
        RECT 772.950 636.600 775.050 637.050 ;
        RECT 838.950 636.600 841.050 637.050 ;
        RECT 772.950 635.400 841.050 636.600 ;
        RECT 772.950 634.950 775.050 635.400 ;
        RECT 838.950 634.950 841.050 635.400 ;
        RECT 139.950 633.600 142.050 634.050 ;
        RECT 148.950 633.600 151.050 634.050 ;
        RECT 157.950 633.600 160.050 634.050 ;
        RECT 139.950 632.400 160.050 633.600 ;
        RECT 139.950 631.950 142.050 632.400 ;
        RECT 148.950 631.950 151.050 632.400 ;
        RECT 157.950 631.950 160.050 632.400 ;
        RECT 160.950 633.600 163.050 634.050 ;
        RECT 166.950 633.600 169.050 634.050 ;
        RECT 160.950 632.400 169.050 633.600 ;
        RECT 160.950 631.950 163.050 632.400 ;
        RECT 166.950 631.950 169.050 632.400 ;
        RECT 178.950 633.600 181.050 634.050 ;
        RECT 217.950 633.600 220.050 634.050 ;
        RECT 178.950 632.400 220.050 633.600 ;
        RECT 178.950 631.950 181.050 632.400 ;
        RECT 217.950 631.950 220.050 632.400 ;
        RECT 223.950 633.600 226.050 634.050 ;
        RECT 232.950 633.600 235.050 634.050 ;
        RECT 235.950 633.600 238.050 634.050 ;
        RECT 223.950 632.400 238.050 633.600 ;
        RECT 223.950 631.950 226.050 632.400 ;
        RECT 232.950 631.950 235.050 632.400 ;
        RECT 235.950 631.950 238.050 632.400 ;
        RECT 241.950 631.950 244.050 634.050 ;
        RECT 277.950 633.600 280.050 634.050 ;
        RECT 286.950 633.600 289.050 634.050 ;
        RECT 277.950 632.400 289.050 633.600 ;
        RECT 277.950 631.950 280.050 632.400 ;
        RECT 286.950 631.950 289.050 632.400 ;
        RECT 289.950 631.950 292.050 634.050 ;
        RECT 292.950 633.600 295.050 634.050 ;
        RECT 298.950 633.600 301.050 634.050 ;
        RECT 307.950 633.600 310.050 634.050 ;
        RECT 292.950 632.400 310.050 633.600 ;
        RECT 292.950 631.950 295.050 632.400 ;
        RECT 298.950 631.950 301.050 632.400 ;
        RECT 307.950 631.950 310.050 632.400 ;
        RECT 349.950 633.600 352.050 634.050 ;
        RECT 367.950 633.600 370.050 634.050 ;
        RECT 349.950 632.400 370.050 633.600 ;
        RECT 349.950 631.950 352.050 632.400 ;
        RECT 367.950 631.950 370.050 632.400 ;
        RECT 400.950 633.600 403.050 634.050 ;
        RECT 448.950 633.600 451.050 634.050 ;
        RECT 400.950 632.400 451.050 633.600 ;
        RECT 400.950 631.950 403.050 632.400 ;
        RECT 448.950 631.950 451.050 632.400 ;
        RECT 463.950 633.600 466.050 634.050 ;
        RECT 475.950 633.600 478.050 634.050 ;
        RECT 463.950 632.400 478.050 633.600 ;
        RECT 463.950 631.950 466.050 632.400 ;
        RECT 475.950 631.950 478.050 632.400 ;
        RECT 490.950 633.600 493.050 634.050 ;
        RECT 499.950 633.600 502.050 634.050 ;
        RECT 490.950 632.400 502.050 633.600 ;
        RECT 490.950 631.950 493.050 632.400 ;
        RECT 499.950 631.950 502.050 632.400 ;
        RECT 505.950 633.600 508.050 634.050 ;
        RECT 514.950 633.600 517.050 634.050 ;
        RECT 520.950 633.600 523.050 634.050 ;
        RECT 505.950 632.400 523.050 633.600 ;
        RECT 505.950 631.950 508.050 632.400 ;
        RECT 514.950 631.950 517.050 632.400 ;
        RECT 520.950 631.950 523.050 632.400 ;
        RECT 532.950 633.600 535.050 634.050 ;
        RECT 562.950 633.600 565.050 634.050 ;
        RECT 532.950 632.400 565.050 633.600 ;
        RECT 532.950 631.950 535.050 632.400 ;
        RECT 562.950 631.950 565.050 632.400 ;
        RECT 628.950 633.600 631.050 634.050 ;
        RECT 643.950 633.600 646.050 634.050 ;
        RECT 628.950 632.400 646.050 633.600 ;
        RECT 628.950 631.950 631.050 632.400 ;
        RECT 643.950 631.950 646.050 632.400 ;
        RECT 763.950 633.600 766.050 634.050 ;
        RECT 790.950 633.600 793.050 634.050 ;
        RECT 835.950 633.600 838.050 634.050 ;
        RECT 763.950 632.400 838.050 633.600 ;
        RECT 763.950 631.950 766.050 632.400 ;
        RECT 790.950 631.950 793.050 632.400 ;
        RECT 835.950 631.950 838.050 632.400 ;
        RECT 847.950 631.950 850.050 634.050 ;
        RECT 94.950 630.600 97.050 631.050 ;
        RECT 86.400 629.400 97.050 630.600 ;
        RECT 86.400 628.050 87.600 629.400 ;
        RECT 94.950 628.950 97.050 629.400 ;
        RECT 115.950 630.600 118.050 631.050 ;
        RECT 127.950 630.600 130.050 631.050 ;
        RECT 115.950 629.400 130.050 630.600 ;
        RECT 115.950 628.950 118.050 629.400 ;
        RECT 127.950 628.950 130.050 629.400 ;
        RECT 142.950 630.600 145.050 631.050 ;
        RECT 160.950 630.600 163.050 631.050 ;
        RECT 142.950 629.400 163.050 630.600 ;
        RECT 142.950 628.950 145.050 629.400 ;
        RECT 160.950 628.950 163.050 629.400 ;
        RECT 196.950 630.600 199.050 631.050 ;
        RECT 208.950 630.600 211.050 631.050 ;
        RECT 196.950 629.400 211.050 630.600 ;
        RECT 196.950 628.950 199.050 629.400 ;
        RECT 208.950 628.950 211.050 629.400 ;
        RECT 238.950 630.600 241.050 631.050 ;
        RECT 280.950 630.600 283.050 631.050 ;
        RECT 238.950 629.400 283.050 630.600 ;
        RECT 238.950 628.950 241.050 629.400 ;
        RECT 280.950 628.950 283.050 629.400 ;
        RECT 25.950 627.600 28.050 628.050 ;
        RECT 79.950 627.600 82.050 628.050 ;
        RECT 25.950 626.400 82.050 627.600 ;
        RECT 25.950 625.950 28.050 626.400 ;
        RECT 79.950 625.950 82.050 626.400 ;
        RECT 85.950 625.950 88.050 628.050 ;
        RECT 130.950 627.600 133.050 628.050 ;
        RECT 145.950 627.600 148.050 628.050 ;
        RECT 130.950 626.400 148.050 627.600 ;
        RECT 130.950 625.950 133.050 626.400 ;
        RECT 145.950 625.950 148.050 626.400 ;
        RECT 151.950 627.600 154.050 628.050 ;
        RECT 190.950 627.600 193.050 628.050 ;
        RECT 151.950 626.400 193.050 627.600 ;
        RECT 151.950 625.950 154.050 626.400 ;
        RECT 190.950 625.950 193.050 626.400 ;
        RECT 193.950 627.600 196.050 628.050 ;
        RECT 202.950 627.600 205.050 628.050 ;
        RECT 193.950 626.400 205.050 627.600 ;
        RECT 193.950 625.950 196.050 626.400 ;
        RECT 202.950 625.950 205.050 626.400 ;
        RECT 283.950 627.600 286.050 628.050 ;
        RECT 290.400 627.600 291.600 631.950 ;
        RECT 310.950 630.600 313.050 631.050 ;
        RECT 337.950 630.600 340.050 631.050 ;
        RECT 310.950 629.400 340.050 630.600 ;
        RECT 310.950 628.950 313.050 629.400 ;
        RECT 337.950 628.950 340.050 629.400 ;
        RECT 358.950 630.600 361.050 631.050 ;
        RECT 445.950 630.600 448.050 631.050 ;
        RECT 508.950 630.600 511.050 631.050 ;
        RECT 358.950 629.400 384.600 630.600 ;
        RECT 358.950 628.950 361.050 629.400 ;
        RECT 283.950 626.400 291.600 627.600 ;
        RECT 295.950 627.600 298.050 628.050 ;
        RECT 319.950 627.600 322.050 628.050 ;
        RECT 295.950 626.400 322.050 627.600 ;
        RECT 283.950 625.950 286.050 626.400 ;
        RECT 295.950 625.950 298.050 626.400 ;
        RECT 319.950 625.950 322.050 626.400 ;
        RECT 358.950 627.600 361.050 628.050 ;
        RECT 364.950 627.600 367.050 628.050 ;
        RECT 358.950 626.400 367.050 627.600 ;
        RECT 358.950 625.950 361.050 626.400 ;
        RECT 364.950 625.950 367.050 626.400 ;
        RECT 373.950 627.600 376.050 628.050 ;
        RECT 379.950 627.600 382.050 628.050 ;
        RECT 373.950 626.400 382.050 627.600 ;
        RECT 383.400 627.600 384.600 629.400 ;
        RECT 445.950 629.400 511.050 630.600 ;
        RECT 445.950 628.950 448.050 629.400 ;
        RECT 508.950 628.950 511.050 629.400 ;
        RECT 535.950 630.600 538.050 631.050 ;
        RECT 544.950 630.600 547.050 631.050 ;
        RECT 535.950 629.400 547.050 630.600 ;
        RECT 535.950 628.950 538.050 629.400 ;
        RECT 544.950 628.950 547.050 629.400 ;
        RECT 550.950 630.600 553.050 631.050 ;
        RECT 595.950 630.600 598.050 631.050 ;
        RECT 550.950 629.400 598.050 630.600 ;
        RECT 550.950 628.950 553.050 629.400 ;
        RECT 595.950 628.950 598.050 629.400 ;
        RECT 598.950 630.600 601.050 631.050 ;
        RECT 631.950 630.600 634.050 631.050 ;
        RECT 646.950 630.600 649.050 631.050 ;
        RECT 598.950 629.400 649.050 630.600 ;
        RECT 598.950 628.950 601.050 629.400 ;
        RECT 631.950 628.950 634.050 629.400 ;
        RECT 646.950 628.950 649.050 629.400 ;
        RECT 652.950 630.600 655.050 631.050 ;
        RECT 658.950 630.600 661.050 631.050 ;
        RECT 676.950 630.600 679.050 631.050 ;
        RECT 652.950 629.400 661.050 630.600 ;
        RECT 652.950 628.950 655.050 629.400 ;
        RECT 658.950 628.950 661.050 629.400 ;
        RECT 671.400 629.400 679.050 630.600 ;
        RECT 388.950 627.600 391.050 628.050 ;
        RECT 403.950 627.600 406.050 628.050 ;
        RECT 383.400 626.400 406.050 627.600 ;
        RECT 373.950 625.950 376.050 626.400 ;
        RECT 379.950 625.950 382.050 626.400 ;
        RECT 388.950 625.950 391.050 626.400 ;
        RECT 403.950 625.950 406.050 626.400 ;
        RECT 412.950 627.600 415.050 628.050 ;
        RECT 427.950 627.600 430.050 628.050 ;
        RECT 412.950 626.400 430.050 627.600 ;
        RECT 412.950 625.950 415.050 626.400 ;
        RECT 427.950 625.950 430.050 626.400 ;
        RECT 436.950 627.600 439.050 628.050 ;
        RECT 442.950 627.600 445.050 628.050 ;
        RECT 436.950 626.400 445.050 627.600 ;
        RECT 436.950 625.950 439.050 626.400 ;
        RECT 442.950 625.950 445.050 626.400 ;
        RECT 469.950 627.600 472.050 628.050 ;
        RECT 478.950 627.600 481.050 628.050 ;
        RECT 496.950 627.600 499.050 628.050 ;
        RECT 469.950 626.400 499.050 627.600 ;
        RECT 469.950 625.950 472.050 626.400 ;
        RECT 478.950 625.950 481.050 626.400 ;
        RECT 496.950 625.950 499.050 626.400 ;
        RECT 526.950 627.600 529.050 628.050 ;
        RECT 532.950 627.600 535.050 628.050 ;
        RECT 526.950 626.400 535.050 627.600 ;
        RECT 526.950 625.950 529.050 626.400 ;
        RECT 532.950 625.950 535.050 626.400 ;
        RECT 565.950 627.600 568.050 628.050 ;
        RECT 604.950 627.600 607.050 628.050 ;
        RECT 565.950 626.400 607.050 627.600 ;
        RECT 565.950 625.950 568.050 626.400 ;
        RECT 604.950 625.950 607.050 626.400 ;
        RECT 616.950 627.600 619.050 628.050 ;
        RECT 637.950 627.600 640.050 628.050 ;
        RECT 616.950 626.400 640.050 627.600 ;
        RECT 616.950 625.950 619.050 626.400 ;
        RECT 637.950 625.950 640.050 626.400 ;
        RECT 655.950 627.600 658.050 628.050 ;
        RECT 671.400 627.600 672.600 629.400 ;
        RECT 676.950 628.950 679.050 629.400 ;
        RECT 685.950 630.600 688.050 631.050 ;
        RECT 700.950 630.600 703.050 631.050 ;
        RECT 685.950 629.400 703.050 630.600 ;
        RECT 685.950 628.950 688.050 629.400 ;
        RECT 700.950 628.950 703.050 629.400 ;
        RECT 718.950 630.600 721.050 631.050 ;
        RECT 739.950 630.600 742.050 631.050 ;
        RECT 718.950 629.400 742.050 630.600 ;
        RECT 718.950 628.950 721.050 629.400 ;
        RECT 739.950 628.950 742.050 629.400 ;
        RECT 778.950 630.600 781.050 631.050 ;
        RECT 811.950 630.600 814.050 631.050 ;
        RECT 778.950 629.400 814.050 630.600 ;
        RECT 778.950 628.950 781.050 629.400 ;
        RECT 811.950 628.950 814.050 629.400 ;
        RECT 655.950 626.400 672.600 627.600 ;
        RECT 673.950 627.600 676.050 628.050 ;
        RECT 688.950 627.600 691.050 628.050 ;
        RECT 673.950 626.400 691.050 627.600 ;
        RECT 655.950 625.950 658.050 626.400 ;
        RECT 673.950 625.950 676.050 626.400 ;
        RECT 688.950 625.950 691.050 626.400 ;
        RECT 715.950 627.600 718.050 628.050 ;
        RECT 784.950 627.600 787.050 628.050 ;
        RECT 715.950 626.400 787.050 627.600 ;
        RECT 715.950 625.950 718.050 626.400 ;
        RECT 784.950 625.950 787.050 626.400 ;
        RECT 70.950 624.600 73.050 625.050 ;
        RECT 97.950 624.600 100.050 625.050 ;
        RECT 70.950 623.400 100.050 624.600 ;
        RECT 70.950 622.950 73.050 623.400 ;
        RECT 97.950 622.950 100.050 623.400 ;
        RECT 109.950 624.600 112.050 625.050 ;
        RECT 112.950 624.600 115.050 625.050 ;
        RECT 118.950 624.600 121.050 625.050 ;
        RECT 127.950 624.600 130.050 625.050 ;
        RECT 109.950 623.400 130.050 624.600 ;
        RECT 109.950 622.950 112.050 623.400 ;
        RECT 112.950 622.950 115.050 623.400 ;
        RECT 118.950 622.950 121.050 623.400 ;
        RECT 127.950 622.950 130.050 623.400 ;
        RECT 157.950 624.600 160.050 625.050 ;
        RECT 223.950 624.600 226.050 625.050 ;
        RECT 157.950 623.400 226.050 624.600 ;
        RECT 157.950 622.950 160.050 623.400 ;
        RECT 223.950 622.950 226.050 623.400 ;
        RECT 235.950 624.600 238.050 625.050 ;
        RECT 265.950 624.600 268.050 625.050 ;
        RECT 235.950 623.400 268.050 624.600 ;
        RECT 235.950 622.950 238.050 623.400 ;
        RECT 265.950 622.950 268.050 623.400 ;
        RECT 301.950 624.600 304.050 625.050 ;
        RECT 310.950 624.600 313.050 625.050 ;
        RECT 301.950 623.400 313.050 624.600 ;
        RECT 301.950 622.950 304.050 623.400 ;
        RECT 310.950 622.950 313.050 623.400 ;
        RECT 343.950 624.600 346.050 625.050 ;
        RECT 364.950 624.600 367.050 625.050 ;
        RECT 343.950 623.400 367.050 624.600 ;
        RECT 343.950 622.950 346.050 623.400 ;
        RECT 364.950 622.950 367.050 623.400 ;
        RECT 367.950 624.600 370.050 625.050 ;
        RECT 376.950 624.600 379.050 625.050 ;
        RECT 382.950 624.600 385.050 625.050 ;
        RECT 367.950 623.400 385.050 624.600 ;
        RECT 367.950 622.950 370.050 623.400 ;
        RECT 376.950 622.950 379.050 623.400 ;
        RECT 382.950 622.950 385.050 623.400 ;
        RECT 430.950 624.600 433.050 625.050 ;
        RECT 460.950 624.600 463.050 625.050 ;
        RECT 469.950 624.600 472.050 625.050 ;
        RECT 430.950 623.400 472.050 624.600 ;
        RECT 430.950 622.950 433.050 623.400 ;
        RECT 460.950 622.950 463.050 623.400 ;
        RECT 469.950 622.950 472.050 623.400 ;
        RECT 484.950 624.600 487.050 625.050 ;
        RECT 508.950 624.600 511.050 625.050 ;
        RECT 484.950 623.400 511.050 624.600 ;
        RECT 484.950 622.950 487.050 623.400 ;
        RECT 508.950 622.950 511.050 623.400 ;
        RECT 523.950 624.600 526.050 625.050 ;
        RECT 538.950 624.600 541.050 625.050 ;
        RECT 523.950 623.400 541.050 624.600 ;
        RECT 523.950 622.950 526.050 623.400 ;
        RECT 538.950 622.950 541.050 623.400 ;
        RECT 553.950 624.600 556.050 625.050 ;
        RECT 559.950 624.600 562.050 625.050 ;
        RECT 562.950 624.600 565.050 625.050 ;
        RECT 553.950 623.400 565.050 624.600 ;
        RECT 553.950 622.950 556.050 623.400 ;
        RECT 559.950 622.950 562.050 623.400 ;
        RECT 562.950 622.950 565.050 623.400 ;
        RECT 583.950 624.600 586.050 625.050 ;
        RECT 592.950 624.600 595.050 625.050 ;
        RECT 613.950 624.600 616.050 625.050 ;
        RECT 583.950 623.400 616.050 624.600 ;
        RECT 583.950 622.950 586.050 623.400 ;
        RECT 592.950 622.950 595.050 623.400 ;
        RECT 613.950 622.950 616.050 623.400 ;
        RECT 634.950 624.600 637.050 625.050 ;
        RECT 649.950 624.600 652.050 625.050 ;
        RECT 634.950 623.400 652.050 624.600 ;
        RECT 634.950 622.950 637.050 623.400 ;
        RECT 649.950 622.950 652.050 623.400 ;
        RECT 658.950 624.600 661.050 625.050 ;
        RECT 667.950 624.600 670.050 625.050 ;
        RECT 658.950 623.400 670.050 624.600 ;
        RECT 658.950 622.950 661.050 623.400 ;
        RECT 667.950 622.950 670.050 623.400 ;
        RECT 670.950 624.600 673.050 625.050 ;
        RECT 739.950 624.600 742.050 625.050 ;
        RECT 670.950 623.400 742.050 624.600 ;
        RECT 848.400 624.600 849.600 631.950 ;
        RECT 856.950 624.600 859.050 625.050 ;
        RECT 848.400 623.400 859.050 624.600 ;
        RECT 670.950 622.950 673.050 623.400 ;
        RECT 739.950 622.950 742.050 623.400 ;
        RECT 856.950 622.950 859.050 623.400 ;
        RECT 28.950 621.600 31.050 622.050 ;
        RECT 82.950 621.600 85.050 622.050 ;
        RECT 28.950 620.400 85.050 621.600 ;
        RECT 28.950 619.950 31.050 620.400 ;
        RECT 82.950 619.950 85.050 620.400 ;
        RECT 100.950 621.600 103.050 622.050 ;
        RECT 181.950 621.600 184.050 622.050 ;
        RECT 100.950 620.400 184.050 621.600 ;
        RECT 100.950 619.950 103.050 620.400 ;
        RECT 181.950 619.950 184.050 620.400 ;
        RECT 205.950 621.600 208.050 622.050 ;
        RECT 235.950 621.600 238.050 622.050 ;
        RECT 205.950 620.400 238.050 621.600 ;
        RECT 205.950 619.950 208.050 620.400 ;
        RECT 235.950 619.950 238.050 620.400 ;
        RECT 280.950 621.600 283.050 622.050 ;
        RECT 352.950 621.600 355.050 622.050 ;
        RECT 280.950 620.400 355.050 621.600 ;
        RECT 280.950 619.950 283.050 620.400 ;
        RECT 352.950 619.950 355.050 620.400 ;
        RECT 361.950 621.600 364.050 622.050 ;
        RECT 379.950 621.600 382.050 622.050 ;
        RECT 361.950 620.400 382.050 621.600 ;
        RECT 361.950 619.950 364.050 620.400 ;
        RECT 379.950 619.950 382.050 620.400 ;
        RECT 547.950 621.600 550.050 622.050 ;
        RECT 571.950 621.600 574.050 622.050 ;
        RECT 589.950 621.600 592.050 622.050 ;
        RECT 547.950 620.400 592.050 621.600 ;
        RECT 547.950 619.950 550.050 620.400 ;
        RECT 571.950 619.950 574.050 620.400 ;
        RECT 589.950 619.950 592.050 620.400 ;
        RECT 637.950 621.600 640.050 622.050 ;
        RECT 754.950 621.600 757.050 622.050 ;
        RECT 637.950 620.400 757.050 621.600 ;
        RECT 637.950 619.950 640.050 620.400 ;
        RECT 754.950 619.950 757.050 620.400 ;
        RECT 109.950 618.600 112.050 619.050 ;
        RECT 124.950 618.600 127.050 619.050 ;
        RECT 109.950 617.400 127.050 618.600 ;
        RECT 109.950 616.950 112.050 617.400 ;
        RECT 124.950 616.950 127.050 617.400 ;
        RECT 127.950 618.600 130.050 619.050 ;
        RECT 151.950 618.600 154.050 619.050 ;
        RECT 127.950 617.400 154.050 618.600 ;
        RECT 127.950 616.950 130.050 617.400 ;
        RECT 151.950 616.950 154.050 617.400 ;
        RECT 220.950 618.600 223.050 619.050 ;
        RECT 232.950 618.600 235.050 619.050 ;
        RECT 244.950 618.600 247.050 619.050 ;
        RECT 220.950 617.400 247.050 618.600 ;
        RECT 220.950 616.950 223.050 617.400 ;
        RECT 232.950 616.950 235.050 617.400 ;
        RECT 244.950 616.950 247.050 617.400 ;
        RECT 265.950 618.600 268.050 619.050 ;
        RECT 271.950 618.600 274.050 619.050 ;
        RECT 265.950 617.400 274.050 618.600 ;
        RECT 265.950 616.950 268.050 617.400 ;
        RECT 271.950 616.950 274.050 617.400 ;
        RECT 325.950 618.600 328.050 619.050 ;
        RECT 415.950 618.600 418.050 619.050 ;
        RECT 325.950 617.400 418.050 618.600 ;
        RECT 325.950 616.950 328.050 617.400 ;
        RECT 415.950 616.950 418.050 617.400 ;
        RECT 577.950 618.600 580.050 619.050 ;
        RECT 634.950 618.600 637.050 619.050 ;
        RECT 577.950 617.400 637.050 618.600 ;
        RECT 577.950 616.950 580.050 617.400 ;
        RECT 634.950 616.950 637.050 617.400 ;
        RECT 643.950 618.600 646.050 619.050 ;
        RECT 664.950 618.600 667.050 619.050 ;
        RECT 643.950 617.400 667.050 618.600 ;
        RECT 643.950 616.950 646.050 617.400 ;
        RECT 664.950 616.950 667.050 617.400 ;
        RECT 787.950 618.600 790.050 619.050 ;
        RECT 811.950 618.600 814.050 619.050 ;
        RECT 823.950 618.600 826.050 619.050 ;
        RECT 787.950 617.400 804.600 618.600 ;
        RECT 787.950 616.950 790.050 617.400 ;
        RECT 112.950 615.600 115.050 616.050 ;
        RECT 208.950 615.600 211.050 616.050 ;
        RECT 112.950 614.400 211.050 615.600 ;
        RECT 112.950 613.950 115.050 614.400 ;
        RECT 208.950 613.950 211.050 614.400 ;
        RECT 340.950 615.600 343.050 616.050 ;
        RECT 367.950 615.600 370.050 616.050 ;
        RECT 340.950 614.400 370.050 615.600 ;
        RECT 340.950 613.950 343.050 614.400 ;
        RECT 367.950 613.950 370.050 614.400 ;
        RECT 442.950 615.600 445.050 616.050 ;
        RECT 454.950 615.600 457.050 616.050 ;
        RECT 520.950 615.600 523.050 616.050 ;
        RECT 442.950 614.400 523.050 615.600 ;
        RECT 442.950 613.950 445.050 614.400 ;
        RECT 454.950 613.950 457.050 614.400 ;
        RECT 520.950 613.950 523.050 614.400 ;
        RECT 565.950 615.600 568.050 616.050 ;
        RECT 610.950 615.600 613.050 616.050 ;
        RECT 619.950 615.600 622.050 616.050 ;
        RECT 565.950 614.400 622.050 615.600 ;
        RECT 565.950 613.950 568.050 614.400 ;
        RECT 610.950 613.950 613.050 614.400 ;
        RECT 619.950 613.950 622.050 614.400 ;
        RECT 622.950 615.600 625.050 616.050 ;
        RECT 634.950 615.600 637.050 616.050 ;
        RECT 622.950 614.400 637.050 615.600 ;
        RECT 622.950 613.950 625.050 614.400 ;
        RECT 634.950 613.950 637.050 614.400 ;
        RECT 679.950 615.600 682.050 616.050 ;
        RECT 733.950 615.600 736.050 616.050 ;
        RECT 679.950 614.400 736.050 615.600 ;
        RECT 679.950 613.950 682.050 614.400 ;
        RECT 733.950 613.950 736.050 614.400 ;
        RECT 772.950 615.600 775.050 616.050 ;
        RECT 778.950 615.600 781.050 616.050 ;
        RECT 772.950 614.400 781.050 615.600 ;
        RECT 772.950 613.950 775.050 614.400 ;
        RECT 778.950 613.950 781.050 614.400 ;
        RECT 787.950 615.600 790.050 616.050 ;
        RECT 799.950 615.600 802.050 616.050 ;
        RECT 787.950 614.400 802.050 615.600 ;
        RECT 803.400 615.600 804.600 617.400 ;
        RECT 811.950 617.400 826.050 618.600 ;
        RECT 811.950 616.950 814.050 617.400 ;
        RECT 823.950 616.950 826.050 617.400 ;
        RECT 811.950 615.600 814.050 616.050 ;
        RECT 803.400 614.400 814.050 615.600 ;
        RECT 787.950 613.950 790.050 614.400 ;
        RECT 799.950 613.950 802.050 614.400 ;
        RECT 811.950 613.950 814.050 614.400 ;
        RECT 124.950 612.600 127.050 613.050 ;
        RECT 133.950 612.600 136.050 613.050 ;
        RECT 124.950 611.400 136.050 612.600 ;
        RECT 124.950 610.950 127.050 611.400 ;
        RECT 133.950 610.950 136.050 611.400 ;
        RECT 151.950 612.600 154.050 613.050 ;
        RECT 190.950 612.600 193.050 613.050 ;
        RECT 238.950 612.600 241.050 613.050 ;
        RECT 151.950 611.400 241.050 612.600 ;
        RECT 151.950 610.950 154.050 611.400 ;
        RECT 190.950 610.950 193.050 611.400 ;
        RECT 238.950 610.950 241.050 611.400 ;
        RECT 241.950 612.600 244.050 613.050 ;
        RECT 289.950 612.600 292.050 613.050 ;
        RECT 409.950 612.600 412.050 613.050 ;
        RECT 241.950 611.400 412.050 612.600 ;
        RECT 241.950 610.950 244.050 611.400 ;
        RECT 289.950 610.950 292.050 611.400 ;
        RECT 409.950 610.950 412.050 611.400 ;
        RECT 448.950 612.600 451.050 613.050 ;
        RECT 454.950 612.600 457.050 613.050 ;
        RECT 448.950 611.400 457.050 612.600 ;
        RECT 448.950 610.950 451.050 611.400 ;
        RECT 454.950 610.950 457.050 611.400 ;
        RECT 460.950 612.600 463.050 613.050 ;
        RECT 493.950 612.600 496.050 613.050 ;
        RECT 460.950 611.400 496.050 612.600 ;
        RECT 460.950 610.950 463.050 611.400 ;
        RECT 493.950 610.950 496.050 611.400 ;
        RECT 520.950 612.600 523.050 613.050 ;
        RECT 532.950 612.600 535.050 613.050 ;
        RECT 520.950 611.400 535.050 612.600 ;
        RECT 520.950 610.950 523.050 611.400 ;
        RECT 532.950 610.950 535.050 611.400 ;
        RECT 538.950 612.600 541.050 613.050 ;
        RECT 562.950 612.600 565.050 613.050 ;
        RECT 538.950 611.400 565.050 612.600 ;
        RECT 538.950 610.950 541.050 611.400 ;
        RECT 562.950 610.950 565.050 611.400 ;
        RECT 643.950 612.600 646.050 613.050 ;
        RECT 703.950 612.600 706.050 613.050 ;
        RECT 643.950 611.400 706.050 612.600 ;
        RECT 643.950 610.950 646.050 611.400 ;
        RECT 703.950 610.950 706.050 611.400 ;
        RECT 718.950 612.600 721.050 613.050 ;
        RECT 736.950 612.600 739.050 613.050 ;
        RECT 718.950 611.400 739.050 612.600 ;
        RECT 718.950 610.950 721.050 611.400 ;
        RECT 736.950 610.950 739.050 611.400 ;
        RECT 769.950 612.600 772.050 613.050 ;
        RECT 784.950 612.600 787.050 613.050 ;
        RECT 796.950 612.600 799.050 613.050 ;
        RECT 769.950 611.400 799.050 612.600 ;
        RECT 769.950 610.950 772.050 611.400 ;
        RECT 784.950 610.950 787.050 611.400 ;
        RECT 796.950 610.950 799.050 611.400 ;
        RECT 118.950 609.600 121.050 610.050 ;
        RECT 136.950 609.600 139.050 610.050 ;
        RECT 118.950 608.400 139.050 609.600 ;
        RECT 118.950 607.950 121.050 608.400 ;
        RECT 136.950 607.950 139.050 608.400 ;
        RECT 145.950 609.600 148.050 610.050 ;
        RECT 154.950 609.600 157.050 610.050 ;
        RECT 145.950 608.400 157.050 609.600 ;
        RECT 145.950 607.950 148.050 608.400 ;
        RECT 154.950 607.950 157.050 608.400 ;
        RECT 238.950 609.600 241.050 610.050 ;
        RECT 304.950 609.600 307.050 610.050 ;
        RECT 238.950 608.400 307.050 609.600 ;
        RECT 238.950 607.950 241.050 608.400 ;
        RECT 304.950 607.950 307.050 608.400 ;
        RECT 334.950 609.600 337.050 610.050 ;
        RECT 343.950 609.600 346.050 610.050 ;
        RECT 334.950 608.400 346.050 609.600 ;
        RECT 334.950 607.950 337.050 608.400 ;
        RECT 343.950 607.950 346.050 608.400 ;
        RECT 346.950 609.600 349.050 610.050 ;
        RECT 361.950 609.600 364.050 610.050 ;
        RECT 346.950 608.400 364.050 609.600 ;
        RECT 346.950 607.950 349.050 608.400 ;
        RECT 361.950 607.950 364.050 608.400 ;
        RECT 385.950 609.600 388.050 610.050 ;
        RECT 625.950 609.600 628.050 610.050 ;
        RECT 649.950 609.600 652.050 610.050 ;
        RECT 694.950 609.600 697.050 610.050 ;
        RECT 385.950 608.400 697.050 609.600 ;
        RECT 385.950 607.950 388.050 608.400 ;
        RECT 625.950 607.950 628.050 608.400 ;
        RECT 649.950 607.950 652.050 608.400 ;
        RECT 694.950 607.950 697.050 608.400 ;
        RECT 706.950 609.600 709.050 610.050 ;
        RECT 712.950 609.600 715.050 610.050 ;
        RECT 748.950 609.600 751.050 610.050 ;
        RECT 706.950 608.400 751.050 609.600 ;
        RECT 706.950 607.950 709.050 608.400 ;
        RECT 712.950 607.950 715.050 608.400 ;
        RECT 748.950 607.950 751.050 608.400 ;
        RECT 766.950 609.600 769.050 610.050 ;
        RECT 775.950 609.600 778.050 610.050 ;
        RECT 808.950 609.600 811.050 610.050 ;
        RECT 766.950 608.400 811.050 609.600 ;
        RECT 766.950 607.950 769.050 608.400 ;
        RECT 775.950 607.950 778.050 608.400 ;
        RECT 808.950 607.950 811.050 608.400 ;
        RECT 829.950 609.600 832.050 610.050 ;
        RECT 850.950 609.600 853.050 610.050 ;
        RECT 829.950 608.400 853.050 609.600 ;
        RECT 829.950 607.950 832.050 608.400 ;
        RECT 850.950 607.950 853.050 608.400 ;
        RECT 121.950 606.600 124.050 607.050 ;
        RECT 127.950 606.600 130.050 607.050 ;
        RECT 121.950 605.400 130.050 606.600 ;
        RECT 121.950 604.950 124.050 605.400 ;
        RECT 127.950 604.950 130.050 605.400 ;
        RECT 133.950 606.600 136.050 607.050 ;
        RECT 139.950 606.600 142.050 607.050 ;
        RECT 133.950 605.400 142.050 606.600 ;
        RECT 133.950 604.950 136.050 605.400 ;
        RECT 139.950 604.950 142.050 605.400 ;
        RECT 217.950 606.600 220.050 607.050 ;
        RECT 259.950 606.600 262.050 607.050 ;
        RECT 217.950 605.400 262.050 606.600 ;
        RECT 217.950 604.950 220.050 605.400 ;
        RECT 259.950 604.950 262.050 605.400 ;
        RECT 274.950 606.600 277.050 607.050 ;
        RECT 316.950 606.600 319.050 607.050 ;
        RECT 274.950 605.400 319.050 606.600 ;
        RECT 274.950 604.950 277.050 605.400 ;
        RECT 316.950 604.950 319.050 605.400 ;
        RECT 319.950 606.600 322.050 607.050 ;
        RECT 346.950 606.600 349.050 607.050 ;
        RECT 319.950 605.400 349.050 606.600 ;
        RECT 319.950 604.950 322.050 605.400 ;
        RECT 346.950 604.950 349.050 605.400 ;
        RECT 364.950 606.600 367.050 607.050 ;
        RECT 406.950 606.600 409.050 607.050 ;
        RECT 364.950 605.400 409.050 606.600 ;
        RECT 364.950 604.950 367.050 605.400 ;
        RECT 406.950 604.950 409.050 605.400 ;
        RECT 484.950 606.600 487.050 607.050 ;
        RECT 496.950 606.600 499.050 607.050 ;
        RECT 484.950 605.400 499.050 606.600 ;
        RECT 484.950 604.950 487.050 605.400 ;
        RECT 496.950 604.950 499.050 605.400 ;
        RECT 508.950 606.600 511.050 607.050 ;
        RECT 520.950 606.600 523.050 607.050 ;
        RECT 508.950 605.400 523.050 606.600 ;
        RECT 508.950 604.950 511.050 605.400 ;
        RECT 520.950 604.950 523.050 605.400 ;
        RECT 535.950 606.600 538.050 607.050 ;
        RECT 547.950 606.600 550.050 607.050 ;
        RECT 535.950 605.400 550.050 606.600 ;
        RECT 535.950 604.950 538.050 605.400 ;
        RECT 547.950 604.950 550.050 605.400 ;
        RECT 553.950 606.600 556.050 607.050 ;
        RECT 568.950 606.600 571.050 607.050 ;
        RECT 553.950 605.400 571.050 606.600 ;
        RECT 553.950 604.950 556.050 605.400 ;
        RECT 568.950 604.950 571.050 605.400 ;
        RECT 604.950 606.600 607.050 607.050 ;
        RECT 691.950 606.600 694.050 607.050 ;
        RECT 604.950 605.400 694.050 606.600 ;
        RECT 604.950 604.950 607.050 605.400 ;
        RECT 691.950 604.950 694.050 605.400 ;
        RECT 694.950 606.600 697.050 607.050 ;
        RECT 778.950 606.600 781.050 607.050 ;
        RECT 802.950 606.600 805.050 607.050 ;
        RECT 832.950 606.600 835.050 607.050 ;
        RECT 835.950 606.600 838.050 607.050 ;
        RECT 694.950 605.400 838.050 606.600 ;
        RECT 694.950 604.950 697.050 605.400 ;
        RECT 778.950 604.950 781.050 605.400 ;
        RECT 802.950 604.950 805.050 605.400 ;
        RECT 832.950 604.950 835.050 605.400 ;
        RECT 835.950 604.950 838.050 605.400 ;
        RECT 841.950 606.600 844.050 607.050 ;
        RECT 850.950 606.600 853.050 607.050 ;
        RECT 841.950 605.400 853.050 606.600 ;
        RECT 841.950 604.950 844.050 605.400 ;
        RECT 850.950 604.950 853.050 605.400 ;
        RECT 28.950 603.600 31.050 604.050 ;
        RECT 82.950 603.600 85.050 604.050 ;
        RECT 28.950 602.400 85.050 603.600 ;
        RECT 28.950 601.950 31.050 602.400 ;
        RECT 82.950 601.950 85.050 602.400 ;
        RECT 112.950 603.600 115.050 604.050 ;
        RECT 133.950 603.600 136.050 604.050 ;
        RECT 112.950 602.400 136.050 603.600 ;
        RECT 112.950 601.950 115.050 602.400 ;
        RECT 133.950 601.950 136.050 602.400 ;
        RECT 136.950 603.600 139.050 604.050 ;
        RECT 154.950 603.600 157.050 604.050 ;
        RECT 136.950 602.400 157.050 603.600 ;
        RECT 136.950 601.950 139.050 602.400 ;
        RECT 154.950 601.950 157.050 602.400 ;
        RECT 163.950 603.600 166.050 604.050 ;
        RECT 181.950 603.600 184.050 604.050 ;
        RECT 163.950 602.400 184.050 603.600 ;
        RECT 163.950 601.950 166.050 602.400 ;
        RECT 181.950 601.950 184.050 602.400 ;
        RECT 202.950 603.600 205.050 604.050 ;
        RECT 211.950 603.600 214.050 604.050 ;
        RECT 202.950 602.400 214.050 603.600 ;
        RECT 202.950 601.950 205.050 602.400 ;
        RECT 211.950 601.950 214.050 602.400 ;
        RECT 214.950 603.600 217.050 604.050 ;
        RECT 220.950 603.600 223.050 604.050 ;
        RECT 229.950 603.600 232.050 604.050 ;
        RECT 214.950 602.400 232.050 603.600 ;
        RECT 214.950 601.950 217.050 602.400 ;
        RECT 220.950 601.950 223.050 602.400 ;
        RECT 229.950 601.950 232.050 602.400 ;
        RECT 259.950 603.600 262.050 604.050 ;
        RECT 295.950 603.600 298.050 604.050 ;
        RECT 259.950 602.400 298.050 603.600 ;
        RECT 259.950 601.950 262.050 602.400 ;
        RECT 295.950 601.950 298.050 602.400 ;
        RECT 340.950 603.600 343.050 604.050 ;
        RECT 346.950 603.600 349.050 604.050 ;
        RECT 340.950 602.400 349.050 603.600 ;
        RECT 340.950 601.950 343.050 602.400 ;
        RECT 346.950 601.950 349.050 602.400 ;
        RECT 370.950 603.600 373.050 604.050 ;
        RECT 388.950 603.600 391.050 604.050 ;
        RECT 370.950 602.400 391.050 603.600 ;
        RECT 370.950 601.950 373.050 602.400 ;
        RECT 388.950 601.950 391.050 602.400 ;
        RECT 397.950 601.950 400.050 604.050 ;
        RECT 424.950 603.600 427.050 604.050 ;
        RECT 430.950 603.600 433.050 604.050 ;
        RECT 448.950 603.600 451.050 604.050 ;
        RECT 556.950 603.600 559.050 604.050 ;
        RECT 424.950 602.400 559.050 603.600 ;
        RECT 424.950 601.950 427.050 602.400 ;
        RECT 430.950 601.950 433.050 602.400 ;
        RECT 448.950 601.950 451.050 602.400 ;
        RECT 556.950 601.950 559.050 602.400 ;
        RECT 562.950 603.600 565.050 604.050 ;
        RECT 571.950 603.600 574.050 604.050 ;
        RECT 562.950 602.400 574.050 603.600 ;
        RECT 562.950 601.950 565.050 602.400 ;
        RECT 571.950 601.950 574.050 602.400 ;
        RECT 598.950 603.600 601.050 604.050 ;
        RECT 604.950 603.600 607.050 604.050 ;
        RECT 607.950 603.600 610.050 604.050 ;
        RECT 598.950 602.400 610.050 603.600 ;
        RECT 598.950 601.950 601.050 602.400 ;
        RECT 604.950 601.950 607.050 602.400 ;
        RECT 607.950 601.950 610.050 602.400 ;
        RECT 622.950 603.600 625.050 604.050 ;
        RECT 640.950 603.600 643.050 604.050 ;
        RECT 655.950 603.600 658.050 604.050 ;
        RECT 622.950 602.400 658.050 603.600 ;
        RECT 622.950 601.950 625.050 602.400 ;
        RECT 640.950 601.950 643.050 602.400 ;
        RECT 655.950 601.950 658.050 602.400 ;
        RECT 712.950 603.600 715.050 604.050 ;
        RECT 805.950 603.600 808.050 604.050 ;
        RECT 712.950 602.400 808.050 603.600 ;
        RECT 712.950 601.950 715.050 602.400 ;
        RECT 805.950 601.950 808.050 602.400 ;
        RECT 838.950 603.600 841.050 604.050 ;
        RECT 844.950 603.600 847.050 604.050 ;
        RECT 838.950 602.400 847.050 603.600 ;
        RECT 838.950 601.950 841.050 602.400 ;
        RECT 844.950 601.950 847.050 602.400 ;
        RECT 7.950 600.600 10.050 601.050 ;
        RECT 103.950 600.600 106.050 601.050 ;
        RECT 106.950 600.600 109.050 601.050 ;
        RECT 7.950 599.400 109.050 600.600 ;
        RECT 7.950 598.950 10.050 599.400 ;
        RECT 103.950 598.950 106.050 599.400 ;
        RECT 106.950 598.950 109.050 599.400 ;
        RECT 130.950 600.600 133.050 601.050 ;
        RECT 145.950 600.600 148.050 601.050 ;
        RECT 130.950 599.400 148.050 600.600 ;
        RECT 130.950 598.950 133.050 599.400 ;
        RECT 145.950 598.950 148.050 599.400 ;
        RECT 157.950 600.600 160.050 601.050 ;
        RECT 241.950 600.600 244.050 601.050 ;
        RECT 157.950 599.400 244.050 600.600 ;
        RECT 157.950 598.950 160.050 599.400 ;
        RECT 241.950 598.950 244.050 599.400 ;
        RECT 259.950 600.600 262.050 601.050 ;
        RECT 265.950 600.600 268.050 601.050 ;
        RECT 292.950 600.600 295.050 601.050 ;
        RECT 307.950 600.600 310.050 601.050 ;
        RECT 343.950 600.600 346.050 601.050 ;
        RECT 259.950 599.400 264.600 600.600 ;
        RECT 259.950 598.950 262.050 599.400 ;
        RECT 55.950 595.950 58.050 598.050 ;
        RECT 67.950 597.600 70.050 598.050 ;
        RECT 88.950 597.600 91.050 598.050 ;
        RECT 154.950 597.600 157.050 598.050 ;
        RECT 67.950 596.400 157.050 597.600 ;
        RECT 67.950 595.950 70.050 596.400 ;
        RECT 88.950 595.950 91.050 596.400 ;
        RECT 154.950 595.950 157.050 596.400 ;
        RECT 184.950 597.600 187.050 598.050 ;
        RECT 196.950 597.600 199.050 598.050 ;
        RECT 184.950 596.400 199.050 597.600 ;
        RECT 184.950 595.950 187.050 596.400 ;
        RECT 196.950 595.950 199.050 596.400 ;
        RECT 235.950 597.600 238.050 598.050 ;
        RECT 241.950 597.600 244.050 598.050 ;
        RECT 235.950 596.400 244.050 597.600 ;
        RECT 235.950 595.950 238.050 596.400 ;
        RECT 241.950 595.950 244.050 596.400 ;
        RECT 250.950 595.950 253.050 598.050 ;
        RECT 263.400 597.600 264.600 599.400 ;
        RECT 265.950 599.400 295.050 600.600 ;
        RECT 265.950 598.950 268.050 599.400 ;
        RECT 292.950 598.950 295.050 599.400 ;
        RECT 296.400 599.400 310.050 600.600 ;
        RECT 296.400 598.050 297.600 599.400 ;
        RECT 307.950 598.950 310.050 599.400 ;
        RECT 335.400 599.400 346.050 600.600 ;
        RECT 274.950 597.600 277.050 598.050 ;
        RECT 263.400 596.400 277.050 597.600 ;
        RECT 274.950 595.950 277.050 596.400 ;
        RECT 280.950 597.600 283.050 598.050 ;
        RECT 289.950 597.600 292.050 598.050 ;
        RECT 280.950 596.400 292.050 597.600 ;
        RECT 280.950 595.950 283.050 596.400 ;
        RECT 289.950 595.950 292.050 596.400 ;
        RECT 295.950 595.950 298.050 598.050 ;
        RECT 322.950 597.600 325.050 598.050 ;
        RECT 335.400 597.600 336.600 599.400 ;
        RECT 343.950 598.950 346.050 599.400 ;
        RECT 352.950 600.600 355.050 601.050 ;
        RECT 373.950 600.600 376.050 601.050 ;
        RECT 352.950 599.400 376.050 600.600 ;
        RECT 398.400 600.600 399.600 601.950 ;
        RECT 421.950 600.600 424.050 601.050 ;
        RECT 433.950 600.600 436.050 601.050 ;
        RECT 398.400 599.400 414.600 600.600 ;
        RECT 352.950 598.950 355.050 599.400 ;
        RECT 373.950 598.950 376.050 599.400 ;
        RECT 322.950 596.400 336.600 597.600 ;
        RECT 337.950 597.600 340.050 598.050 ;
        RECT 376.950 597.600 379.050 598.050 ;
        RECT 382.950 597.600 385.050 598.050 ;
        RECT 337.950 596.400 379.050 597.600 ;
        RECT 322.950 595.950 325.050 596.400 ;
        RECT 337.950 595.950 340.050 596.400 ;
        RECT 376.950 595.950 379.050 596.400 ;
        RECT 380.400 596.400 385.050 597.600 ;
        RECT 56.400 594.600 57.600 595.950 ;
        RECT 136.950 594.600 139.050 595.050 ;
        RECT 56.400 593.400 139.050 594.600 ;
        RECT 136.950 592.950 139.050 593.400 ;
        RECT 178.950 594.600 181.050 595.050 ;
        RECT 220.950 594.600 223.050 595.050 ;
        RECT 178.950 593.400 223.050 594.600 ;
        RECT 178.950 592.950 181.050 593.400 ;
        RECT 220.950 592.950 223.050 593.400 ;
        RECT 226.950 594.600 229.050 595.050 ;
        RECT 251.400 594.600 252.600 595.950 ;
        RECT 226.950 593.400 252.600 594.600 ;
        RECT 304.950 594.600 307.050 595.050 ;
        RECT 313.950 594.600 316.050 595.050 ;
        RECT 304.950 593.400 316.050 594.600 ;
        RECT 226.950 592.950 229.050 593.400 ;
        RECT 304.950 592.950 307.050 593.400 ;
        RECT 313.950 592.950 316.050 593.400 ;
        RECT 355.950 594.600 358.050 595.050 ;
        RECT 380.400 594.600 381.600 596.400 ;
        RECT 382.950 595.950 385.050 596.400 ;
        RECT 397.950 597.600 400.050 598.050 ;
        RECT 409.950 597.600 412.050 598.050 ;
        RECT 397.950 596.400 412.050 597.600 ;
        RECT 397.950 595.950 400.050 596.400 ;
        RECT 409.950 595.950 412.050 596.400 ;
        RECT 355.950 593.400 381.600 594.600 ;
        RECT 406.950 594.600 409.050 595.050 ;
        RECT 413.400 594.600 414.600 599.400 ;
        RECT 421.950 599.400 436.050 600.600 ;
        RECT 421.950 598.950 424.050 599.400 ;
        RECT 433.950 598.950 436.050 599.400 ;
        RECT 490.950 600.600 493.050 601.050 ;
        RECT 559.950 600.600 562.050 601.050 ;
        RECT 568.950 600.600 571.050 601.050 ;
        RECT 577.950 600.600 580.050 601.050 ;
        RECT 601.950 600.600 604.050 601.050 ;
        RECT 490.950 599.400 510.600 600.600 ;
        RECT 490.950 598.950 493.050 599.400 ;
        RECT 415.950 597.600 418.050 598.050 ;
        RECT 442.950 597.600 445.050 598.050 ;
        RECT 445.950 597.600 448.050 598.050 ;
        RECT 415.950 596.400 448.050 597.600 ;
        RECT 415.950 595.950 418.050 596.400 ;
        RECT 442.950 595.950 445.050 596.400 ;
        RECT 445.950 595.950 448.050 596.400 ;
        RECT 454.950 597.600 457.050 598.050 ;
        RECT 469.950 597.600 472.050 598.050 ;
        RECT 454.950 596.400 472.050 597.600 ;
        RECT 454.950 595.950 457.050 596.400 ;
        RECT 469.950 595.950 472.050 596.400 ;
        RECT 472.950 597.600 475.050 598.050 ;
        RECT 487.950 597.600 490.050 598.050 ;
        RECT 472.950 596.400 490.050 597.600 ;
        RECT 472.950 595.950 475.050 596.400 ;
        RECT 487.950 595.950 490.050 596.400 ;
        RECT 490.950 597.600 493.050 598.050 ;
        RECT 505.950 597.600 508.050 598.050 ;
        RECT 490.950 596.400 508.050 597.600 ;
        RECT 490.950 595.950 493.050 596.400 ;
        RECT 505.950 595.950 508.050 596.400 ;
        RECT 406.950 593.400 414.600 594.600 ;
        RECT 424.950 594.600 427.050 595.050 ;
        RECT 448.950 594.600 451.050 595.050 ;
        RECT 457.950 594.600 460.050 595.050 ;
        RECT 424.950 593.400 460.050 594.600 ;
        RECT 355.950 592.950 358.050 593.400 ;
        RECT 406.950 592.950 409.050 593.400 ;
        RECT 424.950 592.950 427.050 593.400 ;
        RECT 448.950 592.950 451.050 593.400 ;
        RECT 457.950 592.950 460.050 593.400 ;
        RECT 460.950 594.600 463.050 595.050 ;
        RECT 481.950 594.600 484.050 595.050 ;
        RECT 460.950 593.400 484.050 594.600 ;
        RECT 460.950 592.950 463.050 593.400 ;
        RECT 481.950 592.950 484.050 593.400 ;
        RECT 505.950 594.600 508.050 595.050 ;
        RECT 509.400 594.600 510.600 599.400 ;
        RECT 559.950 599.400 576.600 600.600 ;
        RECT 559.950 598.950 562.050 599.400 ;
        RECT 568.950 598.950 571.050 599.400 ;
        RECT 575.400 598.050 576.600 599.400 ;
        RECT 577.950 599.400 604.050 600.600 ;
        RECT 577.950 598.950 580.050 599.400 ;
        RECT 601.950 598.950 604.050 599.400 ;
        RECT 628.950 600.600 631.050 601.050 ;
        RECT 643.950 600.600 646.050 601.050 ;
        RECT 628.950 599.400 646.050 600.600 ;
        RECT 628.950 598.950 631.050 599.400 ;
        RECT 643.950 598.950 646.050 599.400 ;
        RECT 652.950 600.600 655.050 601.050 ;
        RECT 658.950 600.600 661.050 601.050 ;
        RECT 685.950 600.600 688.050 601.050 ;
        RECT 769.950 600.600 772.050 601.050 ;
        RECT 775.950 600.600 778.050 601.050 ;
        RECT 790.950 600.600 793.050 601.050 ;
        RECT 817.950 600.600 820.050 601.050 ;
        RECT 652.950 599.400 661.050 600.600 ;
        RECT 652.950 598.950 655.050 599.400 ;
        RECT 658.950 598.950 661.050 599.400 ;
        RECT 680.400 599.400 688.050 600.600 ;
        RECT 574.950 595.950 577.050 598.050 ;
        RECT 580.950 597.600 583.050 598.050 ;
        RECT 592.950 597.600 595.050 598.050 ;
        RECT 595.950 597.600 598.050 598.050 ;
        RECT 580.950 596.400 598.050 597.600 ;
        RECT 580.950 595.950 583.050 596.400 ;
        RECT 592.950 595.950 595.050 596.400 ;
        RECT 595.950 595.950 598.050 596.400 ;
        RECT 610.950 597.600 613.050 598.050 ;
        RECT 610.950 596.400 627.600 597.600 ;
        RECT 610.950 595.950 613.050 596.400 ;
        RECT 626.400 595.050 627.600 596.400 ;
        RECT 637.950 595.950 640.050 598.050 ;
        RECT 640.950 597.600 643.050 598.050 ;
        RECT 652.950 597.600 655.050 598.050 ;
        RECT 640.950 596.400 655.050 597.600 ;
        RECT 640.950 595.950 643.050 596.400 ;
        RECT 652.950 595.950 655.050 596.400 ;
        RECT 664.950 597.600 667.050 598.050 ;
        RECT 680.400 597.600 681.600 599.400 ;
        RECT 685.950 598.950 688.050 599.400 ;
        RECT 758.400 599.400 772.050 600.600 ;
        RECT 664.950 596.400 681.600 597.600 ;
        RECT 682.950 597.600 685.050 598.050 ;
        RECT 697.950 597.600 700.050 598.050 ;
        RECT 682.950 596.400 700.050 597.600 ;
        RECT 664.950 595.950 667.050 596.400 ;
        RECT 682.950 595.950 685.050 596.400 ;
        RECT 697.950 595.950 700.050 596.400 ;
        RECT 505.950 593.400 510.600 594.600 ;
        RECT 523.950 594.600 526.050 595.050 ;
        RECT 529.950 594.600 532.050 595.050 ;
        RECT 523.950 593.400 532.050 594.600 ;
        RECT 505.950 592.950 508.050 593.400 ;
        RECT 523.950 592.950 526.050 593.400 ;
        RECT 529.950 592.950 532.050 593.400 ;
        RECT 613.950 594.600 616.050 595.050 ;
        RECT 619.950 594.600 622.050 595.050 ;
        RECT 613.950 593.400 622.050 594.600 ;
        RECT 613.950 592.950 616.050 593.400 ;
        RECT 619.950 592.950 622.050 593.400 ;
        RECT 625.950 592.950 628.050 595.050 ;
        RECT 638.400 594.600 639.600 595.950 ;
        RECT 658.950 594.600 661.050 595.050 ;
        RECT 638.400 593.400 661.050 594.600 ;
        RECT 658.950 592.950 661.050 593.400 ;
        RECT 758.400 592.050 759.600 599.400 ;
        RECT 769.950 598.950 772.050 599.400 ;
        RECT 773.400 599.400 793.050 600.600 ;
        RECT 760.950 597.600 763.050 598.050 ;
        RECT 773.400 597.600 774.600 599.400 ;
        RECT 775.950 598.950 778.050 599.400 ;
        RECT 790.950 598.950 793.050 599.400 ;
        RECT 812.400 599.400 820.050 600.600 ;
        RECT 760.950 596.400 774.600 597.600 ;
        RECT 793.950 597.600 796.050 598.050 ;
        RECT 812.400 597.600 813.600 599.400 ;
        RECT 817.950 598.950 820.050 599.400 ;
        RECT 826.950 600.600 829.050 601.050 ;
        RECT 841.950 600.600 844.050 601.050 ;
        RECT 826.950 599.400 844.050 600.600 ;
        RECT 826.950 598.950 829.050 599.400 ;
        RECT 841.950 598.950 844.050 599.400 ;
        RECT 793.950 596.400 813.600 597.600 ;
        RECT 814.950 597.600 817.050 598.050 ;
        RECT 820.950 597.600 823.050 598.050 ;
        RECT 814.950 596.400 823.050 597.600 ;
        RECT 760.950 595.950 763.050 596.400 ;
        RECT 793.950 595.950 796.050 596.400 ;
        RECT 814.950 595.950 817.050 596.400 ;
        RECT 820.950 595.950 823.050 596.400 ;
        RECT 793.950 594.600 796.050 595.050 ;
        RECT 811.950 594.600 814.050 595.050 ;
        RECT 793.950 593.400 814.050 594.600 ;
        RECT 793.950 592.950 796.050 593.400 ;
        RECT 811.950 592.950 814.050 593.400 ;
        RECT 127.950 591.600 130.050 592.050 ;
        RECT 172.950 591.600 175.050 592.050 ;
        RECT 127.950 590.400 175.050 591.600 ;
        RECT 127.950 589.950 130.050 590.400 ;
        RECT 172.950 589.950 175.050 590.400 ;
        RECT 223.950 591.600 226.050 592.050 ;
        RECT 403.950 591.600 406.050 592.050 ;
        RECT 424.950 591.600 427.050 592.050 ;
        RECT 223.950 590.400 427.050 591.600 ;
        RECT 223.950 589.950 226.050 590.400 ;
        RECT 403.950 589.950 406.050 590.400 ;
        RECT 424.950 589.950 427.050 590.400 ;
        RECT 469.950 591.600 472.050 592.050 ;
        RECT 484.950 591.600 487.050 592.050 ;
        RECT 469.950 590.400 487.050 591.600 ;
        RECT 469.950 589.950 472.050 590.400 ;
        RECT 484.950 589.950 487.050 590.400 ;
        RECT 601.950 591.600 604.050 592.050 ;
        RECT 631.950 591.600 634.050 592.050 ;
        RECT 601.950 590.400 634.050 591.600 ;
        RECT 601.950 589.950 604.050 590.400 ;
        RECT 631.950 589.950 634.050 590.400 ;
        RECT 646.950 591.600 649.050 592.050 ;
        RECT 667.950 591.600 670.050 592.050 ;
        RECT 646.950 590.400 670.050 591.600 ;
        RECT 646.950 589.950 649.050 590.400 ;
        RECT 667.950 589.950 670.050 590.400 ;
        RECT 673.950 591.600 676.050 592.050 ;
        RECT 676.950 591.600 679.050 592.050 ;
        RECT 712.950 591.600 715.050 592.050 ;
        RECT 673.950 590.400 715.050 591.600 ;
        RECT 673.950 589.950 676.050 590.400 ;
        RECT 676.950 589.950 679.050 590.400 ;
        RECT 712.950 589.950 715.050 590.400 ;
        RECT 757.950 589.950 760.050 592.050 ;
        RECT 766.950 591.600 769.050 592.050 ;
        RECT 838.950 591.600 841.050 592.050 ;
        RECT 766.950 590.400 841.050 591.600 ;
        RECT 766.950 589.950 769.050 590.400 ;
        RECT 838.950 589.950 841.050 590.400 ;
        RECT 229.950 588.600 232.050 589.050 ;
        RECT 616.950 588.600 619.050 589.050 ;
        RECT 229.950 587.400 619.050 588.600 ;
        RECT 229.950 586.950 232.050 587.400 ;
        RECT 616.950 586.950 619.050 587.400 ;
        RECT 688.950 588.600 691.050 589.050 ;
        RECT 694.950 588.600 697.050 589.050 ;
        RECT 688.950 587.400 697.050 588.600 ;
        RECT 688.950 586.950 691.050 587.400 ;
        RECT 694.950 586.950 697.050 587.400 ;
        RECT 703.950 588.600 706.050 589.050 ;
        RECT 799.950 588.600 802.050 589.050 ;
        RECT 703.950 587.400 802.050 588.600 ;
        RECT 703.950 586.950 706.050 587.400 ;
        RECT 799.950 586.950 802.050 587.400 ;
        RECT 244.950 585.600 247.050 586.050 ;
        RECT 286.950 585.600 289.050 586.050 ;
        RECT 301.950 585.600 304.050 586.050 ;
        RECT 418.950 585.600 421.050 586.050 ;
        RECT 463.950 585.600 466.050 586.050 ;
        RECT 670.950 585.600 673.050 586.050 ;
        RECT 244.950 584.400 673.050 585.600 ;
        RECT 244.950 583.950 247.050 584.400 ;
        RECT 286.950 583.950 289.050 584.400 ;
        RECT 301.950 583.950 304.050 584.400 ;
        RECT 418.950 583.950 421.050 584.400 ;
        RECT 463.950 583.950 466.050 584.400 ;
        RECT 670.950 583.950 673.050 584.400 ;
        RECT 202.950 582.600 205.050 583.050 ;
        RECT 208.950 582.600 211.050 583.050 ;
        RECT 433.950 582.600 436.050 583.050 ;
        RECT 451.950 582.600 454.050 583.050 ;
        RECT 472.950 582.600 475.050 583.050 ;
        RECT 202.950 581.400 475.050 582.600 ;
        RECT 202.950 580.950 205.050 581.400 ;
        RECT 208.950 580.950 211.050 581.400 ;
        RECT 433.950 580.950 436.050 581.400 ;
        RECT 451.950 580.950 454.050 581.400 ;
        RECT 472.950 580.950 475.050 581.400 ;
        RECT 649.950 582.600 652.050 583.050 ;
        RECT 655.950 582.600 658.050 583.050 ;
        RECT 649.950 581.400 658.050 582.600 ;
        RECT 649.950 580.950 652.050 581.400 ;
        RECT 655.950 580.950 658.050 581.400 ;
        RECT 142.950 579.600 145.050 580.050 ;
        RECT 256.950 579.600 259.050 580.050 ;
        RECT 268.950 579.600 271.050 580.050 ;
        RECT 142.950 578.400 271.050 579.600 ;
        RECT 142.950 577.950 145.050 578.400 ;
        RECT 256.950 577.950 259.050 578.400 ;
        RECT 268.950 577.950 271.050 578.400 ;
        RECT 310.950 579.600 313.050 580.050 ;
        RECT 331.950 579.600 334.050 580.050 ;
        RECT 310.950 578.400 334.050 579.600 ;
        RECT 310.950 577.950 313.050 578.400 ;
        RECT 331.950 577.950 334.050 578.400 ;
        RECT 448.950 579.600 451.050 580.050 ;
        RECT 649.950 579.600 652.050 580.050 ;
        RECT 448.950 578.400 652.050 579.600 ;
        RECT 448.950 577.950 451.050 578.400 ;
        RECT 649.950 577.950 652.050 578.400 ;
        RECT 847.950 579.600 850.050 580.050 ;
        RECT 859.950 579.600 862.050 580.050 ;
        RECT 847.950 578.400 862.050 579.600 ;
        RECT 847.950 577.950 850.050 578.400 ;
        RECT 859.950 577.950 862.050 578.400 ;
        RECT 256.950 576.600 259.050 577.050 ;
        RECT 337.950 576.600 340.050 577.050 ;
        RECT 340.950 576.600 343.050 577.050 ;
        RECT 634.950 576.600 637.050 577.050 ;
        RECT 640.950 576.600 643.050 577.050 ;
        RECT 256.950 575.400 343.050 576.600 ;
        RECT 256.950 574.950 259.050 575.400 ;
        RECT 337.950 574.950 340.050 575.400 ;
        RECT 340.950 574.950 343.050 575.400 ;
        RECT 365.400 575.400 643.050 576.600 ;
        RECT 238.950 573.600 241.050 574.050 ;
        RECT 265.950 573.600 268.050 574.050 ;
        RECT 307.950 573.600 310.050 574.050 ;
        RECT 238.950 572.400 310.050 573.600 ;
        RECT 238.950 571.950 241.050 572.400 ;
        RECT 265.950 571.950 268.050 572.400 ;
        RECT 307.950 571.950 310.050 572.400 ;
        RECT 337.950 573.600 340.050 574.050 ;
        RECT 365.400 573.600 366.600 575.400 ;
        RECT 634.950 574.950 637.050 575.400 ;
        RECT 640.950 574.950 643.050 575.400 ;
        RECT 337.950 572.400 366.600 573.600 ;
        RECT 439.950 573.600 442.050 574.050 ;
        RECT 445.950 573.600 448.050 574.050 ;
        RECT 439.950 572.400 448.050 573.600 ;
        RECT 337.950 571.950 340.050 572.400 ;
        RECT 439.950 571.950 442.050 572.400 ;
        RECT 445.950 571.950 448.050 572.400 ;
        RECT 490.950 573.600 493.050 574.050 ;
        RECT 499.950 573.600 502.050 574.050 ;
        RECT 490.950 572.400 502.050 573.600 ;
        RECT 490.950 571.950 493.050 572.400 ;
        RECT 499.950 571.950 502.050 572.400 ;
        RECT 526.950 573.600 529.050 574.050 ;
        RECT 577.950 573.600 580.050 574.050 ;
        RECT 526.950 572.400 580.050 573.600 ;
        RECT 526.950 571.950 529.050 572.400 ;
        RECT 577.950 571.950 580.050 572.400 ;
        RECT 754.950 573.600 757.050 574.050 ;
        RECT 796.950 573.600 799.050 574.050 ;
        RECT 754.950 572.400 799.050 573.600 ;
        RECT 754.950 571.950 757.050 572.400 ;
        RECT 796.950 571.950 799.050 572.400 ;
        RECT 250.950 570.600 253.050 571.050 ;
        RECT 370.950 570.600 373.050 571.050 ;
        RECT 250.950 569.400 373.050 570.600 ;
        RECT 250.950 568.950 253.050 569.400 ;
        RECT 370.950 568.950 373.050 569.400 ;
        RECT 400.950 570.600 403.050 571.050 ;
        RECT 490.950 570.600 493.050 571.050 ;
        RECT 400.950 569.400 493.050 570.600 ;
        RECT 400.950 568.950 403.050 569.400 ;
        RECT 490.950 568.950 493.050 569.400 ;
        RECT 496.950 570.600 499.050 571.050 ;
        RECT 526.950 570.600 529.050 571.050 ;
        RECT 496.950 569.400 529.050 570.600 ;
        RECT 496.950 568.950 499.050 569.400 ;
        RECT 526.950 568.950 529.050 569.400 ;
        RECT 82.950 567.600 85.050 568.050 ;
        RECT 94.950 567.600 97.050 568.050 ;
        RECT 100.950 567.600 103.050 568.050 ;
        RECT 82.950 566.400 103.050 567.600 ;
        RECT 82.950 565.950 85.050 566.400 ;
        RECT 94.950 565.950 97.050 566.400 ;
        RECT 100.950 565.950 103.050 566.400 ;
        RECT 199.950 567.600 202.050 568.050 ;
        RECT 211.950 567.600 214.050 568.050 ;
        RECT 199.950 566.400 214.050 567.600 ;
        RECT 199.950 565.950 202.050 566.400 ;
        RECT 211.950 565.950 214.050 566.400 ;
        RECT 364.950 567.600 367.050 568.050 ;
        RECT 541.950 567.600 544.050 568.050 ;
        RECT 364.950 566.400 544.050 567.600 ;
        RECT 364.950 565.950 367.050 566.400 ;
        RECT 541.950 565.950 544.050 566.400 ;
        RECT 619.950 567.600 622.050 568.050 ;
        RECT 658.950 567.600 661.050 568.050 ;
        RECT 679.950 567.600 682.050 568.050 ;
        RECT 619.950 566.400 682.050 567.600 ;
        RECT 619.950 565.950 622.050 566.400 ;
        RECT 658.950 565.950 661.050 566.400 ;
        RECT 679.950 565.950 682.050 566.400 ;
        RECT 730.950 567.600 733.050 568.050 ;
        RECT 736.950 567.600 739.050 568.050 ;
        RECT 730.950 566.400 739.050 567.600 ;
        RECT 730.950 565.950 733.050 566.400 ;
        RECT 736.950 565.950 739.050 566.400 ;
        RECT 763.950 567.600 766.050 568.050 ;
        RECT 784.950 567.600 787.050 568.050 ;
        RECT 763.950 566.400 787.050 567.600 ;
        RECT 763.950 565.950 766.050 566.400 ;
        RECT 784.950 565.950 787.050 566.400 ;
        RECT 106.950 564.600 109.050 565.050 ;
        RECT 118.950 564.600 121.050 565.050 ;
        RECT 106.950 563.400 121.050 564.600 ;
        RECT 106.950 562.950 109.050 563.400 ;
        RECT 118.950 562.950 121.050 563.400 ;
        RECT 196.950 564.600 199.050 565.050 ;
        RECT 208.950 564.600 211.050 565.050 ;
        RECT 265.950 564.600 268.050 565.050 ;
        RECT 295.950 564.600 298.050 565.050 ;
        RECT 475.950 564.600 478.050 565.050 ;
        RECT 487.950 564.600 490.050 565.050 ;
        RECT 196.950 563.400 252.600 564.600 ;
        RECT 196.950 562.950 199.050 563.400 ;
        RECT 208.950 562.950 211.050 563.400 ;
        RECT 19.950 561.600 22.050 562.050 ;
        RECT 34.950 561.600 37.050 562.050 ;
        RECT 19.950 560.400 37.050 561.600 ;
        RECT 19.950 559.950 22.050 560.400 ;
        RECT 34.950 559.950 37.050 560.400 ;
        RECT 40.950 561.600 43.050 562.050 ;
        RECT 109.950 561.600 112.050 562.050 ;
        RECT 40.950 560.400 112.050 561.600 ;
        RECT 40.950 559.950 43.050 560.400 ;
        RECT 109.950 559.950 112.050 560.400 ;
        RECT 115.950 561.600 118.050 562.050 ;
        RECT 124.950 561.600 127.050 562.050 ;
        RECT 115.950 560.400 127.050 561.600 ;
        RECT 115.950 559.950 118.050 560.400 ;
        RECT 124.950 559.950 127.050 560.400 ;
        RECT 178.950 561.600 181.050 562.050 ;
        RECT 187.950 561.600 190.050 562.050 ;
        RECT 178.950 560.400 190.050 561.600 ;
        RECT 178.950 559.950 181.050 560.400 ;
        RECT 187.950 559.950 190.050 560.400 ;
        RECT 193.950 561.600 196.050 562.050 ;
        RECT 226.950 561.600 229.050 562.050 ;
        RECT 193.950 560.400 229.050 561.600 ;
        RECT 251.400 561.600 252.600 563.400 ;
        RECT 265.950 563.400 298.050 564.600 ;
        RECT 265.950 562.950 268.050 563.400 ;
        RECT 295.950 562.950 298.050 563.400 ;
        RECT 368.400 563.400 474.600 564.600 ;
        RECT 298.950 561.600 301.050 562.050 ;
        RECT 310.950 561.600 313.050 562.050 ;
        RECT 251.400 560.400 313.050 561.600 ;
        RECT 193.950 559.950 196.050 560.400 ;
        RECT 22.950 558.600 25.050 559.050 ;
        RECT 37.950 558.600 40.050 559.050 ;
        RECT 22.950 557.400 40.050 558.600 ;
        RECT 22.950 556.950 25.050 557.400 ;
        RECT 37.950 556.950 40.050 557.400 ;
        RECT 52.950 558.600 55.050 559.050 ;
        RECT 70.950 558.600 73.050 559.050 ;
        RECT 52.950 557.400 73.050 558.600 ;
        RECT 52.950 556.950 55.050 557.400 ;
        RECT 70.950 556.950 73.050 557.400 ;
        RECT 136.950 558.600 139.050 559.050 ;
        RECT 151.950 558.600 154.050 559.050 ;
        RECT 136.950 557.400 154.050 558.600 ;
        RECT 136.950 556.950 139.050 557.400 ;
        RECT 151.950 556.950 154.050 557.400 ;
        RECT 205.950 558.600 208.050 559.050 ;
        RECT 211.950 558.600 214.050 559.050 ;
        RECT 205.950 557.400 214.050 558.600 ;
        RECT 215.400 558.600 216.600 560.400 ;
        RECT 226.950 559.950 229.050 560.400 ;
        RECT 298.950 559.950 301.050 560.400 ;
        RECT 310.950 559.950 313.050 560.400 ;
        RECT 313.950 561.600 316.050 562.050 ;
        RECT 352.950 561.600 355.050 562.050 ;
        RECT 368.400 561.600 369.600 563.400 ;
        RECT 313.950 560.400 369.600 561.600 ;
        RECT 370.950 561.600 373.050 562.050 ;
        RECT 376.950 561.600 379.050 562.050 ;
        RECT 370.950 560.400 379.050 561.600 ;
        RECT 313.950 559.950 316.050 560.400 ;
        RECT 352.950 559.950 355.050 560.400 ;
        RECT 370.950 559.950 373.050 560.400 ;
        RECT 376.950 559.950 379.050 560.400 ;
        RECT 385.950 561.600 388.050 562.050 ;
        RECT 391.950 561.600 394.050 562.050 ;
        RECT 385.950 560.400 394.050 561.600 ;
        RECT 385.950 559.950 388.050 560.400 ;
        RECT 391.950 559.950 394.050 560.400 ;
        RECT 394.950 559.950 397.050 562.050 ;
        RECT 473.400 561.600 474.600 563.400 ;
        RECT 475.950 563.400 490.050 564.600 ;
        RECT 475.950 562.950 478.050 563.400 ;
        RECT 487.950 562.950 490.050 563.400 ;
        RECT 496.950 564.600 499.050 565.050 ;
        RECT 517.950 564.600 520.050 565.050 ;
        RECT 496.950 563.400 520.050 564.600 ;
        RECT 496.950 562.950 499.050 563.400 ;
        RECT 517.950 562.950 520.050 563.400 ;
        RECT 616.950 564.600 619.050 565.050 ;
        RECT 736.950 564.600 739.050 565.050 ;
        RECT 739.950 564.600 742.050 565.050 ;
        RECT 616.950 563.400 742.050 564.600 ;
        RECT 616.950 562.950 619.050 563.400 ;
        RECT 736.950 562.950 739.050 563.400 ;
        RECT 739.950 562.950 742.050 563.400 ;
        RECT 748.950 564.600 751.050 565.050 ;
        RECT 787.950 564.600 790.050 565.050 ;
        RECT 748.950 563.400 790.050 564.600 ;
        RECT 748.950 562.950 751.050 563.400 ;
        RECT 787.950 562.950 790.050 563.400 ;
        RECT 790.950 564.600 793.050 565.050 ;
        RECT 841.950 564.600 844.050 565.050 ;
        RECT 790.950 563.400 844.050 564.600 ;
        RECT 790.950 562.950 793.050 563.400 ;
        RECT 841.950 562.950 844.050 563.400 ;
        RECT 475.950 561.600 478.050 562.050 ;
        RECT 473.400 560.400 478.050 561.600 ;
        RECT 475.950 559.950 478.050 560.400 ;
        RECT 481.950 561.600 484.050 562.050 ;
        RECT 502.950 561.600 505.050 562.050 ;
        RECT 481.950 560.400 505.050 561.600 ;
        RECT 481.950 559.950 484.050 560.400 ;
        RECT 502.950 559.950 505.050 560.400 ;
        RECT 508.950 561.600 511.050 562.050 ;
        RECT 514.950 561.600 517.050 562.050 ;
        RECT 508.950 560.400 517.050 561.600 ;
        RECT 508.950 559.950 511.050 560.400 ;
        RECT 514.950 559.950 517.050 560.400 ;
        RECT 517.950 561.600 520.050 562.050 ;
        RECT 550.950 561.600 553.050 562.050 ;
        RECT 517.950 560.400 553.050 561.600 ;
        RECT 517.950 559.950 520.050 560.400 ;
        RECT 550.950 559.950 553.050 560.400 ;
        RECT 565.950 561.600 568.050 562.050 ;
        RECT 628.950 561.600 631.050 562.050 ;
        RECT 565.950 560.400 631.050 561.600 ;
        RECT 565.950 559.950 568.050 560.400 ;
        RECT 628.950 559.950 631.050 560.400 ;
        RECT 634.950 559.950 637.050 562.050 ;
        RECT 664.950 561.600 667.050 562.050 ;
        RECT 745.950 561.600 748.050 562.050 ;
        RECT 778.950 561.600 781.050 562.050 ;
        RECT 664.950 560.400 748.050 561.600 ;
        RECT 664.950 559.950 667.050 560.400 ;
        RECT 745.950 559.950 748.050 560.400 ;
        RECT 773.400 560.400 781.050 561.600 ;
        RECT 241.950 558.600 244.050 559.050 ;
        RECT 215.400 557.400 244.050 558.600 ;
        RECT 205.950 556.950 208.050 557.400 ;
        RECT 211.950 556.950 214.050 557.400 ;
        RECT 241.950 556.950 244.050 557.400 ;
        RECT 253.950 558.600 256.050 559.050 ;
        RECT 265.950 558.600 268.050 559.050 ;
        RECT 253.950 557.400 268.050 558.600 ;
        RECT 253.950 556.950 256.050 557.400 ;
        RECT 265.950 556.950 268.050 557.400 ;
        RECT 286.950 558.600 289.050 559.050 ;
        RECT 316.950 558.600 319.050 559.050 ;
        RECT 286.950 557.400 319.050 558.600 ;
        RECT 286.950 556.950 289.050 557.400 ;
        RECT 316.950 556.950 319.050 557.400 ;
        RECT 331.950 558.600 334.050 559.050 ;
        RECT 364.950 558.600 367.050 559.050 ;
        RECT 373.950 558.600 376.050 559.050 ;
        RECT 331.950 557.400 376.050 558.600 ;
        RECT 331.950 556.950 334.050 557.400 ;
        RECT 364.950 556.950 367.050 557.400 ;
        RECT 373.950 556.950 376.050 557.400 ;
        RECT 376.950 558.600 379.050 559.050 ;
        RECT 395.400 558.600 396.600 559.950 ;
        RECT 376.950 557.400 396.600 558.600 ;
        RECT 496.950 558.600 499.050 559.050 ;
        RECT 523.950 558.600 526.050 559.050 ;
        RECT 496.950 557.400 526.050 558.600 ;
        RECT 376.950 556.950 379.050 557.400 ;
        RECT 496.950 556.950 499.050 557.400 ;
        RECT 523.950 556.950 526.050 557.400 ;
        RECT 544.950 558.600 547.050 559.050 ;
        RECT 559.950 558.600 562.050 559.050 ;
        RECT 544.950 557.400 562.050 558.600 ;
        RECT 544.950 556.950 547.050 557.400 ;
        RECT 559.950 556.950 562.050 557.400 ;
        RECT 562.950 558.600 565.050 559.050 ;
        RECT 574.950 558.600 577.050 559.050 ;
        RECT 580.950 558.600 583.050 559.050 ;
        RECT 562.950 557.400 583.050 558.600 ;
        RECT 562.950 556.950 565.050 557.400 ;
        RECT 574.950 556.950 577.050 557.400 ;
        RECT 580.950 556.950 583.050 557.400 ;
        RECT 598.950 558.600 601.050 559.050 ;
        RECT 616.950 558.600 619.050 559.050 ;
        RECT 598.950 557.400 619.050 558.600 ;
        RECT 598.950 556.950 601.050 557.400 ;
        RECT 616.950 556.950 619.050 557.400 ;
        RECT 635.400 556.050 636.600 559.950 ;
        RECT 655.950 558.600 658.050 559.050 ;
        RECT 676.950 558.600 679.050 559.050 ;
        RECT 638.400 557.400 658.050 558.600 ;
        RECT 638.400 556.050 639.600 557.400 ;
        RECT 655.950 556.950 658.050 557.400 ;
        RECT 668.400 557.400 679.050 558.600 ;
        RECT 668.400 556.050 669.600 557.400 ;
        RECT 676.950 556.950 679.050 557.400 ;
        RECT 773.400 556.050 774.600 560.400 ;
        RECT 778.950 559.950 781.050 560.400 ;
        RECT 778.950 558.600 781.050 559.050 ;
        RECT 784.950 558.600 787.050 559.050 ;
        RECT 778.950 557.400 787.050 558.600 ;
        RECT 778.950 556.950 781.050 557.400 ;
        RECT 784.950 556.950 787.050 557.400 ;
        RECT 28.950 555.600 31.050 556.050 ;
        RECT 43.950 555.600 46.050 556.050 ;
        RECT 28.950 554.400 46.050 555.600 ;
        RECT 28.950 553.950 31.050 554.400 ;
        RECT 43.950 553.950 46.050 554.400 ;
        RECT 106.950 555.600 109.050 556.050 ;
        RECT 121.950 555.600 124.050 556.050 ;
        RECT 106.950 554.400 124.050 555.600 ;
        RECT 106.950 553.950 109.050 554.400 ;
        RECT 121.950 553.950 124.050 554.400 ;
        RECT 181.950 555.600 184.050 556.050 ;
        RECT 190.950 555.600 193.050 556.050 ;
        RECT 181.950 554.400 193.050 555.600 ;
        RECT 181.950 553.950 184.050 554.400 ;
        RECT 190.950 553.950 193.050 554.400 ;
        RECT 220.950 555.600 223.050 556.050 ;
        RECT 247.950 555.600 250.050 556.050 ;
        RECT 262.950 555.600 265.050 556.050 ;
        RECT 220.950 554.400 250.050 555.600 ;
        RECT 220.950 553.950 223.050 554.400 ;
        RECT 247.950 553.950 250.050 554.400 ;
        RECT 251.400 554.400 265.050 555.600 ;
        RECT 1.950 552.600 4.050 553.050 ;
        RECT 31.950 552.600 34.050 553.050 ;
        RECT 1.950 551.400 34.050 552.600 ;
        RECT 1.950 550.950 4.050 551.400 ;
        RECT 31.950 550.950 34.050 551.400 ;
        RECT 76.950 552.600 79.050 553.050 ;
        RECT 85.950 552.600 88.050 553.050 ;
        RECT 103.950 552.600 106.050 553.050 ;
        RECT 76.950 551.400 106.050 552.600 ;
        RECT 76.950 550.950 79.050 551.400 ;
        RECT 85.950 550.950 88.050 551.400 ;
        RECT 103.950 550.950 106.050 551.400 ;
        RECT 130.950 552.600 133.050 553.050 ;
        RECT 145.950 552.600 148.050 553.050 ;
        RECT 196.950 552.600 199.050 553.050 ;
        RECT 130.950 551.400 199.050 552.600 ;
        RECT 130.950 550.950 133.050 551.400 ;
        RECT 145.950 550.950 148.050 551.400 ;
        RECT 196.950 550.950 199.050 551.400 ;
        RECT 235.950 552.600 238.050 553.050 ;
        RECT 251.400 552.600 252.600 554.400 ;
        RECT 262.950 553.950 265.050 554.400 ;
        RECT 268.950 555.600 271.050 556.050 ;
        RECT 277.950 555.600 280.050 556.050 ;
        RECT 268.950 554.400 280.050 555.600 ;
        RECT 268.950 553.950 271.050 554.400 ;
        RECT 277.950 553.950 280.050 554.400 ;
        RECT 307.950 555.600 310.050 556.050 ;
        RECT 313.950 555.600 316.050 556.050 ;
        RECT 307.950 554.400 316.050 555.600 ;
        RECT 307.950 553.950 310.050 554.400 ;
        RECT 313.950 553.950 316.050 554.400 ;
        RECT 343.950 555.600 346.050 556.050 ;
        RECT 352.950 555.600 355.050 556.050 ;
        RECT 343.950 554.400 355.050 555.600 ;
        RECT 343.950 553.950 346.050 554.400 ;
        RECT 352.950 553.950 355.050 554.400 ;
        RECT 355.950 555.600 358.050 556.050 ;
        RECT 373.950 555.600 376.050 556.050 ;
        RECT 379.950 555.600 382.050 556.050 ;
        RECT 355.950 554.400 382.050 555.600 ;
        RECT 355.950 553.950 358.050 554.400 ;
        RECT 373.950 553.950 376.050 554.400 ;
        RECT 379.950 553.950 382.050 554.400 ;
        RECT 484.950 555.600 487.050 556.050 ;
        RECT 514.950 555.600 517.050 556.050 ;
        RECT 484.950 554.400 517.050 555.600 ;
        RECT 484.950 553.950 487.050 554.400 ;
        RECT 514.950 553.950 517.050 554.400 ;
        RECT 520.950 555.600 523.050 556.050 ;
        RECT 532.950 555.600 535.050 556.050 ;
        RECT 520.950 554.400 535.050 555.600 ;
        RECT 520.950 553.950 523.050 554.400 ;
        RECT 532.950 553.950 535.050 554.400 ;
        RECT 538.950 555.600 541.050 556.050 ;
        RECT 586.950 555.600 589.050 556.050 ;
        RECT 538.950 554.400 589.050 555.600 ;
        RECT 538.950 553.950 541.050 554.400 ;
        RECT 586.950 553.950 589.050 554.400 ;
        RECT 595.950 555.600 598.050 556.050 ;
        RECT 604.950 555.600 607.050 556.050 ;
        RECT 595.950 554.400 607.050 555.600 ;
        RECT 595.950 553.950 598.050 554.400 ;
        RECT 604.950 553.950 607.050 554.400 ;
        RECT 613.950 555.600 616.050 556.050 ;
        RECT 625.950 555.600 628.050 556.050 ;
        RECT 613.950 554.400 628.050 555.600 ;
        RECT 613.950 553.950 616.050 554.400 ;
        RECT 625.950 553.950 628.050 554.400 ;
        RECT 634.950 553.950 637.050 556.050 ;
        RECT 637.950 553.950 640.050 556.050 ;
        RECT 643.950 555.600 646.050 556.050 ;
        RECT 658.950 555.600 661.050 556.050 ;
        RECT 643.950 554.400 661.050 555.600 ;
        RECT 643.950 553.950 646.050 554.400 ;
        RECT 658.950 553.950 661.050 554.400 ;
        RECT 667.950 553.950 670.050 556.050 ;
        RECT 733.950 555.600 736.050 556.050 ;
        RECT 742.950 555.600 745.050 556.050 ;
        RECT 733.950 554.400 745.050 555.600 ;
        RECT 733.950 553.950 736.050 554.400 ;
        RECT 742.950 553.950 745.050 554.400 ;
        RECT 751.950 555.600 754.050 556.050 ;
        RECT 766.950 555.600 769.050 556.050 ;
        RECT 751.950 554.400 769.050 555.600 ;
        RECT 751.950 553.950 754.050 554.400 ;
        RECT 766.950 553.950 769.050 554.400 ;
        RECT 772.950 553.950 775.050 556.050 ;
        RECT 235.950 551.400 252.600 552.600 ;
        RECT 253.950 552.600 256.050 553.050 ;
        RECT 259.950 552.600 262.050 553.050 ;
        RECT 253.950 551.400 262.050 552.600 ;
        RECT 235.950 550.950 238.050 551.400 ;
        RECT 253.950 550.950 256.050 551.400 ;
        RECT 259.950 550.950 262.050 551.400 ;
        RECT 301.950 552.600 304.050 553.050 ;
        RECT 307.950 552.600 310.050 553.050 ;
        RECT 301.950 551.400 310.050 552.600 ;
        RECT 301.950 550.950 304.050 551.400 ;
        RECT 307.950 550.950 310.050 551.400 ;
        RECT 328.950 552.600 331.050 553.050 ;
        RECT 346.950 552.600 349.050 553.050 ;
        RECT 328.950 551.400 349.050 552.600 ;
        RECT 328.950 550.950 331.050 551.400 ;
        RECT 346.950 550.950 349.050 551.400 ;
        RECT 367.950 552.600 370.050 553.050 ;
        RECT 400.950 552.600 403.050 553.050 ;
        RECT 367.950 551.400 403.050 552.600 ;
        RECT 367.950 550.950 370.050 551.400 ;
        RECT 400.950 550.950 403.050 551.400 ;
        RECT 460.950 552.600 463.050 553.050 ;
        RECT 472.950 552.600 475.050 553.050 ;
        RECT 460.950 551.400 475.050 552.600 ;
        RECT 460.950 550.950 463.050 551.400 ;
        RECT 472.950 550.950 475.050 551.400 ;
        RECT 523.950 552.600 526.050 553.050 ;
        RECT 565.950 552.600 568.050 553.050 ;
        RECT 523.950 551.400 568.050 552.600 ;
        RECT 523.950 550.950 526.050 551.400 ;
        RECT 565.950 550.950 568.050 551.400 ;
        RECT 574.950 552.600 577.050 553.050 ;
        RECT 610.950 552.600 613.050 553.050 ;
        RECT 574.950 551.400 613.050 552.600 ;
        RECT 574.950 550.950 577.050 551.400 ;
        RECT 610.950 550.950 613.050 551.400 ;
        RECT 613.950 552.600 616.050 553.050 ;
        RECT 688.950 552.600 691.050 553.050 ;
        RECT 613.950 551.400 691.050 552.600 ;
        RECT 613.950 550.950 616.050 551.400 ;
        RECT 688.950 550.950 691.050 551.400 ;
        RECT 751.950 552.600 754.050 553.050 ;
        RECT 757.950 552.600 760.050 553.050 ;
        RECT 751.950 551.400 760.050 552.600 ;
        RECT 751.950 550.950 754.050 551.400 ;
        RECT 757.950 550.950 760.050 551.400 ;
        RECT 31.950 549.600 34.050 550.050 ;
        RECT 103.950 549.600 106.050 550.050 ;
        RECT 31.950 548.400 106.050 549.600 ;
        RECT 31.950 547.950 34.050 548.400 ;
        RECT 103.950 547.950 106.050 548.400 ;
        RECT 160.950 549.600 163.050 550.050 ;
        RECT 181.950 549.600 184.050 550.050 ;
        RECT 160.950 548.400 184.050 549.600 ;
        RECT 160.950 547.950 163.050 548.400 ;
        RECT 181.950 547.950 184.050 548.400 ;
        RECT 226.950 549.600 229.050 550.050 ;
        RECT 271.950 549.600 274.050 550.050 ;
        RECT 451.950 549.600 454.050 550.050 ;
        RECT 226.950 548.400 454.050 549.600 ;
        RECT 226.950 547.950 229.050 548.400 ;
        RECT 271.950 547.950 274.050 548.400 ;
        RECT 451.950 547.950 454.050 548.400 ;
        RECT 631.950 549.600 634.050 550.050 ;
        RECT 652.950 549.600 655.050 550.050 ;
        RECT 631.950 548.400 655.050 549.600 ;
        RECT 631.950 547.950 634.050 548.400 ;
        RECT 652.950 547.950 655.050 548.400 ;
        RECT 685.950 549.600 688.050 550.050 ;
        RECT 754.950 549.600 757.050 550.050 ;
        RECT 685.950 548.400 757.050 549.600 ;
        RECT 685.950 547.950 688.050 548.400 ;
        RECT 754.950 547.950 757.050 548.400 ;
        RECT 100.950 546.600 103.050 547.050 ;
        RECT 112.950 546.600 115.050 547.050 ;
        RECT 100.950 545.400 115.050 546.600 ;
        RECT 100.950 544.950 103.050 545.400 ;
        RECT 112.950 544.950 115.050 545.400 ;
        RECT 163.950 546.600 166.050 547.050 ;
        RECT 187.950 546.600 190.050 547.050 ;
        RECT 235.950 546.600 238.050 547.050 ;
        RECT 163.950 545.400 238.050 546.600 ;
        RECT 163.950 544.950 166.050 545.400 ;
        RECT 187.950 544.950 190.050 545.400 ;
        RECT 235.950 544.950 238.050 545.400 ;
        RECT 238.950 546.600 241.050 547.050 ;
        RECT 355.950 546.600 358.050 547.050 ;
        RECT 238.950 545.400 358.050 546.600 ;
        RECT 238.950 544.950 241.050 545.400 ;
        RECT 355.950 544.950 358.050 545.400 ;
        RECT 403.950 546.600 406.050 547.050 ;
        RECT 442.950 546.600 445.050 547.050 ;
        RECT 403.950 545.400 445.050 546.600 ;
        RECT 403.950 544.950 406.050 545.400 ;
        RECT 442.950 544.950 445.050 545.400 ;
        RECT 472.950 546.600 475.050 547.050 ;
        RECT 580.950 546.600 583.050 547.050 ;
        RECT 613.950 546.600 616.050 547.050 ;
        RECT 472.950 545.400 616.050 546.600 ;
        RECT 472.950 544.950 475.050 545.400 ;
        RECT 580.950 544.950 583.050 545.400 ;
        RECT 613.950 544.950 616.050 545.400 ;
        RECT 634.950 546.600 637.050 547.050 ;
        RECT 646.950 546.600 649.050 547.050 ;
        RECT 634.950 545.400 649.050 546.600 ;
        RECT 634.950 544.950 637.050 545.400 ;
        RECT 646.950 544.950 649.050 545.400 ;
        RECT 649.950 546.600 652.050 547.050 ;
        RECT 655.950 546.600 658.050 547.050 ;
        RECT 682.950 546.600 685.050 547.050 ;
        RECT 649.950 545.400 685.050 546.600 ;
        RECT 649.950 544.950 652.050 545.400 ;
        RECT 655.950 544.950 658.050 545.400 ;
        RECT 682.950 544.950 685.050 545.400 ;
        RECT 748.950 546.600 751.050 547.050 ;
        RECT 817.950 546.600 820.050 547.050 ;
        RECT 748.950 545.400 820.050 546.600 ;
        RECT 748.950 544.950 751.050 545.400 ;
        RECT 817.950 544.950 820.050 545.400 ;
        RECT 7.950 543.600 10.050 544.050 ;
        RECT 16.950 543.600 19.050 544.050 ;
        RECT 127.950 543.600 130.050 544.050 ;
        RECT 7.950 542.400 130.050 543.600 ;
        RECT 7.950 541.950 10.050 542.400 ;
        RECT 16.950 541.950 19.050 542.400 ;
        RECT 127.950 541.950 130.050 542.400 ;
        RECT 169.950 543.600 172.050 544.050 ;
        RECT 253.950 543.600 256.050 544.050 ;
        RECT 169.950 542.400 256.050 543.600 ;
        RECT 169.950 541.950 172.050 542.400 ;
        RECT 253.950 541.950 256.050 542.400 ;
        RECT 265.950 543.600 268.050 544.050 ;
        RECT 328.950 543.600 331.050 544.050 ;
        RECT 265.950 542.400 331.050 543.600 ;
        RECT 265.950 541.950 268.050 542.400 ;
        RECT 328.950 541.950 331.050 542.400 ;
        RECT 343.950 543.600 346.050 544.050 ;
        RECT 358.950 543.600 361.050 544.050 ;
        RECT 343.950 542.400 361.050 543.600 ;
        RECT 343.950 541.950 346.050 542.400 ;
        RECT 358.950 541.950 361.050 542.400 ;
        RECT 493.950 543.600 496.050 544.050 ;
        RECT 499.950 543.600 502.050 544.050 ;
        RECT 493.950 542.400 502.050 543.600 ;
        RECT 493.950 541.950 496.050 542.400 ;
        RECT 499.950 541.950 502.050 542.400 ;
        RECT 535.950 543.600 538.050 544.050 ;
        RECT 568.950 543.600 571.050 544.050 ;
        RECT 535.950 542.400 571.050 543.600 ;
        RECT 535.950 541.950 538.050 542.400 ;
        RECT 568.950 541.950 571.050 542.400 ;
        RECT 625.950 543.600 628.050 544.050 ;
        RECT 658.950 543.600 661.050 544.050 ;
        RECT 625.950 542.400 661.050 543.600 ;
        RECT 625.950 541.950 628.050 542.400 ;
        RECT 658.950 541.950 661.050 542.400 ;
        RECT 97.950 540.600 100.050 541.050 ;
        RECT 256.950 540.600 259.050 541.050 ;
        RECT 97.950 539.400 259.050 540.600 ;
        RECT 97.950 538.950 100.050 539.400 ;
        RECT 256.950 538.950 259.050 539.400 ;
        RECT 298.950 540.600 301.050 541.050 ;
        RECT 361.950 540.600 364.050 541.050 ;
        RECT 298.950 539.400 364.050 540.600 ;
        RECT 298.950 538.950 301.050 539.400 ;
        RECT 361.950 538.950 364.050 539.400 ;
        RECT 466.950 540.600 469.050 541.050 ;
        RECT 475.950 540.600 478.050 541.050 ;
        RECT 466.950 539.400 478.050 540.600 ;
        RECT 466.950 538.950 469.050 539.400 ;
        RECT 475.950 538.950 478.050 539.400 ;
        RECT 487.950 540.600 490.050 541.050 ;
        RECT 514.950 540.600 517.050 541.050 ;
        RECT 487.950 539.400 517.050 540.600 ;
        RECT 487.950 538.950 490.050 539.400 ;
        RECT 514.950 538.950 517.050 539.400 ;
        RECT 541.950 540.600 544.050 541.050 ;
        RECT 559.950 540.600 562.050 541.050 ;
        RECT 541.950 539.400 562.050 540.600 ;
        RECT 541.950 538.950 544.050 539.400 ;
        RECT 559.950 538.950 562.050 539.400 ;
        RECT 583.950 540.600 586.050 541.050 ;
        RECT 601.950 540.600 604.050 541.050 ;
        RECT 649.950 540.600 652.050 541.050 ;
        RECT 583.950 539.400 652.050 540.600 ;
        RECT 583.950 538.950 586.050 539.400 ;
        RECT 601.950 538.950 604.050 539.400 ;
        RECT 649.950 538.950 652.050 539.400 ;
        RECT 199.950 537.600 202.050 538.050 ;
        RECT 250.950 537.600 253.050 538.050 ;
        RECT 199.950 536.400 253.050 537.600 ;
        RECT 199.950 535.950 202.050 536.400 ;
        RECT 250.950 535.950 253.050 536.400 ;
        RECT 280.950 537.600 283.050 538.050 ;
        RECT 304.950 537.600 307.050 538.050 ;
        RECT 280.950 536.400 307.050 537.600 ;
        RECT 280.950 535.950 283.050 536.400 ;
        RECT 304.950 535.950 307.050 536.400 ;
        RECT 316.950 537.600 319.050 538.050 ;
        RECT 325.950 537.600 328.050 538.050 ;
        RECT 316.950 536.400 328.050 537.600 ;
        RECT 316.950 535.950 319.050 536.400 ;
        RECT 325.950 535.950 328.050 536.400 ;
        RECT 328.950 537.600 331.050 538.050 ;
        RECT 364.950 537.600 367.050 538.050 ;
        RECT 388.950 537.600 391.050 538.050 ;
        RECT 328.950 536.400 363.600 537.600 ;
        RECT 328.950 535.950 331.050 536.400 ;
        RECT 55.950 534.600 58.050 535.050 ;
        RECT 160.950 534.600 163.050 535.050 ;
        RECT 55.950 533.400 163.050 534.600 ;
        RECT 55.950 532.950 58.050 533.400 ;
        RECT 160.950 532.950 163.050 533.400 ;
        RECT 220.950 534.600 223.050 535.050 ;
        RECT 238.950 534.600 241.050 535.050 ;
        RECT 220.950 533.400 241.050 534.600 ;
        RECT 220.950 532.950 223.050 533.400 ;
        RECT 238.950 532.950 241.050 533.400 ;
        RECT 280.950 534.600 283.050 535.050 ;
        RECT 331.950 534.600 334.050 535.050 ;
        RECT 280.950 533.400 334.050 534.600 ;
        RECT 280.950 532.950 283.050 533.400 ;
        RECT 331.950 532.950 334.050 533.400 ;
        RECT 352.950 534.600 355.050 535.050 ;
        RECT 358.950 534.600 361.050 535.050 ;
        RECT 352.950 533.400 361.050 534.600 ;
        RECT 362.400 534.600 363.600 536.400 ;
        RECT 364.950 536.400 391.050 537.600 ;
        RECT 364.950 535.950 367.050 536.400 ;
        RECT 388.950 535.950 391.050 536.400 ;
        RECT 478.950 537.600 481.050 538.050 ;
        RECT 499.950 537.600 502.050 538.050 ;
        RECT 478.950 536.400 502.050 537.600 ;
        RECT 478.950 535.950 481.050 536.400 ;
        RECT 499.950 535.950 502.050 536.400 ;
        RECT 547.950 537.600 550.050 538.050 ;
        RECT 616.950 537.600 619.050 538.050 ;
        RECT 640.950 537.600 643.050 538.050 ;
        RECT 547.950 536.400 643.050 537.600 ;
        RECT 547.950 535.950 550.050 536.400 ;
        RECT 616.950 535.950 619.050 536.400 ;
        RECT 640.950 535.950 643.050 536.400 ;
        RECT 367.950 534.600 370.050 535.050 ;
        RECT 362.400 533.400 370.050 534.600 ;
        RECT 352.950 532.950 355.050 533.400 ;
        RECT 358.950 532.950 361.050 533.400 ;
        RECT 367.950 532.950 370.050 533.400 ;
        RECT 379.950 534.600 382.050 535.050 ;
        RECT 385.950 534.600 388.050 535.050 ;
        RECT 379.950 533.400 388.050 534.600 ;
        RECT 379.950 532.950 382.050 533.400 ;
        RECT 385.950 532.950 388.050 533.400 ;
        RECT 415.950 534.600 418.050 535.050 ;
        RECT 427.950 534.600 430.050 535.050 ;
        RECT 415.950 533.400 430.050 534.600 ;
        RECT 415.950 532.950 418.050 533.400 ;
        RECT 427.950 532.950 430.050 533.400 ;
        RECT 508.950 534.600 511.050 535.050 ;
        RECT 529.950 534.600 532.050 535.050 ;
        RECT 508.950 533.400 532.050 534.600 ;
        RECT 508.950 532.950 511.050 533.400 ;
        RECT 529.950 532.950 532.050 533.400 ;
        RECT 556.950 534.600 559.050 535.050 ;
        RECT 589.950 534.600 592.050 535.050 ;
        RECT 625.950 534.600 628.050 535.050 ;
        RECT 556.950 533.400 628.050 534.600 ;
        RECT 556.950 532.950 559.050 533.400 ;
        RECT 589.950 532.950 592.050 533.400 ;
        RECT 625.950 532.950 628.050 533.400 ;
        RECT 25.950 531.600 28.050 532.050 ;
        RECT 43.950 531.600 46.050 532.050 ;
        RECT 25.950 530.400 46.050 531.600 ;
        RECT 25.950 529.950 28.050 530.400 ;
        RECT 43.950 529.950 46.050 530.400 ;
        RECT 91.950 531.600 94.050 532.050 ;
        RECT 172.950 531.600 175.050 532.050 ;
        RECT 190.950 531.600 193.050 532.050 ;
        RECT 193.950 531.600 196.050 532.050 ;
        RECT 91.950 530.400 147.600 531.600 ;
        RECT 91.950 529.950 94.050 530.400 ;
        RECT 10.950 528.600 13.050 529.050 ;
        RECT 28.950 528.600 31.050 529.050 ;
        RECT 85.950 528.600 88.050 529.050 ;
        RECT 88.950 528.600 91.050 529.050 ;
        RECT 10.950 527.400 91.050 528.600 ;
        RECT 10.950 526.950 13.050 527.400 ;
        RECT 28.950 526.950 31.050 527.400 ;
        RECT 85.950 526.950 88.050 527.400 ;
        RECT 88.950 526.950 91.050 527.400 ;
        RECT 109.950 528.600 112.050 529.050 ;
        RECT 109.950 527.400 141.600 528.600 ;
        RECT 109.950 526.950 112.050 527.400 ;
        RECT 140.400 526.050 141.600 527.400 ;
        RECT 146.400 526.050 147.600 530.400 ;
        RECT 172.950 530.400 196.050 531.600 ;
        RECT 172.950 529.950 175.050 530.400 ;
        RECT 190.950 529.950 193.050 530.400 ;
        RECT 193.950 529.950 196.050 530.400 ;
        RECT 214.950 531.600 217.050 532.050 ;
        RECT 226.950 531.600 229.050 532.050 ;
        RECT 214.950 530.400 229.050 531.600 ;
        RECT 214.950 529.950 217.050 530.400 ;
        RECT 226.950 529.950 229.050 530.400 ;
        RECT 244.950 531.600 247.050 532.050 ;
        RECT 259.950 531.600 262.050 532.050 ;
        RECT 244.950 530.400 262.050 531.600 ;
        RECT 244.950 529.950 247.050 530.400 ;
        RECT 259.950 529.950 262.050 530.400 ;
        RECT 265.950 531.600 268.050 532.050 ;
        RECT 271.950 531.600 274.050 532.050 ;
        RECT 265.950 530.400 274.050 531.600 ;
        RECT 265.950 529.950 268.050 530.400 ;
        RECT 271.950 529.950 274.050 530.400 ;
        RECT 274.950 531.600 277.050 532.050 ;
        RECT 382.950 531.600 385.050 532.050 ;
        RECT 274.950 530.400 385.050 531.600 ;
        RECT 274.950 529.950 277.050 530.400 ;
        RECT 382.950 529.950 385.050 530.400 ;
        RECT 388.950 529.950 391.050 532.050 ;
        RECT 403.950 531.600 406.050 532.050 ;
        RECT 472.950 531.600 475.050 532.050 ;
        RECT 403.950 530.400 475.050 531.600 ;
        RECT 403.950 529.950 406.050 530.400 ;
        RECT 472.950 529.950 475.050 530.400 ;
        RECT 487.950 531.600 490.050 532.050 ;
        RECT 502.950 531.600 505.050 532.050 ;
        RECT 487.950 530.400 505.050 531.600 ;
        RECT 487.950 529.950 490.050 530.400 ;
        RECT 502.950 529.950 505.050 530.400 ;
        RECT 511.950 531.600 514.050 532.050 ;
        RECT 541.950 531.600 544.050 532.050 ;
        RECT 511.950 530.400 544.050 531.600 ;
        RECT 511.950 529.950 514.050 530.400 ;
        RECT 541.950 529.950 544.050 530.400 ;
        RECT 553.950 531.600 556.050 532.050 ;
        RECT 562.950 531.600 565.050 532.050 ;
        RECT 571.950 531.600 574.050 532.050 ;
        RECT 553.950 530.400 574.050 531.600 ;
        RECT 553.950 529.950 556.050 530.400 ;
        RECT 562.950 529.950 565.050 530.400 ;
        RECT 571.950 529.950 574.050 530.400 ;
        RECT 595.950 531.600 598.050 532.050 ;
        RECT 619.950 531.600 622.050 532.050 ;
        RECT 595.950 530.400 622.050 531.600 ;
        RECT 595.950 529.950 598.050 530.400 ;
        RECT 619.950 529.950 622.050 530.400 ;
        RECT 661.950 531.600 664.050 532.050 ;
        RECT 724.950 531.600 727.050 532.050 ;
        RECT 661.950 530.400 727.050 531.600 ;
        RECT 661.950 529.950 664.050 530.400 ;
        RECT 724.950 529.950 727.050 530.400 ;
        RECT 778.950 531.600 781.050 532.050 ;
        RECT 829.950 531.600 832.050 532.050 ;
        RECT 847.950 531.600 850.050 532.050 ;
        RECT 778.950 530.400 832.050 531.600 ;
        RECT 778.950 529.950 781.050 530.400 ;
        RECT 829.950 529.950 832.050 530.400 ;
        RECT 842.400 530.400 850.050 531.600 ;
        RECT 148.950 528.600 151.050 529.050 ;
        RECT 163.950 528.600 166.050 529.050 ;
        RECT 148.950 527.400 166.050 528.600 ;
        RECT 148.950 526.950 151.050 527.400 ;
        RECT 163.950 526.950 166.050 527.400 ;
        RECT 184.950 528.600 187.050 529.050 ;
        RECT 247.950 528.600 250.050 529.050 ;
        RECT 184.950 527.400 250.050 528.600 ;
        RECT 184.950 526.950 187.050 527.400 ;
        RECT 247.950 526.950 250.050 527.400 ;
        RECT 274.950 528.600 277.050 529.050 ;
        RECT 292.950 528.600 295.050 529.050 ;
        RECT 274.950 527.400 295.050 528.600 ;
        RECT 274.950 526.950 277.050 527.400 ;
        RECT 292.950 526.950 295.050 527.400 ;
        RECT 295.950 528.600 298.050 529.050 ;
        RECT 322.950 528.600 325.050 529.050 ;
        RECT 295.950 527.400 325.050 528.600 ;
        RECT 295.950 526.950 298.050 527.400 ;
        RECT 322.950 526.950 325.050 527.400 ;
        RECT 325.950 528.600 328.050 529.050 ;
        RECT 346.950 528.600 349.050 529.050 ;
        RECT 325.950 527.400 349.050 528.600 ;
        RECT 325.950 526.950 328.050 527.400 ;
        RECT 346.950 526.950 349.050 527.400 ;
        RECT 370.950 528.600 373.050 529.050 ;
        RECT 389.400 528.600 390.600 529.950 ;
        RECT 370.950 527.400 390.600 528.600 ;
        RECT 370.950 526.950 373.050 527.400 ;
        RECT 397.950 526.950 400.050 529.050 ;
        RECT 406.950 528.600 409.050 529.050 ;
        RECT 421.950 528.600 424.050 529.050 ;
        RECT 406.950 527.400 424.050 528.600 ;
        RECT 406.950 526.950 409.050 527.400 ;
        RECT 421.950 526.950 424.050 527.400 ;
        RECT 445.950 528.600 448.050 529.050 ;
        RECT 532.950 528.600 535.050 529.050 ;
        RECT 445.950 527.400 535.050 528.600 ;
        RECT 445.950 526.950 448.050 527.400 ;
        RECT 532.950 526.950 535.050 527.400 ;
        RECT 553.950 526.950 556.050 529.050 ;
        RECT 598.950 526.950 601.050 529.050 ;
        RECT 604.950 528.600 607.050 529.050 ;
        RECT 673.950 528.600 676.050 529.050 ;
        RECT 688.950 528.600 691.050 529.050 ;
        RECT 604.950 527.400 691.050 528.600 ;
        RECT 604.950 526.950 607.050 527.400 ;
        RECT 673.950 526.950 676.050 527.400 ;
        RECT 688.950 526.950 691.050 527.400 ;
        RECT 763.950 528.600 766.050 529.050 ;
        RECT 787.950 528.600 790.050 529.050 ;
        RECT 763.950 527.400 790.050 528.600 ;
        RECT 763.950 526.950 766.050 527.400 ;
        RECT 787.950 526.950 790.050 527.400 ;
        RECT 16.950 525.600 19.050 526.050 ;
        RECT 22.950 525.600 25.050 526.050 ;
        RECT 16.950 524.400 25.050 525.600 ;
        RECT 16.950 523.950 19.050 524.400 ;
        RECT 22.950 523.950 25.050 524.400 ;
        RECT 37.950 525.600 40.050 526.050 ;
        RECT 55.950 525.600 58.050 526.050 ;
        RECT 37.950 524.400 58.050 525.600 ;
        RECT 37.950 523.950 40.050 524.400 ;
        RECT 55.950 523.950 58.050 524.400 ;
        RECT 61.950 525.600 64.050 526.050 ;
        RECT 76.950 525.600 79.050 526.050 ;
        RECT 82.950 525.600 85.050 526.050 ;
        RECT 61.950 524.400 85.050 525.600 ;
        RECT 61.950 523.950 64.050 524.400 ;
        RECT 76.950 523.950 79.050 524.400 ;
        RECT 82.950 523.950 85.050 524.400 ;
        RECT 94.950 525.600 97.050 526.050 ;
        RECT 100.950 525.600 103.050 526.050 ;
        RECT 94.950 524.400 103.050 525.600 ;
        RECT 94.950 523.950 97.050 524.400 ;
        RECT 100.950 523.950 103.050 524.400 ;
        RECT 109.950 525.600 112.050 526.050 ;
        RECT 115.950 525.600 118.050 526.050 ;
        RECT 130.950 525.600 133.050 526.050 ;
        RECT 109.950 524.400 133.050 525.600 ;
        RECT 109.950 523.950 112.050 524.400 ;
        RECT 115.950 523.950 118.050 524.400 ;
        RECT 130.950 523.950 133.050 524.400 ;
        RECT 139.950 523.950 142.050 526.050 ;
        RECT 145.950 523.950 148.050 526.050 ;
        RECT 160.950 525.600 163.050 526.050 ;
        RECT 169.950 525.600 172.050 526.050 ;
        RECT 160.950 524.400 172.050 525.600 ;
        RECT 160.950 523.950 163.050 524.400 ;
        RECT 169.950 523.950 172.050 524.400 ;
        RECT 241.950 523.950 244.050 526.050 ;
        RECT 286.950 525.600 289.050 526.050 ;
        RECT 301.950 525.600 304.050 526.050 ;
        RECT 286.950 524.400 304.050 525.600 ;
        RECT 286.950 523.950 289.050 524.400 ;
        RECT 301.950 523.950 304.050 524.400 ;
        RECT 379.950 525.600 382.050 526.050 ;
        RECT 385.950 525.600 388.050 526.050 ;
        RECT 379.950 524.400 388.050 525.600 ;
        RECT 379.950 523.950 382.050 524.400 ;
        RECT 385.950 523.950 388.050 524.400 ;
        RECT 388.950 525.600 391.050 526.050 ;
        RECT 398.400 525.600 399.600 526.950 ;
        RECT 388.950 524.400 399.600 525.600 ;
        RECT 424.950 525.600 427.050 526.050 ;
        RECT 433.950 525.600 436.050 526.050 ;
        RECT 424.950 524.400 436.050 525.600 ;
        RECT 388.950 523.950 391.050 524.400 ;
        RECT 424.950 523.950 427.050 524.400 ;
        RECT 433.950 523.950 436.050 524.400 ;
        RECT 493.950 525.600 496.050 526.050 ;
        RECT 511.950 525.600 514.050 526.050 ;
        RECT 493.950 524.400 514.050 525.600 ;
        RECT 493.950 523.950 496.050 524.400 ;
        RECT 511.950 523.950 514.050 524.400 ;
        RECT 520.950 525.600 523.050 526.050 ;
        RECT 526.950 525.600 529.050 526.050 ;
        RECT 520.950 524.400 529.050 525.600 ;
        RECT 520.950 523.950 523.050 524.400 ;
        RECT 526.950 523.950 529.050 524.400 ;
        RECT 19.950 522.600 22.050 523.050 ;
        RECT 34.950 522.600 37.050 523.050 ;
        RECT 19.950 521.400 37.050 522.600 ;
        RECT 19.950 520.950 22.050 521.400 ;
        RECT 34.950 520.950 37.050 521.400 ;
        RECT 46.950 522.600 49.050 523.050 ;
        RECT 64.950 522.600 67.050 523.050 ;
        RECT 46.950 521.400 67.050 522.600 ;
        RECT 46.950 520.950 49.050 521.400 ;
        RECT 64.950 520.950 67.050 521.400 ;
        RECT 73.950 522.600 76.050 523.050 ;
        RECT 85.950 522.600 88.050 523.050 ;
        RECT 73.950 521.400 88.050 522.600 ;
        RECT 73.950 520.950 76.050 521.400 ;
        RECT 85.950 520.950 88.050 521.400 ;
        RECT 91.950 520.950 94.050 523.050 ;
        RECT 97.950 522.600 100.050 523.050 ;
        RECT 106.950 522.600 109.050 523.050 ;
        RECT 127.950 522.600 130.050 523.050 ;
        RECT 97.950 521.400 130.050 522.600 ;
        RECT 97.950 520.950 100.050 521.400 ;
        RECT 106.950 520.950 109.050 521.400 ;
        RECT 127.950 520.950 130.050 521.400 ;
        RECT 184.950 522.600 187.050 523.050 ;
        RECT 196.950 522.600 199.050 523.050 ;
        RECT 184.950 521.400 199.050 522.600 ;
        RECT 184.950 520.950 187.050 521.400 ;
        RECT 196.950 520.950 199.050 521.400 ;
        RECT 211.950 522.600 214.050 523.050 ;
        RECT 223.950 522.600 226.050 523.050 ;
        RECT 211.950 521.400 226.050 522.600 ;
        RECT 242.400 522.600 243.600 523.950 ;
        RECT 554.400 523.050 555.600 526.950 ;
        RECT 556.950 525.600 559.050 526.050 ;
        RECT 562.950 525.600 565.050 526.050 ;
        RECT 556.950 524.400 565.050 525.600 ;
        RECT 556.950 523.950 559.050 524.400 ;
        RECT 562.950 523.950 565.050 524.400 ;
        RECT 565.950 525.600 568.050 526.050 ;
        RECT 574.950 525.600 577.050 526.050 ;
        RECT 599.400 525.600 600.600 526.950 ;
        RECT 565.950 524.400 600.600 525.600 ;
        RECT 628.950 525.600 631.050 526.050 ;
        RECT 643.950 525.600 646.050 526.050 ;
        RECT 628.950 524.400 646.050 525.600 ;
        RECT 565.950 523.950 568.050 524.400 ;
        RECT 574.950 523.950 577.050 524.400 ;
        RECT 628.950 523.950 631.050 524.400 ;
        RECT 643.950 523.950 646.050 524.400 ;
        RECT 649.950 525.600 652.050 526.050 ;
        RECT 676.950 525.600 679.050 526.050 ;
        RECT 649.950 524.400 679.050 525.600 ;
        RECT 649.950 523.950 652.050 524.400 ;
        RECT 676.950 523.950 679.050 524.400 ;
        RECT 697.950 525.600 700.050 526.050 ;
        RECT 796.950 525.600 799.050 526.050 ;
        RECT 802.950 525.600 805.050 526.050 ;
        RECT 697.950 524.400 805.050 525.600 ;
        RECT 697.950 523.950 700.050 524.400 ;
        RECT 796.950 523.950 799.050 524.400 ;
        RECT 802.950 523.950 805.050 524.400 ;
        RECT 319.950 522.600 322.050 523.050 ;
        RECT 328.950 522.600 331.050 523.050 ;
        RECT 242.400 521.400 331.050 522.600 ;
        RECT 211.950 520.950 214.050 521.400 ;
        RECT 223.950 520.950 226.050 521.400 ;
        RECT 319.950 520.950 322.050 521.400 ;
        RECT 328.950 520.950 331.050 521.400 ;
        RECT 355.950 522.600 358.050 523.050 ;
        RECT 373.950 522.600 376.050 523.050 ;
        RECT 355.950 521.400 376.050 522.600 ;
        RECT 355.950 520.950 358.050 521.400 ;
        RECT 373.950 520.950 376.050 521.400 ;
        RECT 391.950 522.600 394.050 523.050 ;
        RECT 412.950 522.600 415.050 523.050 ;
        RECT 544.950 522.600 547.050 523.050 ;
        RECT 391.950 521.400 415.050 522.600 ;
        RECT 391.950 520.950 394.050 521.400 ;
        RECT 412.950 520.950 415.050 521.400 ;
        RECT 449.400 521.400 547.050 522.600 ;
        RECT 40.950 519.600 43.050 520.050 ;
        RECT 70.950 519.600 73.050 520.050 ;
        RECT 40.950 518.400 73.050 519.600 ;
        RECT 40.950 517.950 43.050 518.400 ;
        RECT 70.950 517.950 73.050 518.400 ;
        RECT 79.950 519.600 82.050 520.050 ;
        RECT 92.400 519.600 93.600 520.950 ;
        RECT 79.950 518.400 93.600 519.600 ;
        RECT 253.950 519.600 256.050 520.050 ;
        RECT 283.950 519.600 286.050 520.050 ;
        RECT 253.950 518.400 286.050 519.600 ;
        RECT 79.950 517.950 82.050 518.400 ;
        RECT 253.950 517.950 256.050 518.400 ;
        RECT 283.950 517.950 286.050 518.400 ;
        RECT 301.950 519.600 304.050 520.050 ;
        RECT 316.950 519.600 319.050 520.050 ;
        RECT 301.950 518.400 319.050 519.600 ;
        RECT 301.950 517.950 304.050 518.400 ;
        RECT 316.950 517.950 319.050 518.400 ;
        RECT 322.950 519.600 325.050 520.050 ;
        RECT 391.950 519.600 394.050 520.050 ;
        RECT 322.950 518.400 394.050 519.600 ;
        RECT 322.950 517.950 325.050 518.400 ;
        RECT 391.950 517.950 394.050 518.400 ;
        RECT 412.950 519.600 415.050 520.050 ;
        RECT 449.400 519.600 450.600 521.400 ;
        RECT 544.950 520.950 547.050 521.400 ;
        RECT 553.950 520.950 556.050 523.050 ;
        RECT 652.950 522.600 655.050 523.050 ;
        RECT 664.950 522.600 667.050 523.050 ;
        RECT 673.950 522.600 676.050 523.050 ;
        RECT 652.950 521.400 676.050 522.600 ;
        RECT 652.950 520.950 655.050 521.400 ;
        RECT 664.950 520.950 667.050 521.400 ;
        RECT 673.950 520.950 676.050 521.400 ;
        RECT 754.950 522.600 757.050 523.050 ;
        RECT 760.950 522.600 763.050 523.050 ;
        RECT 754.950 521.400 763.050 522.600 ;
        RECT 754.950 520.950 757.050 521.400 ;
        RECT 760.950 520.950 763.050 521.400 ;
        RECT 781.950 522.600 784.050 523.050 ;
        RECT 787.950 522.600 790.050 523.050 ;
        RECT 781.950 521.400 790.050 522.600 ;
        RECT 781.950 520.950 784.050 521.400 ;
        RECT 787.950 520.950 790.050 521.400 ;
        RECT 412.950 518.400 450.600 519.600 ;
        RECT 451.950 519.600 454.050 520.050 ;
        RECT 496.950 519.600 499.050 520.050 ;
        RECT 451.950 518.400 499.050 519.600 ;
        RECT 412.950 517.950 415.050 518.400 ;
        RECT 451.950 517.950 454.050 518.400 ;
        RECT 496.950 517.950 499.050 518.400 ;
        RECT 544.950 519.600 547.050 520.050 ;
        RECT 550.950 519.600 553.050 520.050 ;
        RECT 544.950 518.400 553.050 519.600 ;
        RECT 544.950 517.950 547.050 518.400 ;
        RECT 550.950 517.950 553.050 518.400 ;
        RECT 580.950 519.600 583.050 520.050 ;
        RECT 592.950 519.600 595.050 520.050 ;
        RECT 580.950 518.400 595.050 519.600 ;
        RECT 580.950 517.950 583.050 518.400 ;
        RECT 592.950 517.950 595.050 518.400 ;
        RECT 13.950 516.600 16.050 517.050 ;
        RECT 22.950 516.600 25.050 517.050 ;
        RECT 13.950 515.400 25.050 516.600 ;
        RECT 13.950 514.950 16.050 515.400 ;
        RECT 22.950 514.950 25.050 515.400 ;
        RECT 49.950 516.600 52.050 517.050 ;
        RECT 112.950 516.600 115.050 517.050 ;
        RECT 49.950 515.400 115.050 516.600 ;
        RECT 49.950 514.950 52.050 515.400 ;
        RECT 112.950 514.950 115.050 515.400 ;
        RECT 295.950 516.600 298.050 517.050 ;
        RECT 304.950 516.600 307.050 517.050 ;
        RECT 295.950 515.400 307.050 516.600 ;
        RECT 295.950 514.950 298.050 515.400 ;
        RECT 304.950 514.950 307.050 515.400 ;
        RECT 367.950 516.600 370.050 517.050 ;
        RECT 622.950 516.600 625.050 517.050 ;
        RECT 640.950 516.600 643.050 517.050 ;
        RECT 367.950 515.400 643.050 516.600 ;
        RECT 367.950 514.950 370.050 515.400 ;
        RECT 622.950 514.950 625.050 515.400 ;
        RECT 640.950 514.950 643.050 515.400 ;
        RECT 787.950 516.600 790.050 517.050 ;
        RECT 793.950 516.600 796.050 517.050 ;
        RECT 787.950 515.400 796.050 516.600 ;
        RECT 842.400 516.600 843.600 530.400 ;
        RECT 847.950 529.950 850.050 530.400 ;
        RECT 853.950 528.600 856.050 529.050 ;
        RECT 845.400 527.400 856.050 528.600 ;
        RECT 845.400 519.600 846.600 527.400 ;
        RECT 853.950 526.950 856.050 527.400 ;
        RECT 847.950 519.600 850.050 520.050 ;
        RECT 845.400 518.400 850.050 519.600 ;
        RECT 847.950 517.950 850.050 518.400 ;
        RECT 842.400 515.400 861.600 516.600 ;
        RECT 787.950 514.950 790.050 515.400 ;
        RECT 793.950 514.950 796.050 515.400 ;
        RECT 7.950 513.600 10.050 514.050 ;
        RECT 13.950 513.600 16.050 514.050 ;
        RECT 7.950 512.400 16.050 513.600 ;
        RECT 7.950 511.950 10.050 512.400 ;
        RECT 13.950 511.950 16.050 512.400 ;
        RECT 154.950 513.600 157.050 514.050 ;
        RECT 331.950 513.600 334.050 514.050 ;
        RECT 154.950 512.400 334.050 513.600 ;
        RECT 154.950 511.950 157.050 512.400 ;
        RECT 331.950 511.950 334.050 512.400 ;
        RECT 391.950 513.600 394.050 514.050 ;
        RECT 433.950 513.600 436.050 514.050 ;
        RECT 391.950 512.400 436.050 513.600 ;
        RECT 391.950 511.950 394.050 512.400 ;
        RECT 433.950 511.950 436.050 512.400 ;
        RECT 442.950 513.600 445.050 514.050 ;
        RECT 538.950 513.600 541.050 514.050 ;
        RECT 442.950 512.400 541.050 513.600 ;
        RECT 442.950 511.950 445.050 512.400 ;
        RECT 538.950 511.950 541.050 512.400 ;
        RECT 166.950 510.600 169.050 511.050 ;
        RECT 238.950 510.600 241.050 511.050 ;
        RECT 400.950 510.600 403.050 511.050 ;
        RECT 424.950 510.600 427.050 511.050 ;
        RECT 469.950 510.600 472.050 511.050 ;
        RECT 166.950 509.400 472.050 510.600 ;
        RECT 166.950 508.950 169.050 509.400 ;
        RECT 238.950 508.950 241.050 509.400 ;
        RECT 400.950 508.950 403.050 509.400 ;
        RECT 424.950 508.950 427.050 509.400 ;
        RECT 469.950 508.950 472.050 509.400 ;
        RECT 571.950 510.600 574.050 511.050 ;
        RECT 586.950 510.600 589.050 511.050 ;
        RECT 595.950 510.600 598.050 511.050 ;
        RECT 571.950 509.400 598.050 510.600 ;
        RECT 571.950 508.950 574.050 509.400 ;
        RECT 586.950 508.950 589.050 509.400 ;
        RECT 595.950 508.950 598.050 509.400 ;
        RECT 730.950 510.600 733.050 511.050 ;
        RECT 769.950 510.600 772.050 511.050 ;
        RECT 790.950 510.600 793.050 511.050 ;
        RECT 730.950 509.400 793.050 510.600 ;
        RECT 730.950 508.950 733.050 509.400 ;
        RECT 769.950 508.950 772.050 509.400 ;
        RECT 790.950 508.950 793.050 509.400 ;
        RECT 841.950 510.600 844.050 511.050 ;
        RECT 847.950 510.600 850.050 511.050 ;
        RECT 841.950 509.400 850.050 510.600 ;
        RECT 841.950 508.950 844.050 509.400 ;
        RECT 847.950 508.950 850.050 509.400 ;
        RECT 178.950 507.600 181.050 508.050 ;
        RECT 520.950 507.600 523.050 508.050 ;
        RECT 178.950 506.400 523.050 507.600 ;
        RECT 178.950 505.950 181.050 506.400 ;
        RECT 520.950 505.950 523.050 506.400 ;
        RECT 736.950 507.600 739.050 508.050 ;
        RECT 751.950 507.600 754.050 508.050 ;
        RECT 736.950 506.400 754.050 507.600 ;
        RECT 736.950 505.950 739.050 506.400 ;
        RECT 751.950 505.950 754.050 506.400 ;
        RECT 860.400 505.050 861.600 515.400 ;
        RECT 16.950 504.600 19.050 505.050 ;
        RECT 25.950 504.600 28.050 505.050 ;
        RECT 79.950 504.600 82.050 505.050 ;
        RECT 16.950 503.400 82.050 504.600 ;
        RECT 16.950 502.950 19.050 503.400 ;
        RECT 25.950 502.950 28.050 503.400 ;
        RECT 79.950 502.950 82.050 503.400 ;
        RECT 151.950 504.600 154.050 505.050 ;
        RECT 172.950 504.600 175.050 505.050 ;
        RECT 151.950 503.400 175.050 504.600 ;
        RECT 151.950 502.950 154.050 503.400 ;
        RECT 172.950 502.950 175.050 503.400 ;
        RECT 175.950 504.600 178.050 505.050 ;
        RECT 190.950 504.600 193.050 505.050 ;
        RECT 175.950 503.400 193.050 504.600 ;
        RECT 175.950 502.950 178.050 503.400 ;
        RECT 190.950 502.950 193.050 503.400 ;
        RECT 244.950 504.600 247.050 505.050 ;
        RECT 250.950 504.600 253.050 505.050 ;
        RECT 343.950 504.600 346.050 505.050 ;
        RECT 406.950 504.600 409.050 505.050 ;
        RECT 244.950 503.400 409.050 504.600 ;
        RECT 244.950 502.950 247.050 503.400 ;
        RECT 250.950 502.950 253.050 503.400 ;
        RECT 343.950 502.950 346.050 503.400 ;
        RECT 406.950 502.950 409.050 503.400 ;
        RECT 415.950 504.600 418.050 505.050 ;
        RECT 430.950 504.600 433.050 505.050 ;
        RECT 415.950 503.400 433.050 504.600 ;
        RECT 415.950 502.950 418.050 503.400 ;
        RECT 430.950 502.950 433.050 503.400 ;
        RECT 688.950 504.600 691.050 505.050 ;
        RECT 706.950 504.600 709.050 505.050 ;
        RECT 688.950 503.400 709.050 504.600 ;
        RECT 688.950 502.950 691.050 503.400 ;
        RECT 706.950 502.950 709.050 503.400 ;
        RECT 769.950 504.600 772.050 505.050 ;
        RECT 775.950 504.600 778.050 505.050 ;
        RECT 769.950 503.400 778.050 504.600 ;
        RECT 769.950 502.950 772.050 503.400 ;
        RECT 775.950 502.950 778.050 503.400 ;
        RECT 859.950 502.950 862.050 505.050 ;
        RECT 46.950 501.600 49.050 502.050 ;
        RECT 64.950 501.600 67.050 502.050 ;
        RECT 46.950 500.400 67.050 501.600 ;
        RECT 46.950 499.950 49.050 500.400 ;
        RECT 64.950 499.950 67.050 500.400 ;
        RECT 211.950 501.600 214.050 502.050 ;
        RECT 304.950 501.600 307.050 502.050 ;
        RECT 394.950 501.600 397.050 502.050 ;
        RECT 211.950 500.400 397.050 501.600 ;
        RECT 211.950 499.950 214.050 500.400 ;
        RECT 304.950 499.950 307.050 500.400 ;
        RECT 394.950 499.950 397.050 500.400 ;
        RECT 430.950 501.600 433.050 502.050 ;
        RECT 478.950 501.600 481.050 502.050 ;
        RECT 496.950 501.600 499.050 502.050 ;
        RECT 430.950 500.400 499.050 501.600 ;
        RECT 430.950 499.950 433.050 500.400 ;
        RECT 478.950 499.950 481.050 500.400 ;
        RECT 496.950 499.950 499.050 500.400 ;
        RECT 823.950 501.600 826.050 502.050 ;
        RECT 832.950 501.600 835.050 502.050 ;
        RECT 823.950 500.400 835.050 501.600 ;
        RECT 823.950 499.950 826.050 500.400 ;
        RECT 832.950 499.950 835.050 500.400 ;
        RECT 115.950 498.600 118.050 499.050 ;
        RECT 121.950 498.600 124.050 499.050 ;
        RECT 115.950 497.400 124.050 498.600 ;
        RECT 115.950 496.950 118.050 497.400 ;
        RECT 121.950 496.950 124.050 497.400 ;
        RECT 181.950 498.600 184.050 499.050 ;
        RECT 262.950 498.600 265.050 499.050 ;
        RECT 427.950 498.600 430.050 499.050 ;
        RECT 181.950 497.400 430.050 498.600 ;
        RECT 181.950 496.950 184.050 497.400 ;
        RECT 262.950 496.950 265.050 497.400 ;
        RECT 427.950 496.950 430.050 497.400 ;
        RECT 118.950 495.600 121.050 496.050 ;
        RECT 124.950 495.600 127.050 496.050 ;
        RECT 127.950 495.600 130.050 496.050 ;
        RECT 118.950 494.400 130.050 495.600 ;
        RECT 118.950 493.950 121.050 494.400 ;
        RECT 124.950 493.950 127.050 494.400 ;
        RECT 127.950 493.950 130.050 494.400 ;
        RECT 397.950 495.600 400.050 496.050 ;
        RECT 439.950 495.600 442.050 496.050 ;
        RECT 523.950 495.600 526.050 496.050 ;
        RECT 397.950 494.400 442.050 495.600 ;
        RECT 397.950 493.950 400.050 494.400 ;
        RECT 439.950 493.950 442.050 494.400 ;
        RECT 458.400 494.400 526.050 495.600 ;
        RECT 82.950 492.600 85.050 493.050 ;
        RECT 118.950 492.600 121.050 493.050 ;
        RECT 82.950 491.400 121.050 492.600 ;
        RECT 82.950 490.950 85.050 491.400 ;
        RECT 118.950 490.950 121.050 491.400 ;
        RECT 289.950 492.600 292.050 493.050 ;
        RECT 391.950 492.600 394.050 493.050 ;
        RECT 289.950 491.400 394.050 492.600 ;
        RECT 289.950 490.950 292.050 491.400 ;
        RECT 391.950 490.950 394.050 491.400 ;
        RECT 406.950 492.600 409.050 493.050 ;
        RECT 418.950 492.600 421.050 493.050 ;
        RECT 448.950 492.600 451.050 493.050 ;
        RECT 458.400 492.600 459.600 494.400 ;
        RECT 523.950 493.950 526.050 494.400 ;
        RECT 745.950 495.600 748.050 496.050 ;
        RECT 844.950 495.600 847.050 496.050 ;
        RECT 853.950 495.600 856.050 496.050 ;
        RECT 745.950 494.400 856.050 495.600 ;
        RECT 745.950 493.950 748.050 494.400 ;
        RECT 844.950 493.950 847.050 494.400 ;
        RECT 853.950 493.950 856.050 494.400 ;
        RECT 406.950 491.400 459.600 492.600 ;
        RECT 460.950 492.600 463.050 493.050 ;
        RECT 475.950 492.600 478.050 493.050 ;
        RECT 460.950 491.400 478.050 492.600 ;
        RECT 406.950 490.950 409.050 491.400 ;
        RECT 418.950 490.950 421.050 491.400 ;
        RECT 448.950 490.950 451.050 491.400 ;
        RECT 460.950 490.950 463.050 491.400 ;
        RECT 475.950 490.950 478.050 491.400 ;
        RECT 535.950 492.600 538.050 493.050 ;
        RECT 541.950 492.600 544.050 493.050 ;
        RECT 553.950 492.600 556.050 493.050 ;
        RECT 535.950 491.400 544.050 492.600 ;
        RECT 535.950 490.950 538.050 491.400 ;
        RECT 541.950 490.950 544.050 491.400 ;
        RECT 551.400 491.400 556.050 492.600 ;
        RECT 551.400 490.050 552.600 491.400 ;
        RECT 553.950 490.950 556.050 491.400 ;
        RECT 691.950 492.600 694.050 493.050 ;
        RECT 781.950 492.600 784.050 493.050 ;
        RECT 691.950 491.400 784.050 492.600 ;
        RECT 691.950 490.950 694.050 491.400 ;
        RECT 781.950 490.950 784.050 491.400 ;
        RECT 841.950 492.600 844.050 493.050 ;
        RECT 853.950 492.600 856.050 493.050 ;
        RECT 841.950 491.400 856.050 492.600 ;
        RECT 841.950 490.950 844.050 491.400 ;
        RECT 853.950 490.950 856.050 491.400 ;
        RECT 7.950 489.600 10.050 490.050 ;
        RECT 55.950 489.600 58.050 490.050 ;
        RECT 7.950 488.400 58.050 489.600 ;
        RECT 7.950 487.950 10.050 488.400 ;
        RECT 55.950 487.950 58.050 488.400 ;
        RECT 97.950 489.600 100.050 490.050 ;
        RECT 133.950 489.600 136.050 490.050 ;
        RECT 97.950 488.400 136.050 489.600 ;
        RECT 97.950 487.950 100.050 488.400 ;
        RECT 133.950 487.950 136.050 488.400 ;
        RECT 229.950 489.600 232.050 490.050 ;
        RECT 238.950 489.600 241.050 490.050 ;
        RECT 229.950 488.400 241.050 489.600 ;
        RECT 229.950 487.950 232.050 488.400 ;
        RECT 238.950 487.950 241.050 488.400 ;
        RECT 259.950 489.600 262.050 490.050 ;
        RECT 319.950 489.600 322.050 490.050 ;
        RECT 259.950 488.400 322.050 489.600 ;
        RECT 259.950 487.950 262.050 488.400 ;
        RECT 319.950 487.950 322.050 488.400 ;
        RECT 358.950 489.600 361.050 490.050 ;
        RECT 382.950 489.600 385.050 490.050 ;
        RECT 358.950 488.400 385.050 489.600 ;
        RECT 358.950 487.950 361.050 488.400 ;
        RECT 382.950 487.950 385.050 488.400 ;
        RECT 427.950 487.950 430.050 490.050 ;
        RECT 457.950 489.600 460.050 490.050 ;
        RECT 541.950 489.600 544.050 490.050 ;
        RECT 457.950 488.400 544.050 489.600 ;
        RECT 457.950 487.950 460.050 488.400 ;
        RECT 541.950 487.950 544.050 488.400 ;
        RECT 550.950 487.950 553.050 490.050 ;
        RECT 628.950 489.600 631.050 490.050 ;
        RECT 634.950 489.600 637.050 490.050 ;
        RECT 628.950 488.400 637.050 489.600 ;
        RECT 628.950 487.950 631.050 488.400 ;
        RECT 634.950 487.950 637.050 488.400 ;
        RECT 739.950 489.600 742.050 490.050 ;
        RECT 739.950 488.400 771.600 489.600 ;
        RECT 739.950 487.950 742.050 488.400 ;
        RECT 43.950 486.600 46.050 487.050 ;
        RECT 49.950 486.600 52.050 487.050 ;
        RECT 43.950 485.400 52.050 486.600 ;
        RECT 43.950 484.950 46.050 485.400 ;
        RECT 49.950 484.950 52.050 485.400 ;
        RECT 70.950 486.600 73.050 487.050 ;
        RECT 94.950 486.600 97.050 487.050 ;
        RECT 70.950 485.400 97.050 486.600 ;
        RECT 70.950 484.950 73.050 485.400 ;
        RECT 94.950 484.950 97.050 485.400 ;
        RECT 100.950 486.600 103.050 487.050 ;
        RECT 109.950 486.600 112.050 487.050 ;
        RECT 100.950 485.400 112.050 486.600 ;
        RECT 100.950 484.950 103.050 485.400 ;
        RECT 109.950 484.950 112.050 485.400 ;
        RECT 187.950 486.600 190.050 487.050 ;
        RECT 256.950 486.600 259.050 487.050 ;
        RECT 289.950 486.600 292.050 487.050 ;
        RECT 187.950 485.400 259.050 486.600 ;
        RECT 187.950 484.950 190.050 485.400 ;
        RECT 256.950 484.950 259.050 485.400 ;
        RECT 275.400 485.400 292.050 486.600 ;
        RECT 275.400 484.050 276.600 485.400 ;
        RECT 289.950 484.950 292.050 485.400 ;
        RECT 325.950 486.600 328.050 487.050 ;
        RECT 337.950 486.600 340.050 487.050 ;
        RECT 349.950 486.600 352.050 487.050 ;
        RECT 325.950 485.400 352.050 486.600 ;
        RECT 325.950 484.950 328.050 485.400 ;
        RECT 337.950 484.950 340.050 485.400 ;
        RECT 349.950 484.950 352.050 485.400 ;
        RECT 355.950 486.600 358.050 487.050 ;
        RECT 361.950 486.600 364.050 487.050 ;
        RECT 370.950 486.600 373.050 487.050 ;
        RECT 355.950 485.400 373.050 486.600 ;
        RECT 355.950 484.950 358.050 485.400 ;
        RECT 361.950 484.950 364.050 485.400 ;
        RECT 370.950 484.950 373.050 485.400 ;
        RECT 382.950 486.600 385.050 487.050 ;
        RECT 394.950 486.600 397.050 487.050 ;
        RECT 400.950 486.600 403.050 487.050 ;
        RECT 418.950 486.600 421.050 487.050 ;
        RECT 382.950 485.400 403.050 486.600 ;
        RECT 382.950 484.950 385.050 485.400 ;
        RECT 394.950 484.950 397.050 485.400 ;
        RECT 400.950 484.950 403.050 485.400 ;
        RECT 407.400 485.400 421.050 486.600 ;
        RECT 19.950 483.600 22.050 484.050 ;
        RECT 22.950 483.600 25.050 484.050 ;
        RECT 40.950 483.600 43.050 484.050 ;
        RECT 19.950 482.400 43.050 483.600 ;
        RECT 19.950 481.950 22.050 482.400 ;
        RECT 22.950 481.950 25.050 482.400 ;
        RECT 40.950 481.950 43.050 482.400 ;
        RECT 58.950 483.600 61.050 484.050 ;
        RECT 64.950 483.600 67.050 484.050 ;
        RECT 91.950 483.600 94.050 484.050 ;
        RECT 58.950 482.400 94.050 483.600 ;
        RECT 58.950 481.950 61.050 482.400 ;
        RECT 64.950 481.950 67.050 482.400 ;
        RECT 91.950 481.950 94.050 482.400 ;
        RECT 112.950 483.600 115.050 484.050 ;
        RECT 121.950 483.600 124.050 484.050 ;
        RECT 112.950 482.400 124.050 483.600 ;
        RECT 112.950 481.950 115.050 482.400 ;
        RECT 121.950 481.950 124.050 482.400 ;
        RECT 193.950 483.600 196.050 484.050 ;
        RECT 202.950 483.600 205.050 484.050 ;
        RECT 193.950 482.400 205.050 483.600 ;
        RECT 193.950 481.950 196.050 482.400 ;
        RECT 202.950 481.950 205.050 482.400 ;
        RECT 208.950 483.600 211.050 484.050 ;
        RECT 220.950 483.600 223.050 484.050 ;
        RECT 208.950 482.400 223.050 483.600 ;
        RECT 208.950 481.950 211.050 482.400 ;
        RECT 220.950 481.950 223.050 482.400 ;
        RECT 247.950 483.600 250.050 484.050 ;
        RECT 262.950 483.600 265.050 484.050 ;
        RECT 268.950 483.600 271.050 484.050 ;
        RECT 247.950 482.400 265.050 483.600 ;
        RECT 247.950 481.950 250.050 482.400 ;
        RECT 262.950 481.950 265.050 482.400 ;
        RECT 266.400 482.400 271.050 483.600 ;
        RECT 46.950 480.600 49.050 481.050 ;
        RECT 61.950 480.600 64.050 481.050 ;
        RECT 70.950 480.600 73.050 481.050 ;
        RECT 46.950 479.400 73.050 480.600 ;
        RECT 46.950 478.950 49.050 479.400 ;
        RECT 61.950 478.950 64.050 479.400 ;
        RECT 70.950 478.950 73.050 479.400 ;
        RECT 73.950 480.600 76.050 481.050 ;
        RECT 100.950 480.600 103.050 481.050 ;
        RECT 73.950 479.400 103.050 480.600 ;
        RECT 73.950 478.950 76.050 479.400 ;
        RECT 100.950 478.950 103.050 479.400 ;
        RECT 175.950 480.600 178.050 481.050 ;
        RECT 193.950 480.600 196.050 481.050 ;
        RECT 175.950 479.400 196.050 480.600 ;
        RECT 175.950 478.950 178.050 479.400 ;
        RECT 193.950 478.950 196.050 479.400 ;
        RECT 217.950 480.600 220.050 481.050 ;
        RECT 223.950 480.600 226.050 481.050 ;
        RECT 217.950 479.400 226.050 480.600 ;
        RECT 217.950 478.950 220.050 479.400 ;
        RECT 223.950 478.950 226.050 479.400 ;
        RECT 232.950 480.600 235.050 481.050 ;
        RECT 253.950 480.600 256.050 481.050 ;
        RECT 232.950 479.400 256.050 480.600 ;
        RECT 232.950 478.950 235.050 479.400 ;
        RECT 253.950 478.950 256.050 479.400 ;
        RECT 262.950 480.600 265.050 481.050 ;
        RECT 266.400 480.600 267.600 482.400 ;
        RECT 268.950 481.950 271.050 482.400 ;
        RECT 274.950 481.950 277.050 484.050 ;
        RECT 316.950 483.600 319.050 484.050 ;
        RECT 290.400 482.400 319.050 483.600 ;
        RECT 290.400 481.050 291.600 482.400 ;
        RECT 316.950 481.950 319.050 482.400 ;
        RECT 322.950 483.600 325.050 484.050 ;
        RECT 385.950 483.600 388.050 484.050 ;
        RECT 397.950 483.600 400.050 484.050 ;
        RECT 322.950 482.400 400.050 483.600 ;
        RECT 322.950 481.950 325.050 482.400 ;
        RECT 385.950 481.950 388.050 482.400 ;
        RECT 397.950 481.950 400.050 482.400 ;
        RECT 403.950 483.600 406.050 484.050 ;
        RECT 407.400 483.600 408.600 485.400 ;
        RECT 418.950 484.950 421.050 485.400 ;
        RECT 403.950 482.400 408.600 483.600 ;
        RECT 409.950 483.600 412.050 484.050 ;
        RECT 428.400 483.600 429.600 487.950 ;
        RECT 770.400 487.050 771.600 488.400 ;
        RECT 469.950 486.600 472.050 487.050 ;
        RECT 475.950 486.600 478.050 487.050 ;
        RECT 469.950 485.400 478.050 486.600 ;
        RECT 469.950 484.950 472.050 485.400 ;
        RECT 475.950 484.950 478.050 485.400 ;
        RECT 502.950 484.950 505.050 487.050 ;
        RECT 535.950 486.600 538.050 487.050 ;
        RECT 547.950 486.600 550.050 487.050 ;
        RECT 643.950 486.600 646.050 487.050 ;
        RECT 535.950 485.400 550.050 486.600 ;
        RECT 535.950 484.950 538.050 485.400 ;
        RECT 547.950 484.950 550.050 485.400 ;
        RECT 620.400 485.400 646.050 486.600 ;
        RECT 445.950 483.600 448.050 484.050 ;
        RECT 409.950 482.400 448.050 483.600 ;
        RECT 403.950 481.950 406.050 482.400 ;
        RECT 409.950 481.950 412.050 482.400 ;
        RECT 445.950 481.950 448.050 482.400 ;
        RECT 451.950 483.600 454.050 484.050 ;
        RECT 463.950 483.600 466.050 484.050 ;
        RECT 451.950 482.400 466.050 483.600 ;
        RECT 451.950 481.950 454.050 482.400 ;
        RECT 463.950 481.950 466.050 482.400 ;
        RECT 484.950 483.600 487.050 484.050 ;
        RECT 503.400 483.600 504.600 484.950 ;
        RECT 620.400 484.050 621.600 485.400 ;
        RECT 643.950 484.950 646.050 485.400 ;
        RECT 664.950 486.600 667.050 487.050 ;
        RECT 694.950 486.600 697.050 487.050 ;
        RECT 664.950 485.400 697.050 486.600 ;
        RECT 664.950 484.950 667.050 485.400 ;
        RECT 694.950 484.950 697.050 485.400 ;
        RECT 724.950 486.600 727.050 487.050 ;
        RECT 730.950 486.600 733.050 487.050 ;
        RECT 724.950 485.400 733.050 486.600 ;
        RECT 724.950 484.950 727.050 485.400 ;
        RECT 730.950 484.950 733.050 485.400 ;
        RECT 769.950 484.950 772.050 487.050 ;
        RECT 484.950 482.400 504.600 483.600 ;
        RECT 529.950 483.600 532.050 484.050 ;
        RECT 538.950 483.600 541.050 484.050 ;
        RECT 574.950 483.600 577.050 484.050 ;
        RECT 529.950 482.400 577.050 483.600 ;
        RECT 484.950 481.950 487.050 482.400 ;
        RECT 529.950 481.950 532.050 482.400 ;
        RECT 538.950 481.950 541.050 482.400 ;
        RECT 574.950 481.950 577.050 482.400 ;
        RECT 619.950 481.950 622.050 484.050 ;
        RECT 718.950 483.600 721.050 484.050 ;
        RECT 739.950 483.600 742.050 484.050 ;
        RECT 745.950 483.600 748.050 484.050 ;
        RECT 718.950 482.400 748.050 483.600 ;
        RECT 718.950 481.950 721.050 482.400 ;
        RECT 739.950 481.950 742.050 482.400 ;
        RECT 745.950 481.950 748.050 482.400 ;
        RECT 262.950 479.400 267.600 480.600 ;
        RECT 271.950 480.600 274.050 481.050 ;
        RECT 280.950 480.600 283.050 481.050 ;
        RECT 271.950 479.400 283.050 480.600 ;
        RECT 262.950 478.950 265.050 479.400 ;
        RECT 271.950 478.950 274.050 479.400 ;
        RECT 280.950 478.950 283.050 479.400 ;
        RECT 289.950 478.950 292.050 481.050 ;
        RECT 292.950 480.600 295.050 481.050 ;
        RECT 316.950 480.600 319.050 481.050 ;
        RECT 292.950 479.400 319.050 480.600 ;
        RECT 292.950 478.950 295.050 479.400 ;
        RECT 316.950 478.950 319.050 479.400 ;
        RECT 340.950 480.600 343.050 481.050 ;
        RECT 346.950 480.600 349.050 481.050 ;
        RECT 340.950 479.400 349.050 480.600 ;
        RECT 340.950 478.950 343.050 479.400 ;
        RECT 346.950 478.950 349.050 479.400 ;
        RECT 367.950 480.600 370.050 481.050 ;
        RECT 391.950 480.600 394.050 481.050 ;
        RECT 367.950 479.400 394.050 480.600 ;
        RECT 367.950 478.950 370.050 479.400 ;
        RECT 391.950 478.950 394.050 479.400 ;
        RECT 418.950 480.600 421.050 481.050 ;
        RECT 430.950 480.600 433.050 481.050 ;
        RECT 418.950 479.400 433.050 480.600 ;
        RECT 418.950 478.950 421.050 479.400 ;
        RECT 430.950 478.950 433.050 479.400 ;
        RECT 472.950 480.600 475.050 481.050 ;
        RECT 478.950 480.600 481.050 481.050 ;
        RECT 472.950 479.400 481.050 480.600 ;
        RECT 472.950 478.950 475.050 479.400 ;
        RECT 478.950 478.950 481.050 479.400 ;
        RECT 661.950 480.600 664.050 481.050 ;
        RECT 691.950 480.600 694.050 481.050 ;
        RECT 661.950 479.400 694.050 480.600 ;
        RECT 661.950 478.950 664.050 479.400 ;
        RECT 691.950 478.950 694.050 479.400 ;
        RECT 727.950 480.600 730.050 481.050 ;
        RECT 748.950 480.600 751.050 481.050 ;
        RECT 763.950 480.600 766.050 481.050 ;
        RECT 727.950 479.400 766.050 480.600 ;
        RECT 727.950 478.950 730.050 479.400 ;
        RECT 748.950 478.950 751.050 479.400 ;
        RECT 763.950 478.950 766.050 479.400 ;
        RECT 25.950 477.600 28.050 478.050 ;
        RECT 49.950 477.600 52.050 478.050 ;
        RECT 52.950 477.600 55.050 478.050 ;
        RECT 25.950 476.400 55.050 477.600 ;
        RECT 25.950 475.950 28.050 476.400 ;
        RECT 49.950 475.950 52.050 476.400 ;
        RECT 52.950 475.950 55.050 476.400 ;
        RECT 148.950 477.600 151.050 478.050 ;
        RECT 235.950 477.600 238.050 478.050 ;
        RECT 148.950 476.400 238.050 477.600 ;
        RECT 148.950 475.950 151.050 476.400 ;
        RECT 235.950 475.950 238.050 476.400 ;
        RECT 241.950 477.600 244.050 478.050 ;
        RECT 259.950 477.600 262.050 478.050 ;
        RECT 241.950 476.400 262.050 477.600 ;
        RECT 241.950 475.950 244.050 476.400 ;
        RECT 259.950 475.950 262.050 476.400 ;
        RECT 307.950 477.600 310.050 478.050 ;
        RECT 319.950 477.600 322.050 478.050 ;
        RECT 334.950 477.600 337.050 478.050 ;
        RECT 307.950 476.400 337.050 477.600 ;
        RECT 307.950 475.950 310.050 476.400 ;
        RECT 319.950 475.950 322.050 476.400 ;
        RECT 334.950 475.950 337.050 476.400 ;
        RECT 379.950 477.600 382.050 478.050 ;
        RECT 472.950 477.600 475.050 478.050 ;
        RECT 379.950 476.400 475.050 477.600 ;
        RECT 379.950 475.950 382.050 476.400 ;
        RECT 472.950 475.950 475.050 476.400 ;
        RECT 565.950 477.600 568.050 478.050 ;
        RECT 727.950 477.600 730.050 478.050 ;
        RECT 565.950 476.400 730.050 477.600 ;
        RECT 565.950 475.950 568.050 476.400 ;
        RECT 727.950 475.950 730.050 476.400 ;
        RECT 64.950 474.600 67.050 475.050 ;
        RECT 133.950 474.600 136.050 475.050 ;
        RECT 196.950 474.600 199.050 475.050 ;
        RECT 211.950 474.600 214.050 475.050 ;
        RECT 64.950 473.400 214.050 474.600 ;
        RECT 64.950 472.950 67.050 473.400 ;
        RECT 133.950 472.950 136.050 473.400 ;
        RECT 196.950 472.950 199.050 473.400 ;
        RECT 211.950 472.950 214.050 473.400 ;
        RECT 229.950 474.600 232.050 475.050 ;
        RECT 235.950 474.600 238.050 475.050 ;
        RECT 274.950 474.600 277.050 475.050 ;
        RECT 229.950 473.400 238.050 474.600 ;
        RECT 229.950 472.950 232.050 473.400 ;
        RECT 235.950 472.950 238.050 473.400 ;
        RECT 239.400 473.400 277.050 474.600 ;
        RECT 88.950 471.600 91.050 472.050 ;
        RECT 94.950 471.600 97.050 472.050 ;
        RECT 106.950 471.600 109.050 472.050 ;
        RECT 88.950 470.400 109.050 471.600 ;
        RECT 88.950 469.950 91.050 470.400 ;
        RECT 94.950 469.950 97.050 470.400 ;
        RECT 106.950 469.950 109.050 470.400 ;
        RECT 220.950 471.600 223.050 472.050 ;
        RECT 239.400 471.600 240.600 473.400 ;
        RECT 274.950 472.950 277.050 473.400 ;
        RECT 286.950 474.600 289.050 475.050 ;
        RECT 310.950 474.600 313.050 475.050 ;
        RECT 286.950 473.400 313.050 474.600 ;
        RECT 286.950 472.950 289.050 473.400 ;
        RECT 310.950 472.950 313.050 473.400 ;
        RECT 334.950 474.600 337.050 475.050 ;
        RECT 379.950 474.600 382.050 475.050 ;
        RECT 334.950 473.400 382.050 474.600 ;
        RECT 334.950 472.950 337.050 473.400 ;
        RECT 379.950 472.950 382.050 473.400 ;
        RECT 385.950 474.600 388.050 475.050 ;
        RECT 409.950 474.600 412.050 475.050 ;
        RECT 385.950 473.400 412.050 474.600 ;
        RECT 385.950 472.950 388.050 473.400 ;
        RECT 409.950 472.950 412.050 473.400 ;
        RECT 427.950 474.600 430.050 475.050 ;
        RECT 436.950 474.600 439.050 475.050 ;
        RECT 427.950 473.400 439.050 474.600 ;
        RECT 427.950 472.950 430.050 473.400 ;
        RECT 436.950 472.950 439.050 473.400 ;
        RECT 445.950 474.600 448.050 475.050 ;
        RECT 466.950 474.600 469.050 475.050 ;
        RECT 502.950 474.600 505.050 475.050 ;
        RECT 445.950 473.400 465.600 474.600 ;
        RECT 445.950 472.950 448.050 473.400 ;
        RECT 220.950 470.400 240.600 471.600 ;
        RECT 262.950 471.600 265.050 472.050 ;
        RECT 292.950 471.600 295.050 472.050 ;
        RECT 262.950 470.400 295.050 471.600 ;
        RECT 220.950 469.950 223.050 470.400 ;
        RECT 262.950 469.950 265.050 470.400 ;
        RECT 292.950 469.950 295.050 470.400 ;
        RECT 295.950 471.600 298.050 472.050 ;
        RECT 304.950 471.600 307.050 472.050 ;
        RECT 295.950 470.400 307.050 471.600 ;
        RECT 295.950 469.950 298.050 470.400 ;
        RECT 304.950 469.950 307.050 470.400 ;
        RECT 316.950 471.600 319.050 472.050 ;
        RECT 361.950 471.600 364.050 472.050 ;
        RECT 400.950 471.600 403.050 472.050 ;
        RECT 406.950 471.600 409.050 472.050 ;
        RECT 316.950 470.400 360.600 471.600 ;
        RECT 316.950 469.950 319.050 470.400 ;
        RECT 232.950 468.600 235.050 469.050 ;
        RECT 355.950 468.600 358.050 469.050 ;
        RECT 232.950 467.400 358.050 468.600 ;
        RECT 359.400 468.600 360.600 470.400 ;
        RECT 361.950 470.400 409.050 471.600 ;
        RECT 361.950 469.950 364.050 470.400 ;
        RECT 400.950 469.950 403.050 470.400 ;
        RECT 406.950 469.950 409.050 470.400 ;
        RECT 412.950 471.600 415.050 472.050 ;
        RECT 427.950 471.600 430.050 472.050 ;
        RECT 412.950 470.400 430.050 471.600 ;
        RECT 464.400 471.600 465.600 473.400 ;
        RECT 466.950 473.400 505.050 474.600 ;
        RECT 466.950 472.950 469.050 473.400 ;
        RECT 502.950 472.950 505.050 473.400 ;
        RECT 616.950 474.600 619.050 475.050 ;
        RECT 634.950 474.600 637.050 475.050 ;
        RECT 616.950 473.400 637.050 474.600 ;
        RECT 616.950 472.950 619.050 473.400 ;
        RECT 634.950 472.950 637.050 473.400 ;
        RECT 481.950 471.600 484.050 472.050 ;
        RECT 464.400 470.400 484.050 471.600 ;
        RECT 412.950 469.950 415.050 470.400 ;
        RECT 427.950 469.950 430.050 470.400 ;
        RECT 481.950 469.950 484.050 470.400 ;
        RECT 487.950 471.600 490.050 472.050 ;
        RECT 502.950 471.600 505.050 472.050 ;
        RECT 487.950 470.400 505.050 471.600 ;
        RECT 487.950 469.950 490.050 470.400 ;
        RECT 502.950 469.950 505.050 470.400 ;
        RECT 697.950 471.600 700.050 472.050 ;
        RECT 718.950 471.600 721.050 472.050 ;
        RECT 697.950 470.400 721.050 471.600 ;
        RECT 697.950 469.950 700.050 470.400 ;
        RECT 718.950 469.950 721.050 470.400 ;
        RECT 766.950 471.600 769.050 472.050 ;
        RECT 772.950 471.600 775.050 472.050 ;
        RECT 766.950 470.400 775.050 471.600 ;
        RECT 766.950 469.950 769.050 470.400 ;
        RECT 772.950 469.950 775.050 470.400 ;
        RECT 391.950 468.600 394.050 469.050 ;
        RECT 359.400 467.400 394.050 468.600 ;
        RECT 232.950 466.950 235.050 467.400 ;
        RECT 355.950 466.950 358.050 467.400 ;
        RECT 391.950 466.950 394.050 467.400 ;
        RECT 397.950 468.600 400.050 469.050 ;
        RECT 478.950 468.600 481.050 469.050 ;
        RECT 520.950 468.600 523.050 469.050 ;
        RECT 397.950 467.400 477.600 468.600 ;
        RECT 397.950 466.950 400.050 467.400 ;
        RECT 217.950 465.600 220.050 466.050 ;
        RECT 247.950 465.600 250.050 466.050 ;
        RECT 217.950 464.400 250.050 465.600 ;
        RECT 217.950 463.950 220.050 464.400 ;
        RECT 247.950 463.950 250.050 464.400 ;
        RECT 265.950 465.600 268.050 466.050 ;
        RECT 274.950 465.600 277.050 466.050 ;
        RECT 265.950 464.400 277.050 465.600 ;
        RECT 265.950 463.950 268.050 464.400 ;
        RECT 274.950 463.950 277.050 464.400 ;
        RECT 376.950 465.600 379.050 466.050 ;
        RECT 394.950 465.600 397.050 466.050 ;
        RECT 376.950 464.400 397.050 465.600 ;
        RECT 376.950 463.950 379.050 464.400 ;
        RECT 394.950 463.950 397.050 464.400 ;
        RECT 451.950 465.600 454.050 466.050 ;
        RECT 463.950 465.600 466.050 466.050 ;
        RECT 451.950 464.400 466.050 465.600 ;
        RECT 476.400 465.600 477.600 467.400 ;
        RECT 478.950 467.400 523.050 468.600 ;
        RECT 478.950 466.950 481.050 467.400 ;
        RECT 520.950 466.950 523.050 467.400 ;
        RECT 580.950 468.600 583.050 469.050 ;
        RECT 667.950 468.600 670.050 469.050 ;
        RECT 580.950 467.400 670.050 468.600 ;
        RECT 580.950 466.950 583.050 467.400 ;
        RECT 667.950 466.950 670.050 467.400 ;
        RECT 673.950 468.600 676.050 469.050 ;
        RECT 820.950 468.600 823.050 469.050 ;
        RECT 673.950 467.400 823.050 468.600 ;
        RECT 673.950 466.950 676.050 467.400 ;
        RECT 820.950 466.950 823.050 467.400 ;
        RECT 490.950 465.600 493.050 466.050 ;
        RECT 476.400 464.400 493.050 465.600 ;
        RECT 451.950 463.950 454.050 464.400 ;
        RECT 463.950 463.950 466.050 464.400 ;
        RECT 490.950 463.950 493.050 464.400 ;
        RECT 169.950 462.600 172.050 463.050 ;
        RECT 226.950 462.600 229.050 463.050 ;
        RECT 169.950 461.400 229.050 462.600 ;
        RECT 169.950 460.950 172.050 461.400 ;
        RECT 226.950 460.950 229.050 461.400 ;
        RECT 238.950 462.600 241.050 463.050 ;
        RECT 244.950 462.600 247.050 463.050 ;
        RECT 238.950 461.400 247.050 462.600 ;
        RECT 238.950 460.950 241.050 461.400 ;
        RECT 244.950 460.950 247.050 461.400 ;
        RECT 262.950 462.600 265.050 463.050 ;
        RECT 277.950 462.600 280.050 463.050 ;
        RECT 262.950 461.400 280.050 462.600 ;
        RECT 262.950 460.950 265.050 461.400 ;
        RECT 277.950 460.950 280.050 461.400 ;
        RECT 280.950 462.600 283.050 463.050 ;
        RECT 316.950 462.600 319.050 463.050 ;
        RECT 325.950 462.600 328.050 463.050 ;
        RECT 280.950 461.400 328.050 462.600 ;
        RECT 280.950 460.950 283.050 461.400 ;
        RECT 316.950 460.950 319.050 461.400 ;
        RECT 325.950 460.950 328.050 461.400 ;
        RECT 364.950 462.600 367.050 463.050 ;
        RECT 388.950 462.600 391.050 463.050 ;
        RECT 364.950 461.400 391.050 462.600 ;
        RECT 364.950 460.950 367.050 461.400 ;
        RECT 388.950 460.950 391.050 461.400 ;
        RECT 403.950 462.600 406.050 463.050 ;
        RECT 442.950 462.600 445.050 463.050 ;
        RECT 403.950 461.400 445.050 462.600 ;
        RECT 403.950 460.950 406.050 461.400 ;
        RECT 442.950 460.950 445.050 461.400 ;
        RECT 460.950 462.600 463.050 463.050 ;
        RECT 466.950 462.600 469.050 463.050 ;
        RECT 460.950 461.400 469.050 462.600 ;
        RECT 460.950 460.950 463.050 461.400 ;
        RECT 466.950 460.950 469.050 461.400 ;
        RECT 484.950 462.600 487.050 463.050 ;
        RECT 496.950 462.600 499.050 463.050 ;
        RECT 484.950 461.400 499.050 462.600 ;
        RECT 484.950 460.950 487.050 461.400 ;
        RECT 496.950 460.950 499.050 461.400 ;
        RECT 598.950 462.600 601.050 463.050 ;
        RECT 652.950 462.600 655.050 463.050 ;
        RECT 598.950 461.400 655.050 462.600 ;
        RECT 598.950 460.950 601.050 461.400 ;
        RECT 652.950 460.950 655.050 461.400 ;
        RECT 58.950 459.600 61.050 460.050 ;
        RECT 88.950 459.600 91.050 460.050 ;
        RECT 58.950 458.400 91.050 459.600 ;
        RECT 58.950 457.950 61.050 458.400 ;
        RECT 88.950 457.950 91.050 458.400 ;
        RECT 91.950 459.600 94.050 460.050 ;
        RECT 109.950 459.600 112.050 460.050 ;
        RECT 91.950 458.400 112.050 459.600 ;
        RECT 91.950 457.950 94.050 458.400 ;
        RECT 109.950 457.950 112.050 458.400 ;
        RECT 223.950 459.600 226.050 460.050 ;
        RECT 244.950 459.600 247.050 460.050 ;
        RECT 223.950 458.400 247.050 459.600 ;
        RECT 223.950 457.950 226.050 458.400 ;
        RECT 244.950 457.950 247.050 458.400 ;
        RECT 256.950 459.600 259.050 460.050 ;
        RECT 265.950 459.600 268.050 460.050 ;
        RECT 268.950 459.600 271.050 460.050 ;
        RECT 289.950 459.600 292.050 460.050 ;
        RECT 298.950 459.600 301.050 460.050 ;
        RECT 256.950 458.400 301.050 459.600 ;
        RECT 256.950 457.950 259.050 458.400 ;
        RECT 265.950 457.950 268.050 458.400 ;
        RECT 268.950 457.950 271.050 458.400 ;
        RECT 289.950 457.950 292.050 458.400 ;
        RECT 298.950 457.950 301.050 458.400 ;
        RECT 307.950 459.600 310.050 460.050 ;
        RECT 352.950 459.600 355.050 460.050 ;
        RECT 358.950 459.600 361.050 460.050 ;
        RECT 307.950 458.400 361.050 459.600 ;
        RECT 307.950 457.950 310.050 458.400 ;
        RECT 352.950 457.950 355.050 458.400 ;
        RECT 358.950 457.950 361.050 458.400 ;
        RECT 361.950 459.600 364.050 460.050 ;
        RECT 376.950 459.600 379.050 460.050 ;
        RECT 361.950 458.400 379.050 459.600 ;
        RECT 361.950 457.950 364.050 458.400 ;
        RECT 376.950 457.950 379.050 458.400 ;
        RECT 391.950 459.600 394.050 460.050 ;
        RECT 424.950 459.600 427.050 460.050 ;
        RECT 430.950 459.600 433.050 460.050 ;
        RECT 454.950 459.600 457.050 460.050 ;
        RECT 475.950 459.600 478.050 460.050 ;
        RECT 484.950 459.600 487.050 460.050 ;
        RECT 391.950 458.400 420.600 459.600 ;
        RECT 391.950 457.950 394.050 458.400 ;
        RECT 10.950 456.600 13.050 457.050 ;
        RECT 34.950 456.600 37.050 457.050 ;
        RECT 37.950 456.600 40.050 457.050 ;
        RECT 10.950 455.400 40.050 456.600 ;
        RECT 10.950 454.950 13.050 455.400 ;
        RECT 34.950 454.950 37.050 455.400 ;
        RECT 37.950 454.950 40.050 455.400 ;
        RECT 43.950 456.600 46.050 457.050 ;
        RECT 55.950 456.600 58.050 457.050 ;
        RECT 43.950 455.400 58.050 456.600 ;
        RECT 43.950 454.950 46.050 455.400 ;
        RECT 55.950 454.950 58.050 455.400 ;
        RECT 64.950 456.600 67.050 457.050 ;
        RECT 70.950 456.600 73.050 457.050 ;
        RECT 85.950 456.600 88.050 457.050 ;
        RECT 64.950 455.400 88.050 456.600 ;
        RECT 64.950 454.950 67.050 455.400 ;
        RECT 70.950 454.950 73.050 455.400 ;
        RECT 85.950 454.950 88.050 455.400 ;
        RECT 241.950 456.600 244.050 457.050 ;
        RECT 253.950 456.600 256.050 457.050 ;
        RECT 286.950 456.600 289.050 457.050 ;
        RECT 241.950 455.400 289.050 456.600 ;
        RECT 241.950 454.950 244.050 455.400 ;
        RECT 253.950 454.950 256.050 455.400 ;
        RECT 286.950 454.950 289.050 455.400 ;
        RECT 319.950 454.950 322.050 457.050 ;
        RECT 322.950 456.600 325.050 457.050 ;
        RECT 346.950 456.600 349.050 457.050 ;
        RECT 322.950 455.400 349.050 456.600 ;
        RECT 322.950 454.950 325.050 455.400 ;
        RECT 346.950 454.950 349.050 455.400 ;
        RECT 349.950 456.600 352.050 457.050 ;
        RECT 367.950 456.600 370.050 457.050 ;
        RECT 349.950 455.400 370.050 456.600 ;
        RECT 349.950 454.950 352.050 455.400 ;
        RECT 367.950 454.950 370.050 455.400 ;
        RECT 370.950 456.600 373.050 457.050 ;
        RECT 385.950 456.600 388.050 457.050 ;
        RECT 370.950 455.400 388.050 456.600 ;
        RECT 370.950 454.950 373.050 455.400 ;
        RECT 385.950 454.950 388.050 455.400 ;
        RECT 394.950 456.600 397.050 457.050 ;
        RECT 415.950 456.600 418.050 457.050 ;
        RECT 394.950 455.400 418.050 456.600 ;
        RECT 419.400 456.600 420.600 458.400 ;
        RECT 424.950 458.400 433.050 459.600 ;
        RECT 424.950 457.950 427.050 458.400 ;
        RECT 430.950 457.950 433.050 458.400 ;
        RECT 434.400 458.400 487.050 459.600 ;
        RECT 434.400 456.600 435.600 458.400 ;
        RECT 454.950 457.950 457.050 458.400 ;
        RECT 475.950 457.950 478.050 458.400 ;
        RECT 484.950 457.950 487.050 458.400 ;
        RECT 517.950 459.600 520.050 460.050 ;
        RECT 526.950 459.600 529.050 460.050 ;
        RECT 517.950 458.400 529.050 459.600 ;
        RECT 517.950 457.950 520.050 458.400 ;
        RECT 526.950 457.950 529.050 458.400 ;
        RECT 553.950 459.600 556.050 460.050 ;
        RECT 559.950 459.600 562.050 460.050 ;
        RECT 553.950 458.400 562.050 459.600 ;
        RECT 553.950 457.950 556.050 458.400 ;
        RECT 559.950 457.950 562.050 458.400 ;
        RECT 562.950 459.600 565.050 460.050 ;
        RECT 571.950 459.600 574.050 460.050 ;
        RECT 631.950 459.600 634.050 460.050 ;
        RECT 562.950 458.400 634.050 459.600 ;
        RECT 562.950 457.950 565.050 458.400 ;
        RECT 571.950 457.950 574.050 458.400 ;
        RECT 631.950 457.950 634.050 458.400 ;
        RECT 637.950 459.600 640.050 460.050 ;
        RECT 646.950 459.600 649.050 460.050 ;
        RECT 637.950 458.400 649.050 459.600 ;
        RECT 637.950 457.950 640.050 458.400 ;
        RECT 646.950 457.950 649.050 458.400 ;
        RECT 700.950 459.600 703.050 460.050 ;
        RECT 724.950 459.600 727.050 460.050 ;
        RECT 700.950 458.400 727.050 459.600 ;
        RECT 700.950 457.950 703.050 458.400 ;
        RECT 724.950 457.950 727.050 458.400 ;
        RECT 733.950 459.600 736.050 460.050 ;
        RECT 739.950 459.600 742.050 460.050 ;
        RECT 733.950 458.400 742.050 459.600 ;
        RECT 733.950 457.950 736.050 458.400 ;
        RECT 739.950 457.950 742.050 458.400 ;
        RECT 760.950 459.600 763.050 460.050 ;
        RECT 817.950 459.600 820.050 460.050 ;
        RECT 760.950 458.400 820.050 459.600 ;
        RECT 760.950 457.950 763.050 458.400 ;
        RECT 817.950 457.950 820.050 458.400 ;
        RECT 419.400 455.400 435.600 456.600 ;
        RECT 439.950 456.600 442.050 457.050 ;
        RECT 445.950 456.600 448.050 457.050 ;
        RECT 439.950 455.400 448.050 456.600 ;
        RECT 394.950 454.950 397.050 455.400 ;
        RECT 415.950 454.950 418.050 455.400 ;
        RECT 439.950 454.950 442.050 455.400 ;
        RECT 445.950 454.950 448.050 455.400 ;
        RECT 454.950 454.950 457.050 457.050 ;
        RECT 460.950 456.600 463.050 457.050 ;
        RECT 496.950 456.600 499.050 457.050 ;
        RECT 499.950 456.600 502.050 457.050 ;
        RECT 526.950 456.600 529.050 457.050 ;
        RECT 460.950 455.400 495.600 456.600 ;
        RECT 460.950 454.950 463.050 455.400 ;
        RECT 61.950 453.600 64.050 454.050 ;
        RECT 79.950 453.600 82.050 454.050 ;
        RECT 61.950 452.400 82.050 453.600 ;
        RECT 61.950 451.950 64.050 452.400 ;
        RECT 79.950 451.950 82.050 452.400 ;
        RECT 97.950 453.600 100.050 454.050 ;
        RECT 103.950 453.600 106.050 454.050 ;
        RECT 97.950 452.400 106.050 453.600 ;
        RECT 97.950 451.950 100.050 452.400 ;
        RECT 103.950 451.950 106.050 452.400 ;
        RECT 124.950 453.600 127.050 454.050 ;
        RECT 199.950 453.600 202.050 454.050 ;
        RECT 124.950 452.400 202.050 453.600 ;
        RECT 124.950 451.950 127.050 452.400 ;
        RECT 199.950 451.950 202.050 452.400 ;
        RECT 208.950 453.600 211.050 454.050 ;
        RECT 241.950 453.600 244.050 454.050 ;
        RECT 295.950 453.600 298.050 454.050 ;
        RECT 208.950 452.400 244.050 453.600 ;
        RECT 208.950 451.950 211.050 452.400 ;
        RECT 241.950 451.950 244.050 452.400 ;
        RECT 290.400 452.400 298.050 453.600 ;
        RECT 13.950 450.600 16.050 451.050 ;
        RECT 31.950 450.600 34.050 451.050 ;
        RECT 13.950 449.400 34.050 450.600 ;
        RECT 13.950 448.950 16.050 449.400 ;
        RECT 31.950 448.950 34.050 449.400 ;
        RECT 40.950 450.600 43.050 451.050 ;
        RECT 49.950 450.600 52.050 451.050 ;
        RECT 40.950 449.400 52.050 450.600 ;
        RECT 40.950 448.950 43.050 449.400 ;
        RECT 49.950 448.950 52.050 449.400 ;
        RECT 94.950 450.600 97.050 451.050 ;
        RECT 106.950 450.600 109.050 451.050 ;
        RECT 94.950 449.400 109.050 450.600 ;
        RECT 94.950 448.950 97.050 449.400 ;
        RECT 106.950 448.950 109.050 449.400 ;
        RECT 127.950 450.600 130.050 451.050 ;
        RECT 145.950 450.600 148.050 451.050 ;
        RECT 127.950 449.400 148.050 450.600 ;
        RECT 127.950 448.950 130.050 449.400 ;
        RECT 145.950 448.950 148.050 449.400 ;
        RECT 238.950 450.600 241.050 451.050 ;
        RECT 247.950 450.600 250.050 451.050 ;
        RECT 238.950 449.400 250.050 450.600 ;
        RECT 238.950 448.950 241.050 449.400 ;
        RECT 247.950 448.950 250.050 449.400 ;
        RECT 277.950 450.600 280.050 451.050 ;
        RECT 290.400 450.600 291.600 452.400 ;
        RECT 295.950 451.950 298.050 452.400 ;
        RECT 313.950 453.600 316.050 454.050 ;
        RECT 320.400 453.600 321.600 454.950 ;
        RECT 364.950 453.600 367.050 454.050 ;
        RECT 395.400 453.600 396.600 454.950 ;
        RECT 313.950 452.400 336.600 453.600 ;
        RECT 313.950 451.950 316.050 452.400 ;
        RECT 277.950 449.400 291.600 450.600 ;
        RECT 292.950 450.600 295.050 451.050 ;
        RECT 301.950 450.600 304.050 451.050 ;
        RECT 292.950 449.400 304.050 450.600 ;
        RECT 277.950 448.950 280.050 449.400 ;
        RECT 292.950 448.950 295.050 449.400 ;
        RECT 301.950 448.950 304.050 449.400 ;
        RECT 307.950 450.600 310.050 451.050 ;
        RECT 319.950 450.600 322.050 451.050 ;
        RECT 307.950 449.400 322.050 450.600 ;
        RECT 307.950 448.950 310.050 449.400 ;
        RECT 319.950 448.950 322.050 449.400 ;
        RECT 325.950 450.600 328.050 451.050 ;
        RECT 331.950 450.600 334.050 451.050 ;
        RECT 325.950 449.400 334.050 450.600 ;
        RECT 335.400 450.600 336.600 452.400 ;
        RECT 364.950 452.400 396.600 453.600 ;
        RECT 409.950 453.600 412.050 454.050 ;
        RECT 412.950 453.600 415.050 454.050 ;
        RECT 433.950 453.600 436.050 454.050 ;
        RECT 455.400 453.600 456.600 454.950 ;
        RECT 409.950 452.400 456.600 453.600 ;
        RECT 463.950 453.600 466.050 454.050 ;
        RECT 478.950 453.600 481.050 454.050 ;
        RECT 463.950 452.400 481.050 453.600 ;
        RECT 494.400 453.600 495.600 455.400 ;
        RECT 496.950 455.400 529.050 456.600 ;
        RECT 496.950 454.950 499.050 455.400 ;
        RECT 499.950 454.950 502.050 455.400 ;
        RECT 526.950 454.950 529.050 455.400 ;
        RECT 532.950 454.950 535.050 457.050 ;
        RECT 643.950 456.600 646.050 457.050 ;
        RECT 655.950 456.600 658.050 457.050 ;
        RECT 676.950 456.600 679.050 457.050 ;
        RECT 643.950 455.400 679.050 456.600 ;
        RECT 643.950 454.950 646.050 455.400 ;
        RECT 655.950 454.950 658.050 455.400 ;
        RECT 676.950 454.950 679.050 455.400 ;
        RECT 679.950 456.600 682.050 457.050 ;
        RECT 691.950 456.600 694.050 457.050 ;
        RECT 679.950 455.400 694.050 456.600 ;
        RECT 679.950 454.950 682.050 455.400 ;
        RECT 691.950 454.950 694.050 455.400 ;
        RECT 730.950 456.600 733.050 457.050 ;
        RECT 751.950 456.600 754.050 457.050 ;
        RECT 730.950 455.400 754.050 456.600 ;
        RECT 730.950 454.950 733.050 455.400 ;
        RECT 751.950 454.950 754.050 455.400 ;
        RECT 508.950 453.600 511.050 454.050 ;
        RECT 494.400 452.400 511.050 453.600 ;
        RECT 364.950 451.950 367.050 452.400 ;
        RECT 409.950 451.950 412.050 452.400 ;
        RECT 412.950 451.950 415.050 452.400 ;
        RECT 433.950 451.950 436.050 452.400 ;
        RECT 463.950 451.950 466.050 452.400 ;
        RECT 478.950 451.950 481.050 452.400 ;
        RECT 508.950 451.950 511.050 452.400 ;
        RECT 511.950 453.600 514.050 454.050 ;
        RECT 511.950 452.400 531.600 453.600 ;
        RECT 511.950 451.950 514.050 452.400 ;
        RECT 530.400 451.050 531.600 452.400 ;
        RECT 337.950 450.600 340.050 451.050 ;
        RECT 335.400 449.400 340.050 450.600 ;
        RECT 325.950 448.950 328.050 449.400 ;
        RECT 331.950 448.950 334.050 449.400 ;
        RECT 337.950 448.950 340.050 449.400 ;
        RECT 343.950 450.600 346.050 451.050 ;
        RECT 355.950 450.600 358.050 451.050 ;
        RECT 343.950 449.400 358.050 450.600 ;
        RECT 343.950 448.950 346.050 449.400 ;
        RECT 355.950 448.950 358.050 449.400 ;
        RECT 409.950 450.600 412.050 451.050 ;
        RECT 427.950 450.600 430.050 451.050 ;
        RECT 409.950 449.400 430.050 450.600 ;
        RECT 409.950 448.950 412.050 449.400 ;
        RECT 427.950 448.950 430.050 449.400 ;
        RECT 493.950 450.600 496.050 451.050 ;
        RECT 502.950 450.600 505.050 451.050 ;
        RECT 493.950 449.400 505.050 450.600 ;
        RECT 493.950 448.950 496.050 449.400 ;
        RECT 502.950 448.950 505.050 449.400 ;
        RECT 514.950 450.600 517.050 451.050 ;
        RECT 520.950 450.600 523.050 451.050 ;
        RECT 514.950 449.400 523.050 450.600 ;
        RECT 514.950 448.950 517.050 449.400 ;
        RECT 520.950 448.950 523.050 449.400 ;
        RECT 529.950 448.950 532.050 451.050 ;
        RECT 7.950 447.600 10.050 448.050 ;
        RECT 19.950 447.600 22.050 448.050 ;
        RECT 22.950 447.600 25.050 448.050 ;
        RECT 7.950 446.400 25.050 447.600 ;
        RECT 7.950 445.950 10.050 446.400 ;
        RECT 19.950 445.950 22.050 446.400 ;
        RECT 22.950 445.950 25.050 446.400 ;
        RECT 190.950 447.600 193.050 448.050 ;
        RECT 196.950 447.600 199.050 448.050 ;
        RECT 190.950 446.400 199.050 447.600 ;
        RECT 190.950 445.950 193.050 446.400 ;
        RECT 196.950 445.950 199.050 446.400 ;
        RECT 298.950 447.600 301.050 448.050 ;
        RECT 310.950 447.600 313.050 448.050 ;
        RECT 364.950 447.600 367.050 448.050 ;
        RECT 298.950 446.400 367.050 447.600 ;
        RECT 298.950 445.950 301.050 446.400 ;
        RECT 310.950 445.950 313.050 446.400 ;
        RECT 364.950 445.950 367.050 446.400 ;
        RECT 379.950 447.600 382.050 448.050 ;
        RECT 436.950 447.600 439.050 448.050 ;
        RECT 379.950 446.400 439.050 447.600 ;
        RECT 379.950 445.950 382.050 446.400 ;
        RECT 436.950 445.950 439.050 446.400 ;
        RECT 457.950 447.600 460.050 448.050 ;
        RECT 472.950 447.600 475.050 448.050 ;
        RECT 457.950 446.400 475.050 447.600 ;
        RECT 457.950 445.950 460.050 446.400 ;
        RECT 472.950 445.950 475.050 446.400 ;
        RECT 499.950 447.600 502.050 448.050 ;
        RECT 505.950 447.600 508.050 448.050 ;
        RECT 499.950 446.400 508.050 447.600 ;
        RECT 499.950 445.950 502.050 446.400 ;
        RECT 505.950 445.950 508.050 446.400 ;
        RECT 526.950 447.600 529.050 448.050 ;
        RECT 530.400 447.600 531.600 448.950 ;
        RECT 533.400 448.050 534.600 454.950 ;
        RECT 616.950 453.600 619.050 454.050 ;
        RECT 631.950 453.600 634.050 454.050 ;
        RECT 616.950 452.400 634.050 453.600 ;
        RECT 616.950 451.950 619.050 452.400 ;
        RECT 631.950 451.950 634.050 452.400 ;
        RECT 649.950 453.600 652.050 454.050 ;
        RECT 670.950 453.600 673.050 454.050 ;
        RECT 649.950 452.400 673.050 453.600 ;
        RECT 649.950 451.950 652.050 452.400 ;
        RECT 670.950 451.950 673.050 452.400 ;
        RECT 688.950 453.600 691.050 454.050 ;
        RECT 709.950 453.600 712.050 454.050 ;
        RECT 727.950 453.600 730.050 454.050 ;
        RECT 688.950 452.400 730.050 453.600 ;
        RECT 688.950 451.950 691.050 452.400 ;
        RECT 709.950 451.950 712.050 452.400 ;
        RECT 727.950 451.950 730.050 452.400 ;
        RECT 733.950 453.600 736.050 454.050 ;
        RECT 745.950 453.600 748.050 454.050 ;
        RECT 733.950 452.400 748.050 453.600 ;
        RECT 733.950 451.950 736.050 452.400 ;
        RECT 745.950 451.950 748.050 452.400 ;
        RECT 766.950 453.600 769.050 454.050 ;
        RECT 778.950 453.600 781.050 454.050 ;
        RECT 766.950 452.400 781.050 453.600 ;
        RECT 766.950 451.950 769.050 452.400 ;
        RECT 778.950 451.950 781.050 452.400 ;
        RECT 712.950 450.600 715.050 451.050 ;
        RECT 724.950 450.600 727.050 451.050 ;
        RECT 712.950 449.400 727.050 450.600 ;
        RECT 712.950 448.950 715.050 449.400 ;
        RECT 724.950 448.950 727.050 449.400 ;
        RECT 754.950 450.600 757.050 451.050 ;
        RECT 763.950 450.600 766.050 451.050 ;
        RECT 769.950 450.600 772.050 451.050 ;
        RECT 754.950 449.400 772.050 450.600 ;
        RECT 754.950 448.950 757.050 449.400 ;
        RECT 763.950 448.950 766.050 449.400 ;
        RECT 769.950 448.950 772.050 449.400 ;
        RECT 526.950 446.400 531.600 447.600 ;
        RECT 526.950 445.950 529.050 446.400 ;
        RECT 532.950 445.950 535.050 448.050 ;
        RECT 616.950 447.600 619.050 448.050 ;
        RECT 661.950 447.600 664.050 448.050 ;
        RECT 616.950 446.400 664.050 447.600 ;
        RECT 616.950 445.950 619.050 446.400 ;
        RECT 661.950 445.950 664.050 446.400 ;
        RECT 718.950 447.600 721.050 448.050 ;
        RECT 733.950 447.600 736.050 448.050 ;
        RECT 763.950 447.600 766.050 448.050 ;
        RECT 718.950 446.400 766.050 447.600 ;
        RECT 718.950 445.950 721.050 446.400 ;
        RECT 733.950 445.950 736.050 446.400 ;
        RECT 763.950 445.950 766.050 446.400 ;
        RECT 835.950 447.600 838.050 448.050 ;
        RECT 856.950 447.600 859.050 448.050 ;
        RECT 835.950 446.400 859.050 447.600 ;
        RECT 835.950 445.950 838.050 446.400 ;
        RECT 856.950 445.950 859.050 446.400 ;
        RECT 136.950 444.600 139.050 445.050 ;
        RECT 256.950 444.600 259.050 445.050 ;
        RECT 136.950 443.400 259.050 444.600 ;
        RECT 136.950 442.950 139.050 443.400 ;
        RECT 256.950 442.950 259.050 443.400 ;
        RECT 271.950 444.600 274.050 445.050 ;
        RECT 385.950 444.600 388.050 445.050 ;
        RECT 415.950 444.600 418.050 445.050 ;
        RECT 271.950 443.400 418.050 444.600 ;
        RECT 271.950 442.950 274.050 443.400 ;
        RECT 385.950 442.950 388.050 443.400 ;
        RECT 415.950 442.950 418.050 443.400 ;
        RECT 502.950 444.600 505.050 445.050 ;
        RECT 511.950 444.600 514.050 445.050 ;
        RECT 502.950 443.400 514.050 444.600 ;
        RECT 502.950 442.950 505.050 443.400 ;
        RECT 511.950 442.950 514.050 443.400 ;
        RECT 718.950 444.600 721.050 445.050 ;
        RECT 757.950 444.600 760.050 445.050 ;
        RECT 718.950 443.400 760.050 444.600 ;
        RECT 718.950 442.950 721.050 443.400 ;
        RECT 757.950 442.950 760.050 443.400 ;
        RECT 7.950 441.600 10.050 442.050 ;
        RECT 16.950 441.600 19.050 442.050 ;
        RECT 88.950 441.600 91.050 442.050 ;
        RECT 97.950 441.600 100.050 442.050 ;
        RECT 7.950 440.400 100.050 441.600 ;
        RECT 7.950 439.950 10.050 440.400 ;
        RECT 16.950 439.950 19.050 440.400 ;
        RECT 88.950 439.950 91.050 440.400 ;
        RECT 97.950 439.950 100.050 440.400 ;
        RECT 292.950 441.600 295.050 442.050 ;
        RECT 304.950 441.600 307.050 442.050 ;
        RECT 292.950 440.400 307.050 441.600 ;
        RECT 292.950 439.950 295.050 440.400 ;
        RECT 304.950 439.950 307.050 440.400 ;
        RECT 307.950 441.600 310.050 442.050 ;
        RECT 316.950 441.600 319.050 442.050 ;
        RECT 307.950 440.400 319.050 441.600 ;
        RECT 307.950 439.950 310.050 440.400 ;
        RECT 316.950 439.950 319.050 440.400 ;
        RECT 346.950 441.600 349.050 442.050 ;
        RECT 424.950 441.600 427.050 442.050 ;
        RECT 346.950 440.400 427.050 441.600 ;
        RECT 346.950 439.950 349.050 440.400 ;
        RECT 424.950 439.950 427.050 440.400 ;
        RECT 64.950 438.600 67.050 439.050 ;
        RECT 118.950 438.600 121.050 439.050 ;
        RECT 181.950 438.600 184.050 439.050 ;
        RECT 64.950 437.400 184.050 438.600 ;
        RECT 64.950 436.950 67.050 437.400 ;
        RECT 118.950 436.950 121.050 437.400 ;
        RECT 181.950 436.950 184.050 437.400 ;
        RECT 184.950 438.600 187.050 439.050 ;
        RECT 220.950 438.600 223.050 439.050 ;
        RECT 184.950 437.400 223.050 438.600 ;
        RECT 184.950 436.950 187.050 437.400 ;
        RECT 220.950 436.950 223.050 437.400 ;
        RECT 247.950 438.600 250.050 439.050 ;
        RECT 256.950 438.600 259.050 439.050 ;
        RECT 247.950 437.400 259.050 438.600 ;
        RECT 247.950 436.950 250.050 437.400 ;
        RECT 256.950 436.950 259.050 437.400 ;
        RECT 289.950 438.600 292.050 439.050 ;
        RECT 340.950 438.600 343.050 439.050 ;
        RECT 343.950 438.600 346.050 439.050 ;
        RECT 415.950 438.600 418.050 439.050 ;
        RECT 637.950 438.600 640.050 439.050 ;
        RECT 736.950 438.600 739.050 439.050 ;
        RECT 289.950 437.400 346.050 438.600 ;
        RECT 289.950 436.950 292.050 437.400 ;
        RECT 340.950 436.950 343.050 437.400 ;
        RECT 343.950 436.950 346.050 437.400 ;
        RECT 347.400 437.400 393.600 438.600 ;
        RECT 175.950 435.600 178.050 436.050 ;
        RECT 214.950 435.600 217.050 436.050 ;
        RECT 175.950 434.400 217.050 435.600 ;
        RECT 175.950 433.950 178.050 434.400 ;
        RECT 214.950 433.950 217.050 434.400 ;
        RECT 250.950 435.600 253.050 436.050 ;
        RECT 347.400 435.600 348.600 437.400 ;
        RECT 250.950 434.400 348.600 435.600 ;
        RECT 361.950 435.600 364.050 436.050 ;
        RECT 388.950 435.600 391.050 436.050 ;
        RECT 361.950 434.400 391.050 435.600 ;
        RECT 392.400 435.600 393.600 437.400 ;
        RECT 415.950 437.400 739.050 438.600 ;
        RECT 415.950 436.950 418.050 437.400 ;
        RECT 637.950 436.950 640.050 437.400 ;
        RECT 736.950 436.950 739.050 437.400 ;
        RECT 550.950 435.600 553.050 436.050 ;
        RECT 392.400 434.400 553.050 435.600 ;
        RECT 250.950 433.950 253.050 434.400 ;
        RECT 361.950 433.950 364.050 434.400 ;
        RECT 388.950 433.950 391.050 434.400 ;
        RECT 550.950 433.950 553.050 434.400 ;
        RECT 562.950 435.600 565.050 436.050 ;
        RECT 574.950 435.600 577.050 436.050 ;
        RECT 586.950 435.600 589.050 436.050 ;
        RECT 562.950 434.400 589.050 435.600 ;
        RECT 562.950 433.950 565.050 434.400 ;
        RECT 574.950 433.950 577.050 434.400 ;
        RECT 586.950 433.950 589.050 434.400 ;
        RECT 229.950 432.600 232.050 433.050 ;
        RECT 235.950 432.600 238.050 433.050 ;
        RECT 280.950 432.600 283.050 433.050 ;
        RECT 229.950 431.400 283.050 432.600 ;
        RECT 229.950 430.950 232.050 431.400 ;
        RECT 235.950 430.950 238.050 431.400 ;
        RECT 280.950 430.950 283.050 431.400 ;
        RECT 304.950 432.600 307.050 433.050 ;
        RECT 322.950 432.600 325.050 433.050 ;
        RECT 304.950 431.400 325.050 432.600 ;
        RECT 304.950 430.950 307.050 431.400 ;
        RECT 322.950 430.950 325.050 431.400 ;
        RECT 358.950 432.600 361.050 433.050 ;
        RECT 448.950 432.600 451.050 433.050 ;
        RECT 358.950 431.400 451.050 432.600 ;
        RECT 358.950 430.950 361.050 431.400 ;
        RECT 448.950 430.950 451.050 431.400 ;
        RECT 217.950 429.600 220.050 430.050 ;
        RECT 247.950 429.600 250.050 430.050 ;
        RECT 217.950 428.400 250.050 429.600 ;
        RECT 217.950 427.950 220.050 428.400 ;
        RECT 247.950 427.950 250.050 428.400 ;
        RECT 325.950 429.600 328.050 430.050 ;
        RECT 340.950 429.600 343.050 430.050 ;
        RECT 364.950 429.600 367.050 430.050 ;
        RECT 379.950 429.600 382.050 430.050 ;
        RECT 325.950 428.400 382.050 429.600 ;
        RECT 325.950 427.950 328.050 428.400 ;
        RECT 340.950 427.950 343.050 428.400 ;
        RECT 364.950 427.950 367.050 428.400 ;
        RECT 379.950 427.950 382.050 428.400 ;
        RECT 682.950 429.600 685.050 430.050 ;
        RECT 736.950 429.600 739.050 430.050 ;
        RECT 682.950 428.400 739.050 429.600 ;
        RECT 682.950 427.950 685.050 428.400 ;
        RECT 736.950 427.950 739.050 428.400 ;
        RECT 31.950 426.600 34.050 427.050 ;
        RECT 100.950 426.600 103.050 427.050 ;
        RECT 31.950 425.400 103.050 426.600 ;
        RECT 31.950 424.950 34.050 425.400 ;
        RECT 100.950 424.950 103.050 425.400 ;
        RECT 283.950 426.600 286.050 427.050 ;
        RECT 298.950 426.600 301.050 427.050 ;
        RECT 283.950 425.400 301.050 426.600 ;
        RECT 283.950 424.950 286.050 425.400 ;
        RECT 298.950 424.950 301.050 425.400 ;
        RECT 373.950 426.600 376.050 427.050 ;
        RECT 379.950 426.600 382.050 427.050 ;
        RECT 373.950 425.400 382.050 426.600 ;
        RECT 373.950 424.950 376.050 425.400 ;
        RECT 379.950 424.950 382.050 425.400 ;
        RECT 424.950 426.600 427.050 427.050 ;
        RECT 484.950 426.600 487.050 427.050 ;
        RECT 424.950 425.400 487.050 426.600 ;
        RECT 424.950 424.950 427.050 425.400 ;
        RECT 484.950 424.950 487.050 425.400 ;
        RECT 733.950 426.600 736.050 427.050 ;
        RECT 742.950 426.600 745.050 427.050 ;
        RECT 733.950 425.400 745.050 426.600 ;
        RECT 733.950 424.950 736.050 425.400 ;
        RECT 742.950 424.950 745.050 425.400 ;
        RECT 49.950 423.600 52.050 424.050 ;
        RECT 97.950 423.600 100.050 424.050 ;
        RECT 49.950 422.400 100.050 423.600 ;
        RECT 49.950 421.950 52.050 422.400 ;
        RECT 97.950 421.950 100.050 422.400 ;
        RECT 127.950 423.600 130.050 424.050 ;
        RECT 133.950 423.600 136.050 424.050 ;
        RECT 136.950 423.600 139.050 424.050 ;
        RECT 127.950 422.400 139.050 423.600 ;
        RECT 127.950 421.950 130.050 422.400 ;
        RECT 133.950 421.950 136.050 422.400 ;
        RECT 136.950 421.950 139.050 422.400 ;
        RECT 253.950 423.600 256.050 424.050 ;
        RECT 295.950 423.600 298.050 424.050 ;
        RECT 346.950 423.600 349.050 424.050 ;
        RECT 376.950 423.600 379.050 424.050 ;
        RECT 253.950 422.400 349.050 423.600 ;
        RECT 253.950 421.950 256.050 422.400 ;
        RECT 295.950 421.950 298.050 422.400 ;
        RECT 346.950 421.950 349.050 422.400 ;
        RECT 350.400 422.400 379.050 423.600 ;
        RECT 61.950 420.600 64.050 421.050 ;
        RECT 67.950 420.600 70.050 421.050 ;
        RECT 61.950 419.400 70.050 420.600 ;
        RECT 61.950 418.950 64.050 419.400 ;
        RECT 67.950 418.950 70.050 419.400 ;
        RECT 100.950 420.600 103.050 421.050 ;
        RECT 103.950 420.600 106.050 421.050 ;
        RECT 136.950 420.600 139.050 421.050 ;
        RECT 100.950 419.400 139.050 420.600 ;
        RECT 100.950 418.950 103.050 419.400 ;
        RECT 103.950 418.950 106.050 419.400 ;
        RECT 136.950 418.950 139.050 419.400 ;
        RECT 244.950 420.600 247.050 421.050 ;
        RECT 274.950 420.600 277.050 421.050 ;
        RECT 244.950 419.400 277.050 420.600 ;
        RECT 244.950 418.950 247.050 419.400 ;
        RECT 274.950 418.950 277.050 419.400 ;
        RECT 304.950 418.950 307.050 421.050 ;
        RECT 331.950 420.600 334.050 421.050 ;
        RECT 350.400 420.600 351.600 422.400 ;
        RECT 376.950 421.950 379.050 422.400 ;
        RECT 481.950 423.600 484.050 424.050 ;
        RECT 499.950 423.600 502.050 424.050 ;
        RECT 481.950 422.400 502.050 423.600 ;
        RECT 481.950 421.950 484.050 422.400 ;
        RECT 499.950 421.950 502.050 422.400 ;
        RECT 326.400 419.400 334.050 420.600 ;
        RECT 46.950 417.600 49.050 418.050 ;
        RECT 58.950 417.600 61.050 418.050 ;
        RECT 46.950 416.400 61.050 417.600 ;
        RECT 46.950 415.950 49.050 416.400 ;
        RECT 58.950 415.950 61.050 416.400 ;
        RECT 73.950 417.600 76.050 418.050 ;
        RECT 82.950 417.600 85.050 418.050 ;
        RECT 73.950 416.400 85.050 417.600 ;
        RECT 73.950 415.950 76.050 416.400 ;
        RECT 82.950 415.950 85.050 416.400 ;
        RECT 118.950 417.600 121.050 418.050 ;
        RECT 124.950 417.600 127.050 418.050 ;
        RECT 118.950 416.400 127.050 417.600 ;
        RECT 118.950 415.950 121.050 416.400 ;
        RECT 124.950 415.950 127.050 416.400 ;
        RECT 130.950 417.600 133.050 418.050 ;
        RECT 172.950 417.600 175.050 418.050 ;
        RECT 178.950 417.600 181.050 418.050 ;
        RECT 130.950 416.400 156.600 417.600 ;
        RECT 130.950 415.950 133.050 416.400 ;
        RECT 22.950 414.600 25.050 415.050 ;
        RECT 34.950 414.600 37.050 415.050 ;
        RECT 22.950 413.400 37.050 414.600 ;
        RECT 22.950 412.950 25.050 413.400 ;
        RECT 34.950 412.950 37.050 413.400 ;
        RECT 43.950 414.600 46.050 415.050 ;
        RECT 49.950 414.600 52.050 415.050 ;
        RECT 43.950 413.400 52.050 414.600 ;
        RECT 43.950 412.950 46.050 413.400 ;
        RECT 49.950 412.950 52.050 413.400 ;
        RECT 58.950 414.600 61.050 415.050 ;
        RECT 148.950 414.600 151.050 415.050 ;
        RECT 151.950 414.600 154.050 415.050 ;
        RECT 58.950 413.400 154.050 414.600 ;
        RECT 155.400 414.600 156.600 416.400 ;
        RECT 172.950 416.400 181.050 417.600 ;
        RECT 172.950 415.950 175.050 416.400 ;
        RECT 178.950 415.950 181.050 416.400 ;
        RECT 181.950 417.600 184.050 418.050 ;
        RECT 199.950 417.600 202.050 418.050 ;
        RECT 277.950 417.600 280.050 418.050 ;
        RECT 301.950 417.600 304.050 418.050 ;
        RECT 181.950 416.400 280.050 417.600 ;
        RECT 181.950 415.950 184.050 416.400 ;
        RECT 199.950 415.950 202.050 416.400 ;
        RECT 169.950 414.600 172.050 415.050 ;
        RECT 155.400 413.400 172.050 414.600 ;
        RECT 251.400 414.600 252.600 416.400 ;
        RECT 277.950 415.950 280.050 416.400 ;
        RECT 284.400 416.400 304.050 417.600 ;
        RECT 262.950 414.600 265.050 415.050 ;
        RECT 251.400 413.400 265.050 414.600 ;
        RECT 58.950 412.950 61.050 413.400 ;
        RECT 148.950 412.950 151.050 413.400 ;
        RECT 151.950 412.950 154.050 413.400 ;
        RECT 169.950 412.950 172.050 413.400 ;
        RECT 262.950 412.950 265.050 413.400 ;
        RECT 265.950 414.600 268.050 415.050 ;
        RECT 274.950 414.600 277.050 415.050 ;
        RECT 265.950 413.400 277.050 414.600 ;
        RECT 265.950 412.950 268.050 413.400 ;
        RECT 274.950 412.950 277.050 413.400 ;
        RECT 284.400 412.050 285.600 416.400 ;
        RECT 301.950 415.950 304.050 416.400 ;
        RECT 305.400 415.050 306.600 418.950 ;
        RECT 289.950 414.600 292.050 415.050 ;
        RECT 289.950 413.400 303.600 414.600 ;
        RECT 289.950 412.950 292.050 413.400 ;
        RECT 13.950 411.600 16.050 412.050 ;
        RECT 19.950 411.600 22.050 412.050 ;
        RECT 13.950 410.400 22.050 411.600 ;
        RECT 13.950 409.950 16.050 410.400 ;
        RECT 19.950 409.950 22.050 410.400 ;
        RECT 25.950 411.600 28.050 412.050 ;
        RECT 52.950 411.600 55.050 412.050 ;
        RECT 25.950 410.400 55.050 411.600 ;
        RECT 25.950 409.950 28.050 410.400 ;
        RECT 52.950 409.950 55.050 410.400 ;
        RECT 55.950 411.600 58.050 412.050 ;
        RECT 70.950 411.600 73.050 412.050 ;
        RECT 55.950 410.400 73.050 411.600 ;
        RECT 55.950 409.950 58.050 410.400 ;
        RECT 70.950 409.950 73.050 410.400 ;
        RECT 82.950 411.600 85.050 412.050 ;
        RECT 91.950 411.600 94.050 412.050 ;
        RECT 82.950 410.400 94.050 411.600 ;
        RECT 82.950 409.950 85.050 410.400 ;
        RECT 91.950 409.950 94.050 410.400 ;
        RECT 106.950 411.600 109.050 412.050 ;
        RECT 121.950 411.600 124.050 412.050 ;
        RECT 106.950 410.400 124.050 411.600 ;
        RECT 106.950 409.950 109.050 410.400 ;
        RECT 121.950 409.950 124.050 410.400 ;
        RECT 133.950 411.600 136.050 412.050 ;
        RECT 139.950 411.600 142.050 412.050 ;
        RECT 163.950 411.600 166.050 412.050 ;
        RECT 133.950 410.400 142.050 411.600 ;
        RECT 133.950 409.950 136.050 410.400 ;
        RECT 139.950 409.950 142.050 410.400 ;
        RECT 143.400 410.400 166.050 411.600 ;
        RECT 25.950 408.600 28.050 409.050 ;
        RECT 37.950 408.600 40.050 409.050 ;
        RECT 61.950 408.600 64.050 409.050 ;
        RECT 25.950 407.400 64.050 408.600 ;
        RECT 25.950 406.950 28.050 407.400 ;
        RECT 37.950 406.950 40.050 407.400 ;
        RECT 61.950 406.950 64.050 407.400 ;
        RECT 124.950 408.600 127.050 409.050 ;
        RECT 143.400 408.600 144.600 410.400 ;
        RECT 163.950 409.950 166.050 410.400 ;
        RECT 166.950 411.600 169.050 412.050 ;
        RECT 172.950 411.600 175.050 412.050 ;
        RECT 166.950 410.400 175.050 411.600 ;
        RECT 166.950 409.950 169.050 410.400 ;
        RECT 172.950 409.950 175.050 410.400 ;
        RECT 247.950 411.600 250.050 412.050 ;
        RECT 253.950 411.600 256.050 412.050 ;
        RECT 277.950 411.600 280.050 412.050 ;
        RECT 247.950 410.400 256.050 411.600 ;
        RECT 247.950 409.950 250.050 410.400 ;
        RECT 253.950 409.950 256.050 410.400 ;
        RECT 260.400 410.400 280.050 411.600 ;
        RECT 124.950 407.400 144.600 408.600 ;
        RECT 145.950 408.600 148.050 409.050 ;
        RECT 151.950 408.600 154.050 409.050 ;
        RECT 145.950 407.400 154.050 408.600 ;
        RECT 124.950 406.950 127.050 407.400 ;
        RECT 145.950 406.950 148.050 407.400 ;
        RECT 151.950 406.950 154.050 407.400 ;
        RECT 220.950 408.600 223.050 409.050 ;
        RECT 260.400 408.600 261.600 410.400 ;
        RECT 277.950 409.950 280.050 410.400 ;
        RECT 283.950 409.950 286.050 412.050 ;
        RECT 302.400 411.600 303.600 413.400 ;
        RECT 304.950 412.950 307.050 415.050 ;
        RECT 326.400 414.600 327.600 419.400 ;
        RECT 331.950 418.950 334.050 419.400 ;
        RECT 347.400 419.400 351.600 420.600 ;
        RECT 358.950 420.600 361.050 421.050 ;
        RECT 391.950 420.600 394.050 421.050 ;
        RECT 406.950 420.600 409.050 421.050 ;
        RECT 412.950 420.600 415.050 421.050 ;
        RECT 358.950 419.400 405.600 420.600 ;
        RECT 328.950 417.600 331.050 418.050 ;
        RECT 328.950 416.400 342.600 417.600 ;
        RECT 328.950 415.950 331.050 416.400 ;
        RECT 337.950 414.600 340.050 415.050 ;
        RECT 326.400 413.400 340.050 414.600 ;
        RECT 337.950 412.950 340.050 413.400 ;
        RECT 341.400 412.050 342.600 416.400 ;
        RECT 347.400 415.050 348.600 419.400 ;
        RECT 358.950 418.950 361.050 419.400 ;
        RECT 391.950 418.950 394.050 419.400 ;
        RECT 355.950 417.600 358.050 418.050 ;
        RECT 364.950 417.600 367.050 418.050 ;
        RECT 370.950 417.600 373.050 418.050 ;
        RECT 355.950 416.400 363.600 417.600 ;
        RECT 355.950 415.950 358.050 416.400 ;
        RECT 346.950 412.950 349.050 415.050 ;
        RECT 362.400 414.600 363.600 416.400 ;
        RECT 364.950 416.400 373.050 417.600 ;
        RECT 364.950 415.950 367.050 416.400 ;
        RECT 370.950 415.950 373.050 416.400 ;
        RECT 376.950 417.600 379.050 418.050 ;
        RECT 385.950 417.600 388.050 418.050 ;
        RECT 376.950 416.400 388.050 417.600 ;
        RECT 404.400 417.600 405.600 419.400 ;
        RECT 406.950 419.400 415.050 420.600 ;
        RECT 406.950 418.950 409.050 419.400 ;
        RECT 412.950 418.950 415.050 419.400 ;
        RECT 460.950 420.600 463.050 421.050 ;
        RECT 466.950 420.600 469.050 421.050 ;
        RECT 460.950 419.400 469.050 420.600 ;
        RECT 460.950 418.950 463.050 419.400 ;
        RECT 466.950 418.950 469.050 419.400 ;
        RECT 481.950 420.600 484.050 421.050 ;
        RECT 487.950 420.600 490.050 421.050 ;
        RECT 523.950 420.600 526.050 421.050 ;
        RECT 481.950 419.400 526.050 420.600 ;
        RECT 481.950 418.950 484.050 419.400 ;
        RECT 487.950 418.950 490.050 419.400 ;
        RECT 523.950 418.950 526.050 419.400 ;
        RECT 610.950 420.600 613.050 421.050 ;
        RECT 634.950 420.600 637.050 421.050 ;
        RECT 610.950 419.400 637.050 420.600 ;
        RECT 610.950 418.950 613.050 419.400 ;
        RECT 634.950 418.950 637.050 419.400 ;
        RECT 703.950 420.600 706.050 421.050 ;
        RECT 727.950 420.600 730.050 421.050 ;
        RECT 703.950 419.400 730.050 420.600 ;
        RECT 703.950 418.950 706.050 419.400 ;
        RECT 727.950 418.950 730.050 419.400 ;
        RECT 427.950 417.600 430.050 418.050 ;
        RECT 404.400 416.400 430.050 417.600 ;
        RECT 376.950 415.950 379.050 416.400 ;
        RECT 385.950 415.950 388.050 416.400 ;
        RECT 427.950 415.950 430.050 416.400 ;
        RECT 439.950 417.600 442.050 418.050 ;
        RECT 448.950 417.600 451.050 418.050 ;
        RECT 439.950 416.400 451.050 417.600 ;
        RECT 439.950 415.950 442.050 416.400 ;
        RECT 448.950 415.950 451.050 416.400 ;
        RECT 454.950 417.600 457.050 418.050 ;
        RECT 466.950 417.600 469.050 418.050 ;
        RECT 526.950 417.600 529.050 418.050 ;
        RECT 454.950 416.400 469.050 417.600 ;
        RECT 454.950 415.950 457.050 416.400 ;
        RECT 466.950 415.950 469.050 416.400 ;
        RECT 497.400 416.400 529.050 417.600 ;
        RECT 421.950 414.600 424.050 415.050 ;
        RECT 430.950 414.600 433.050 415.050 ;
        RECT 362.400 413.400 366.600 414.600 ;
        RECT 319.950 411.600 322.050 412.050 ;
        RECT 302.400 410.400 322.050 411.600 ;
        RECT 319.950 409.950 322.050 410.400 ;
        RECT 340.950 409.950 343.050 412.050 ;
        RECT 343.950 411.600 346.050 412.050 ;
        RECT 349.950 411.600 352.050 412.050 ;
        RECT 343.950 410.400 352.050 411.600 ;
        RECT 365.400 411.600 366.600 413.400 ;
        RECT 421.950 413.400 433.050 414.600 ;
        RECT 421.950 412.950 424.050 413.400 ;
        RECT 430.950 412.950 433.050 413.400 ;
        RECT 445.950 414.600 448.050 415.050 ;
        RECT 497.400 414.600 498.600 416.400 ;
        RECT 526.950 415.950 529.050 416.400 ;
        RECT 538.950 417.600 541.050 418.050 ;
        RECT 559.950 417.600 562.050 418.050 ;
        RECT 538.950 416.400 562.050 417.600 ;
        RECT 538.950 415.950 541.050 416.400 ;
        RECT 559.950 415.950 562.050 416.400 ;
        RECT 634.950 417.600 637.050 418.050 ;
        RECT 706.950 417.600 709.050 418.050 ;
        RECT 634.950 416.400 709.050 417.600 ;
        RECT 634.950 415.950 637.050 416.400 ;
        RECT 706.950 415.950 709.050 416.400 ;
        RECT 712.950 417.600 715.050 418.050 ;
        RECT 715.950 417.600 718.050 418.050 ;
        RECT 754.950 417.600 757.050 418.050 ;
        RECT 772.950 417.600 775.050 418.050 ;
        RECT 712.950 416.400 775.050 417.600 ;
        RECT 712.950 415.950 715.050 416.400 ;
        RECT 715.950 415.950 718.050 416.400 ;
        RECT 754.950 415.950 757.050 416.400 ;
        RECT 772.950 415.950 775.050 416.400 ;
        RECT 445.950 413.400 498.600 414.600 ;
        RECT 499.950 414.600 502.050 415.050 ;
        RECT 508.950 414.600 511.050 415.050 ;
        RECT 517.950 414.600 520.050 415.050 ;
        RECT 499.950 413.400 504.600 414.600 ;
        RECT 445.950 412.950 448.050 413.400 ;
        RECT 499.950 412.950 502.050 413.400 ;
        RECT 503.400 412.050 504.600 413.400 ;
        RECT 508.950 413.400 520.050 414.600 ;
        RECT 508.950 412.950 511.050 413.400 ;
        RECT 517.950 412.950 520.050 413.400 ;
        RECT 529.950 414.600 532.050 415.050 ;
        RECT 535.950 414.600 538.050 415.050 ;
        RECT 529.950 413.400 538.050 414.600 ;
        RECT 529.950 412.950 532.050 413.400 ;
        RECT 535.950 412.950 538.050 413.400 ;
        RECT 556.950 412.950 559.050 415.050 ;
        RECT 625.950 412.950 628.050 415.050 ;
        RECT 703.950 414.600 706.050 415.050 ;
        RECT 742.950 414.600 745.050 415.050 ;
        RECT 703.950 413.400 745.050 414.600 ;
        RECT 703.950 412.950 706.050 413.400 ;
        RECT 742.950 412.950 745.050 413.400 ;
        RECT 766.950 414.600 769.050 415.050 ;
        RECT 775.950 414.600 778.050 415.050 ;
        RECT 766.950 413.400 778.050 414.600 ;
        RECT 766.950 412.950 769.050 413.400 ;
        RECT 775.950 412.950 778.050 413.400 ;
        RECT 382.950 411.600 385.050 412.050 ;
        RECT 365.400 410.400 385.050 411.600 ;
        RECT 343.950 409.950 346.050 410.400 ;
        RECT 349.950 409.950 352.050 410.400 ;
        RECT 382.950 409.950 385.050 410.400 ;
        RECT 436.950 411.600 439.050 412.050 ;
        RECT 451.950 411.600 454.050 412.050 ;
        RECT 436.950 410.400 454.050 411.600 ;
        RECT 436.950 409.950 439.050 410.400 ;
        RECT 451.950 409.950 454.050 410.400 ;
        RECT 463.950 411.600 466.050 412.050 ;
        RECT 475.950 411.600 478.050 412.050 ;
        RECT 463.950 410.400 478.050 411.600 ;
        RECT 463.950 409.950 466.050 410.400 ;
        RECT 475.950 409.950 478.050 410.400 ;
        RECT 484.950 411.600 487.050 412.050 ;
        RECT 502.950 411.600 505.050 412.050 ;
        RECT 484.950 410.400 505.050 411.600 ;
        RECT 484.950 409.950 487.050 410.400 ;
        RECT 502.950 409.950 505.050 410.400 ;
        RECT 220.950 407.400 261.600 408.600 ;
        RECT 262.950 408.600 265.050 409.050 ;
        RECT 286.950 408.600 289.050 409.050 ;
        RECT 262.950 407.400 289.050 408.600 ;
        RECT 220.950 406.950 223.050 407.400 ;
        RECT 262.950 406.950 265.050 407.400 ;
        RECT 286.950 406.950 289.050 407.400 ;
        RECT 307.950 408.600 310.050 409.050 ;
        RECT 322.950 408.600 325.050 409.050 ;
        RECT 307.950 407.400 325.050 408.600 ;
        RECT 307.950 406.950 310.050 407.400 ;
        RECT 322.950 406.950 325.050 407.400 ;
        RECT 340.950 408.600 343.050 409.050 ;
        RECT 385.950 408.600 388.050 409.050 ;
        RECT 340.950 407.400 388.050 408.600 ;
        RECT 340.950 406.950 343.050 407.400 ;
        RECT 385.950 406.950 388.050 407.400 ;
        RECT 415.950 408.600 418.050 409.050 ;
        RECT 424.950 408.600 427.050 409.050 ;
        RECT 415.950 407.400 427.050 408.600 ;
        RECT 415.950 406.950 418.050 407.400 ;
        RECT 424.950 406.950 427.050 407.400 ;
        RECT 472.950 408.600 475.050 409.050 ;
        RECT 490.950 408.600 493.050 409.050 ;
        RECT 472.950 407.400 493.050 408.600 ;
        RECT 472.950 406.950 475.050 407.400 ;
        RECT 490.950 406.950 493.050 407.400 ;
        RECT 529.950 408.600 532.050 409.050 ;
        RECT 547.950 408.600 550.050 409.050 ;
        RECT 529.950 407.400 550.050 408.600 ;
        RECT 529.950 406.950 532.050 407.400 ;
        RECT 547.950 406.950 550.050 407.400 ;
        RECT 557.400 406.050 558.600 412.950 ;
        RECT 616.950 411.600 619.050 412.050 ;
        RECT 626.400 411.600 627.600 412.950 ;
        RECT 616.950 410.400 627.600 411.600 ;
        RECT 709.950 411.600 712.050 412.050 ;
        RECT 721.950 411.600 724.050 412.050 ;
        RECT 709.950 410.400 724.050 411.600 ;
        RECT 616.950 409.950 619.050 410.400 ;
        RECT 709.950 409.950 712.050 410.400 ;
        RECT 721.950 409.950 724.050 410.400 ;
        RECT 724.950 411.600 727.050 412.050 ;
        RECT 733.950 411.600 736.050 412.050 ;
        RECT 724.950 410.400 736.050 411.600 ;
        RECT 724.950 409.950 727.050 410.400 ;
        RECT 733.950 409.950 736.050 410.400 ;
        RECT 736.950 411.600 739.050 412.050 ;
        RECT 751.950 411.600 754.050 412.050 ;
        RECT 736.950 410.400 754.050 411.600 ;
        RECT 736.950 409.950 739.050 410.400 ;
        RECT 751.950 409.950 754.050 410.400 ;
        RECT 763.950 411.600 766.050 412.050 ;
        RECT 784.950 411.600 787.050 412.050 ;
        RECT 763.950 410.400 787.050 411.600 ;
        RECT 763.950 409.950 766.050 410.400 ;
        RECT 784.950 409.950 787.050 410.400 ;
        RECT 787.950 411.600 790.050 412.050 ;
        RECT 793.950 411.600 796.050 412.050 ;
        RECT 787.950 410.400 796.050 411.600 ;
        RECT 787.950 409.950 790.050 410.400 ;
        RECT 793.950 409.950 796.050 410.400 ;
        RECT 841.950 411.600 844.050 412.050 ;
        RECT 853.950 411.600 856.050 412.050 ;
        RECT 841.950 410.400 856.050 411.600 ;
        RECT 841.950 409.950 844.050 410.400 ;
        RECT 853.950 409.950 856.050 410.400 ;
        RECT 634.950 408.600 637.050 409.050 ;
        RECT 649.950 408.600 652.050 409.050 ;
        RECT 634.950 407.400 652.050 408.600 ;
        RECT 634.950 406.950 637.050 407.400 ;
        RECT 649.950 406.950 652.050 407.400 ;
        RECT 748.950 408.600 751.050 409.050 ;
        RECT 775.950 408.600 778.050 409.050 ;
        RECT 748.950 407.400 778.050 408.600 ;
        RECT 748.950 406.950 751.050 407.400 ;
        RECT 775.950 406.950 778.050 407.400 ;
        RECT 835.950 408.600 838.050 409.050 ;
        RECT 847.950 408.600 850.050 409.050 ;
        RECT 835.950 407.400 850.050 408.600 ;
        RECT 835.950 406.950 838.050 407.400 ;
        RECT 847.950 406.950 850.050 407.400 ;
        RECT 34.950 405.600 37.050 406.050 ;
        RECT 154.950 405.600 157.050 406.050 ;
        RECT 34.950 404.400 157.050 405.600 ;
        RECT 34.950 403.950 37.050 404.400 ;
        RECT 154.950 403.950 157.050 404.400 ;
        RECT 262.950 405.600 265.050 406.050 ;
        RECT 271.950 405.600 274.050 406.050 ;
        RECT 262.950 404.400 274.050 405.600 ;
        RECT 262.950 403.950 265.050 404.400 ;
        RECT 271.950 403.950 274.050 404.400 ;
        RECT 274.950 405.600 277.050 406.050 ;
        RECT 298.950 405.600 301.050 406.050 ;
        RECT 319.950 405.600 322.050 406.050 ;
        RECT 274.950 404.400 322.050 405.600 ;
        RECT 274.950 403.950 277.050 404.400 ;
        RECT 298.950 403.950 301.050 404.400 ;
        RECT 319.950 403.950 322.050 404.400 ;
        RECT 328.950 405.600 331.050 406.050 ;
        RECT 367.950 405.600 370.050 406.050 ;
        RECT 328.950 404.400 370.050 405.600 ;
        RECT 328.950 403.950 331.050 404.400 ;
        RECT 367.950 403.950 370.050 404.400 ;
        RECT 391.950 405.600 394.050 406.050 ;
        RECT 403.950 405.600 406.050 406.050 ;
        RECT 484.950 405.600 487.050 406.050 ;
        RECT 499.950 405.600 502.050 406.050 ;
        RECT 511.950 405.600 514.050 406.050 ;
        RECT 391.950 404.400 514.050 405.600 ;
        RECT 391.950 403.950 394.050 404.400 ;
        RECT 403.950 403.950 406.050 404.400 ;
        RECT 484.950 403.950 487.050 404.400 ;
        RECT 499.950 403.950 502.050 404.400 ;
        RECT 511.950 403.950 514.050 404.400 ;
        RECT 556.950 403.950 559.050 406.050 ;
        RECT 694.950 405.600 697.050 406.050 ;
        RECT 820.950 405.600 823.050 406.050 ;
        RECT 694.950 404.400 823.050 405.600 ;
        RECT 694.950 403.950 697.050 404.400 ;
        RECT 820.950 403.950 823.050 404.400 ;
        RECT 61.950 402.600 64.050 403.050 ;
        RECT 121.950 402.600 124.050 403.050 ;
        RECT 130.950 402.600 133.050 403.050 ;
        RECT 187.950 402.600 190.050 403.050 ;
        RECT 244.950 402.600 247.050 403.050 ;
        RECT 61.950 401.400 133.050 402.600 ;
        RECT 61.950 400.950 64.050 401.400 ;
        RECT 121.950 400.950 124.050 401.400 ;
        RECT 130.950 400.950 133.050 401.400 ;
        RECT 134.400 401.400 247.050 402.600 ;
        RECT 109.950 399.600 112.050 400.050 ;
        RECT 134.400 399.600 135.600 401.400 ;
        RECT 187.950 400.950 190.050 401.400 ;
        RECT 244.950 400.950 247.050 401.400 ;
        RECT 259.950 402.600 262.050 403.050 ;
        RECT 265.950 402.600 268.050 403.050 ;
        RECT 259.950 401.400 268.050 402.600 ;
        RECT 259.950 400.950 262.050 401.400 ;
        RECT 265.950 400.950 268.050 401.400 ;
        RECT 487.950 402.600 490.050 403.050 ;
        RECT 493.950 402.600 496.050 403.050 ;
        RECT 487.950 401.400 496.050 402.600 ;
        RECT 487.950 400.950 490.050 401.400 ;
        RECT 493.950 400.950 496.050 401.400 ;
        RECT 523.950 402.600 526.050 403.050 ;
        RECT 571.950 402.600 574.050 403.050 ;
        RECT 523.950 401.400 574.050 402.600 ;
        RECT 523.950 400.950 526.050 401.400 ;
        RECT 571.950 400.950 574.050 401.400 ;
        RECT 631.950 402.600 634.050 403.050 ;
        RECT 676.950 402.600 679.050 403.050 ;
        RECT 631.950 401.400 679.050 402.600 ;
        RECT 631.950 400.950 634.050 401.400 ;
        RECT 676.950 400.950 679.050 401.400 ;
        RECT 109.950 398.400 135.600 399.600 ;
        RECT 142.950 399.600 145.050 400.050 ;
        RECT 175.950 399.600 178.050 400.050 ;
        RECT 142.950 398.400 178.050 399.600 ;
        RECT 109.950 397.950 112.050 398.400 ;
        RECT 142.950 397.950 145.050 398.400 ;
        RECT 175.950 397.950 178.050 398.400 ;
        RECT 199.950 399.600 202.050 400.050 ;
        RECT 205.950 399.600 208.050 400.050 ;
        RECT 199.950 398.400 208.050 399.600 ;
        RECT 199.950 397.950 202.050 398.400 ;
        RECT 205.950 397.950 208.050 398.400 ;
        RECT 214.950 399.600 217.050 400.050 ;
        RECT 274.950 399.600 277.050 400.050 ;
        RECT 214.950 398.400 277.050 399.600 ;
        RECT 214.950 397.950 217.050 398.400 ;
        RECT 274.950 397.950 277.050 398.400 ;
        RECT 283.950 399.600 286.050 400.050 ;
        RECT 295.950 399.600 298.050 400.050 ;
        RECT 352.950 399.600 355.050 400.050 ;
        RECT 283.950 398.400 355.050 399.600 ;
        RECT 283.950 397.950 286.050 398.400 ;
        RECT 295.950 397.950 298.050 398.400 ;
        RECT 352.950 397.950 355.050 398.400 ;
        RECT 370.950 399.600 373.050 400.050 ;
        RECT 535.950 399.600 538.050 400.050 ;
        RECT 370.950 398.400 538.050 399.600 ;
        RECT 370.950 397.950 373.050 398.400 ;
        RECT 535.950 397.950 538.050 398.400 ;
        RECT 568.950 399.600 571.050 400.050 ;
        RECT 607.950 399.600 610.050 400.050 ;
        RECT 619.950 399.600 622.050 400.050 ;
        RECT 568.950 398.400 622.050 399.600 ;
        RECT 568.950 397.950 571.050 398.400 ;
        RECT 607.950 397.950 610.050 398.400 ;
        RECT 619.950 397.950 622.050 398.400 ;
        RECT 643.950 399.600 646.050 400.050 ;
        RECT 661.950 399.600 664.050 400.050 ;
        RECT 643.950 398.400 664.050 399.600 ;
        RECT 643.950 397.950 646.050 398.400 ;
        RECT 661.950 397.950 664.050 398.400 ;
        RECT 664.950 399.600 667.050 400.050 ;
        RECT 718.950 399.600 721.050 400.050 ;
        RECT 664.950 398.400 721.050 399.600 ;
        RECT 664.950 397.950 667.050 398.400 ;
        RECT 718.950 397.950 721.050 398.400 ;
        RECT 76.950 396.600 79.050 397.050 ;
        RECT 103.950 396.600 106.050 397.050 ;
        RECT 76.950 395.400 106.050 396.600 ;
        RECT 76.950 394.950 79.050 395.400 ;
        RECT 103.950 394.950 106.050 395.400 ;
        RECT 112.950 396.600 115.050 397.050 ;
        RECT 265.950 396.600 268.050 397.050 ;
        RECT 112.950 395.400 268.050 396.600 ;
        RECT 112.950 394.950 115.050 395.400 ;
        RECT 265.950 394.950 268.050 395.400 ;
        RECT 304.950 396.600 307.050 397.050 ;
        RECT 388.950 396.600 391.050 397.050 ;
        RECT 445.950 396.600 448.050 397.050 ;
        RECT 304.950 395.400 448.050 396.600 ;
        RECT 304.950 394.950 307.050 395.400 ;
        RECT 388.950 394.950 391.050 395.400 ;
        RECT 445.950 394.950 448.050 395.400 ;
        RECT 481.950 396.600 484.050 397.050 ;
        RECT 490.950 396.600 493.050 397.050 ;
        RECT 481.950 395.400 493.050 396.600 ;
        RECT 481.950 394.950 484.050 395.400 ;
        RECT 490.950 394.950 493.050 395.400 ;
        RECT 628.950 396.600 631.050 397.050 ;
        RECT 670.950 396.600 673.050 397.050 ;
        RECT 628.950 395.400 673.050 396.600 ;
        RECT 628.950 394.950 631.050 395.400 ;
        RECT 670.950 394.950 673.050 395.400 ;
        RECT 700.950 396.600 703.050 397.050 ;
        RECT 715.950 396.600 718.050 397.050 ;
        RECT 700.950 395.400 718.050 396.600 ;
        RECT 700.950 394.950 703.050 395.400 ;
        RECT 715.950 394.950 718.050 395.400 ;
        RECT 10.950 393.600 13.050 394.050 ;
        RECT 37.950 393.600 40.050 394.050 ;
        RECT 10.950 392.400 40.050 393.600 ;
        RECT 10.950 391.950 13.050 392.400 ;
        RECT 37.950 391.950 40.050 392.400 ;
        RECT 97.950 393.600 100.050 394.050 ;
        RECT 112.950 393.600 115.050 394.050 ;
        RECT 97.950 392.400 115.050 393.600 ;
        RECT 97.950 391.950 100.050 392.400 ;
        RECT 112.950 391.950 115.050 392.400 ;
        RECT 163.950 393.600 166.050 394.050 ;
        RECT 166.950 393.600 169.050 394.050 ;
        RECT 184.950 393.600 187.050 394.050 ;
        RECT 163.950 392.400 187.050 393.600 ;
        RECT 163.950 391.950 166.050 392.400 ;
        RECT 166.950 391.950 169.050 392.400 ;
        RECT 184.950 391.950 187.050 392.400 ;
        RECT 196.950 393.600 199.050 394.050 ;
        RECT 250.950 393.600 253.050 394.050 ;
        RECT 196.950 392.400 253.050 393.600 ;
        RECT 196.950 391.950 199.050 392.400 ;
        RECT 250.950 391.950 253.050 392.400 ;
        RECT 280.950 393.600 283.050 394.050 ;
        RECT 301.950 393.600 304.050 394.050 ;
        RECT 280.950 392.400 304.050 393.600 ;
        RECT 280.950 391.950 283.050 392.400 ;
        RECT 301.950 391.950 304.050 392.400 ;
        RECT 325.950 393.600 328.050 394.050 ;
        RECT 409.950 393.600 412.050 394.050 ;
        RECT 325.950 392.400 412.050 393.600 ;
        RECT 325.950 391.950 328.050 392.400 ;
        RECT 409.950 391.950 412.050 392.400 ;
        RECT 415.950 393.600 418.050 394.050 ;
        RECT 562.950 393.600 565.050 394.050 ;
        RECT 415.950 392.400 565.050 393.600 ;
        RECT 415.950 391.950 418.050 392.400 ;
        RECT 562.950 391.950 565.050 392.400 ;
        RECT 637.950 393.600 640.050 394.050 ;
        RECT 682.950 393.600 685.050 394.050 ;
        RECT 715.950 393.600 718.050 394.050 ;
        RECT 637.950 392.400 718.050 393.600 ;
        RECT 637.950 391.950 640.050 392.400 ;
        RECT 682.950 391.950 685.050 392.400 ;
        RECT 715.950 391.950 718.050 392.400 ;
        RECT 730.950 393.600 733.050 394.050 ;
        RECT 808.950 393.600 811.050 394.050 ;
        RECT 730.950 392.400 811.050 393.600 ;
        RECT 730.950 391.950 733.050 392.400 ;
        RECT 808.950 391.950 811.050 392.400 ;
        RECT 16.950 390.600 19.050 391.050 ;
        RECT 19.950 390.600 22.050 391.050 ;
        RECT 193.950 390.600 196.050 391.050 ;
        RECT 16.950 389.400 196.050 390.600 ;
        RECT 16.950 388.950 19.050 389.400 ;
        RECT 19.950 388.950 22.050 389.400 ;
        RECT 193.950 388.950 196.050 389.400 ;
        RECT 196.950 390.600 199.050 391.050 ;
        RECT 202.950 390.600 205.050 391.050 ;
        RECT 196.950 389.400 205.050 390.600 ;
        RECT 196.950 388.950 199.050 389.400 ;
        RECT 202.950 388.950 205.050 389.400 ;
        RECT 226.950 390.600 229.050 391.050 ;
        RECT 232.950 390.600 235.050 391.050 ;
        RECT 226.950 389.400 235.050 390.600 ;
        RECT 226.950 388.950 229.050 389.400 ;
        RECT 232.950 388.950 235.050 389.400 ;
        RECT 238.950 390.600 241.050 391.050 ;
        RECT 316.950 390.600 319.050 391.050 ;
        RECT 337.950 390.600 340.050 391.050 ;
        RECT 238.950 389.400 315.600 390.600 ;
        RECT 238.950 388.950 241.050 389.400 ;
        RECT 10.950 387.600 13.050 388.050 ;
        RECT 19.950 387.600 22.050 388.050 ;
        RECT 10.950 386.400 22.050 387.600 ;
        RECT 10.950 385.950 13.050 386.400 ;
        RECT 19.950 385.950 22.050 386.400 ;
        RECT 82.950 387.600 85.050 388.050 ;
        RECT 97.950 387.600 100.050 388.050 ;
        RECT 109.950 387.600 112.050 388.050 ;
        RECT 127.950 387.600 130.050 388.050 ;
        RECT 82.950 386.400 96.600 387.600 ;
        RECT 82.950 385.950 85.050 386.400 ;
        RECT 43.950 384.600 46.050 385.050 ;
        RECT 52.950 384.600 55.050 385.050 ;
        RECT 43.950 383.400 55.050 384.600 ;
        RECT 43.950 382.950 46.050 383.400 ;
        RECT 52.950 382.950 55.050 383.400 ;
        RECT 58.950 384.600 61.050 385.050 ;
        RECT 64.950 384.600 67.050 385.050 ;
        RECT 58.950 383.400 67.050 384.600 ;
        RECT 58.950 382.950 61.050 383.400 ;
        RECT 64.950 382.950 67.050 383.400 ;
        RECT 76.950 384.600 79.050 385.050 ;
        RECT 88.950 384.600 91.050 385.050 ;
        RECT 76.950 383.400 91.050 384.600 ;
        RECT 76.950 382.950 79.050 383.400 ;
        RECT 88.950 382.950 91.050 383.400 ;
        RECT 91.950 382.950 94.050 385.050 ;
        RECT 95.400 384.600 96.600 386.400 ;
        RECT 97.950 386.400 130.050 387.600 ;
        RECT 97.950 385.950 100.050 386.400 ;
        RECT 109.950 385.950 112.050 386.400 ;
        RECT 127.950 385.950 130.050 386.400 ;
        RECT 193.950 387.600 196.050 388.050 ;
        RECT 268.950 387.600 271.050 388.050 ;
        RECT 310.950 387.600 313.050 388.050 ;
        RECT 193.950 386.400 313.050 387.600 ;
        RECT 314.400 387.600 315.600 389.400 ;
        RECT 316.950 389.400 340.050 390.600 ;
        RECT 316.950 388.950 319.050 389.400 ;
        RECT 337.950 388.950 340.050 389.400 ;
        RECT 373.950 390.600 376.050 391.050 ;
        RECT 391.950 390.600 394.050 391.050 ;
        RECT 397.950 390.600 400.050 391.050 ;
        RECT 373.950 389.400 400.050 390.600 ;
        RECT 373.950 388.950 376.050 389.400 ;
        RECT 391.950 388.950 394.050 389.400 ;
        RECT 397.950 388.950 400.050 389.400 ;
        RECT 442.950 390.600 445.050 391.050 ;
        RECT 469.950 390.600 472.050 391.050 ;
        RECT 442.950 389.400 472.050 390.600 ;
        RECT 442.950 388.950 445.050 389.400 ;
        RECT 469.950 388.950 472.050 389.400 ;
        RECT 481.950 390.600 484.050 391.050 ;
        RECT 493.950 390.600 496.050 391.050 ;
        RECT 481.950 389.400 496.050 390.600 ;
        RECT 481.950 388.950 484.050 389.400 ;
        RECT 493.950 388.950 496.050 389.400 ;
        RECT 628.950 390.600 631.050 391.050 ;
        RECT 640.950 390.600 643.050 391.050 ;
        RECT 628.950 389.400 643.050 390.600 ;
        RECT 628.950 388.950 631.050 389.400 ;
        RECT 640.950 388.950 643.050 389.400 ;
        RECT 646.950 390.600 649.050 391.050 ;
        RECT 757.950 390.600 760.050 391.050 ;
        RECT 820.950 390.600 823.050 391.050 ;
        RECT 856.950 390.600 859.050 391.050 ;
        RECT 646.950 389.400 735.600 390.600 ;
        RECT 646.950 388.950 649.050 389.400 ;
        RECT 376.950 387.600 379.050 388.050 ;
        RECT 314.400 386.400 379.050 387.600 ;
        RECT 193.950 385.950 196.050 386.400 ;
        RECT 268.950 385.950 271.050 386.400 ;
        RECT 310.950 385.950 313.050 386.400 ;
        RECT 376.950 385.950 379.050 386.400 ;
        RECT 397.950 387.600 400.050 388.050 ;
        RECT 475.950 387.600 478.050 388.050 ;
        RECT 610.950 387.600 613.050 388.050 ;
        RECT 397.950 386.400 613.050 387.600 ;
        RECT 397.950 385.950 400.050 386.400 ;
        RECT 475.950 385.950 478.050 386.400 ;
        RECT 610.950 385.950 613.050 386.400 ;
        RECT 625.950 387.600 628.050 388.050 ;
        RECT 640.950 387.600 643.050 388.050 ;
        RECT 655.950 387.600 658.050 388.050 ;
        RECT 625.950 386.400 658.050 387.600 ;
        RECT 625.950 385.950 628.050 386.400 ;
        RECT 640.950 385.950 643.050 386.400 ;
        RECT 655.950 385.950 658.050 386.400 ;
        RECT 730.950 385.950 733.050 388.050 ;
        RECT 734.400 387.600 735.600 389.400 ;
        RECT 757.950 389.400 859.050 390.600 ;
        RECT 757.950 388.950 760.050 389.400 ;
        RECT 820.950 388.950 823.050 389.400 ;
        RECT 856.950 388.950 859.050 389.400 ;
        RECT 790.950 387.600 793.050 388.050 ;
        RECT 734.400 386.400 793.050 387.600 ;
        RECT 106.950 384.600 109.050 385.050 ;
        RECT 115.950 384.600 118.050 385.050 ;
        RECT 95.400 383.400 118.050 384.600 ;
        RECT 106.950 382.950 109.050 383.400 ;
        RECT 115.950 382.950 118.050 383.400 ;
        RECT 124.950 384.600 127.050 385.050 ;
        RECT 157.950 384.600 160.050 385.050 ;
        RECT 124.950 383.400 160.050 384.600 ;
        RECT 124.950 382.950 127.050 383.400 ;
        RECT 157.950 382.950 160.050 383.400 ;
        RECT 211.950 384.600 214.050 385.050 ;
        RECT 256.950 384.600 259.050 385.050 ;
        RECT 274.950 384.600 277.050 385.050 ;
        RECT 295.950 384.600 298.050 385.050 ;
        RECT 211.950 383.400 231.600 384.600 ;
        RECT 211.950 382.950 214.050 383.400 ;
        RECT 64.950 381.600 67.050 382.050 ;
        RECT 92.400 381.600 93.600 382.950 ;
        RECT 230.400 382.050 231.600 383.400 ;
        RECT 256.950 383.400 277.050 384.600 ;
        RECT 256.950 382.950 259.050 383.400 ;
        RECT 274.950 382.950 277.050 383.400 ;
        RECT 278.400 383.400 298.050 384.600 ;
        RECT 35.400 380.400 93.600 381.600 ;
        RECT 118.950 381.600 121.050 382.050 ;
        RECT 163.950 381.600 166.050 382.050 ;
        RECT 220.950 381.600 223.050 382.050 ;
        RECT 118.950 380.400 166.050 381.600 ;
        RECT 35.400 379.050 36.600 380.400 ;
        RECT 64.950 379.950 67.050 380.400 ;
        RECT 118.950 379.950 121.050 380.400 ;
        RECT 163.950 379.950 166.050 380.400 ;
        RECT 209.400 380.400 223.050 381.600 ;
        RECT 209.400 379.050 210.600 380.400 ;
        RECT 220.950 379.950 223.050 380.400 ;
        RECT 229.950 379.950 232.050 382.050 ;
        RECT 235.950 381.600 238.050 382.050 ;
        RECT 278.400 381.600 279.600 383.400 ;
        RECT 295.950 382.950 298.050 383.400 ;
        RECT 301.950 384.600 304.050 385.050 ;
        RECT 325.950 384.600 328.050 385.050 ;
        RECT 301.950 383.400 328.050 384.600 ;
        RECT 301.950 382.950 304.050 383.400 ;
        RECT 325.950 382.950 328.050 383.400 ;
        RECT 358.950 384.600 361.050 385.050 ;
        RECT 367.950 384.600 370.050 385.050 ;
        RECT 358.950 383.400 370.050 384.600 ;
        RECT 358.950 382.950 361.050 383.400 ;
        RECT 367.950 382.950 370.050 383.400 ;
        RECT 394.950 382.950 397.050 385.050 ;
        RECT 418.950 384.600 421.050 385.050 ;
        RECT 457.950 384.600 460.050 385.050 ;
        RECT 418.950 383.400 460.050 384.600 ;
        RECT 418.950 382.950 421.050 383.400 ;
        RECT 457.950 382.950 460.050 383.400 ;
        RECT 460.950 384.600 463.050 385.050 ;
        RECT 469.950 384.600 472.050 385.050 ;
        RECT 460.950 383.400 472.050 384.600 ;
        RECT 460.950 382.950 463.050 383.400 ;
        RECT 469.950 382.950 472.050 383.400 ;
        RECT 478.950 384.600 481.050 385.050 ;
        RECT 496.950 384.600 499.050 385.050 ;
        RECT 478.950 383.400 499.050 384.600 ;
        RECT 478.950 382.950 481.050 383.400 ;
        RECT 496.950 382.950 499.050 383.400 ;
        RECT 499.950 384.600 502.050 385.050 ;
        RECT 520.950 384.600 523.050 385.050 ;
        RECT 499.950 383.400 523.050 384.600 ;
        RECT 499.950 382.950 502.050 383.400 ;
        RECT 520.950 382.950 523.050 383.400 ;
        RECT 523.950 384.600 526.050 385.050 ;
        RECT 541.950 384.600 544.050 385.050 ;
        RECT 523.950 383.400 544.050 384.600 ;
        RECT 523.950 382.950 526.050 383.400 ;
        RECT 541.950 382.950 544.050 383.400 ;
        RECT 646.950 384.600 649.050 385.050 ;
        RECT 652.950 384.600 655.050 385.050 ;
        RECT 646.950 383.400 655.050 384.600 ;
        RECT 646.950 382.950 649.050 383.400 ;
        RECT 652.950 382.950 655.050 383.400 ;
        RECT 658.950 384.600 661.050 385.050 ;
        RECT 664.950 384.600 667.050 385.050 ;
        RECT 658.950 383.400 667.050 384.600 ;
        RECT 731.400 384.600 732.600 385.950 ;
        RECT 758.400 385.050 759.600 386.400 ;
        RECT 790.950 385.950 793.050 386.400 ;
        RECT 814.950 387.600 817.050 388.050 ;
        RECT 844.950 387.600 847.050 388.050 ;
        RECT 814.950 386.400 847.050 387.600 ;
        RECT 814.950 385.950 817.050 386.400 ;
        RECT 844.950 385.950 847.050 386.400 ;
        RECT 754.950 384.600 757.050 385.050 ;
        RECT 731.400 383.400 757.050 384.600 ;
        RECT 658.950 382.950 661.050 383.400 ;
        RECT 664.950 382.950 667.050 383.400 ;
        RECT 754.950 382.950 757.050 383.400 ;
        RECT 757.950 382.950 760.050 385.050 ;
        RECT 760.950 384.600 763.050 385.050 ;
        RECT 787.950 384.600 790.050 385.050 ;
        RECT 760.950 383.400 790.050 384.600 ;
        RECT 760.950 382.950 763.050 383.400 ;
        RECT 787.950 382.950 790.050 383.400 ;
        RECT 802.950 384.600 805.050 385.050 ;
        RECT 802.950 383.400 834.600 384.600 ;
        RECT 802.950 382.950 805.050 383.400 ;
        RECT 235.950 380.400 279.600 381.600 ;
        RECT 313.950 381.600 316.050 382.050 ;
        RECT 328.950 381.600 331.050 382.050 ;
        RECT 313.950 380.400 331.050 381.600 ;
        RECT 235.950 379.950 238.050 380.400 ;
        RECT 313.950 379.950 316.050 380.400 ;
        RECT 328.950 379.950 331.050 380.400 ;
        RECT 361.950 381.600 364.050 382.050 ;
        RECT 373.950 381.600 376.050 382.050 ;
        RECT 361.950 380.400 376.050 381.600 ;
        RECT 361.950 379.950 364.050 380.400 ;
        RECT 373.950 379.950 376.050 380.400 ;
        RECT 376.950 381.600 379.050 382.050 ;
        RECT 382.950 381.600 385.050 382.050 ;
        RECT 395.400 381.600 396.600 382.950 ;
        RECT 529.950 381.600 532.050 382.050 ;
        RECT 376.950 380.400 385.050 381.600 ;
        RECT 376.950 379.950 379.050 380.400 ;
        RECT 382.950 379.950 385.050 380.400 ;
        RECT 392.400 380.400 532.050 381.600 ;
        RECT 34.950 376.950 37.050 379.050 ;
        RECT 70.950 378.600 73.050 379.050 ;
        RECT 190.950 378.600 193.050 379.050 ;
        RECT 202.950 378.600 205.050 379.050 ;
        RECT 70.950 377.400 205.050 378.600 ;
        RECT 70.950 376.950 73.050 377.400 ;
        RECT 190.950 376.950 193.050 377.400 ;
        RECT 202.950 376.950 205.050 377.400 ;
        RECT 208.950 376.950 211.050 379.050 ;
        RECT 238.950 378.600 241.050 379.050 ;
        RECT 253.950 378.600 256.050 379.050 ;
        RECT 238.950 377.400 256.050 378.600 ;
        RECT 238.950 376.950 241.050 377.400 ;
        RECT 253.950 376.950 256.050 377.400 ;
        RECT 322.950 378.600 325.050 379.050 ;
        RECT 392.400 378.600 393.600 380.400 ;
        RECT 529.950 379.950 532.050 380.400 ;
        RECT 535.950 381.600 538.050 382.050 ;
        RECT 541.950 381.600 544.050 382.050 ;
        RECT 535.950 380.400 544.050 381.600 ;
        RECT 535.950 379.950 538.050 380.400 ;
        RECT 541.950 379.950 544.050 380.400 ;
        RECT 637.950 381.600 640.050 382.050 ;
        RECT 673.950 381.600 676.050 382.050 ;
        RECT 637.950 380.400 676.050 381.600 ;
        RECT 637.950 379.950 640.050 380.400 ;
        RECT 673.950 379.950 676.050 380.400 ;
        RECT 754.950 381.600 757.050 382.050 ;
        RECT 784.950 381.600 787.050 382.050 ;
        RECT 808.950 381.600 811.050 382.050 ;
        RECT 829.950 381.600 832.050 382.050 ;
        RECT 754.950 380.400 811.050 381.600 ;
        RECT 754.950 379.950 757.050 380.400 ;
        RECT 784.950 379.950 787.050 380.400 ;
        RECT 808.950 379.950 811.050 380.400 ;
        RECT 812.400 380.400 832.050 381.600 ;
        RECT 833.400 381.600 834.600 383.400 ;
        RECT 853.950 382.950 856.050 385.050 ;
        RECT 847.950 381.600 850.050 382.050 ;
        RECT 833.400 380.400 850.050 381.600 ;
        RECT 854.400 381.600 855.600 382.950 ;
        RECT 856.950 381.600 859.050 382.050 ;
        RECT 854.400 380.400 859.050 381.600 ;
        RECT 812.400 379.050 813.600 380.400 ;
        RECT 829.950 379.950 832.050 380.400 ;
        RECT 847.950 379.950 850.050 380.400 ;
        RECT 856.950 379.950 859.050 380.400 ;
        RECT 322.950 377.400 393.600 378.600 ;
        RECT 394.950 378.600 397.050 379.050 ;
        RECT 463.950 378.600 466.050 379.050 ;
        RECT 394.950 377.400 466.050 378.600 ;
        RECT 322.950 376.950 325.050 377.400 ;
        RECT 394.950 376.950 397.050 377.400 ;
        RECT 463.950 376.950 466.050 377.400 ;
        RECT 475.950 378.600 478.050 379.050 ;
        RECT 481.950 378.600 484.050 379.050 ;
        RECT 475.950 377.400 484.050 378.600 ;
        RECT 475.950 376.950 478.050 377.400 ;
        RECT 481.950 376.950 484.050 377.400 ;
        RECT 526.950 378.600 529.050 379.050 ;
        RECT 532.950 378.600 535.050 379.050 ;
        RECT 526.950 377.400 535.050 378.600 ;
        RECT 526.950 376.950 529.050 377.400 ;
        RECT 532.950 376.950 535.050 377.400 ;
        RECT 538.950 378.600 541.050 379.050 ;
        RECT 556.950 378.600 559.050 379.050 ;
        RECT 538.950 377.400 559.050 378.600 ;
        RECT 538.950 376.950 541.050 377.400 ;
        RECT 556.950 376.950 559.050 377.400 ;
        RECT 610.950 378.600 613.050 379.050 ;
        RECT 679.950 378.600 682.050 379.050 ;
        RECT 706.950 378.600 709.050 379.050 ;
        RECT 610.950 377.400 709.050 378.600 ;
        RECT 610.950 376.950 613.050 377.400 ;
        RECT 679.950 376.950 682.050 377.400 ;
        RECT 706.950 376.950 709.050 377.400 ;
        RECT 727.950 378.600 730.050 379.050 ;
        RECT 769.950 378.600 772.050 379.050 ;
        RECT 787.950 378.600 790.050 379.050 ;
        RECT 793.950 378.600 796.050 379.050 ;
        RECT 727.950 377.400 796.050 378.600 ;
        RECT 727.950 376.950 730.050 377.400 ;
        RECT 769.950 376.950 772.050 377.400 ;
        RECT 787.950 376.950 790.050 377.400 ;
        RECT 793.950 376.950 796.050 377.400 ;
        RECT 805.950 378.600 808.050 379.050 ;
        RECT 811.950 378.600 814.050 379.050 ;
        RECT 805.950 377.400 814.050 378.600 ;
        RECT 805.950 376.950 808.050 377.400 ;
        RECT 811.950 376.950 814.050 377.400 ;
        RECT 820.950 378.600 823.050 379.050 ;
        RECT 832.950 378.600 835.050 379.050 ;
        RECT 820.950 377.400 835.050 378.600 ;
        RECT 820.950 376.950 823.050 377.400 ;
        RECT 832.950 376.950 835.050 377.400 ;
        RECT 841.950 378.600 844.050 379.050 ;
        RECT 853.950 378.600 856.050 379.050 ;
        RECT 841.950 377.400 856.050 378.600 ;
        RECT 841.950 376.950 844.050 377.400 ;
        RECT 853.950 376.950 856.050 377.400 ;
        RECT 13.950 375.600 16.050 376.050 ;
        RECT 64.950 375.600 67.050 376.050 ;
        RECT 85.950 375.600 88.050 376.050 ;
        RECT 13.950 374.400 88.050 375.600 ;
        RECT 13.950 373.950 16.050 374.400 ;
        RECT 64.950 373.950 67.050 374.400 ;
        RECT 85.950 373.950 88.050 374.400 ;
        RECT 94.950 375.600 97.050 376.050 ;
        RECT 154.950 375.600 157.050 376.050 ;
        RECT 184.950 375.600 187.050 376.050 ;
        RECT 457.950 375.600 460.050 376.050 ;
        RECT 751.950 375.600 754.050 376.050 ;
        RECT 94.950 374.400 754.050 375.600 ;
        RECT 94.950 373.950 97.050 374.400 ;
        RECT 154.950 373.950 157.050 374.400 ;
        RECT 184.950 373.950 187.050 374.400 ;
        RECT 457.950 373.950 460.050 374.400 ;
        RECT 751.950 373.950 754.050 374.400 ;
        RECT 835.950 375.600 838.050 376.050 ;
        RECT 847.950 375.600 850.050 376.050 ;
        RECT 835.950 374.400 850.050 375.600 ;
        RECT 835.950 373.950 838.050 374.400 ;
        RECT 847.950 373.950 850.050 374.400 ;
        RECT 67.950 372.600 70.050 373.050 ;
        RECT 118.950 372.600 121.050 373.050 ;
        RECT 67.950 371.400 121.050 372.600 ;
        RECT 67.950 370.950 70.050 371.400 ;
        RECT 118.950 370.950 121.050 371.400 ;
        RECT 121.950 372.600 124.050 373.050 ;
        RECT 139.950 372.600 142.050 373.050 ;
        RECT 121.950 371.400 142.050 372.600 ;
        RECT 121.950 370.950 124.050 371.400 ;
        RECT 139.950 370.950 142.050 371.400 ;
        RECT 151.950 372.600 154.050 373.050 ;
        RECT 172.950 372.600 175.050 373.050 ;
        RECT 151.950 371.400 175.050 372.600 ;
        RECT 151.950 370.950 154.050 371.400 ;
        RECT 172.950 370.950 175.050 371.400 ;
        RECT 175.950 372.600 178.050 373.050 ;
        RECT 187.950 372.600 190.050 373.050 ;
        RECT 175.950 371.400 190.050 372.600 ;
        RECT 175.950 370.950 178.050 371.400 ;
        RECT 187.950 370.950 190.050 371.400 ;
        RECT 298.950 372.600 301.050 373.050 ;
        RECT 391.950 372.600 394.050 373.050 ;
        RECT 298.950 371.400 394.050 372.600 ;
        RECT 298.950 370.950 301.050 371.400 ;
        RECT 391.950 370.950 394.050 371.400 ;
        RECT 403.950 372.600 406.050 373.050 ;
        RECT 412.950 372.600 415.050 373.050 ;
        RECT 475.950 372.600 478.050 373.050 ;
        RECT 487.950 372.600 490.050 373.050 ;
        RECT 403.950 371.400 490.050 372.600 ;
        RECT 403.950 370.950 406.050 371.400 ;
        RECT 412.950 370.950 415.050 371.400 ;
        RECT 475.950 370.950 478.050 371.400 ;
        RECT 487.950 370.950 490.050 371.400 ;
        RECT 565.950 370.950 568.050 373.050 ;
        RECT 649.950 372.600 652.050 373.050 ;
        RECT 661.950 372.600 664.050 373.050 ;
        RECT 649.950 371.400 664.050 372.600 ;
        RECT 649.950 370.950 652.050 371.400 ;
        RECT 661.950 370.950 664.050 371.400 ;
        RECT 673.950 372.600 676.050 373.050 ;
        RECT 700.950 372.600 703.050 373.050 ;
        RECT 673.950 371.400 703.050 372.600 ;
        RECT 673.950 370.950 676.050 371.400 ;
        RECT 700.950 370.950 703.050 371.400 ;
        RECT 769.950 372.600 772.050 373.050 ;
        RECT 778.950 372.600 781.050 373.050 ;
        RECT 769.950 371.400 781.050 372.600 ;
        RECT 769.950 370.950 772.050 371.400 ;
        RECT 778.950 370.950 781.050 371.400 ;
        RECT 826.950 372.600 829.050 373.050 ;
        RECT 856.950 372.600 859.050 373.050 ;
        RECT 826.950 371.400 859.050 372.600 ;
        RECT 826.950 370.950 829.050 371.400 ;
        RECT 856.950 370.950 859.050 371.400 ;
        RECT 61.950 369.600 64.050 370.050 ;
        RECT 142.950 369.600 145.050 370.050 ;
        RECT 163.950 369.600 166.050 370.050 ;
        RECT 61.950 368.400 135.600 369.600 ;
        RECT 61.950 367.950 64.050 368.400 ;
        RECT 134.400 366.600 135.600 368.400 ;
        RECT 142.950 368.400 166.050 369.600 ;
        RECT 142.950 367.950 145.050 368.400 ;
        RECT 163.950 367.950 166.050 368.400 ;
        RECT 244.950 369.600 247.050 370.050 ;
        RECT 259.950 369.600 262.050 370.050 ;
        RECT 244.950 368.400 262.050 369.600 ;
        RECT 244.950 367.950 247.050 368.400 ;
        RECT 259.950 367.950 262.050 368.400 ;
        RECT 325.950 369.600 328.050 370.050 ;
        RECT 553.950 369.600 556.050 370.050 ;
        RECT 325.950 368.400 556.050 369.600 ;
        RECT 325.950 367.950 328.050 368.400 ;
        RECT 553.950 367.950 556.050 368.400 ;
        RECT 556.950 369.600 559.050 370.050 ;
        RECT 566.400 369.600 567.600 370.950 ;
        RECT 556.950 368.400 567.600 369.600 ;
        RECT 673.950 369.600 676.050 370.050 ;
        RECT 685.950 369.600 688.050 370.050 ;
        RECT 673.950 368.400 688.050 369.600 ;
        RECT 556.950 367.950 559.050 368.400 ;
        RECT 673.950 367.950 676.050 368.400 ;
        RECT 685.950 367.950 688.050 368.400 ;
        RECT 838.950 369.600 841.050 370.050 ;
        RECT 856.950 369.600 859.050 370.050 ;
        RECT 838.950 368.400 859.050 369.600 ;
        RECT 838.950 367.950 841.050 368.400 ;
        RECT 856.950 367.950 859.050 368.400 ;
        RECT 325.950 366.600 328.050 367.050 ;
        RECT 134.400 365.400 328.050 366.600 ;
        RECT 325.950 364.950 328.050 365.400 ;
        RECT 373.950 366.600 376.050 367.050 ;
        RECT 379.950 366.600 382.050 367.050 ;
        RECT 373.950 365.400 382.050 366.600 ;
        RECT 373.950 364.950 376.050 365.400 ;
        RECT 379.950 364.950 382.050 365.400 ;
        RECT 382.950 366.600 385.050 367.050 ;
        RECT 406.950 366.600 409.050 367.050 ;
        RECT 382.950 365.400 409.050 366.600 ;
        RECT 382.950 364.950 385.050 365.400 ;
        RECT 406.950 364.950 409.050 365.400 ;
        RECT 463.950 366.600 466.050 367.050 ;
        RECT 589.950 366.600 592.050 367.050 ;
        RECT 595.950 366.600 598.050 367.050 ;
        RECT 463.950 365.400 537.600 366.600 ;
        RECT 463.950 364.950 466.050 365.400 ;
        RECT 121.950 363.600 124.050 364.050 ;
        RECT 196.950 363.600 199.050 364.050 ;
        RECT 121.950 362.400 199.050 363.600 ;
        RECT 121.950 361.950 124.050 362.400 ;
        RECT 196.950 361.950 199.050 362.400 ;
        RECT 202.950 363.600 205.050 364.050 ;
        RECT 532.950 363.600 535.050 364.050 ;
        RECT 202.950 362.400 535.050 363.600 ;
        RECT 536.400 363.600 537.600 365.400 ;
        RECT 589.950 365.400 598.050 366.600 ;
        RECT 589.950 364.950 592.050 365.400 ;
        RECT 595.950 364.950 598.050 365.400 ;
        RECT 643.950 366.600 646.050 367.050 ;
        RECT 661.950 366.600 664.050 367.050 ;
        RECT 643.950 365.400 664.050 366.600 ;
        RECT 643.950 364.950 646.050 365.400 ;
        RECT 661.950 364.950 664.050 365.400 ;
        RECT 751.950 366.600 754.050 367.050 ;
        RECT 850.950 366.600 853.050 367.050 ;
        RECT 751.950 365.400 853.050 366.600 ;
        RECT 751.950 364.950 754.050 365.400 ;
        RECT 850.950 364.950 853.050 365.400 ;
        RECT 682.950 363.600 685.050 364.050 ;
        RECT 536.400 362.400 685.050 363.600 ;
        RECT 202.950 361.950 205.050 362.400 ;
        RECT 532.950 361.950 535.050 362.400 ;
        RECT 682.950 361.950 685.050 362.400 ;
        RECT 220.950 360.600 223.050 361.050 ;
        RECT 226.950 360.600 229.050 361.050 ;
        RECT 220.950 359.400 229.050 360.600 ;
        RECT 220.950 358.950 223.050 359.400 ;
        RECT 226.950 358.950 229.050 359.400 ;
        RECT 385.950 360.600 388.050 361.050 ;
        RECT 436.950 360.600 439.050 361.050 ;
        RECT 385.950 359.400 439.050 360.600 ;
        RECT 385.950 358.950 388.050 359.400 ;
        RECT 436.950 358.950 439.050 359.400 ;
        RECT 445.950 360.600 448.050 361.050 ;
        RECT 628.950 360.600 631.050 361.050 ;
        RECT 739.950 360.600 742.050 361.050 ;
        RECT 445.950 359.400 564.600 360.600 ;
        RECT 445.950 358.950 448.050 359.400 ;
        RECT 1.950 357.600 4.050 358.050 ;
        RECT 196.950 357.600 199.050 358.050 ;
        RECT 1.950 356.400 199.050 357.600 ;
        RECT 1.950 355.950 4.050 356.400 ;
        RECT 196.950 355.950 199.050 356.400 ;
        RECT 331.950 357.600 334.050 358.050 ;
        RECT 385.950 357.600 388.050 358.050 ;
        RECT 433.950 357.600 436.050 358.050 ;
        RECT 331.950 356.400 436.050 357.600 ;
        RECT 331.950 355.950 334.050 356.400 ;
        RECT 385.950 355.950 388.050 356.400 ;
        RECT 433.950 355.950 436.050 356.400 ;
        RECT 526.950 357.600 529.050 358.050 ;
        RECT 559.950 357.600 562.050 358.050 ;
        RECT 526.950 356.400 562.050 357.600 ;
        RECT 563.400 357.600 564.600 359.400 ;
        RECT 628.950 359.400 742.050 360.600 ;
        RECT 628.950 358.950 631.050 359.400 ;
        RECT 739.950 358.950 742.050 359.400 ;
        RECT 769.950 357.600 772.050 358.050 ;
        RECT 563.400 356.400 772.050 357.600 ;
        RECT 526.950 355.950 529.050 356.400 ;
        RECT 559.950 355.950 562.050 356.400 ;
        RECT 769.950 355.950 772.050 356.400 ;
        RECT 49.950 354.600 52.050 355.050 ;
        RECT 445.950 354.600 448.050 355.050 ;
        RECT 49.950 353.400 448.050 354.600 ;
        RECT 49.950 352.950 52.050 353.400 ;
        RECT 445.950 352.950 448.050 353.400 ;
        RECT 487.950 354.600 490.050 355.050 ;
        RECT 505.950 354.600 508.050 355.050 ;
        RECT 487.950 353.400 508.050 354.600 ;
        RECT 487.950 352.950 490.050 353.400 ;
        RECT 505.950 352.950 508.050 353.400 ;
        RECT 520.950 354.600 523.050 355.050 ;
        RECT 538.950 354.600 541.050 355.050 ;
        RECT 547.950 354.600 550.050 355.050 ;
        RECT 577.950 354.600 580.050 355.050 ;
        RECT 604.950 354.600 607.050 355.050 ;
        RECT 520.950 353.400 541.050 354.600 ;
        RECT 520.950 352.950 523.050 353.400 ;
        RECT 538.950 352.950 541.050 353.400 ;
        RECT 542.400 353.400 607.050 354.600 ;
        RECT 127.950 351.600 130.050 352.050 ;
        RECT 208.950 351.600 211.050 352.050 ;
        RECT 127.950 350.400 211.050 351.600 ;
        RECT 127.950 349.950 130.050 350.400 ;
        RECT 208.950 349.950 211.050 350.400 ;
        RECT 277.950 351.600 280.050 352.050 ;
        RECT 542.400 351.600 543.600 353.400 ;
        RECT 547.950 352.950 550.050 353.400 ;
        RECT 577.950 352.950 580.050 353.400 ;
        RECT 604.950 352.950 607.050 353.400 ;
        RECT 715.950 354.600 718.050 355.050 ;
        RECT 736.950 354.600 739.050 355.050 ;
        RECT 715.950 353.400 739.050 354.600 ;
        RECT 715.950 352.950 718.050 353.400 ;
        RECT 736.950 352.950 739.050 353.400 ;
        RECT 784.950 354.600 787.050 355.050 ;
        RECT 826.950 354.600 829.050 355.050 ;
        RECT 784.950 353.400 829.050 354.600 ;
        RECT 784.950 352.950 787.050 353.400 ;
        RECT 826.950 352.950 829.050 353.400 ;
        RECT 601.950 351.600 604.050 352.050 ;
        RECT 676.950 351.600 679.050 352.050 ;
        RECT 277.950 350.400 543.600 351.600 ;
        RECT 545.400 350.400 679.050 351.600 ;
        RECT 277.950 349.950 280.050 350.400 ;
        RECT 31.950 348.600 34.050 349.050 ;
        RECT 37.950 348.600 40.050 349.050 ;
        RECT 31.950 347.400 40.050 348.600 ;
        RECT 31.950 346.950 34.050 347.400 ;
        RECT 37.950 346.950 40.050 347.400 ;
        RECT 130.950 348.600 133.050 349.050 ;
        RECT 148.950 348.600 151.050 349.050 ;
        RECT 157.950 348.600 160.050 349.050 ;
        RECT 130.950 347.400 147.600 348.600 ;
        RECT 130.950 346.950 133.050 347.400 ;
        RECT 25.950 345.600 28.050 346.050 ;
        RECT 34.950 345.600 37.050 346.050 ;
        RECT 25.950 344.400 37.050 345.600 ;
        RECT 25.950 343.950 28.050 344.400 ;
        RECT 34.950 343.950 37.050 344.400 ;
        RECT 58.950 345.600 61.050 346.050 ;
        RECT 67.950 345.600 70.050 346.050 ;
        RECT 58.950 344.400 70.050 345.600 ;
        RECT 58.950 343.950 61.050 344.400 ;
        RECT 67.950 343.950 70.050 344.400 ;
        RECT 133.950 343.950 136.050 346.050 ;
        RECT 146.400 345.600 147.600 347.400 ;
        RECT 148.950 347.400 160.050 348.600 ;
        RECT 148.950 346.950 151.050 347.400 ;
        RECT 157.950 346.950 160.050 347.400 ;
        RECT 160.950 348.600 163.050 349.050 ;
        RECT 166.950 348.600 169.050 349.050 ;
        RECT 160.950 347.400 169.050 348.600 ;
        RECT 160.950 346.950 163.050 347.400 ;
        RECT 166.950 346.950 169.050 347.400 ;
        RECT 265.950 348.600 268.050 349.050 ;
        RECT 283.950 348.600 286.050 349.050 ;
        RECT 265.950 347.400 286.050 348.600 ;
        RECT 265.950 346.950 268.050 347.400 ;
        RECT 283.950 346.950 286.050 347.400 ;
        RECT 340.950 348.600 343.050 349.050 ;
        RECT 397.950 348.600 400.050 349.050 ;
        RECT 340.950 347.400 400.050 348.600 ;
        RECT 340.950 346.950 343.050 347.400 ;
        RECT 397.950 346.950 400.050 347.400 ;
        RECT 451.950 348.600 454.050 349.050 ;
        RECT 499.950 348.600 502.050 349.050 ;
        RECT 545.400 348.600 546.600 350.400 ;
        RECT 601.950 349.950 604.050 350.400 ;
        RECT 676.950 349.950 679.050 350.400 ;
        RECT 802.950 351.600 805.050 352.050 ;
        RECT 820.950 351.600 823.050 352.050 ;
        RECT 802.950 350.400 823.050 351.600 ;
        RECT 802.950 349.950 805.050 350.400 ;
        RECT 820.950 349.950 823.050 350.400 ;
        RECT 451.950 347.400 546.600 348.600 ;
        RECT 559.950 348.600 562.050 349.050 ;
        RECT 568.950 348.600 571.050 349.050 ;
        RECT 559.950 347.400 571.050 348.600 ;
        RECT 451.950 346.950 454.050 347.400 ;
        RECT 499.950 346.950 502.050 347.400 ;
        RECT 559.950 346.950 562.050 347.400 ;
        RECT 568.950 346.950 571.050 347.400 ;
        RECT 571.950 348.600 574.050 349.050 ;
        RECT 727.950 348.600 730.050 349.050 ;
        RECT 571.950 347.400 730.050 348.600 ;
        RECT 571.950 346.950 574.050 347.400 ;
        RECT 727.950 346.950 730.050 347.400 ;
        RECT 799.950 348.600 802.050 349.050 ;
        RECT 829.950 348.600 832.050 349.050 ;
        RECT 799.950 347.400 832.050 348.600 ;
        RECT 799.950 346.950 802.050 347.400 ;
        RECT 829.950 346.950 832.050 347.400 ;
        RECT 148.950 345.600 151.050 346.050 ;
        RECT 146.400 344.400 151.050 345.600 ;
        RECT 148.950 343.950 151.050 344.400 ;
        RECT 154.950 343.950 157.050 346.050 ;
        RECT 160.950 345.600 163.050 346.050 ;
        RECT 280.950 345.600 283.050 346.050 ;
        RECT 307.950 345.600 310.050 346.050 ;
        RECT 160.950 344.400 168.600 345.600 ;
        RECT 160.950 343.950 163.050 344.400 ;
        RECT 22.950 342.600 25.050 343.050 ;
        RECT 52.950 342.600 55.050 343.050 ;
        RECT 73.950 342.600 76.050 343.050 ;
        RECT 22.950 341.400 76.050 342.600 ;
        RECT 22.950 340.950 25.050 341.400 ;
        RECT 52.950 340.950 55.050 341.400 ;
        RECT 73.950 340.950 76.050 341.400 ;
        RECT 100.950 342.600 103.050 343.050 ;
        RECT 115.950 342.600 118.050 343.050 ;
        RECT 100.950 341.400 118.050 342.600 ;
        RECT 100.950 340.950 103.050 341.400 ;
        RECT 115.950 340.950 118.050 341.400 ;
        RECT 118.950 342.600 121.050 343.050 ;
        RECT 127.950 342.600 130.050 343.050 ;
        RECT 118.950 341.400 130.050 342.600 ;
        RECT 134.400 342.600 135.600 343.950 ;
        RECT 155.400 342.600 156.600 343.950 ;
        RECT 163.950 342.600 166.050 343.050 ;
        RECT 134.400 341.400 150.600 342.600 ;
        RECT 155.400 341.400 166.050 342.600 ;
        RECT 118.950 340.950 121.050 341.400 ;
        RECT 127.950 340.950 130.050 341.400 ;
        RECT 13.950 339.600 16.050 340.050 ;
        RECT 28.950 339.600 31.050 340.050 ;
        RECT 13.950 338.400 31.050 339.600 ;
        RECT 13.950 337.950 16.050 338.400 ;
        RECT 28.950 337.950 31.050 338.400 ;
        RECT 34.950 339.600 37.050 340.050 ;
        RECT 40.950 339.600 43.050 340.050 ;
        RECT 34.950 338.400 43.050 339.600 ;
        RECT 34.950 337.950 37.050 338.400 ;
        RECT 40.950 337.950 43.050 338.400 ;
        RECT 64.950 339.600 67.050 340.050 ;
        RECT 85.950 339.600 88.050 340.050 ;
        RECT 64.950 338.400 88.050 339.600 ;
        RECT 64.950 337.950 67.050 338.400 ;
        RECT 85.950 337.950 88.050 338.400 ;
        RECT 130.950 339.600 133.050 340.050 ;
        RECT 136.950 339.600 139.050 340.050 ;
        RECT 130.950 338.400 139.050 339.600 ;
        RECT 149.400 339.600 150.600 341.400 ;
        RECT 163.950 340.950 166.050 341.400 ;
        RECT 160.950 339.600 163.050 340.050 ;
        RECT 149.400 338.400 163.050 339.600 ;
        RECT 130.950 337.950 133.050 338.400 ;
        RECT 136.950 337.950 139.050 338.400 ;
        RECT 160.950 337.950 163.050 338.400 ;
        RECT 163.950 339.600 166.050 340.050 ;
        RECT 167.400 339.600 168.600 344.400 ;
        RECT 280.950 344.400 310.050 345.600 ;
        RECT 280.950 343.950 283.050 344.400 ;
        RECT 307.950 343.950 310.050 344.400 ;
        RECT 313.950 345.600 316.050 346.050 ;
        RECT 322.950 345.600 325.050 346.050 ;
        RECT 313.950 344.400 325.050 345.600 ;
        RECT 313.950 343.950 316.050 344.400 ;
        RECT 322.950 343.950 325.050 344.400 ;
        RECT 352.950 345.600 355.050 346.050 ;
        RECT 355.950 345.600 358.050 346.050 ;
        RECT 403.950 345.600 406.050 346.050 ;
        RECT 352.950 344.400 406.050 345.600 ;
        RECT 352.950 343.950 355.050 344.400 ;
        RECT 355.950 343.950 358.050 344.400 ;
        RECT 403.950 343.950 406.050 344.400 ;
        RECT 409.950 345.600 412.050 346.050 ;
        RECT 418.950 345.600 421.050 346.050 ;
        RECT 493.950 345.600 496.050 346.050 ;
        RECT 409.950 344.400 496.050 345.600 ;
        RECT 409.950 343.950 412.050 344.400 ;
        RECT 418.950 343.950 421.050 344.400 ;
        RECT 493.950 343.950 496.050 344.400 ;
        RECT 541.950 345.600 544.050 346.050 ;
        RECT 562.950 345.600 565.050 346.050 ;
        RECT 574.950 345.600 577.050 346.050 ;
        RECT 541.950 344.400 577.050 345.600 ;
        RECT 541.950 343.950 544.050 344.400 ;
        RECT 562.950 343.950 565.050 344.400 ;
        RECT 574.950 343.950 577.050 344.400 ;
        RECT 607.950 345.600 610.050 346.050 ;
        RECT 625.950 345.600 628.050 346.050 ;
        RECT 607.950 344.400 628.050 345.600 ;
        RECT 607.950 343.950 610.050 344.400 ;
        RECT 625.950 343.950 628.050 344.400 ;
        RECT 670.950 345.600 673.050 346.050 ;
        RECT 679.950 345.600 682.050 346.050 ;
        RECT 670.950 344.400 682.050 345.600 ;
        RECT 670.950 343.950 673.050 344.400 ;
        RECT 679.950 343.950 682.050 344.400 ;
        RECT 682.950 345.600 685.050 346.050 ;
        RECT 703.950 345.600 706.050 346.050 ;
        RECT 682.950 344.400 706.050 345.600 ;
        RECT 682.950 343.950 685.050 344.400 ;
        RECT 703.950 343.950 706.050 344.400 ;
        RECT 781.950 345.600 784.050 346.050 ;
        RECT 793.950 345.600 796.050 346.050 ;
        RECT 781.950 344.400 796.050 345.600 ;
        RECT 781.950 343.950 784.050 344.400 ;
        RECT 793.950 343.950 796.050 344.400 ;
        RECT 805.950 345.600 808.050 346.050 ;
        RECT 811.950 345.600 814.050 346.050 ;
        RECT 805.950 344.400 814.050 345.600 ;
        RECT 805.950 343.950 808.050 344.400 ;
        RECT 811.950 343.950 814.050 344.400 ;
        RECT 817.950 345.600 820.050 346.050 ;
        RECT 823.950 345.600 826.050 346.050 ;
        RECT 817.950 344.400 826.050 345.600 ;
        RECT 817.950 343.950 820.050 344.400 ;
        RECT 823.950 343.950 826.050 344.400 ;
        RECT 826.950 345.600 829.050 346.050 ;
        RECT 835.950 345.600 838.050 346.050 ;
        RECT 826.950 344.400 838.050 345.600 ;
        RECT 826.950 343.950 829.050 344.400 ;
        RECT 835.950 343.950 838.050 344.400 ;
        RECT 178.950 340.950 181.050 343.050 ;
        RECT 184.950 340.950 187.050 343.050 ;
        RECT 229.950 342.600 232.050 343.050 ;
        RECT 197.400 341.400 232.050 342.600 ;
        RECT 163.950 338.400 168.600 339.600 ;
        RECT 163.950 337.950 166.050 338.400 ;
        RECT 179.400 337.050 180.600 340.950 ;
        RECT 185.400 339.600 186.600 340.950 ;
        RECT 185.400 338.400 189.600 339.600 ;
        RECT 16.950 336.600 19.050 337.050 ;
        RECT 22.950 336.600 25.050 337.050 ;
        RECT 16.950 335.400 25.050 336.600 ;
        RECT 16.950 334.950 19.050 335.400 ;
        RECT 22.950 334.950 25.050 335.400 ;
        RECT 34.950 336.600 37.050 337.050 ;
        RECT 37.950 336.600 40.050 337.050 ;
        RECT 46.950 336.600 49.050 337.050 ;
        RECT 34.950 335.400 49.050 336.600 ;
        RECT 34.950 334.950 37.050 335.400 ;
        RECT 37.950 334.950 40.050 335.400 ;
        RECT 46.950 334.950 49.050 335.400 ;
        RECT 76.950 336.600 79.050 337.050 ;
        RECT 79.950 336.600 82.050 337.050 ;
        RECT 112.950 336.600 115.050 337.050 ;
        RECT 76.950 335.400 115.050 336.600 ;
        RECT 76.950 334.950 79.050 335.400 ;
        RECT 79.950 334.950 82.050 335.400 ;
        RECT 112.950 334.950 115.050 335.400 ;
        RECT 154.950 336.600 157.050 337.050 ;
        RECT 166.950 336.600 169.050 337.050 ;
        RECT 154.950 335.400 169.050 336.600 ;
        RECT 154.950 334.950 157.050 335.400 ;
        RECT 166.950 334.950 169.050 335.400 ;
        RECT 178.950 334.950 181.050 337.050 ;
        RECT 188.400 336.600 189.600 338.400 ;
        RECT 190.950 336.600 193.050 337.050 ;
        RECT 188.400 335.400 193.050 336.600 ;
        RECT 190.950 334.950 193.050 335.400 ;
        RECT 28.950 333.600 31.050 334.050 ;
        RECT 55.950 333.600 58.050 334.050 ;
        RECT 28.950 332.400 58.050 333.600 ;
        RECT 28.950 331.950 31.050 332.400 ;
        RECT 55.950 331.950 58.050 332.400 ;
        RECT 88.950 333.600 91.050 334.050 ;
        RECT 163.950 333.600 166.050 334.050 ;
        RECT 88.950 332.400 166.050 333.600 ;
        RECT 88.950 331.950 91.050 332.400 ;
        RECT 163.950 331.950 166.050 332.400 ;
        RECT 175.950 333.600 178.050 334.050 ;
        RECT 197.400 333.600 198.600 341.400 ;
        RECT 229.950 340.950 232.050 341.400 ;
        RECT 250.950 342.600 253.050 343.050 ;
        RECT 256.950 342.600 259.050 343.050 ;
        RECT 250.950 341.400 259.050 342.600 ;
        RECT 250.950 340.950 253.050 341.400 ;
        RECT 256.950 340.950 259.050 341.400 ;
        RECT 271.950 342.600 274.050 343.050 ;
        RECT 283.950 342.600 286.050 343.050 ;
        RECT 271.950 341.400 286.050 342.600 ;
        RECT 271.950 340.950 274.050 341.400 ;
        RECT 283.950 340.950 286.050 341.400 ;
        RECT 289.950 342.600 292.050 343.050 ;
        RECT 301.950 342.600 304.050 343.050 ;
        RECT 289.950 341.400 304.050 342.600 ;
        RECT 289.950 340.950 292.050 341.400 ;
        RECT 301.950 340.950 304.050 341.400 ;
        RECT 307.950 342.600 310.050 343.050 ;
        RECT 307.950 341.400 336.600 342.600 ;
        RECT 307.950 340.950 310.050 341.400 ;
        RECT 199.950 339.600 202.050 340.050 ;
        RECT 211.950 339.600 214.050 340.050 ;
        RECT 199.950 338.400 214.050 339.600 ;
        RECT 199.950 337.950 202.050 338.400 ;
        RECT 211.950 337.950 214.050 338.400 ;
        RECT 223.950 339.600 226.050 340.050 ;
        RECT 331.950 339.600 334.050 340.050 ;
        RECT 223.950 338.400 334.050 339.600 ;
        RECT 335.400 339.600 336.600 341.400 ;
        RECT 346.950 340.950 349.050 343.050 ;
        RECT 361.950 342.600 364.050 343.050 ;
        RECT 421.950 342.600 424.050 343.050 ;
        RECT 361.950 341.400 424.050 342.600 ;
        RECT 361.950 340.950 364.050 341.400 ;
        RECT 421.950 340.950 424.050 341.400 ;
        RECT 451.950 342.600 454.050 343.050 ;
        RECT 457.950 342.600 460.050 343.050 ;
        RECT 451.950 341.400 460.050 342.600 ;
        RECT 451.950 340.950 454.050 341.400 ;
        RECT 457.950 340.950 460.050 341.400 ;
        RECT 508.950 340.950 511.050 343.050 ;
        RECT 523.950 342.600 526.050 343.050 ;
        RECT 586.950 342.600 589.050 343.050 ;
        RECT 592.950 342.600 595.050 343.050 ;
        RECT 523.950 341.400 531.600 342.600 ;
        RECT 523.950 340.950 526.050 341.400 ;
        RECT 343.950 339.600 346.050 340.050 ;
        RECT 335.400 338.400 346.050 339.600 ;
        RECT 223.950 337.950 226.050 338.400 ;
        RECT 331.950 337.950 334.050 338.400 ;
        RECT 343.950 337.950 346.050 338.400 ;
        RECT 347.400 337.050 348.600 340.950 ;
        RECT 362.400 339.600 363.600 340.950 ;
        RECT 350.400 338.400 363.600 339.600 ;
        RECT 367.950 339.600 370.050 340.050 ;
        RECT 388.950 339.600 391.050 340.050 ;
        RECT 367.950 338.400 391.050 339.600 ;
        RECT 350.400 337.050 351.600 338.400 ;
        RECT 367.950 337.950 370.050 338.400 ;
        RECT 388.950 337.950 391.050 338.400 ;
        RECT 397.950 339.600 400.050 340.050 ;
        RECT 415.950 339.600 418.050 340.050 ;
        RECT 430.950 339.600 433.050 340.050 ;
        RECT 397.950 338.400 402.600 339.600 ;
        RECT 397.950 337.950 400.050 338.400 ;
        RECT 208.950 336.600 211.050 337.050 ;
        RECT 214.950 336.600 217.050 337.050 ;
        RECT 208.950 335.400 217.050 336.600 ;
        RECT 208.950 334.950 211.050 335.400 ;
        RECT 214.950 334.950 217.050 335.400 ;
        RECT 220.950 336.600 223.050 337.050 ;
        RECT 232.950 336.600 235.050 337.050 ;
        RECT 220.950 335.400 235.050 336.600 ;
        RECT 220.950 334.950 223.050 335.400 ;
        RECT 232.950 334.950 235.050 335.400 ;
        RECT 238.950 336.600 241.050 337.050 ;
        RECT 253.950 336.600 256.050 337.050 ;
        RECT 238.950 335.400 256.050 336.600 ;
        RECT 238.950 334.950 241.050 335.400 ;
        RECT 253.950 334.950 256.050 335.400 ;
        RECT 262.950 336.600 265.050 337.050 ;
        RECT 274.950 336.600 277.050 337.050 ;
        RECT 262.950 335.400 277.050 336.600 ;
        RECT 262.950 334.950 265.050 335.400 ;
        RECT 274.950 334.950 277.050 335.400 ;
        RECT 346.950 334.950 349.050 337.050 ;
        RECT 349.950 334.950 352.050 337.050 ;
        RECT 373.950 336.600 376.050 337.050 ;
        RECT 397.950 336.600 400.050 337.050 ;
        RECT 373.950 335.400 400.050 336.600 ;
        RECT 401.400 336.600 402.600 338.400 ;
        RECT 415.950 338.400 433.050 339.600 ;
        RECT 415.950 337.950 418.050 338.400 ;
        RECT 430.950 337.950 433.050 338.400 ;
        RECT 436.950 339.600 439.050 340.050 ;
        RECT 454.950 339.600 457.050 340.050 ;
        RECT 436.950 338.400 457.050 339.600 ;
        RECT 436.950 337.950 439.050 338.400 ;
        RECT 454.950 337.950 457.050 338.400 ;
        RECT 490.950 339.600 493.050 340.050 ;
        RECT 509.400 339.600 510.600 340.950 ;
        RECT 530.400 340.050 531.600 341.400 ;
        RECT 586.950 341.400 595.050 342.600 ;
        RECT 586.950 340.950 589.050 341.400 ;
        RECT 592.950 340.950 595.050 341.400 ;
        RECT 601.950 342.600 604.050 343.050 ;
        RECT 607.950 342.600 610.050 343.050 ;
        RECT 601.950 341.400 610.050 342.600 ;
        RECT 601.950 340.950 604.050 341.400 ;
        RECT 607.950 340.950 610.050 341.400 ;
        RECT 619.950 342.600 622.050 343.050 ;
        RECT 742.950 342.600 745.050 343.050 ;
        RECT 760.950 342.600 763.050 343.050 ;
        RECT 619.950 341.400 624.600 342.600 ;
        RECT 619.950 340.950 622.050 341.400 ;
        RECT 490.950 338.400 510.600 339.600 ;
        RECT 490.950 337.950 493.050 338.400 ;
        RECT 529.950 337.950 532.050 340.050 ;
        RECT 559.950 339.600 562.050 340.050 ;
        RECT 583.950 339.600 586.050 340.050 ;
        RECT 559.950 338.400 586.050 339.600 ;
        RECT 559.950 337.950 562.050 338.400 ;
        RECT 583.950 337.950 586.050 338.400 ;
        RECT 589.950 339.600 592.050 340.050 ;
        RECT 598.950 339.600 601.050 340.050 ;
        RECT 619.950 339.600 622.050 340.050 ;
        RECT 589.950 338.400 622.050 339.600 ;
        RECT 589.950 337.950 592.050 338.400 ;
        RECT 598.950 337.950 601.050 338.400 ;
        RECT 619.950 337.950 622.050 338.400 ;
        RECT 412.950 336.600 415.050 337.050 ;
        RECT 401.400 335.400 415.050 336.600 ;
        RECT 373.950 334.950 376.050 335.400 ;
        RECT 397.950 334.950 400.050 335.400 ;
        RECT 412.950 334.950 415.050 335.400 ;
        RECT 442.950 336.600 445.050 337.050 ;
        RECT 484.950 336.600 487.050 337.050 ;
        RECT 442.950 335.400 487.050 336.600 ;
        RECT 442.950 334.950 445.050 335.400 ;
        RECT 484.950 334.950 487.050 335.400 ;
        RECT 487.950 336.600 490.050 337.050 ;
        RECT 502.950 336.600 505.050 337.050 ;
        RECT 487.950 335.400 505.050 336.600 ;
        RECT 487.950 334.950 490.050 335.400 ;
        RECT 502.950 334.950 505.050 335.400 ;
        RECT 529.950 336.600 532.050 337.050 ;
        RECT 532.950 336.600 535.050 337.050 ;
        RECT 556.950 336.600 559.050 337.050 ;
        RECT 529.950 335.400 559.050 336.600 ;
        RECT 529.950 334.950 532.050 335.400 ;
        RECT 532.950 334.950 535.050 335.400 ;
        RECT 556.950 334.950 559.050 335.400 ;
        RECT 580.950 336.600 583.050 337.050 ;
        RECT 592.950 336.600 595.050 337.050 ;
        RECT 580.950 335.400 595.050 336.600 ;
        RECT 623.400 336.600 624.600 341.400 ;
        RECT 742.950 341.400 763.050 342.600 ;
        RECT 742.950 340.950 745.050 341.400 ;
        RECT 758.400 340.050 759.600 341.400 ;
        RECT 760.950 340.950 763.050 341.400 ;
        RECT 766.950 342.600 769.050 343.050 ;
        RECT 814.950 342.600 817.050 343.050 ;
        RECT 766.950 341.400 817.050 342.600 ;
        RECT 766.950 340.950 769.050 341.400 ;
        RECT 814.950 340.950 817.050 341.400 ;
        RECT 829.950 340.950 832.050 343.050 ;
        RECT 841.950 340.950 844.050 343.050 ;
        RECT 757.950 339.600 760.050 340.050 ;
        RECT 826.950 339.600 829.050 340.050 ;
        RECT 757.950 338.400 829.050 339.600 ;
        RECT 757.950 337.950 760.050 338.400 ;
        RECT 826.950 337.950 829.050 338.400 ;
        RECT 730.950 336.600 733.050 337.050 ;
        RECT 623.400 335.400 733.050 336.600 ;
        RECT 580.950 334.950 583.050 335.400 ;
        RECT 592.950 334.950 595.050 335.400 ;
        RECT 730.950 334.950 733.050 335.400 ;
        RECT 751.950 336.600 754.050 337.050 ;
        RECT 763.950 336.600 766.050 337.050 ;
        RECT 751.950 335.400 766.050 336.600 ;
        RECT 751.950 334.950 754.050 335.400 ;
        RECT 763.950 334.950 766.050 335.400 ;
        RECT 775.950 336.600 778.050 337.050 ;
        RECT 781.950 336.600 784.050 337.050 ;
        RECT 775.950 335.400 784.050 336.600 ;
        RECT 775.950 334.950 778.050 335.400 ;
        RECT 781.950 334.950 784.050 335.400 ;
        RECT 793.950 336.600 796.050 337.050 ;
        RECT 823.950 336.600 826.050 337.050 ;
        RECT 793.950 335.400 826.050 336.600 ;
        RECT 793.950 334.950 796.050 335.400 ;
        RECT 823.950 334.950 826.050 335.400 ;
        RECT 826.950 336.600 829.050 337.050 ;
        RECT 830.400 336.600 831.600 340.950 ;
        RECT 826.950 335.400 831.600 336.600 ;
        RECT 842.400 336.600 843.600 340.950 ;
        RECT 844.950 339.600 847.050 340.050 ;
        RECT 850.950 339.600 853.050 340.050 ;
        RECT 844.950 338.400 853.050 339.600 ;
        RECT 844.950 337.950 847.050 338.400 ;
        RECT 850.950 337.950 853.050 338.400 ;
        RECT 844.950 336.600 847.050 337.050 ;
        RECT 842.400 335.400 847.050 336.600 ;
        RECT 826.950 334.950 829.050 335.400 ;
        RECT 844.950 334.950 847.050 335.400 ;
        RECT 175.950 332.400 198.600 333.600 ;
        RECT 217.950 333.600 220.050 334.050 ;
        RECT 226.950 333.600 229.050 334.050 ;
        RECT 277.950 333.600 280.050 334.050 ;
        RECT 217.950 332.400 280.050 333.600 ;
        RECT 175.950 331.950 178.050 332.400 ;
        RECT 217.950 331.950 220.050 332.400 ;
        RECT 226.950 331.950 229.050 332.400 ;
        RECT 277.950 331.950 280.050 332.400 ;
        RECT 337.950 333.600 340.050 334.050 ;
        RECT 376.950 333.600 379.050 334.050 ;
        RECT 409.950 333.600 412.050 334.050 ;
        RECT 337.950 332.400 412.050 333.600 ;
        RECT 337.950 331.950 340.050 332.400 ;
        RECT 376.950 331.950 379.050 332.400 ;
        RECT 409.950 331.950 412.050 332.400 ;
        RECT 421.950 333.600 424.050 334.050 ;
        RECT 466.950 333.600 469.050 334.050 ;
        RECT 574.950 333.600 577.050 334.050 ;
        RECT 421.950 332.400 577.050 333.600 ;
        RECT 421.950 331.950 424.050 332.400 ;
        RECT 466.950 331.950 469.050 332.400 ;
        RECT 574.950 331.950 577.050 332.400 ;
        RECT 586.950 333.600 589.050 334.050 ;
        RECT 595.950 333.600 598.050 334.050 ;
        RECT 586.950 332.400 598.050 333.600 ;
        RECT 586.950 331.950 589.050 332.400 ;
        RECT 595.950 331.950 598.050 332.400 ;
        RECT 760.950 333.600 763.050 334.050 ;
        RECT 772.950 333.600 775.050 334.050 ;
        RECT 760.950 332.400 775.050 333.600 ;
        RECT 760.950 331.950 763.050 332.400 ;
        RECT 772.950 331.950 775.050 332.400 ;
        RECT 811.950 333.600 814.050 334.050 ;
        RECT 823.950 333.600 826.050 334.050 ;
        RECT 811.950 332.400 826.050 333.600 ;
        RECT 811.950 331.950 814.050 332.400 ;
        RECT 823.950 331.950 826.050 332.400 ;
        RECT 835.950 333.600 838.050 334.050 ;
        RECT 841.950 333.600 844.050 334.050 ;
        RECT 835.950 332.400 844.050 333.600 ;
        RECT 835.950 331.950 838.050 332.400 ;
        RECT 841.950 331.950 844.050 332.400 ;
        RECT 10.950 330.600 13.050 331.050 ;
        RECT 37.950 330.600 40.050 331.050 ;
        RECT 91.950 330.600 94.050 331.050 ;
        RECT 10.950 329.400 94.050 330.600 ;
        RECT 10.950 328.950 13.050 329.400 ;
        RECT 37.950 328.950 40.050 329.400 ;
        RECT 91.950 328.950 94.050 329.400 ;
        RECT 190.950 330.600 193.050 331.050 ;
        RECT 202.950 330.600 205.050 331.050 ;
        RECT 190.950 329.400 205.050 330.600 ;
        RECT 190.950 328.950 193.050 329.400 ;
        RECT 202.950 328.950 205.050 329.400 ;
        RECT 241.950 330.600 244.050 331.050 ;
        RECT 295.950 330.600 298.050 331.050 ;
        RECT 241.950 329.400 298.050 330.600 ;
        RECT 241.950 328.950 244.050 329.400 ;
        RECT 295.950 328.950 298.050 329.400 ;
        RECT 346.950 330.600 349.050 331.050 ;
        RECT 364.950 330.600 367.050 331.050 ;
        RECT 346.950 329.400 367.050 330.600 ;
        RECT 346.950 328.950 349.050 329.400 ;
        RECT 364.950 328.950 367.050 329.400 ;
        RECT 367.950 330.600 370.050 331.050 ;
        RECT 379.950 330.600 382.050 331.050 ;
        RECT 367.950 329.400 382.050 330.600 ;
        RECT 367.950 328.950 370.050 329.400 ;
        RECT 379.950 328.950 382.050 329.400 ;
        RECT 382.950 330.600 385.050 331.050 ;
        RECT 400.950 330.600 403.050 331.050 ;
        RECT 382.950 329.400 403.050 330.600 ;
        RECT 382.950 328.950 385.050 329.400 ;
        RECT 400.950 328.950 403.050 329.400 ;
        RECT 403.950 330.600 406.050 331.050 ;
        RECT 424.950 330.600 427.050 331.050 ;
        RECT 457.950 330.600 460.050 331.050 ;
        RECT 403.950 329.400 460.050 330.600 ;
        RECT 403.950 328.950 406.050 329.400 ;
        RECT 424.950 328.950 427.050 329.400 ;
        RECT 457.950 328.950 460.050 329.400 ;
        RECT 475.950 330.600 478.050 331.050 ;
        RECT 523.950 330.600 526.050 331.050 ;
        RECT 475.950 329.400 526.050 330.600 ;
        RECT 475.950 328.950 478.050 329.400 ;
        RECT 523.950 328.950 526.050 329.400 ;
        RECT 646.950 330.600 649.050 331.050 ;
        RECT 652.950 330.600 655.050 331.050 ;
        RECT 646.950 329.400 655.050 330.600 ;
        RECT 646.950 328.950 649.050 329.400 ;
        RECT 652.950 328.950 655.050 329.400 ;
        RECT 769.950 330.600 772.050 331.050 ;
        RECT 811.950 330.600 814.050 331.050 ;
        RECT 817.950 330.600 820.050 331.050 ;
        RECT 769.950 329.400 820.050 330.600 ;
        RECT 769.950 328.950 772.050 329.400 ;
        RECT 811.950 328.950 814.050 329.400 ;
        RECT 817.950 328.950 820.050 329.400 ;
        RECT 829.950 330.600 832.050 331.050 ;
        RECT 838.950 330.600 841.050 331.050 ;
        RECT 829.950 329.400 841.050 330.600 ;
        RECT 829.950 328.950 832.050 329.400 ;
        RECT 838.950 328.950 841.050 329.400 ;
        RECT 841.950 330.600 844.050 331.050 ;
        RECT 853.950 330.600 856.050 331.050 ;
        RECT 841.950 329.400 856.050 330.600 ;
        RECT 841.950 328.950 844.050 329.400 ;
        RECT 853.950 328.950 856.050 329.400 ;
        RECT 43.950 327.600 46.050 328.050 ;
        RECT 67.950 327.600 70.050 328.050 ;
        RECT 97.950 327.600 100.050 328.050 ;
        RECT 43.950 326.400 100.050 327.600 ;
        RECT 43.950 325.950 46.050 326.400 ;
        RECT 67.950 325.950 70.050 326.400 ;
        RECT 97.950 325.950 100.050 326.400 ;
        RECT 103.950 327.600 106.050 328.050 ;
        RECT 247.950 327.600 250.050 328.050 ;
        RECT 103.950 326.400 250.050 327.600 ;
        RECT 103.950 325.950 106.050 326.400 ;
        RECT 247.950 325.950 250.050 326.400 ;
        RECT 256.950 327.600 259.050 328.050 ;
        RECT 316.950 327.600 319.050 328.050 ;
        RECT 256.950 326.400 319.050 327.600 ;
        RECT 256.950 325.950 259.050 326.400 ;
        RECT 316.950 325.950 319.050 326.400 ;
        RECT 322.950 327.600 325.050 328.050 ;
        RECT 364.950 327.600 367.050 328.050 ;
        RECT 322.950 326.400 367.050 327.600 ;
        RECT 322.950 325.950 325.050 326.400 ;
        RECT 364.950 325.950 367.050 326.400 ;
        RECT 370.950 327.600 373.050 328.050 ;
        RECT 376.950 327.600 379.050 328.050 ;
        RECT 370.950 326.400 379.050 327.600 ;
        RECT 370.950 325.950 373.050 326.400 ;
        RECT 376.950 325.950 379.050 326.400 ;
        RECT 379.950 327.600 382.050 328.050 ;
        RECT 406.950 327.600 409.050 328.050 ;
        RECT 379.950 326.400 409.050 327.600 ;
        RECT 379.950 325.950 382.050 326.400 ;
        RECT 406.950 325.950 409.050 326.400 ;
        RECT 433.950 327.600 436.050 328.050 ;
        RECT 460.950 327.600 463.050 328.050 ;
        RECT 463.950 327.600 466.050 328.050 ;
        RECT 556.950 327.600 559.050 328.050 ;
        RECT 589.950 327.600 592.050 328.050 ;
        RECT 433.950 326.400 453.600 327.600 ;
        RECT 433.950 325.950 436.050 326.400 ;
        RECT 61.950 324.600 64.050 325.050 ;
        RECT 181.950 324.600 184.050 325.050 ;
        RECT 61.950 323.400 184.050 324.600 ;
        RECT 61.950 322.950 64.050 323.400 ;
        RECT 181.950 322.950 184.050 323.400 ;
        RECT 319.950 324.600 322.050 325.050 ;
        RECT 382.950 324.600 385.050 325.050 ;
        RECT 319.950 323.400 385.050 324.600 ;
        RECT 319.950 322.950 322.050 323.400 ;
        RECT 382.950 322.950 385.050 323.400 ;
        RECT 388.950 324.600 391.050 325.050 ;
        RECT 427.950 324.600 430.050 325.050 ;
        RECT 388.950 323.400 430.050 324.600 ;
        RECT 388.950 322.950 391.050 323.400 ;
        RECT 427.950 322.950 430.050 323.400 ;
        RECT 430.950 324.600 433.050 325.050 ;
        RECT 445.950 324.600 448.050 325.050 ;
        RECT 430.950 323.400 448.050 324.600 ;
        RECT 452.400 324.600 453.600 326.400 ;
        RECT 460.950 326.400 592.050 327.600 ;
        RECT 460.950 325.950 463.050 326.400 ;
        RECT 463.950 325.950 466.050 326.400 ;
        RECT 556.950 325.950 559.050 326.400 ;
        RECT 589.950 325.950 592.050 326.400 ;
        RECT 616.950 327.600 619.050 328.050 ;
        RECT 631.950 327.600 634.050 328.050 ;
        RECT 616.950 326.400 634.050 327.600 ;
        RECT 616.950 325.950 619.050 326.400 ;
        RECT 631.950 325.950 634.050 326.400 ;
        RECT 649.950 327.600 652.050 328.050 ;
        RECT 658.950 327.600 661.050 328.050 ;
        RECT 649.950 326.400 661.050 327.600 ;
        RECT 649.950 325.950 652.050 326.400 ;
        RECT 658.950 325.950 661.050 326.400 ;
        RECT 769.950 327.600 772.050 328.050 ;
        RECT 778.950 327.600 781.050 328.050 ;
        RECT 769.950 326.400 781.050 327.600 ;
        RECT 769.950 325.950 772.050 326.400 ;
        RECT 778.950 325.950 781.050 326.400 ;
        RECT 787.950 327.600 790.050 328.050 ;
        RECT 832.950 327.600 835.050 328.050 ;
        RECT 787.950 326.400 835.050 327.600 ;
        RECT 787.950 325.950 790.050 326.400 ;
        RECT 832.950 325.950 835.050 326.400 ;
        RECT 472.950 324.600 475.050 325.050 ;
        RECT 493.950 324.600 496.050 325.050 ;
        RECT 452.400 323.400 496.050 324.600 ;
        RECT 430.950 322.950 433.050 323.400 ;
        RECT 445.950 322.950 448.050 323.400 ;
        RECT 472.950 322.950 475.050 323.400 ;
        RECT 493.950 322.950 496.050 323.400 ;
        RECT 553.950 324.600 556.050 325.050 ;
        RECT 571.950 324.600 574.050 325.050 ;
        RECT 553.950 323.400 574.050 324.600 ;
        RECT 553.950 322.950 556.050 323.400 ;
        RECT 571.950 322.950 574.050 323.400 ;
        RECT 598.950 324.600 601.050 325.050 ;
        RECT 637.950 324.600 640.050 325.050 ;
        RECT 598.950 323.400 640.050 324.600 ;
        RECT 598.950 322.950 601.050 323.400 ;
        RECT 637.950 322.950 640.050 323.400 ;
        RECT 766.950 324.600 769.050 325.050 ;
        RECT 853.950 324.600 856.050 325.050 ;
        RECT 766.950 323.400 856.050 324.600 ;
        RECT 766.950 322.950 769.050 323.400 ;
        RECT 853.950 322.950 856.050 323.400 ;
        RECT 43.950 321.600 46.050 322.050 ;
        RECT 64.950 321.600 67.050 322.050 ;
        RECT 43.950 320.400 67.050 321.600 ;
        RECT 43.950 319.950 46.050 320.400 ;
        RECT 64.950 319.950 67.050 320.400 ;
        RECT 115.950 321.600 118.050 322.050 ;
        RECT 145.950 321.600 148.050 322.050 ;
        RECT 115.950 320.400 148.050 321.600 ;
        RECT 115.950 319.950 118.050 320.400 ;
        RECT 145.950 319.950 148.050 320.400 ;
        RECT 193.950 321.600 196.050 322.050 ;
        RECT 223.950 321.600 226.050 322.050 ;
        RECT 193.950 320.400 226.050 321.600 ;
        RECT 193.950 319.950 196.050 320.400 ;
        RECT 223.950 319.950 226.050 320.400 ;
        RECT 289.950 321.600 292.050 322.050 ;
        RECT 301.950 321.600 304.050 322.050 ;
        RECT 334.950 321.600 337.050 322.050 ;
        RECT 289.950 320.400 337.050 321.600 ;
        RECT 289.950 319.950 292.050 320.400 ;
        RECT 301.950 319.950 304.050 320.400 ;
        RECT 334.950 319.950 337.050 320.400 ;
        RECT 358.950 321.600 361.050 322.050 ;
        RECT 394.950 321.600 397.050 322.050 ;
        RECT 358.950 320.400 397.050 321.600 ;
        RECT 358.950 319.950 361.050 320.400 ;
        RECT 394.950 319.950 397.050 320.400 ;
        RECT 412.950 321.600 415.050 322.050 ;
        RECT 475.950 321.600 478.050 322.050 ;
        RECT 412.950 320.400 478.050 321.600 ;
        RECT 412.950 319.950 415.050 320.400 ;
        RECT 475.950 319.950 478.050 320.400 ;
        RECT 496.950 321.600 499.050 322.050 ;
        RECT 517.950 321.600 520.050 322.050 ;
        RECT 565.950 321.600 568.050 322.050 ;
        RECT 496.950 320.400 568.050 321.600 ;
        RECT 496.950 319.950 499.050 320.400 ;
        RECT 517.950 319.950 520.050 320.400 ;
        RECT 565.950 319.950 568.050 320.400 ;
        RECT 595.950 321.600 598.050 322.050 ;
        RECT 616.950 321.600 619.050 322.050 ;
        RECT 595.950 320.400 619.050 321.600 ;
        RECT 595.950 319.950 598.050 320.400 ;
        RECT 616.950 319.950 619.050 320.400 ;
        RECT 676.950 321.600 679.050 322.050 ;
        RECT 691.950 321.600 694.050 322.050 ;
        RECT 676.950 320.400 694.050 321.600 ;
        RECT 676.950 319.950 679.050 320.400 ;
        RECT 691.950 319.950 694.050 320.400 ;
        RECT 718.950 321.600 721.050 322.050 ;
        RECT 736.950 321.600 739.050 322.050 ;
        RECT 718.950 320.400 739.050 321.600 ;
        RECT 718.950 319.950 721.050 320.400 ;
        RECT 736.950 319.950 739.050 320.400 ;
        RECT 754.950 321.600 757.050 322.050 ;
        RECT 760.950 321.600 763.050 322.050 ;
        RECT 754.950 320.400 763.050 321.600 ;
        RECT 754.950 319.950 757.050 320.400 ;
        RECT 760.950 319.950 763.050 320.400 ;
        RECT 820.950 321.600 823.050 322.050 ;
        RECT 832.950 321.600 835.050 322.050 ;
        RECT 820.950 320.400 835.050 321.600 ;
        RECT 820.950 319.950 823.050 320.400 ;
        RECT 832.950 319.950 835.050 320.400 ;
        RECT 13.950 318.600 16.050 319.050 ;
        RECT 67.950 318.600 70.050 319.050 ;
        RECT 13.950 317.400 70.050 318.600 ;
        RECT 13.950 316.950 16.050 317.400 ;
        RECT 67.950 316.950 70.050 317.400 ;
        RECT 70.950 318.600 73.050 319.050 ;
        RECT 79.950 318.600 82.050 319.050 ;
        RECT 70.950 317.400 82.050 318.600 ;
        RECT 70.950 316.950 73.050 317.400 ;
        RECT 79.950 316.950 82.050 317.400 ;
        RECT 88.950 318.600 91.050 319.050 ;
        RECT 106.950 318.600 109.050 319.050 ;
        RECT 88.950 317.400 109.050 318.600 ;
        RECT 88.950 316.950 91.050 317.400 ;
        RECT 106.950 316.950 109.050 317.400 ;
        RECT 157.950 318.600 160.050 319.050 ;
        RECT 166.950 318.600 169.050 319.050 ;
        RECT 157.950 317.400 169.050 318.600 ;
        RECT 157.950 316.950 160.050 317.400 ;
        RECT 166.950 316.950 169.050 317.400 ;
        RECT 172.950 318.600 175.050 319.050 ;
        RECT 193.950 318.600 196.050 319.050 ;
        RECT 259.950 318.600 262.050 319.050 ;
        RECT 172.950 317.400 196.050 318.600 ;
        RECT 172.950 316.950 175.050 317.400 ;
        RECT 193.950 316.950 196.050 317.400 ;
        RECT 203.400 317.400 262.050 318.600 ;
        RECT 28.950 315.600 31.050 316.050 ;
        RECT 31.950 315.600 34.050 316.050 ;
        RECT 40.950 315.600 43.050 316.050 ;
        RECT 28.950 314.400 43.050 315.600 ;
        RECT 28.950 313.950 31.050 314.400 ;
        RECT 31.950 313.950 34.050 314.400 ;
        RECT 40.950 313.950 43.050 314.400 ;
        RECT 55.950 313.950 58.050 316.050 ;
        RECT 73.950 315.600 76.050 316.050 ;
        RECT 97.950 315.600 100.050 316.050 ;
        RECT 73.950 314.400 100.050 315.600 ;
        RECT 73.950 313.950 76.050 314.400 ;
        RECT 97.950 313.950 100.050 314.400 ;
        RECT 109.950 313.950 112.050 316.050 ;
        RECT 118.950 315.600 121.050 316.050 ;
        RECT 124.950 315.600 127.050 316.050 ;
        RECT 113.400 314.400 121.050 315.600 ;
        RECT 43.950 312.600 46.050 313.050 ;
        RECT 17.400 311.400 46.050 312.600 ;
        RECT 17.400 310.050 18.600 311.400 ;
        RECT 43.950 310.950 46.050 311.400 ;
        RECT 16.950 307.950 19.050 310.050 ;
        RECT 43.950 309.600 46.050 310.050 ;
        RECT 52.950 309.600 55.050 310.050 ;
        RECT 43.950 308.400 55.050 309.600 ;
        RECT 43.950 307.950 46.050 308.400 ;
        RECT 52.950 307.950 55.050 308.400 ;
        RECT 1.950 306.600 4.050 307.050 ;
        RECT 7.950 306.600 10.050 307.050 ;
        RECT 1.950 305.400 10.050 306.600 ;
        RECT 1.950 304.950 4.050 305.400 ;
        RECT 7.950 304.950 10.050 305.400 ;
        RECT 31.950 306.600 34.050 307.050 ;
        RECT 40.950 306.600 43.050 307.050 ;
        RECT 31.950 305.400 43.050 306.600 ;
        RECT 56.400 306.600 57.600 313.950 ;
        RECT 76.950 312.600 79.050 313.050 ;
        RECT 103.950 312.600 106.050 313.050 ;
        RECT 110.400 312.600 111.600 313.950 ;
        RECT 59.400 311.400 79.050 312.600 ;
        RECT 59.400 310.050 60.600 311.400 ;
        RECT 76.950 310.950 79.050 311.400 ;
        RECT 80.400 311.400 106.050 312.600 ;
        RECT 58.950 307.950 61.050 310.050 ;
        RECT 76.950 309.600 79.050 310.050 ;
        RECT 80.400 309.600 81.600 311.400 ;
        RECT 103.950 310.950 106.050 311.400 ;
        RECT 107.400 311.400 111.600 312.600 ;
        RECT 76.950 308.400 81.600 309.600 ;
        RECT 76.950 307.950 79.050 308.400 ;
        RECT 58.950 306.600 61.050 307.050 ;
        RECT 56.400 305.400 61.050 306.600 ;
        RECT 31.950 304.950 34.050 305.400 ;
        RECT 40.950 304.950 43.050 305.400 ;
        RECT 58.950 304.950 61.050 305.400 ;
        RECT 103.950 306.600 106.050 307.050 ;
        RECT 107.400 306.600 108.600 311.400 ;
        RECT 109.950 309.600 112.050 310.050 ;
        RECT 113.400 309.600 114.600 314.400 ;
        RECT 118.950 313.950 121.050 314.400 ;
        RECT 122.400 314.400 127.050 315.600 ;
        RECT 122.400 312.600 123.600 314.400 ;
        RECT 124.950 313.950 127.050 314.400 ;
        RECT 163.950 315.600 166.050 316.050 ;
        RECT 178.950 315.600 181.050 316.050 ;
        RECT 203.400 315.600 204.600 317.400 ;
        RECT 259.950 316.950 262.050 317.400 ;
        RECT 265.950 318.600 268.050 319.050 ;
        RECT 271.950 318.600 274.050 319.050 ;
        RECT 304.950 318.600 307.050 319.050 ;
        RECT 265.950 317.400 307.050 318.600 ;
        RECT 265.950 316.950 268.050 317.400 ;
        RECT 271.950 316.950 274.050 317.400 ;
        RECT 304.950 316.950 307.050 317.400 ;
        RECT 307.950 318.600 310.050 319.050 ;
        RECT 325.950 318.600 328.050 319.050 ;
        RECT 307.950 317.400 328.050 318.600 ;
        RECT 307.950 316.950 310.050 317.400 ;
        RECT 325.950 316.950 328.050 317.400 ;
        RECT 394.950 318.600 397.050 319.050 ;
        RECT 418.950 318.600 421.050 319.050 ;
        RECT 427.950 318.600 430.050 319.050 ;
        RECT 394.950 317.400 417.600 318.600 ;
        RECT 394.950 316.950 397.050 317.400 ;
        RECT 163.950 314.400 204.600 315.600 ;
        RECT 163.950 313.950 166.050 314.400 ;
        RECT 178.950 313.950 181.050 314.400 ;
        RECT 136.950 312.600 139.050 313.050 ;
        RECT 119.400 311.400 123.600 312.600 ;
        RECT 125.400 311.400 139.050 312.600 ;
        RECT 119.400 310.050 120.600 311.400 ;
        RECT 109.950 308.400 114.600 309.600 ;
        RECT 109.950 307.950 112.050 308.400 ;
        RECT 118.950 307.950 121.050 310.050 ;
        RECT 125.400 309.600 126.600 311.400 ;
        RECT 136.950 310.950 139.050 311.400 ;
        RECT 151.950 312.600 154.050 313.050 ;
        RECT 196.950 312.600 199.050 313.050 ;
        RECT 151.950 311.400 199.050 312.600 ;
        RECT 151.950 310.950 154.050 311.400 ;
        RECT 196.950 310.950 199.050 311.400 ;
        RECT 199.950 310.950 202.050 313.050 ;
        RECT 122.400 308.400 126.600 309.600 ;
        RECT 127.950 309.600 130.050 310.050 ;
        RECT 142.950 309.600 145.050 310.050 ;
        RECT 157.950 309.600 160.050 310.050 ;
        RECT 127.950 308.400 160.050 309.600 ;
        RECT 103.950 305.400 108.600 306.600 ;
        RECT 112.950 306.600 115.050 307.050 ;
        RECT 122.400 306.600 123.600 308.400 ;
        RECT 127.950 307.950 130.050 308.400 ;
        RECT 142.950 307.950 145.050 308.400 ;
        RECT 157.950 307.950 160.050 308.400 ;
        RECT 160.950 309.600 163.050 310.050 ;
        RECT 175.950 309.600 178.050 310.050 ;
        RECT 160.950 308.400 178.050 309.600 ;
        RECT 160.950 307.950 163.050 308.400 ;
        RECT 175.950 307.950 178.050 308.400 ;
        RECT 112.950 305.400 123.600 306.600 ;
        RECT 130.950 306.600 133.050 307.050 ;
        RECT 154.950 306.600 157.050 307.050 ;
        RECT 200.400 306.600 201.600 310.950 ;
        RECT 203.400 309.600 204.600 314.400 ;
        RECT 205.950 315.600 208.050 316.050 ;
        RECT 217.950 315.600 220.050 316.050 ;
        RECT 220.950 315.600 223.050 316.050 ;
        RECT 205.950 314.400 223.050 315.600 ;
        RECT 205.950 313.950 208.050 314.400 ;
        RECT 217.950 313.950 220.050 314.400 ;
        RECT 220.950 313.950 223.050 314.400 ;
        RECT 223.950 315.600 226.050 316.050 ;
        RECT 238.950 315.600 241.050 316.050 ;
        RECT 223.950 314.400 241.050 315.600 ;
        RECT 223.950 313.950 226.050 314.400 ;
        RECT 238.950 313.950 241.050 314.400 ;
        RECT 268.950 315.600 271.050 316.050 ;
        RECT 274.950 315.600 277.050 316.050 ;
        RECT 268.950 314.400 277.050 315.600 ;
        RECT 268.950 313.950 271.050 314.400 ;
        RECT 274.950 313.950 277.050 314.400 ;
        RECT 298.950 315.600 301.050 316.050 ;
        RECT 310.950 315.600 313.050 316.050 ;
        RECT 298.950 314.400 313.050 315.600 ;
        RECT 298.950 313.950 301.050 314.400 ;
        RECT 310.950 313.950 313.050 314.400 ;
        RECT 319.950 315.600 322.050 316.050 ;
        RECT 325.950 315.600 328.050 316.050 ;
        RECT 319.950 314.400 328.050 315.600 ;
        RECT 319.950 313.950 322.050 314.400 ;
        RECT 325.950 313.950 328.050 314.400 ;
        RECT 361.950 315.600 364.050 316.050 ;
        RECT 367.950 315.600 370.050 316.050 ;
        RECT 361.950 314.400 370.050 315.600 ;
        RECT 361.950 313.950 364.050 314.400 ;
        RECT 367.950 313.950 370.050 314.400 ;
        RECT 370.950 315.600 373.050 316.050 ;
        RECT 373.950 315.600 376.050 316.050 ;
        RECT 385.950 315.600 388.050 316.050 ;
        RECT 412.950 315.600 415.050 316.050 ;
        RECT 370.950 314.400 388.050 315.600 ;
        RECT 370.950 313.950 373.050 314.400 ;
        RECT 373.950 313.950 376.050 314.400 ;
        RECT 385.950 313.950 388.050 314.400 ;
        RECT 389.400 314.400 415.050 315.600 ;
        RECT 416.400 315.600 417.600 317.400 ;
        RECT 418.950 317.400 430.050 318.600 ;
        RECT 418.950 316.950 421.050 317.400 ;
        RECT 427.950 316.950 430.050 317.400 ;
        RECT 514.950 318.600 517.050 319.050 ;
        RECT 541.950 318.600 544.050 319.050 ;
        RECT 514.950 317.400 544.050 318.600 ;
        RECT 514.950 316.950 517.050 317.400 ;
        RECT 541.950 316.950 544.050 317.400 ;
        RECT 610.950 318.600 613.050 319.050 ;
        RECT 625.950 318.600 628.050 319.050 ;
        RECT 610.950 317.400 628.050 318.600 ;
        RECT 610.950 316.950 613.050 317.400 ;
        RECT 625.950 316.950 628.050 317.400 ;
        RECT 682.950 318.600 685.050 319.050 ;
        RECT 715.950 318.600 718.050 319.050 ;
        RECT 682.950 317.400 718.050 318.600 ;
        RECT 682.950 316.950 685.050 317.400 ;
        RECT 715.950 316.950 718.050 317.400 ;
        RECT 736.950 318.600 739.050 319.050 ;
        RECT 754.950 318.600 757.050 319.050 ;
        RECT 736.950 317.400 757.050 318.600 ;
        RECT 736.950 316.950 739.050 317.400 ;
        RECT 754.950 316.950 757.050 317.400 ;
        RECT 757.950 318.600 760.050 319.050 ;
        RECT 775.950 318.600 778.050 319.050 ;
        RECT 757.950 317.400 778.050 318.600 ;
        RECT 757.950 316.950 760.050 317.400 ;
        RECT 775.950 316.950 778.050 317.400 ;
        RECT 805.950 318.600 808.050 319.050 ;
        RECT 835.950 318.600 838.050 319.050 ;
        RECT 805.950 317.400 838.050 318.600 ;
        RECT 805.950 316.950 808.050 317.400 ;
        RECT 835.950 316.950 838.050 317.400 ;
        RECT 418.950 315.600 421.050 316.050 ;
        RECT 416.400 314.400 421.050 315.600 ;
        RECT 205.950 312.600 208.050 313.050 ;
        RECT 265.950 312.600 268.050 313.050 ;
        RECT 205.950 311.400 246.600 312.600 ;
        RECT 205.950 310.950 208.050 311.400 ;
        RECT 229.950 309.600 232.050 310.050 ;
        RECT 203.400 308.400 232.050 309.600 ;
        RECT 229.950 307.950 232.050 308.400 ;
        RECT 130.950 305.400 201.600 306.600 ;
        RECT 245.400 306.600 246.600 311.400 ;
        RECT 248.400 311.400 268.050 312.600 ;
        RECT 248.400 310.050 249.600 311.400 ;
        RECT 265.950 310.950 268.050 311.400 ;
        RECT 328.950 312.600 331.050 313.050 ;
        RECT 331.950 312.600 334.050 313.050 ;
        RECT 389.400 312.600 390.600 314.400 ;
        RECT 412.950 313.950 415.050 314.400 ;
        RECT 418.950 313.950 421.050 314.400 ;
        RECT 436.950 315.600 439.050 316.050 ;
        RECT 448.950 315.600 451.050 316.050 ;
        RECT 454.950 315.600 457.050 316.050 ;
        RECT 436.950 314.400 447.600 315.600 ;
        RECT 436.950 313.950 439.050 314.400 ;
        RECT 328.950 311.400 390.600 312.600 ;
        RECT 391.950 312.600 394.050 313.050 ;
        RECT 412.950 312.600 415.050 313.050 ;
        RECT 391.950 311.400 415.050 312.600 ;
        RECT 328.950 310.950 331.050 311.400 ;
        RECT 331.950 310.950 334.050 311.400 ;
        RECT 391.950 310.950 394.050 311.400 ;
        RECT 412.950 310.950 415.050 311.400 ;
        RECT 424.950 312.600 427.050 313.050 ;
        RECT 442.950 312.600 445.050 313.050 ;
        RECT 424.950 311.400 445.050 312.600 ;
        RECT 446.400 312.600 447.600 314.400 ;
        RECT 448.950 314.400 457.050 315.600 ;
        RECT 448.950 313.950 451.050 314.400 ;
        RECT 454.950 313.950 457.050 314.400 ;
        RECT 460.950 315.600 463.050 316.050 ;
        RECT 466.950 315.600 469.050 316.050 ;
        RECT 460.950 314.400 469.050 315.600 ;
        RECT 460.950 313.950 463.050 314.400 ;
        RECT 466.950 313.950 469.050 314.400 ;
        RECT 469.950 315.600 472.050 316.050 ;
        RECT 502.950 315.600 505.050 316.050 ;
        RECT 469.950 314.400 505.050 315.600 ;
        RECT 469.950 313.950 472.050 314.400 ;
        RECT 502.950 313.950 505.050 314.400 ;
        RECT 514.950 315.600 517.050 316.050 ;
        RECT 535.950 315.600 538.050 316.050 ;
        RECT 514.950 314.400 538.050 315.600 ;
        RECT 514.950 313.950 517.050 314.400 ;
        RECT 535.950 313.950 538.050 314.400 ;
        RECT 565.950 315.600 568.050 316.050 ;
        RECT 571.950 315.600 574.050 316.050 ;
        RECT 622.950 315.600 625.050 316.050 ;
        RECT 670.950 315.600 673.050 316.050 ;
        RECT 565.950 314.400 673.050 315.600 ;
        RECT 565.950 313.950 568.050 314.400 ;
        RECT 571.950 313.950 574.050 314.400 ;
        RECT 622.950 313.950 625.050 314.400 ;
        RECT 670.950 313.950 673.050 314.400 ;
        RECT 673.950 315.600 676.050 316.050 ;
        RECT 679.950 315.600 682.050 316.050 ;
        RECT 700.950 315.600 703.050 316.050 ;
        RECT 673.950 314.400 703.050 315.600 ;
        RECT 673.950 313.950 676.050 314.400 ;
        RECT 679.950 313.950 682.050 314.400 ;
        RECT 700.950 313.950 703.050 314.400 ;
        RECT 709.950 315.600 712.050 316.050 ;
        RECT 733.950 315.600 736.050 316.050 ;
        RECT 766.950 315.600 769.050 316.050 ;
        RECT 709.950 314.400 769.050 315.600 ;
        RECT 709.950 313.950 712.050 314.400 ;
        RECT 733.950 313.950 736.050 314.400 ;
        RECT 766.950 313.950 769.050 314.400 ;
        RECT 781.950 315.600 784.050 316.050 ;
        RECT 820.950 315.600 823.050 316.050 ;
        RECT 847.950 315.600 850.050 316.050 ;
        RECT 781.950 314.400 823.050 315.600 ;
        RECT 781.950 313.950 784.050 314.400 ;
        RECT 820.950 313.950 823.050 314.400 ;
        RECT 830.400 314.400 850.050 315.600 ;
        RECT 446.400 311.400 459.600 312.600 ;
        RECT 424.950 310.950 427.050 311.400 ;
        RECT 442.950 310.950 445.050 311.400 ;
        RECT 247.950 307.950 250.050 310.050 ;
        RECT 310.950 309.600 313.050 310.050 ;
        RECT 316.950 309.600 319.050 310.050 ;
        RECT 349.950 309.600 352.050 310.050 ;
        RECT 310.950 308.400 319.050 309.600 ;
        RECT 310.950 307.950 313.050 308.400 ;
        RECT 316.950 307.950 319.050 308.400 ;
        RECT 338.400 308.400 352.050 309.600 ;
        RECT 338.400 307.050 339.600 308.400 ;
        RECT 349.950 307.950 352.050 308.400 ;
        RECT 250.950 306.600 253.050 307.050 ;
        RECT 245.400 305.400 253.050 306.600 ;
        RECT 103.950 304.950 106.050 305.400 ;
        RECT 112.950 304.950 115.050 305.400 ;
        RECT 130.950 304.950 133.050 305.400 ;
        RECT 154.950 304.950 157.050 305.400 ;
        RECT 250.950 304.950 253.050 305.400 ;
        RECT 277.950 306.600 280.050 307.050 ;
        RECT 283.950 306.600 286.050 307.050 ;
        RECT 277.950 305.400 286.050 306.600 ;
        RECT 277.950 304.950 280.050 305.400 ;
        RECT 283.950 304.950 286.050 305.400 ;
        RECT 337.950 304.950 340.050 307.050 ;
        RECT 367.950 306.600 370.050 307.050 ;
        RECT 385.950 306.600 388.050 307.050 ;
        RECT 367.950 305.400 388.050 306.600 ;
        RECT 413.400 306.600 414.600 310.950 ;
        RECT 415.950 309.600 418.050 310.050 ;
        RECT 427.950 309.600 430.050 310.050 ;
        RECT 415.950 308.400 430.050 309.600 ;
        RECT 443.400 309.600 444.600 310.950 ;
        RECT 458.400 310.050 459.600 311.400 ;
        RECT 466.950 310.950 469.050 313.050 ;
        RECT 472.950 312.600 475.050 313.050 ;
        RECT 508.950 312.600 511.050 313.050 ;
        RECT 523.950 312.600 526.050 313.050 ;
        RECT 568.950 312.600 571.050 313.050 ;
        RECT 595.950 312.600 598.050 313.050 ;
        RECT 472.950 311.400 480.600 312.600 ;
        RECT 472.950 310.950 475.050 311.400 ;
        RECT 454.950 309.600 457.050 310.050 ;
        RECT 443.400 308.400 457.050 309.600 ;
        RECT 415.950 307.950 418.050 308.400 ;
        RECT 427.950 307.950 430.050 308.400 ;
        RECT 454.950 307.950 457.050 308.400 ;
        RECT 457.950 307.950 460.050 310.050 ;
        RECT 467.400 307.050 468.600 310.950 ;
        RECT 415.950 306.600 418.050 307.050 ;
        RECT 413.400 305.400 418.050 306.600 ;
        RECT 367.950 304.950 370.050 305.400 ;
        RECT 385.950 304.950 388.050 305.400 ;
        RECT 415.950 304.950 418.050 305.400 ;
        RECT 427.950 306.600 430.050 307.050 ;
        RECT 433.950 306.600 436.050 307.050 ;
        RECT 427.950 305.400 436.050 306.600 ;
        RECT 427.950 304.950 430.050 305.400 ;
        RECT 433.950 304.950 436.050 305.400 ;
        RECT 466.950 304.950 469.050 307.050 ;
        RECT 479.400 306.600 480.600 311.400 ;
        RECT 508.950 311.400 522.600 312.600 ;
        RECT 508.950 310.950 511.050 311.400 ;
        RECT 521.400 310.050 522.600 311.400 ;
        RECT 523.950 311.400 598.050 312.600 ;
        RECT 523.950 310.950 526.050 311.400 ;
        RECT 568.950 310.950 571.050 311.400 ;
        RECT 595.950 310.950 598.050 311.400 ;
        RECT 619.950 312.600 622.050 313.050 ;
        RECT 646.950 312.600 649.050 313.050 ;
        RECT 667.950 312.600 670.050 313.050 ;
        RECT 619.950 311.400 670.050 312.600 ;
        RECT 619.950 310.950 622.050 311.400 ;
        RECT 646.950 310.950 649.050 311.400 ;
        RECT 667.950 310.950 670.050 311.400 ;
        RECT 685.950 312.600 688.050 313.050 ;
        RECT 697.950 312.600 700.050 313.050 ;
        RECT 685.950 311.400 700.050 312.600 ;
        RECT 685.950 310.950 688.050 311.400 ;
        RECT 697.950 310.950 700.050 311.400 ;
        RECT 724.950 312.600 727.050 313.050 ;
        RECT 748.950 312.600 751.050 313.050 ;
        RECT 724.950 311.400 751.050 312.600 ;
        RECT 724.950 310.950 727.050 311.400 ;
        RECT 748.950 310.950 751.050 311.400 ;
        RECT 772.950 312.600 775.050 313.050 ;
        RECT 778.950 312.600 781.050 313.050 ;
        RECT 772.950 311.400 781.050 312.600 ;
        RECT 772.950 310.950 775.050 311.400 ;
        RECT 778.950 310.950 781.050 311.400 ;
        RECT 787.950 312.600 790.050 313.050 ;
        RECT 796.950 312.600 799.050 313.050 ;
        RECT 787.950 311.400 799.050 312.600 ;
        RECT 787.950 310.950 790.050 311.400 ;
        RECT 796.950 310.950 799.050 311.400 ;
        RECT 811.950 312.600 814.050 313.050 ;
        RECT 811.950 311.400 819.600 312.600 ;
        RECT 811.950 310.950 814.050 311.400 ;
        RECT 508.950 309.600 511.050 310.050 ;
        RECT 517.950 309.600 520.050 310.050 ;
        RECT 508.950 308.400 520.050 309.600 ;
        RECT 508.950 307.950 511.050 308.400 ;
        RECT 517.950 307.950 520.050 308.400 ;
        RECT 520.950 307.950 523.050 310.050 ;
        RECT 535.950 309.600 538.050 310.050 ;
        RECT 538.950 309.600 541.050 310.050 ;
        RECT 565.950 309.600 568.050 310.050 ;
        RECT 535.950 308.400 568.050 309.600 ;
        RECT 535.950 307.950 538.050 308.400 ;
        RECT 538.950 307.950 541.050 308.400 ;
        RECT 565.950 307.950 568.050 308.400 ;
        RECT 628.950 309.600 631.050 310.050 ;
        RECT 634.950 309.600 637.050 310.050 ;
        RECT 628.950 308.400 637.050 309.600 ;
        RECT 628.950 307.950 631.050 308.400 ;
        RECT 634.950 307.950 637.050 308.400 ;
        RECT 655.950 309.600 658.050 310.050 ;
        RECT 712.950 309.600 715.050 310.050 ;
        RECT 760.950 309.600 763.050 310.050 ;
        RECT 784.950 309.600 787.050 310.050 ;
        RECT 655.950 308.400 711.600 309.600 ;
        RECT 655.950 307.950 658.050 308.400 ;
        RECT 484.950 306.600 487.050 307.050 ;
        RECT 479.400 305.400 487.050 306.600 ;
        RECT 484.950 304.950 487.050 305.400 ;
        RECT 505.950 306.600 508.050 307.050 ;
        RECT 562.950 306.600 565.050 307.050 ;
        RECT 505.950 305.400 565.050 306.600 ;
        RECT 505.950 304.950 508.050 305.400 ;
        RECT 562.950 304.950 565.050 305.400 ;
        RECT 583.950 306.600 586.050 307.050 ;
        RECT 601.950 306.600 604.050 307.050 ;
        RECT 583.950 305.400 604.050 306.600 ;
        RECT 583.950 304.950 586.050 305.400 ;
        RECT 601.950 304.950 604.050 305.400 ;
        RECT 604.950 306.600 607.050 307.050 ;
        RECT 613.950 306.600 616.050 307.050 ;
        RECT 604.950 305.400 616.050 306.600 ;
        RECT 604.950 304.950 607.050 305.400 ;
        RECT 613.950 304.950 616.050 305.400 ;
        RECT 619.950 306.600 622.050 307.050 ;
        RECT 625.950 306.600 628.050 307.050 ;
        RECT 673.950 306.600 676.050 307.050 ;
        RECT 619.950 305.400 676.050 306.600 ;
        RECT 619.950 304.950 622.050 305.400 ;
        RECT 625.950 304.950 628.050 305.400 ;
        RECT 673.950 304.950 676.050 305.400 ;
        RECT 697.950 306.600 700.050 307.050 ;
        RECT 706.950 306.600 709.050 307.050 ;
        RECT 697.950 305.400 709.050 306.600 ;
        RECT 710.400 306.600 711.600 308.400 ;
        RECT 712.950 308.400 787.050 309.600 ;
        RECT 712.950 307.950 715.050 308.400 ;
        RECT 760.950 307.950 763.050 308.400 ;
        RECT 784.950 307.950 787.050 308.400 ;
        RECT 790.950 307.950 793.050 310.050 ;
        RECT 802.950 309.600 805.050 310.050 ;
        RECT 814.950 309.600 817.050 310.050 ;
        RECT 802.950 308.400 817.050 309.600 ;
        RECT 802.950 307.950 805.050 308.400 ;
        RECT 814.950 307.950 817.050 308.400 ;
        RECT 751.950 306.600 754.050 307.050 ;
        RECT 710.400 305.400 754.050 306.600 ;
        RECT 697.950 304.950 700.050 305.400 ;
        RECT 706.950 304.950 709.050 305.400 ;
        RECT 751.950 304.950 754.050 305.400 ;
        RECT 757.950 306.600 760.050 307.050 ;
        RECT 766.950 306.600 769.050 307.050 ;
        RECT 757.950 305.400 769.050 306.600 ;
        RECT 791.400 306.600 792.600 307.950 ;
        RECT 799.950 306.600 802.050 307.050 ;
        RECT 791.400 305.400 802.050 306.600 ;
        RECT 818.400 306.600 819.600 311.400 ;
        RECT 823.950 309.600 826.050 310.050 ;
        RECT 830.400 309.600 831.600 314.400 ;
        RECT 847.950 313.950 850.050 314.400 ;
        RECT 832.950 310.950 835.050 313.050 ;
        RECT 847.950 310.950 850.050 313.050 ;
        RECT 823.950 308.400 831.600 309.600 ;
        RECT 823.950 307.950 826.050 308.400 ;
        RECT 833.400 307.050 834.600 310.950 ;
        RECT 820.950 306.600 823.050 307.050 ;
        RECT 818.400 305.400 823.050 306.600 ;
        RECT 757.950 304.950 760.050 305.400 ;
        RECT 766.950 304.950 769.050 305.400 ;
        RECT 799.950 304.950 802.050 305.400 ;
        RECT 820.950 304.950 823.050 305.400 ;
        RECT 832.950 304.950 835.050 307.050 ;
        RECT 848.400 306.600 849.600 310.950 ;
        RECT 853.950 306.600 856.050 307.050 ;
        RECT 848.400 305.400 856.050 306.600 ;
        RECT 853.950 304.950 856.050 305.400 ;
        RECT 139.950 303.600 142.050 304.050 ;
        RECT 145.950 303.600 148.050 304.050 ;
        RECT 139.950 302.400 148.050 303.600 ;
        RECT 139.950 301.950 142.050 302.400 ;
        RECT 145.950 301.950 148.050 302.400 ;
        RECT 148.950 303.600 151.050 304.050 ;
        RECT 163.950 303.600 166.050 304.050 ;
        RECT 148.950 302.400 166.050 303.600 ;
        RECT 148.950 301.950 151.050 302.400 ;
        RECT 163.950 301.950 166.050 302.400 ;
        RECT 187.950 303.600 190.050 304.050 ;
        RECT 202.950 303.600 205.050 304.050 ;
        RECT 223.950 303.600 226.050 304.050 ;
        RECT 187.950 302.400 226.050 303.600 ;
        RECT 187.950 301.950 190.050 302.400 ;
        RECT 202.950 301.950 205.050 302.400 ;
        RECT 223.950 301.950 226.050 302.400 ;
        RECT 304.950 303.600 307.050 304.050 ;
        RECT 313.950 303.600 316.050 304.050 ;
        RECT 304.950 302.400 316.050 303.600 ;
        RECT 304.950 301.950 307.050 302.400 ;
        RECT 313.950 301.950 316.050 302.400 ;
        RECT 325.950 303.600 328.050 304.050 ;
        RECT 352.950 303.600 355.050 304.050 ;
        RECT 325.950 302.400 355.050 303.600 ;
        RECT 325.950 301.950 328.050 302.400 ;
        RECT 352.950 301.950 355.050 302.400 ;
        RECT 361.950 303.600 364.050 304.050 ;
        RECT 367.950 303.600 370.050 304.050 ;
        RECT 361.950 302.400 370.050 303.600 ;
        RECT 361.950 301.950 364.050 302.400 ;
        RECT 367.950 301.950 370.050 302.400 ;
        RECT 373.950 303.600 376.050 304.050 ;
        RECT 379.950 303.600 382.050 304.050 ;
        RECT 385.950 303.600 388.050 304.050 ;
        RECT 373.950 302.400 388.050 303.600 ;
        RECT 373.950 301.950 376.050 302.400 ;
        RECT 379.950 301.950 382.050 302.400 ;
        RECT 385.950 301.950 388.050 302.400 ;
        RECT 394.950 303.600 397.050 304.050 ;
        RECT 421.950 303.600 424.050 304.050 ;
        RECT 394.950 302.400 424.050 303.600 ;
        RECT 394.950 301.950 397.050 302.400 ;
        RECT 421.950 301.950 424.050 302.400 ;
        RECT 478.950 303.600 481.050 304.050 ;
        RECT 508.950 303.600 511.050 304.050 ;
        RECT 478.950 302.400 511.050 303.600 ;
        RECT 478.950 301.950 481.050 302.400 ;
        RECT 508.950 301.950 511.050 302.400 ;
        RECT 583.950 303.600 586.050 304.050 ;
        RECT 598.950 303.600 601.050 304.050 ;
        RECT 583.950 302.400 601.050 303.600 ;
        RECT 583.950 301.950 586.050 302.400 ;
        RECT 598.950 301.950 601.050 302.400 ;
        RECT 640.950 303.600 643.050 304.050 ;
        RECT 694.950 303.600 697.050 304.050 ;
        RECT 640.950 302.400 697.050 303.600 ;
        RECT 640.950 301.950 643.050 302.400 ;
        RECT 694.950 301.950 697.050 302.400 ;
        RECT 778.950 303.600 781.050 304.050 ;
        RECT 850.950 303.600 853.050 304.050 ;
        RECT 778.950 302.400 853.050 303.600 ;
        RECT 778.950 301.950 781.050 302.400 ;
        RECT 850.950 301.950 853.050 302.400 ;
        RECT 37.950 300.600 40.050 301.050 ;
        RECT 61.950 300.600 64.050 301.050 ;
        RECT 37.950 299.400 64.050 300.600 ;
        RECT 37.950 298.950 40.050 299.400 ;
        RECT 61.950 298.950 64.050 299.400 ;
        RECT 124.950 300.600 127.050 301.050 ;
        RECT 133.950 300.600 136.050 301.050 ;
        RECT 172.950 300.600 175.050 301.050 ;
        RECT 124.950 299.400 175.050 300.600 ;
        RECT 124.950 298.950 127.050 299.400 ;
        RECT 133.950 298.950 136.050 299.400 ;
        RECT 172.950 298.950 175.050 299.400 ;
        RECT 190.950 300.600 193.050 301.050 ;
        RECT 205.950 300.600 208.050 301.050 ;
        RECT 190.950 299.400 208.050 300.600 ;
        RECT 190.950 298.950 193.050 299.400 ;
        RECT 205.950 298.950 208.050 299.400 ;
        RECT 256.950 300.600 259.050 301.050 ;
        RECT 319.950 300.600 322.050 301.050 ;
        RECT 256.950 299.400 322.050 300.600 ;
        RECT 256.950 298.950 259.050 299.400 ;
        RECT 319.950 298.950 322.050 299.400 ;
        RECT 322.950 300.600 325.050 301.050 ;
        RECT 346.950 300.600 349.050 301.050 ;
        RECT 322.950 299.400 349.050 300.600 ;
        RECT 322.950 298.950 325.050 299.400 ;
        RECT 346.950 298.950 349.050 299.400 ;
        RECT 364.950 300.600 367.050 301.050 ;
        RECT 400.950 300.600 403.050 301.050 ;
        RECT 364.950 299.400 403.050 300.600 ;
        RECT 364.950 298.950 367.050 299.400 ;
        RECT 400.950 298.950 403.050 299.400 ;
        RECT 418.950 300.600 421.050 301.050 ;
        RECT 445.950 300.600 448.050 301.050 ;
        RECT 418.950 299.400 448.050 300.600 ;
        RECT 418.950 298.950 421.050 299.400 ;
        RECT 445.950 298.950 448.050 299.400 ;
        RECT 490.950 300.600 493.050 301.050 ;
        RECT 535.950 300.600 538.050 301.050 ;
        RECT 490.950 299.400 538.050 300.600 ;
        RECT 490.950 298.950 493.050 299.400 ;
        RECT 535.950 298.950 538.050 299.400 ;
        RECT 649.950 300.600 652.050 301.050 ;
        RECT 712.950 300.600 715.050 301.050 ;
        RECT 649.950 299.400 715.050 300.600 ;
        RECT 649.950 298.950 652.050 299.400 ;
        RECT 712.950 298.950 715.050 299.400 ;
        RECT 739.950 300.600 742.050 301.050 ;
        RECT 808.950 300.600 811.050 301.050 ;
        RECT 811.950 300.600 814.050 301.050 ;
        RECT 739.950 299.400 814.050 300.600 ;
        RECT 739.950 298.950 742.050 299.400 ;
        RECT 808.950 298.950 811.050 299.400 ;
        RECT 811.950 298.950 814.050 299.400 ;
        RECT 826.950 300.600 829.050 301.050 ;
        RECT 838.950 300.600 841.050 301.050 ;
        RECT 826.950 299.400 841.050 300.600 ;
        RECT 826.950 298.950 829.050 299.400 ;
        RECT 838.950 298.950 841.050 299.400 ;
        RECT 46.950 297.600 49.050 298.050 ;
        RECT 73.950 297.600 76.050 298.050 ;
        RECT 46.950 296.400 76.050 297.600 ;
        RECT 46.950 295.950 49.050 296.400 ;
        RECT 73.950 295.950 76.050 296.400 ;
        RECT 160.950 297.600 163.050 298.050 ;
        RECT 202.950 297.600 205.050 298.050 ;
        RECT 208.950 297.600 211.050 298.050 ;
        RECT 160.950 296.400 211.050 297.600 ;
        RECT 160.950 295.950 163.050 296.400 ;
        RECT 202.950 295.950 205.050 296.400 ;
        RECT 208.950 295.950 211.050 296.400 ;
        RECT 304.950 297.600 307.050 298.050 ;
        RECT 388.950 297.600 391.050 298.050 ;
        RECT 304.950 296.400 391.050 297.600 ;
        RECT 304.950 295.950 307.050 296.400 ;
        RECT 388.950 295.950 391.050 296.400 ;
        RECT 421.950 297.600 424.050 298.050 ;
        RECT 439.950 297.600 442.050 298.050 ;
        RECT 472.950 297.600 475.050 298.050 ;
        RECT 421.950 296.400 475.050 297.600 ;
        RECT 421.950 295.950 424.050 296.400 ;
        RECT 439.950 295.950 442.050 296.400 ;
        RECT 472.950 295.950 475.050 296.400 ;
        RECT 511.950 297.600 514.050 298.050 ;
        RECT 601.950 297.600 604.050 298.050 ;
        RECT 511.950 296.400 604.050 297.600 ;
        RECT 511.950 295.950 514.050 296.400 ;
        RECT 601.950 295.950 604.050 296.400 ;
        RECT 637.950 297.600 640.050 298.050 ;
        RECT 661.950 297.600 664.050 298.050 ;
        RECT 637.950 296.400 664.050 297.600 ;
        RECT 637.950 295.950 640.050 296.400 ;
        RECT 661.950 295.950 664.050 296.400 ;
        RECT 727.950 297.600 730.050 298.050 ;
        RECT 787.950 297.600 790.050 298.050 ;
        RECT 727.950 296.400 790.050 297.600 ;
        RECT 727.950 295.950 730.050 296.400 ;
        RECT 787.950 295.950 790.050 296.400 ;
        RECT 823.950 297.600 826.050 298.050 ;
        RECT 832.950 297.600 835.050 298.050 ;
        RECT 823.950 296.400 835.050 297.600 ;
        RECT 823.950 295.950 826.050 296.400 ;
        RECT 832.950 295.950 835.050 296.400 ;
        RECT 34.950 294.600 37.050 295.050 ;
        RECT 67.950 294.600 70.050 295.050 ;
        RECT 34.950 293.400 70.050 294.600 ;
        RECT 34.950 292.950 37.050 293.400 ;
        RECT 67.950 292.950 70.050 293.400 ;
        RECT 70.950 294.600 73.050 295.050 ;
        RECT 139.950 294.600 142.050 295.050 ;
        RECT 70.950 293.400 142.050 294.600 ;
        RECT 70.950 292.950 73.050 293.400 ;
        RECT 139.950 292.950 142.050 293.400 ;
        RECT 163.950 294.600 166.050 295.050 ;
        RECT 175.950 294.600 178.050 295.050 ;
        RECT 163.950 293.400 178.050 294.600 ;
        RECT 163.950 292.950 166.050 293.400 ;
        RECT 175.950 292.950 178.050 293.400 ;
        RECT 214.950 294.600 217.050 295.050 ;
        RECT 235.950 294.600 238.050 295.050 ;
        RECT 262.950 294.600 265.050 295.050 ;
        RECT 412.950 294.600 415.050 295.050 ;
        RECT 214.950 293.400 415.050 294.600 ;
        RECT 214.950 292.950 217.050 293.400 ;
        RECT 235.950 292.950 238.050 293.400 ;
        RECT 262.950 292.950 265.050 293.400 ;
        RECT 412.950 292.950 415.050 293.400 ;
        RECT 415.950 294.600 418.050 295.050 ;
        RECT 520.950 294.600 523.050 295.050 ;
        RECT 682.950 294.600 685.050 295.050 ;
        RECT 415.950 293.400 501.600 294.600 ;
        RECT 415.950 292.950 418.050 293.400 ;
        RECT 10.950 291.600 13.050 292.050 ;
        RECT 70.950 291.600 73.050 292.050 ;
        RECT 10.950 290.400 73.050 291.600 ;
        RECT 10.950 289.950 13.050 290.400 ;
        RECT 70.950 289.950 73.050 290.400 ;
        RECT 181.950 291.600 184.050 292.050 ;
        RECT 247.950 291.600 250.050 292.050 ;
        RECT 367.950 291.600 370.050 292.050 ;
        RECT 181.950 290.400 370.050 291.600 ;
        RECT 181.950 289.950 184.050 290.400 ;
        RECT 247.950 289.950 250.050 290.400 ;
        RECT 367.950 289.950 370.050 290.400 ;
        RECT 406.950 291.600 409.050 292.050 ;
        RECT 457.950 291.600 460.050 292.050 ;
        RECT 406.950 290.400 460.050 291.600 ;
        RECT 406.950 289.950 409.050 290.400 ;
        RECT 457.950 289.950 460.050 290.400 ;
        RECT 475.950 291.600 478.050 292.050 ;
        RECT 496.950 291.600 499.050 292.050 ;
        RECT 475.950 290.400 499.050 291.600 ;
        RECT 500.400 291.600 501.600 293.400 ;
        RECT 520.950 293.400 685.050 294.600 ;
        RECT 520.950 292.950 523.050 293.400 ;
        RECT 682.950 292.950 685.050 293.400 ;
        RECT 688.950 294.600 691.050 295.050 ;
        RECT 724.950 294.600 727.050 295.050 ;
        RECT 688.950 293.400 727.050 294.600 ;
        RECT 688.950 292.950 691.050 293.400 ;
        RECT 724.950 292.950 727.050 293.400 ;
        RECT 763.950 294.600 766.050 295.050 ;
        RECT 838.950 294.600 841.050 295.050 ;
        RECT 763.950 293.400 841.050 294.600 ;
        RECT 763.950 292.950 766.050 293.400 ;
        RECT 838.950 292.950 841.050 293.400 ;
        RECT 532.950 291.600 535.050 292.050 ;
        RECT 500.400 290.400 535.050 291.600 ;
        RECT 475.950 289.950 478.050 290.400 ;
        RECT 496.950 289.950 499.050 290.400 ;
        RECT 532.950 289.950 535.050 290.400 ;
        RECT 580.950 291.600 583.050 292.050 ;
        RECT 607.950 291.600 610.050 292.050 ;
        RECT 580.950 290.400 610.050 291.600 ;
        RECT 580.950 289.950 583.050 290.400 ;
        RECT 607.950 289.950 610.050 290.400 ;
        RECT 709.950 291.600 712.050 292.050 ;
        RECT 820.950 291.600 823.050 292.050 ;
        RECT 853.950 291.600 856.050 292.050 ;
        RECT 709.950 290.400 856.050 291.600 ;
        RECT 709.950 289.950 712.050 290.400 ;
        RECT 820.950 289.950 823.050 290.400 ;
        RECT 853.950 289.950 856.050 290.400 ;
        RECT 1.950 288.600 4.050 289.050 ;
        RECT 49.950 288.600 52.050 289.050 ;
        RECT 1.950 287.400 52.050 288.600 ;
        RECT 1.950 286.950 4.050 287.400 ;
        RECT 49.950 286.950 52.050 287.400 ;
        RECT 82.950 288.600 85.050 289.050 ;
        RECT 169.950 288.600 172.050 289.050 ;
        RECT 82.950 287.400 172.050 288.600 ;
        RECT 82.950 286.950 85.050 287.400 ;
        RECT 169.950 286.950 172.050 287.400 ;
        RECT 175.950 288.600 178.050 289.050 ;
        RECT 193.950 288.600 196.050 289.050 ;
        RECT 232.950 288.600 235.050 289.050 ;
        RECT 175.950 287.400 235.050 288.600 ;
        RECT 175.950 286.950 178.050 287.400 ;
        RECT 193.950 286.950 196.050 287.400 ;
        RECT 232.950 286.950 235.050 287.400 ;
        RECT 253.950 288.600 256.050 289.050 ;
        RECT 469.950 288.600 472.050 289.050 ;
        RECT 253.950 287.400 472.050 288.600 ;
        RECT 253.950 286.950 256.050 287.400 ;
        RECT 469.950 286.950 472.050 287.400 ;
        RECT 472.950 288.600 475.050 289.050 ;
        RECT 547.950 288.600 550.050 289.050 ;
        RECT 598.950 288.600 601.050 289.050 ;
        RECT 472.950 287.400 495.600 288.600 ;
        RECT 472.950 286.950 475.050 287.400 ;
        RECT 4.950 285.600 7.050 286.050 ;
        RECT 13.950 285.600 16.050 286.050 ;
        RECT 253.950 285.600 256.050 286.050 ;
        RECT 4.950 284.400 256.050 285.600 ;
        RECT 4.950 283.950 7.050 284.400 ;
        RECT 13.950 283.950 16.050 284.400 ;
        RECT 253.950 283.950 256.050 284.400 ;
        RECT 277.950 285.600 280.050 286.050 ;
        RECT 337.950 285.600 340.050 286.050 ;
        RECT 358.950 285.600 361.050 286.050 ;
        RECT 277.950 284.400 361.050 285.600 ;
        RECT 277.950 283.950 280.050 284.400 ;
        RECT 337.950 283.950 340.050 284.400 ;
        RECT 358.950 283.950 361.050 284.400 ;
        RECT 415.950 285.600 418.050 286.050 ;
        RECT 448.950 285.600 451.050 286.050 ;
        RECT 484.950 285.600 487.050 286.050 ;
        RECT 415.950 284.400 487.050 285.600 ;
        RECT 494.400 285.600 495.600 287.400 ;
        RECT 547.950 287.400 601.050 288.600 ;
        RECT 547.950 286.950 550.050 287.400 ;
        RECT 598.950 286.950 601.050 287.400 ;
        RECT 601.950 288.600 604.050 289.050 ;
        RECT 700.950 288.600 703.050 289.050 ;
        RECT 601.950 287.400 703.050 288.600 ;
        RECT 601.950 286.950 604.050 287.400 ;
        RECT 700.950 286.950 703.050 287.400 ;
        RECT 781.950 288.600 784.050 289.050 ;
        RECT 817.950 288.600 820.050 289.050 ;
        RECT 781.950 287.400 820.050 288.600 ;
        RECT 781.950 286.950 784.050 287.400 ;
        RECT 817.950 286.950 820.050 287.400 ;
        RECT 559.950 285.600 562.050 286.050 ;
        RECT 494.400 284.400 562.050 285.600 ;
        RECT 415.950 283.950 418.050 284.400 ;
        RECT 448.950 283.950 451.050 284.400 ;
        RECT 484.950 283.950 487.050 284.400 ;
        RECT 559.950 283.950 562.050 284.400 ;
        RECT 574.950 285.600 577.050 286.050 ;
        RECT 697.950 285.600 700.050 286.050 ;
        RECT 574.950 284.400 700.050 285.600 ;
        RECT 574.950 283.950 577.050 284.400 ;
        RECT 697.950 283.950 700.050 284.400 ;
        RECT 733.950 285.600 736.050 286.050 ;
        RECT 760.950 285.600 763.050 286.050 ;
        RECT 733.950 284.400 763.050 285.600 ;
        RECT 733.950 283.950 736.050 284.400 ;
        RECT 760.950 283.950 763.050 284.400 ;
        RECT 796.950 285.600 799.050 286.050 ;
        RECT 805.950 285.600 808.050 286.050 ;
        RECT 796.950 284.400 808.050 285.600 ;
        RECT 796.950 283.950 799.050 284.400 ;
        RECT 805.950 283.950 808.050 284.400 ;
        RECT 829.950 285.600 832.050 286.050 ;
        RECT 835.950 285.600 838.050 286.050 ;
        RECT 829.950 284.400 838.050 285.600 ;
        RECT 829.950 283.950 832.050 284.400 ;
        RECT 835.950 283.950 838.050 284.400 ;
        RECT 79.950 282.600 82.050 283.050 ;
        RECT 100.950 282.600 103.050 283.050 ;
        RECT 79.950 281.400 103.050 282.600 ;
        RECT 79.950 280.950 82.050 281.400 ;
        RECT 100.950 280.950 103.050 281.400 ;
        RECT 112.950 282.600 115.050 283.050 ;
        RECT 121.950 282.600 124.050 283.050 ;
        RECT 178.950 282.600 181.050 283.050 ;
        RECT 112.950 281.400 181.050 282.600 ;
        RECT 112.950 280.950 115.050 281.400 ;
        RECT 121.950 280.950 124.050 281.400 ;
        RECT 178.950 280.950 181.050 281.400 ;
        RECT 199.950 282.600 202.050 283.050 ;
        RECT 229.950 282.600 232.050 283.050 ;
        RECT 199.950 281.400 232.050 282.600 ;
        RECT 199.950 280.950 202.050 281.400 ;
        RECT 229.950 280.950 232.050 281.400 ;
        RECT 232.950 282.600 235.050 283.050 ;
        RECT 277.950 282.600 280.050 283.050 ;
        RECT 232.950 281.400 280.050 282.600 ;
        RECT 232.950 280.950 235.050 281.400 ;
        RECT 277.950 280.950 280.050 281.400 ;
        RECT 301.950 282.600 304.050 283.050 ;
        RECT 325.950 282.600 328.050 283.050 ;
        RECT 301.950 281.400 328.050 282.600 ;
        RECT 301.950 280.950 304.050 281.400 ;
        RECT 325.950 280.950 328.050 281.400 ;
        RECT 355.950 282.600 358.050 283.050 ;
        RECT 391.950 282.600 394.050 283.050 ;
        RECT 448.950 282.600 451.050 283.050 ;
        RECT 355.950 281.400 451.050 282.600 ;
        RECT 355.950 280.950 358.050 281.400 ;
        RECT 391.950 280.950 394.050 281.400 ;
        RECT 448.950 280.950 451.050 281.400 ;
        RECT 451.950 282.600 454.050 283.050 ;
        RECT 490.950 282.600 493.050 283.050 ;
        RECT 451.950 281.400 493.050 282.600 ;
        RECT 451.950 280.950 454.050 281.400 ;
        RECT 490.950 280.950 493.050 281.400 ;
        RECT 499.950 282.600 502.050 283.050 ;
        RECT 574.950 282.600 577.050 283.050 ;
        RECT 499.950 281.400 577.050 282.600 ;
        RECT 499.950 280.950 502.050 281.400 ;
        RECT 574.950 280.950 577.050 281.400 ;
        RECT 577.950 282.600 580.050 283.050 ;
        RECT 640.950 282.600 643.050 283.050 ;
        RECT 577.950 281.400 643.050 282.600 ;
        RECT 577.950 280.950 580.050 281.400 ;
        RECT 640.950 280.950 643.050 281.400 ;
        RECT 691.950 282.600 694.050 283.050 ;
        RECT 739.950 282.600 742.050 283.050 ;
        RECT 691.950 281.400 742.050 282.600 ;
        RECT 691.950 280.950 694.050 281.400 ;
        RECT 739.950 280.950 742.050 281.400 ;
        RECT 742.950 282.600 745.050 283.050 ;
        RECT 775.950 282.600 778.050 283.050 ;
        RECT 742.950 281.400 778.050 282.600 ;
        RECT 742.950 280.950 745.050 281.400 ;
        RECT 775.950 280.950 778.050 281.400 ;
        RECT 166.950 279.600 169.050 280.050 ;
        RECT 187.950 279.600 190.050 280.050 ;
        RECT 292.950 279.600 295.050 280.050 ;
        RECT 298.950 279.600 301.050 280.050 ;
        RECT 379.950 279.600 382.050 280.050 ;
        RECT 166.950 278.400 279.600 279.600 ;
        RECT 166.950 277.950 169.050 278.400 ;
        RECT 187.950 277.950 190.050 278.400 ;
        RECT 61.950 276.600 64.050 277.050 ;
        RECT 88.950 276.600 91.050 277.050 ;
        RECT 94.950 276.600 97.050 277.050 ;
        RECT 61.950 275.400 84.600 276.600 ;
        RECT 61.950 274.950 64.050 275.400 ;
        RECT 83.400 274.050 84.600 275.400 ;
        RECT 88.950 275.400 97.050 276.600 ;
        RECT 88.950 274.950 91.050 275.400 ;
        RECT 94.950 274.950 97.050 275.400 ;
        RECT 112.950 276.600 115.050 277.050 ;
        RECT 130.950 276.600 133.050 277.050 ;
        RECT 112.950 275.400 133.050 276.600 ;
        RECT 112.950 274.950 115.050 275.400 ;
        RECT 130.950 274.950 133.050 275.400 ;
        RECT 166.950 276.600 169.050 277.050 ;
        RECT 175.950 276.600 178.050 277.050 ;
        RECT 166.950 275.400 178.050 276.600 ;
        RECT 166.950 274.950 169.050 275.400 ;
        RECT 175.950 274.950 178.050 275.400 ;
        RECT 196.950 276.600 199.050 277.050 ;
        RECT 220.950 276.600 223.050 277.050 ;
        RECT 196.950 275.400 223.050 276.600 ;
        RECT 196.950 274.950 199.050 275.400 ;
        RECT 220.950 274.950 223.050 275.400 ;
        RECT 253.950 276.600 256.050 277.050 ;
        RECT 274.950 276.600 277.050 277.050 ;
        RECT 253.950 275.400 277.050 276.600 ;
        RECT 253.950 274.950 256.050 275.400 ;
        RECT 274.950 274.950 277.050 275.400 ;
        RECT 278.400 276.600 279.600 278.400 ;
        RECT 292.950 278.400 382.050 279.600 ;
        RECT 292.950 277.950 295.050 278.400 ;
        RECT 298.950 277.950 301.050 278.400 ;
        RECT 379.950 277.950 382.050 278.400 ;
        RECT 385.950 279.600 388.050 280.050 ;
        RECT 424.950 279.600 427.050 280.050 ;
        RECT 460.950 279.600 463.050 280.050 ;
        RECT 385.950 278.400 427.050 279.600 ;
        RECT 385.950 277.950 388.050 278.400 ;
        RECT 424.950 277.950 427.050 278.400 ;
        RECT 431.400 278.400 463.050 279.600 ;
        RECT 340.950 276.600 343.050 277.050 ;
        RECT 346.950 276.600 349.050 277.050 ;
        RECT 278.400 275.400 349.050 276.600 ;
        RECT 76.950 273.600 79.050 274.050 ;
        RECT 76.950 272.400 81.600 273.600 ;
        RECT 76.950 271.950 79.050 272.400 ;
        RECT 25.950 270.600 28.050 271.050 ;
        RECT 52.950 270.600 55.050 271.050 ;
        RECT 25.950 269.400 55.050 270.600 ;
        RECT 25.950 268.950 28.050 269.400 ;
        RECT 52.950 268.950 55.050 269.400 ;
        RECT 67.950 268.950 70.050 271.050 ;
        RECT 25.950 267.600 28.050 268.050 ;
        RECT 68.400 267.600 69.600 268.950 ;
        RECT 80.400 268.050 81.600 272.400 ;
        RECT 82.950 271.950 85.050 274.050 ;
        RECT 118.950 273.600 121.050 274.050 ;
        RECT 133.950 273.600 136.050 274.050 ;
        RECT 154.950 273.600 157.050 274.050 ;
        RECT 118.950 272.400 136.050 273.600 ;
        RECT 118.950 271.950 121.050 272.400 ;
        RECT 133.950 271.950 136.050 272.400 ;
        RECT 143.400 272.400 157.050 273.600 ;
        RECT 143.400 271.050 144.600 272.400 ;
        RECT 154.950 271.950 157.050 272.400 ;
        RECT 160.950 273.600 163.050 274.050 ;
        RECT 181.950 273.600 184.050 274.050 ;
        RECT 160.950 272.400 184.050 273.600 ;
        RECT 160.950 271.950 163.050 272.400 ;
        RECT 181.950 271.950 184.050 272.400 ;
        RECT 214.950 273.600 217.050 274.050 ;
        RECT 214.950 272.400 261.600 273.600 ;
        RECT 214.950 271.950 217.050 272.400 ;
        RECT 85.950 270.600 88.050 271.050 ;
        RECT 91.950 270.600 94.050 271.050 ;
        RECT 112.950 270.600 115.050 271.050 ;
        RECT 85.950 269.400 115.050 270.600 ;
        RECT 85.950 268.950 88.050 269.400 ;
        RECT 91.950 268.950 94.050 269.400 ;
        RECT 112.950 268.950 115.050 269.400 ;
        RECT 121.950 270.600 124.050 271.050 ;
        RECT 121.950 269.400 135.600 270.600 ;
        RECT 121.950 268.950 124.050 269.400 ;
        RECT 25.950 266.400 69.600 267.600 ;
        RECT 25.950 265.950 28.050 266.400 ;
        RECT 79.950 265.950 82.050 268.050 ;
        RECT 115.950 267.600 118.050 268.050 ;
        RECT 127.950 267.600 130.050 268.050 ;
        RECT 115.950 266.400 130.050 267.600 ;
        RECT 134.400 267.600 135.600 269.400 ;
        RECT 142.950 268.950 145.050 271.050 ;
        RECT 145.950 270.600 148.050 271.050 ;
        RECT 196.950 270.600 199.050 271.050 ;
        RECT 145.950 269.400 199.050 270.600 ;
        RECT 145.950 268.950 148.050 269.400 ;
        RECT 196.950 268.950 199.050 269.400 ;
        RECT 211.950 268.950 214.050 271.050 ;
        RECT 217.950 268.950 220.050 271.050 ;
        RECT 220.950 270.600 223.050 271.050 ;
        RECT 226.950 270.600 229.050 271.050 ;
        RECT 238.950 270.600 241.050 271.050 ;
        RECT 220.950 269.400 225.600 270.600 ;
        RECT 220.950 268.950 223.050 269.400 ;
        RECT 148.950 267.600 151.050 268.050 ;
        RECT 134.400 266.400 151.050 267.600 ;
        RECT 115.950 265.950 118.050 266.400 ;
        RECT 127.950 265.950 130.050 266.400 ;
        RECT 148.950 265.950 151.050 266.400 ;
        RECT 157.950 267.600 160.050 268.050 ;
        RECT 163.950 267.600 166.050 268.050 ;
        RECT 157.950 266.400 166.050 267.600 ;
        RECT 157.950 265.950 160.050 266.400 ;
        RECT 163.950 265.950 166.050 266.400 ;
        RECT 184.950 267.600 187.050 268.050 ;
        RECT 196.950 267.600 199.050 268.050 ;
        RECT 184.950 266.400 199.050 267.600 ;
        RECT 184.950 265.950 187.050 266.400 ;
        RECT 196.950 265.950 199.050 266.400 ;
        RECT 7.950 264.600 10.050 265.050 ;
        RECT 82.950 264.600 85.050 265.050 ;
        RECT 7.950 263.400 85.050 264.600 ;
        RECT 7.950 262.950 10.050 263.400 ;
        RECT 82.950 262.950 85.050 263.400 ;
        RECT 100.950 264.600 103.050 265.050 ;
        RECT 115.950 264.600 118.050 265.050 ;
        RECT 100.950 263.400 118.050 264.600 ;
        RECT 100.950 262.950 103.050 263.400 ;
        RECT 115.950 262.950 118.050 263.400 ;
        RECT 121.950 264.600 124.050 265.050 ;
        RECT 139.950 264.600 142.050 265.050 ;
        RECT 121.950 263.400 142.050 264.600 ;
        RECT 121.950 262.950 124.050 263.400 ;
        RECT 139.950 262.950 142.050 263.400 ;
        RECT 142.950 264.600 145.050 265.050 ;
        RECT 190.950 264.600 193.050 265.050 ;
        RECT 142.950 263.400 193.050 264.600 ;
        RECT 212.400 264.600 213.600 268.950 ;
        RECT 218.400 267.600 219.600 268.950 ;
        RECT 220.950 267.600 223.050 268.050 ;
        RECT 218.400 266.400 223.050 267.600 ;
        RECT 224.400 267.600 225.600 269.400 ;
        RECT 226.950 269.400 241.050 270.600 ;
        RECT 260.400 270.600 261.600 272.400 ;
        RECT 265.950 271.950 268.050 274.050 ;
        RECT 271.950 273.600 274.050 274.050 ;
        RECT 278.400 273.600 279.600 275.400 ;
        RECT 340.950 274.950 343.050 275.400 ;
        RECT 346.950 274.950 349.050 275.400 ;
        RECT 349.950 276.600 352.050 277.050 ;
        RECT 418.950 276.600 421.050 277.050 ;
        RECT 427.950 276.600 430.050 277.050 ;
        RECT 349.950 275.400 421.050 276.600 ;
        RECT 349.950 274.950 352.050 275.400 ;
        RECT 418.950 274.950 421.050 275.400 ;
        RECT 422.400 275.400 430.050 276.600 ;
        RECT 286.950 273.600 289.050 274.050 ;
        RECT 271.950 272.400 279.600 273.600 ;
        RECT 281.400 272.400 289.050 273.600 ;
        RECT 271.950 271.950 274.050 272.400 ;
        RECT 266.400 270.600 267.600 271.950 ;
        RECT 274.950 270.600 277.050 271.050 ;
        RECT 281.400 270.600 282.600 272.400 ;
        RECT 286.950 271.950 289.050 272.400 ;
        RECT 322.950 273.600 325.050 274.050 ;
        RECT 358.950 273.600 361.050 274.050 ;
        RECT 364.950 273.600 367.050 274.050 ;
        RECT 400.950 273.600 403.050 274.050 ;
        RECT 322.950 272.400 348.600 273.600 ;
        RECT 322.950 271.950 325.050 272.400 ;
        RECT 260.400 269.400 264.600 270.600 ;
        RECT 266.400 269.400 277.050 270.600 ;
        RECT 226.950 268.950 229.050 269.400 ;
        RECT 238.950 268.950 241.050 269.400 ;
        RECT 232.950 267.600 235.050 268.050 ;
        RECT 224.400 266.400 235.050 267.600 ;
        RECT 263.400 267.600 264.600 269.400 ;
        RECT 274.950 268.950 277.050 269.400 ;
        RECT 278.400 269.400 282.600 270.600 ;
        RECT 283.950 270.600 286.050 271.050 ;
        RECT 289.950 270.600 292.050 271.050 ;
        RECT 301.950 270.600 304.050 271.050 ;
        RECT 283.950 269.400 292.050 270.600 ;
        RECT 271.950 267.600 274.050 268.050 ;
        RECT 263.400 266.400 274.050 267.600 ;
        RECT 220.950 265.950 223.050 266.400 ;
        RECT 232.950 265.950 235.050 266.400 ;
        RECT 271.950 265.950 274.050 266.400 ;
        RECT 274.950 267.600 277.050 268.050 ;
        RECT 278.400 267.600 279.600 269.400 ;
        RECT 283.950 268.950 286.050 269.400 ;
        RECT 289.950 268.950 292.050 269.400 ;
        RECT 293.400 269.400 304.050 270.600 ;
        RECT 274.950 266.400 279.600 267.600 ;
        RECT 280.950 267.600 283.050 268.050 ;
        RECT 286.950 267.600 289.050 268.050 ;
        RECT 280.950 266.400 289.050 267.600 ;
        RECT 274.950 265.950 277.050 266.400 ;
        RECT 280.950 265.950 283.050 266.400 ;
        RECT 286.950 265.950 289.050 266.400 ;
        RECT 289.950 267.600 292.050 268.050 ;
        RECT 293.400 267.600 294.600 269.400 ;
        RECT 301.950 268.950 304.050 269.400 ;
        RECT 310.950 270.600 313.050 271.050 ;
        RECT 343.950 270.600 346.050 271.050 ;
        RECT 310.950 269.400 346.050 270.600 ;
        RECT 347.400 270.600 348.600 272.400 ;
        RECT 358.950 272.400 367.050 273.600 ;
        RECT 358.950 271.950 361.050 272.400 ;
        RECT 364.950 271.950 367.050 272.400 ;
        RECT 374.400 272.400 403.050 273.600 ;
        RECT 355.950 270.600 358.050 271.050 ;
        RECT 367.950 270.600 370.050 271.050 ;
        RECT 347.400 269.400 351.600 270.600 ;
        RECT 310.950 268.950 313.050 269.400 ;
        RECT 343.950 268.950 346.050 269.400 ;
        RECT 289.950 266.400 294.600 267.600 ;
        RECT 310.950 267.600 313.050 268.050 ;
        RECT 316.950 267.600 319.050 268.050 ;
        RECT 310.950 266.400 319.050 267.600 ;
        RECT 289.950 265.950 292.050 266.400 ;
        RECT 310.950 265.950 313.050 266.400 ;
        RECT 316.950 265.950 319.050 266.400 ;
        RECT 334.950 267.600 337.050 268.050 ;
        RECT 346.950 267.600 349.050 268.050 ;
        RECT 334.950 266.400 349.050 267.600 ;
        RECT 350.400 267.600 351.600 269.400 ;
        RECT 355.950 269.400 370.050 270.600 ;
        RECT 355.950 268.950 358.050 269.400 ;
        RECT 367.950 268.950 370.050 269.400 ;
        RECT 370.950 267.600 373.050 268.050 ;
        RECT 350.400 266.400 373.050 267.600 ;
        RECT 334.950 265.950 337.050 266.400 ;
        RECT 346.950 265.950 349.050 266.400 ;
        RECT 370.950 265.950 373.050 266.400 ;
        RECT 229.950 264.600 232.050 265.050 ;
        RECT 212.400 263.400 232.050 264.600 ;
        RECT 142.950 262.950 145.050 263.400 ;
        RECT 190.950 262.950 193.050 263.400 ;
        RECT 229.950 262.950 232.050 263.400 ;
        RECT 235.950 264.600 238.050 265.050 ;
        RECT 307.950 264.600 310.050 265.050 ;
        RECT 235.950 263.400 310.050 264.600 ;
        RECT 235.950 262.950 238.050 263.400 ;
        RECT 307.950 262.950 310.050 263.400 ;
        RECT 358.950 264.600 361.050 265.050 ;
        RECT 364.950 264.600 367.050 265.050 ;
        RECT 358.950 263.400 367.050 264.600 ;
        RECT 374.400 264.600 375.600 272.400 ;
        RECT 400.950 271.950 403.050 272.400 ;
        RECT 415.950 273.600 418.050 274.050 ;
        RECT 415.950 272.400 420.600 273.600 ;
        RECT 415.950 271.950 418.050 272.400 ;
        RECT 376.950 270.600 379.050 271.050 ;
        RECT 385.950 270.600 388.050 271.050 ;
        RECT 376.950 269.400 388.050 270.600 ;
        RECT 376.950 268.950 379.050 269.400 ;
        RECT 385.950 268.950 388.050 269.400 ;
        RECT 388.950 268.950 391.050 271.050 ;
        RECT 406.950 270.600 409.050 271.050 ;
        RECT 415.950 270.600 418.050 271.050 ;
        RECT 406.950 269.400 418.050 270.600 ;
        RECT 406.950 268.950 409.050 269.400 ;
        RECT 415.950 268.950 418.050 269.400 ;
        RECT 385.950 264.600 388.050 265.050 ;
        RECT 374.400 263.400 388.050 264.600 ;
        RECT 389.400 264.600 390.600 268.950 ;
        RECT 419.400 268.050 420.600 272.400 ;
        RECT 397.950 267.600 400.050 268.050 ;
        RECT 397.950 266.400 405.600 267.600 ;
        RECT 397.950 265.950 400.050 266.400 ;
        RECT 404.400 265.050 405.600 266.400 ;
        RECT 418.950 265.950 421.050 268.050 ;
        RECT 394.950 264.600 397.050 265.050 ;
        RECT 389.400 263.400 397.050 264.600 ;
        RECT 358.950 262.950 361.050 263.400 ;
        RECT 364.950 262.950 367.050 263.400 ;
        RECT 385.950 262.950 388.050 263.400 ;
        RECT 394.950 262.950 397.050 263.400 ;
        RECT 403.950 262.950 406.050 265.050 ;
        RECT 422.400 264.600 423.600 275.400 ;
        RECT 427.950 274.950 430.050 275.400 ;
        RECT 431.400 274.050 432.600 278.400 ;
        RECT 460.950 277.950 463.050 278.400 ;
        RECT 595.950 279.600 598.050 280.050 ;
        RECT 616.950 279.600 619.050 280.050 ;
        RECT 595.950 278.400 619.050 279.600 ;
        RECT 595.950 277.950 598.050 278.400 ;
        RECT 616.950 277.950 619.050 278.400 ;
        RECT 643.950 279.600 646.050 280.050 ;
        RECT 652.950 279.600 655.050 280.050 ;
        RECT 643.950 278.400 655.050 279.600 ;
        RECT 643.950 277.950 646.050 278.400 ;
        RECT 652.950 277.950 655.050 278.400 ;
        RECT 715.950 279.600 718.050 280.050 ;
        RECT 733.950 279.600 736.050 280.050 ;
        RECT 715.950 278.400 736.050 279.600 ;
        RECT 715.950 277.950 718.050 278.400 ;
        RECT 733.950 277.950 736.050 278.400 ;
        RECT 757.950 279.600 760.050 280.050 ;
        RECT 775.950 279.600 778.050 280.050 ;
        RECT 757.950 278.400 778.050 279.600 ;
        RECT 757.950 277.950 760.050 278.400 ;
        RECT 775.950 277.950 778.050 278.400 ;
        RECT 445.950 276.600 448.050 277.050 ;
        RECT 454.950 276.600 457.050 277.050 ;
        RECT 445.950 275.400 457.050 276.600 ;
        RECT 445.950 274.950 448.050 275.400 ;
        RECT 454.950 274.950 457.050 275.400 ;
        RECT 469.950 276.600 472.050 277.050 ;
        RECT 469.950 275.400 477.600 276.600 ;
        RECT 469.950 274.950 472.050 275.400 ;
        RECT 424.950 273.600 427.050 274.050 ;
        RECT 424.950 272.400 429.600 273.600 ;
        RECT 424.950 271.950 427.050 272.400 ;
        RECT 428.400 270.600 429.600 272.400 ;
        RECT 430.950 271.950 433.050 274.050 ;
        RECT 451.950 273.600 454.050 274.050 ;
        RECT 472.950 273.600 475.050 274.050 ;
        RECT 451.950 272.400 475.050 273.600 ;
        RECT 451.950 271.950 454.050 272.400 ;
        RECT 472.950 271.950 475.050 272.400 ;
        RECT 439.950 270.600 442.050 271.050 ;
        RECT 469.950 270.600 472.050 271.050 ;
        RECT 428.400 269.400 438.600 270.600 ;
        RECT 437.400 267.600 438.600 269.400 ;
        RECT 439.950 269.400 472.050 270.600 ;
        RECT 439.950 268.950 442.050 269.400 ;
        RECT 469.950 268.950 472.050 269.400 ;
        RECT 445.950 267.600 448.050 268.050 ;
        RECT 437.400 266.400 448.050 267.600 ;
        RECT 445.950 265.950 448.050 266.400 ;
        RECT 451.950 267.600 454.050 268.050 ;
        RECT 457.950 267.600 460.050 268.050 ;
        RECT 451.950 266.400 460.050 267.600 ;
        RECT 451.950 265.950 454.050 266.400 ;
        RECT 457.950 265.950 460.050 266.400 ;
        RECT 463.950 267.600 466.050 268.050 ;
        RECT 472.950 267.600 475.050 268.050 ;
        RECT 463.950 266.400 475.050 267.600 ;
        RECT 476.400 267.600 477.600 275.400 ;
        RECT 484.950 274.950 487.050 277.050 ;
        RECT 496.950 276.600 499.050 277.050 ;
        RECT 541.950 276.600 544.050 277.050 ;
        RECT 496.950 275.400 544.050 276.600 ;
        RECT 496.950 274.950 499.050 275.400 ;
        RECT 541.950 274.950 544.050 275.400 ;
        RECT 568.950 276.600 571.050 277.050 ;
        RECT 613.950 276.600 616.050 277.050 ;
        RECT 568.950 275.400 616.050 276.600 ;
        RECT 568.950 274.950 571.050 275.400 ;
        RECT 613.950 274.950 616.050 275.400 ;
        RECT 634.950 276.600 637.050 277.050 ;
        RECT 646.950 276.600 649.050 277.050 ;
        RECT 634.950 275.400 649.050 276.600 ;
        RECT 634.950 274.950 637.050 275.400 ;
        RECT 646.950 274.950 649.050 275.400 ;
        RECT 658.950 276.600 661.050 277.050 ;
        RECT 664.950 276.600 667.050 277.050 ;
        RECT 658.950 275.400 667.050 276.600 ;
        RECT 658.950 274.950 661.050 275.400 ;
        RECT 664.950 274.950 667.050 275.400 ;
        RECT 667.950 276.600 670.050 277.050 ;
        RECT 706.950 276.600 709.050 277.050 ;
        RECT 667.950 275.400 709.050 276.600 ;
        RECT 667.950 274.950 670.050 275.400 ;
        RECT 706.950 274.950 709.050 275.400 ;
        RECT 739.950 276.600 742.050 277.050 ;
        RECT 745.950 276.600 748.050 277.050 ;
        RECT 754.950 276.600 757.050 277.050 ;
        RECT 739.950 275.400 744.600 276.600 ;
        RECT 739.950 274.950 742.050 275.400 ;
        RECT 481.950 273.600 484.050 274.050 ;
        RECT 485.400 273.600 486.600 274.950 ;
        RECT 493.950 273.600 496.050 274.050 ;
        RECT 502.950 273.600 505.050 274.050 ;
        RECT 481.950 272.400 492.600 273.600 ;
        RECT 481.950 271.950 484.050 272.400 ;
        RECT 491.400 270.600 492.600 272.400 ;
        RECT 493.950 272.400 505.050 273.600 ;
        RECT 493.950 271.950 496.050 272.400 ;
        RECT 502.950 271.950 505.050 272.400 ;
        RECT 514.950 273.600 517.050 274.050 ;
        RECT 529.950 273.600 532.050 274.050 ;
        RECT 514.950 272.400 532.050 273.600 ;
        RECT 514.950 271.950 517.050 272.400 ;
        RECT 529.950 271.950 532.050 272.400 ;
        RECT 547.950 273.600 550.050 274.050 ;
        RECT 553.950 273.600 556.050 274.050 ;
        RECT 547.950 272.400 556.050 273.600 ;
        RECT 547.950 271.950 550.050 272.400 ;
        RECT 553.950 271.950 556.050 272.400 ;
        RECT 556.950 273.600 559.050 274.050 ;
        RECT 598.950 273.600 601.050 274.050 ;
        RECT 610.950 273.600 613.050 274.050 ;
        RECT 628.950 273.600 631.050 274.050 ;
        RECT 640.950 273.600 643.050 274.050 ;
        RECT 670.950 273.600 673.050 274.050 ;
        RECT 688.950 273.600 691.050 274.050 ;
        RECT 556.950 272.400 561.600 273.600 ;
        RECT 556.950 271.950 559.050 272.400 ;
        RECT 491.400 269.400 519.600 270.600 ;
        RECT 518.400 268.050 519.600 269.400 ;
        RECT 526.950 268.950 529.050 271.050 ;
        RECT 538.950 270.600 541.050 271.050 ;
        RECT 530.400 269.400 541.050 270.600 ;
        RECT 481.950 267.600 484.050 268.050 ;
        RECT 476.400 266.400 484.050 267.600 ;
        RECT 463.950 265.950 466.050 266.400 ;
        RECT 472.950 265.950 475.050 266.400 ;
        RECT 481.950 265.950 484.050 266.400 ;
        RECT 505.950 267.600 508.050 268.050 ;
        RECT 511.950 267.600 514.050 268.050 ;
        RECT 505.950 266.400 514.050 267.600 ;
        RECT 505.950 265.950 508.050 266.400 ;
        RECT 511.950 265.950 514.050 266.400 ;
        RECT 517.950 265.950 520.050 268.050 ;
        RECT 457.950 264.600 460.050 265.050 ;
        RECT 422.400 263.400 460.050 264.600 ;
        RECT 457.950 262.950 460.050 263.400 ;
        RECT 466.950 264.600 469.050 265.050 ;
        RECT 484.950 264.600 487.050 265.050 ;
        RECT 466.950 263.400 487.050 264.600 ;
        RECT 466.950 262.950 469.050 263.400 ;
        RECT 484.950 262.950 487.050 263.400 ;
        RECT 499.950 264.600 502.050 265.050 ;
        RECT 508.950 264.600 511.050 265.050 ;
        RECT 520.950 264.600 523.050 265.050 ;
        RECT 527.400 264.600 528.600 268.950 ;
        RECT 530.400 268.050 531.600 269.400 ;
        RECT 538.950 268.950 541.050 269.400 ;
        RECT 541.950 268.950 544.050 271.050 ;
        RECT 553.950 268.950 556.050 271.050 ;
        RECT 560.400 270.600 561.600 272.400 ;
        RECT 598.950 272.400 603.600 273.600 ;
        RECT 598.950 271.950 601.050 272.400 ;
        RECT 602.400 271.050 603.600 272.400 ;
        RECT 610.950 272.400 639.600 273.600 ;
        RECT 610.950 271.950 613.050 272.400 ;
        RECT 628.950 271.950 631.050 272.400 ;
        RECT 586.950 270.600 589.050 271.050 ;
        RECT 595.950 270.600 598.050 271.050 ;
        RECT 560.400 269.400 564.600 270.600 ;
        RECT 529.950 265.950 532.050 268.050 ;
        RECT 499.950 263.400 511.050 264.600 ;
        RECT 518.400 263.400 528.600 264.600 ;
        RECT 529.950 264.600 532.050 265.050 ;
        RECT 542.400 264.600 543.600 268.950 ;
        RECT 554.400 267.600 555.600 268.950 ;
        RECT 563.400 268.050 564.600 269.400 ;
        RECT 586.950 269.400 598.050 270.600 ;
        RECT 586.950 268.950 589.050 269.400 ;
        RECT 595.950 268.950 598.050 269.400 ;
        RECT 601.950 268.950 604.050 271.050 ;
        RECT 638.400 270.600 639.600 272.400 ;
        RECT 640.950 272.400 691.050 273.600 ;
        RECT 640.950 271.950 643.050 272.400 ;
        RECT 670.950 271.950 673.050 272.400 ;
        RECT 688.950 271.950 691.050 272.400 ;
        RECT 703.950 273.600 706.050 274.050 ;
        RECT 718.950 273.600 721.050 274.050 ;
        RECT 703.950 272.400 721.050 273.600 ;
        RECT 703.950 271.950 706.050 272.400 ;
        RECT 718.950 271.950 721.050 272.400 ;
        RECT 727.950 273.600 730.050 274.050 ;
        RECT 736.950 273.600 739.050 274.050 ;
        RECT 727.950 272.400 739.050 273.600 ;
        RECT 727.950 271.950 730.050 272.400 ;
        RECT 736.950 271.950 739.050 272.400 ;
        RECT 688.950 270.600 691.050 271.050 ;
        RECT 700.950 270.600 703.050 271.050 ;
        RECT 638.400 269.400 687.600 270.600 ;
        RECT 554.400 266.400 558.600 267.600 ;
        RECT 553.950 264.600 556.050 265.050 ;
        RECT 529.950 263.400 556.050 264.600 ;
        RECT 557.400 264.600 558.600 266.400 ;
        RECT 562.950 265.950 565.050 268.050 ;
        RECT 577.950 267.600 580.050 268.050 ;
        RECT 583.950 267.600 586.050 268.050 ;
        RECT 598.950 267.600 601.050 268.050 ;
        RECT 643.950 267.600 646.050 268.050 ;
        RECT 577.950 266.400 597.600 267.600 ;
        RECT 577.950 265.950 580.050 266.400 ;
        RECT 583.950 265.950 586.050 266.400 ;
        RECT 559.950 264.600 562.050 265.050 ;
        RECT 557.400 263.400 562.050 264.600 ;
        RECT 499.950 262.950 502.050 263.400 ;
        RECT 508.950 262.950 511.050 263.400 ;
        RECT 520.950 262.950 523.050 263.400 ;
        RECT 529.950 262.950 532.050 263.400 ;
        RECT 553.950 262.950 556.050 263.400 ;
        RECT 559.950 262.950 562.050 263.400 ;
        RECT 565.950 264.600 568.050 265.050 ;
        RECT 592.950 264.600 595.050 265.050 ;
        RECT 565.950 263.400 595.050 264.600 ;
        RECT 565.950 262.950 568.050 263.400 ;
        RECT 592.950 262.950 595.050 263.400 ;
        RECT 64.950 261.600 67.050 262.050 ;
        RECT 151.950 261.600 154.050 262.050 ;
        RECT 64.950 260.400 154.050 261.600 ;
        RECT 64.950 259.950 67.050 260.400 ;
        RECT 151.950 259.950 154.050 260.400 ;
        RECT 154.950 261.600 157.050 262.050 ;
        RECT 175.950 261.600 178.050 262.050 ;
        RECT 154.950 260.400 178.050 261.600 ;
        RECT 154.950 259.950 157.050 260.400 ;
        RECT 175.950 259.950 178.050 260.400 ;
        RECT 253.950 261.600 256.050 262.050 ;
        RECT 280.950 261.600 283.050 262.050 ;
        RECT 253.950 260.400 283.050 261.600 ;
        RECT 253.950 259.950 256.050 260.400 ;
        RECT 280.950 259.950 283.050 260.400 ;
        RECT 301.950 261.600 304.050 262.050 ;
        RECT 307.950 261.600 310.050 262.050 ;
        RECT 301.950 260.400 310.050 261.600 ;
        RECT 301.950 259.950 304.050 260.400 ;
        RECT 307.950 259.950 310.050 260.400 ;
        RECT 352.950 261.600 355.050 262.050 ;
        RECT 370.950 261.600 373.050 262.050 ;
        RECT 352.950 260.400 373.050 261.600 ;
        RECT 352.950 259.950 355.050 260.400 ;
        RECT 370.950 259.950 373.050 260.400 ;
        RECT 379.950 261.600 382.050 262.050 ;
        RECT 409.950 261.600 412.050 262.050 ;
        RECT 379.950 260.400 412.050 261.600 ;
        RECT 379.950 259.950 382.050 260.400 ;
        RECT 409.950 259.950 412.050 260.400 ;
        RECT 412.950 261.600 415.050 262.050 ;
        RECT 550.950 261.600 553.050 262.050 ;
        RECT 412.950 260.400 553.050 261.600 ;
        RECT 412.950 259.950 415.050 260.400 ;
        RECT 550.950 259.950 553.050 260.400 ;
        RECT 556.950 261.600 559.050 262.050 ;
        RECT 571.950 261.600 574.050 262.050 ;
        RECT 589.950 261.600 592.050 262.050 ;
        RECT 556.950 260.400 592.050 261.600 ;
        RECT 596.400 261.600 597.600 266.400 ;
        RECT 598.950 266.400 646.050 267.600 ;
        RECT 598.950 265.950 601.050 266.400 ;
        RECT 643.950 265.950 646.050 266.400 ;
        RECT 649.950 267.600 652.050 268.050 ;
        RECT 661.950 267.600 664.050 268.050 ;
        RECT 649.950 266.400 664.050 267.600 ;
        RECT 649.950 265.950 652.050 266.400 ;
        RECT 661.950 265.950 664.050 266.400 ;
        RECT 670.950 267.600 673.050 268.050 ;
        RECT 686.400 267.600 687.600 269.400 ;
        RECT 688.950 269.400 703.050 270.600 ;
        RECT 688.950 268.950 691.050 269.400 ;
        RECT 700.950 268.950 703.050 269.400 ;
        RECT 743.400 268.050 744.600 275.400 ;
        RECT 745.950 275.400 757.050 276.600 ;
        RECT 745.950 274.950 748.050 275.400 ;
        RECT 754.950 274.950 757.050 275.400 ;
        RECT 829.950 276.600 832.050 277.050 ;
        RECT 835.950 276.600 838.050 277.050 ;
        RECT 829.950 275.400 838.050 276.600 ;
        RECT 829.950 274.950 832.050 275.400 ;
        RECT 835.950 274.950 838.050 275.400 ;
        RECT 748.950 273.600 751.050 274.050 ;
        RECT 784.950 273.600 787.050 274.050 ;
        RECT 748.950 272.400 787.050 273.600 ;
        RECT 748.950 271.950 751.050 272.400 ;
        RECT 784.950 271.950 787.050 272.400 ;
        RECT 757.950 270.600 760.050 271.050 ;
        RECT 760.950 270.600 763.050 271.050 ;
        RECT 757.950 269.400 763.050 270.600 ;
        RECT 757.950 268.950 760.050 269.400 ;
        RECT 760.950 268.950 763.050 269.400 ;
        RECT 766.950 270.600 769.050 271.050 ;
        RECT 766.950 269.400 771.600 270.600 ;
        RECT 766.950 268.950 769.050 269.400 ;
        RECT 715.950 267.600 718.050 268.050 ;
        RECT 670.950 266.400 718.050 267.600 ;
        RECT 670.950 265.950 673.050 266.400 ;
        RECT 715.950 265.950 718.050 266.400 ;
        RECT 742.950 265.950 745.050 268.050 ;
        RECT 761.400 267.600 762.600 268.950 ;
        RECT 766.950 267.600 769.050 268.050 ;
        RECT 761.400 266.400 769.050 267.600 ;
        RECT 770.400 267.600 771.600 269.400 ;
        RECT 808.950 268.950 811.050 271.050 ;
        RECT 838.950 270.600 841.050 271.050 ;
        RECT 847.950 270.600 850.050 271.050 ;
        RECT 838.950 269.400 850.050 270.600 ;
        RECT 838.950 268.950 841.050 269.400 ;
        RECT 847.950 268.950 850.050 269.400 ;
        RECT 790.950 267.600 793.050 268.050 ;
        RECT 770.400 266.400 793.050 267.600 ;
        RECT 766.950 265.950 769.050 266.400 ;
        RECT 790.950 265.950 793.050 266.400 ;
        RECT 598.950 264.600 601.050 265.050 ;
        RECT 628.950 264.600 631.050 265.050 ;
        RECT 598.950 263.400 631.050 264.600 ;
        RECT 598.950 262.950 601.050 263.400 ;
        RECT 628.950 262.950 631.050 263.400 ;
        RECT 646.950 264.600 649.050 265.050 ;
        RECT 661.950 264.600 664.050 265.050 ;
        RECT 646.950 263.400 664.050 264.600 ;
        RECT 646.950 262.950 649.050 263.400 ;
        RECT 661.950 262.950 664.050 263.400 ;
        RECT 673.950 264.600 676.050 265.050 ;
        RECT 772.950 264.600 775.050 265.050 ;
        RECT 673.950 263.400 775.050 264.600 ;
        RECT 673.950 262.950 676.050 263.400 ;
        RECT 772.950 262.950 775.050 263.400 ;
        RECT 809.400 262.050 810.600 268.950 ;
        RECT 616.950 261.600 619.050 262.050 ;
        RECT 596.400 260.400 619.050 261.600 ;
        RECT 556.950 259.950 559.050 260.400 ;
        RECT 571.950 259.950 574.050 260.400 ;
        RECT 589.950 259.950 592.050 260.400 ;
        RECT 616.950 259.950 619.050 260.400 ;
        RECT 619.950 261.600 622.050 262.050 ;
        RECT 640.950 261.600 643.050 262.050 ;
        RECT 652.950 261.600 655.050 262.050 ;
        RECT 619.950 260.400 655.050 261.600 ;
        RECT 619.950 259.950 622.050 260.400 ;
        RECT 640.950 259.950 643.050 260.400 ;
        RECT 652.950 259.950 655.050 260.400 ;
        RECT 676.950 261.600 679.050 262.050 ;
        RECT 682.950 261.600 685.050 262.050 ;
        RECT 676.950 260.400 685.050 261.600 ;
        RECT 676.950 259.950 679.050 260.400 ;
        RECT 682.950 259.950 685.050 260.400 ;
        RECT 688.950 261.600 691.050 262.050 ;
        RECT 694.950 261.600 697.050 262.050 ;
        RECT 688.950 260.400 697.050 261.600 ;
        RECT 688.950 259.950 691.050 260.400 ;
        RECT 694.950 259.950 697.050 260.400 ;
        RECT 697.950 261.600 700.050 262.050 ;
        RECT 736.950 261.600 739.050 262.050 ;
        RECT 697.950 260.400 739.050 261.600 ;
        RECT 697.950 259.950 700.050 260.400 ;
        RECT 736.950 259.950 739.050 260.400 ;
        RECT 751.950 261.600 754.050 262.050 ;
        RECT 769.950 261.600 772.050 262.050 ;
        RECT 751.950 260.400 772.050 261.600 ;
        RECT 751.950 259.950 754.050 260.400 ;
        RECT 769.950 259.950 772.050 260.400 ;
        RECT 808.950 259.950 811.050 262.050 ;
        RECT 49.950 258.600 52.050 259.050 ;
        RECT 85.950 258.600 88.050 259.050 ;
        RECT 49.950 257.400 88.050 258.600 ;
        RECT 49.950 256.950 52.050 257.400 ;
        RECT 85.950 256.950 88.050 257.400 ;
        RECT 103.950 258.600 106.050 259.050 ;
        RECT 112.950 258.600 115.050 259.050 ;
        RECT 124.950 258.600 127.050 259.050 ;
        RECT 103.950 257.400 127.050 258.600 ;
        RECT 103.950 256.950 106.050 257.400 ;
        RECT 112.950 256.950 115.050 257.400 ;
        RECT 124.950 256.950 127.050 257.400 ;
        RECT 130.950 258.600 133.050 259.050 ;
        RECT 136.950 258.600 139.050 259.050 ;
        RECT 130.950 257.400 139.050 258.600 ;
        RECT 130.950 256.950 133.050 257.400 ;
        RECT 136.950 256.950 139.050 257.400 ;
        RECT 169.950 258.600 172.050 259.050 ;
        RECT 220.950 258.600 223.050 259.050 ;
        RECT 169.950 257.400 223.050 258.600 ;
        RECT 169.950 256.950 172.050 257.400 ;
        RECT 220.950 256.950 223.050 257.400 ;
        RECT 268.950 258.600 271.050 259.050 ;
        RECT 316.950 258.600 319.050 259.050 ;
        RECT 268.950 257.400 319.050 258.600 ;
        RECT 268.950 256.950 271.050 257.400 ;
        RECT 316.950 256.950 319.050 257.400 ;
        RECT 346.950 258.600 349.050 259.050 ;
        RECT 391.950 258.600 394.050 259.050 ;
        RECT 346.950 257.400 394.050 258.600 ;
        RECT 346.950 256.950 349.050 257.400 ;
        RECT 391.950 256.950 394.050 257.400 ;
        RECT 394.950 258.600 397.050 259.050 ;
        RECT 424.950 258.600 427.050 259.050 ;
        RECT 394.950 257.400 427.050 258.600 ;
        RECT 394.950 256.950 397.050 257.400 ;
        RECT 424.950 256.950 427.050 257.400 ;
        RECT 430.950 258.600 433.050 259.050 ;
        RECT 436.950 258.600 439.050 259.050 ;
        RECT 460.950 258.600 463.050 259.050 ;
        RECT 430.950 257.400 463.050 258.600 ;
        RECT 430.950 256.950 433.050 257.400 ;
        RECT 436.950 256.950 439.050 257.400 ;
        RECT 460.950 256.950 463.050 257.400 ;
        RECT 469.950 258.600 472.050 259.050 ;
        RECT 487.950 258.600 490.050 259.050 ;
        RECT 499.950 258.600 502.050 259.050 ;
        RECT 469.950 257.400 490.050 258.600 ;
        RECT 469.950 256.950 472.050 257.400 ;
        RECT 487.950 256.950 490.050 257.400 ;
        RECT 491.400 257.400 502.050 258.600 ;
        RECT 25.950 255.600 28.050 256.050 ;
        RECT 34.950 255.600 37.050 256.050 ;
        RECT 25.950 254.400 37.050 255.600 ;
        RECT 25.950 253.950 28.050 254.400 ;
        RECT 34.950 253.950 37.050 254.400 ;
        RECT 61.950 255.600 64.050 256.050 ;
        RECT 67.950 255.600 70.050 256.050 ;
        RECT 61.950 254.400 70.050 255.600 ;
        RECT 61.950 253.950 64.050 254.400 ;
        RECT 67.950 253.950 70.050 254.400 ;
        RECT 76.950 255.600 79.050 256.050 ;
        RECT 97.950 255.600 100.050 256.050 ;
        RECT 76.950 254.400 100.050 255.600 ;
        RECT 76.950 253.950 79.050 254.400 ;
        RECT 97.950 253.950 100.050 254.400 ;
        RECT 100.950 255.600 103.050 256.050 ;
        RECT 118.950 255.600 121.050 256.050 ;
        RECT 100.950 254.400 121.050 255.600 ;
        RECT 100.950 253.950 103.050 254.400 ;
        RECT 118.950 253.950 121.050 254.400 ;
        RECT 133.950 255.600 136.050 256.050 ;
        RECT 325.950 255.600 328.050 256.050 ;
        RECT 367.950 255.600 370.050 256.050 ;
        RECT 133.950 254.400 370.050 255.600 ;
        RECT 133.950 253.950 136.050 254.400 ;
        RECT 325.950 253.950 328.050 254.400 ;
        RECT 367.950 253.950 370.050 254.400 ;
        RECT 376.950 255.600 379.050 256.050 ;
        RECT 406.950 255.600 409.050 256.050 ;
        RECT 376.950 254.400 409.050 255.600 ;
        RECT 376.950 253.950 379.050 254.400 ;
        RECT 406.950 253.950 409.050 254.400 ;
        RECT 445.950 255.600 448.050 256.050 ;
        RECT 491.400 255.600 492.600 257.400 ;
        RECT 499.950 256.950 502.050 257.400 ;
        RECT 523.950 258.600 526.050 259.050 ;
        RECT 547.950 258.600 550.050 259.050 ;
        RECT 523.950 257.400 550.050 258.600 ;
        RECT 523.950 256.950 526.050 257.400 ;
        RECT 547.950 256.950 550.050 257.400 ;
        RECT 559.950 258.600 562.050 259.050 ;
        RECT 574.950 258.600 577.050 259.050 ;
        RECT 559.950 257.400 577.050 258.600 ;
        RECT 559.950 256.950 562.050 257.400 ;
        RECT 574.950 256.950 577.050 257.400 ;
        RECT 628.950 258.600 631.050 259.050 ;
        RECT 709.950 258.600 712.050 259.050 ;
        RECT 628.950 257.400 712.050 258.600 ;
        RECT 628.950 256.950 631.050 257.400 ;
        RECT 709.950 256.950 712.050 257.400 ;
        RECT 739.950 258.600 742.050 259.050 ;
        RECT 757.950 258.600 760.050 259.050 ;
        RECT 739.950 257.400 760.050 258.600 ;
        RECT 739.950 256.950 742.050 257.400 ;
        RECT 757.950 256.950 760.050 257.400 ;
        RECT 787.950 258.600 790.050 259.050 ;
        RECT 802.950 258.600 805.050 259.050 ;
        RECT 787.950 257.400 805.050 258.600 ;
        RECT 787.950 256.950 790.050 257.400 ;
        RECT 802.950 256.950 805.050 257.400 ;
        RECT 805.950 258.600 808.050 259.050 ;
        RECT 844.950 258.600 847.050 259.050 ;
        RECT 805.950 257.400 847.050 258.600 ;
        RECT 805.950 256.950 808.050 257.400 ;
        RECT 844.950 256.950 847.050 257.400 ;
        RECT 445.950 254.400 492.600 255.600 ;
        RECT 493.950 255.600 496.050 256.050 ;
        RECT 514.950 255.600 517.050 256.050 ;
        RECT 493.950 254.400 517.050 255.600 ;
        RECT 445.950 253.950 448.050 254.400 ;
        RECT 493.950 253.950 496.050 254.400 ;
        RECT 514.950 253.950 517.050 254.400 ;
        RECT 526.950 255.600 529.050 256.050 ;
        RECT 535.950 255.600 538.050 256.050 ;
        RECT 526.950 254.400 538.050 255.600 ;
        RECT 526.950 253.950 529.050 254.400 ;
        RECT 535.950 253.950 538.050 254.400 ;
        RECT 541.950 255.600 544.050 256.050 ;
        RECT 547.950 255.600 550.050 256.050 ;
        RECT 541.950 254.400 550.050 255.600 ;
        RECT 541.950 253.950 544.050 254.400 ;
        RECT 547.950 253.950 550.050 254.400 ;
        RECT 571.950 255.600 574.050 256.050 ;
        RECT 634.950 255.600 637.050 256.050 ;
        RECT 733.950 255.600 736.050 256.050 ;
        RECT 571.950 254.400 736.050 255.600 ;
        RECT 571.950 253.950 574.050 254.400 ;
        RECT 634.950 253.950 637.050 254.400 ;
        RECT 733.950 253.950 736.050 254.400 ;
        RECT 766.950 255.600 769.050 256.050 ;
        RECT 814.950 255.600 817.050 256.050 ;
        RECT 766.950 254.400 817.050 255.600 ;
        RECT 766.950 253.950 769.050 254.400 ;
        RECT 814.950 253.950 817.050 254.400 ;
        RECT 817.950 255.600 820.050 256.050 ;
        RECT 832.950 255.600 835.050 256.050 ;
        RECT 817.950 254.400 835.050 255.600 ;
        RECT 817.950 253.950 820.050 254.400 ;
        RECT 832.950 253.950 835.050 254.400 ;
        RECT 25.950 252.600 28.050 253.050 ;
        RECT 103.950 252.600 106.050 253.050 ;
        RECT 25.950 251.400 106.050 252.600 ;
        RECT 25.950 250.950 28.050 251.400 ;
        RECT 103.950 250.950 106.050 251.400 ;
        RECT 121.950 252.600 124.050 253.050 ;
        RECT 133.950 252.600 136.050 253.050 ;
        RECT 121.950 251.400 136.050 252.600 ;
        RECT 121.950 250.950 124.050 251.400 ;
        RECT 133.950 250.950 136.050 251.400 ;
        RECT 151.950 252.600 154.050 253.050 ;
        RECT 166.950 252.600 169.050 253.050 ;
        RECT 151.950 251.400 169.050 252.600 ;
        RECT 151.950 250.950 154.050 251.400 ;
        RECT 166.950 250.950 169.050 251.400 ;
        RECT 181.950 252.600 184.050 253.050 ;
        RECT 346.950 252.600 349.050 253.050 ;
        RECT 412.950 252.600 415.050 253.050 ;
        RECT 181.950 251.400 349.050 252.600 ;
        RECT 181.950 250.950 184.050 251.400 ;
        RECT 346.950 250.950 349.050 251.400 ;
        RECT 350.400 251.400 415.050 252.600 ;
        RECT 16.950 249.600 19.050 250.050 ;
        RECT 28.950 249.600 31.050 250.050 ;
        RECT 16.950 248.400 31.050 249.600 ;
        RECT 16.950 247.950 19.050 248.400 ;
        RECT 28.950 247.950 31.050 248.400 ;
        RECT 31.950 249.600 34.050 250.050 ;
        RECT 43.950 249.600 46.050 250.050 ;
        RECT 91.950 249.600 94.050 250.050 ;
        RECT 31.950 248.400 94.050 249.600 ;
        RECT 31.950 247.950 34.050 248.400 ;
        RECT 43.950 247.950 46.050 248.400 ;
        RECT 91.950 247.950 94.050 248.400 ;
        RECT 112.950 249.600 115.050 250.050 ;
        RECT 160.950 249.600 163.050 250.050 ;
        RECT 112.950 248.400 163.050 249.600 ;
        RECT 112.950 247.950 115.050 248.400 ;
        RECT 160.950 247.950 163.050 248.400 ;
        RECT 163.950 249.600 166.050 250.050 ;
        RECT 214.950 249.600 217.050 250.050 ;
        RECT 238.950 249.600 241.050 250.050 ;
        RECT 163.950 248.400 241.050 249.600 ;
        RECT 163.950 247.950 166.050 248.400 ;
        RECT 214.950 247.950 217.050 248.400 ;
        RECT 238.950 247.950 241.050 248.400 ;
        RECT 268.950 249.600 271.050 250.050 ;
        RECT 328.950 249.600 331.050 250.050 ;
        RECT 268.950 248.400 331.050 249.600 ;
        RECT 268.950 247.950 271.050 248.400 ;
        RECT 328.950 247.950 331.050 248.400 ;
        RECT 331.950 249.600 334.050 250.050 ;
        RECT 350.400 249.600 351.600 251.400 ;
        RECT 412.950 250.950 415.050 251.400 ;
        RECT 415.950 252.600 418.050 253.050 ;
        RECT 439.950 252.600 442.050 253.050 ;
        RECT 415.950 251.400 442.050 252.600 ;
        RECT 415.950 250.950 418.050 251.400 ;
        RECT 439.950 250.950 442.050 251.400 ;
        RECT 448.950 252.600 451.050 253.050 ;
        RECT 508.950 252.600 511.050 253.050 ;
        RECT 448.950 251.400 511.050 252.600 ;
        RECT 448.950 250.950 451.050 251.400 ;
        RECT 508.950 250.950 511.050 251.400 ;
        RECT 514.950 252.600 517.050 253.050 ;
        RECT 529.950 252.600 532.050 253.050 ;
        RECT 514.950 251.400 532.050 252.600 ;
        RECT 514.950 250.950 517.050 251.400 ;
        RECT 529.950 250.950 532.050 251.400 ;
        RECT 532.950 252.600 535.050 253.050 ;
        RECT 541.950 252.600 544.050 253.050 ;
        RECT 532.950 251.400 544.050 252.600 ;
        RECT 532.950 250.950 535.050 251.400 ;
        RECT 541.950 250.950 544.050 251.400 ;
        RECT 559.950 252.600 562.050 253.050 ;
        RECT 700.950 252.600 703.050 253.050 ;
        RECT 559.950 251.400 703.050 252.600 ;
        RECT 559.950 250.950 562.050 251.400 ;
        RECT 700.950 250.950 703.050 251.400 ;
        RECT 727.950 252.600 730.050 253.050 ;
        RECT 733.950 252.600 736.050 253.050 ;
        RECT 727.950 251.400 736.050 252.600 ;
        RECT 727.950 250.950 730.050 251.400 ;
        RECT 733.950 250.950 736.050 251.400 ;
        RECT 745.950 252.600 748.050 253.050 ;
        RECT 784.950 252.600 787.050 253.050 ;
        RECT 745.950 251.400 787.050 252.600 ;
        RECT 745.950 250.950 748.050 251.400 ;
        RECT 784.950 250.950 787.050 251.400 ;
        RECT 823.950 252.600 826.050 253.050 ;
        RECT 850.950 252.600 853.050 253.050 ;
        RECT 823.950 251.400 853.050 252.600 ;
        RECT 823.950 250.950 826.050 251.400 ;
        RECT 850.950 250.950 853.050 251.400 ;
        RECT 331.950 248.400 351.600 249.600 ;
        RECT 409.950 249.600 412.050 250.050 ;
        RECT 427.950 249.600 430.050 250.050 ;
        RECT 409.950 248.400 430.050 249.600 ;
        RECT 331.950 247.950 334.050 248.400 ;
        RECT 409.950 247.950 412.050 248.400 ;
        RECT 427.950 247.950 430.050 248.400 ;
        RECT 454.950 249.600 457.050 250.050 ;
        RECT 565.950 249.600 568.050 250.050 ;
        RECT 454.950 248.400 568.050 249.600 ;
        RECT 454.950 247.950 457.050 248.400 ;
        RECT 565.950 247.950 568.050 248.400 ;
        RECT 568.950 249.600 571.050 250.050 ;
        RECT 574.950 249.600 577.050 250.050 ;
        RECT 670.950 249.600 673.050 250.050 ;
        RECT 568.950 248.400 673.050 249.600 ;
        RECT 568.950 247.950 571.050 248.400 ;
        RECT 574.950 247.950 577.050 248.400 ;
        RECT 670.950 247.950 673.050 248.400 ;
        RECT 691.950 249.600 694.050 250.050 ;
        RECT 700.950 249.600 703.050 250.050 ;
        RECT 691.950 248.400 703.050 249.600 ;
        RECT 691.950 247.950 694.050 248.400 ;
        RECT 700.950 247.950 703.050 248.400 ;
        RECT 742.950 249.600 745.050 250.050 ;
        RECT 751.950 249.600 754.050 250.050 ;
        RECT 742.950 248.400 754.050 249.600 ;
        RECT 742.950 247.950 745.050 248.400 ;
        RECT 751.950 247.950 754.050 248.400 ;
        RECT 754.950 249.600 757.050 250.050 ;
        RECT 808.950 249.600 811.050 250.050 ;
        RECT 754.950 248.400 811.050 249.600 ;
        RECT 754.950 247.950 757.050 248.400 ;
        RECT 808.950 247.950 811.050 248.400 ;
        RECT 13.950 246.600 16.050 247.050 ;
        RECT 8.400 245.400 16.050 246.600 ;
        RECT 8.400 235.050 9.600 245.400 ;
        RECT 13.950 244.950 16.050 245.400 ;
        RECT 28.950 246.600 31.050 247.050 ;
        RECT 49.950 246.600 52.050 247.050 ;
        RECT 94.950 246.600 97.050 247.050 ;
        RECT 106.950 246.600 109.050 247.050 ;
        RECT 28.950 245.400 109.050 246.600 ;
        RECT 28.950 244.950 31.050 245.400 ;
        RECT 49.950 244.950 52.050 245.400 ;
        RECT 94.950 244.950 97.050 245.400 ;
        RECT 106.950 244.950 109.050 245.400 ;
        RECT 109.950 246.600 112.050 247.050 ;
        RECT 118.950 246.600 121.050 247.050 ;
        RECT 109.950 245.400 121.050 246.600 ;
        RECT 109.950 244.950 112.050 245.400 ;
        RECT 118.950 244.950 121.050 245.400 ;
        RECT 133.950 246.600 136.050 247.050 ;
        RECT 139.950 246.600 142.050 247.050 ;
        RECT 133.950 245.400 142.050 246.600 ;
        RECT 133.950 244.950 136.050 245.400 ;
        RECT 139.950 244.950 142.050 245.400 ;
        RECT 148.950 246.600 151.050 247.050 ;
        RECT 154.950 246.600 157.050 247.050 ;
        RECT 169.950 246.600 172.050 247.050 ;
        RECT 175.950 246.600 178.050 247.050 ;
        RECT 148.950 245.400 178.050 246.600 ;
        RECT 148.950 244.950 151.050 245.400 ;
        RECT 154.950 244.950 157.050 245.400 ;
        RECT 169.950 244.950 172.050 245.400 ;
        RECT 175.950 244.950 178.050 245.400 ;
        RECT 187.950 246.600 190.050 247.050 ;
        RECT 199.950 246.600 202.050 247.050 ;
        RECT 187.950 245.400 202.050 246.600 ;
        RECT 187.950 244.950 190.050 245.400 ;
        RECT 199.950 244.950 202.050 245.400 ;
        RECT 232.950 246.600 235.050 247.050 ;
        RECT 250.950 246.600 253.050 247.050 ;
        RECT 232.950 245.400 253.050 246.600 ;
        RECT 232.950 244.950 235.050 245.400 ;
        RECT 250.950 244.950 253.050 245.400 ;
        RECT 253.950 246.600 256.050 247.050 ;
        RECT 262.950 246.600 265.050 247.050 ;
        RECT 253.950 245.400 265.050 246.600 ;
        RECT 253.950 244.950 256.050 245.400 ;
        RECT 262.950 244.950 265.050 245.400 ;
        RECT 382.950 246.600 385.050 247.050 ;
        RECT 406.950 246.600 409.050 247.050 ;
        RECT 382.950 245.400 409.050 246.600 ;
        RECT 382.950 244.950 385.050 245.400 ;
        RECT 406.950 244.950 409.050 245.400 ;
        RECT 511.950 246.600 514.050 247.050 ;
        RECT 538.950 246.600 541.050 247.050 ;
        RECT 511.950 245.400 541.050 246.600 ;
        RECT 511.950 244.950 514.050 245.400 ;
        RECT 538.950 244.950 541.050 245.400 ;
        RECT 541.950 246.600 544.050 247.050 ;
        RECT 562.950 246.600 565.050 247.050 ;
        RECT 541.950 245.400 565.050 246.600 ;
        RECT 541.950 244.950 544.050 245.400 ;
        RECT 562.950 244.950 565.050 245.400 ;
        RECT 565.950 246.600 568.050 247.050 ;
        RECT 580.950 246.600 583.050 247.050 ;
        RECT 583.950 246.600 586.050 247.050 ;
        RECT 565.950 245.400 586.050 246.600 ;
        RECT 565.950 244.950 568.050 245.400 ;
        RECT 580.950 244.950 583.050 245.400 ;
        RECT 583.950 244.950 586.050 245.400 ;
        RECT 589.950 246.600 592.050 247.050 ;
        RECT 595.950 246.600 598.050 247.050 ;
        RECT 589.950 245.400 598.050 246.600 ;
        RECT 589.950 244.950 592.050 245.400 ;
        RECT 595.950 244.950 598.050 245.400 ;
        RECT 616.950 246.600 619.050 247.050 ;
        RECT 643.950 246.600 646.050 247.050 ;
        RECT 616.950 245.400 646.050 246.600 ;
        RECT 616.950 244.950 619.050 245.400 ;
        RECT 643.950 244.950 646.050 245.400 ;
        RECT 655.950 246.600 658.050 247.050 ;
        RECT 691.950 246.600 694.050 247.050 ;
        RECT 655.950 245.400 694.050 246.600 ;
        RECT 655.950 244.950 658.050 245.400 ;
        RECT 691.950 244.950 694.050 245.400 ;
        RECT 712.950 246.600 715.050 247.050 ;
        RECT 718.950 246.600 721.050 247.050 ;
        RECT 712.950 245.400 721.050 246.600 ;
        RECT 712.950 244.950 715.050 245.400 ;
        RECT 718.950 244.950 721.050 245.400 ;
        RECT 730.950 246.600 733.050 247.050 ;
        RECT 835.950 246.600 838.050 247.050 ;
        RECT 730.950 245.400 838.050 246.600 ;
        RECT 730.950 244.950 733.050 245.400 ;
        RECT 835.950 244.950 838.050 245.400 ;
        RECT 37.950 243.600 40.050 244.050 ;
        RECT 145.950 243.600 148.050 244.050 ;
        RECT 37.950 242.400 148.050 243.600 ;
        RECT 37.950 241.950 40.050 242.400 ;
        RECT 145.950 241.950 148.050 242.400 ;
        RECT 163.950 241.950 166.050 244.050 ;
        RECT 166.950 243.600 169.050 244.050 ;
        RECT 181.950 243.600 184.050 244.050 ;
        RECT 166.950 242.400 184.050 243.600 ;
        RECT 166.950 241.950 169.050 242.400 ;
        RECT 181.950 241.950 184.050 242.400 ;
        RECT 193.950 243.600 196.050 244.050 ;
        RECT 208.950 243.600 211.050 244.050 ;
        RECT 193.950 242.400 211.050 243.600 ;
        RECT 193.950 241.950 196.050 242.400 ;
        RECT 208.950 241.950 211.050 242.400 ;
        RECT 214.950 243.600 217.050 244.050 ;
        RECT 256.950 243.600 259.050 244.050 ;
        RECT 214.950 242.400 259.050 243.600 ;
        RECT 214.950 241.950 217.050 242.400 ;
        RECT 256.950 241.950 259.050 242.400 ;
        RECT 274.950 241.950 277.050 244.050 ;
        RECT 277.950 243.600 280.050 244.050 ;
        RECT 289.950 243.600 292.050 244.050 ;
        RECT 277.950 242.400 292.050 243.600 ;
        RECT 277.950 241.950 280.050 242.400 ;
        RECT 289.950 241.950 292.050 242.400 ;
        RECT 310.950 243.600 313.050 244.050 ;
        RECT 310.950 242.400 318.600 243.600 ;
        RECT 310.950 241.950 313.050 242.400 ;
        RECT 19.950 240.600 22.050 241.050 ;
        RECT 37.950 240.600 40.050 241.050 ;
        RECT 19.950 239.400 40.050 240.600 ;
        RECT 19.950 238.950 22.050 239.400 ;
        RECT 37.950 238.950 40.050 239.400 ;
        RECT 55.950 238.950 58.050 241.050 ;
        RECT 64.950 240.600 67.050 241.050 ;
        RECT 85.950 240.600 88.050 241.050 ;
        RECT 106.950 240.600 109.050 241.050 ;
        RECT 164.400 240.600 165.600 241.950 ;
        RECT 64.950 239.400 105.600 240.600 ;
        RECT 64.950 238.950 67.050 239.400 ;
        RECT 85.950 238.950 88.050 239.400 ;
        RECT 10.950 237.600 13.050 238.050 ;
        RECT 22.950 237.600 25.050 238.050 ;
        RECT 10.950 236.400 25.050 237.600 ;
        RECT 38.400 237.600 39.600 238.950 ;
        RECT 38.400 236.400 45.600 237.600 ;
        RECT 10.950 235.950 13.050 236.400 ;
        RECT 22.950 235.950 25.050 236.400 ;
        RECT 44.400 235.050 45.600 236.400 ;
        RECT 7.950 232.950 10.050 235.050 ;
        RECT 43.950 232.950 46.050 235.050 ;
        RECT 52.950 234.600 55.050 235.050 ;
        RECT 56.400 234.600 57.600 238.950 ;
        RECT 70.950 237.600 73.050 238.050 ;
        RECT 62.400 236.400 73.050 237.600 ;
        RECT 52.950 233.400 57.600 234.600 ;
        RECT 58.950 234.600 61.050 235.050 ;
        RECT 62.400 234.600 63.600 236.400 ;
        RECT 70.950 235.950 73.050 236.400 ;
        RECT 73.950 235.950 76.050 238.050 ;
        RECT 76.950 237.600 79.050 238.050 ;
        RECT 94.950 237.600 97.050 238.050 ;
        RECT 76.950 236.400 97.050 237.600 ;
        RECT 104.400 237.600 105.600 239.400 ;
        RECT 106.950 239.400 165.600 240.600 ;
        RECT 196.950 240.600 199.050 241.050 ;
        RECT 205.950 240.600 208.050 241.050 ;
        RECT 226.950 240.600 229.050 241.050 ;
        RECT 196.950 239.400 229.050 240.600 ;
        RECT 106.950 238.950 109.050 239.400 ;
        RECT 196.950 238.950 199.050 239.400 ;
        RECT 205.950 238.950 208.050 239.400 ;
        RECT 226.950 238.950 229.050 239.400 ;
        RECT 235.950 240.600 238.050 241.050 ;
        RECT 241.950 240.600 244.050 241.050 ;
        RECT 235.950 239.400 244.050 240.600 ;
        RECT 235.950 238.950 238.050 239.400 ;
        RECT 241.950 238.950 244.050 239.400 ;
        RECT 250.950 240.600 253.050 241.050 ;
        RECT 259.950 240.600 262.050 241.050 ;
        RECT 250.950 239.400 262.050 240.600 ;
        RECT 250.950 238.950 253.050 239.400 ;
        RECT 259.950 238.950 262.050 239.400 ;
        RECT 265.950 238.950 268.050 241.050 ;
        RECT 124.950 237.600 127.050 238.050 ;
        RECT 104.400 236.400 127.050 237.600 ;
        RECT 76.950 235.950 79.050 236.400 ;
        RECT 94.950 235.950 97.050 236.400 ;
        RECT 124.950 235.950 127.050 236.400 ;
        RECT 136.950 237.600 139.050 238.050 ;
        RECT 148.950 237.600 151.050 238.050 ;
        RECT 136.950 236.400 151.050 237.600 ;
        RECT 136.950 235.950 139.050 236.400 ;
        RECT 148.950 235.950 151.050 236.400 ;
        RECT 178.950 237.600 181.050 238.050 ;
        RECT 184.950 237.600 187.050 238.050 ;
        RECT 266.400 237.600 267.600 238.950 ;
        RECT 178.950 236.400 187.050 237.600 ;
        RECT 178.950 235.950 181.050 236.400 ;
        RECT 184.950 235.950 187.050 236.400 ;
        RECT 227.400 236.400 267.600 237.600 ;
        RECT 271.950 237.600 274.050 238.050 ;
        RECT 275.400 237.600 276.600 241.950 ;
        RECT 283.950 240.600 286.050 241.050 ;
        RECT 301.950 240.600 304.050 241.050 ;
        RECT 283.950 239.400 304.050 240.600 ;
        RECT 283.950 238.950 286.050 239.400 ;
        RECT 301.950 238.950 304.050 239.400 ;
        RECT 271.950 236.400 276.600 237.600 ;
        RECT 280.950 237.600 283.050 238.050 ;
        RECT 280.950 236.400 315.600 237.600 ;
        RECT 58.950 233.400 63.600 234.600 ;
        RECT 64.950 234.600 67.050 235.050 ;
        RECT 74.400 234.600 75.600 235.950 ;
        RECT 64.950 233.400 75.600 234.600 ;
        RECT 76.950 234.600 79.050 235.050 ;
        RECT 103.950 234.600 106.050 235.050 ;
        RECT 76.950 233.400 106.050 234.600 ;
        RECT 52.950 232.950 55.050 233.400 ;
        RECT 58.950 232.950 61.050 233.400 ;
        RECT 64.950 232.950 67.050 233.400 ;
        RECT 76.950 232.950 79.050 233.400 ;
        RECT 103.950 232.950 106.050 233.400 ;
        RECT 124.950 234.600 127.050 235.050 ;
        RECT 130.950 234.600 133.050 235.050 ;
        RECT 124.950 233.400 133.050 234.600 ;
        RECT 124.950 232.950 127.050 233.400 ;
        RECT 130.950 232.950 133.050 233.400 ;
        RECT 160.950 234.600 163.050 235.050 ;
        RECT 181.950 234.600 184.050 235.050 ;
        RECT 211.950 234.600 214.050 235.050 ;
        RECT 160.950 233.400 214.050 234.600 ;
        RECT 160.950 232.950 163.050 233.400 ;
        RECT 181.950 232.950 184.050 233.400 ;
        RECT 211.950 232.950 214.050 233.400 ;
        RECT 223.950 234.600 226.050 235.050 ;
        RECT 227.400 234.600 228.600 236.400 ;
        RECT 271.950 235.950 274.050 236.400 ;
        RECT 280.950 235.950 283.050 236.400 ;
        RECT 314.400 235.050 315.600 236.400 ;
        RECT 223.950 233.400 228.600 234.600 ;
        RECT 229.950 234.600 232.050 235.050 ;
        RECT 253.950 234.600 256.050 235.050 ;
        RECT 262.950 234.600 265.050 235.050 ;
        RECT 229.950 233.400 265.050 234.600 ;
        RECT 223.950 232.950 226.050 233.400 ;
        RECT 229.950 232.950 232.050 233.400 ;
        RECT 253.950 232.950 256.050 233.400 ;
        RECT 262.950 232.950 265.050 233.400 ;
        RECT 280.950 234.600 283.050 235.050 ;
        RECT 298.950 234.600 301.050 235.050 ;
        RECT 310.950 234.600 313.050 235.050 ;
        RECT 280.950 233.400 313.050 234.600 ;
        RECT 280.950 232.950 283.050 233.400 ;
        RECT 298.950 232.950 301.050 233.400 ;
        RECT 310.950 232.950 313.050 233.400 ;
        RECT 313.950 232.950 316.050 235.050 ;
        RECT 317.400 234.600 318.600 242.400 ;
        RECT 337.950 241.950 340.050 244.050 ;
        RECT 397.950 243.600 400.050 244.050 ;
        RECT 418.950 243.600 421.050 244.050 ;
        RECT 397.950 242.400 421.050 243.600 ;
        RECT 397.950 241.950 400.050 242.400 ;
        RECT 418.950 241.950 421.050 242.400 ;
        RECT 421.950 243.600 424.050 244.050 ;
        RECT 430.950 243.600 433.050 244.050 ;
        RECT 421.950 242.400 433.050 243.600 ;
        RECT 421.950 241.950 424.050 242.400 ;
        RECT 430.950 241.950 433.050 242.400 ;
        RECT 439.950 243.600 442.050 244.050 ;
        RECT 466.950 243.600 469.050 244.050 ;
        RECT 439.950 242.400 469.050 243.600 ;
        RECT 439.950 241.950 442.050 242.400 ;
        RECT 466.950 241.950 469.050 242.400 ;
        RECT 469.950 241.950 472.050 244.050 ;
        RECT 487.950 243.600 490.050 244.050 ;
        RECT 493.950 243.600 496.050 244.050 ;
        RECT 487.950 242.400 496.050 243.600 ;
        RECT 487.950 241.950 490.050 242.400 ;
        RECT 493.950 241.950 496.050 242.400 ;
        RECT 505.950 243.600 508.050 244.050 ;
        RECT 505.950 242.400 513.600 243.600 ;
        RECT 505.950 241.950 508.050 242.400 ;
        RECT 338.400 238.050 339.600 241.950 ;
        RECT 364.950 240.600 367.050 241.050 ;
        RECT 382.950 240.600 385.050 241.050 ;
        RECT 397.950 240.600 400.050 241.050 ;
        RECT 364.950 239.400 369.600 240.600 ;
        RECT 364.950 238.950 367.050 239.400 ;
        RECT 337.950 235.950 340.050 238.050 ;
        RECT 364.950 235.950 367.050 238.050 ;
        RECT 317.400 233.400 321.600 234.600 ;
        RECT 320.400 232.050 321.600 233.400 ;
        RECT 16.950 231.600 19.050 232.050 ;
        RECT 67.950 231.600 70.050 232.050 ;
        RECT 118.950 231.600 121.050 232.050 ;
        RECT 16.950 230.400 121.050 231.600 ;
        RECT 16.950 229.950 19.050 230.400 ;
        RECT 67.950 229.950 70.050 230.400 ;
        RECT 118.950 229.950 121.050 230.400 ;
        RECT 157.950 231.600 160.050 232.050 ;
        RECT 211.950 231.600 214.050 232.050 ;
        RECT 238.950 231.600 241.050 232.050 ;
        RECT 157.950 230.400 241.050 231.600 ;
        RECT 157.950 229.950 160.050 230.400 ;
        RECT 211.950 229.950 214.050 230.400 ;
        RECT 238.950 229.950 241.050 230.400 ;
        RECT 244.950 231.600 247.050 232.050 ;
        RECT 274.950 231.600 277.050 232.050 ;
        RECT 244.950 230.400 277.050 231.600 ;
        RECT 244.950 229.950 247.050 230.400 ;
        RECT 274.950 229.950 277.050 230.400 ;
        RECT 307.950 231.600 310.050 232.050 ;
        RECT 313.950 231.600 316.050 232.050 ;
        RECT 307.950 230.400 316.050 231.600 ;
        RECT 307.950 229.950 310.050 230.400 ;
        RECT 313.950 229.950 316.050 230.400 ;
        RECT 319.950 229.950 322.050 232.050 ;
        RECT 70.950 228.600 73.050 229.050 ;
        RECT 76.950 228.600 79.050 229.050 ;
        RECT 70.950 227.400 79.050 228.600 ;
        RECT 70.950 226.950 73.050 227.400 ;
        RECT 76.950 226.950 79.050 227.400 ;
        RECT 103.950 228.600 106.050 229.050 ;
        RECT 199.950 228.600 202.050 229.050 ;
        RECT 103.950 227.400 202.050 228.600 ;
        RECT 103.950 226.950 106.050 227.400 ;
        RECT 199.950 226.950 202.050 227.400 ;
        RECT 205.950 228.600 208.050 229.050 ;
        RECT 223.950 228.600 226.050 229.050 ;
        RECT 205.950 227.400 226.050 228.600 ;
        RECT 205.950 226.950 208.050 227.400 ;
        RECT 223.950 226.950 226.050 227.400 ;
        RECT 298.950 228.600 301.050 229.050 ;
        RECT 316.950 228.600 319.050 229.050 ;
        RECT 298.950 227.400 319.050 228.600 ;
        RECT 365.400 228.600 366.600 235.950 ;
        RECT 368.400 234.600 369.600 239.400 ;
        RECT 382.950 239.400 400.050 240.600 ;
        RECT 382.950 238.950 385.050 239.400 ;
        RECT 397.950 238.950 400.050 239.400 ;
        RECT 424.950 240.600 427.050 241.050 ;
        RECT 442.950 240.600 445.050 241.050 ;
        RECT 470.400 240.600 471.600 241.950 ;
        RECT 424.950 239.400 471.600 240.600 ;
        RECT 478.950 240.600 481.050 241.050 ;
        RECT 493.950 240.600 496.050 241.050 ;
        RECT 508.950 240.600 511.050 241.050 ;
        RECT 478.950 239.400 492.600 240.600 ;
        RECT 424.950 238.950 427.050 239.400 ;
        RECT 442.950 238.950 445.050 239.400 ;
        RECT 478.950 238.950 481.050 239.400 ;
        RECT 385.950 237.600 388.050 238.050 ;
        RECT 394.950 237.600 397.050 238.050 ;
        RECT 457.950 237.600 460.050 238.050 ;
        RECT 463.950 237.600 466.050 238.050 ;
        RECT 385.950 236.400 397.050 237.600 ;
        RECT 385.950 235.950 388.050 236.400 ;
        RECT 394.950 235.950 397.050 236.400 ;
        RECT 422.400 236.400 466.050 237.600 ;
        RECT 491.400 237.600 492.600 239.400 ;
        RECT 493.950 239.400 511.050 240.600 ;
        RECT 512.400 240.600 513.600 242.400 ;
        RECT 529.950 241.950 532.050 244.050 ;
        RECT 568.950 243.600 571.050 244.050 ;
        RECT 533.400 242.400 571.050 243.600 ;
        RECT 514.950 240.600 517.050 241.050 ;
        RECT 512.400 239.400 517.050 240.600 ;
        RECT 493.950 238.950 496.050 239.400 ;
        RECT 508.950 238.950 511.050 239.400 ;
        RECT 514.950 238.950 517.050 239.400 ;
        RECT 530.400 238.050 531.600 241.950 ;
        RECT 533.400 238.050 534.600 242.400 ;
        RECT 568.950 241.950 571.050 242.400 ;
        RECT 607.950 243.600 610.050 244.050 ;
        RECT 619.950 243.600 622.050 244.050 ;
        RECT 607.950 242.400 622.050 243.600 ;
        RECT 607.950 241.950 610.050 242.400 ;
        RECT 619.950 241.950 622.050 242.400 ;
        RECT 625.950 241.950 628.050 244.050 ;
        RECT 634.950 241.950 637.050 244.050 ;
        RECT 658.950 243.600 661.050 244.050 ;
        RECT 667.950 243.600 670.050 244.050 ;
        RECT 658.950 242.400 670.050 243.600 ;
        RECT 658.950 241.950 661.050 242.400 ;
        RECT 667.950 241.950 670.050 242.400 ;
        RECT 706.950 243.600 709.050 244.050 ;
        RECT 739.950 243.600 742.050 244.050 ;
        RECT 706.950 242.400 742.050 243.600 ;
        RECT 706.950 241.950 709.050 242.400 ;
        RECT 739.950 241.950 742.050 242.400 ;
        RECT 742.950 243.600 745.050 244.050 ;
        RECT 778.950 243.600 781.050 244.050 ;
        RECT 742.950 242.400 781.050 243.600 ;
        RECT 742.950 241.950 745.050 242.400 ;
        RECT 778.950 241.950 781.050 242.400 ;
        RECT 793.950 243.600 796.050 244.050 ;
        RECT 799.950 243.600 802.050 244.050 ;
        RECT 793.950 242.400 802.050 243.600 ;
        RECT 793.950 241.950 796.050 242.400 ;
        RECT 799.950 241.950 802.050 242.400 ;
        RECT 802.950 243.600 805.050 244.050 ;
        RECT 835.950 243.600 838.050 244.050 ;
        RECT 853.950 243.600 856.050 244.050 ;
        RECT 802.950 242.400 813.600 243.600 ;
        RECT 802.950 241.950 805.050 242.400 ;
        RECT 541.950 240.600 544.050 241.050 ;
        RECT 547.950 240.600 550.050 241.050 ;
        RECT 583.950 240.600 586.050 241.050 ;
        RECT 541.950 239.400 550.050 240.600 ;
        RECT 541.950 238.950 544.050 239.400 ;
        RECT 547.950 238.950 550.050 239.400 ;
        RECT 581.400 239.400 586.050 240.600 ;
        RECT 581.400 238.050 582.600 239.400 ;
        RECT 583.950 238.950 586.050 239.400 ;
        RECT 601.950 240.600 604.050 241.050 ;
        RECT 613.950 240.600 616.050 241.050 ;
        RECT 601.950 239.400 616.050 240.600 ;
        RECT 601.950 238.950 604.050 239.400 ;
        RECT 613.950 238.950 616.050 239.400 ;
        RECT 626.400 238.050 627.600 241.950 ;
        RECT 635.400 240.600 636.600 241.950 ;
        RECT 637.950 240.600 640.050 241.050 ;
        RECT 635.400 239.400 640.050 240.600 ;
        RECT 637.950 238.950 640.050 239.400 ;
        RECT 640.950 240.600 643.050 241.050 ;
        RECT 652.950 240.600 655.050 241.050 ;
        RECT 640.950 239.400 655.050 240.600 ;
        RECT 640.950 238.950 643.050 239.400 ;
        RECT 652.950 238.950 655.050 239.400 ;
        RECT 670.950 240.600 673.050 241.050 ;
        RECT 697.950 240.600 700.050 241.050 ;
        RECT 670.950 239.400 700.050 240.600 ;
        RECT 670.950 238.950 673.050 239.400 ;
        RECT 697.950 238.950 700.050 239.400 ;
        RECT 712.950 240.600 715.050 241.050 ;
        RECT 721.950 240.600 724.050 241.050 ;
        RECT 712.950 239.400 724.050 240.600 ;
        RECT 712.950 238.950 715.050 239.400 ;
        RECT 721.950 238.950 724.050 239.400 ;
        RECT 727.950 238.950 730.050 241.050 ;
        RECT 760.950 240.600 763.050 241.050 ;
        RECT 766.950 240.600 769.050 241.050 ;
        RECT 760.950 239.400 769.050 240.600 ;
        RECT 760.950 238.950 763.050 239.400 ;
        RECT 766.950 238.950 769.050 239.400 ;
        RECT 778.950 240.600 781.050 241.050 ;
        RECT 796.950 240.600 799.050 241.050 ;
        RECT 802.950 240.600 805.050 241.050 ;
        RECT 808.950 240.600 811.050 241.050 ;
        RECT 778.950 239.400 805.050 240.600 ;
        RECT 778.950 238.950 781.050 239.400 ;
        RECT 796.950 238.950 799.050 239.400 ;
        RECT 802.950 238.950 805.050 239.400 ;
        RECT 806.400 239.400 811.050 240.600 ;
        RECT 520.950 237.600 523.050 238.050 ;
        RECT 491.400 236.400 523.050 237.600 ;
        RECT 376.950 234.600 379.050 235.050 ;
        RECT 368.400 233.400 379.050 234.600 ;
        RECT 376.950 232.950 379.050 233.400 ;
        RECT 397.950 234.600 400.050 235.050 ;
        RECT 422.400 234.600 423.600 236.400 ;
        RECT 457.950 235.950 460.050 236.400 ;
        RECT 463.950 235.950 466.050 236.400 ;
        RECT 520.950 235.950 523.050 236.400 ;
        RECT 529.950 235.950 532.050 238.050 ;
        RECT 532.950 235.950 535.050 238.050 ;
        RECT 580.950 235.950 583.050 238.050 ;
        RECT 610.950 237.600 613.050 238.050 ;
        RECT 608.400 236.400 613.050 237.600 ;
        RECT 397.950 233.400 423.600 234.600 ;
        RECT 448.950 234.600 451.050 235.050 ;
        RECT 502.950 234.600 505.050 235.050 ;
        RECT 517.950 234.600 520.050 235.050 ;
        RECT 526.950 234.600 529.050 235.050 ;
        RECT 448.950 233.400 505.050 234.600 ;
        RECT 397.950 232.950 400.050 233.400 ;
        RECT 448.950 232.950 451.050 233.400 ;
        RECT 502.950 232.950 505.050 233.400 ;
        RECT 506.400 233.400 529.050 234.600 ;
        RECT 367.950 231.600 370.050 232.050 ;
        RECT 388.950 231.600 391.050 232.050 ;
        RECT 367.950 230.400 391.050 231.600 ;
        RECT 367.950 229.950 370.050 230.400 ;
        RECT 388.950 229.950 391.050 230.400 ;
        RECT 391.950 231.600 394.050 232.050 ;
        RECT 400.950 231.600 403.050 232.050 ;
        RECT 412.950 231.600 415.050 232.050 ;
        RECT 391.950 230.400 399.600 231.600 ;
        RECT 391.950 229.950 394.050 230.400 ;
        RECT 394.950 228.600 397.050 229.050 ;
        RECT 365.400 227.400 397.050 228.600 ;
        RECT 398.400 228.600 399.600 230.400 ;
        RECT 400.950 230.400 415.050 231.600 ;
        RECT 400.950 229.950 403.050 230.400 ;
        RECT 412.950 229.950 415.050 230.400 ;
        RECT 433.950 231.600 436.050 232.050 ;
        RECT 506.400 231.600 507.600 233.400 ;
        RECT 517.950 232.950 520.050 233.400 ;
        RECT 526.950 232.950 529.050 233.400 ;
        RECT 553.950 234.600 556.050 235.050 ;
        RECT 559.950 234.600 562.050 235.050 ;
        RECT 562.950 234.600 565.050 235.050 ;
        RECT 553.950 233.400 565.050 234.600 ;
        RECT 553.950 232.950 556.050 233.400 ;
        RECT 559.950 232.950 562.050 233.400 ;
        RECT 562.950 232.950 565.050 233.400 ;
        RECT 568.950 232.950 571.050 235.050 ;
        RECT 601.950 234.600 604.050 235.050 ;
        RECT 608.400 234.600 609.600 236.400 ;
        RECT 610.950 235.950 613.050 236.400 ;
        RECT 613.950 237.600 616.050 238.050 ;
        RECT 622.950 237.600 625.050 238.050 ;
        RECT 613.950 236.400 625.050 237.600 ;
        RECT 613.950 235.950 616.050 236.400 ;
        RECT 622.950 235.950 625.050 236.400 ;
        RECT 625.950 235.950 628.050 238.050 ;
        RECT 655.950 237.600 658.050 238.050 ;
        RECT 653.400 236.400 658.050 237.600 ;
        RECT 653.400 235.050 654.600 236.400 ;
        RECT 655.950 235.950 658.050 236.400 ;
        RECT 667.950 237.600 670.050 238.050 ;
        RECT 671.400 237.600 672.600 238.950 ;
        RECT 667.950 236.400 672.600 237.600 ;
        RECT 679.950 237.600 682.050 238.050 ;
        RECT 685.950 237.600 688.050 238.050 ;
        RECT 679.950 236.400 688.050 237.600 ;
        RECT 667.950 235.950 670.050 236.400 ;
        RECT 679.950 235.950 682.050 236.400 ;
        RECT 685.950 235.950 688.050 236.400 ;
        RECT 724.950 237.600 727.050 238.050 ;
        RECT 728.400 237.600 729.600 238.950 ;
        RECT 724.950 236.400 729.600 237.600 ;
        RECT 763.950 237.600 766.050 238.050 ;
        RECT 769.950 237.600 772.050 238.050 ;
        RECT 763.950 236.400 772.050 237.600 ;
        RECT 724.950 235.950 727.050 236.400 ;
        RECT 763.950 235.950 766.050 236.400 ;
        RECT 769.950 235.950 772.050 236.400 ;
        RECT 775.950 235.950 778.050 238.050 ;
        RECT 787.950 237.600 790.050 238.050 ;
        RECT 793.950 237.600 796.050 238.050 ;
        RECT 806.400 237.600 807.600 239.400 ;
        RECT 808.950 238.950 811.050 239.400 ;
        RECT 787.950 236.400 792.600 237.600 ;
        RECT 787.950 235.950 790.050 236.400 ;
        RECT 601.950 233.400 609.600 234.600 ;
        RECT 610.950 234.600 613.050 235.050 ;
        RECT 625.950 234.600 628.050 235.050 ;
        RECT 610.950 233.400 628.050 234.600 ;
        RECT 601.950 232.950 604.050 233.400 ;
        RECT 610.950 232.950 613.050 233.400 ;
        RECT 625.950 232.950 628.050 233.400 ;
        RECT 652.950 232.950 655.050 235.050 ;
        RECT 655.950 234.600 658.050 235.050 ;
        RECT 706.950 234.600 709.050 235.050 ;
        RECT 715.950 234.600 718.050 235.050 ;
        RECT 655.950 233.400 718.050 234.600 ;
        RECT 655.950 232.950 658.050 233.400 ;
        RECT 706.950 232.950 709.050 233.400 ;
        RECT 715.950 232.950 718.050 233.400 ;
        RECT 433.950 230.400 507.600 231.600 ;
        RECT 511.950 231.600 514.050 232.050 ;
        RECT 526.950 231.600 529.050 232.050 ;
        RECT 529.950 231.600 532.050 232.050 ;
        RECT 541.950 231.600 544.050 232.050 ;
        RECT 511.950 230.400 532.050 231.600 ;
        RECT 433.950 229.950 436.050 230.400 ;
        RECT 511.950 229.950 514.050 230.400 ;
        RECT 526.950 229.950 529.050 230.400 ;
        RECT 529.950 229.950 532.050 230.400 ;
        RECT 533.400 230.400 544.050 231.600 ;
        RECT 409.950 228.600 412.050 229.050 ;
        RECT 398.400 227.400 412.050 228.600 ;
        RECT 298.950 226.950 301.050 227.400 ;
        RECT 316.950 226.950 319.050 227.400 ;
        RECT 394.950 226.950 397.050 227.400 ;
        RECT 409.950 226.950 412.050 227.400 ;
        RECT 415.950 228.600 418.050 229.050 ;
        RECT 427.950 228.600 430.050 229.050 ;
        RECT 415.950 227.400 430.050 228.600 ;
        RECT 415.950 226.950 418.050 227.400 ;
        RECT 427.950 226.950 430.050 227.400 ;
        RECT 433.950 228.600 436.050 229.050 ;
        RECT 445.950 228.600 448.050 229.050 ;
        RECT 433.950 227.400 448.050 228.600 ;
        RECT 433.950 226.950 436.050 227.400 ;
        RECT 445.950 226.950 448.050 227.400 ;
        RECT 481.950 228.600 484.050 229.050 ;
        RECT 487.950 228.600 490.050 229.050 ;
        RECT 481.950 227.400 490.050 228.600 ;
        RECT 481.950 226.950 484.050 227.400 ;
        RECT 487.950 226.950 490.050 227.400 ;
        RECT 502.950 228.600 505.050 229.050 ;
        RECT 533.400 228.600 534.600 230.400 ;
        RECT 541.950 229.950 544.050 230.400 ;
        RECT 550.950 231.600 553.050 232.050 ;
        RECT 556.950 231.600 559.050 232.050 ;
        RECT 550.950 230.400 559.050 231.600 ;
        RECT 569.400 231.600 570.600 232.950 ;
        RECT 571.950 231.600 574.050 232.050 ;
        RECT 706.950 231.600 709.050 232.050 ;
        RECT 569.400 230.400 574.050 231.600 ;
        RECT 550.950 229.950 553.050 230.400 ;
        RECT 556.950 229.950 559.050 230.400 ;
        RECT 571.950 229.950 574.050 230.400 ;
        RECT 632.400 230.400 709.050 231.600 ;
        RECT 502.950 227.400 534.600 228.600 ;
        RECT 535.950 228.600 538.050 229.050 ;
        RECT 580.950 228.600 583.050 229.050 ;
        RECT 535.950 227.400 583.050 228.600 ;
        RECT 502.950 226.950 505.050 227.400 ;
        RECT 535.950 226.950 538.050 227.400 ;
        RECT 580.950 226.950 583.050 227.400 ;
        RECT 598.950 228.600 601.050 229.050 ;
        RECT 632.400 228.600 633.600 230.400 ;
        RECT 706.950 229.950 709.050 230.400 ;
        RECT 709.950 231.600 712.050 232.050 ;
        RECT 736.950 231.600 739.050 232.050 ;
        RECT 760.950 231.600 763.050 232.050 ;
        RECT 709.950 230.400 763.050 231.600 ;
        RECT 776.400 231.600 777.600 235.950 ;
        RECT 791.400 234.600 792.600 236.400 ;
        RECT 793.950 236.400 807.600 237.600 ;
        RECT 812.400 237.600 813.600 242.400 ;
        RECT 835.950 242.400 856.050 243.600 ;
        RECT 835.950 241.950 838.050 242.400 ;
        RECT 853.950 241.950 856.050 242.400 ;
        RECT 832.950 237.600 835.050 238.050 ;
        RECT 812.400 236.400 835.050 237.600 ;
        RECT 793.950 235.950 796.050 236.400 ;
        RECT 832.950 235.950 835.050 236.400 ;
        RECT 841.950 237.600 844.050 238.050 ;
        RECT 847.950 237.600 850.050 238.050 ;
        RECT 853.950 237.600 856.050 238.050 ;
        RECT 841.950 236.400 856.050 237.600 ;
        RECT 841.950 235.950 844.050 236.400 ;
        RECT 847.950 235.950 850.050 236.400 ;
        RECT 853.950 235.950 856.050 236.400 ;
        RECT 808.950 234.600 811.050 235.050 ;
        RECT 791.400 233.400 811.050 234.600 ;
        RECT 808.950 232.950 811.050 233.400 ;
        RECT 814.950 234.600 817.050 235.050 ;
        RECT 823.950 234.600 826.050 235.050 ;
        RECT 814.950 233.400 826.050 234.600 ;
        RECT 814.950 232.950 817.050 233.400 ;
        RECT 823.950 232.950 826.050 233.400 ;
        RECT 829.950 234.600 832.050 235.050 ;
        RECT 844.950 234.600 847.050 235.050 ;
        RECT 829.950 233.400 847.050 234.600 ;
        RECT 829.950 232.950 832.050 233.400 ;
        RECT 844.950 232.950 847.050 233.400 ;
        RECT 850.950 234.600 853.050 235.050 ;
        RECT 859.950 234.600 862.050 235.050 ;
        RECT 850.950 233.400 862.050 234.600 ;
        RECT 850.950 232.950 853.050 233.400 ;
        RECT 859.950 232.950 862.050 233.400 ;
        RECT 787.950 231.600 790.050 232.050 ;
        RECT 776.400 230.400 790.050 231.600 ;
        RECT 709.950 229.950 712.050 230.400 ;
        RECT 736.950 229.950 739.050 230.400 ;
        RECT 760.950 229.950 763.050 230.400 ;
        RECT 787.950 229.950 790.050 230.400 ;
        RECT 598.950 227.400 633.600 228.600 ;
        RECT 634.950 228.600 637.050 229.050 ;
        RECT 673.950 228.600 676.050 229.050 ;
        RECT 688.950 228.600 691.050 229.050 ;
        RECT 634.950 227.400 691.050 228.600 ;
        RECT 598.950 226.950 601.050 227.400 ;
        RECT 634.950 226.950 637.050 227.400 ;
        RECT 673.950 226.950 676.050 227.400 ;
        RECT 688.950 226.950 691.050 227.400 ;
        RECT 733.950 228.600 736.050 229.050 ;
        RECT 805.950 228.600 808.050 229.050 ;
        RECT 733.950 227.400 808.050 228.600 ;
        RECT 733.950 226.950 736.050 227.400 ;
        RECT 805.950 226.950 808.050 227.400 ;
        RECT 61.950 225.600 64.050 226.050 ;
        RECT 124.950 225.600 127.050 226.050 ;
        RECT 61.950 224.400 127.050 225.600 ;
        RECT 61.950 223.950 64.050 224.400 ;
        RECT 124.950 223.950 127.050 224.400 ;
        RECT 139.950 225.600 142.050 226.050 ;
        RECT 193.950 225.600 196.050 226.050 ;
        RECT 139.950 224.400 196.050 225.600 ;
        RECT 139.950 223.950 142.050 224.400 ;
        RECT 193.950 223.950 196.050 224.400 ;
        RECT 349.950 225.600 352.050 226.050 ;
        RECT 373.950 225.600 376.050 226.050 ;
        RECT 349.950 224.400 376.050 225.600 ;
        RECT 349.950 223.950 352.050 224.400 ;
        RECT 373.950 223.950 376.050 224.400 ;
        RECT 379.950 225.600 382.050 226.050 ;
        RECT 430.950 225.600 433.050 226.050 ;
        RECT 379.950 224.400 433.050 225.600 ;
        RECT 379.950 223.950 382.050 224.400 ;
        RECT 430.950 223.950 433.050 224.400 ;
        RECT 439.950 225.600 442.050 226.050 ;
        RECT 451.950 225.600 454.050 226.050 ;
        RECT 574.950 225.600 577.050 226.050 ;
        RECT 439.950 224.400 454.050 225.600 ;
        RECT 439.950 223.950 442.050 224.400 ;
        RECT 451.950 223.950 454.050 224.400 ;
        RECT 455.400 224.400 577.050 225.600 ;
        RECT 1.950 222.600 4.050 223.050 ;
        RECT 64.950 222.600 67.050 223.050 ;
        RECT 1.950 221.400 67.050 222.600 ;
        RECT 1.950 220.950 4.050 221.400 ;
        RECT 64.950 220.950 67.050 221.400 ;
        RECT 88.950 222.600 91.050 223.050 ;
        RECT 148.950 222.600 151.050 223.050 ;
        RECT 88.950 221.400 151.050 222.600 ;
        RECT 88.950 220.950 91.050 221.400 ;
        RECT 148.950 220.950 151.050 221.400 ;
        RECT 220.950 222.600 223.050 223.050 ;
        RECT 274.950 222.600 277.050 223.050 ;
        RECT 455.400 222.600 456.600 224.400 ;
        RECT 574.950 223.950 577.050 224.400 ;
        RECT 577.950 225.600 580.050 226.050 ;
        RECT 604.950 225.600 607.050 226.050 ;
        RECT 616.950 225.600 619.050 226.050 ;
        RECT 577.950 224.400 619.050 225.600 ;
        RECT 577.950 223.950 580.050 224.400 ;
        RECT 604.950 223.950 607.050 224.400 ;
        RECT 616.950 223.950 619.050 224.400 ;
        RECT 628.950 225.600 631.050 226.050 ;
        RECT 661.950 225.600 664.050 226.050 ;
        RECT 628.950 224.400 664.050 225.600 ;
        RECT 628.950 223.950 631.050 224.400 ;
        RECT 661.950 223.950 664.050 224.400 ;
        RECT 670.950 225.600 673.050 226.050 ;
        RECT 682.950 225.600 685.050 226.050 ;
        RECT 670.950 224.400 685.050 225.600 ;
        RECT 670.950 223.950 673.050 224.400 ;
        RECT 682.950 223.950 685.050 224.400 ;
        RECT 706.950 225.600 709.050 226.050 ;
        RECT 826.950 225.600 829.050 226.050 ;
        RECT 838.950 225.600 841.050 226.050 ;
        RECT 706.950 224.400 841.050 225.600 ;
        RECT 706.950 223.950 709.050 224.400 ;
        RECT 826.950 223.950 829.050 224.400 ;
        RECT 838.950 223.950 841.050 224.400 ;
        RECT 220.950 221.400 456.600 222.600 ;
        RECT 457.950 222.600 460.050 223.050 ;
        RECT 541.950 222.600 544.050 223.050 ;
        RECT 457.950 221.400 544.050 222.600 ;
        RECT 220.950 220.950 223.050 221.400 ;
        RECT 274.950 220.950 277.050 221.400 ;
        RECT 457.950 220.950 460.050 221.400 ;
        RECT 541.950 220.950 544.050 221.400 ;
        RECT 571.950 222.600 574.050 223.050 ;
        RECT 589.950 222.600 592.050 223.050 ;
        RECT 571.950 221.400 592.050 222.600 ;
        RECT 571.950 220.950 574.050 221.400 ;
        RECT 589.950 220.950 592.050 221.400 ;
        RECT 616.950 222.600 619.050 223.050 ;
        RECT 634.950 222.600 637.050 223.050 ;
        RECT 616.950 221.400 637.050 222.600 ;
        RECT 616.950 220.950 619.050 221.400 ;
        RECT 634.950 220.950 637.050 221.400 ;
        RECT 706.950 222.600 709.050 223.050 ;
        RECT 724.950 222.600 727.050 223.050 ;
        RECT 841.950 222.600 844.050 223.050 ;
        RECT 706.950 221.400 844.050 222.600 ;
        RECT 706.950 220.950 709.050 221.400 ;
        RECT 724.950 220.950 727.050 221.400 ;
        RECT 841.950 220.950 844.050 221.400 ;
        RECT 49.950 219.600 52.050 220.050 ;
        RECT 61.950 219.600 64.050 220.050 ;
        RECT 49.950 218.400 64.050 219.600 ;
        RECT 49.950 217.950 52.050 218.400 ;
        RECT 61.950 217.950 64.050 218.400 ;
        RECT 64.950 219.600 67.050 220.050 ;
        RECT 91.950 219.600 94.050 220.050 ;
        RECT 64.950 218.400 94.050 219.600 ;
        RECT 64.950 217.950 67.050 218.400 ;
        RECT 91.950 217.950 94.050 218.400 ;
        RECT 277.950 219.600 280.050 220.050 ;
        RECT 316.950 219.600 319.050 220.050 ;
        RECT 406.950 219.600 409.050 220.050 ;
        RECT 277.950 218.400 315.600 219.600 ;
        RECT 277.950 217.950 280.050 218.400 ;
        RECT 94.950 216.600 97.050 217.050 ;
        RECT 286.950 216.600 289.050 217.050 ;
        RECT 94.950 215.400 289.050 216.600 ;
        RECT 314.400 216.600 315.600 218.400 ;
        RECT 316.950 218.400 409.050 219.600 ;
        RECT 316.950 217.950 319.050 218.400 ;
        RECT 406.950 217.950 409.050 218.400 ;
        RECT 418.950 219.600 421.050 220.050 ;
        RECT 442.950 219.600 445.050 220.050 ;
        RECT 469.950 219.600 472.050 220.050 ;
        RECT 418.950 218.400 472.050 219.600 ;
        RECT 418.950 217.950 421.050 218.400 ;
        RECT 442.950 217.950 445.050 218.400 ;
        RECT 469.950 217.950 472.050 218.400 ;
        RECT 508.950 219.600 511.050 220.050 ;
        RECT 571.950 219.600 574.050 220.050 ;
        RECT 508.950 218.400 574.050 219.600 ;
        RECT 508.950 217.950 511.050 218.400 ;
        RECT 571.950 217.950 574.050 218.400 ;
        RECT 574.950 219.600 577.050 220.050 ;
        RECT 595.950 219.600 598.050 220.050 ;
        RECT 820.950 219.600 823.050 220.050 ;
        RECT 574.950 218.400 823.050 219.600 ;
        RECT 574.950 217.950 577.050 218.400 ;
        RECT 595.950 217.950 598.050 218.400 ;
        RECT 820.950 217.950 823.050 218.400 ;
        RECT 331.950 216.600 334.050 217.050 ;
        RECT 314.400 215.400 334.050 216.600 ;
        RECT 94.950 214.950 97.050 215.400 ;
        RECT 286.950 214.950 289.050 215.400 ;
        RECT 331.950 214.950 334.050 215.400 ;
        RECT 358.950 216.600 361.050 217.050 ;
        RECT 382.950 216.600 385.050 217.050 ;
        RECT 358.950 215.400 385.050 216.600 ;
        RECT 358.950 214.950 361.050 215.400 ;
        RECT 382.950 214.950 385.050 215.400 ;
        RECT 388.950 216.600 391.050 217.050 ;
        RECT 424.950 216.600 427.050 217.050 ;
        RECT 388.950 215.400 427.050 216.600 ;
        RECT 388.950 214.950 391.050 215.400 ;
        RECT 424.950 214.950 427.050 215.400 ;
        RECT 430.950 216.600 433.050 217.050 ;
        RECT 439.950 216.600 442.050 217.050 ;
        RECT 430.950 215.400 442.050 216.600 ;
        RECT 430.950 214.950 433.050 215.400 ;
        RECT 439.950 214.950 442.050 215.400 ;
        RECT 445.950 216.600 448.050 217.050 ;
        RECT 451.950 216.600 454.050 217.050 ;
        RECT 445.950 215.400 454.050 216.600 ;
        RECT 445.950 214.950 448.050 215.400 ;
        RECT 451.950 214.950 454.050 215.400 ;
        RECT 493.950 216.600 496.050 217.050 ;
        RECT 505.950 216.600 508.050 217.050 ;
        RECT 493.950 215.400 508.050 216.600 ;
        RECT 493.950 214.950 496.050 215.400 ;
        RECT 505.950 214.950 508.050 215.400 ;
        RECT 523.950 216.600 526.050 217.050 ;
        RECT 529.950 216.600 532.050 217.050 ;
        RECT 523.950 215.400 532.050 216.600 ;
        RECT 523.950 214.950 526.050 215.400 ;
        RECT 529.950 214.950 532.050 215.400 ;
        RECT 538.950 216.600 541.050 217.050 ;
        RECT 601.950 216.600 604.050 217.050 ;
        RECT 538.950 215.400 604.050 216.600 ;
        RECT 538.950 214.950 541.050 215.400 ;
        RECT 601.950 214.950 604.050 215.400 ;
        RECT 85.950 213.600 88.050 214.050 ;
        RECT 94.950 213.600 97.050 214.050 ;
        RECT 319.950 213.600 322.050 214.050 ;
        RECT 85.950 212.400 97.050 213.600 ;
        RECT 85.950 211.950 88.050 212.400 ;
        RECT 94.950 211.950 97.050 212.400 ;
        RECT 206.400 212.400 322.050 213.600 ;
        RECT 31.950 210.600 34.050 211.050 ;
        RECT 70.950 210.600 73.050 211.050 ;
        RECT 31.950 209.400 73.050 210.600 ;
        RECT 31.950 208.950 34.050 209.400 ;
        RECT 70.950 208.950 73.050 209.400 ;
        RECT 73.950 210.600 76.050 211.050 ;
        RECT 206.400 210.600 207.600 212.400 ;
        RECT 319.950 211.950 322.050 212.400 ;
        RECT 361.950 213.600 364.050 214.050 ;
        RECT 472.950 213.600 475.050 214.050 ;
        RECT 484.950 213.600 487.050 214.050 ;
        RECT 505.950 213.600 508.050 214.050 ;
        RECT 556.950 213.600 559.050 214.050 ;
        RECT 361.950 212.400 559.050 213.600 ;
        RECT 361.950 211.950 364.050 212.400 ;
        RECT 472.950 211.950 475.050 212.400 ;
        RECT 484.950 211.950 487.050 212.400 ;
        RECT 505.950 211.950 508.050 212.400 ;
        RECT 556.950 211.950 559.050 212.400 ;
        RECT 571.950 213.600 574.050 214.050 ;
        RECT 637.950 213.600 640.050 214.050 ;
        RECT 571.950 212.400 640.050 213.600 ;
        RECT 571.950 211.950 574.050 212.400 ;
        RECT 637.950 211.950 640.050 212.400 ;
        RECT 748.950 213.600 751.050 214.050 ;
        RECT 820.950 213.600 823.050 214.050 ;
        RECT 748.950 212.400 823.050 213.600 ;
        RECT 748.950 211.950 751.050 212.400 ;
        RECT 820.950 211.950 823.050 212.400 ;
        RECT 73.950 209.400 207.600 210.600 ;
        RECT 229.950 210.600 232.050 211.050 ;
        RECT 268.950 210.600 271.050 211.050 ;
        RECT 229.950 209.400 271.050 210.600 ;
        RECT 73.950 208.950 76.050 209.400 ;
        RECT 229.950 208.950 232.050 209.400 ;
        RECT 268.950 208.950 271.050 209.400 ;
        RECT 322.950 210.600 325.050 211.050 ;
        RECT 547.950 210.600 550.050 211.050 ;
        RECT 604.950 210.600 607.050 211.050 ;
        RECT 322.950 209.400 607.050 210.600 ;
        RECT 322.950 208.950 325.050 209.400 ;
        RECT 547.950 208.950 550.050 209.400 ;
        RECT 604.950 208.950 607.050 209.400 ;
        RECT 613.950 210.600 616.050 211.050 ;
        RECT 664.950 210.600 667.050 211.050 ;
        RECT 667.950 210.600 670.050 211.050 ;
        RECT 613.950 209.400 670.050 210.600 ;
        RECT 613.950 208.950 616.050 209.400 ;
        RECT 664.950 208.950 667.050 209.400 ;
        RECT 667.950 208.950 670.050 209.400 ;
        RECT 673.950 210.600 676.050 211.050 ;
        RECT 748.950 210.600 751.050 211.050 ;
        RECT 673.950 209.400 751.050 210.600 ;
        RECT 673.950 208.950 676.050 209.400 ;
        RECT 748.950 208.950 751.050 209.400 ;
        RECT 22.950 207.600 25.050 208.050 ;
        RECT 25.950 207.600 28.050 208.050 ;
        RECT 34.950 207.600 37.050 208.050 ;
        RECT 40.950 207.600 43.050 208.050 ;
        RECT 22.950 206.400 43.050 207.600 ;
        RECT 22.950 205.950 25.050 206.400 ;
        RECT 25.950 205.950 28.050 206.400 ;
        RECT 34.950 205.950 37.050 206.400 ;
        RECT 40.950 205.950 43.050 206.400 ;
        RECT 46.950 207.600 49.050 208.050 ;
        RECT 79.950 207.600 82.050 208.050 ;
        RECT 46.950 206.400 82.050 207.600 ;
        RECT 46.950 205.950 49.050 206.400 ;
        RECT 79.950 205.950 82.050 206.400 ;
        RECT 97.950 207.600 100.050 208.050 ;
        RECT 217.950 207.600 220.050 208.050 ;
        RECT 97.950 206.400 220.050 207.600 ;
        RECT 97.950 205.950 100.050 206.400 ;
        RECT 217.950 205.950 220.050 206.400 ;
        RECT 256.950 207.600 259.050 208.050 ;
        RECT 295.950 207.600 298.050 208.050 ;
        RECT 256.950 206.400 298.050 207.600 ;
        RECT 256.950 205.950 259.050 206.400 ;
        RECT 295.950 205.950 298.050 206.400 ;
        RECT 301.950 207.600 304.050 208.050 ;
        RECT 352.950 207.600 355.050 208.050 ;
        RECT 385.950 207.600 388.050 208.050 ;
        RECT 301.950 206.400 355.050 207.600 ;
        RECT 301.950 205.950 304.050 206.400 ;
        RECT 352.950 205.950 355.050 206.400 ;
        RECT 368.400 206.400 388.050 207.600 ;
        RECT 49.950 202.950 52.050 205.050 ;
        RECT 70.950 204.600 73.050 205.050 ;
        RECT 53.400 203.400 73.050 204.600 ;
        RECT 1.950 201.600 4.050 202.050 ;
        RECT 7.950 201.600 10.050 202.050 ;
        RECT 1.950 200.400 10.050 201.600 ;
        RECT 1.950 199.950 4.050 200.400 ;
        RECT 7.950 199.950 10.050 200.400 ;
        RECT 10.950 201.600 13.050 202.050 ;
        RECT 31.950 201.600 34.050 202.050 ;
        RECT 40.950 201.600 43.050 202.050 ;
        RECT 43.950 201.600 46.050 202.050 ;
        RECT 10.950 200.400 46.050 201.600 ;
        RECT 10.950 199.950 13.050 200.400 ;
        RECT 31.950 199.950 34.050 200.400 ;
        RECT 40.950 199.950 43.050 200.400 ;
        RECT 43.950 199.950 46.050 200.400 ;
        RECT 25.950 196.950 28.050 199.050 ;
        RECT 22.950 195.600 25.050 196.050 ;
        RECT 26.400 195.600 27.600 196.950 ;
        RECT 22.950 194.400 27.600 195.600 ;
        RECT 50.400 195.600 51.600 202.950 ;
        RECT 53.400 202.050 54.600 203.400 ;
        RECT 70.950 202.950 73.050 203.400 ;
        RECT 82.950 204.600 85.050 205.050 ;
        RECT 88.950 204.600 91.050 205.050 ;
        RECT 97.950 204.600 100.050 205.050 ;
        RECT 82.950 203.400 100.050 204.600 ;
        RECT 82.950 202.950 85.050 203.400 ;
        RECT 88.950 202.950 91.050 203.400 ;
        RECT 97.950 202.950 100.050 203.400 ;
        RECT 127.950 204.600 130.050 205.050 ;
        RECT 136.950 204.600 139.050 205.050 ;
        RECT 178.950 204.600 181.050 205.050 ;
        RECT 127.950 203.400 181.050 204.600 ;
        RECT 127.950 202.950 130.050 203.400 ;
        RECT 136.950 202.950 139.050 203.400 ;
        RECT 167.400 202.050 168.600 203.400 ;
        RECT 178.950 202.950 181.050 203.400 ;
        RECT 187.950 204.600 190.050 205.050 ;
        RECT 190.950 204.600 193.050 205.050 ;
        RECT 199.950 204.600 202.050 205.050 ;
        RECT 187.950 203.400 202.050 204.600 ;
        RECT 187.950 202.950 190.050 203.400 ;
        RECT 190.950 202.950 193.050 203.400 ;
        RECT 199.950 202.950 202.050 203.400 ;
        RECT 226.950 204.600 229.050 205.050 ;
        RECT 232.950 204.600 235.050 205.050 ;
        RECT 226.950 203.400 235.050 204.600 ;
        RECT 226.950 202.950 229.050 203.400 ;
        RECT 232.950 202.950 235.050 203.400 ;
        RECT 238.950 204.600 241.050 205.050 ;
        RECT 247.950 204.600 250.050 205.050 ;
        RECT 238.950 203.400 250.050 204.600 ;
        RECT 238.950 202.950 241.050 203.400 ;
        RECT 247.950 202.950 250.050 203.400 ;
        RECT 292.950 202.950 295.050 205.050 ;
        RECT 304.950 202.950 307.050 205.050 ;
        RECT 346.950 204.600 349.050 205.050 ;
        RECT 368.400 204.600 369.600 206.400 ;
        RECT 385.950 205.950 388.050 206.400 ;
        RECT 391.950 207.600 394.050 208.050 ;
        RECT 421.950 207.600 424.050 208.050 ;
        RECT 391.950 206.400 424.050 207.600 ;
        RECT 391.950 205.950 394.050 206.400 ;
        RECT 421.950 205.950 424.050 206.400 ;
        RECT 427.950 207.600 430.050 208.050 ;
        RECT 502.950 207.600 505.050 208.050 ;
        RECT 427.950 206.400 505.050 207.600 ;
        RECT 427.950 205.950 430.050 206.400 ;
        RECT 502.950 205.950 505.050 206.400 ;
        RECT 511.950 207.600 514.050 208.050 ;
        RECT 517.950 207.600 520.050 208.050 ;
        RECT 523.950 207.600 526.050 208.050 ;
        RECT 511.950 206.400 516.600 207.600 ;
        RECT 511.950 205.950 514.050 206.400 ;
        RECT 346.950 203.400 369.600 204.600 ;
        RECT 370.950 204.600 373.050 205.050 ;
        RECT 379.950 204.600 382.050 205.050 ;
        RECT 415.950 204.600 418.050 205.050 ;
        RECT 370.950 203.400 382.050 204.600 ;
        RECT 346.950 202.950 349.050 203.400 ;
        RECT 370.950 202.950 373.050 203.400 ;
        RECT 379.950 202.950 382.050 203.400 ;
        RECT 383.400 203.400 418.050 204.600 ;
        RECT 52.950 199.950 55.050 202.050 ;
        RECT 73.950 201.600 76.050 202.050 ;
        RECT 56.400 200.400 76.050 201.600 ;
        RECT 56.400 199.050 57.600 200.400 ;
        RECT 73.950 199.950 76.050 200.400 ;
        RECT 118.950 201.600 121.050 202.050 ;
        RECT 133.950 201.600 136.050 202.050 ;
        RECT 139.950 201.600 142.050 202.050 ;
        RECT 118.950 200.400 142.050 201.600 ;
        RECT 118.950 199.950 121.050 200.400 ;
        RECT 133.950 199.950 136.050 200.400 ;
        RECT 139.950 199.950 142.050 200.400 ;
        RECT 166.950 199.950 169.050 202.050 ;
        RECT 172.950 201.600 175.050 202.050 ;
        RECT 184.950 201.600 187.050 202.050 ;
        RECT 172.950 200.400 180.600 201.600 ;
        RECT 172.950 199.950 175.050 200.400 ;
        RECT 55.950 196.950 58.050 199.050 ;
        RECT 103.950 198.600 106.050 199.050 ;
        RECT 109.950 198.600 112.050 199.050 ;
        RECT 103.950 197.400 112.050 198.600 ;
        RECT 103.950 196.950 106.050 197.400 ;
        RECT 109.950 196.950 112.050 197.400 ;
        RECT 130.950 198.600 133.050 199.050 ;
        RECT 151.950 198.600 154.050 199.050 ;
        RECT 130.950 197.400 154.050 198.600 ;
        RECT 130.950 196.950 133.050 197.400 ;
        RECT 151.950 196.950 154.050 197.400 ;
        RECT 160.950 198.600 163.050 199.050 ;
        RECT 169.950 198.600 172.050 199.050 ;
        RECT 160.950 197.400 172.050 198.600 ;
        RECT 160.950 196.950 163.050 197.400 ;
        RECT 169.950 196.950 172.050 197.400 ;
        RECT 179.400 196.050 180.600 200.400 ;
        RECT 184.950 200.400 192.600 201.600 ;
        RECT 184.950 199.950 187.050 200.400 ;
        RECT 191.400 196.050 192.600 200.400 ;
        RECT 211.950 199.950 214.050 202.050 ;
        RECT 214.950 201.600 217.050 202.050 ;
        RECT 250.950 201.600 253.050 202.050 ;
        RECT 259.950 201.600 262.050 202.050 ;
        RECT 214.950 200.400 262.050 201.600 ;
        RECT 214.950 199.950 217.050 200.400 ;
        RECT 250.950 199.950 253.050 200.400 ;
        RECT 259.950 199.950 262.050 200.400 ;
        RECT 277.950 201.600 280.050 202.050 ;
        RECT 283.950 201.600 286.050 202.050 ;
        RECT 289.950 201.600 292.050 202.050 ;
        RECT 277.950 200.400 292.050 201.600 ;
        RECT 277.950 199.950 280.050 200.400 ;
        RECT 283.950 199.950 286.050 200.400 ;
        RECT 289.950 199.950 292.050 200.400 ;
        RECT 55.950 195.600 58.050 196.050 ;
        RECT 50.400 194.400 58.050 195.600 ;
        RECT 22.950 193.950 25.050 194.400 ;
        RECT 55.950 193.950 58.050 194.400 ;
        RECT 76.950 195.600 79.050 196.050 ;
        RECT 82.950 195.600 85.050 196.050 ;
        RECT 115.950 195.600 118.050 196.050 ;
        RECT 76.950 194.400 118.050 195.600 ;
        RECT 76.950 193.950 79.050 194.400 ;
        RECT 82.950 193.950 85.050 194.400 ;
        RECT 115.950 193.950 118.050 194.400 ;
        RECT 178.950 193.950 181.050 196.050 ;
        RECT 190.950 193.950 193.050 196.050 ;
        RECT 67.950 192.600 70.050 193.050 ;
        RECT 73.950 192.600 76.050 193.050 ;
        RECT 106.950 192.600 109.050 193.050 ;
        RECT 67.950 191.400 109.050 192.600 ;
        RECT 67.950 190.950 70.050 191.400 ;
        RECT 73.950 190.950 76.050 191.400 ;
        RECT 106.950 190.950 109.050 191.400 ;
        RECT 127.950 192.600 130.050 193.050 ;
        RECT 142.950 192.600 145.050 193.050 ;
        RECT 127.950 191.400 145.050 192.600 ;
        RECT 127.950 190.950 130.050 191.400 ;
        RECT 142.950 190.950 145.050 191.400 ;
        RECT 145.950 192.600 148.050 193.050 ;
        RECT 163.950 192.600 166.050 193.050 ;
        RECT 196.950 192.600 199.050 193.050 ;
        RECT 145.950 191.400 199.050 192.600 ;
        RECT 212.400 192.600 213.600 199.950 ;
        RECT 293.400 199.050 294.600 202.950 ;
        RECT 220.950 198.600 223.050 199.050 ;
        RECT 232.950 198.600 235.050 199.050 ;
        RECT 220.950 197.400 235.050 198.600 ;
        RECT 220.950 196.950 223.050 197.400 ;
        RECT 232.950 196.950 235.050 197.400 ;
        RECT 235.950 198.600 238.050 199.050 ;
        RECT 238.950 198.600 241.050 199.050 ;
        RECT 247.950 198.600 250.050 199.050 ;
        RECT 235.950 197.400 250.050 198.600 ;
        RECT 235.950 196.950 238.050 197.400 ;
        RECT 238.950 196.950 241.050 197.400 ;
        RECT 247.950 196.950 250.050 197.400 ;
        RECT 280.950 196.950 283.050 199.050 ;
        RECT 292.950 196.950 295.050 199.050 ;
        RECT 305.400 198.600 306.600 202.950 ;
        RECT 307.950 201.600 310.050 202.050 ;
        RECT 364.950 201.600 367.050 202.050 ;
        RECT 383.400 201.600 384.600 203.400 ;
        RECT 415.950 202.950 418.050 203.400 ;
        RECT 424.950 204.600 427.050 205.050 ;
        RECT 424.950 203.400 513.600 204.600 ;
        RECT 424.950 202.950 427.050 203.400 ;
        RECT 512.400 202.050 513.600 203.400 ;
        RECT 307.950 200.400 315.600 201.600 ;
        RECT 307.950 199.950 310.050 200.400 ;
        RECT 307.950 198.600 310.050 199.050 ;
        RECT 305.400 197.400 310.050 198.600 ;
        RECT 307.950 196.950 310.050 197.400 ;
        RECT 226.950 195.600 229.050 196.050 ;
        RECT 241.950 195.600 244.050 196.050 ;
        RECT 226.950 194.400 244.050 195.600 ;
        RECT 226.950 193.950 229.050 194.400 ;
        RECT 241.950 193.950 244.050 194.400 ;
        RECT 253.950 195.600 256.050 196.050 ;
        RECT 268.950 195.600 271.050 196.050 ;
        RECT 253.950 194.400 271.050 195.600 ;
        RECT 253.950 193.950 256.050 194.400 ;
        RECT 268.950 193.950 271.050 194.400 ;
        RECT 281.400 193.050 282.600 196.950 ;
        RECT 286.950 195.600 289.050 196.050 ;
        RECT 304.950 195.600 307.050 196.050 ;
        RECT 286.950 194.400 307.050 195.600 ;
        RECT 314.400 195.600 315.600 200.400 ;
        RECT 364.950 200.400 384.600 201.600 ;
        RECT 412.950 201.600 415.050 202.050 ;
        RECT 445.950 201.600 448.050 202.050 ;
        RECT 412.950 200.400 448.050 201.600 ;
        RECT 364.950 199.950 367.050 200.400 ;
        RECT 412.950 199.950 415.050 200.400 ;
        RECT 445.950 199.950 448.050 200.400 ;
        RECT 484.950 201.600 487.050 202.050 ;
        RECT 496.950 201.600 499.050 202.050 ;
        RECT 484.950 200.400 499.050 201.600 ;
        RECT 484.950 199.950 487.050 200.400 ;
        RECT 496.950 199.950 499.050 200.400 ;
        RECT 511.950 199.950 514.050 202.050 ;
        RECT 515.400 201.600 516.600 206.400 ;
        RECT 517.950 206.400 526.050 207.600 ;
        RECT 517.950 205.950 520.050 206.400 ;
        RECT 523.950 205.950 526.050 206.400 ;
        RECT 622.950 207.600 625.050 208.050 ;
        RECT 631.950 207.600 634.050 208.050 ;
        RECT 622.950 206.400 634.050 207.600 ;
        RECT 622.950 205.950 625.050 206.400 ;
        RECT 631.950 205.950 634.050 206.400 ;
        RECT 634.950 207.600 637.050 208.050 ;
        RECT 673.950 207.600 676.050 208.050 ;
        RECT 634.950 206.400 676.050 207.600 ;
        RECT 634.950 205.950 637.050 206.400 ;
        RECT 673.950 205.950 676.050 206.400 ;
        RECT 520.950 204.600 523.050 205.050 ;
        RECT 535.950 204.600 538.050 205.050 ;
        RECT 520.950 203.400 538.050 204.600 ;
        RECT 520.950 202.950 523.050 203.400 ;
        RECT 535.950 202.950 538.050 203.400 ;
        RECT 580.950 204.600 583.050 205.050 ;
        RECT 625.950 204.600 628.050 205.050 ;
        RECT 580.950 203.400 628.050 204.600 ;
        RECT 580.950 202.950 583.050 203.400 ;
        RECT 520.950 201.600 523.050 202.050 ;
        RECT 515.400 200.400 523.050 201.600 ;
        RECT 520.950 199.950 523.050 200.400 ;
        RECT 529.950 199.950 532.050 202.050 ;
        RECT 538.950 199.950 541.050 202.050 ;
        RECT 559.950 201.600 562.050 202.050 ;
        RECT 554.400 200.400 562.050 201.600 ;
        RECT 325.950 198.600 328.050 199.050 ;
        RECT 337.950 198.600 340.050 199.050 ;
        RECT 325.950 197.400 340.050 198.600 ;
        RECT 325.950 196.950 328.050 197.400 ;
        RECT 337.950 196.950 340.050 197.400 ;
        RECT 364.950 198.600 367.050 199.050 ;
        RECT 379.950 198.600 382.050 199.050 ;
        RECT 364.950 197.400 382.050 198.600 ;
        RECT 364.950 196.950 367.050 197.400 ;
        RECT 379.950 196.950 382.050 197.400 ;
        RECT 385.950 198.600 388.050 199.050 ;
        RECT 397.950 198.600 400.050 199.050 ;
        RECT 436.950 198.600 439.050 199.050 ;
        RECT 457.950 198.600 460.050 199.050 ;
        RECT 385.950 197.400 400.050 198.600 ;
        RECT 385.950 196.950 388.050 197.400 ;
        RECT 397.950 196.950 400.050 197.400 ;
        RECT 401.400 197.400 439.050 198.600 ;
        RECT 319.950 195.600 322.050 196.050 ;
        RECT 314.400 194.400 322.050 195.600 ;
        RECT 286.950 193.950 289.050 194.400 ;
        RECT 304.950 193.950 307.050 194.400 ;
        RECT 319.950 193.950 322.050 194.400 ;
        RECT 328.950 195.600 331.050 196.050 ;
        RECT 340.950 195.600 343.050 196.050 ;
        RECT 328.950 194.400 343.050 195.600 ;
        RECT 328.950 193.950 331.050 194.400 ;
        RECT 340.950 193.950 343.050 194.400 ;
        RECT 361.950 195.600 364.050 196.050 ;
        RECT 373.950 195.600 376.050 196.050 ;
        RECT 361.950 194.400 376.050 195.600 ;
        RECT 361.950 193.950 364.050 194.400 ;
        RECT 373.950 193.950 376.050 194.400 ;
        RECT 388.950 195.600 391.050 196.050 ;
        RECT 401.400 195.600 402.600 197.400 ;
        RECT 436.950 196.950 439.050 197.400 ;
        RECT 443.400 197.400 460.050 198.600 ;
        RECT 388.950 194.400 402.600 195.600 ;
        RECT 415.950 195.600 418.050 196.050 ;
        RECT 443.400 195.600 444.600 197.400 ;
        RECT 457.950 196.950 460.050 197.400 ;
        RECT 463.950 198.600 466.050 199.050 ;
        RECT 469.950 198.600 472.050 199.050 ;
        RECT 475.950 198.600 478.050 199.050 ;
        RECT 463.950 197.400 472.050 198.600 ;
        RECT 463.950 196.950 466.050 197.400 ;
        RECT 469.950 196.950 472.050 197.400 ;
        RECT 473.400 197.400 478.050 198.600 ;
        RECT 415.950 194.400 444.600 195.600 ;
        RECT 388.950 193.950 391.050 194.400 ;
        RECT 415.950 193.950 418.050 194.400 ;
        RECT 214.950 192.600 217.050 193.050 ;
        RECT 212.400 191.400 217.050 192.600 ;
        RECT 145.950 190.950 148.050 191.400 ;
        RECT 163.950 190.950 166.050 191.400 ;
        RECT 196.950 190.950 199.050 191.400 ;
        RECT 214.950 190.950 217.050 191.400 ;
        RECT 280.950 192.600 283.050 193.050 ;
        RECT 286.950 192.600 289.050 193.050 ;
        RECT 280.950 191.400 289.050 192.600 ;
        RECT 280.950 190.950 283.050 191.400 ;
        RECT 286.950 190.950 289.050 191.400 ;
        RECT 313.950 192.600 316.050 193.050 ;
        RECT 319.950 192.600 322.050 193.050 ;
        RECT 343.950 192.600 346.050 193.050 ;
        RECT 313.950 191.400 346.050 192.600 ;
        RECT 313.950 190.950 316.050 191.400 ;
        RECT 319.950 190.950 322.050 191.400 ;
        RECT 343.950 190.950 346.050 191.400 ;
        RECT 352.950 192.600 355.050 193.050 ;
        RECT 367.950 192.600 370.050 193.050 ;
        RECT 352.950 191.400 370.050 192.600 ;
        RECT 352.950 190.950 355.050 191.400 ;
        RECT 367.950 190.950 370.050 191.400 ;
        RECT 370.950 192.600 373.050 193.050 ;
        RECT 382.950 192.600 385.050 193.050 ;
        RECT 370.950 191.400 385.050 192.600 ;
        RECT 370.950 190.950 373.050 191.400 ;
        RECT 382.950 190.950 385.050 191.400 ;
        RECT 397.950 192.600 400.050 193.050 ;
        RECT 403.950 192.600 406.050 193.050 ;
        RECT 397.950 191.400 406.050 192.600 ;
        RECT 443.400 192.600 444.600 194.400 ;
        RECT 445.950 195.600 448.050 196.050 ;
        RECT 454.950 195.600 457.050 196.050 ;
        RECT 445.950 194.400 457.050 195.600 ;
        RECT 445.950 193.950 448.050 194.400 ;
        RECT 454.950 193.950 457.050 194.400 ;
        RECT 466.950 195.600 469.050 196.050 ;
        RECT 473.400 195.600 474.600 197.400 ;
        RECT 475.950 196.950 478.050 197.400 ;
        RECT 478.950 198.600 481.050 199.050 ;
        RECT 508.950 198.600 511.050 199.050 ;
        RECT 478.950 197.400 511.050 198.600 ;
        RECT 478.950 196.950 481.050 197.400 ;
        RECT 508.950 196.950 511.050 197.400 ;
        RECT 530.400 196.050 531.600 199.950 ;
        RECT 484.950 195.600 487.050 196.050 ;
        RECT 490.950 195.600 493.050 196.050 ;
        RECT 466.950 194.400 474.600 195.600 ;
        RECT 479.400 194.400 493.050 195.600 ;
        RECT 466.950 193.950 469.050 194.400 ;
        RECT 445.950 192.600 448.050 193.050 ;
        RECT 443.400 191.400 448.050 192.600 ;
        RECT 397.950 190.950 400.050 191.400 ;
        RECT 403.950 190.950 406.050 191.400 ;
        RECT 445.950 190.950 448.050 191.400 ;
        RECT 451.950 192.600 454.050 193.050 ;
        RECT 463.950 192.600 466.050 193.050 ;
        RECT 451.950 191.400 466.050 192.600 ;
        RECT 451.950 190.950 454.050 191.400 ;
        RECT 463.950 190.950 466.050 191.400 ;
        RECT 28.950 189.600 31.050 190.050 ;
        RECT 79.950 189.600 82.050 190.050 ;
        RECT 91.950 189.600 94.050 190.050 ;
        RECT 28.950 188.400 94.050 189.600 ;
        RECT 28.950 187.950 31.050 188.400 ;
        RECT 79.950 187.950 82.050 188.400 ;
        RECT 91.950 187.950 94.050 188.400 ;
        RECT 94.950 189.600 97.050 190.050 ;
        RECT 109.950 189.600 112.050 190.050 ;
        RECT 94.950 188.400 112.050 189.600 ;
        RECT 94.950 187.950 97.050 188.400 ;
        RECT 109.950 187.950 112.050 188.400 ;
        RECT 112.950 189.600 115.050 190.050 ;
        RECT 118.950 189.600 121.050 190.050 ;
        RECT 112.950 188.400 121.050 189.600 ;
        RECT 112.950 187.950 115.050 188.400 ;
        RECT 118.950 187.950 121.050 188.400 ;
        RECT 133.950 189.600 136.050 190.050 ;
        RECT 148.950 189.600 151.050 190.050 ;
        RECT 133.950 188.400 151.050 189.600 ;
        RECT 133.950 187.950 136.050 188.400 ;
        RECT 148.950 187.950 151.050 188.400 ;
        RECT 166.950 189.600 169.050 190.050 ;
        RECT 193.950 189.600 196.050 190.050 ;
        RECT 166.950 188.400 196.050 189.600 ;
        RECT 166.950 187.950 169.050 188.400 ;
        RECT 193.950 187.950 196.050 188.400 ;
        RECT 346.950 189.600 349.050 190.050 ;
        RECT 355.950 189.600 358.050 190.050 ;
        RECT 346.950 188.400 358.050 189.600 ;
        RECT 346.950 187.950 349.050 188.400 ;
        RECT 355.950 187.950 358.050 188.400 ;
        RECT 364.950 189.600 367.050 190.050 ;
        RECT 370.950 189.600 373.050 190.050 ;
        RECT 364.950 188.400 373.050 189.600 ;
        RECT 364.950 187.950 367.050 188.400 ;
        RECT 370.950 187.950 373.050 188.400 ;
        RECT 409.950 189.600 412.050 190.050 ;
        RECT 424.950 189.600 427.050 190.050 ;
        RECT 409.950 188.400 427.050 189.600 ;
        RECT 409.950 187.950 412.050 188.400 ;
        RECT 424.950 187.950 427.050 188.400 ;
        RECT 451.950 189.600 454.050 190.050 ;
        RECT 479.400 189.600 480.600 194.400 ;
        RECT 484.950 193.950 487.050 194.400 ;
        RECT 490.950 193.950 493.050 194.400 ;
        RECT 505.950 195.600 508.050 196.050 ;
        RECT 514.950 195.600 517.050 196.050 ;
        RECT 505.950 194.400 517.050 195.600 ;
        RECT 505.950 193.950 508.050 194.400 ;
        RECT 514.950 193.950 517.050 194.400 ;
        RECT 529.950 193.950 532.050 196.050 ;
        RECT 481.950 192.600 484.050 193.050 ;
        RECT 490.950 192.600 493.050 193.050 ;
        RECT 481.950 191.400 493.050 192.600 ;
        RECT 481.950 190.950 484.050 191.400 ;
        RECT 490.950 190.950 493.050 191.400 ;
        RECT 499.950 192.600 502.050 193.050 ;
        RECT 511.950 192.600 514.050 193.050 ;
        RECT 499.950 191.400 514.050 192.600 ;
        RECT 499.950 190.950 502.050 191.400 ;
        RECT 511.950 190.950 514.050 191.400 ;
        RECT 514.950 192.600 517.050 193.050 ;
        RECT 539.400 192.600 540.600 199.950 ;
        RECT 544.950 196.950 547.050 199.050 ;
        RECT 545.400 193.050 546.600 196.950 ;
        RECT 554.400 195.600 555.600 200.400 ;
        RECT 559.950 199.950 562.050 200.400 ;
        RECT 565.950 201.600 568.050 202.050 ;
        RECT 580.950 201.600 583.050 202.050 ;
        RECT 565.950 200.400 583.050 201.600 ;
        RECT 565.950 199.950 568.050 200.400 ;
        RECT 580.950 199.950 583.050 200.400 ;
        RECT 616.950 199.950 619.050 202.050 ;
        RECT 556.950 198.600 559.050 199.050 ;
        RECT 562.950 198.600 565.050 199.050 ;
        RECT 556.950 197.400 565.050 198.600 ;
        RECT 556.950 196.950 559.050 197.400 ;
        RECT 562.950 196.950 565.050 197.400 ;
        RECT 568.950 198.600 571.050 199.050 ;
        RECT 598.950 198.600 601.050 199.050 ;
        RECT 568.950 197.400 601.050 198.600 ;
        RECT 568.950 196.950 571.050 197.400 ;
        RECT 598.950 196.950 601.050 197.400 ;
        RECT 617.400 196.050 618.600 199.950 ;
        RECT 620.400 199.050 621.600 203.400 ;
        RECT 625.950 202.950 628.050 203.400 ;
        RECT 733.950 204.600 736.050 205.050 ;
        RECT 787.950 204.600 790.050 205.050 ;
        RECT 733.950 203.400 790.050 204.600 ;
        RECT 733.950 202.950 736.050 203.400 ;
        RECT 787.950 202.950 790.050 203.400 ;
        RECT 853.950 204.600 856.050 205.050 ;
        RECT 859.950 204.600 862.050 205.050 ;
        RECT 853.950 203.400 862.050 204.600 ;
        RECT 853.950 202.950 856.050 203.400 ;
        RECT 859.950 202.950 862.050 203.400 ;
        RECT 634.950 201.600 637.050 202.050 ;
        RECT 623.400 200.400 637.050 201.600 ;
        RECT 619.950 196.950 622.050 199.050 ;
        RECT 562.950 195.600 565.050 196.050 ;
        RECT 554.400 194.400 565.050 195.600 ;
        RECT 562.950 193.950 565.050 194.400 ;
        RECT 616.950 193.950 619.050 196.050 ;
        RECT 619.950 195.600 622.050 196.050 ;
        RECT 623.400 195.600 624.600 200.400 ;
        RECT 634.950 199.950 637.050 200.400 ;
        RECT 640.950 201.600 643.050 202.050 ;
        RECT 661.950 201.600 664.050 202.050 ;
        RECT 676.950 201.600 679.050 202.050 ;
        RECT 640.950 200.400 645.600 201.600 ;
        RECT 640.950 199.950 643.050 200.400 ;
        RECT 625.950 198.600 628.050 199.050 ;
        RECT 631.950 198.600 634.050 199.050 ;
        RECT 625.950 197.400 634.050 198.600 ;
        RECT 625.950 196.950 628.050 197.400 ;
        RECT 631.950 196.950 634.050 197.400 ;
        RECT 634.950 198.600 637.050 199.050 ;
        RECT 640.950 198.600 643.050 199.050 ;
        RECT 634.950 197.400 643.050 198.600 ;
        RECT 634.950 196.950 637.050 197.400 ;
        RECT 640.950 196.950 643.050 197.400 ;
        RECT 644.400 196.050 645.600 200.400 ;
        RECT 661.950 200.400 679.050 201.600 ;
        RECT 661.950 199.950 664.050 200.400 ;
        RECT 676.950 199.950 679.050 200.400 ;
        RECT 712.950 201.600 715.050 202.050 ;
        RECT 736.950 201.600 739.050 202.050 ;
        RECT 712.950 200.400 739.050 201.600 ;
        RECT 712.950 199.950 715.050 200.400 ;
        RECT 736.950 199.950 739.050 200.400 ;
        RECT 778.950 201.600 781.050 202.050 ;
        RECT 811.950 201.600 814.050 202.050 ;
        RECT 778.950 200.400 814.050 201.600 ;
        RECT 778.950 199.950 781.050 200.400 ;
        RECT 811.950 199.950 814.050 200.400 ;
        RECT 847.950 201.600 850.050 202.050 ;
        RECT 853.950 201.600 856.050 202.050 ;
        RECT 847.950 200.400 856.050 201.600 ;
        RECT 847.950 199.950 850.050 200.400 ;
        RECT 853.950 199.950 856.050 200.400 ;
        RECT 646.950 198.600 649.050 199.050 ;
        RECT 652.950 198.600 655.050 199.050 ;
        RECT 646.950 197.400 655.050 198.600 ;
        RECT 646.950 196.950 649.050 197.400 ;
        RECT 652.950 196.950 655.050 197.400 ;
        RECT 664.950 196.950 667.050 199.050 ;
        RECT 679.950 198.600 682.050 199.050 ;
        RECT 668.400 197.400 682.050 198.600 ;
        RECT 619.950 194.400 624.600 195.600 ;
        RECT 619.950 193.950 622.050 194.400 ;
        RECT 643.950 193.950 646.050 196.050 ;
        RECT 652.950 195.600 655.050 196.050 ;
        RECT 661.950 195.600 664.050 196.050 ;
        RECT 652.950 194.400 664.050 195.600 ;
        RECT 652.950 193.950 655.050 194.400 ;
        RECT 661.950 193.950 664.050 194.400 ;
        RECT 665.400 193.050 666.600 196.950 ;
        RECT 668.400 196.050 669.600 197.400 ;
        RECT 679.950 196.950 682.050 197.400 ;
        RECT 718.950 198.600 721.050 199.050 ;
        RECT 727.950 198.600 730.050 199.050 ;
        RECT 745.950 198.600 748.050 199.050 ;
        RECT 718.950 197.400 748.050 198.600 ;
        RECT 718.950 196.950 721.050 197.400 ;
        RECT 727.950 196.950 730.050 197.400 ;
        RECT 745.950 196.950 748.050 197.400 ;
        RECT 751.950 198.600 754.050 199.050 ;
        RECT 760.950 198.600 763.050 199.050 ;
        RECT 751.950 197.400 763.050 198.600 ;
        RECT 751.950 196.950 754.050 197.400 ;
        RECT 760.950 196.950 763.050 197.400 ;
        RECT 826.950 198.600 829.050 199.050 ;
        RECT 859.950 198.600 862.050 199.050 ;
        RECT 826.950 197.400 862.050 198.600 ;
        RECT 826.950 196.950 829.050 197.400 ;
        RECT 859.950 196.950 862.050 197.400 ;
        RECT 667.950 195.600 670.050 196.050 ;
        RECT 709.950 195.600 712.050 196.050 ;
        RECT 715.950 195.600 718.050 196.050 ;
        RECT 667.950 194.400 718.050 195.600 ;
        RECT 667.950 193.950 670.050 194.400 ;
        RECT 709.950 193.950 712.050 194.400 ;
        RECT 715.950 193.950 718.050 194.400 ;
        RECT 733.950 195.600 736.050 196.050 ;
        RECT 739.950 195.600 742.050 196.050 ;
        RECT 733.950 194.400 742.050 195.600 ;
        RECT 733.950 193.950 736.050 194.400 ;
        RECT 739.950 193.950 742.050 194.400 ;
        RECT 742.950 195.600 745.050 196.050 ;
        RECT 757.950 195.600 760.050 196.050 ;
        RECT 742.950 194.400 760.050 195.600 ;
        RECT 742.950 193.950 745.050 194.400 ;
        RECT 757.950 193.950 760.050 194.400 ;
        RECT 763.950 195.600 766.050 196.050 ;
        RECT 769.950 195.600 772.050 196.050 ;
        RECT 763.950 194.400 772.050 195.600 ;
        RECT 763.950 193.950 766.050 194.400 ;
        RECT 769.950 193.950 772.050 194.400 ;
        RECT 784.950 195.600 787.050 196.050 ;
        RECT 838.950 195.600 841.050 196.050 ;
        RECT 784.950 194.400 841.050 195.600 ;
        RECT 784.950 193.950 787.050 194.400 ;
        RECT 838.950 193.950 841.050 194.400 ;
        RECT 850.950 195.600 853.050 196.050 ;
        RECT 859.950 195.600 862.050 196.050 ;
        RECT 850.950 194.400 862.050 195.600 ;
        RECT 850.950 193.950 853.050 194.400 ;
        RECT 859.950 193.950 862.050 194.400 ;
        RECT 514.950 191.400 540.600 192.600 ;
        RECT 514.950 190.950 517.050 191.400 ;
        RECT 544.950 190.950 547.050 193.050 ;
        RECT 664.950 190.950 667.050 193.050 ;
        RECT 694.950 192.600 697.050 193.050 ;
        RECT 703.950 192.600 706.050 193.050 ;
        RECT 694.950 191.400 706.050 192.600 ;
        RECT 694.950 190.950 697.050 191.400 ;
        RECT 703.950 190.950 706.050 191.400 ;
        RECT 712.950 192.600 715.050 193.050 ;
        RECT 724.950 192.600 727.050 193.050 ;
        RECT 712.950 191.400 727.050 192.600 ;
        RECT 712.950 190.950 715.050 191.400 ;
        RECT 724.950 190.950 727.050 191.400 ;
        RECT 730.950 192.600 733.050 193.050 ;
        RECT 745.950 192.600 748.050 193.050 ;
        RECT 730.950 191.400 748.050 192.600 ;
        RECT 730.950 190.950 733.050 191.400 ;
        RECT 745.950 190.950 748.050 191.400 ;
        RECT 754.950 192.600 757.050 193.050 ;
        RECT 796.950 192.600 799.050 193.050 ;
        RECT 754.950 191.400 799.050 192.600 ;
        RECT 754.950 190.950 757.050 191.400 ;
        RECT 796.950 190.950 799.050 191.400 ;
        RECT 808.950 192.600 811.050 193.050 ;
        RECT 814.950 192.600 817.050 193.050 ;
        RECT 808.950 191.400 817.050 192.600 ;
        RECT 808.950 190.950 811.050 191.400 ;
        RECT 814.950 190.950 817.050 191.400 ;
        RECT 451.950 188.400 480.600 189.600 ;
        RECT 481.950 189.600 484.050 190.050 ;
        RECT 520.950 189.600 523.050 190.050 ;
        RECT 601.950 189.600 604.050 190.050 ;
        RECT 607.950 189.600 610.050 190.050 ;
        RECT 481.950 188.400 610.050 189.600 ;
        RECT 451.950 187.950 454.050 188.400 ;
        RECT 481.950 187.950 484.050 188.400 ;
        RECT 520.950 187.950 523.050 188.400 ;
        RECT 601.950 187.950 604.050 188.400 ;
        RECT 607.950 187.950 610.050 188.400 ;
        RECT 622.950 189.600 625.050 190.050 ;
        RECT 658.950 189.600 661.050 190.050 ;
        RECT 622.950 188.400 661.050 189.600 ;
        RECT 622.950 187.950 625.050 188.400 ;
        RECT 658.950 187.950 661.050 188.400 ;
        RECT 697.950 189.600 700.050 190.050 ;
        RECT 724.950 189.600 727.050 190.050 ;
        RECT 697.950 188.400 727.050 189.600 ;
        RECT 697.950 187.950 700.050 188.400 ;
        RECT 724.950 187.950 727.050 188.400 ;
        RECT 796.950 189.600 799.050 190.050 ;
        RECT 844.950 189.600 847.050 190.050 ;
        RECT 796.950 188.400 847.050 189.600 ;
        RECT 796.950 187.950 799.050 188.400 ;
        RECT 844.950 187.950 847.050 188.400 ;
        RECT 58.950 186.600 61.050 187.050 ;
        RECT 70.950 186.600 73.050 187.050 ;
        RECT 58.950 185.400 73.050 186.600 ;
        RECT 58.950 184.950 61.050 185.400 ;
        RECT 70.950 184.950 73.050 185.400 ;
        RECT 91.950 186.600 94.050 187.050 ;
        RECT 148.950 186.600 151.050 187.050 ;
        RECT 202.950 186.600 205.050 187.050 ;
        RECT 91.950 185.400 147.600 186.600 ;
        RECT 91.950 184.950 94.050 185.400 ;
        RECT 25.950 183.600 28.050 184.050 ;
        RECT 64.950 183.600 67.050 184.050 ;
        RECT 94.950 183.600 97.050 184.050 ;
        RECT 25.950 182.400 97.050 183.600 ;
        RECT 25.950 181.950 28.050 182.400 ;
        RECT 64.950 181.950 67.050 182.400 ;
        RECT 94.950 181.950 97.050 182.400 ;
        RECT 100.950 183.600 103.050 184.050 ;
        RECT 112.950 183.600 115.050 184.050 ;
        RECT 100.950 182.400 115.050 183.600 ;
        RECT 100.950 181.950 103.050 182.400 ;
        RECT 112.950 181.950 115.050 182.400 ;
        RECT 121.950 183.600 124.050 184.050 ;
        RECT 136.950 183.600 139.050 184.050 ;
        RECT 121.950 182.400 139.050 183.600 ;
        RECT 146.400 183.600 147.600 185.400 ;
        RECT 148.950 185.400 205.050 186.600 ;
        RECT 148.950 184.950 151.050 185.400 ;
        RECT 202.950 184.950 205.050 185.400 ;
        RECT 223.950 186.600 226.050 187.050 ;
        RECT 376.950 186.600 379.050 187.050 ;
        RECT 223.950 185.400 379.050 186.600 ;
        RECT 223.950 184.950 226.050 185.400 ;
        RECT 376.950 184.950 379.050 185.400 ;
        RECT 391.950 186.600 394.050 187.050 ;
        RECT 406.950 186.600 409.050 187.050 ;
        RECT 418.950 186.600 421.050 187.050 ;
        RECT 427.950 186.600 430.050 187.050 ;
        RECT 391.950 185.400 430.050 186.600 ;
        RECT 391.950 184.950 394.050 185.400 ;
        RECT 406.950 184.950 409.050 185.400 ;
        RECT 418.950 184.950 421.050 185.400 ;
        RECT 427.950 184.950 430.050 185.400 ;
        RECT 439.950 186.600 442.050 187.050 ;
        RECT 469.950 186.600 472.050 187.050 ;
        RECT 472.950 186.600 475.050 187.050 ;
        RECT 439.950 185.400 475.050 186.600 ;
        RECT 439.950 184.950 442.050 185.400 ;
        RECT 469.950 184.950 472.050 185.400 ;
        RECT 472.950 184.950 475.050 185.400 ;
        RECT 487.950 186.600 490.050 187.050 ;
        RECT 496.950 186.600 499.050 187.050 ;
        RECT 487.950 185.400 499.050 186.600 ;
        RECT 487.950 184.950 490.050 185.400 ;
        RECT 496.950 184.950 499.050 185.400 ;
        RECT 538.950 186.600 541.050 187.050 ;
        RECT 571.950 186.600 574.050 187.050 ;
        RECT 538.950 185.400 574.050 186.600 ;
        RECT 538.950 184.950 541.050 185.400 ;
        RECT 571.950 184.950 574.050 185.400 ;
        RECT 589.950 186.600 592.050 187.050 ;
        RECT 634.950 186.600 637.050 187.050 ;
        RECT 589.950 185.400 637.050 186.600 ;
        RECT 589.950 184.950 592.050 185.400 ;
        RECT 634.950 184.950 637.050 185.400 ;
        RECT 664.950 186.600 667.050 187.050 ;
        RECT 685.950 186.600 688.050 187.050 ;
        RECT 664.950 185.400 688.050 186.600 ;
        RECT 664.950 184.950 667.050 185.400 ;
        RECT 685.950 184.950 688.050 185.400 ;
        RECT 691.950 186.600 694.050 187.050 ;
        RECT 760.950 186.600 763.050 187.050 ;
        RECT 691.950 185.400 763.050 186.600 ;
        RECT 691.950 184.950 694.050 185.400 ;
        RECT 760.950 184.950 763.050 185.400 ;
        RECT 799.950 186.600 802.050 187.050 ;
        RECT 811.950 186.600 814.050 187.050 ;
        RECT 799.950 185.400 814.050 186.600 ;
        RECT 799.950 184.950 802.050 185.400 ;
        RECT 811.950 184.950 814.050 185.400 ;
        RECT 172.950 183.600 175.050 184.050 ;
        RECT 146.400 182.400 175.050 183.600 ;
        RECT 121.950 181.950 124.050 182.400 ;
        RECT 136.950 181.950 139.050 182.400 ;
        RECT 172.950 181.950 175.050 182.400 ;
        RECT 208.950 183.600 211.050 184.050 ;
        RECT 304.950 183.600 307.050 184.050 ;
        RECT 208.950 182.400 307.050 183.600 ;
        RECT 208.950 181.950 211.050 182.400 ;
        RECT 304.950 181.950 307.050 182.400 ;
        RECT 403.950 183.600 406.050 184.050 ;
        RECT 421.950 183.600 424.050 184.050 ;
        RECT 403.950 182.400 424.050 183.600 ;
        RECT 403.950 181.950 406.050 182.400 ;
        RECT 421.950 181.950 424.050 182.400 ;
        RECT 484.950 183.600 487.050 184.050 ;
        RECT 508.950 183.600 511.050 184.050 ;
        RECT 484.950 182.400 511.050 183.600 ;
        RECT 484.950 181.950 487.050 182.400 ;
        RECT 508.950 181.950 511.050 182.400 ;
        RECT 526.950 183.600 529.050 184.050 ;
        RECT 532.950 183.600 535.050 184.050 ;
        RECT 526.950 182.400 535.050 183.600 ;
        RECT 526.950 181.950 529.050 182.400 ;
        RECT 532.950 181.950 535.050 182.400 ;
        RECT 538.950 183.600 541.050 184.050 ;
        RECT 544.950 183.600 547.050 184.050 ;
        RECT 568.950 183.600 571.050 184.050 ;
        RECT 538.950 182.400 571.050 183.600 ;
        RECT 538.950 181.950 541.050 182.400 ;
        RECT 544.950 181.950 547.050 182.400 ;
        RECT 568.950 181.950 571.050 182.400 ;
        RECT 571.950 183.600 574.050 184.050 ;
        RECT 619.950 183.600 622.050 184.050 ;
        RECT 571.950 182.400 622.050 183.600 ;
        RECT 571.950 181.950 574.050 182.400 ;
        RECT 619.950 181.950 622.050 182.400 ;
        RECT 676.950 183.600 679.050 184.050 ;
        RECT 703.950 183.600 706.050 184.050 ;
        RECT 676.950 182.400 706.050 183.600 ;
        RECT 676.950 181.950 679.050 182.400 ;
        RECT 703.950 181.950 706.050 182.400 ;
        RECT 751.950 183.600 754.050 184.050 ;
        RECT 754.950 183.600 757.050 184.050 ;
        RECT 775.950 183.600 778.050 184.050 ;
        RECT 751.950 182.400 778.050 183.600 ;
        RECT 751.950 181.950 754.050 182.400 ;
        RECT 754.950 181.950 757.050 182.400 ;
        RECT 775.950 181.950 778.050 182.400 ;
        RECT 793.950 183.600 796.050 184.050 ;
        RECT 862.950 183.600 865.050 184.050 ;
        RECT 793.950 182.400 865.050 183.600 ;
        RECT 793.950 181.950 796.050 182.400 ;
        RECT 862.950 181.950 865.050 182.400 ;
        RECT 85.950 180.600 88.050 181.050 ;
        RECT 163.950 180.600 166.050 181.050 ;
        RECT 211.950 180.600 214.050 181.050 ;
        RECT 85.950 179.400 166.050 180.600 ;
        RECT 85.950 178.950 88.050 179.400 ;
        RECT 163.950 178.950 166.050 179.400 ;
        RECT 176.400 179.400 214.050 180.600 ;
        RECT 46.950 177.600 49.050 178.050 ;
        RECT 176.400 177.600 177.600 179.400 ;
        RECT 211.950 178.950 214.050 179.400 ;
        RECT 265.950 180.600 268.050 181.050 ;
        RECT 595.950 180.600 598.050 181.050 ;
        RECT 676.950 180.600 679.050 181.050 ;
        RECT 265.950 179.400 679.050 180.600 ;
        RECT 265.950 178.950 268.050 179.400 ;
        RECT 595.950 178.950 598.050 179.400 ;
        RECT 676.950 178.950 679.050 179.400 ;
        RECT 721.950 180.600 724.050 181.050 ;
        RECT 772.950 180.600 775.050 181.050 ;
        RECT 817.950 180.600 820.050 181.050 ;
        RECT 829.950 180.600 832.050 181.050 ;
        RECT 721.950 179.400 771.600 180.600 ;
        RECT 721.950 178.950 724.050 179.400 ;
        RECT 46.950 176.400 177.600 177.600 ;
        RECT 178.950 177.600 181.050 178.050 ;
        RECT 226.950 177.600 229.050 178.050 ;
        RECT 232.950 177.600 235.050 178.050 ;
        RECT 178.950 176.400 235.050 177.600 ;
        RECT 46.950 175.950 49.050 176.400 ;
        RECT 178.950 175.950 181.050 176.400 ;
        RECT 226.950 175.950 229.050 176.400 ;
        RECT 232.950 175.950 235.050 176.400 ;
        RECT 265.950 177.600 268.050 178.050 ;
        RECT 271.950 177.600 274.050 178.050 ;
        RECT 265.950 176.400 274.050 177.600 ;
        RECT 265.950 175.950 268.050 176.400 ;
        RECT 271.950 175.950 274.050 176.400 ;
        RECT 298.950 177.600 301.050 178.050 ;
        RECT 355.950 177.600 358.050 178.050 ;
        RECT 298.950 176.400 358.050 177.600 ;
        RECT 298.950 175.950 301.050 176.400 ;
        RECT 355.950 175.950 358.050 176.400 ;
        RECT 400.950 177.600 403.050 178.050 ;
        RECT 415.950 177.600 418.050 178.050 ;
        RECT 400.950 176.400 418.050 177.600 ;
        RECT 400.950 175.950 403.050 176.400 ;
        RECT 415.950 175.950 418.050 176.400 ;
        RECT 418.950 177.600 421.050 178.050 ;
        RECT 433.950 177.600 436.050 178.050 ;
        RECT 418.950 176.400 436.050 177.600 ;
        RECT 418.950 175.950 421.050 176.400 ;
        RECT 433.950 175.950 436.050 176.400 ;
        RECT 475.950 177.600 478.050 178.050 ;
        RECT 505.950 177.600 508.050 178.050 ;
        RECT 475.950 176.400 508.050 177.600 ;
        RECT 475.950 175.950 478.050 176.400 ;
        RECT 505.950 175.950 508.050 176.400 ;
        RECT 520.950 177.600 523.050 178.050 ;
        RECT 526.950 177.600 529.050 178.050 ;
        RECT 520.950 176.400 529.050 177.600 ;
        RECT 520.950 175.950 523.050 176.400 ;
        RECT 526.950 175.950 529.050 176.400 ;
        RECT 541.950 177.600 544.050 178.050 ;
        RECT 571.950 177.600 574.050 178.050 ;
        RECT 541.950 176.400 574.050 177.600 ;
        RECT 541.950 175.950 544.050 176.400 ;
        RECT 571.950 175.950 574.050 176.400 ;
        RECT 589.950 177.600 592.050 178.050 ;
        RECT 613.950 177.600 616.050 178.050 ;
        RECT 589.950 176.400 616.050 177.600 ;
        RECT 589.950 175.950 592.050 176.400 ;
        RECT 613.950 175.950 616.050 176.400 ;
        RECT 700.950 177.600 703.050 178.050 ;
        RECT 721.950 177.600 724.050 178.050 ;
        RECT 700.950 176.400 724.050 177.600 ;
        RECT 770.400 177.600 771.600 179.400 ;
        RECT 772.950 179.400 832.050 180.600 ;
        RECT 772.950 178.950 775.050 179.400 ;
        RECT 817.950 178.950 820.050 179.400 ;
        RECT 829.950 178.950 832.050 179.400 ;
        RECT 817.950 177.600 820.050 178.050 ;
        RECT 770.400 176.400 820.050 177.600 ;
        RECT 700.950 175.950 703.050 176.400 ;
        RECT 721.950 175.950 724.050 176.400 ;
        RECT 817.950 175.950 820.050 176.400 ;
        RECT 31.950 174.600 34.050 175.050 ;
        RECT 91.950 174.600 94.050 175.050 ;
        RECT 106.950 174.600 109.050 175.050 ;
        RECT 31.950 173.400 109.050 174.600 ;
        RECT 31.950 172.950 34.050 173.400 ;
        RECT 91.950 172.950 94.050 173.400 ;
        RECT 106.950 172.950 109.050 173.400 ;
        RECT 160.950 174.600 163.050 175.050 ;
        RECT 190.950 174.600 193.050 175.050 ;
        RECT 244.950 174.600 247.050 175.050 ;
        RECT 160.950 173.400 247.050 174.600 ;
        RECT 160.950 172.950 163.050 173.400 ;
        RECT 190.950 172.950 193.050 173.400 ;
        RECT 244.950 172.950 247.050 173.400 ;
        RECT 250.950 174.600 253.050 175.050 ;
        RECT 409.950 174.600 412.050 175.050 ;
        RECT 250.950 173.400 412.050 174.600 ;
        RECT 250.950 172.950 253.050 173.400 ;
        RECT 409.950 172.950 412.050 173.400 ;
        RECT 424.950 174.600 427.050 175.050 ;
        RECT 439.950 174.600 442.050 175.050 ;
        RECT 424.950 173.400 442.050 174.600 ;
        RECT 424.950 172.950 427.050 173.400 ;
        RECT 439.950 172.950 442.050 173.400 ;
        RECT 457.950 174.600 460.050 175.050 ;
        RECT 469.950 174.600 472.050 175.050 ;
        RECT 457.950 173.400 472.050 174.600 ;
        RECT 457.950 172.950 460.050 173.400 ;
        RECT 469.950 172.950 472.050 173.400 ;
        RECT 478.950 174.600 481.050 175.050 ;
        RECT 502.950 174.600 505.050 175.050 ;
        RECT 478.950 173.400 505.050 174.600 ;
        RECT 478.950 172.950 481.050 173.400 ;
        RECT 502.950 172.950 505.050 173.400 ;
        RECT 505.950 174.600 508.050 175.050 ;
        RECT 565.950 174.600 568.050 175.050 ;
        RECT 598.950 174.600 601.050 175.050 ;
        RECT 505.950 173.400 568.050 174.600 ;
        RECT 505.950 172.950 508.050 173.400 ;
        RECT 565.950 172.950 568.050 173.400 ;
        RECT 590.400 173.400 601.050 174.600 ;
        RECT 22.950 171.600 25.050 172.050 ;
        RECT 40.950 171.600 43.050 172.050 ;
        RECT 22.950 170.400 43.050 171.600 ;
        RECT 22.950 169.950 25.050 170.400 ;
        RECT 40.950 169.950 43.050 170.400 ;
        RECT 43.950 171.600 46.050 172.050 ;
        RECT 49.950 171.600 52.050 172.050 ;
        RECT 43.950 170.400 52.050 171.600 ;
        RECT 43.950 169.950 46.050 170.400 ;
        RECT 49.950 169.950 52.050 170.400 ;
        RECT 61.950 171.600 64.050 172.050 ;
        RECT 67.950 171.600 70.050 172.050 ;
        RECT 73.950 171.600 76.050 172.050 ;
        RECT 61.950 170.400 70.050 171.600 ;
        RECT 61.950 169.950 64.050 170.400 ;
        RECT 67.950 169.950 70.050 170.400 ;
        RECT 71.400 170.400 76.050 171.600 ;
        RECT 7.950 168.600 10.050 169.050 ;
        RECT 16.950 168.600 19.050 169.050 ;
        RECT 7.950 167.400 19.050 168.600 ;
        RECT 7.950 166.950 10.050 167.400 ;
        RECT 16.950 166.950 19.050 167.400 ;
        RECT 10.950 165.600 13.050 166.050 ;
        RECT 28.950 165.600 31.050 166.050 ;
        RECT 10.950 164.400 31.050 165.600 ;
        RECT 10.950 163.950 13.050 164.400 ;
        RECT 28.950 163.950 31.050 164.400 ;
        RECT 31.950 165.600 34.050 166.050 ;
        RECT 37.950 165.600 40.050 166.050 ;
        RECT 31.950 164.400 40.050 165.600 ;
        RECT 31.950 163.950 34.050 164.400 ;
        RECT 37.950 163.950 40.050 164.400 ;
        RECT 40.950 165.600 43.050 166.050 ;
        RECT 67.950 165.600 70.050 166.050 ;
        RECT 40.950 164.400 70.050 165.600 ;
        RECT 40.950 163.950 43.050 164.400 ;
        RECT 67.950 163.950 70.050 164.400 ;
        RECT 64.950 162.600 67.050 163.050 ;
        RECT 64.950 161.400 69.600 162.600 ;
        RECT 64.950 160.950 67.050 161.400 ;
        RECT 68.400 160.050 69.600 161.400 ;
        RECT 19.950 159.600 22.050 160.050 ;
        RECT 61.950 159.600 64.050 160.050 ;
        RECT 19.950 158.400 64.050 159.600 ;
        RECT 19.950 157.950 22.050 158.400 ;
        RECT 61.950 157.950 64.050 158.400 ;
        RECT 67.950 157.950 70.050 160.050 ;
        RECT 71.400 159.600 72.600 170.400 ;
        RECT 73.950 169.950 76.050 170.400 ;
        RECT 79.950 171.600 82.050 172.050 ;
        RECT 88.950 171.600 91.050 172.050 ;
        RECT 79.950 170.400 91.050 171.600 ;
        RECT 79.950 169.950 82.050 170.400 ;
        RECT 88.950 169.950 91.050 170.400 ;
        RECT 97.950 171.600 100.050 172.050 ;
        RECT 142.950 171.600 145.050 172.050 ;
        RECT 97.950 170.400 145.050 171.600 ;
        RECT 97.950 169.950 100.050 170.400 ;
        RECT 142.950 169.950 145.050 170.400 ;
        RECT 145.950 171.600 148.050 172.050 ;
        RECT 154.950 171.600 157.050 172.050 ;
        RECT 145.950 170.400 157.050 171.600 ;
        RECT 145.950 169.950 148.050 170.400 ;
        RECT 154.950 169.950 157.050 170.400 ;
        RECT 175.950 169.950 178.050 172.050 ;
        RECT 205.950 171.600 208.050 172.050 ;
        RECT 238.950 171.600 241.050 172.050 ;
        RECT 205.950 170.400 241.050 171.600 ;
        RECT 205.950 169.950 208.050 170.400 ;
        RECT 238.950 169.950 241.050 170.400 ;
        RECT 259.950 171.600 262.050 172.050 ;
        RECT 283.950 171.600 286.050 172.050 ;
        RECT 259.950 170.400 286.050 171.600 ;
        RECT 259.950 169.950 262.050 170.400 ;
        RECT 283.950 169.950 286.050 170.400 ;
        RECT 298.950 171.600 301.050 172.050 ;
        RECT 310.950 171.600 313.050 172.050 ;
        RECT 298.950 170.400 313.050 171.600 ;
        RECT 298.950 169.950 301.050 170.400 ;
        RECT 310.950 169.950 313.050 170.400 ;
        RECT 334.950 171.600 337.050 172.050 ;
        RECT 340.950 171.600 343.050 172.050 ;
        RECT 334.950 170.400 343.050 171.600 ;
        RECT 334.950 169.950 337.050 170.400 ;
        RECT 340.950 169.950 343.050 170.400 ;
        RECT 379.950 171.600 382.050 172.050 ;
        RECT 406.950 171.600 409.050 172.050 ;
        RECT 451.950 171.600 454.050 172.050 ;
        RECT 379.950 170.400 409.050 171.600 ;
        RECT 379.950 169.950 382.050 170.400 ;
        RECT 406.950 169.950 409.050 170.400 ;
        RECT 410.400 170.400 454.050 171.600 ;
        RECT 73.950 166.950 76.050 169.050 ;
        RECT 77.400 167.400 105.600 168.600 ;
        RECT 74.400 163.050 75.600 166.950 ;
        RECT 77.400 166.050 78.600 167.400 ;
        RECT 104.400 166.050 105.600 167.400 ;
        RECT 76.950 163.950 79.050 166.050 ;
        RECT 82.950 165.600 85.050 166.050 ;
        RECT 97.950 165.600 100.050 166.050 ;
        RECT 82.950 164.400 100.050 165.600 ;
        RECT 82.950 163.950 85.050 164.400 ;
        RECT 97.950 163.950 100.050 164.400 ;
        RECT 103.950 163.950 106.050 166.050 ;
        RECT 109.950 165.600 112.050 166.050 ;
        RECT 127.950 165.600 130.050 166.050 ;
        RECT 107.400 164.400 112.050 165.600 ;
        RECT 73.950 160.950 76.050 163.050 ;
        RECT 79.950 162.600 82.050 163.050 ;
        RECT 88.950 162.600 91.050 163.050 ;
        RECT 100.950 162.600 103.050 163.050 ;
        RECT 79.950 161.400 103.050 162.600 ;
        RECT 79.950 160.950 82.050 161.400 ;
        RECT 88.950 160.950 91.050 161.400 ;
        RECT 100.950 160.950 103.050 161.400 ;
        RECT 104.400 160.050 105.600 163.950 ;
        RECT 107.400 160.050 108.600 164.400 ;
        RECT 109.950 163.950 112.050 164.400 ;
        RECT 122.400 164.400 130.050 165.600 ;
        RECT 109.950 160.950 112.050 163.050 ;
        RECT 76.950 159.600 79.050 160.050 ;
        RECT 71.400 158.400 79.050 159.600 ;
        RECT 76.950 157.950 79.050 158.400 ;
        RECT 103.950 157.950 106.050 160.050 ;
        RECT 106.950 157.950 109.050 160.050 ;
        RECT 110.400 159.600 111.600 160.950 ;
        RECT 112.950 159.600 115.050 160.050 ;
        RECT 110.400 158.400 115.050 159.600 ;
        RECT 122.400 159.600 123.600 164.400 ;
        RECT 127.950 163.950 130.050 164.400 ;
        RECT 136.950 165.600 139.050 166.050 ;
        RECT 166.950 165.600 169.050 166.050 ;
        RECT 136.950 164.400 169.050 165.600 ;
        RECT 176.400 165.600 177.600 169.950 ;
        RECT 178.950 168.600 181.050 169.050 ;
        RECT 184.950 168.600 187.050 169.050 ;
        RECT 202.950 168.600 205.050 169.050 ;
        RECT 178.950 167.400 183.600 168.600 ;
        RECT 178.950 166.950 181.050 167.400 ;
        RECT 182.400 165.600 183.600 167.400 ;
        RECT 184.950 167.400 205.050 168.600 ;
        RECT 184.950 166.950 187.050 167.400 ;
        RECT 202.950 166.950 205.050 167.400 ;
        RECT 220.950 166.950 223.050 169.050 ;
        RECT 241.950 168.600 244.050 169.050 ;
        RECT 262.950 168.600 265.050 169.050 ;
        RECT 241.950 167.400 265.050 168.600 ;
        RECT 241.950 166.950 244.050 167.400 ;
        RECT 262.950 166.950 265.050 167.400 ;
        RECT 268.950 168.600 271.050 169.050 ;
        RECT 277.950 168.600 280.050 169.050 ;
        RECT 268.950 167.400 280.050 168.600 ;
        RECT 268.950 166.950 271.050 167.400 ;
        RECT 277.950 166.950 280.050 167.400 ;
        RECT 310.950 168.600 313.050 169.050 ;
        RECT 316.950 168.600 319.050 169.050 ;
        RECT 349.950 168.600 352.050 169.050 ;
        RECT 367.950 168.600 370.050 169.050 ;
        RECT 410.400 168.600 411.600 170.400 ;
        RECT 451.950 169.950 454.050 170.400 ;
        RECT 454.950 171.600 457.050 172.050 ;
        RECT 472.950 171.600 475.050 172.050 ;
        RECT 496.950 171.600 499.050 172.050 ;
        RECT 590.400 171.600 591.600 173.400 ;
        RECT 598.950 172.950 601.050 173.400 ;
        RECT 604.950 174.600 607.050 175.050 ;
        RECT 607.950 174.600 610.050 175.050 ;
        RECT 619.950 174.600 622.050 175.050 ;
        RECT 604.950 173.400 622.050 174.600 ;
        RECT 604.950 172.950 607.050 173.400 ;
        RECT 607.950 172.950 610.050 173.400 ;
        RECT 619.950 172.950 622.050 173.400 ;
        RECT 631.950 174.600 634.050 175.050 ;
        RECT 661.950 174.600 664.050 175.050 ;
        RECT 730.950 174.600 733.050 175.050 ;
        RECT 757.950 174.600 760.050 175.050 ;
        RECT 631.950 173.400 760.050 174.600 ;
        RECT 631.950 172.950 634.050 173.400 ;
        RECT 661.950 172.950 664.050 173.400 ;
        RECT 730.950 172.950 733.050 173.400 ;
        RECT 757.950 172.950 760.050 173.400 ;
        RECT 763.950 174.600 766.050 175.050 ;
        RECT 772.950 174.600 775.050 175.050 ;
        RECT 763.950 173.400 775.050 174.600 ;
        RECT 763.950 172.950 766.050 173.400 ;
        RECT 772.950 172.950 775.050 173.400 ;
        RECT 781.950 174.600 784.050 175.050 ;
        RECT 787.950 174.600 790.050 175.050 ;
        RECT 781.950 173.400 790.050 174.600 ;
        RECT 781.950 172.950 784.050 173.400 ;
        RECT 787.950 172.950 790.050 173.400 ;
        RECT 454.950 170.400 468.600 171.600 ;
        RECT 454.950 169.950 457.050 170.400 ;
        RECT 310.950 167.400 319.050 168.600 ;
        RECT 310.950 166.950 313.050 167.400 ;
        RECT 316.950 166.950 319.050 167.400 ;
        RECT 320.400 167.400 411.600 168.600 ;
        RECT 412.950 168.600 415.050 169.050 ;
        RECT 424.950 168.600 427.050 169.050 ;
        RECT 412.950 167.400 427.050 168.600 ;
        RECT 193.950 165.600 196.050 166.050 ;
        RECT 176.400 164.400 180.600 165.600 ;
        RECT 182.400 164.400 196.050 165.600 ;
        RECT 136.950 163.950 139.050 164.400 ;
        RECT 166.950 163.950 169.050 164.400 ;
        RECT 179.400 163.050 180.600 164.400 ;
        RECT 193.950 163.950 196.050 164.400 ;
        RECT 205.950 165.600 208.050 166.050 ;
        RECT 221.400 165.600 222.600 166.950 ;
        RECT 205.950 164.400 222.600 165.600 ;
        RECT 277.950 165.600 280.050 166.050 ;
        RECT 295.950 165.600 298.050 166.050 ;
        RECT 301.950 165.600 304.050 166.050 ;
        RECT 316.950 165.600 319.050 166.050 ;
        RECT 277.950 164.400 298.050 165.600 ;
        RECT 205.950 163.950 208.050 164.400 ;
        RECT 277.950 163.950 280.050 164.400 ;
        RECT 295.950 163.950 298.050 164.400 ;
        RECT 299.400 164.400 319.050 165.600 ;
        RECT 124.950 162.600 127.050 163.050 ;
        RECT 139.950 162.600 142.050 163.050 ;
        RECT 124.950 161.400 142.050 162.600 ;
        RECT 124.950 160.950 127.050 161.400 ;
        RECT 139.950 160.950 142.050 161.400 ;
        RECT 145.950 162.600 148.050 163.050 ;
        RECT 151.950 162.600 154.050 163.050 ;
        RECT 145.950 161.400 154.050 162.600 ;
        RECT 145.950 160.950 148.050 161.400 ;
        RECT 151.950 160.950 154.050 161.400 ;
        RECT 157.950 162.600 160.050 163.050 ;
        RECT 163.950 162.600 166.050 163.050 ;
        RECT 157.950 161.400 166.050 162.600 ;
        RECT 157.950 160.950 160.050 161.400 ;
        RECT 163.950 160.950 166.050 161.400 ;
        RECT 178.950 160.950 181.050 163.050 ;
        RECT 184.950 162.600 187.050 163.050 ;
        RECT 193.950 162.600 196.050 163.050 ;
        RECT 184.950 161.400 196.050 162.600 ;
        RECT 184.950 160.950 187.050 161.400 ;
        RECT 193.950 160.950 196.050 161.400 ;
        RECT 235.950 162.600 238.050 163.050 ;
        RECT 253.950 162.600 256.050 163.050 ;
        RECT 235.950 161.400 256.050 162.600 ;
        RECT 235.950 160.950 238.050 161.400 ;
        RECT 253.950 160.950 256.050 161.400 ;
        RECT 280.950 162.600 283.050 163.050 ;
        RECT 299.400 162.600 300.600 164.400 ;
        RECT 301.950 163.950 304.050 164.400 ;
        RECT 316.950 163.950 319.050 164.400 ;
        RECT 280.950 161.400 300.600 162.600 ;
        RECT 313.950 162.600 316.050 163.050 ;
        RECT 320.400 162.600 321.600 167.400 ;
        RECT 349.950 166.950 352.050 167.400 ;
        RECT 367.950 166.950 370.050 167.400 ;
        RECT 412.950 166.950 415.050 167.400 ;
        RECT 424.950 166.950 427.050 167.400 ;
        RECT 439.950 168.600 442.050 169.050 ;
        RECT 451.950 168.600 454.050 169.050 ;
        RECT 439.950 167.400 454.050 168.600 ;
        RECT 439.950 166.950 442.050 167.400 ;
        RECT 451.950 166.950 454.050 167.400 ;
        RECT 331.950 165.600 334.050 166.050 ;
        RECT 349.950 165.600 352.050 166.050 ;
        RECT 331.950 164.400 352.050 165.600 ;
        RECT 331.950 163.950 334.050 164.400 ;
        RECT 349.950 163.950 352.050 164.400 ;
        RECT 361.950 165.600 364.050 166.050 ;
        RECT 391.950 165.600 394.050 166.050 ;
        RECT 361.950 164.400 394.050 165.600 ;
        RECT 361.950 163.950 364.050 164.400 ;
        RECT 391.950 163.950 394.050 164.400 ;
        RECT 406.950 165.600 409.050 166.050 ;
        RECT 454.950 165.600 457.050 166.050 ;
        RECT 406.950 164.400 457.050 165.600 ;
        RECT 406.950 163.950 409.050 164.400 ;
        RECT 454.950 163.950 457.050 164.400 ;
        RECT 313.950 161.400 321.600 162.600 ;
        RECT 334.950 162.600 337.050 163.050 ;
        RECT 358.950 162.600 361.050 163.050 ;
        RECT 334.950 161.400 361.050 162.600 ;
        RECT 280.950 160.950 283.050 161.400 ;
        RECT 313.950 160.950 316.050 161.400 ;
        RECT 334.950 160.950 337.050 161.400 ;
        RECT 358.950 160.950 361.050 161.400 ;
        RECT 364.950 160.950 367.050 163.050 ;
        RECT 388.950 162.600 391.050 163.050 ;
        RECT 403.950 162.600 406.050 163.050 ;
        RECT 388.950 161.400 406.050 162.600 ;
        RECT 388.950 160.950 391.050 161.400 ;
        RECT 403.950 160.950 406.050 161.400 ;
        RECT 412.950 162.600 415.050 163.050 ;
        RECT 436.950 162.600 439.050 163.050 ;
        RECT 412.950 161.400 439.050 162.600 ;
        RECT 412.950 160.950 415.050 161.400 ;
        RECT 436.950 160.950 439.050 161.400 ;
        RECT 442.950 162.600 445.050 163.050 ;
        RECT 467.400 162.600 468.600 170.400 ;
        RECT 472.950 170.400 499.050 171.600 ;
        RECT 472.950 169.950 475.050 170.400 ;
        RECT 496.950 169.950 499.050 170.400 ;
        RECT 569.400 170.400 591.600 171.600 ;
        RECT 598.950 171.600 601.050 172.050 ;
        RECT 604.950 171.600 607.050 172.050 ;
        RECT 598.950 170.400 607.050 171.600 ;
        RECT 475.950 168.600 478.050 169.050 ;
        RECT 487.950 168.600 490.050 169.050 ;
        RECT 475.950 167.400 490.050 168.600 ;
        RECT 475.950 166.950 478.050 167.400 ;
        RECT 487.950 166.950 490.050 167.400 ;
        RECT 490.950 168.600 493.050 169.050 ;
        RECT 499.950 168.600 502.050 169.050 ;
        RECT 505.950 168.600 508.050 169.050 ;
        RECT 514.950 168.600 517.050 169.050 ;
        RECT 490.950 167.400 508.050 168.600 ;
        RECT 490.950 166.950 493.050 167.400 ;
        RECT 499.950 166.950 502.050 167.400 ;
        RECT 505.950 166.950 508.050 167.400 ;
        RECT 512.400 167.400 517.050 168.600 ;
        RECT 469.950 165.600 472.050 166.050 ;
        RECT 512.400 165.600 513.600 167.400 ;
        RECT 514.950 166.950 517.050 167.400 ;
        RECT 523.950 166.950 526.050 169.050 ;
        RECT 535.950 168.600 538.050 169.050 ;
        RECT 544.950 168.600 547.050 169.050 ;
        RECT 535.950 167.400 547.050 168.600 ;
        RECT 535.950 166.950 538.050 167.400 ;
        RECT 544.950 166.950 547.050 167.400 ;
        RECT 550.950 168.600 553.050 169.050 ;
        RECT 569.400 168.600 570.600 170.400 ;
        RECT 598.950 169.950 601.050 170.400 ;
        RECT 604.950 169.950 607.050 170.400 ;
        RECT 628.950 171.600 631.050 172.050 ;
        RECT 634.950 171.600 637.050 172.050 ;
        RECT 628.950 170.400 637.050 171.600 ;
        RECT 628.950 169.950 631.050 170.400 ;
        RECT 634.950 169.950 637.050 170.400 ;
        RECT 637.950 171.600 640.050 172.050 ;
        RECT 679.950 171.600 682.050 172.050 ;
        RECT 685.950 171.600 688.050 172.050 ;
        RECT 697.950 171.600 700.050 172.050 ;
        RECT 637.950 170.400 645.600 171.600 ;
        RECT 637.950 169.950 640.050 170.400 ;
        RECT 583.950 168.600 586.050 169.050 ;
        RECT 622.950 168.600 625.050 169.050 ;
        RECT 640.950 168.600 643.050 169.050 ;
        RECT 550.950 167.400 573.600 168.600 ;
        RECT 550.950 166.950 553.050 167.400 ;
        RECT 469.950 164.400 513.600 165.600 ;
        RECT 469.950 163.950 472.050 164.400 ;
        RECT 514.950 163.950 517.050 166.050 ;
        RECT 469.950 162.600 472.050 163.050 ;
        RECT 442.950 161.400 472.050 162.600 ;
        RECT 442.950 160.950 445.050 161.400 ;
        RECT 469.950 160.950 472.050 161.400 ;
        RECT 487.950 162.600 490.050 163.050 ;
        RECT 515.400 162.600 516.600 163.950 ;
        RECT 524.400 163.050 525.600 166.950 ;
        RECT 572.400 166.050 573.600 167.400 ;
        RECT 583.950 167.400 643.050 168.600 ;
        RECT 583.950 166.950 586.050 167.400 ;
        RECT 617.400 166.050 618.600 167.400 ;
        RECT 622.950 166.950 625.050 167.400 ;
        RECT 640.950 166.950 643.050 167.400 ;
        RECT 541.950 163.950 544.050 166.050 ;
        RECT 571.950 163.950 574.050 166.050 ;
        RECT 616.950 163.950 619.050 166.050 ;
        RECT 487.950 161.400 516.600 162.600 ;
        RECT 487.950 160.950 490.050 161.400 ;
        RECT 523.950 160.950 526.050 163.050 ;
        RECT 529.950 162.600 532.050 163.050 ;
        RECT 535.950 162.600 538.050 163.050 ;
        RECT 529.950 161.400 538.050 162.600 ;
        RECT 542.400 162.600 543.600 163.950 ;
        RECT 580.950 162.600 583.050 163.050 ;
        RECT 542.400 161.400 583.050 162.600 ;
        RECT 529.950 160.950 532.050 161.400 ;
        RECT 535.950 160.950 538.050 161.400 ;
        RECT 580.950 160.950 583.050 161.400 ;
        RECT 604.950 162.600 607.050 163.050 ;
        RECT 625.950 162.600 628.050 163.050 ;
        RECT 604.950 161.400 628.050 162.600 ;
        RECT 604.950 160.950 607.050 161.400 ;
        RECT 625.950 160.950 628.050 161.400 ;
        RECT 628.950 162.600 631.050 163.050 ;
        RECT 637.950 162.600 640.050 163.050 ;
        RECT 628.950 161.400 640.050 162.600 ;
        RECT 628.950 160.950 631.050 161.400 ;
        RECT 637.950 160.950 640.050 161.400 ;
        RECT 145.950 159.600 148.050 160.050 ;
        RECT 122.400 158.400 148.050 159.600 ;
        RECT 112.950 157.950 115.050 158.400 ;
        RECT 145.950 157.950 148.050 158.400 ;
        RECT 175.950 159.600 178.050 160.050 ;
        RECT 190.950 159.600 193.050 160.050 ;
        RECT 175.950 158.400 193.050 159.600 ;
        RECT 175.950 157.950 178.050 158.400 ;
        RECT 190.950 157.950 193.050 158.400 ;
        RECT 277.950 159.600 280.050 160.050 ;
        RECT 310.950 159.600 313.050 160.050 ;
        RECT 277.950 158.400 313.050 159.600 ;
        RECT 277.950 157.950 280.050 158.400 ;
        RECT 310.950 157.950 313.050 158.400 ;
        RECT 313.950 159.600 316.050 160.050 ;
        RECT 325.950 159.600 328.050 160.050 ;
        RECT 313.950 158.400 328.050 159.600 ;
        RECT 313.950 157.950 316.050 158.400 ;
        RECT 325.950 157.950 328.050 158.400 ;
        RECT 328.950 159.600 331.050 160.050 ;
        RECT 343.950 159.600 346.050 160.050 ;
        RECT 328.950 158.400 346.050 159.600 ;
        RECT 328.950 157.950 331.050 158.400 ;
        RECT 343.950 157.950 346.050 158.400 ;
        RECT 361.950 159.600 364.050 160.050 ;
        RECT 365.400 159.600 366.600 160.950 ;
        RECT 361.950 158.400 366.600 159.600 ;
        RECT 367.950 159.600 370.050 160.050 ;
        RECT 394.950 159.600 397.050 160.050 ;
        RECT 367.950 158.400 397.050 159.600 ;
        RECT 361.950 157.950 364.050 158.400 ;
        RECT 367.950 157.950 370.050 158.400 ;
        RECT 394.950 157.950 397.050 158.400 ;
        RECT 409.950 159.600 412.050 160.050 ;
        RECT 427.950 159.600 430.050 160.050 ;
        RECT 514.950 159.600 517.050 160.050 ;
        RECT 409.950 158.400 430.050 159.600 ;
        RECT 409.950 157.950 412.050 158.400 ;
        RECT 427.950 157.950 430.050 158.400 ;
        RECT 431.400 158.400 517.050 159.600 ;
        RECT 58.950 156.600 61.050 157.050 ;
        RECT 79.950 156.600 82.050 157.050 ;
        RECT 58.950 155.400 82.050 156.600 ;
        RECT 58.950 154.950 61.050 155.400 ;
        RECT 79.950 154.950 82.050 155.400 ;
        RECT 82.950 156.600 85.050 157.050 ;
        RECT 127.950 156.600 130.050 157.050 ;
        RECT 82.950 155.400 130.050 156.600 ;
        RECT 82.950 154.950 85.050 155.400 ;
        RECT 127.950 154.950 130.050 155.400 ;
        RECT 133.950 156.600 136.050 157.050 ;
        RECT 187.950 156.600 190.050 157.050 ;
        RECT 133.950 155.400 190.050 156.600 ;
        RECT 133.950 154.950 136.050 155.400 ;
        RECT 187.950 154.950 190.050 155.400 ;
        RECT 319.950 156.600 322.050 157.050 ;
        RECT 337.950 156.600 340.050 157.050 ;
        RECT 319.950 155.400 340.050 156.600 ;
        RECT 319.950 154.950 322.050 155.400 ;
        RECT 337.950 154.950 340.050 155.400 ;
        RECT 355.950 156.600 358.050 157.050 ;
        RECT 431.400 156.600 432.600 158.400 ;
        RECT 514.950 157.950 517.050 158.400 ;
        RECT 565.950 159.600 568.050 160.050 ;
        RECT 568.950 159.600 571.050 160.050 ;
        RECT 592.950 159.600 595.050 160.050 ;
        RECT 565.950 158.400 595.050 159.600 ;
        RECT 565.950 157.950 568.050 158.400 ;
        RECT 568.950 157.950 571.050 158.400 ;
        RECT 592.950 157.950 595.050 158.400 ;
        RECT 640.950 159.600 643.050 160.050 ;
        RECT 644.400 159.600 645.600 170.400 ;
        RECT 679.950 170.400 700.050 171.600 ;
        RECT 679.950 169.950 682.050 170.400 ;
        RECT 685.950 169.950 688.050 170.400 ;
        RECT 697.950 169.950 700.050 170.400 ;
        RECT 715.950 171.600 718.050 172.050 ;
        RECT 730.950 171.600 733.050 172.050 ;
        RECT 715.950 170.400 733.050 171.600 ;
        RECT 715.950 169.950 718.050 170.400 ;
        RECT 730.950 169.950 733.050 170.400 ;
        RECT 736.950 171.600 739.050 172.050 ;
        RECT 742.950 171.600 745.050 172.050 ;
        RECT 736.950 170.400 745.050 171.600 ;
        RECT 736.950 169.950 739.050 170.400 ;
        RECT 742.950 169.950 745.050 170.400 ;
        RECT 751.950 171.600 754.050 172.050 ;
        RECT 766.950 171.600 769.050 172.050 ;
        RECT 775.950 171.600 778.050 172.050 ;
        RECT 751.950 170.400 778.050 171.600 ;
        RECT 751.950 169.950 754.050 170.400 ;
        RECT 766.950 169.950 769.050 170.400 ;
        RECT 775.950 169.950 778.050 170.400 ;
        RECT 655.950 168.600 658.050 169.050 ;
        RECT 739.950 168.600 742.050 169.050 ;
        RECT 655.950 167.400 742.050 168.600 ;
        RECT 655.950 166.950 658.050 167.400 ;
        RECT 739.950 166.950 742.050 167.400 ;
        RECT 766.950 168.600 769.050 169.050 ;
        RECT 784.950 168.600 787.050 169.050 ;
        RECT 766.950 167.400 787.050 168.600 ;
        RECT 766.950 166.950 769.050 167.400 ;
        RECT 784.950 166.950 787.050 167.400 ;
        RECT 844.950 168.600 847.050 169.050 ;
        RECT 856.950 168.600 859.050 169.050 ;
        RECT 844.950 167.400 859.050 168.600 ;
        RECT 844.950 166.950 847.050 167.400 ;
        RECT 856.950 166.950 859.050 167.400 ;
        RECT 673.950 165.600 676.050 166.050 ;
        RECT 691.950 165.600 694.050 166.050 ;
        RECT 715.950 165.600 718.050 166.050 ;
        RECT 673.950 164.400 694.050 165.600 ;
        RECT 673.950 163.950 676.050 164.400 ;
        RECT 691.950 163.950 694.050 164.400 ;
        RECT 710.400 164.400 718.050 165.600 ;
        RECT 688.950 162.600 691.050 163.050 ;
        RECT 694.950 162.600 697.050 163.050 ;
        RECT 688.950 161.400 697.050 162.600 ;
        RECT 688.950 160.950 691.050 161.400 ;
        RECT 694.950 160.950 697.050 161.400 ;
        RECT 700.950 162.600 703.050 163.050 ;
        RECT 710.400 162.600 711.600 164.400 ;
        RECT 715.950 163.950 718.050 164.400 ;
        RECT 745.950 165.600 748.050 166.050 ;
        RECT 790.950 165.600 793.050 166.050 ;
        RECT 745.950 164.400 793.050 165.600 ;
        RECT 745.950 163.950 748.050 164.400 ;
        RECT 790.950 163.950 793.050 164.400 ;
        RECT 832.950 165.600 835.050 166.050 ;
        RECT 847.950 165.600 850.050 166.050 ;
        RECT 853.950 165.600 856.050 166.050 ;
        RECT 832.950 164.400 856.050 165.600 ;
        RECT 832.950 163.950 835.050 164.400 ;
        RECT 847.950 163.950 850.050 164.400 ;
        RECT 853.950 163.950 856.050 164.400 ;
        RECT 700.950 161.400 711.600 162.600 ;
        RECT 700.950 160.950 703.050 161.400 ;
        RECT 712.950 160.950 715.050 163.050 ;
        RECT 748.950 162.600 751.050 163.050 ;
        RECT 763.950 162.600 766.050 163.050 ;
        RECT 778.950 162.600 781.050 163.050 ;
        RECT 748.950 161.400 781.050 162.600 ;
        RECT 748.950 160.950 751.050 161.400 ;
        RECT 763.950 160.950 766.050 161.400 ;
        RECT 778.950 160.950 781.050 161.400 ;
        RECT 820.950 162.600 823.050 163.050 ;
        RECT 841.950 162.600 844.050 163.050 ;
        RECT 853.950 162.600 856.050 163.050 ;
        RECT 820.950 161.400 856.050 162.600 ;
        RECT 820.950 160.950 823.050 161.400 ;
        RECT 841.950 160.950 844.050 161.400 ;
        RECT 853.950 160.950 856.050 161.400 ;
        RECT 640.950 158.400 645.600 159.600 ;
        RECT 673.950 159.600 676.050 160.050 ;
        RECT 682.950 159.600 685.050 160.050 ;
        RECT 673.950 158.400 685.050 159.600 ;
        RECT 640.950 157.950 643.050 158.400 ;
        RECT 673.950 157.950 676.050 158.400 ;
        RECT 682.950 157.950 685.050 158.400 ;
        RECT 700.950 159.600 703.050 160.050 ;
        RECT 713.400 159.600 714.600 160.950 ;
        RECT 700.950 158.400 714.600 159.600 ;
        RECT 700.950 157.950 703.050 158.400 ;
        RECT 355.950 155.400 432.600 156.600 ;
        RECT 439.950 156.600 442.050 157.050 ;
        RECT 487.950 156.600 490.050 157.050 ;
        RECT 439.950 155.400 490.050 156.600 ;
        RECT 355.950 154.950 358.050 155.400 ;
        RECT 439.950 154.950 442.050 155.400 ;
        RECT 487.950 154.950 490.050 155.400 ;
        RECT 493.950 156.600 496.050 157.050 ;
        RECT 508.950 156.600 511.050 157.050 ;
        RECT 562.950 156.600 565.050 157.050 ;
        RECT 493.950 155.400 565.050 156.600 ;
        RECT 493.950 154.950 496.050 155.400 ;
        RECT 508.950 154.950 511.050 155.400 ;
        RECT 562.950 154.950 565.050 155.400 ;
        RECT 592.950 156.600 595.050 157.050 ;
        RECT 652.950 156.600 655.050 157.050 ;
        RECT 733.950 156.600 736.050 157.050 ;
        RECT 592.950 155.400 736.050 156.600 ;
        RECT 592.950 154.950 595.050 155.400 ;
        RECT 652.950 154.950 655.050 155.400 ;
        RECT 733.950 154.950 736.050 155.400 ;
        RECT 43.950 153.600 46.050 154.050 ;
        RECT 73.950 153.600 76.050 154.050 ;
        RECT 43.950 152.400 76.050 153.600 ;
        RECT 43.950 151.950 46.050 152.400 ;
        RECT 73.950 151.950 76.050 152.400 ;
        RECT 88.950 153.600 91.050 154.050 ;
        RECT 124.950 153.600 127.050 154.050 ;
        RECT 88.950 152.400 127.050 153.600 ;
        RECT 88.950 151.950 91.050 152.400 ;
        RECT 124.950 151.950 127.050 152.400 ;
        RECT 178.950 153.600 181.050 154.050 ;
        RECT 187.950 153.600 190.050 154.050 ;
        RECT 178.950 152.400 190.050 153.600 ;
        RECT 178.950 151.950 181.050 152.400 ;
        RECT 187.950 151.950 190.050 152.400 ;
        RECT 247.950 153.600 250.050 154.050 ;
        RECT 289.950 153.600 292.050 154.050 ;
        RECT 247.950 152.400 292.050 153.600 ;
        RECT 247.950 151.950 250.050 152.400 ;
        RECT 289.950 151.950 292.050 152.400 ;
        RECT 349.950 153.600 352.050 154.050 ;
        RECT 364.950 153.600 367.050 154.050 ;
        RECT 349.950 152.400 367.050 153.600 ;
        RECT 349.950 151.950 352.050 152.400 ;
        RECT 364.950 151.950 367.050 152.400 ;
        RECT 382.950 153.600 385.050 154.050 ;
        RECT 397.950 153.600 400.050 154.050 ;
        RECT 382.950 152.400 400.050 153.600 ;
        RECT 382.950 151.950 385.050 152.400 ;
        RECT 397.950 151.950 400.050 152.400 ;
        RECT 406.950 153.600 409.050 154.050 ;
        RECT 436.950 153.600 439.050 154.050 ;
        RECT 406.950 152.400 439.050 153.600 ;
        RECT 406.950 151.950 409.050 152.400 ;
        RECT 436.950 151.950 439.050 152.400 ;
        RECT 442.950 153.600 445.050 154.050 ;
        RECT 481.950 153.600 484.050 154.050 ;
        RECT 442.950 152.400 484.050 153.600 ;
        RECT 442.950 151.950 445.050 152.400 ;
        RECT 481.950 151.950 484.050 152.400 ;
        RECT 538.950 153.600 541.050 154.050 ;
        RECT 547.950 153.600 550.050 154.050 ;
        RECT 538.950 152.400 550.050 153.600 ;
        RECT 538.950 151.950 541.050 152.400 ;
        RECT 547.950 151.950 550.050 152.400 ;
        RECT 562.950 153.600 565.050 154.050 ;
        RECT 607.950 153.600 610.050 154.050 ;
        RECT 562.950 152.400 610.050 153.600 ;
        RECT 562.950 151.950 565.050 152.400 ;
        RECT 607.950 151.950 610.050 152.400 ;
        RECT 610.950 153.600 613.050 154.050 ;
        RECT 781.950 153.600 784.050 154.050 ;
        RECT 610.950 152.400 784.050 153.600 ;
        RECT 610.950 151.950 613.050 152.400 ;
        RECT 781.950 151.950 784.050 152.400 ;
        RECT 40.950 150.600 43.050 151.050 ;
        RECT 97.950 150.600 100.050 151.050 ;
        RECT 121.950 150.600 124.050 151.050 ;
        RECT 40.950 149.400 66.600 150.600 ;
        RECT 40.950 148.950 43.050 149.400 ;
        RECT 52.950 147.600 55.050 148.050 ;
        RECT 58.950 147.600 61.050 148.050 ;
        RECT 52.950 146.400 61.050 147.600 ;
        RECT 65.400 147.600 66.600 149.400 ;
        RECT 97.950 149.400 124.050 150.600 ;
        RECT 97.950 148.950 100.050 149.400 ;
        RECT 121.950 148.950 124.050 149.400 ;
        RECT 151.950 150.600 154.050 151.050 ;
        RECT 214.950 150.600 217.050 151.050 ;
        RECT 151.950 149.400 217.050 150.600 ;
        RECT 151.950 148.950 154.050 149.400 ;
        RECT 214.950 148.950 217.050 149.400 ;
        RECT 229.950 150.600 232.050 151.050 ;
        RECT 490.950 150.600 493.050 151.050 ;
        RECT 229.950 149.400 493.050 150.600 ;
        RECT 229.950 148.950 232.050 149.400 ;
        RECT 490.950 148.950 493.050 149.400 ;
        RECT 652.950 150.600 655.050 151.050 ;
        RECT 664.950 150.600 667.050 151.050 ;
        RECT 652.950 149.400 667.050 150.600 ;
        RECT 652.950 148.950 655.050 149.400 ;
        RECT 664.950 148.950 667.050 149.400 ;
        RECT 109.950 147.600 112.050 148.050 ;
        RECT 65.400 146.400 112.050 147.600 ;
        RECT 52.950 145.950 55.050 146.400 ;
        RECT 58.950 145.950 61.050 146.400 ;
        RECT 109.950 145.950 112.050 146.400 ;
        RECT 115.950 147.600 118.050 148.050 ;
        RECT 205.950 147.600 208.050 148.050 ;
        RECT 115.950 146.400 208.050 147.600 ;
        RECT 115.950 145.950 118.050 146.400 ;
        RECT 205.950 145.950 208.050 146.400 ;
        RECT 217.950 147.600 220.050 148.050 ;
        RECT 673.950 147.600 676.050 148.050 ;
        RECT 688.950 147.600 691.050 148.050 ;
        RECT 217.950 146.400 691.050 147.600 ;
        RECT 217.950 145.950 220.050 146.400 ;
        RECT 673.950 145.950 676.050 146.400 ;
        RECT 688.950 145.950 691.050 146.400 ;
        RECT 34.950 144.600 37.050 145.050 ;
        RECT 88.950 144.600 91.050 145.050 ;
        RECT 118.950 144.600 121.050 145.050 ;
        RECT 130.950 144.600 133.050 145.050 ;
        RECT 34.950 143.400 133.050 144.600 ;
        RECT 34.950 142.950 37.050 143.400 ;
        RECT 88.950 142.950 91.050 143.400 ;
        RECT 118.950 142.950 121.050 143.400 ;
        RECT 130.950 142.950 133.050 143.400 ;
        RECT 154.950 144.600 157.050 145.050 ;
        RECT 271.950 144.600 274.050 145.050 ;
        RECT 154.950 143.400 274.050 144.600 ;
        RECT 154.950 142.950 157.050 143.400 ;
        RECT 271.950 142.950 274.050 143.400 ;
        RECT 304.950 144.600 307.050 145.050 ;
        RECT 376.950 144.600 379.050 145.050 ;
        RECT 304.950 143.400 379.050 144.600 ;
        RECT 304.950 142.950 307.050 143.400 ;
        RECT 376.950 142.950 379.050 143.400 ;
        RECT 379.950 144.600 382.050 145.050 ;
        RECT 439.950 144.600 442.050 145.050 ;
        RECT 379.950 143.400 442.050 144.600 ;
        RECT 379.950 142.950 382.050 143.400 ;
        RECT 439.950 142.950 442.050 143.400 ;
        RECT 460.950 144.600 463.050 145.050 ;
        RECT 475.950 144.600 478.050 145.050 ;
        RECT 460.950 143.400 478.050 144.600 ;
        RECT 460.950 142.950 463.050 143.400 ;
        RECT 475.950 142.950 478.050 143.400 ;
        RECT 478.950 144.600 481.050 145.050 ;
        RECT 502.950 144.600 505.050 145.050 ;
        RECT 478.950 143.400 505.050 144.600 ;
        RECT 478.950 142.950 481.050 143.400 ;
        RECT 502.950 142.950 505.050 143.400 ;
        RECT 574.950 144.600 577.050 145.050 ;
        RECT 610.950 144.600 613.050 145.050 ;
        RECT 574.950 143.400 613.050 144.600 ;
        RECT 574.950 142.950 577.050 143.400 ;
        RECT 610.950 142.950 613.050 143.400 ;
        RECT 643.950 144.600 646.050 145.050 ;
        RECT 748.950 144.600 751.050 145.050 ;
        RECT 760.950 144.600 763.050 145.050 ;
        RECT 643.950 143.400 763.050 144.600 ;
        RECT 643.950 142.950 646.050 143.400 ;
        RECT 748.950 142.950 751.050 143.400 ;
        RECT 760.950 142.950 763.050 143.400 ;
        RECT 49.950 141.600 52.050 142.050 ;
        RECT 73.950 141.600 76.050 142.050 ;
        RECT 49.950 140.400 76.050 141.600 ;
        RECT 49.950 139.950 52.050 140.400 ;
        RECT 73.950 139.950 76.050 140.400 ;
        RECT 112.950 141.600 115.050 142.050 ;
        RECT 193.950 141.600 196.050 142.050 ;
        RECT 112.950 140.400 196.050 141.600 ;
        RECT 112.950 139.950 115.050 140.400 ;
        RECT 193.950 139.950 196.050 140.400 ;
        RECT 199.950 141.600 202.050 142.050 ;
        RECT 421.950 141.600 424.050 142.050 ;
        RECT 199.950 140.400 424.050 141.600 ;
        RECT 199.950 139.950 202.050 140.400 ;
        RECT 421.950 139.950 424.050 140.400 ;
        RECT 424.950 141.600 427.050 142.050 ;
        RECT 445.950 141.600 448.050 142.050 ;
        RECT 424.950 140.400 448.050 141.600 ;
        RECT 424.950 139.950 427.050 140.400 ;
        RECT 445.950 139.950 448.050 140.400 ;
        RECT 457.950 141.600 460.050 142.050 ;
        RECT 478.950 141.600 481.050 142.050 ;
        RECT 457.950 140.400 481.050 141.600 ;
        RECT 457.950 139.950 460.050 140.400 ;
        RECT 478.950 139.950 481.050 140.400 ;
        RECT 511.950 141.600 514.050 142.050 ;
        RECT 562.950 141.600 565.050 142.050 ;
        RECT 595.950 141.600 598.050 142.050 ;
        RECT 511.950 140.400 565.050 141.600 ;
        RECT 511.950 139.950 514.050 140.400 ;
        RECT 562.950 139.950 565.050 140.400 ;
        RECT 566.400 140.400 598.050 141.600 ;
        RECT 346.950 138.600 349.050 139.050 ;
        RECT 379.950 138.600 382.050 139.050 ;
        RECT 346.950 137.400 382.050 138.600 ;
        RECT 346.950 136.950 349.050 137.400 ;
        RECT 379.950 136.950 382.050 137.400 ;
        RECT 394.950 138.600 397.050 139.050 ;
        RECT 412.950 138.600 415.050 139.050 ;
        RECT 394.950 137.400 415.050 138.600 ;
        RECT 394.950 136.950 397.050 137.400 ;
        RECT 412.950 136.950 415.050 137.400 ;
        RECT 448.950 138.600 451.050 139.050 ;
        RECT 463.950 138.600 466.050 139.050 ;
        RECT 448.950 137.400 466.050 138.600 ;
        RECT 448.950 136.950 451.050 137.400 ;
        RECT 463.950 136.950 466.050 137.400 ;
        RECT 481.950 138.600 484.050 139.050 ;
        RECT 499.950 138.600 502.050 139.050 ;
        RECT 481.950 137.400 502.050 138.600 ;
        RECT 481.950 136.950 484.050 137.400 ;
        RECT 499.950 136.950 502.050 137.400 ;
        RECT 508.950 138.600 511.050 139.050 ;
        RECT 523.950 138.600 526.050 139.050 ;
        RECT 508.950 137.400 526.050 138.600 ;
        RECT 508.950 136.950 511.050 137.400 ;
        RECT 523.950 136.950 526.050 137.400 ;
        RECT 541.950 138.600 544.050 139.050 ;
        RECT 559.950 138.600 562.050 139.050 ;
        RECT 566.400 138.600 567.600 140.400 ;
        RECT 595.950 139.950 598.050 140.400 ;
        RECT 601.950 141.600 604.050 142.050 ;
        RECT 616.950 141.600 619.050 142.050 ;
        RECT 601.950 140.400 619.050 141.600 ;
        RECT 601.950 139.950 604.050 140.400 ;
        RECT 616.950 139.950 619.050 140.400 ;
        RECT 664.950 141.600 667.050 142.050 ;
        RECT 697.950 141.600 700.050 142.050 ;
        RECT 706.950 141.600 709.050 142.050 ;
        RECT 664.950 140.400 709.050 141.600 ;
        RECT 664.950 139.950 667.050 140.400 ;
        RECT 697.950 139.950 700.050 140.400 ;
        RECT 706.950 139.950 709.050 140.400 ;
        RECT 541.950 137.400 567.600 138.600 ;
        RECT 628.950 138.600 631.050 139.050 ;
        RECT 724.950 138.600 727.050 139.050 ;
        RECT 736.950 138.600 739.050 139.050 ;
        RECT 754.950 138.600 757.050 139.050 ;
        RECT 628.950 137.400 757.050 138.600 ;
        RECT 541.950 136.950 544.050 137.400 ;
        RECT 559.950 136.950 562.050 137.400 ;
        RECT 628.950 136.950 631.050 137.400 ;
        RECT 724.950 136.950 727.050 137.400 ;
        RECT 736.950 136.950 739.050 137.400 ;
        RECT 754.950 136.950 757.050 137.400 ;
        RECT 106.950 135.600 109.050 136.050 ;
        RECT 205.950 135.600 208.050 136.050 ;
        RECT 106.950 134.400 208.050 135.600 ;
        RECT 106.950 133.950 109.050 134.400 ;
        RECT 205.950 133.950 208.050 134.400 ;
        RECT 259.950 135.600 262.050 136.050 ;
        RECT 289.950 135.600 292.050 136.050 ;
        RECT 259.950 134.400 292.050 135.600 ;
        RECT 259.950 133.950 262.050 134.400 ;
        RECT 289.950 133.950 292.050 134.400 ;
        RECT 307.950 135.600 310.050 136.050 ;
        RECT 328.950 135.600 331.050 136.050 ;
        RECT 580.950 135.600 583.050 136.050 ;
        RECT 751.950 135.600 754.050 136.050 ;
        RECT 307.950 134.400 754.050 135.600 ;
        RECT 307.950 133.950 310.050 134.400 ;
        RECT 328.950 133.950 331.050 134.400 ;
        RECT 580.950 133.950 583.050 134.400 ;
        RECT 751.950 133.950 754.050 134.400 ;
        RECT 28.950 132.600 31.050 133.050 ;
        RECT 82.950 132.600 85.050 133.050 ;
        RECT 85.950 132.600 88.050 133.050 ;
        RECT 118.950 132.600 121.050 133.050 ;
        RECT 136.950 132.600 139.050 133.050 ;
        RECT 28.950 131.400 139.050 132.600 ;
        RECT 28.950 130.950 31.050 131.400 ;
        RECT 82.950 130.950 85.050 131.400 ;
        RECT 85.950 130.950 88.050 131.400 ;
        RECT 118.950 130.950 121.050 131.400 ;
        RECT 136.950 130.950 139.050 131.400 ;
        RECT 166.950 132.600 169.050 133.050 ;
        RECT 175.950 132.600 178.050 133.050 ;
        RECT 166.950 131.400 178.050 132.600 ;
        RECT 166.950 130.950 169.050 131.400 ;
        RECT 175.950 130.950 178.050 131.400 ;
        RECT 241.950 130.950 244.050 133.050 ;
        RECT 256.950 132.600 259.050 133.050 ;
        RECT 265.950 132.600 268.050 133.050 ;
        RECT 256.950 131.400 268.050 132.600 ;
        RECT 256.950 130.950 259.050 131.400 ;
        RECT 265.950 130.950 268.050 131.400 ;
        RECT 274.950 130.950 277.050 133.050 ;
        RECT 283.950 132.600 286.050 133.050 ;
        RECT 292.950 132.600 295.050 133.050 ;
        RECT 346.950 132.600 349.050 133.050 ;
        RECT 283.950 131.400 349.050 132.600 ;
        RECT 283.950 130.950 286.050 131.400 ;
        RECT 292.950 130.950 295.050 131.400 ;
        RECT 346.950 130.950 349.050 131.400 ;
        RECT 349.950 132.600 352.050 133.050 ;
        RECT 358.950 132.600 361.050 133.050 ;
        RECT 382.950 132.600 385.050 133.050 ;
        RECT 349.950 131.400 361.050 132.600 ;
        RECT 349.950 130.950 352.050 131.400 ;
        RECT 358.950 130.950 361.050 131.400 ;
        RECT 365.400 131.400 385.050 132.600 ;
        RECT 49.950 129.600 52.050 130.050 ;
        RECT 67.950 129.600 70.050 130.050 ;
        RECT 73.950 129.600 76.050 130.050 ;
        RECT 49.950 128.400 76.050 129.600 ;
        RECT 49.950 127.950 52.050 128.400 ;
        RECT 67.950 127.950 70.050 128.400 ;
        RECT 73.950 127.950 76.050 128.400 ;
        RECT 163.950 129.600 166.050 130.050 ;
        RECT 199.950 129.600 202.050 130.050 ;
        RECT 217.950 129.600 220.050 130.050 ;
        RECT 163.950 128.400 220.050 129.600 ;
        RECT 163.950 127.950 166.050 128.400 ;
        RECT 199.950 127.950 202.050 128.400 ;
        RECT 217.950 127.950 220.050 128.400 ;
        RECT 94.950 126.600 97.050 127.050 ;
        RECT 103.950 126.600 106.050 127.050 ;
        RECT 154.950 126.600 157.050 127.050 ;
        RECT 166.950 126.600 169.050 127.050 ;
        RECT 94.950 125.400 102.600 126.600 ;
        RECT 94.950 124.950 97.050 125.400 ;
        RECT 101.400 124.050 102.600 125.400 ;
        RECT 103.950 125.400 169.050 126.600 ;
        RECT 103.950 124.950 106.050 125.400 ;
        RECT 154.950 124.950 157.050 125.400 ;
        RECT 166.950 124.950 169.050 125.400 ;
        RECT 175.950 126.600 178.050 127.050 ;
        RECT 202.950 126.600 205.050 127.050 ;
        RECT 175.950 125.400 205.050 126.600 ;
        RECT 175.950 124.950 178.050 125.400 ;
        RECT 202.950 124.950 205.050 125.400 ;
        RECT 214.950 126.600 217.050 127.050 ;
        RECT 220.950 126.600 223.050 127.050 ;
        RECT 214.950 125.400 223.050 126.600 ;
        RECT 242.400 126.600 243.600 130.950 ;
        RECT 247.950 127.950 250.050 130.050 ;
        RECT 244.950 126.600 247.050 127.050 ;
        RECT 242.400 125.400 247.050 126.600 ;
        RECT 248.400 126.600 249.600 127.950 ;
        RECT 275.400 127.050 276.600 130.950 ;
        RECT 277.950 129.600 280.050 130.050 ;
        RECT 304.950 129.600 307.050 130.050 ;
        RECT 310.950 129.600 313.050 130.050 ;
        RECT 277.950 128.400 303.600 129.600 ;
        RECT 277.950 127.950 280.050 128.400 ;
        RECT 256.950 126.600 259.050 127.050 ;
        RECT 248.400 125.400 259.050 126.600 ;
        RECT 214.950 124.950 217.050 125.400 ;
        RECT 220.950 124.950 223.050 125.400 ;
        RECT 244.950 124.950 247.050 125.400 ;
        RECT 256.950 124.950 259.050 125.400 ;
        RECT 274.950 124.950 277.050 127.050 ;
        RECT 302.400 126.600 303.600 128.400 ;
        RECT 304.950 128.400 313.050 129.600 ;
        RECT 304.950 127.950 307.050 128.400 ;
        RECT 310.950 127.950 313.050 128.400 ;
        RECT 331.950 129.600 334.050 130.050 ;
        RECT 340.950 129.600 343.050 130.050 ;
        RECT 331.950 128.400 343.050 129.600 ;
        RECT 331.950 127.950 334.050 128.400 ;
        RECT 340.950 127.950 343.050 128.400 ;
        RECT 352.950 129.600 355.050 130.050 ;
        RECT 358.950 129.600 361.050 130.050 ;
        RECT 365.400 129.600 366.600 131.400 ;
        RECT 382.950 130.950 385.050 131.400 ;
        RECT 391.950 132.600 394.050 133.050 ;
        RECT 397.950 132.600 400.050 133.050 ;
        RECT 391.950 131.400 400.050 132.600 ;
        RECT 391.950 130.950 394.050 131.400 ;
        RECT 397.950 130.950 400.050 131.400 ;
        RECT 412.950 132.600 415.050 133.050 ;
        RECT 478.950 132.600 481.050 133.050 ;
        RECT 556.950 132.600 559.050 133.050 ;
        RECT 580.950 132.600 583.050 133.050 ;
        RECT 412.950 131.400 477.600 132.600 ;
        RECT 412.950 130.950 415.050 131.400 ;
        RECT 352.950 128.400 361.050 129.600 ;
        RECT 352.950 127.950 355.050 128.400 ;
        RECT 358.950 127.950 361.050 128.400 ;
        RECT 362.400 128.400 366.600 129.600 ;
        RECT 373.950 129.600 376.050 130.050 ;
        RECT 385.950 129.600 388.050 130.050 ;
        RECT 400.950 129.600 403.050 130.050 ;
        RECT 373.950 128.400 381.600 129.600 ;
        RECT 334.950 126.600 337.050 127.050 ;
        RECT 355.950 126.600 358.050 127.050 ;
        RECT 302.400 125.400 337.050 126.600 ;
        RECT 334.950 124.950 337.050 125.400 ;
        RECT 350.400 125.400 358.050 126.600 ;
        RECT 70.950 123.600 73.050 124.050 ;
        RECT 100.950 123.600 103.050 124.050 ;
        RECT 70.950 122.400 103.050 123.600 ;
        RECT 70.950 121.950 73.050 122.400 ;
        RECT 100.950 121.950 103.050 122.400 ;
        RECT 106.950 123.600 109.050 124.050 ;
        RECT 112.950 123.600 115.050 124.050 ;
        RECT 106.950 122.400 115.050 123.600 ;
        RECT 106.950 121.950 109.050 122.400 ;
        RECT 112.950 121.950 115.050 122.400 ;
        RECT 115.950 123.600 118.050 124.050 ;
        RECT 133.950 123.600 136.050 124.050 ;
        RECT 169.950 123.600 172.050 124.050 ;
        RECT 115.950 122.400 172.050 123.600 ;
        RECT 115.950 121.950 118.050 122.400 ;
        RECT 133.950 121.950 136.050 122.400 ;
        RECT 169.950 121.950 172.050 122.400 ;
        RECT 187.950 123.600 190.050 124.050 ;
        RECT 214.950 123.600 217.050 124.050 ;
        RECT 187.950 122.400 217.050 123.600 ;
        RECT 187.950 121.950 190.050 122.400 ;
        RECT 214.950 121.950 217.050 122.400 ;
        RECT 217.950 123.600 220.050 124.050 ;
        RECT 223.950 123.600 226.050 124.050 ;
        RECT 217.950 122.400 226.050 123.600 ;
        RECT 217.950 121.950 220.050 122.400 ;
        RECT 223.950 121.950 226.050 122.400 ;
        RECT 238.950 123.600 241.050 124.050 ;
        RECT 262.950 123.600 265.050 124.050 ;
        RECT 238.950 122.400 265.050 123.600 ;
        RECT 238.950 121.950 241.050 122.400 ;
        RECT 262.950 121.950 265.050 122.400 ;
        RECT 286.950 123.600 289.050 124.050 ;
        RECT 298.950 123.600 301.050 124.050 ;
        RECT 286.950 122.400 301.050 123.600 ;
        RECT 286.950 121.950 289.050 122.400 ;
        RECT 298.950 121.950 301.050 122.400 ;
        RECT 307.950 123.600 310.050 124.050 ;
        RECT 313.950 123.600 316.050 124.050 ;
        RECT 307.950 122.400 316.050 123.600 ;
        RECT 307.950 121.950 310.050 122.400 ;
        RECT 313.950 121.950 316.050 122.400 ;
        RECT 328.950 123.600 331.050 124.050 ;
        RECT 346.950 123.600 349.050 124.050 ;
        RECT 328.950 122.400 349.050 123.600 ;
        RECT 328.950 121.950 331.050 122.400 ;
        RECT 346.950 121.950 349.050 122.400 ;
        RECT 61.950 120.600 64.050 121.050 ;
        RECT 73.950 120.600 76.050 121.050 ;
        RECT 61.950 119.400 76.050 120.600 ;
        RECT 61.950 118.950 64.050 119.400 ;
        RECT 73.950 118.950 76.050 119.400 ;
        RECT 82.950 120.600 85.050 121.050 ;
        RECT 85.950 120.600 88.050 121.050 ;
        RECT 91.950 120.600 94.050 121.050 ;
        RECT 82.950 119.400 94.050 120.600 ;
        RECT 82.950 118.950 85.050 119.400 ;
        RECT 85.950 118.950 88.050 119.400 ;
        RECT 91.950 118.950 94.050 119.400 ;
        RECT 121.950 120.600 124.050 121.050 ;
        RECT 127.950 120.600 130.050 121.050 ;
        RECT 121.950 119.400 130.050 120.600 ;
        RECT 121.950 118.950 124.050 119.400 ;
        RECT 127.950 118.950 130.050 119.400 ;
        RECT 139.950 120.600 142.050 121.050 ;
        RECT 160.950 120.600 163.050 121.050 ;
        RECT 184.950 120.600 187.050 121.050 ;
        RECT 196.950 120.600 199.050 121.050 ;
        RECT 208.950 120.600 211.050 121.050 ;
        RECT 139.950 119.400 211.050 120.600 ;
        RECT 139.950 118.950 142.050 119.400 ;
        RECT 160.950 118.950 163.050 119.400 ;
        RECT 184.950 118.950 187.050 119.400 ;
        RECT 196.950 118.950 199.050 119.400 ;
        RECT 208.950 118.950 211.050 119.400 ;
        RECT 322.950 120.600 325.050 121.050 ;
        RECT 337.950 120.600 340.050 121.050 ;
        RECT 322.950 119.400 340.050 120.600 ;
        RECT 350.400 120.600 351.600 125.400 ;
        RECT 355.950 124.950 358.050 125.400 ;
        RECT 352.950 123.600 355.050 124.050 ;
        RECT 362.400 123.600 363.600 128.400 ;
        RECT 373.950 127.950 376.050 128.400 ;
        RECT 364.950 126.600 367.050 127.050 ;
        RECT 376.950 126.600 379.050 127.050 ;
        RECT 364.950 125.400 379.050 126.600 ;
        RECT 380.400 126.600 381.600 128.400 ;
        RECT 385.950 128.400 403.050 129.600 ;
        RECT 385.950 127.950 388.050 128.400 ;
        RECT 400.950 127.950 403.050 128.400 ;
        RECT 427.950 129.600 430.050 130.050 ;
        RECT 457.950 129.600 460.050 130.050 ;
        RECT 427.950 128.400 460.050 129.600 ;
        RECT 476.400 129.600 477.600 131.400 ;
        RECT 478.950 131.400 555.600 132.600 ;
        RECT 478.950 130.950 481.050 131.400 ;
        RECT 484.950 129.600 487.050 130.050 ;
        RECT 508.950 129.600 511.050 130.050 ;
        RECT 476.400 128.400 480.600 129.600 ;
        RECT 427.950 127.950 430.050 128.400 ;
        RECT 457.950 127.950 460.050 128.400 ;
        RECT 479.400 127.050 480.600 128.400 ;
        RECT 484.950 128.400 511.050 129.600 ;
        RECT 484.950 127.950 487.050 128.400 ;
        RECT 508.950 127.950 511.050 128.400 ;
        RECT 517.950 127.950 520.050 130.050 ;
        RECT 554.400 129.600 555.600 131.400 ;
        RECT 556.950 131.400 583.050 132.600 ;
        RECT 556.950 130.950 559.050 131.400 ;
        RECT 580.950 130.950 583.050 131.400 ;
        RECT 598.950 132.600 601.050 133.050 ;
        RECT 613.950 132.600 616.050 133.050 ;
        RECT 625.950 132.600 628.050 133.050 ;
        RECT 598.950 131.400 628.050 132.600 ;
        RECT 598.950 130.950 601.050 131.400 ;
        RECT 613.950 130.950 616.050 131.400 ;
        RECT 625.950 130.950 628.050 131.400 ;
        RECT 649.950 130.950 652.050 133.050 ;
        RECT 721.950 132.600 724.050 133.050 ;
        RECT 733.950 132.600 736.050 133.050 ;
        RECT 742.950 132.600 745.050 133.050 ;
        RECT 721.950 131.400 729.600 132.600 ;
        RECT 721.950 130.950 724.050 131.400 ;
        RECT 628.950 129.600 631.050 130.050 ;
        RECT 554.400 128.400 631.050 129.600 ;
        RECT 650.400 129.600 651.600 130.950 ;
        RECT 728.400 130.050 729.600 131.400 ;
        RECT 733.950 131.400 745.050 132.600 ;
        RECT 733.950 130.950 736.050 131.400 ;
        RECT 742.950 130.950 745.050 131.400 ;
        RECT 679.950 129.600 682.050 130.050 ;
        RECT 691.950 129.600 694.050 130.050 ;
        RECT 700.950 129.600 703.050 130.050 ;
        RECT 650.400 128.400 675.600 129.600 ;
        RECT 628.950 127.950 631.050 128.400 ;
        RECT 394.950 126.600 397.050 127.050 ;
        RECT 442.950 126.600 445.050 127.050 ;
        RECT 380.400 125.400 397.050 126.600 ;
        RECT 364.950 124.950 367.050 125.400 ;
        RECT 376.950 124.950 379.050 125.400 ;
        RECT 394.950 124.950 397.050 125.400 ;
        RECT 419.400 125.400 445.050 126.600 ;
        RECT 419.400 124.050 420.600 125.400 ;
        RECT 442.950 124.950 445.050 125.400 ;
        RECT 466.950 126.600 469.050 127.050 ;
        RECT 472.950 126.600 475.050 127.050 ;
        RECT 466.950 125.400 475.050 126.600 ;
        RECT 466.950 124.950 469.050 125.400 ;
        RECT 472.950 124.950 475.050 125.400 ;
        RECT 478.950 124.950 481.050 127.050 ;
        RECT 505.950 126.600 508.050 127.050 ;
        RECT 511.950 126.600 514.050 127.050 ;
        RECT 518.400 126.600 519.600 127.950 ;
        RECT 505.950 125.400 514.050 126.600 ;
        RECT 505.950 124.950 508.050 125.400 ;
        RECT 511.950 124.950 514.050 125.400 ;
        RECT 515.400 125.400 519.600 126.600 ;
        RECT 520.950 126.600 523.050 127.050 ;
        RECT 535.950 126.600 538.050 127.050 ;
        RECT 520.950 125.400 538.050 126.600 ;
        RECT 352.950 122.400 363.600 123.600 ;
        RECT 373.950 123.600 376.050 124.050 ;
        RECT 382.950 123.600 385.050 124.050 ;
        RECT 373.950 122.400 385.050 123.600 ;
        RECT 352.950 121.950 355.050 122.400 ;
        RECT 373.950 121.950 376.050 122.400 ;
        RECT 382.950 121.950 385.050 122.400 ;
        RECT 418.950 121.950 421.050 124.050 ;
        RECT 439.950 123.600 442.050 124.050 ;
        RECT 445.950 123.600 448.050 124.050 ;
        RECT 439.950 122.400 448.050 123.600 ;
        RECT 439.950 121.950 442.050 122.400 ;
        RECT 445.950 121.950 448.050 122.400 ;
        RECT 451.950 123.600 454.050 124.050 ;
        RECT 463.950 123.600 466.050 124.050 ;
        RECT 451.950 122.400 466.050 123.600 ;
        RECT 451.950 121.950 454.050 122.400 ;
        RECT 463.950 121.950 466.050 122.400 ;
        RECT 481.950 123.600 484.050 124.050 ;
        RECT 496.950 123.600 499.050 124.050 ;
        RECT 481.950 122.400 499.050 123.600 ;
        RECT 481.950 121.950 484.050 122.400 ;
        RECT 496.950 121.950 499.050 122.400 ;
        RECT 505.950 123.600 508.050 124.050 ;
        RECT 515.400 123.600 516.600 125.400 ;
        RECT 520.950 124.950 523.050 125.400 ;
        RECT 535.950 124.950 538.050 125.400 ;
        RECT 550.950 126.600 553.050 127.050 ;
        RECT 559.950 126.600 562.050 127.050 ;
        RECT 550.950 125.400 562.050 126.600 ;
        RECT 550.950 124.950 553.050 125.400 ;
        RECT 559.950 124.950 562.050 125.400 ;
        RECT 571.950 126.600 574.050 127.050 ;
        RECT 592.950 126.600 595.050 127.050 ;
        RECT 631.950 126.600 634.050 127.050 ;
        RECT 571.950 125.400 634.050 126.600 ;
        RECT 571.950 124.950 574.050 125.400 ;
        RECT 592.950 124.950 595.050 125.400 ;
        RECT 631.950 124.950 634.050 125.400 ;
        RECT 643.950 126.600 646.050 127.050 ;
        RECT 670.950 126.600 673.050 127.050 ;
        RECT 643.950 125.400 673.050 126.600 ;
        RECT 643.950 124.950 646.050 125.400 ;
        RECT 670.950 124.950 673.050 125.400 ;
        RECT 505.950 122.400 516.600 123.600 ;
        RECT 553.950 123.600 556.050 124.050 ;
        RECT 562.950 123.600 565.050 124.050 ;
        RECT 553.950 122.400 565.050 123.600 ;
        RECT 505.950 121.950 508.050 122.400 ;
        RECT 553.950 121.950 556.050 122.400 ;
        RECT 562.950 121.950 565.050 122.400 ;
        RECT 586.950 123.600 589.050 124.050 ;
        RECT 598.950 123.600 601.050 124.050 ;
        RECT 586.950 122.400 601.050 123.600 ;
        RECT 586.950 121.950 589.050 122.400 ;
        RECT 598.950 121.950 601.050 122.400 ;
        RECT 604.950 123.600 607.050 124.050 ;
        RECT 619.950 123.600 622.050 124.050 ;
        RECT 604.950 122.400 622.050 123.600 ;
        RECT 604.950 121.950 607.050 122.400 ;
        RECT 619.950 121.950 622.050 122.400 ;
        RECT 628.950 123.600 631.050 124.050 ;
        RECT 649.950 123.600 652.050 124.050 ;
        RECT 658.950 123.600 661.050 124.050 ;
        RECT 628.950 122.400 661.050 123.600 ;
        RECT 674.400 123.600 675.600 128.400 ;
        RECT 679.950 128.400 690.600 129.600 ;
        RECT 679.950 127.950 682.050 128.400 ;
        RECT 685.950 124.950 688.050 127.050 ;
        RECT 689.400 126.600 690.600 128.400 ;
        RECT 691.950 128.400 703.050 129.600 ;
        RECT 691.950 127.950 694.050 128.400 ;
        RECT 700.950 127.950 703.050 128.400 ;
        RECT 706.950 127.950 709.050 130.050 ;
        RECT 727.950 127.950 730.050 130.050 ;
        RECT 742.950 129.600 745.050 130.050 ;
        RECT 784.950 129.600 787.050 130.050 ;
        RECT 850.950 129.600 853.050 130.050 ;
        RECT 742.950 128.400 787.050 129.600 ;
        RECT 742.950 127.950 745.050 128.400 ;
        RECT 784.950 127.950 787.050 128.400 ;
        RECT 800.400 128.400 853.050 129.600 ;
        RECT 694.950 126.600 697.050 127.050 ;
        RECT 689.400 125.400 697.050 126.600 ;
        RECT 707.400 126.600 708.600 127.950 ;
        RECT 800.400 127.050 801.600 128.400 ;
        RECT 850.950 127.950 853.050 128.400 ;
        RECT 775.950 126.600 778.050 127.050 ;
        RECT 707.400 125.400 778.050 126.600 ;
        RECT 694.950 124.950 697.050 125.400 ;
        RECT 676.950 123.600 679.050 124.050 ;
        RECT 674.400 122.400 679.050 123.600 ;
        RECT 628.950 121.950 631.050 122.400 ;
        RECT 649.950 121.950 652.050 122.400 ;
        RECT 658.950 121.950 661.050 122.400 ;
        RECT 676.950 121.950 679.050 122.400 ;
        RECT 373.950 120.600 376.050 121.050 ;
        RECT 350.400 119.400 376.050 120.600 ;
        RECT 322.950 118.950 325.050 119.400 ;
        RECT 337.950 118.950 340.050 119.400 ;
        RECT 373.950 118.950 376.050 119.400 ;
        RECT 376.950 120.600 379.050 121.050 ;
        RECT 388.950 120.600 391.050 121.050 ;
        RECT 376.950 119.400 391.050 120.600 ;
        RECT 376.950 118.950 379.050 119.400 ;
        RECT 388.950 118.950 391.050 119.400 ;
        RECT 418.950 120.600 421.050 121.050 ;
        RECT 424.950 120.600 427.050 121.050 ;
        RECT 418.950 119.400 427.050 120.600 ;
        RECT 418.950 118.950 421.050 119.400 ;
        RECT 424.950 118.950 427.050 119.400 ;
        RECT 430.950 120.600 433.050 121.050 ;
        RECT 472.950 120.600 475.050 121.050 ;
        RECT 430.950 119.400 475.050 120.600 ;
        RECT 430.950 118.950 433.050 119.400 ;
        RECT 472.950 118.950 475.050 119.400 ;
        RECT 475.950 120.600 478.050 121.050 ;
        RECT 532.950 120.600 535.050 121.050 ;
        RECT 475.950 119.400 535.050 120.600 ;
        RECT 475.950 118.950 478.050 119.400 ;
        RECT 532.950 118.950 535.050 119.400 ;
        RECT 538.950 120.600 541.050 121.050 ;
        RECT 592.950 120.600 595.050 121.050 ;
        RECT 538.950 119.400 595.050 120.600 ;
        RECT 538.950 118.950 541.050 119.400 ;
        RECT 592.950 118.950 595.050 119.400 ;
        RECT 595.950 120.600 598.050 121.050 ;
        RECT 625.950 120.600 628.050 121.050 ;
        RECT 634.950 120.600 637.050 121.050 ;
        RECT 595.950 119.400 637.050 120.600 ;
        RECT 595.950 118.950 598.050 119.400 ;
        RECT 625.950 118.950 628.050 119.400 ;
        RECT 634.950 118.950 637.050 119.400 ;
        RECT 646.950 120.600 649.050 121.050 ;
        RECT 658.950 120.600 661.050 121.050 ;
        RECT 646.950 119.400 661.050 120.600 ;
        RECT 646.950 118.950 649.050 119.400 ;
        RECT 658.950 118.950 661.050 119.400 ;
        RECT 673.950 120.600 676.050 121.050 ;
        RECT 682.950 120.600 685.050 121.050 ;
        RECT 673.950 119.400 685.050 120.600 ;
        RECT 686.400 120.600 687.600 124.950 ;
        RECT 758.400 124.050 759.600 125.400 ;
        RECT 775.950 124.950 778.050 125.400 ;
        RECT 781.950 126.600 784.050 127.050 ;
        RECT 787.950 126.600 790.050 127.050 ;
        RECT 781.950 125.400 790.050 126.600 ;
        RECT 781.950 124.950 784.050 125.400 ;
        RECT 787.950 124.950 790.050 125.400 ;
        RECT 799.950 124.950 802.050 127.050 ;
        RECT 829.950 126.600 832.050 127.050 ;
        RECT 838.950 126.600 841.050 127.050 ;
        RECT 850.950 126.600 853.050 127.050 ;
        RECT 829.950 125.400 853.050 126.600 ;
        RECT 829.950 124.950 832.050 125.400 ;
        RECT 838.950 124.950 841.050 125.400 ;
        RECT 850.950 124.950 853.050 125.400 ;
        RECT 688.950 123.600 691.050 124.050 ;
        RECT 694.950 123.600 697.050 124.050 ;
        RECT 688.950 122.400 697.050 123.600 ;
        RECT 688.950 121.950 691.050 122.400 ;
        RECT 694.950 121.950 697.050 122.400 ;
        RECT 709.950 123.600 712.050 124.050 ;
        RECT 718.950 123.600 721.050 124.050 ;
        RECT 709.950 122.400 721.050 123.600 ;
        RECT 709.950 121.950 712.050 122.400 ;
        RECT 718.950 121.950 721.050 122.400 ;
        RECT 757.950 121.950 760.050 124.050 ;
        RECT 796.950 123.600 799.050 124.050 ;
        RECT 805.950 123.600 808.050 124.050 ;
        RECT 796.950 122.400 808.050 123.600 ;
        RECT 796.950 121.950 799.050 122.400 ;
        RECT 805.950 121.950 808.050 122.400 ;
        RECT 817.950 123.600 820.050 124.050 ;
        RECT 823.950 123.600 826.050 124.050 ;
        RECT 817.950 122.400 826.050 123.600 ;
        RECT 817.950 121.950 820.050 122.400 ;
        RECT 823.950 121.950 826.050 122.400 ;
        RECT 706.950 120.600 709.050 121.050 ;
        RECT 686.400 119.400 709.050 120.600 ;
        RECT 673.950 118.950 676.050 119.400 ;
        RECT 682.950 118.950 685.050 119.400 ;
        RECT 706.950 118.950 709.050 119.400 ;
        RECT 715.950 120.600 718.050 121.050 ;
        RECT 757.950 120.600 760.050 121.050 ;
        RECT 715.950 119.400 760.050 120.600 ;
        RECT 715.950 118.950 718.050 119.400 ;
        RECT 757.950 118.950 760.050 119.400 ;
        RECT 784.950 120.600 787.050 121.050 ;
        RECT 814.950 120.600 817.050 121.050 ;
        RECT 784.950 119.400 817.050 120.600 ;
        RECT 784.950 118.950 787.050 119.400 ;
        RECT 814.950 118.950 817.050 119.400 ;
        RECT 52.950 117.600 55.050 118.050 ;
        RECT 58.950 117.600 61.050 118.050 ;
        RECT 52.950 116.400 61.050 117.600 ;
        RECT 52.950 115.950 55.050 116.400 ;
        RECT 58.950 115.950 61.050 116.400 ;
        RECT 109.950 117.600 112.050 118.050 ;
        RECT 142.950 117.600 145.050 118.050 ;
        RECT 148.950 117.600 151.050 118.050 ;
        RECT 166.950 117.600 169.050 118.050 ;
        RECT 109.950 116.400 169.050 117.600 ;
        RECT 109.950 115.950 112.050 116.400 ;
        RECT 142.950 115.950 145.050 116.400 ;
        RECT 148.950 115.950 151.050 116.400 ;
        RECT 166.950 115.950 169.050 116.400 ;
        RECT 172.950 117.600 175.050 118.050 ;
        RECT 190.950 117.600 193.050 118.050 ;
        RECT 172.950 116.400 193.050 117.600 ;
        RECT 172.950 115.950 175.050 116.400 ;
        RECT 190.950 115.950 193.050 116.400 ;
        RECT 265.950 117.600 268.050 118.050 ;
        RECT 286.950 117.600 289.050 118.050 ;
        RECT 265.950 116.400 289.050 117.600 ;
        RECT 265.950 115.950 268.050 116.400 ;
        RECT 286.950 115.950 289.050 116.400 ;
        RECT 331.950 117.600 334.050 118.050 ;
        RECT 364.950 117.600 367.050 118.050 ;
        RECT 403.950 117.600 406.050 118.050 ;
        RECT 331.950 116.400 406.050 117.600 ;
        RECT 331.950 115.950 334.050 116.400 ;
        RECT 364.950 115.950 367.050 116.400 ;
        RECT 403.950 115.950 406.050 116.400 ;
        RECT 409.950 117.600 412.050 118.050 ;
        RECT 415.950 117.600 418.050 118.050 ;
        RECT 499.950 117.600 502.050 118.050 ;
        RECT 715.950 117.600 718.050 118.050 ;
        RECT 409.950 116.400 718.050 117.600 ;
        RECT 409.950 115.950 412.050 116.400 ;
        RECT 415.950 115.950 418.050 116.400 ;
        RECT 499.950 115.950 502.050 116.400 ;
        RECT 715.950 115.950 718.050 116.400 ;
        RECT 718.950 117.600 721.050 118.050 ;
        RECT 739.950 117.600 742.050 118.050 ;
        RECT 718.950 116.400 742.050 117.600 ;
        RECT 718.950 115.950 721.050 116.400 ;
        RECT 739.950 115.950 742.050 116.400 ;
        RECT 760.950 117.600 763.050 118.050 ;
        RECT 820.950 117.600 823.050 118.050 ;
        RECT 760.950 116.400 823.050 117.600 ;
        RECT 760.950 115.950 763.050 116.400 ;
        RECT 820.950 115.950 823.050 116.400 ;
        RECT 163.950 114.600 166.050 115.050 ;
        RECT 178.950 114.600 181.050 115.050 ;
        RECT 163.950 113.400 181.050 114.600 ;
        RECT 163.950 112.950 166.050 113.400 ;
        RECT 178.950 112.950 181.050 113.400 ;
        RECT 199.950 114.600 202.050 115.050 ;
        RECT 289.950 114.600 292.050 115.050 ;
        RECT 199.950 113.400 292.050 114.600 ;
        RECT 199.950 112.950 202.050 113.400 ;
        RECT 289.950 112.950 292.050 113.400 ;
        RECT 295.950 114.600 298.050 115.050 ;
        RECT 361.950 114.600 364.050 115.050 ;
        RECT 406.950 114.600 409.050 115.050 ;
        RECT 430.950 114.600 433.050 115.050 ;
        RECT 433.950 114.600 436.050 115.050 ;
        RECT 466.950 114.600 469.050 115.050 ;
        RECT 481.950 114.600 484.050 115.050 ;
        RECT 295.950 113.400 484.050 114.600 ;
        RECT 295.950 112.950 298.050 113.400 ;
        RECT 361.950 112.950 364.050 113.400 ;
        RECT 406.950 112.950 409.050 113.400 ;
        RECT 430.950 112.950 433.050 113.400 ;
        RECT 433.950 112.950 436.050 113.400 ;
        RECT 466.950 112.950 469.050 113.400 ;
        RECT 481.950 112.950 484.050 113.400 ;
        RECT 487.950 114.600 490.050 115.050 ;
        RECT 496.950 114.600 499.050 115.050 ;
        RECT 487.950 113.400 499.050 114.600 ;
        RECT 487.950 112.950 490.050 113.400 ;
        RECT 496.950 112.950 499.050 113.400 ;
        RECT 508.950 114.600 511.050 115.050 ;
        RECT 586.950 114.600 589.050 115.050 ;
        RECT 589.950 114.600 592.050 115.050 ;
        RECT 508.950 113.400 592.050 114.600 ;
        RECT 508.950 112.950 511.050 113.400 ;
        RECT 586.950 112.950 589.050 113.400 ;
        RECT 589.950 112.950 592.050 113.400 ;
        RECT 592.950 114.600 595.050 115.050 ;
        RECT 655.950 114.600 658.050 115.050 ;
        RECT 592.950 113.400 658.050 114.600 ;
        RECT 592.950 112.950 595.050 113.400 ;
        RECT 655.950 112.950 658.050 113.400 ;
        RECT 685.950 114.600 688.050 115.050 ;
        RECT 700.950 114.600 703.050 115.050 ;
        RECT 685.950 113.400 703.050 114.600 ;
        RECT 685.950 112.950 688.050 113.400 ;
        RECT 700.950 112.950 703.050 113.400 ;
        RECT 727.950 114.600 730.050 115.050 ;
        RECT 751.950 114.600 754.050 115.050 ;
        RECT 763.950 114.600 766.050 115.050 ;
        RECT 772.950 114.600 775.050 115.050 ;
        RECT 775.950 114.600 778.050 115.050 ;
        RECT 727.950 113.400 778.050 114.600 ;
        RECT 727.950 112.950 730.050 113.400 ;
        RECT 751.950 112.950 754.050 113.400 ;
        RECT 763.950 112.950 766.050 113.400 ;
        RECT 772.950 112.950 775.050 113.400 ;
        RECT 775.950 112.950 778.050 113.400 ;
        RECT 787.950 114.600 790.050 115.050 ;
        RECT 802.950 114.600 805.050 115.050 ;
        RECT 787.950 113.400 805.050 114.600 ;
        RECT 787.950 112.950 790.050 113.400 ;
        RECT 802.950 112.950 805.050 113.400 ;
        RECT 46.950 111.600 49.050 112.050 ;
        RECT 55.950 111.600 58.050 112.050 ;
        RECT 46.950 110.400 58.050 111.600 ;
        RECT 46.950 109.950 49.050 110.400 ;
        RECT 55.950 109.950 58.050 110.400 ;
        RECT 67.950 111.600 70.050 112.050 ;
        RECT 235.950 111.600 238.050 112.050 ;
        RECT 271.950 111.600 274.050 112.050 ;
        RECT 67.950 110.400 274.050 111.600 ;
        RECT 67.950 109.950 70.050 110.400 ;
        RECT 235.950 109.950 238.050 110.400 ;
        RECT 271.950 109.950 274.050 110.400 ;
        RECT 343.950 111.600 346.050 112.050 ;
        RECT 379.950 111.600 382.050 112.050 ;
        RECT 406.950 111.600 409.050 112.050 ;
        RECT 418.950 111.600 421.050 112.050 ;
        RECT 343.950 110.400 421.050 111.600 ;
        RECT 343.950 109.950 346.050 110.400 ;
        RECT 379.950 109.950 382.050 110.400 ;
        RECT 406.950 109.950 409.050 110.400 ;
        RECT 418.950 109.950 421.050 110.400 ;
        RECT 421.950 111.600 424.050 112.050 ;
        RECT 436.950 111.600 439.050 112.050 ;
        RECT 421.950 110.400 439.050 111.600 ;
        RECT 421.950 109.950 424.050 110.400 ;
        RECT 436.950 109.950 439.050 110.400 ;
        RECT 484.950 111.600 487.050 112.050 ;
        RECT 502.950 111.600 505.050 112.050 ;
        RECT 511.950 111.600 514.050 112.050 ;
        RECT 484.950 110.400 514.050 111.600 ;
        RECT 484.950 109.950 487.050 110.400 ;
        RECT 502.950 109.950 505.050 110.400 ;
        RECT 511.950 109.950 514.050 110.400 ;
        RECT 526.950 111.600 529.050 112.050 ;
        RECT 580.950 111.600 583.050 112.050 ;
        RECT 526.950 110.400 583.050 111.600 ;
        RECT 526.950 109.950 529.050 110.400 ;
        RECT 580.950 109.950 583.050 110.400 ;
        RECT 604.950 111.600 607.050 112.050 ;
        RECT 616.950 111.600 619.050 112.050 ;
        RECT 604.950 110.400 619.050 111.600 ;
        RECT 604.950 109.950 607.050 110.400 ;
        RECT 616.950 109.950 619.050 110.400 ;
        RECT 52.950 108.600 55.050 109.050 ;
        RECT 184.950 108.600 187.050 109.050 ;
        RECT 52.950 107.400 187.050 108.600 ;
        RECT 52.950 106.950 55.050 107.400 ;
        RECT 184.950 106.950 187.050 107.400 ;
        RECT 202.950 108.600 205.050 109.050 ;
        RECT 319.950 108.600 322.050 109.050 ;
        RECT 334.950 108.600 337.050 109.050 ;
        RECT 202.950 107.400 337.050 108.600 ;
        RECT 202.950 106.950 205.050 107.400 ;
        RECT 319.950 106.950 322.050 107.400 ;
        RECT 334.950 106.950 337.050 107.400 ;
        RECT 400.950 108.600 403.050 109.050 ;
        RECT 433.950 108.600 436.050 109.050 ;
        RECT 400.950 107.400 436.050 108.600 ;
        RECT 400.950 106.950 403.050 107.400 ;
        RECT 433.950 106.950 436.050 107.400 ;
        RECT 439.950 108.600 442.050 109.050 ;
        RECT 484.950 108.600 487.050 109.050 ;
        RECT 439.950 107.400 487.050 108.600 ;
        RECT 439.950 106.950 442.050 107.400 ;
        RECT 484.950 106.950 487.050 107.400 ;
        RECT 79.950 105.600 82.050 106.050 ;
        RECT 94.950 105.600 97.050 106.050 ;
        RECT 79.950 104.400 97.050 105.600 ;
        RECT 79.950 103.950 82.050 104.400 ;
        RECT 94.950 103.950 97.050 104.400 ;
        RECT 133.950 105.600 136.050 106.050 ;
        RECT 145.950 105.600 148.050 106.050 ;
        RECT 133.950 104.400 148.050 105.600 ;
        RECT 133.950 103.950 136.050 104.400 ;
        RECT 145.950 103.950 148.050 104.400 ;
        RECT 148.950 105.600 151.050 106.050 ;
        RECT 160.950 105.600 163.050 106.050 ;
        RECT 148.950 104.400 163.050 105.600 ;
        RECT 148.950 103.950 151.050 104.400 ;
        RECT 160.950 103.950 163.050 104.400 ;
        RECT 226.950 105.600 229.050 106.050 ;
        RECT 235.950 105.600 238.050 106.050 ;
        RECT 280.950 105.600 283.050 106.050 ;
        RECT 301.950 105.600 304.050 106.050 ;
        RECT 355.950 105.600 358.050 106.050 ;
        RECT 226.950 104.400 358.050 105.600 ;
        RECT 226.950 103.950 229.050 104.400 ;
        RECT 235.950 103.950 238.050 104.400 ;
        RECT 280.950 103.950 283.050 104.400 ;
        RECT 301.950 103.950 304.050 104.400 ;
        RECT 355.950 103.950 358.050 104.400 ;
        RECT 358.950 105.600 361.050 106.050 ;
        RECT 364.950 105.600 367.050 106.050 ;
        RECT 358.950 104.400 367.050 105.600 ;
        RECT 358.950 103.950 361.050 104.400 ;
        RECT 364.950 103.950 367.050 104.400 ;
        RECT 400.950 105.600 403.050 106.050 ;
        RECT 442.950 105.600 445.050 106.050 ;
        RECT 400.950 104.400 445.050 105.600 ;
        RECT 400.950 103.950 403.050 104.400 ;
        RECT 442.950 103.950 445.050 104.400 ;
        RECT 457.950 105.600 460.050 106.050 ;
        RECT 547.950 105.600 550.050 106.050 ;
        RECT 568.950 105.600 571.050 106.050 ;
        RECT 457.950 104.400 571.050 105.600 ;
        RECT 457.950 103.950 460.050 104.400 ;
        RECT 547.950 103.950 550.050 104.400 ;
        RECT 568.950 103.950 571.050 104.400 ;
        RECT 610.950 105.600 613.050 106.050 ;
        RECT 691.950 105.600 694.050 106.050 ;
        RECT 709.950 105.600 712.050 106.050 ;
        RECT 610.950 104.400 712.050 105.600 ;
        RECT 610.950 103.950 613.050 104.400 ;
        RECT 691.950 103.950 694.050 104.400 ;
        RECT 709.950 103.950 712.050 104.400 ;
        RECT 724.950 105.600 727.050 106.050 ;
        RECT 811.950 105.600 814.050 106.050 ;
        RECT 829.950 105.600 832.050 106.050 ;
        RECT 844.950 105.600 847.050 106.050 ;
        RECT 724.950 104.400 847.050 105.600 ;
        RECT 724.950 103.950 727.050 104.400 ;
        RECT 811.950 103.950 814.050 104.400 ;
        RECT 829.950 103.950 832.050 104.400 ;
        RECT 844.950 103.950 847.050 104.400 ;
        RECT 79.950 102.600 82.050 103.050 ;
        RECT 85.950 102.600 88.050 103.050 ;
        RECT 79.950 101.400 88.050 102.600 ;
        RECT 79.950 100.950 82.050 101.400 ;
        RECT 85.950 100.950 88.050 101.400 ;
        RECT 124.950 102.600 127.050 103.050 ;
        RECT 151.950 102.600 154.050 103.050 ;
        RECT 163.950 102.600 166.050 103.050 ;
        RECT 124.950 101.400 166.050 102.600 ;
        RECT 124.950 100.950 127.050 101.400 ;
        RECT 151.950 100.950 154.050 101.400 ;
        RECT 163.950 100.950 166.050 101.400 ;
        RECT 232.950 102.600 235.050 103.050 ;
        RECT 274.950 102.600 277.050 103.050 ;
        RECT 304.950 102.600 307.050 103.050 ;
        RECT 232.950 101.400 307.050 102.600 ;
        RECT 232.950 100.950 235.050 101.400 ;
        RECT 274.950 100.950 277.050 101.400 ;
        RECT 304.950 100.950 307.050 101.400 ;
        RECT 325.950 102.600 328.050 103.050 ;
        RECT 331.950 102.600 334.050 103.050 ;
        RECT 418.950 102.600 421.050 103.050 ;
        RECT 325.950 101.400 421.050 102.600 ;
        RECT 325.950 100.950 328.050 101.400 ;
        RECT 331.950 100.950 334.050 101.400 ;
        RECT 418.950 100.950 421.050 101.400 ;
        RECT 490.950 102.600 493.050 103.050 ;
        RECT 553.950 102.600 556.050 103.050 ;
        RECT 490.950 101.400 556.050 102.600 ;
        RECT 490.950 100.950 493.050 101.400 ;
        RECT 553.950 100.950 556.050 101.400 ;
        RECT 592.950 102.600 595.050 103.050 ;
        RECT 643.950 102.600 646.050 103.050 ;
        RECT 592.950 101.400 646.050 102.600 ;
        RECT 592.950 100.950 595.050 101.400 ;
        RECT 643.950 100.950 646.050 101.400 ;
        RECT 673.950 102.600 676.050 103.050 ;
        RECT 718.950 102.600 721.050 103.050 ;
        RECT 673.950 101.400 721.050 102.600 ;
        RECT 673.950 100.950 676.050 101.400 ;
        RECT 718.950 100.950 721.050 101.400 ;
        RECT 760.950 102.600 763.050 103.050 ;
        RECT 766.950 102.600 769.050 103.050 ;
        RECT 760.950 101.400 769.050 102.600 ;
        RECT 760.950 100.950 763.050 101.400 ;
        RECT 766.950 100.950 769.050 101.400 ;
        RECT 769.950 102.600 772.050 103.050 ;
        RECT 799.950 102.600 802.050 103.050 ;
        RECT 769.950 101.400 802.050 102.600 ;
        RECT 769.950 100.950 772.050 101.400 ;
        RECT 799.950 100.950 802.050 101.400 ;
        RECT 805.950 102.600 808.050 103.050 ;
        RECT 814.950 102.600 817.050 103.050 ;
        RECT 805.950 101.400 817.050 102.600 ;
        RECT 805.950 100.950 808.050 101.400 ;
        RECT 814.950 100.950 817.050 101.400 ;
        RECT 7.950 99.600 10.050 100.050 ;
        RECT 58.950 99.600 61.050 100.050 ;
        RECT 7.950 98.400 61.050 99.600 ;
        RECT 7.950 97.950 10.050 98.400 ;
        RECT 58.950 97.950 61.050 98.400 ;
        RECT 64.950 99.600 67.050 100.050 ;
        RECT 154.950 99.600 157.050 100.050 ;
        RECT 64.950 98.400 157.050 99.600 ;
        RECT 64.950 97.950 67.050 98.400 ;
        RECT 154.950 97.950 157.050 98.400 ;
        RECT 184.950 99.600 187.050 100.050 ;
        RECT 211.950 99.600 214.050 100.050 ;
        RECT 283.950 99.600 286.050 100.050 ;
        RECT 292.950 99.600 295.050 100.050 ;
        RECT 316.950 99.600 319.050 100.050 ;
        RECT 184.950 98.400 273.600 99.600 ;
        RECT 184.950 97.950 187.050 98.400 ;
        RECT 211.950 97.950 214.050 98.400 ;
        RECT 13.950 96.600 16.050 97.050 ;
        RECT 19.950 96.600 22.050 97.050 ;
        RECT 13.950 95.400 22.050 96.600 ;
        RECT 13.950 94.950 16.050 95.400 ;
        RECT 19.950 94.950 22.050 95.400 ;
        RECT 31.950 96.600 34.050 97.050 ;
        RECT 40.950 96.600 43.050 97.050 ;
        RECT 31.950 95.400 43.050 96.600 ;
        RECT 31.950 94.950 34.050 95.400 ;
        RECT 40.950 94.950 43.050 95.400 ;
        RECT 58.950 96.600 61.050 97.050 ;
        RECT 67.950 96.600 70.050 97.050 ;
        RECT 58.950 95.400 70.050 96.600 ;
        RECT 58.950 94.950 61.050 95.400 ;
        RECT 67.950 94.950 70.050 95.400 ;
        RECT 76.950 96.600 79.050 97.050 ;
        RECT 106.950 96.600 109.050 97.050 ;
        RECT 76.950 95.400 109.050 96.600 ;
        RECT 76.950 94.950 79.050 95.400 ;
        RECT 106.950 94.950 109.050 95.400 ;
        RECT 130.950 96.600 133.050 97.050 ;
        RECT 163.950 96.600 166.050 97.050 ;
        RECT 175.950 96.600 178.050 97.050 ;
        RECT 199.950 96.600 202.050 97.050 ;
        RECT 130.950 95.400 159.600 96.600 ;
        RECT 130.950 94.950 133.050 95.400 ;
        RECT 158.400 94.050 159.600 95.400 ;
        RECT 163.950 95.400 178.050 96.600 ;
        RECT 163.950 94.950 166.050 95.400 ;
        RECT 175.950 94.950 178.050 95.400 ;
        RECT 179.400 95.400 202.050 96.600 ;
        RECT 272.400 96.600 273.600 98.400 ;
        RECT 283.950 98.400 319.050 99.600 ;
        RECT 283.950 97.950 286.050 98.400 ;
        RECT 292.950 97.950 295.050 98.400 ;
        RECT 316.950 97.950 319.050 98.400 ;
        RECT 352.950 99.600 355.050 100.050 ;
        RECT 361.950 99.600 364.050 100.050 ;
        RECT 352.950 98.400 364.050 99.600 ;
        RECT 352.950 97.950 355.050 98.400 ;
        RECT 361.950 97.950 364.050 98.400 ;
        RECT 382.950 99.600 385.050 100.050 ;
        RECT 412.950 99.600 415.050 100.050 ;
        RECT 382.950 98.400 415.050 99.600 ;
        RECT 382.950 97.950 385.050 98.400 ;
        RECT 412.950 97.950 415.050 98.400 ;
        RECT 421.950 99.600 424.050 100.050 ;
        RECT 454.950 99.600 457.050 100.050 ;
        RECT 421.950 98.400 457.050 99.600 ;
        RECT 421.950 97.950 424.050 98.400 ;
        RECT 454.950 97.950 457.050 98.400 ;
        RECT 484.950 99.600 487.050 100.050 ;
        RECT 508.950 99.600 511.050 100.050 ;
        RECT 484.950 98.400 511.050 99.600 ;
        RECT 484.950 97.950 487.050 98.400 ;
        RECT 508.950 97.950 511.050 98.400 ;
        RECT 535.950 99.600 538.050 100.050 ;
        RECT 577.950 99.600 580.050 100.050 ;
        RECT 535.950 98.400 580.050 99.600 ;
        RECT 535.950 97.950 538.050 98.400 ;
        RECT 577.950 97.950 580.050 98.400 ;
        RECT 589.950 99.600 592.050 100.050 ;
        RECT 598.950 99.600 601.050 100.050 ;
        RECT 589.950 98.400 601.050 99.600 ;
        RECT 589.950 97.950 592.050 98.400 ;
        RECT 598.950 97.950 601.050 98.400 ;
        RECT 631.950 99.600 634.050 100.050 ;
        RECT 643.950 99.600 646.050 100.050 ;
        RECT 631.950 98.400 646.050 99.600 ;
        RECT 631.950 97.950 634.050 98.400 ;
        RECT 643.950 97.950 646.050 98.400 ;
        RECT 670.950 99.600 673.050 100.050 ;
        RECT 679.950 99.600 682.050 100.050 ;
        RECT 670.950 98.400 682.050 99.600 ;
        RECT 670.950 97.950 673.050 98.400 ;
        RECT 679.950 97.950 682.050 98.400 ;
        RECT 754.950 99.600 757.050 100.050 ;
        RECT 772.950 99.600 775.050 100.050 ;
        RECT 754.950 98.400 775.050 99.600 ;
        RECT 754.950 97.950 757.050 98.400 ;
        RECT 772.950 97.950 775.050 98.400 ;
        RECT 778.950 99.600 781.050 100.050 ;
        RECT 817.950 99.600 820.050 100.050 ;
        RECT 826.950 99.600 829.050 100.050 ;
        RECT 778.950 98.400 829.050 99.600 ;
        RECT 778.950 97.950 781.050 98.400 ;
        RECT 817.950 97.950 820.050 98.400 ;
        RECT 826.950 97.950 829.050 98.400 ;
        RECT 307.950 96.600 310.050 97.050 ;
        RECT 322.950 96.600 325.050 97.050 ;
        RECT 272.400 95.400 294.600 96.600 ;
        RECT 179.400 94.050 180.600 95.400 ;
        RECT 199.950 94.950 202.050 95.400 ;
        RECT 293.400 94.050 294.600 95.400 ;
        RECT 307.950 95.400 325.050 96.600 ;
        RECT 307.950 94.950 310.050 95.400 ;
        RECT 322.950 94.950 325.050 95.400 ;
        RECT 337.950 96.600 340.050 97.050 ;
        RECT 358.950 96.600 361.050 97.050 ;
        RECT 412.950 96.600 415.050 97.050 ;
        RECT 337.950 95.400 361.050 96.600 ;
        RECT 337.950 94.950 340.050 95.400 ;
        RECT 358.950 94.950 361.050 95.400 ;
        RECT 398.400 95.400 415.050 96.600 ;
        RECT 398.400 94.050 399.600 95.400 ;
        RECT 412.950 94.950 415.050 95.400 ;
        RECT 424.950 96.600 427.050 97.050 ;
        RECT 439.950 96.600 442.050 97.050 ;
        RECT 424.950 95.400 442.050 96.600 ;
        RECT 424.950 94.950 427.050 95.400 ;
        RECT 439.950 94.950 442.050 95.400 ;
        RECT 448.950 94.950 451.050 97.050 ;
        RECT 475.950 96.600 478.050 97.050 ;
        RECT 490.950 96.600 493.050 97.050 ;
        RECT 475.950 95.400 493.050 96.600 ;
        RECT 475.950 94.950 478.050 95.400 ;
        RECT 490.950 94.950 493.050 95.400 ;
        RECT 547.950 94.950 550.050 97.050 ;
        RECT 553.950 96.600 556.050 97.050 ;
        RECT 577.950 96.600 580.050 97.050 ;
        RECT 553.950 95.400 580.050 96.600 ;
        RECT 553.950 94.950 556.050 95.400 ;
        RECT 577.950 94.950 580.050 95.400 ;
        RECT 580.950 96.600 583.050 97.050 ;
        RECT 628.950 96.600 631.050 97.050 ;
        RECT 634.950 96.600 637.050 97.050 ;
        RECT 580.950 95.400 624.600 96.600 ;
        RECT 580.950 94.950 583.050 95.400 ;
        RECT 13.950 93.600 16.050 94.050 ;
        RECT 19.950 93.600 22.050 94.050 ;
        RECT 61.950 93.600 64.050 94.050 ;
        RECT 13.950 92.400 18.600 93.600 ;
        RECT 13.950 91.950 16.050 92.400 ;
        RECT 17.400 90.600 18.600 92.400 ;
        RECT 19.950 92.400 64.050 93.600 ;
        RECT 19.950 91.950 22.050 92.400 ;
        RECT 61.950 91.950 64.050 92.400 ;
        RECT 79.950 93.600 82.050 94.050 ;
        RECT 103.950 93.600 106.050 94.050 ;
        RECT 79.950 92.400 106.050 93.600 ;
        RECT 79.950 91.950 82.050 92.400 ;
        RECT 103.950 91.950 106.050 92.400 ;
        RECT 109.950 91.950 112.050 94.050 ;
        RECT 112.950 93.600 115.050 94.050 ;
        RECT 136.950 93.600 139.050 94.050 ;
        RECT 112.950 92.400 139.050 93.600 ;
        RECT 112.950 91.950 115.050 92.400 ;
        RECT 136.950 91.950 139.050 92.400 ;
        RECT 142.950 91.950 145.050 94.050 ;
        RECT 157.950 91.950 160.050 94.050 ;
        RECT 166.950 93.600 169.050 94.050 ;
        RECT 178.950 93.600 181.050 94.050 ;
        RECT 166.950 92.400 181.050 93.600 ;
        RECT 166.950 91.950 169.050 92.400 ;
        RECT 178.950 91.950 181.050 92.400 ;
        RECT 184.950 93.600 187.050 94.050 ;
        RECT 196.950 93.600 199.050 94.050 ;
        RECT 184.950 92.400 199.050 93.600 ;
        RECT 184.950 91.950 187.050 92.400 ;
        RECT 196.950 91.950 199.050 92.400 ;
        RECT 205.950 93.600 208.050 94.050 ;
        RECT 247.950 93.600 250.050 94.050 ;
        RECT 205.950 92.400 250.050 93.600 ;
        RECT 205.950 91.950 208.050 92.400 ;
        RECT 247.950 91.950 250.050 92.400 ;
        RECT 250.950 93.600 253.050 94.050 ;
        RECT 277.950 93.600 280.050 94.050 ;
        RECT 250.950 92.400 280.050 93.600 ;
        RECT 250.950 91.950 253.050 92.400 ;
        RECT 277.950 91.950 280.050 92.400 ;
        RECT 292.950 91.950 295.050 94.050 ;
        RECT 298.950 91.950 301.050 94.050 ;
        RECT 355.950 93.600 358.050 94.050 ;
        RECT 382.950 93.600 385.050 94.050 ;
        RECT 355.950 92.400 385.050 93.600 ;
        RECT 355.950 91.950 358.050 92.400 ;
        RECT 382.950 91.950 385.050 92.400 ;
        RECT 397.950 91.950 400.050 94.050 ;
        RECT 403.950 93.600 406.050 94.050 ;
        RECT 409.950 93.600 412.050 94.050 ;
        RECT 403.950 92.400 412.050 93.600 ;
        RECT 403.950 91.950 406.050 92.400 ;
        RECT 409.950 91.950 412.050 92.400 ;
        RECT 427.950 91.950 430.050 94.050 ;
        RECT 433.950 93.600 436.050 94.050 ;
        RECT 439.950 93.600 442.050 94.050 ;
        RECT 433.950 92.400 442.050 93.600 ;
        RECT 433.950 91.950 436.050 92.400 ;
        RECT 439.950 91.950 442.050 92.400 ;
        RECT 22.950 90.600 25.050 91.050 ;
        RECT 17.400 89.400 25.050 90.600 ;
        RECT 22.950 88.950 25.050 89.400 ;
        RECT 37.950 90.600 40.050 91.050 ;
        RECT 49.950 90.600 52.050 91.050 ;
        RECT 37.950 89.400 52.050 90.600 ;
        RECT 37.950 88.950 40.050 89.400 ;
        RECT 49.950 88.950 52.050 89.400 ;
        RECT 106.950 90.600 109.050 91.050 ;
        RECT 110.400 90.600 111.600 91.950 ;
        RECT 106.950 89.400 111.600 90.600 ;
        RECT 143.400 90.600 144.600 91.950 ;
        RECT 154.950 90.600 157.050 91.050 ;
        RECT 143.400 89.400 157.050 90.600 ;
        RECT 106.950 88.950 109.050 89.400 ;
        RECT 154.950 88.950 157.050 89.400 ;
        RECT 220.950 90.600 223.050 91.050 ;
        RECT 238.950 90.600 241.050 91.050 ;
        RECT 244.950 90.600 247.050 91.050 ;
        RECT 220.950 89.400 237.600 90.600 ;
        RECT 220.950 88.950 223.050 89.400 ;
        RECT 190.950 87.600 193.050 88.050 ;
        RECT 232.950 87.600 235.050 88.050 ;
        RECT 190.950 86.400 235.050 87.600 ;
        RECT 236.400 87.600 237.600 89.400 ;
        RECT 238.950 89.400 247.050 90.600 ;
        RECT 238.950 88.950 241.050 89.400 ;
        RECT 244.950 88.950 247.050 89.400 ;
        RECT 250.950 88.950 253.050 91.050 ;
        RECT 299.400 90.600 300.600 91.950 ;
        RECT 340.950 90.600 343.050 91.050 ;
        RECT 299.400 89.400 343.050 90.600 ;
        RECT 340.950 88.950 343.050 89.400 ;
        RECT 343.950 90.600 346.050 91.050 ;
        RECT 349.950 90.600 352.050 91.050 ;
        RECT 343.950 89.400 352.050 90.600 ;
        RECT 343.950 88.950 346.050 89.400 ;
        RECT 349.950 88.950 352.050 89.400 ;
        RECT 370.950 90.600 373.050 91.050 ;
        RECT 428.400 90.600 429.600 91.950 ;
        RECT 370.950 89.400 429.600 90.600 ;
        RECT 436.950 90.600 439.050 91.050 ;
        RECT 442.950 90.600 445.050 91.050 ;
        RECT 436.950 89.400 445.050 90.600 ;
        RECT 449.400 90.600 450.600 94.950 ;
        RECT 451.950 93.600 454.050 94.050 ;
        RECT 460.950 93.600 463.050 94.050 ;
        RECT 451.950 92.400 463.050 93.600 ;
        RECT 451.950 91.950 454.050 92.400 ;
        RECT 460.950 91.950 463.050 92.400 ;
        RECT 463.950 93.600 466.050 94.050 ;
        RECT 469.950 93.600 472.050 94.050 ;
        RECT 463.950 92.400 472.050 93.600 ;
        RECT 463.950 91.950 466.050 92.400 ;
        RECT 469.950 91.950 472.050 92.400 ;
        RECT 481.950 93.600 484.050 94.050 ;
        RECT 487.950 93.600 490.050 94.050 ;
        RECT 481.950 92.400 490.050 93.600 ;
        RECT 481.950 91.950 484.050 92.400 ;
        RECT 487.950 91.950 490.050 92.400 ;
        RECT 493.950 93.600 496.050 94.050 ;
        RECT 499.950 93.600 502.050 94.050 ;
        RECT 493.950 92.400 502.050 93.600 ;
        RECT 493.950 91.950 496.050 92.400 ;
        RECT 499.950 91.950 502.050 92.400 ;
        RECT 508.950 93.600 511.050 94.050 ;
        RECT 523.950 93.600 526.050 94.050 ;
        RECT 508.950 92.400 526.050 93.600 ;
        RECT 508.950 91.950 511.050 92.400 ;
        RECT 523.950 91.950 526.050 92.400 ;
        RECT 538.950 93.600 541.050 94.050 ;
        RECT 544.950 93.600 547.050 94.050 ;
        RECT 538.950 92.400 547.050 93.600 ;
        RECT 538.950 91.950 541.050 92.400 ;
        RECT 544.950 91.950 547.050 92.400 ;
        RECT 451.950 90.600 454.050 91.050 ;
        RECT 449.400 89.400 454.050 90.600 ;
        RECT 370.950 88.950 373.050 89.400 ;
        RECT 436.950 88.950 439.050 89.400 ;
        RECT 442.950 88.950 445.050 89.400 ;
        RECT 451.950 88.950 454.050 89.400 ;
        RECT 484.950 90.600 487.050 91.050 ;
        RECT 496.950 90.600 499.050 91.050 ;
        RECT 484.950 89.400 499.050 90.600 ;
        RECT 484.950 88.950 487.050 89.400 ;
        RECT 496.950 88.950 499.050 89.400 ;
        RECT 502.950 90.600 505.050 91.050 ;
        RECT 526.950 90.600 529.050 91.050 ;
        RECT 502.950 89.400 529.050 90.600 ;
        RECT 502.950 88.950 505.050 89.400 ;
        RECT 526.950 88.950 529.050 89.400 ;
        RECT 541.950 90.600 544.050 91.050 ;
        RECT 548.400 90.600 549.600 94.950 ;
        RECT 574.950 91.950 577.050 94.050 ;
        RECT 610.950 93.600 613.050 94.050 ;
        RECT 619.950 93.600 622.050 94.050 ;
        RECT 610.950 92.400 622.050 93.600 ;
        RECT 610.950 91.950 613.050 92.400 ;
        RECT 619.950 91.950 622.050 92.400 ;
        RECT 541.950 89.400 549.600 90.600 ;
        RECT 559.950 90.600 562.050 91.050 ;
        RECT 575.400 90.600 576.600 91.950 ;
        RECT 559.950 89.400 576.600 90.600 ;
        RECT 589.950 90.600 592.050 91.050 ;
        RECT 613.950 90.600 616.050 91.050 ;
        RECT 589.950 89.400 616.050 90.600 ;
        RECT 623.400 90.600 624.600 95.400 ;
        RECT 628.950 95.400 637.050 96.600 ;
        RECT 628.950 94.950 631.050 95.400 ;
        RECT 634.950 94.950 637.050 95.400 ;
        RECT 649.950 96.600 652.050 97.050 ;
        RECT 661.950 96.600 664.050 97.050 ;
        RECT 649.950 95.400 664.050 96.600 ;
        RECT 649.950 94.950 652.050 95.400 ;
        RECT 661.950 94.950 664.050 95.400 ;
        RECT 664.950 96.600 667.050 97.050 ;
        RECT 676.950 96.600 679.050 97.050 ;
        RECT 664.950 95.400 679.050 96.600 ;
        RECT 664.950 94.950 667.050 95.400 ;
        RECT 676.950 94.950 679.050 95.400 ;
        RECT 688.950 96.600 691.050 97.050 ;
        RECT 739.950 96.600 742.050 97.050 ;
        RECT 688.950 95.400 742.050 96.600 ;
        RECT 688.950 94.950 691.050 95.400 ;
        RECT 739.950 94.950 742.050 95.400 ;
        RECT 781.950 96.600 784.050 97.050 ;
        RECT 787.950 96.600 790.050 97.050 ;
        RECT 835.950 96.600 838.050 97.050 ;
        RECT 781.950 95.400 790.050 96.600 ;
        RECT 781.950 94.950 784.050 95.400 ;
        RECT 787.950 94.950 790.050 95.400 ;
        RECT 803.400 95.400 838.050 96.600 ;
        RECT 803.400 94.050 804.600 95.400 ;
        RECT 835.950 94.950 838.050 95.400 ;
        RECT 625.950 93.600 628.050 94.050 ;
        RECT 640.950 93.600 643.050 94.050 ;
        RECT 625.950 92.400 643.050 93.600 ;
        RECT 625.950 91.950 628.050 92.400 ;
        RECT 640.950 91.950 643.050 92.400 ;
        RECT 706.950 93.600 709.050 94.050 ;
        RECT 724.950 93.600 727.050 94.050 ;
        RECT 706.950 92.400 727.050 93.600 ;
        RECT 706.950 91.950 709.050 92.400 ;
        RECT 724.950 91.950 727.050 92.400 ;
        RECT 730.950 93.600 733.050 94.050 ;
        RECT 763.950 93.600 766.050 94.050 ;
        RECT 778.950 93.600 781.050 94.050 ;
        RECT 796.950 93.600 799.050 94.050 ;
        RECT 730.950 92.400 799.050 93.600 ;
        RECT 730.950 91.950 733.050 92.400 ;
        RECT 763.950 91.950 766.050 92.400 ;
        RECT 778.950 91.950 781.050 92.400 ;
        RECT 796.950 91.950 799.050 92.400 ;
        RECT 802.950 91.950 805.050 94.050 ;
        RECT 625.950 90.600 628.050 91.050 ;
        RECT 623.400 89.400 628.050 90.600 ;
        RECT 541.950 88.950 544.050 89.400 ;
        RECT 559.950 88.950 562.050 89.400 ;
        RECT 589.950 88.950 592.050 89.400 ;
        RECT 613.950 88.950 616.050 89.400 ;
        RECT 625.950 88.950 628.050 89.400 ;
        RECT 652.950 90.600 655.050 91.050 ;
        RECT 667.950 90.600 670.050 91.050 ;
        RECT 736.950 90.600 739.050 91.050 ;
        RECT 652.950 89.400 739.050 90.600 ;
        RECT 652.950 88.950 655.050 89.400 ;
        RECT 667.950 88.950 670.050 89.400 ;
        RECT 736.950 88.950 739.050 89.400 ;
        RECT 748.950 90.600 751.050 91.050 ;
        RECT 766.950 90.600 769.050 91.050 ;
        RECT 808.950 90.600 811.050 91.050 ;
        RECT 748.950 89.400 811.050 90.600 ;
        RECT 748.950 88.950 751.050 89.400 ;
        RECT 766.950 88.950 769.050 89.400 ;
        RECT 808.950 88.950 811.050 89.400 ;
        RECT 251.400 87.600 252.600 88.950 ;
        RECT 236.400 86.400 252.600 87.600 ;
        RECT 259.950 87.600 262.050 88.050 ;
        RECT 283.950 87.600 286.050 88.050 ;
        RECT 259.950 86.400 286.050 87.600 ;
        RECT 190.950 85.950 193.050 86.400 ;
        RECT 232.950 85.950 235.050 86.400 ;
        RECT 259.950 85.950 262.050 86.400 ;
        RECT 283.950 85.950 286.050 86.400 ;
        RECT 298.950 87.600 301.050 88.050 ;
        RECT 439.950 87.600 442.050 88.050 ;
        RECT 298.950 86.400 442.050 87.600 ;
        RECT 298.950 85.950 301.050 86.400 ;
        RECT 439.950 85.950 442.050 86.400 ;
        RECT 478.950 87.600 481.050 88.050 ;
        RECT 523.950 87.600 526.050 88.050 ;
        RECT 478.950 86.400 526.050 87.600 ;
        RECT 478.950 85.950 481.050 86.400 ;
        RECT 523.950 85.950 526.050 86.400 ;
        RECT 547.950 87.600 550.050 88.050 ;
        RECT 562.950 87.600 565.050 88.050 ;
        RECT 547.950 86.400 565.050 87.600 ;
        RECT 547.950 85.950 550.050 86.400 ;
        RECT 562.950 85.950 565.050 86.400 ;
        RECT 583.950 87.600 586.050 88.050 ;
        RECT 595.950 87.600 598.050 88.050 ;
        RECT 583.950 86.400 598.050 87.600 ;
        RECT 583.950 85.950 586.050 86.400 ;
        RECT 595.950 85.950 598.050 86.400 ;
        RECT 601.950 87.600 604.050 88.050 ;
        RECT 607.950 87.600 610.050 88.050 ;
        RECT 601.950 86.400 610.050 87.600 ;
        RECT 601.950 85.950 604.050 86.400 ;
        RECT 607.950 85.950 610.050 86.400 ;
        RECT 631.950 87.600 634.050 88.050 ;
        RECT 673.950 87.600 676.050 88.050 ;
        RECT 631.950 86.400 676.050 87.600 ;
        RECT 631.950 85.950 634.050 86.400 ;
        RECT 673.950 85.950 676.050 86.400 ;
        RECT 682.950 87.600 685.050 88.050 ;
        RECT 688.950 87.600 691.050 88.050 ;
        RECT 697.950 87.600 700.050 88.050 ;
        RECT 682.950 86.400 700.050 87.600 ;
        RECT 682.950 85.950 685.050 86.400 ;
        RECT 688.950 85.950 691.050 86.400 ;
        RECT 697.950 85.950 700.050 86.400 ;
        RECT 10.950 84.600 13.050 85.050 ;
        RECT 70.950 84.600 73.050 85.050 ;
        RECT 10.950 83.400 73.050 84.600 ;
        RECT 10.950 82.950 13.050 83.400 ;
        RECT 70.950 82.950 73.050 83.400 ;
        RECT 133.950 84.600 136.050 85.050 ;
        RECT 208.950 84.600 211.050 85.050 ;
        RECT 133.950 83.400 211.050 84.600 ;
        RECT 133.950 82.950 136.050 83.400 ;
        RECT 208.950 82.950 211.050 83.400 ;
        RECT 214.950 84.600 217.050 85.050 ;
        RECT 268.950 84.600 271.050 85.050 ;
        RECT 358.950 84.600 361.050 85.050 ;
        RECT 463.950 84.600 466.050 85.050 ;
        RECT 214.950 83.400 466.050 84.600 ;
        RECT 214.950 82.950 217.050 83.400 ;
        RECT 268.950 82.950 271.050 83.400 ;
        RECT 358.950 82.950 361.050 83.400 ;
        RECT 463.950 82.950 466.050 83.400 ;
        RECT 526.950 84.600 529.050 85.050 ;
        RECT 538.950 84.600 541.050 85.050 ;
        RECT 526.950 83.400 541.050 84.600 ;
        RECT 526.950 82.950 529.050 83.400 ;
        RECT 538.950 82.950 541.050 83.400 ;
        RECT 565.950 84.600 568.050 85.050 ;
        RECT 634.950 84.600 637.050 85.050 ;
        RECT 565.950 83.400 637.050 84.600 ;
        RECT 565.950 82.950 568.050 83.400 ;
        RECT 634.950 82.950 637.050 83.400 ;
        RECT 43.950 81.600 46.050 82.050 ;
        RECT 52.950 81.600 55.050 82.050 ;
        RECT 43.950 80.400 55.050 81.600 ;
        RECT 43.950 79.950 46.050 80.400 ;
        RECT 52.950 79.950 55.050 80.400 ;
        RECT 250.950 81.600 253.050 82.050 ;
        RECT 256.950 81.600 259.050 82.050 ;
        RECT 250.950 80.400 259.050 81.600 ;
        RECT 250.950 79.950 253.050 80.400 ;
        RECT 256.950 79.950 259.050 80.400 ;
        RECT 310.950 81.600 313.050 82.050 ;
        RECT 322.950 81.600 325.050 82.050 ;
        RECT 310.950 80.400 325.050 81.600 ;
        RECT 310.950 79.950 313.050 80.400 ;
        RECT 322.950 79.950 325.050 80.400 ;
        RECT 325.950 81.600 328.050 82.050 ;
        RECT 373.950 81.600 376.050 82.050 ;
        RECT 385.950 81.600 388.050 82.050 ;
        RECT 325.950 80.400 388.050 81.600 ;
        RECT 325.950 79.950 328.050 80.400 ;
        RECT 373.950 79.950 376.050 80.400 ;
        RECT 385.950 79.950 388.050 80.400 ;
        RECT 388.950 81.600 391.050 82.050 ;
        RECT 538.950 81.600 541.050 82.050 ;
        RECT 388.950 80.400 541.050 81.600 ;
        RECT 388.950 79.950 391.050 80.400 ;
        RECT 538.950 79.950 541.050 80.400 ;
        RECT 547.950 81.600 550.050 82.050 ;
        RECT 679.950 81.600 682.050 82.050 ;
        RECT 742.950 81.600 745.050 82.050 ;
        RECT 751.950 81.600 754.050 82.050 ;
        RECT 547.950 80.400 754.050 81.600 ;
        RECT 547.950 79.950 550.050 80.400 ;
        RECT 679.950 79.950 682.050 80.400 ;
        RECT 742.950 79.950 745.050 80.400 ;
        RECT 751.950 79.950 754.050 80.400 ;
        RECT 283.950 78.600 286.050 79.050 ;
        RECT 379.950 78.600 382.050 79.050 ;
        RECT 391.950 78.600 394.050 79.050 ;
        RECT 283.950 77.400 394.050 78.600 ;
        RECT 283.950 76.950 286.050 77.400 ;
        RECT 379.950 76.950 382.050 77.400 ;
        RECT 391.950 76.950 394.050 77.400 ;
        RECT 418.950 78.600 421.050 79.050 ;
        RECT 442.950 78.600 445.050 79.050 ;
        RECT 418.950 77.400 445.050 78.600 ;
        RECT 418.950 76.950 421.050 77.400 ;
        RECT 442.950 76.950 445.050 77.400 ;
        RECT 532.950 78.600 535.050 79.050 ;
        RECT 559.950 78.600 562.050 79.050 ;
        RECT 532.950 77.400 562.050 78.600 ;
        RECT 532.950 76.950 535.050 77.400 ;
        RECT 559.950 76.950 562.050 77.400 ;
        RECT 562.950 78.600 565.050 79.050 ;
        RECT 730.950 78.600 733.050 79.050 ;
        RECT 562.950 77.400 733.050 78.600 ;
        RECT 562.950 76.950 565.050 77.400 ;
        RECT 730.950 76.950 733.050 77.400 ;
        RECT 46.950 75.600 49.050 76.050 ;
        RECT 58.950 75.600 61.050 76.050 ;
        RECT 235.950 75.600 238.050 76.050 ;
        RECT 367.950 75.600 370.050 76.050 ;
        RECT 388.950 75.600 391.050 76.050 ;
        RECT 46.950 74.400 391.050 75.600 ;
        RECT 46.950 73.950 49.050 74.400 ;
        RECT 58.950 73.950 61.050 74.400 ;
        RECT 235.950 73.950 238.050 74.400 ;
        RECT 367.950 73.950 370.050 74.400 ;
        RECT 388.950 73.950 391.050 74.400 ;
        RECT 394.950 75.600 397.050 76.050 ;
        RECT 433.950 75.600 436.050 76.050 ;
        RECT 469.950 75.600 472.050 76.050 ;
        RECT 394.950 74.400 472.050 75.600 ;
        RECT 394.950 73.950 397.050 74.400 ;
        RECT 433.950 73.950 436.050 74.400 ;
        RECT 469.950 73.950 472.050 74.400 ;
        RECT 586.950 75.600 589.050 76.050 ;
        RECT 646.950 75.600 649.050 76.050 ;
        RECT 694.950 75.600 697.050 76.050 ;
        RECT 586.950 74.400 697.050 75.600 ;
        RECT 586.950 73.950 589.050 74.400 ;
        RECT 646.950 73.950 649.050 74.400 ;
        RECT 694.950 73.950 697.050 74.400 ;
        RECT 280.950 72.600 283.050 73.050 ;
        RECT 460.950 72.600 463.050 73.050 ;
        RECT 280.950 71.400 463.050 72.600 ;
        RECT 280.950 70.950 283.050 71.400 ;
        RECT 460.950 70.950 463.050 71.400 ;
        RECT 772.950 72.600 775.050 73.050 ;
        RECT 778.950 72.600 781.050 73.050 ;
        RECT 772.950 71.400 781.050 72.600 ;
        RECT 772.950 70.950 775.050 71.400 ;
        RECT 778.950 70.950 781.050 71.400 ;
        RECT 304.950 69.600 307.050 70.050 ;
        RECT 355.950 69.600 358.050 70.050 ;
        RECT 304.950 68.400 358.050 69.600 ;
        RECT 304.950 67.950 307.050 68.400 ;
        RECT 355.950 67.950 358.050 68.400 ;
        RECT 364.950 69.600 367.050 70.050 ;
        RECT 412.950 69.600 415.050 70.050 ;
        RECT 364.950 68.400 415.050 69.600 ;
        RECT 364.950 67.950 367.050 68.400 ;
        RECT 412.950 67.950 415.050 68.400 ;
        RECT 430.950 69.600 433.050 70.050 ;
        RECT 445.950 69.600 448.050 70.050 ;
        RECT 469.950 69.600 472.050 70.050 ;
        RECT 430.950 68.400 472.050 69.600 ;
        RECT 430.950 67.950 433.050 68.400 ;
        RECT 445.950 67.950 448.050 68.400 ;
        RECT 469.950 67.950 472.050 68.400 ;
        RECT 700.950 69.600 703.050 70.050 ;
        RECT 709.950 69.600 712.050 70.050 ;
        RECT 715.950 69.600 718.050 70.050 ;
        RECT 700.950 68.400 718.050 69.600 ;
        RECT 700.950 67.950 703.050 68.400 ;
        RECT 709.950 67.950 712.050 68.400 ;
        RECT 715.950 67.950 718.050 68.400 ;
        RECT 97.950 66.600 100.050 67.050 ;
        RECT 109.950 66.600 112.050 67.050 ;
        RECT 118.950 66.600 121.050 67.050 ;
        RECT 124.950 66.600 127.050 67.050 ;
        RECT 97.950 65.400 127.050 66.600 ;
        RECT 97.950 64.950 100.050 65.400 ;
        RECT 109.950 64.950 112.050 65.400 ;
        RECT 118.950 64.950 121.050 65.400 ;
        RECT 124.950 64.950 127.050 65.400 ;
        RECT 178.950 66.600 181.050 67.050 ;
        RECT 187.950 66.600 190.050 67.050 ;
        RECT 226.950 66.600 229.050 67.050 ;
        RECT 256.950 66.600 259.050 67.050 ;
        RECT 265.950 66.600 268.050 67.050 ;
        RECT 364.950 66.600 367.050 67.050 ;
        RECT 439.950 66.600 442.050 67.050 ;
        RECT 508.950 66.600 511.050 67.050 ;
        RECT 178.950 65.400 511.050 66.600 ;
        RECT 178.950 64.950 181.050 65.400 ;
        RECT 187.950 64.950 190.050 65.400 ;
        RECT 226.950 64.950 229.050 65.400 ;
        RECT 256.950 64.950 259.050 65.400 ;
        RECT 265.950 64.950 268.050 65.400 ;
        RECT 364.950 64.950 367.050 65.400 ;
        RECT 439.950 64.950 442.050 65.400 ;
        RECT 508.950 64.950 511.050 65.400 ;
        RECT 529.950 66.600 532.050 67.050 ;
        RECT 604.950 66.600 607.050 67.050 ;
        RECT 619.950 66.600 622.050 67.050 ;
        RECT 529.950 65.400 622.050 66.600 ;
        RECT 529.950 64.950 532.050 65.400 ;
        RECT 604.950 64.950 607.050 65.400 ;
        RECT 619.950 64.950 622.050 65.400 ;
        RECT 658.950 66.600 661.050 67.050 ;
        RECT 772.950 66.600 775.050 67.050 ;
        RECT 658.950 65.400 775.050 66.600 ;
        RECT 658.950 64.950 661.050 65.400 ;
        RECT 772.950 64.950 775.050 65.400 ;
        RECT 97.950 63.600 100.050 64.050 ;
        RECT 253.950 63.600 256.050 64.050 ;
        RECT 466.950 63.600 469.050 64.050 ;
        RECT 478.950 63.600 481.050 64.050 ;
        RECT 97.950 62.400 481.050 63.600 ;
        RECT 97.950 61.950 100.050 62.400 ;
        RECT 253.950 61.950 256.050 62.400 ;
        RECT 466.950 61.950 469.050 62.400 ;
        RECT 478.950 61.950 481.050 62.400 ;
        RECT 70.950 60.600 73.050 61.050 ;
        RECT 85.950 60.600 88.050 61.050 ;
        RECT 97.950 60.600 100.050 61.050 ;
        RECT 70.950 59.400 100.050 60.600 ;
        RECT 70.950 58.950 73.050 59.400 ;
        RECT 85.950 58.950 88.050 59.400 ;
        RECT 97.950 58.950 100.050 59.400 ;
        RECT 103.950 60.600 106.050 61.050 ;
        RECT 145.950 60.600 148.050 61.050 ;
        RECT 103.950 59.400 148.050 60.600 ;
        RECT 103.950 58.950 106.050 59.400 ;
        RECT 145.950 58.950 148.050 59.400 ;
        RECT 232.950 60.600 235.050 61.050 ;
        RECT 265.950 60.600 268.050 61.050 ;
        RECT 232.950 59.400 268.050 60.600 ;
        RECT 232.950 58.950 235.050 59.400 ;
        RECT 265.950 58.950 268.050 59.400 ;
        RECT 286.950 60.600 289.050 61.050 ;
        RECT 295.950 60.600 298.050 61.050 ;
        RECT 286.950 59.400 298.050 60.600 ;
        RECT 286.950 58.950 289.050 59.400 ;
        RECT 295.950 58.950 298.050 59.400 ;
        RECT 319.950 60.600 322.050 61.050 ;
        RECT 328.950 60.600 331.050 61.050 ;
        RECT 319.950 59.400 331.050 60.600 ;
        RECT 319.950 58.950 322.050 59.400 ;
        RECT 328.950 58.950 331.050 59.400 ;
        RECT 355.950 60.600 358.050 61.050 ;
        RECT 355.950 59.400 432.600 60.600 ;
        RECT 355.950 58.950 358.050 59.400 ;
        RECT 67.950 57.600 70.050 58.050 ;
        RECT 115.950 57.600 118.050 58.050 ;
        RECT 130.950 57.600 133.050 58.050 ;
        RECT 67.950 56.400 99.600 57.600 ;
        RECT 67.950 55.950 70.050 56.400 ;
        RECT 76.950 54.600 79.050 55.050 ;
        RECT 85.950 54.600 88.050 55.050 ;
        RECT 76.950 53.400 88.050 54.600 ;
        RECT 98.400 54.600 99.600 56.400 ;
        RECT 115.950 56.400 133.050 57.600 ;
        RECT 115.950 55.950 118.050 56.400 ;
        RECT 130.950 55.950 133.050 56.400 ;
        RECT 148.950 57.600 151.050 58.050 ;
        RECT 160.950 57.600 163.050 58.050 ;
        RECT 148.950 56.400 163.050 57.600 ;
        RECT 148.950 55.950 151.050 56.400 ;
        RECT 160.950 55.950 163.050 56.400 ;
        RECT 205.950 57.600 208.050 58.050 ;
        RECT 217.950 57.600 220.050 58.050 ;
        RECT 205.950 56.400 220.050 57.600 ;
        RECT 205.950 55.950 208.050 56.400 ;
        RECT 217.950 55.950 220.050 56.400 ;
        RECT 247.950 55.950 250.050 58.050 ;
        RECT 265.950 57.600 268.050 58.050 ;
        RECT 310.950 57.600 313.050 58.050 ;
        RECT 346.950 57.600 349.050 58.050 ;
        RECT 361.950 57.600 364.050 58.050 ;
        RECT 265.950 56.400 313.050 57.600 ;
        RECT 265.950 55.950 268.050 56.400 ;
        RECT 310.950 55.950 313.050 56.400 ;
        RECT 323.400 56.400 349.050 57.600 ;
        RECT 175.950 54.600 178.050 55.050 ;
        RECT 202.950 54.600 205.050 55.050 ;
        RECT 208.950 54.600 211.050 55.050 ;
        RECT 98.400 53.400 192.600 54.600 ;
        RECT 76.950 52.950 79.050 53.400 ;
        RECT 85.950 52.950 88.050 53.400 ;
        RECT 175.950 52.950 178.050 53.400 ;
        RECT 79.950 51.600 82.050 52.050 ;
        RECT 100.950 51.600 103.050 52.050 ;
        RECT 145.950 51.600 148.050 52.050 ;
        RECT 151.950 51.600 154.050 52.050 ;
        RECT 79.950 50.400 103.050 51.600 ;
        RECT 79.950 49.950 82.050 50.400 ;
        RECT 100.950 49.950 103.050 50.400 ;
        RECT 104.400 50.400 154.050 51.600 ;
        RECT 28.950 48.600 31.050 49.050 ;
        RECT 82.950 48.600 85.050 49.050 ;
        RECT 28.950 47.400 85.050 48.600 ;
        RECT 28.950 46.950 31.050 47.400 ;
        RECT 82.950 46.950 85.050 47.400 ;
        RECT 88.950 48.600 91.050 49.050 ;
        RECT 104.400 48.600 105.600 50.400 ;
        RECT 145.950 49.950 148.050 50.400 ;
        RECT 151.950 49.950 154.050 50.400 ;
        RECT 157.950 51.600 160.050 52.050 ;
        RECT 172.950 51.600 175.050 52.050 ;
        RECT 178.950 51.600 181.050 52.050 ;
        RECT 187.950 51.600 190.050 52.050 ;
        RECT 157.950 50.400 177.600 51.600 ;
        RECT 157.950 49.950 160.050 50.400 ;
        RECT 172.950 49.950 175.050 50.400 ;
        RECT 88.950 47.400 105.600 48.600 ;
        RECT 136.950 48.600 139.050 49.050 ;
        RECT 145.950 48.600 148.050 49.050 ;
        RECT 163.950 48.600 166.050 49.050 ;
        RECT 172.950 48.600 175.050 49.050 ;
        RECT 136.950 47.400 175.050 48.600 ;
        RECT 176.400 48.600 177.600 50.400 ;
        RECT 178.950 50.400 190.050 51.600 ;
        RECT 191.400 51.600 192.600 53.400 ;
        RECT 202.950 53.400 211.050 54.600 ;
        RECT 202.950 52.950 205.050 53.400 ;
        RECT 208.950 52.950 211.050 53.400 ;
        RECT 214.950 54.600 217.050 55.050 ;
        RECT 220.950 54.600 223.050 55.050 ;
        RECT 241.950 54.600 244.050 55.050 ;
        RECT 214.950 53.400 244.050 54.600 ;
        RECT 214.950 52.950 217.050 53.400 ;
        RECT 220.950 52.950 223.050 53.400 ;
        RECT 241.950 52.950 244.050 53.400 ;
        RECT 248.400 52.050 249.600 55.950 ;
        RECT 323.400 55.050 324.600 56.400 ;
        RECT 346.950 55.950 349.050 56.400 ;
        RECT 359.400 56.400 364.050 57.600 ;
        RECT 259.950 54.600 262.050 55.050 ;
        RECT 271.950 54.600 274.050 55.050 ;
        RECT 298.950 54.600 301.050 55.050 ;
        RECT 259.950 53.400 270.600 54.600 ;
        RECT 259.950 52.950 262.050 53.400 ;
        RECT 199.950 51.600 202.050 52.050 ;
        RECT 191.400 50.400 202.050 51.600 ;
        RECT 178.950 49.950 181.050 50.400 ;
        RECT 187.950 49.950 190.050 50.400 ;
        RECT 199.950 49.950 202.050 50.400 ;
        RECT 217.950 51.600 220.050 52.050 ;
        RECT 244.950 51.600 247.050 52.050 ;
        RECT 217.950 50.400 247.050 51.600 ;
        RECT 217.950 49.950 220.050 50.400 ;
        RECT 244.950 49.950 247.050 50.400 ;
        RECT 247.950 49.950 250.050 52.050 ;
        RECT 269.400 51.600 270.600 53.400 ;
        RECT 271.950 53.400 301.050 54.600 ;
        RECT 271.950 52.950 274.050 53.400 ;
        RECT 298.950 52.950 301.050 53.400 ;
        RECT 301.950 54.600 304.050 55.050 ;
        RECT 307.950 54.600 310.050 55.050 ;
        RECT 316.950 54.600 319.050 55.050 ;
        RECT 301.950 53.400 319.050 54.600 ;
        RECT 301.950 52.950 304.050 53.400 ;
        RECT 307.950 52.950 310.050 53.400 ;
        RECT 316.950 52.950 319.050 53.400 ;
        RECT 322.950 52.950 325.050 55.050 ;
        RECT 277.950 51.600 280.050 52.050 ;
        RECT 286.950 51.600 289.050 52.050 ;
        RECT 269.400 50.400 289.050 51.600 ;
        RECT 277.950 49.950 280.050 50.400 ;
        RECT 286.950 49.950 289.050 50.400 ;
        RECT 295.950 51.600 298.050 52.050 ;
        RECT 307.950 51.600 310.050 52.050 ;
        RECT 295.950 50.400 310.050 51.600 ;
        RECT 295.950 49.950 298.050 50.400 ;
        RECT 307.950 49.950 310.050 50.400 ;
        RECT 319.950 51.600 322.050 52.050 ;
        RECT 325.950 51.600 328.050 52.050 ;
        RECT 319.950 50.400 328.050 51.600 ;
        RECT 319.950 49.950 322.050 50.400 ;
        RECT 325.950 49.950 328.050 50.400 ;
        RECT 337.950 51.600 340.050 52.050 ;
        RECT 355.950 51.600 358.050 52.050 ;
        RECT 337.950 50.400 358.050 51.600 ;
        RECT 359.400 51.600 360.600 56.400 ;
        RECT 361.950 55.950 364.050 56.400 ;
        RECT 379.950 57.600 382.050 58.050 ;
        RECT 421.950 57.600 424.050 58.050 ;
        RECT 379.950 56.400 424.050 57.600 ;
        RECT 379.950 55.950 382.050 56.400 ;
        RECT 421.950 55.950 424.050 56.400 ;
        RECT 424.950 57.600 427.050 58.050 ;
        RECT 424.950 56.400 429.600 57.600 ;
        RECT 424.950 55.950 427.050 56.400 ;
        RECT 361.950 54.600 364.050 55.050 ;
        RECT 370.950 54.600 373.050 55.050 ;
        RECT 361.950 53.400 373.050 54.600 ;
        RECT 361.950 52.950 364.050 53.400 ;
        RECT 370.950 52.950 373.050 53.400 ;
        RECT 376.950 54.600 379.050 55.050 ;
        RECT 382.950 54.600 385.050 55.050 ;
        RECT 376.950 53.400 385.050 54.600 ;
        RECT 376.950 52.950 379.050 53.400 ;
        RECT 382.950 52.950 385.050 53.400 ;
        RECT 400.950 54.600 403.050 55.050 ;
        RECT 409.950 54.600 412.050 55.050 ;
        RECT 400.950 53.400 412.050 54.600 ;
        RECT 400.950 52.950 403.050 53.400 ;
        RECT 409.950 52.950 412.050 53.400 ;
        RECT 412.950 54.600 415.050 55.050 ;
        RECT 418.950 54.600 421.050 55.050 ;
        RECT 412.950 53.400 421.050 54.600 ;
        RECT 412.950 52.950 415.050 53.400 ;
        RECT 418.950 52.950 421.050 53.400 ;
        RECT 424.950 52.950 427.050 55.050 ;
        RECT 367.950 51.600 370.050 52.050 ;
        RECT 359.400 50.400 370.050 51.600 ;
        RECT 337.950 49.950 340.050 50.400 ;
        RECT 355.950 49.950 358.050 50.400 ;
        RECT 367.950 49.950 370.050 50.400 ;
        RECT 388.950 51.600 391.050 52.050 ;
        RECT 394.950 51.600 397.050 52.050 ;
        RECT 388.950 50.400 397.050 51.600 ;
        RECT 388.950 49.950 391.050 50.400 ;
        RECT 394.950 49.950 397.050 50.400 ;
        RECT 406.950 51.600 409.050 52.050 ;
        RECT 415.950 51.600 418.050 52.050 ;
        RECT 406.950 50.400 418.050 51.600 ;
        RECT 406.950 49.950 409.050 50.400 ;
        RECT 415.950 49.950 418.050 50.400 ;
        RECT 418.950 51.600 421.050 52.050 ;
        RECT 425.400 51.600 426.600 52.950 ;
        RECT 428.400 52.050 429.600 56.400 ;
        RECT 418.950 50.400 426.600 51.600 ;
        RECT 418.950 49.950 421.050 50.400 ;
        RECT 427.950 49.950 430.050 52.050 ;
        RECT 431.400 51.600 432.600 59.400 ;
        RECT 433.950 58.950 436.050 61.050 ;
        RECT 442.950 60.600 445.050 61.050 ;
        RECT 490.950 60.600 493.050 61.050 ;
        RECT 553.950 60.600 556.050 61.050 ;
        RECT 601.950 60.600 604.050 61.050 ;
        RECT 442.950 59.400 604.050 60.600 ;
        RECT 442.950 58.950 445.050 59.400 ;
        RECT 490.950 58.950 493.050 59.400 ;
        RECT 553.950 58.950 556.050 59.400 ;
        RECT 601.950 58.950 604.050 59.400 ;
        RECT 610.950 60.600 613.050 61.050 ;
        RECT 661.950 60.600 664.050 61.050 ;
        RECT 682.950 60.600 685.050 61.050 ;
        RECT 841.950 60.600 844.050 61.050 ;
        RECT 610.950 59.400 844.050 60.600 ;
        RECT 610.950 58.950 613.050 59.400 ;
        RECT 661.950 58.950 664.050 59.400 ;
        RECT 682.950 58.950 685.050 59.400 ;
        RECT 841.950 58.950 844.050 59.400 ;
        RECT 434.400 55.050 435.600 58.950 ;
        RECT 436.950 57.600 439.050 58.050 ;
        RECT 445.950 57.600 448.050 58.050 ;
        RECT 436.950 56.400 448.050 57.600 ;
        RECT 436.950 55.950 439.050 56.400 ;
        RECT 445.950 55.950 448.050 56.400 ;
        RECT 469.950 57.600 472.050 58.050 ;
        RECT 505.950 57.600 508.050 58.050 ;
        RECT 511.950 57.600 514.050 58.050 ;
        RECT 469.950 56.400 514.050 57.600 ;
        RECT 469.950 55.950 472.050 56.400 ;
        RECT 505.950 55.950 508.050 56.400 ;
        RECT 511.950 55.950 514.050 56.400 ;
        RECT 538.950 57.600 541.050 58.050 ;
        RECT 706.950 57.600 709.050 58.050 ;
        RECT 721.950 57.600 724.050 58.050 ;
        RECT 538.950 56.400 561.600 57.600 ;
        RECT 538.950 55.950 541.050 56.400 ;
        RECT 560.400 55.050 561.600 56.400 ;
        RECT 706.950 56.400 724.050 57.600 ;
        RECT 706.950 55.950 709.050 56.400 ;
        RECT 721.950 55.950 724.050 56.400 ;
        RECT 841.950 57.600 844.050 58.050 ;
        RECT 853.950 57.600 856.050 58.050 ;
        RECT 841.950 56.400 856.050 57.600 ;
        RECT 841.950 55.950 844.050 56.400 ;
        RECT 853.950 55.950 856.050 56.400 ;
        RECT 433.950 52.950 436.050 55.050 ;
        RECT 439.950 54.600 442.050 55.050 ;
        RECT 457.950 54.600 460.050 55.050 ;
        RECT 439.950 53.400 460.050 54.600 ;
        RECT 439.950 52.950 442.050 53.400 ;
        RECT 457.950 52.950 460.050 53.400 ;
        RECT 460.950 54.600 463.050 55.050 ;
        RECT 463.950 54.600 466.050 55.050 ;
        RECT 469.950 54.600 472.050 55.050 ;
        RECT 502.950 54.600 505.050 55.050 ;
        RECT 460.950 53.400 472.050 54.600 ;
        RECT 460.950 52.950 463.050 53.400 ;
        RECT 463.950 52.950 466.050 53.400 ;
        RECT 469.950 52.950 472.050 53.400 ;
        RECT 491.400 53.400 505.050 54.600 ;
        RECT 448.950 51.600 451.050 52.050 ;
        RECT 431.400 50.400 451.050 51.600 ;
        RECT 448.950 49.950 451.050 50.400 ;
        RECT 475.950 51.600 478.050 52.050 ;
        RECT 491.400 51.600 492.600 53.400 ;
        RECT 502.950 52.950 505.050 53.400 ;
        RECT 511.950 54.600 514.050 55.050 ;
        RECT 547.950 54.600 550.050 55.050 ;
        RECT 511.950 53.400 550.050 54.600 ;
        RECT 511.950 52.950 514.050 53.400 ;
        RECT 547.950 52.950 550.050 53.400 ;
        RECT 559.950 54.600 562.050 55.050 ;
        RECT 601.950 54.600 604.050 55.050 ;
        RECT 559.950 53.400 604.050 54.600 ;
        RECT 559.950 52.950 562.050 53.400 ;
        RECT 601.950 52.950 604.050 53.400 ;
        RECT 619.950 54.600 622.050 55.050 ;
        RECT 673.950 54.600 676.050 55.050 ;
        RECT 619.950 53.400 676.050 54.600 ;
        RECT 619.950 52.950 622.050 53.400 ;
        RECT 673.950 52.950 676.050 53.400 ;
        RECT 700.950 54.600 703.050 55.050 ;
        RECT 709.950 54.600 712.050 55.050 ;
        RECT 700.950 53.400 712.050 54.600 ;
        RECT 700.950 52.950 703.050 53.400 ;
        RECT 709.950 52.950 712.050 53.400 ;
        RECT 730.950 54.600 733.050 55.050 ;
        RECT 745.950 54.600 748.050 55.050 ;
        RECT 757.950 54.600 760.050 55.050 ;
        RECT 790.950 54.600 793.050 55.050 ;
        RECT 796.950 54.600 799.050 55.050 ;
        RECT 730.950 53.400 799.050 54.600 ;
        RECT 730.950 52.950 733.050 53.400 ;
        RECT 745.950 52.950 748.050 53.400 ;
        RECT 757.950 52.950 760.050 53.400 ;
        RECT 790.950 52.950 793.050 53.400 ;
        RECT 796.950 52.950 799.050 53.400 ;
        RECT 475.950 50.400 492.600 51.600 ;
        RECT 493.950 51.600 496.050 52.050 ;
        RECT 541.950 51.600 544.050 52.050 ;
        RECT 550.950 51.600 553.050 52.050 ;
        RECT 493.950 50.400 553.050 51.600 ;
        RECT 475.950 49.950 478.050 50.400 ;
        RECT 493.950 49.950 496.050 50.400 ;
        RECT 541.950 49.950 544.050 50.400 ;
        RECT 550.950 49.950 553.050 50.400 ;
        RECT 727.950 51.600 730.050 52.050 ;
        RECT 769.950 51.600 772.050 52.050 ;
        RECT 727.950 50.400 772.050 51.600 ;
        RECT 727.950 49.950 730.050 50.400 ;
        RECT 769.950 49.950 772.050 50.400 ;
        RECT 181.950 48.600 184.050 49.050 ;
        RECT 176.400 47.400 184.050 48.600 ;
        RECT 88.950 46.950 91.050 47.400 ;
        RECT 136.950 46.950 139.050 47.400 ;
        RECT 145.950 46.950 148.050 47.400 ;
        RECT 163.950 46.950 166.050 47.400 ;
        RECT 172.950 46.950 175.050 47.400 ;
        RECT 181.950 46.950 184.050 47.400 ;
        RECT 196.950 48.600 199.050 49.050 ;
        RECT 214.950 48.600 217.050 49.050 ;
        RECT 196.950 47.400 217.050 48.600 ;
        RECT 196.950 46.950 199.050 47.400 ;
        RECT 214.950 46.950 217.050 47.400 ;
        RECT 217.950 48.600 220.050 49.050 ;
        RECT 223.950 48.600 226.050 49.050 ;
        RECT 217.950 47.400 226.050 48.600 ;
        RECT 217.950 46.950 220.050 47.400 ;
        RECT 223.950 46.950 226.050 47.400 ;
        RECT 238.950 48.600 241.050 49.050 ;
        RECT 256.950 48.600 259.050 49.050 ;
        RECT 238.950 47.400 259.050 48.600 ;
        RECT 238.950 46.950 241.050 47.400 ;
        RECT 256.950 46.950 259.050 47.400 ;
        RECT 286.950 48.600 289.050 49.050 ;
        RECT 352.950 48.600 355.050 49.050 ;
        RECT 373.950 48.600 376.050 49.050 ;
        RECT 379.950 48.600 382.050 49.050 ;
        RECT 448.950 48.600 451.050 49.050 ;
        RECT 286.950 47.400 451.050 48.600 ;
        RECT 286.950 46.950 289.050 47.400 ;
        RECT 352.950 46.950 355.050 47.400 ;
        RECT 373.950 46.950 376.050 47.400 ;
        RECT 379.950 46.950 382.050 47.400 ;
        RECT 448.950 46.950 451.050 47.400 ;
        RECT 481.950 48.600 484.050 49.050 ;
        RECT 502.950 48.600 505.050 49.050 ;
        RECT 586.950 48.600 589.050 49.050 ;
        RECT 481.950 47.400 492.600 48.600 ;
        RECT 481.950 46.950 484.050 47.400 ;
        RECT 491.400 46.050 492.600 47.400 ;
        RECT 502.950 47.400 589.050 48.600 ;
        RECT 502.950 46.950 505.050 47.400 ;
        RECT 586.950 46.950 589.050 47.400 ;
        RECT 631.950 48.600 634.050 49.050 ;
        RECT 730.950 48.600 733.050 49.050 ;
        RECT 631.950 47.400 733.050 48.600 ;
        RECT 631.950 46.950 634.050 47.400 ;
        RECT 730.950 46.950 733.050 47.400 ;
        RECT 760.950 48.600 763.050 49.050 ;
        RECT 817.950 48.600 820.050 49.050 ;
        RECT 760.950 47.400 820.050 48.600 ;
        RECT 760.950 46.950 763.050 47.400 ;
        RECT 817.950 46.950 820.050 47.400 ;
        RECT 112.950 45.600 115.050 46.050 ;
        RECT 133.950 45.600 136.050 46.050 ;
        RECT 139.950 45.600 142.050 46.050 ;
        RECT 112.950 44.400 142.050 45.600 ;
        RECT 112.950 43.950 115.050 44.400 ;
        RECT 133.950 43.950 136.050 44.400 ;
        RECT 139.950 43.950 142.050 44.400 ;
        RECT 250.950 45.600 253.050 46.050 ;
        RECT 334.950 45.600 337.050 46.050 ;
        RECT 385.950 45.600 388.050 46.050 ;
        RECT 484.950 45.600 487.050 46.050 ;
        RECT 250.950 44.400 487.050 45.600 ;
        RECT 250.950 43.950 253.050 44.400 ;
        RECT 334.950 43.950 337.050 44.400 ;
        RECT 385.950 43.950 388.050 44.400 ;
        RECT 484.950 43.950 487.050 44.400 ;
        RECT 490.950 45.600 493.050 46.050 ;
        RECT 499.950 45.600 502.050 46.050 ;
        RECT 508.950 45.600 511.050 46.050 ;
        RECT 718.950 45.600 721.050 46.050 ;
        RECT 733.950 45.600 736.050 46.050 ;
        RECT 745.950 45.600 748.050 46.050 ;
        RECT 757.950 45.600 760.050 46.050 ;
        RECT 490.950 44.400 543.600 45.600 ;
        RECT 490.950 43.950 493.050 44.400 ;
        RECT 499.950 43.950 502.050 44.400 ;
        RECT 508.950 43.950 511.050 44.400 ;
        RECT 106.950 42.600 109.050 43.050 ;
        RECT 274.950 42.600 277.050 43.050 ;
        RECT 343.950 42.600 346.050 43.050 ;
        RECT 535.950 42.600 538.050 43.050 ;
        RECT 106.950 41.400 538.050 42.600 ;
        RECT 542.400 42.600 543.600 44.400 ;
        RECT 718.950 44.400 760.050 45.600 ;
        RECT 718.950 43.950 721.050 44.400 ;
        RECT 733.950 43.950 736.050 44.400 ;
        RECT 745.950 43.950 748.050 44.400 ;
        RECT 757.950 43.950 760.050 44.400 ;
        RECT 706.950 42.600 709.050 43.050 ;
        RECT 724.950 42.600 727.050 43.050 ;
        RECT 542.400 41.400 727.050 42.600 ;
        RECT 106.950 40.950 109.050 41.400 ;
        RECT 274.950 40.950 277.050 41.400 ;
        RECT 343.950 40.950 346.050 41.400 ;
        RECT 535.950 40.950 538.050 41.400 ;
        RECT 706.950 40.950 709.050 41.400 ;
        RECT 724.950 40.950 727.050 41.400 ;
        RECT 142.950 39.600 145.050 40.050 ;
        RECT 166.950 39.600 169.050 40.050 ;
        RECT 142.950 38.400 169.050 39.600 ;
        RECT 142.950 37.950 145.050 38.400 ;
        RECT 166.950 37.950 169.050 38.400 ;
        RECT 172.950 39.600 175.050 40.050 ;
        RECT 286.950 39.600 289.050 40.050 ;
        RECT 172.950 38.400 289.050 39.600 ;
        RECT 172.950 37.950 175.050 38.400 ;
        RECT 286.950 37.950 289.050 38.400 ;
        RECT 289.950 39.600 292.050 40.050 ;
        RECT 298.950 39.600 301.050 40.050 ;
        RECT 289.950 38.400 301.050 39.600 ;
        RECT 289.950 37.950 292.050 38.400 ;
        RECT 298.950 37.950 301.050 38.400 ;
        RECT 307.950 39.600 310.050 40.050 ;
        RECT 337.950 39.600 340.050 40.050 ;
        RECT 307.950 38.400 340.050 39.600 ;
        RECT 307.950 37.950 310.050 38.400 ;
        RECT 337.950 37.950 340.050 38.400 ;
        RECT 349.950 39.600 352.050 40.050 ;
        RECT 361.950 39.600 364.050 40.050 ;
        RECT 349.950 38.400 364.050 39.600 ;
        RECT 349.950 37.950 352.050 38.400 ;
        RECT 361.950 37.950 364.050 38.400 ;
        RECT 391.950 39.600 394.050 40.050 ;
        RECT 397.950 39.600 400.050 40.050 ;
        RECT 409.950 39.600 412.050 40.050 ;
        RECT 418.950 39.600 421.050 40.050 ;
        RECT 391.950 38.400 421.050 39.600 ;
        RECT 391.950 37.950 394.050 38.400 ;
        RECT 397.950 37.950 400.050 38.400 ;
        RECT 409.950 37.950 412.050 38.400 ;
        RECT 418.950 37.950 421.050 38.400 ;
        RECT 445.950 39.600 448.050 40.050 ;
        RECT 496.950 39.600 499.050 40.050 ;
        RECT 517.950 39.600 520.050 40.050 ;
        RECT 529.950 39.600 532.050 40.050 ;
        RECT 445.950 38.400 532.050 39.600 ;
        RECT 445.950 37.950 448.050 38.400 ;
        RECT 496.950 37.950 499.050 38.400 ;
        RECT 517.950 37.950 520.050 38.400 ;
        RECT 529.950 37.950 532.050 38.400 ;
        RECT 91.950 36.600 94.050 37.050 ;
        RECT 166.950 36.600 169.050 37.050 ;
        RECT 322.950 36.600 325.050 37.050 ;
        RECT 91.950 35.400 132.600 36.600 ;
        RECT 91.950 34.950 94.050 35.400 ;
        RECT 85.950 33.600 88.050 34.050 ;
        RECT 127.950 33.600 130.050 34.050 ;
        RECT 85.950 32.400 130.050 33.600 ;
        RECT 131.400 33.600 132.600 35.400 ;
        RECT 166.950 35.400 325.050 36.600 ;
        RECT 166.950 34.950 169.050 35.400 ;
        RECT 322.950 34.950 325.050 35.400 ;
        RECT 361.950 36.600 364.050 37.050 ;
        RECT 463.950 36.600 466.050 37.050 ;
        RECT 361.950 35.400 466.050 36.600 ;
        RECT 361.950 34.950 364.050 35.400 ;
        RECT 463.950 34.950 466.050 35.400 ;
        RECT 469.950 36.600 472.050 37.050 ;
        RECT 493.950 36.600 496.050 37.050 ;
        RECT 469.950 35.400 496.050 36.600 ;
        RECT 469.950 34.950 472.050 35.400 ;
        RECT 493.950 34.950 496.050 35.400 ;
        RECT 658.950 36.600 661.050 37.050 ;
        RECT 682.950 36.600 685.050 37.050 ;
        RECT 658.950 35.400 685.050 36.600 ;
        RECT 658.950 34.950 661.050 35.400 ;
        RECT 682.950 34.950 685.050 35.400 ;
        RECT 166.950 33.600 169.050 34.050 ;
        RECT 131.400 32.400 169.050 33.600 ;
        RECT 85.950 31.950 88.050 32.400 ;
        RECT 127.950 31.950 130.050 32.400 ;
        RECT 166.950 31.950 169.050 32.400 ;
        RECT 208.950 33.600 211.050 34.050 ;
        RECT 262.950 33.600 265.050 34.050 ;
        RECT 208.950 32.400 265.050 33.600 ;
        RECT 208.950 31.950 211.050 32.400 ;
        RECT 262.950 31.950 265.050 32.400 ;
        RECT 298.950 33.600 301.050 34.050 ;
        RECT 370.950 33.600 373.050 34.050 ;
        RECT 298.950 32.400 373.050 33.600 ;
        RECT 298.950 31.950 301.050 32.400 ;
        RECT 370.950 31.950 373.050 32.400 ;
        RECT 382.950 33.600 385.050 34.050 ;
        RECT 394.950 33.600 397.050 34.050 ;
        RECT 382.950 32.400 397.050 33.600 ;
        RECT 382.950 31.950 385.050 32.400 ;
        RECT 394.950 31.950 397.050 32.400 ;
        RECT 406.950 33.600 409.050 34.050 ;
        RECT 664.950 33.600 667.050 34.050 ;
        RECT 703.950 33.600 706.050 34.050 ;
        RECT 406.950 32.400 706.050 33.600 ;
        RECT 406.950 31.950 409.050 32.400 ;
        RECT 664.950 31.950 667.050 32.400 ;
        RECT 703.950 31.950 706.050 32.400 ;
        RECT 94.950 30.600 97.050 31.050 ;
        RECT 115.950 30.600 118.050 31.050 ;
        RECT 94.950 29.400 118.050 30.600 ;
        RECT 94.950 28.950 97.050 29.400 ;
        RECT 115.950 28.950 118.050 29.400 ;
        RECT 127.950 30.600 130.050 31.050 ;
        RECT 193.950 30.600 196.050 31.050 ;
        RECT 127.950 29.400 196.050 30.600 ;
        RECT 127.950 28.950 130.050 29.400 ;
        RECT 193.950 28.950 196.050 29.400 ;
        RECT 247.950 30.600 250.050 31.050 ;
        RECT 289.950 30.600 292.050 31.050 ;
        RECT 247.950 29.400 292.050 30.600 ;
        RECT 247.950 28.950 250.050 29.400 ;
        RECT 289.950 28.950 292.050 29.400 ;
        RECT 298.950 30.600 301.050 31.050 ;
        RECT 376.950 30.600 379.050 31.050 ;
        RECT 400.950 30.600 403.050 31.050 ;
        RECT 418.950 30.600 421.050 31.050 ;
        RECT 298.950 29.400 421.050 30.600 ;
        RECT 298.950 28.950 301.050 29.400 ;
        RECT 376.950 28.950 379.050 29.400 ;
        RECT 400.950 28.950 403.050 29.400 ;
        RECT 418.950 28.950 421.050 29.400 ;
        RECT 430.950 30.600 433.050 31.050 ;
        RECT 439.950 30.600 442.050 31.050 ;
        RECT 484.950 30.600 487.050 31.050 ;
        RECT 514.950 30.600 517.050 31.050 ;
        RECT 430.950 29.400 487.050 30.600 ;
        RECT 430.950 28.950 433.050 29.400 ;
        RECT 439.950 28.950 442.050 29.400 ;
        RECT 484.950 28.950 487.050 29.400 ;
        RECT 488.400 29.400 517.050 30.600 ;
        RECT 28.950 27.600 31.050 28.050 ;
        RECT 106.950 27.600 109.050 28.050 ;
        RECT 28.950 26.400 109.050 27.600 ;
        RECT 28.950 25.950 31.050 26.400 ;
        RECT 106.950 25.950 109.050 26.400 ;
        RECT 124.950 27.600 127.050 28.050 ;
        RECT 136.950 27.600 139.050 28.050 ;
        RECT 124.950 26.400 139.050 27.600 ;
        RECT 124.950 25.950 127.050 26.400 ;
        RECT 136.950 25.950 139.050 26.400 ;
        RECT 139.950 27.600 142.050 28.050 ;
        RECT 163.950 27.600 166.050 28.050 ;
        RECT 139.950 26.400 166.050 27.600 ;
        RECT 139.950 25.950 142.050 26.400 ;
        RECT 163.950 25.950 166.050 26.400 ;
        RECT 184.950 27.600 187.050 28.050 ;
        RECT 292.950 27.600 295.050 28.050 ;
        RECT 184.950 26.400 295.050 27.600 ;
        RECT 184.950 25.950 187.050 26.400 ;
        RECT 292.950 25.950 295.050 26.400 ;
        RECT 295.950 27.600 298.050 28.050 ;
        RECT 301.950 27.600 304.050 28.050 ;
        RECT 295.950 26.400 304.050 27.600 ;
        RECT 295.950 25.950 298.050 26.400 ;
        RECT 301.950 25.950 304.050 26.400 ;
        RECT 313.950 27.600 316.050 28.050 ;
        RECT 328.950 27.600 331.050 28.050 ;
        RECT 313.950 26.400 331.050 27.600 ;
        RECT 313.950 25.950 316.050 26.400 ;
        RECT 328.950 25.950 331.050 26.400 ;
        RECT 340.950 27.600 343.050 28.050 ;
        RECT 352.950 27.600 355.050 28.050 ;
        RECT 361.950 27.600 364.050 28.050 ;
        RECT 340.950 26.400 364.050 27.600 ;
        RECT 340.950 25.950 343.050 26.400 ;
        RECT 352.950 25.950 355.050 26.400 ;
        RECT 361.950 25.950 364.050 26.400 ;
        RECT 370.950 27.600 373.050 28.050 ;
        RECT 436.950 27.600 439.050 28.050 ;
        RECT 370.950 26.400 439.050 27.600 ;
        RECT 370.950 25.950 373.050 26.400 ;
        RECT 436.950 25.950 439.050 26.400 ;
        RECT 454.950 27.600 457.050 28.050 ;
        RECT 488.400 27.600 489.600 29.400 ;
        RECT 514.950 28.950 517.050 29.400 ;
        RECT 454.950 26.400 489.600 27.600 ;
        RECT 493.950 27.600 496.050 28.050 ;
        RECT 526.950 27.600 529.050 28.050 ;
        RECT 493.950 26.400 529.050 27.600 ;
        RECT 454.950 25.950 457.050 26.400 ;
        RECT 493.950 25.950 496.050 26.400 ;
        RECT 526.950 25.950 529.050 26.400 ;
        RECT 532.950 27.600 535.050 28.050 ;
        RECT 559.950 27.600 562.050 28.050 ;
        RECT 532.950 26.400 562.050 27.600 ;
        RECT 532.950 25.950 535.050 26.400 ;
        RECT 559.950 25.950 562.050 26.400 ;
        RECT 577.950 27.600 580.050 28.050 ;
        RECT 628.950 27.600 631.050 28.050 ;
        RECT 577.950 26.400 631.050 27.600 ;
        RECT 577.950 25.950 580.050 26.400 ;
        RECT 628.950 25.950 631.050 26.400 ;
        RECT 655.950 27.600 658.050 28.050 ;
        RECT 661.950 27.600 664.050 28.050 ;
        RECT 655.950 26.400 664.050 27.600 ;
        RECT 655.950 25.950 658.050 26.400 ;
        RECT 661.950 25.950 664.050 26.400 ;
        RECT 670.950 27.600 673.050 28.050 ;
        RECT 679.950 27.600 682.050 28.050 ;
        RECT 670.950 26.400 682.050 27.600 ;
        RECT 670.950 25.950 673.050 26.400 ;
        RECT 679.950 25.950 682.050 26.400 ;
        RECT 685.950 27.600 688.050 28.050 ;
        RECT 697.950 27.600 700.050 28.050 ;
        RECT 685.950 26.400 700.050 27.600 ;
        RECT 685.950 25.950 688.050 26.400 ;
        RECT 697.950 25.950 700.050 26.400 ;
        RECT 787.950 27.600 790.050 28.050 ;
        RECT 823.950 27.600 826.050 28.050 ;
        RECT 787.950 26.400 826.050 27.600 ;
        RECT 787.950 25.950 790.050 26.400 ;
        RECT 823.950 25.950 826.050 26.400 ;
        RECT 91.950 24.600 94.050 25.050 ;
        RECT 103.950 24.600 106.050 25.050 ;
        RECT 91.950 23.400 106.050 24.600 ;
        RECT 91.950 22.950 94.050 23.400 ;
        RECT 103.950 22.950 106.050 23.400 ;
        RECT 112.950 24.600 115.050 25.050 ;
        RECT 127.950 24.600 130.050 25.050 ;
        RECT 142.950 24.600 145.050 25.050 ;
        RECT 298.950 24.600 301.050 25.050 ;
        RECT 112.950 23.400 130.050 24.600 ;
        RECT 112.950 22.950 115.050 23.400 ;
        RECT 127.950 22.950 130.050 23.400 ;
        RECT 131.400 23.400 145.050 24.600 ;
        RECT 124.950 21.600 127.050 22.050 ;
        RECT 131.400 21.600 132.600 23.400 ;
        RECT 142.950 22.950 145.050 23.400 ;
        RECT 251.400 23.400 301.050 24.600 ;
        RECT 124.950 20.400 132.600 21.600 ;
        RECT 139.950 21.600 142.050 22.050 ;
        RECT 160.950 21.600 163.050 22.050 ;
        RECT 139.950 20.400 163.050 21.600 ;
        RECT 124.950 19.950 127.050 20.400 ;
        RECT 139.950 19.950 142.050 20.400 ;
        RECT 160.950 19.950 163.050 20.400 ;
        RECT 166.950 21.600 169.050 22.050 ;
        RECT 175.950 21.600 178.050 22.050 ;
        RECT 251.400 21.600 252.600 23.400 ;
        RECT 298.950 22.950 301.050 23.400 ;
        RECT 310.950 24.600 313.050 25.050 ;
        RECT 316.950 24.600 319.050 25.050 ;
        RECT 310.950 23.400 319.050 24.600 ;
        RECT 310.950 22.950 313.050 23.400 ;
        RECT 316.950 22.950 319.050 23.400 ;
        RECT 319.950 24.600 322.050 25.050 ;
        RECT 325.950 24.600 328.050 25.050 ;
        RECT 319.950 23.400 328.050 24.600 ;
        RECT 319.950 22.950 322.050 23.400 ;
        RECT 325.950 22.950 328.050 23.400 ;
        RECT 364.950 24.600 367.050 25.050 ;
        RECT 391.950 24.600 394.050 25.050 ;
        RECT 364.950 23.400 394.050 24.600 ;
        RECT 364.950 22.950 367.050 23.400 ;
        RECT 391.950 22.950 394.050 23.400 ;
        RECT 409.950 24.600 412.050 25.050 ;
        RECT 451.950 24.600 454.050 25.050 ;
        RECT 409.950 23.400 454.050 24.600 ;
        RECT 409.950 22.950 412.050 23.400 ;
        RECT 451.950 22.950 454.050 23.400 ;
        RECT 457.950 24.600 460.050 25.050 ;
        RECT 466.950 24.600 469.050 25.050 ;
        RECT 478.950 24.600 481.050 25.050 ;
        RECT 457.950 23.400 465.600 24.600 ;
        RECT 457.950 22.950 460.050 23.400 ;
        RECT 166.950 20.400 252.600 21.600 ;
        RECT 253.950 21.600 256.050 22.050 ;
        RECT 259.950 21.600 262.050 22.050 ;
        RECT 253.950 20.400 262.050 21.600 ;
        RECT 166.950 19.950 169.050 20.400 ;
        RECT 175.950 19.950 178.050 20.400 ;
        RECT 253.950 19.950 256.050 20.400 ;
        RECT 259.950 19.950 262.050 20.400 ;
        RECT 265.950 21.600 268.050 22.050 ;
        RECT 280.950 21.600 283.050 22.050 ;
        RECT 265.950 20.400 283.050 21.600 ;
        RECT 265.950 19.950 268.050 20.400 ;
        RECT 280.950 19.950 283.050 20.400 ;
        RECT 286.950 21.600 289.050 22.050 ;
        RECT 307.950 21.600 310.050 22.050 ;
        RECT 286.950 20.400 310.050 21.600 ;
        RECT 286.950 19.950 289.050 20.400 ;
        RECT 307.950 19.950 310.050 20.400 ;
        RECT 322.950 21.600 325.050 22.050 ;
        RECT 331.950 21.600 334.050 22.050 ;
        RECT 340.950 21.600 343.050 22.050 ;
        RECT 322.950 20.400 343.050 21.600 ;
        RECT 322.950 19.950 325.050 20.400 ;
        RECT 331.950 19.950 334.050 20.400 ;
        RECT 340.950 19.950 343.050 20.400 ;
        RECT 346.950 21.600 349.050 22.050 ;
        RECT 397.950 21.600 400.050 22.050 ;
        RECT 403.950 21.600 406.050 22.050 ;
        RECT 346.950 20.400 406.050 21.600 ;
        RECT 346.950 19.950 349.050 20.400 ;
        RECT 397.950 19.950 400.050 20.400 ;
        RECT 403.950 19.950 406.050 20.400 ;
        RECT 409.950 21.600 412.050 22.050 ;
        RECT 424.950 21.600 427.050 22.050 ;
        RECT 409.950 20.400 427.050 21.600 ;
        RECT 409.950 19.950 412.050 20.400 ;
        RECT 424.950 19.950 427.050 20.400 ;
        RECT 448.950 21.600 451.050 22.050 ;
        RECT 454.950 21.600 457.050 22.050 ;
        RECT 448.950 20.400 457.050 21.600 ;
        RECT 464.400 21.600 465.600 23.400 ;
        RECT 466.950 23.400 481.050 24.600 ;
        RECT 466.950 22.950 469.050 23.400 ;
        RECT 478.950 22.950 481.050 23.400 ;
        RECT 481.950 24.600 484.050 25.050 ;
        RECT 502.950 24.600 505.050 25.050 ;
        RECT 481.950 23.400 505.050 24.600 ;
        RECT 481.950 22.950 484.050 23.400 ;
        RECT 502.950 22.950 505.050 23.400 ;
        RECT 505.950 24.600 508.050 25.050 ;
        RECT 511.950 24.600 514.050 25.050 ;
        RECT 505.950 23.400 514.050 24.600 ;
        RECT 505.950 22.950 508.050 23.400 ;
        RECT 511.950 22.950 514.050 23.400 ;
        RECT 526.950 24.600 529.050 25.050 ;
        RECT 535.950 24.600 538.050 25.050 ;
        RECT 547.950 24.600 550.050 25.050 ;
        RECT 526.950 23.400 550.050 24.600 ;
        RECT 526.950 22.950 529.050 23.400 ;
        RECT 535.950 22.950 538.050 23.400 ;
        RECT 547.950 22.950 550.050 23.400 ;
        RECT 565.950 24.600 568.050 25.050 ;
        RECT 583.950 24.600 586.050 25.050 ;
        RECT 565.950 23.400 586.050 24.600 ;
        RECT 565.950 22.950 568.050 23.400 ;
        RECT 583.950 22.950 586.050 23.400 ;
        RECT 700.950 24.600 703.050 25.050 ;
        RECT 712.950 24.600 715.050 25.050 ;
        RECT 700.950 23.400 715.050 24.600 ;
        RECT 700.950 22.950 703.050 23.400 ;
        RECT 712.950 22.950 715.050 23.400 ;
        RECT 727.950 24.600 730.050 25.050 ;
        RECT 766.950 24.600 769.050 25.050 ;
        RECT 727.950 23.400 769.050 24.600 ;
        RECT 727.950 22.950 730.050 23.400 ;
        RECT 766.950 22.950 769.050 23.400 ;
        RECT 466.950 21.600 469.050 22.050 ;
        RECT 464.400 20.400 469.050 21.600 ;
        RECT 448.950 19.950 451.050 20.400 ;
        RECT 454.950 19.950 457.050 20.400 ;
        RECT 466.950 19.950 469.050 20.400 ;
        RECT 487.950 21.600 490.050 22.050 ;
        RECT 499.950 21.600 502.050 22.050 ;
        RECT 487.950 20.400 502.050 21.600 ;
        RECT 487.950 19.950 490.050 20.400 ;
        RECT 499.950 19.950 502.050 20.400 ;
        RECT 547.950 21.600 550.050 22.050 ;
        RECT 661.950 21.600 664.050 22.050 ;
        RECT 547.950 20.400 664.050 21.600 ;
        RECT 547.950 19.950 550.050 20.400 ;
        RECT 661.950 19.950 664.050 20.400 ;
        RECT 667.950 21.600 670.050 22.050 ;
        RECT 673.950 21.600 676.050 22.050 ;
        RECT 718.950 21.600 721.050 22.050 ;
        RECT 667.950 20.400 676.050 21.600 ;
        RECT 667.950 19.950 670.050 20.400 ;
        RECT 673.950 19.950 676.050 20.400 ;
        RECT 704.400 20.400 721.050 21.600 ;
        RECT 67.950 18.600 70.050 19.050 ;
        RECT 85.950 18.600 88.050 19.050 ;
        RECT 67.950 17.400 88.050 18.600 ;
        RECT 67.950 16.950 70.050 17.400 ;
        RECT 85.950 16.950 88.050 17.400 ;
        RECT 94.950 18.600 97.050 19.050 ;
        RECT 127.950 18.600 130.050 19.050 ;
        RECT 493.950 18.600 496.050 19.050 ;
        RECT 94.950 17.400 496.050 18.600 ;
        RECT 94.950 16.950 97.050 17.400 ;
        RECT 127.950 16.950 130.050 17.400 ;
        RECT 493.950 16.950 496.050 17.400 ;
        RECT 535.950 18.600 538.050 19.050 ;
        RECT 544.950 18.600 547.050 19.050 ;
        RECT 535.950 17.400 547.050 18.600 ;
        RECT 535.950 16.950 538.050 17.400 ;
        RECT 544.950 16.950 547.050 17.400 ;
        RECT 553.950 18.600 556.050 19.050 ;
        RECT 568.950 18.600 571.050 19.050 ;
        RECT 589.950 18.600 592.050 19.050 ;
        RECT 553.950 17.400 592.050 18.600 ;
        RECT 553.950 16.950 556.050 17.400 ;
        RECT 568.950 16.950 571.050 17.400 ;
        RECT 589.950 16.950 592.050 17.400 ;
        RECT 661.950 18.600 664.050 19.050 ;
        RECT 704.400 18.600 705.600 20.400 ;
        RECT 718.950 19.950 721.050 20.400 ;
        RECT 733.950 21.600 736.050 22.050 ;
        RECT 739.950 21.600 742.050 22.050 ;
        RECT 733.950 20.400 742.050 21.600 ;
        RECT 733.950 19.950 736.050 20.400 ;
        RECT 739.950 19.950 742.050 20.400 ;
        RECT 661.950 17.400 705.600 18.600 ;
        RECT 706.950 18.600 709.050 19.050 ;
        RECT 724.950 18.600 727.050 19.050 ;
        RECT 706.950 17.400 727.050 18.600 ;
        RECT 661.950 16.950 664.050 17.400 ;
        RECT 706.950 16.950 709.050 17.400 ;
        RECT 724.950 16.950 727.050 17.400 ;
        RECT 736.950 18.600 739.050 19.050 ;
        RECT 754.950 18.600 757.050 19.050 ;
        RECT 736.950 17.400 757.050 18.600 ;
        RECT 736.950 16.950 739.050 17.400 ;
        RECT 754.950 16.950 757.050 17.400 ;
        RECT 760.950 18.600 763.050 19.050 ;
        RECT 769.950 18.600 772.050 19.050 ;
        RECT 760.950 17.400 772.050 18.600 ;
        RECT 760.950 16.950 763.050 17.400 ;
        RECT 769.950 16.950 772.050 17.400 ;
        RECT 847.950 18.600 850.050 19.050 ;
        RECT 853.950 18.600 856.050 19.050 ;
        RECT 847.950 17.400 856.050 18.600 ;
        RECT 847.950 16.950 850.050 17.400 ;
        RECT 853.950 16.950 856.050 17.400 ;
        RECT 52.950 15.600 55.050 16.050 ;
        RECT 73.950 15.600 76.050 16.050 ;
        RECT 94.950 15.600 97.050 16.050 ;
        RECT 52.950 14.400 97.050 15.600 ;
        RECT 52.950 13.950 55.050 14.400 ;
        RECT 73.950 13.950 76.050 14.400 ;
        RECT 94.950 13.950 97.050 14.400 ;
        RECT 118.950 15.600 121.050 16.050 ;
        RECT 148.950 15.600 151.050 16.050 ;
        RECT 118.950 14.400 151.050 15.600 ;
        RECT 118.950 13.950 121.050 14.400 ;
        RECT 148.950 13.950 151.050 14.400 ;
        RECT 301.950 15.600 304.050 16.050 ;
        RECT 319.950 15.600 322.050 16.050 ;
        RECT 379.950 15.600 382.050 16.050 ;
        RECT 301.950 14.400 382.050 15.600 ;
        RECT 301.950 13.950 304.050 14.400 ;
        RECT 319.950 13.950 322.050 14.400 ;
        RECT 379.950 13.950 382.050 14.400 ;
        RECT 394.950 15.600 397.050 16.050 ;
        RECT 535.950 15.600 538.050 16.050 ;
        RECT 394.950 14.400 538.050 15.600 ;
        RECT 394.950 13.950 397.050 14.400 ;
        RECT 535.950 13.950 538.050 14.400 ;
        RECT 550.950 15.600 553.050 16.050 ;
        RECT 574.950 15.600 577.050 16.050 ;
        RECT 550.950 14.400 577.050 15.600 ;
        RECT 550.950 13.950 553.050 14.400 ;
        RECT 574.950 13.950 577.050 14.400 ;
        RECT 703.950 15.600 706.050 16.050 ;
        RECT 709.950 15.600 712.050 16.050 ;
        RECT 703.950 14.400 712.050 15.600 ;
        RECT 703.950 13.950 706.050 14.400 ;
        RECT 709.950 13.950 712.050 14.400 ;
        RECT 721.950 15.600 724.050 16.050 ;
        RECT 736.950 15.600 739.050 16.050 ;
        RECT 721.950 14.400 739.050 15.600 ;
        RECT 721.950 13.950 724.050 14.400 ;
        RECT 736.950 13.950 739.050 14.400 ;
        RECT 766.950 15.600 769.050 16.050 ;
        RECT 775.950 15.600 778.050 16.050 ;
        RECT 766.950 14.400 778.050 15.600 ;
        RECT 766.950 13.950 769.050 14.400 ;
        RECT 775.950 13.950 778.050 14.400 ;
        RECT 109.950 12.600 112.050 13.050 ;
        RECT 130.950 12.600 133.050 13.050 ;
        RECT 109.950 11.400 133.050 12.600 ;
        RECT 109.950 10.950 112.050 11.400 ;
        RECT 130.950 10.950 133.050 11.400 ;
        RECT 283.950 12.600 286.050 13.050 ;
        RECT 316.950 12.600 319.050 13.050 ;
        RECT 283.950 11.400 319.050 12.600 ;
        RECT 283.950 10.950 286.050 11.400 ;
        RECT 316.950 10.950 319.050 11.400 ;
        RECT 460.950 12.600 463.050 13.050 ;
        RECT 481.950 12.600 484.050 13.050 ;
        RECT 460.950 11.400 484.050 12.600 ;
        RECT 460.950 10.950 463.050 11.400 ;
        RECT 481.950 10.950 484.050 11.400 ;
        RECT 4.950 9.600 7.050 10.050 ;
        RECT 184.950 9.600 187.050 10.050 ;
        RECT 4.950 8.400 187.050 9.600 ;
        RECT 4.950 7.950 7.050 8.400 ;
        RECT 184.950 7.950 187.050 8.400 ;
        RECT 412.950 9.600 415.050 10.050 ;
        RECT 490.950 9.600 493.050 10.050 ;
        RECT 763.950 9.600 766.050 10.050 ;
        RECT 784.950 9.600 787.050 10.050 ;
        RECT 412.950 8.400 493.050 9.600 ;
        RECT 412.950 7.950 415.050 8.400 ;
        RECT 490.950 7.950 493.050 8.400 ;
        RECT 536.400 8.400 787.050 9.600 ;
        RECT 337.950 6.600 340.050 7.050 ;
        RECT 523.950 6.600 526.050 7.050 ;
        RECT 536.400 6.600 537.600 8.400 ;
        RECT 763.950 7.950 766.050 8.400 ;
        RECT 784.950 7.950 787.050 8.400 ;
        RECT 337.950 5.400 537.600 6.600 ;
        RECT 337.950 4.950 340.050 5.400 ;
        RECT 523.950 4.950 526.050 5.400 ;
  END
END pong_pt1
END LIBRARY

