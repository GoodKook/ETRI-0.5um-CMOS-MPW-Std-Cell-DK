magic
tech scmos
magscale 1 60
timestamp 1709422372
<< checkpaint >>
rect 147100 672200 952620 677000
rect 140100 605700 952620 672200
rect 140100 600900 663108 605700
rect 147040 596560 663108 600900
rect 141400 596320 663108 596560
rect 135220 585368 663108 596320
rect 128800 584900 663108 585368
rect 128800 573954 663400 584900
rect 674260 577720 726780 590260
rect 128800 561414 666414 573954
rect 128800 555112 663400 561414
rect 110500 462584 663400 555112
rect 110500 444584 767640 462584
rect 110500 404530 663400 444584
rect 110500 316292 672200 404530
rect 82768 315260 672200 316292
rect 59274 288860 672200 315260
rect 62160 288654 672200 288860
rect 75556 278350 672200 288654
rect 110500 238750 672200 278350
rect 124042 235112 672200 238750
rect 110500 206750 672200 235112
rect 124042 173948 672200 206750
rect 101586 147100 672200 173948
rect 101586 128800 553500 147100
rect 558558 146716 645594 147100
rect 558558 130540 611800 146716
rect 558558 130300 611500 130540
rect 558558 130000 610540 130300
rect 558558 128800 587340 130000
rect 101586 127840 552958 128800
rect 101586 126030 182410 127840
rect 110910 113416 182410 126030
rect 109300 109300 111702 111702
rect 204796 110500 232958 127840
rect 236796 110500 265158 127840
rect 268796 110500 297158 127840
rect 300796 110500 552958 127840
<< metal1 >>
rect 208600 557700 226300 559300
rect 208600 539260 210400 557700
rect 530700 556300 552580 558700
rect 550780 538060 552580 556300
rect 208500 379700 209300 381300
rect 208600 201900 210400 207100
rect 550780 202900 552580 207238
rect 208596 200900 226300 201900
rect 208596 200700 213100 200900
rect 213100 198882 226300 198900
rect 530700 200900 552580 202900
<< m2contact >>
rect 213100 559300 226300 561100
rect 530700 558700 548900 561100
rect 213100 198900 226300 200900
rect 530700 198700 548900 200900
<< metal2 >>
rect 240900 549100 241600 561100
rect 272900 550300 273600 561100
rect 304900 551500 305600 561100
rect 336900 552700 337600 561100
rect 368900 556900 369600 561100
rect 363300 556300 369600 556900
rect 336900 552100 356700 552700
rect 304900 550900 354700 551500
rect 272900 549700 352500 550300
rect 240900 548500 341700 549100
rect 201900 547300 274400 547900
rect 201900 529400 202500 547300
rect 198800 528700 202500 529400
rect 203100 546100 270700 546700
rect 203100 519000 203700 546100
rect 198800 518300 203700 519000
rect 204300 544900 263200 545500
rect 204300 465400 204900 544900
rect 198800 464700 204900 465400
rect 205500 543700 252700 544300
rect 205500 433400 206100 543700
rect 198800 432700 206100 433400
rect 206700 542500 222100 543100
rect 252100 542500 252700 543700
rect 262500 542600 263200 544900
rect 270100 542500 270700 546100
rect 206700 401500 207300 542500
rect 221500 542300 222100 542500
rect 273800 542400 274400 547300
rect 341000 542500 341700 548500
rect 351700 542500 352500 549700
rect 353900 542500 354700 550900
rect 355900 542500 356700 552100
rect 363300 542500 363900 556300
rect 400900 555700 401600 561100
rect 365700 555100 401600 555700
rect 365700 542500 366300 555100
rect 432900 554500 433600 561000
rect 370900 553900 433600 554500
rect 370900 542500 371500 553900
rect 464900 553300 465600 561100
rect 374030 552700 465600 553300
rect 374030 542498 374592 552700
rect 496900 552100 497600 561100
rect 379972 551500 497600 552100
rect 379978 542476 380578 551500
rect 381260 550312 560500 550900
rect 381260 550300 383992 550312
rect 385150 550300 560500 550312
rect 381266 542432 381866 550300
rect 385150 549656 559300 549700
rect 384196 549110 559300 549656
rect 384196 549100 387112 549110
rect 387918 549100 559300 549110
rect 384200 548600 384800 549100
rect 384200 548500 384788 548600
rect 384196 547900 384788 548500
rect 384200 547300 384788 547900
rect 384196 546700 384788 547300
rect 384200 546100 384788 546700
rect 384196 545500 384788 546100
rect 384200 544900 384788 545500
rect 384196 544300 384788 544900
rect 384200 543700 384788 544300
rect 384196 543100 384788 543700
rect 384200 542400 384788 543100
rect 387208 548500 387800 548528
rect 387208 547900 558100 548500
rect 387208 547450 387800 547900
rect 387208 542400 387776 547450
rect 389602 546700 556900 547300
rect 389602 546690 390200 546700
rect 389614 546322 390200 546690
rect 389614 542400 390196 546322
rect 392602 545500 555700 546100
rect 392602 545030 393200 545500
rect 392602 543868 393194 545030
rect 399194 544300 554500 544900
rect 392602 542802 393184 543868
rect 399200 543726 399800 544300
rect 399200 543700 399798 543726
rect 399194 543100 399798 543700
rect 402182 543100 553300 543700
rect 392602 542400 393194 542802
rect 399200 542600 399798 543100
rect 399200 542400 399800 542600
rect 402200 542400 402800 543100
rect 198800 400700 207300 401500
rect 204300 387500 208500 388300
rect 198800 368700 200100 369400
rect 198800 358300 200600 359000
rect 198800 326300 201700 327000
rect 198800 294300 200800 295000
rect 198800 262300 201100 263100
rect 198800 230300 201500 231000
rect 204304 202500 204896 387500
rect 205500 379700 208500 380500
rect 205500 203700 206100 379700
rect 206700 362900 208500 363700
rect 206700 204900 207300 362900
rect 552700 337600 553300 543100
rect 553900 369600 554500 544300
rect 555100 401600 555700 545500
rect 556300 455200 556900 546700
rect 557500 465600 558100 547900
rect 558700 497600 559300 549100
rect 559900 529600 560500 550300
rect 559900 528880 561100 529600
rect 558700 496900 561100 497600
rect 557500 464900 561100 465600
rect 556300 454500 561100 455200
rect 555100 400900 561100 401600
rect 553900 368900 561100 369600
rect 552700 336900 561100 337600
rect 558700 326500 561100 327200
rect 557500 272900 561100 273600
rect 556300 262500 561100 263200
rect 555100 230500 561100 231200
rect 206700 204300 359200 204900
rect 205500 203100 305600 203700
rect 204300 201900 273600 202500
rect 262500 198800 263200 200000
rect 272900 198800 273600 201900
rect 304900 198800 305600 203100
rect 358500 198800 359200 204300
rect 370300 201700 370900 204700
rect 368900 201100 370900 201700
rect 368900 198800 369600 201100
rect 417100 200500 417700 204900
rect 417100 199900 423200 200500
rect 422500 198800 423200 199900
rect 518500 198800 519300 204500
<< m3contact >>
rect 208500 387500 209300 389100
rect 200100 368700 200700 370100
rect 200600 358300 201900 359000
rect 201700 326300 203100 327000
rect 200800 294300 202400 295000
rect 201100 262300 202600 263100
rect 201500 230300 202900 231000
rect 208500 379700 209300 381300
rect 208500 362900 209300 364500
rect 558100 326500 558700 328000
rect 556900 272900 557500 274300
rect 555700 262500 556300 263900
rect 554500 230500 555100 231800
rect 262500 200000 263200 201200
rect 518500 204500 520000 205100
<< metal3 >>
rect 200100 538510 208900 538700
rect 200100 538270 210820 538510
rect 200100 538100 208900 538270
rect 200100 370100 200700 538100
rect 201300 484300 208700 484900
rect 201300 359000 201900 484300
rect 202500 482900 208700 483500
rect 202500 327000 203100 482900
rect 203700 466700 208900 467300
rect 203700 295000 204300 466700
rect 202400 294300 204300 295000
rect 204900 443300 208700 443900
rect 204900 263100 205500 443300
rect 202600 262300 205500 263100
rect 206100 421500 208700 422300
rect 206100 231000 206700 421500
rect 202900 230300 206700 231000
rect 207300 419700 208700 420500
rect 552300 419700 558700 420500
rect 207300 203100 207900 419700
rect 552300 411900 557500 412700
rect 552300 404100 556300 404900
rect 552300 387300 555100 388100
rect 552300 357900 553900 358700
rect 553300 205100 553900 357900
rect 554500 231800 555100 387300
rect 555700 263900 556300 404100
rect 556900 274300 557500 411900
rect 558100 328000 558700 419700
rect 520000 204500 553900 205100
rect 207300 202500 263200 203100
rect 262500 201200 263200 202500
<< comment >>
rect 0 0 760000 760000
use POB8  AB[0] ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/chip_top/pads_ETRI050
timestamp 1537935238
transform 0 -1 611610 1 0 271950
box -200 -18300 24200 50600
use POB8  AB[1]
timestamp 1537935238
transform 1 0 271958 0 -1 611560
box -200 -18300 24200 50600
use POB8  AB[2]
timestamp 1537935238
transform 1 0 303958 0 -1 611560
box -200 -18300 24200 50600
use POB8  AB[3]
timestamp 1537935238
transform 1 0 463958 0 -1 611560
box -200 -18300 24200 50600
use POB8  AB[4]
timestamp 1537935238
transform 1 0 239958 0 -1 611560
box -200 -18300 24200 50600
use POB8  AB[5]
timestamp 1537935238
transform 1 0 399958 0 -1 611560
box -200 -18300 24200 50600
use POB8  AB[6]
timestamp 1537935238
transform 1 0 495958 0 -1 611560
box -200 -18300 24200 50600
use POB8  AB[7]
timestamp 1537935238
transform 1 0 431958 0 -1 611560
box -200 -18300 24200 50600
use POB8  AB[8]
timestamp 1537935238
transform 1 0 303958 0 1 148300
box -200 -18300 24200 50600
use POB8  AB[9]
timestamp 1537935238
transform 0 1 148300 -1 0 231950
box -200 -18300 24200 50600
use POB8  AB[10]
timestamp 1537935238
transform 1 0 271958 0 1 148300
box -200 -18300 24200 50600
use POB8  AB[11]
timestamp 1537935238
transform 0 1 148300 -1 0 263950
box -200 -18300 24200 50600
use POB8  AB[12]
timestamp 1537935238
transform 0 1 148300 -1 0 295950
box -200 -18300 24200 50600
use POB8  AB[13]
timestamp 1537935238
transform 0 1 148300 -1 0 327950
box -200 -18300 24200 50600
use POB8  AB[14]
timestamp 1537935238
transform 0 1 148300 -1 0 519950
box -200 -18300 24200 50600
use POB8  AB[15]
timestamp 1537935238
transform 0 1 148300 -1 0 359950
box -200 -18300 24200 50600
use PIC  CLK ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/chip_top/pads_ETRI050
timestamp 1537935238
transform 0 -1 611610 1 0 303950
box -200 -18300 24200 50600
use cpu6502_Core  cpu6502_Core_0
timestamp 1709127331
transform 1 0 210490 0 1 205360
box -1890 -720 342090 337290
use PIC  DI[0]
timestamp 1537935238
transform 1 0 399958 0 1 148300
box -200 -18300 24200 50600
use PIC  DI[1]
timestamp 1537935238
transform 0 -1 611610 1 0 431950
box -200 -18300 24200 50600
use PIC  DI[2]
timestamp 1537935238
transform 1 0 335958 0 1 148300
box -200 -18300 24200 50600
use PIC  DI[3]
timestamp 1537935238
transform 0 1 148300 -1 0 423950
box -200 -18300 24200 50600
use PIC  DI[4]
timestamp 1537935238
transform 1 0 239958 0 1 148300
box -200 -18300 24200 50600
use PIC  DI[5]
timestamp 1537935238
transform 0 1 148300 -1 0 455950
box -200 -18300 24200 50600
use PIC  DI[6]
timestamp 1537935238
transform 0 1 148300 -1 0 487950
box -200 -18300 24200 50600
use PIC  DI[7]
timestamp 1537935238
transform 0 1 148300 -1 0 551950
box -200 -18300 24200 50600
use POB8  DO[0]
timestamp 1537935238
transform 1 0 367958 0 -1 611560
box -200 -18300 24200 50600
use POB8  DO[1]
timestamp 1537935238
transform 0 -1 611610 1 0 335950
box -200 -18300 24200 50600
use POB8  DO[2]
timestamp 1537935238
transform 0 -1 611610 1 0 495950
box -200 -18300 24200 50600
use POB8  DO[3]
timestamp 1537935238
transform 0 -1 611610 1 0 367950
box -200 -18300 24200 50600
use POB8  DO[4]
timestamp 1537935238
transform 1 0 335958 0 -1 611560
box -200 -18300 24200 50600
use POB8  DO[5]
timestamp 1537935238
transform 0 -1 611610 1 0 527950
box -200 -18300 24200 50600
use POB8  DO[6]
timestamp 1537935238
transform 0 -1 611610 1 0 399950
box -200 -18300 24200 50600
use POB8  DO[7]
timestamp 1537935238
transform 0 -1 611610 1 0 463950
box -200 -18300 24200 50600
use IOFILLER10  IOFILLER10_0 ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/chip_top/pads_ETRI050
timestamp 1537935238
transform 1 0 444678 0 1 148301
box -70 0 2070 50120
use IOFILLER10  IOFILLER10_1
timestamp 1537935238
transform 1 0 473438 0 1 148301
box -70 0 2070 50120
use IOFILLER10  IOFILLER10_2
timestamp 1537935238
transform 1 0 443038 0 1 148301
box -70 0 2070 50120
use IOFILLER10  IOFILLER10_3
timestamp 1537935238
transform 1 0 441438 0 1 148301
box -70 0 2070 50120
use IOFILLER10  IOFILLER10_4
timestamp 1537935238
transform 1 0 476678 0 1 148301
box -70 0 2070 50120
use IOFILLER10  IOFILLER10_5
timestamp 1537935238
transform 1 0 475038 0 1 148301
box -70 0 2070 50120
use IOFILLER40  IOFILLER40_0 ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/chip_top/pads_ETRI050
timestamp 1709340318
transform 1 0 263648 0 1 148300
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_1
timestamp 1709340318
transform 1 0 231648 0 1 148300
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_2
timestamp 1709340318
transform 1 0 327648 0 1 148300
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_3
timestamp 1709340318
transform 1 0 295648 0 1 148300
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_4
timestamp 1709340318
transform 1 0 391648 0 1 148300
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_5
timestamp 1709340318
transform 1 0 359648 0 1 148300
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_6
timestamp 1709340318
transform 1 0 455648 0 1 148300
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_7
timestamp 1709340318
transform 1 0 423648 0 1 148300
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_8
timestamp 1709340318
transform 1 0 519648 0 1 148300
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_9
timestamp 1709340318
transform 1 0 487648 0 1 148300
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_11
timestamp 1709340318
transform 1 0 263648 0 -1 611560
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_12
timestamp 1709340318
transform 1 0 231648 0 -1 611560
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_13
timestamp 1709340318
transform 1 0 327648 0 -1 611560
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_14
timestamp 1709340318
transform 1 0 295648 0 -1 611560
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_15
timestamp 1709340318
transform 1 0 391648 0 -1 611560
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_16
timestamp 1709340318
transform 1 0 359648 0 -1 611560
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_17
timestamp 1709340318
transform 1 0 455648 0 -1 611560
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_18
timestamp 1709340318
transform 1 0 423648 0 -1 611560
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_19
timestamp 1709340318
transform 1 0 519648 0 -1 611560
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_20
timestamp 1709340318
transform 1 0 487648 0 -1 611560
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_22
timestamp 1709340318
transform 0 1 148300 -1 0 304380
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_23
timestamp 1709340318
transform 0 1 148300 -1 0 240380
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_24
timestamp 1709340318
transform 0 1 148300 -1 0 272380
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_25
timestamp 1709340318
transform 0 1 148300 -1 0 400380
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_26
timestamp 1709340318
transform 0 1 148300 -1 0 336380
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_27
timestamp 1709340318
transform 0 1 148300 -1 0 368380
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_28
timestamp 1709340318
transform 0 1 148300 -1 0 464380
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_29
timestamp 1709340318
transform 0 1 148300 -1 0 432380
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_31
timestamp 1709340318
transform 0 1 148300 -1 0 496380
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_32
timestamp 1709340318
transform 0 1 148300 -1 0 528380
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_33
timestamp 1709340318
transform 0 -1 611610 1 0 295640
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_34
timestamp 1709340318
transform 0 -1 611610 1 0 231640
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_35
timestamp 1709340318
transform 0 -1 611610 1 0 263640
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_36
timestamp 1709340318
transform 0 -1 611610 1 0 391640
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_37
timestamp 1709340318
transform 0 -1 611610 1 0 327640
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_38
timestamp 1709340318
transform 0 -1 611610 1 0 359640
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_39
timestamp 1709340318
transform 0 -1 611610 1 0 455640
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_40
timestamp 1709340318
transform 0 -1 611610 1 0 423640
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_42
timestamp 1709340318
transform 0 -1 611610 1 0 487640
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_43
timestamp 1709340318
transform 0 -1 611610 1 0 519640
box 0 0 8720 50120
use IOFILLER50  IOFILLER50_0 ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/chip_top/pads_ETRI050
timestamp 1537935238
transform 1 0 198120 0 1 148300
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_1
timestamp 1537935238
transform 1 0 551650 0 1 148300
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_2
timestamp 1537935238
transform 1 0 551650 0 -1 611560
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_3
timestamp 1537935238
transform 1 0 198128 0 -1 611560
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_4
timestamp 1537935238
transform 0 1 148300 -1 0 208260
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_5
timestamp 1537935238
transform 0 1 148300 -1 0 561780
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_6
timestamp 1537935238
transform 0 -1 611610 -1 0 208260
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_7
timestamp 1537935238
transform 0 -1 611608 -1 0 561832
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_8
timestamp 1537935238
transform 1 0 463818 0 1 148301
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_9
timestamp 1537935238
transform 1 0 446198 0 1 148300
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_10
timestamp 1537935238
transform 1 0 431818 0 1 148301
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_11
timestamp 1537935238
transform 1 0 478198 0 1 148300
box -70 0 10070 50120
use PIC  IRQ
timestamp 1537935238
transform 0 -1 611610 1 0 207950
box -200 -18300 24200 50600
use MY_LOGO  MY_LOGO_0
timestamp 1706263538
transform 1 0 555820 0 1 131500
box 14100 240 54780 15240
use PIC  NMI
timestamp 1537935238
transform 1 0 495958 0 1 148300
box -200 -18300 24200 50600
use PAD80  PAD80_0 ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/chip_top/pads_ETRI050
timestamp 1709379016
transform 1 0 467458 0 1 130000
box 0 0 17000 17000
use PAD80  PAD80_1
timestamp 1709379016
transform 1 0 435458 0 1 130000
box 0 0 17000 17000
use PCORNER  PCORNER_0 ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/chip_top/pads_ETRI050
timestamp 1537935238
transform 1 0 148300 0 1 148300
box 0 0 50600 50600
use PCORNER  PCORNER_1
timestamp 1537935238
transform 1 0 148302 0 -1 611560
box 0 0 50600 50600
use PCORNER  PCORNER_2
timestamp 1537935238
transform 0 -1 611610 1 0 148300
box 0 0 50600 50600
use PCORNER  PCORNER_3
timestamp 1537935238
transform -1 0 611608 0 -1 611560
box 0 0 50600 50600
use PVDD  PVDD_0 ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/chip_top/pads_ETRI050
timestamp 1537935238
transform 1 0 207958 0 -1 611560
box 0 -18300 24000 50600
use PVDD  PVDD_1
timestamp 1537935238
transform 1 0 207758 0 1 148300
box 0 -18300 24000 50600
use PVSS  PVSS_0 ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/chip_top/pads_ETRI050
timestamp 1537935238
transform 1 0 527958 0 -1 611560
box 0 -18300 24000 50600
use PVSS  PVSS_1
timestamp 1537935238
transform 1 0 527958 0 1 148300
box 0 -18300 24000 50600
use PIC  RDY
timestamp 1537935238
transform 0 1 148300 -1 0 391950
box -200 -18300 24200 50600
use PIC  RESET
timestamp 1537935238
transform 0 -1 611610 1 0 239950
box -200 -18300 24200 50600
use POB8  WE
timestamp 1537935238
transform 1 0 367958 0 1 148300
box -200 -18300 24200 50600
<< end >>
