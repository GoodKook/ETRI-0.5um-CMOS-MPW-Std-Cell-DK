/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */

module fir8(
    inout vdd,
    inout gnd,
    input [7:0] Xin,
    output [7:0] Xout,
    input [15:0] Yin,
    output [15:0] Yout,
    input clk
);

wire _4972_ ;
wire _4552_ ;
wire _4132_ ;
wire _5757_ ;
wire _5337_ ;
wire _1677_ ;
wire _1257_ ;
wire _5090_ ;
wire _588_ ;
wire _168_ ;
wire _3823_ ;
wire _3403_ ;
wire _6295_ ;
wire _4608_ ;
wire [15:0] _4781_ ;
wire _4361_ ;
wire _800_ ;
wire _5986_ ;
wire _5566_ ;
wire _5146_ ;
wire _60_ ;
wire _1486_ ;
wire _1066_ ;
wire _397_ ;
wire _3632_ ;
wire _3212_ ;
wire _4837_ ;
wire _4417_ ;
wire _4590_ ;
wire _4170_ ;
wire _2903_ ;
wire _5795_ ;
wire _5375_ ;
wire [15:0] \u_fir_pe2.mul  ;
wire _1295_ ;
wire _3861_ ;
wire _3441_ ;
wire _3021_ ;
wire _4646_ ;
wire _4226_ ;
wire _2712_ ;
wire _5184_ ;
wire \X[1]_5_bF$buf0  ;
wire _3917_ ;
wire _3670_ ;
wire _3250_ ;
wire _4875_ ;
wire _4455_ ;
wire _4035_ ;
wire _2941_ ;
wire _2521_ ;
wire _2101_ ;
wire _3726_ ;
wire _3306_ ;
wire _6198_ ;
wire _4684_ ;
wire _4264_ ;
wire _703_ ;
wire _5889_ ;
wire _5469_ ;
wire _5049_ ;
wire _1389_ ;
wire _2750_ ;
wire _2330_ ;
wire _3955_ ;
wire _3535_ ;
wire _3115_ ;
wire _19_ ;
wire _1601_ ;
wire _4493_ ;
wire _4073_ ;
wire _932_ ;
wire _512_ ;
wire _2806_ ;
wire _5698_ ;
wire _5278_ ;
wire _1198_ ;
wire _3764_ ;
wire _3344_ ;
wire _4969_ ;
wire _4549_ ;
wire _4129_ ;
wire _5910_ ;
wire _1830_ ;
wire _1410_ ;
wire _741_ ;
wire _321_ ;
wire _2615_ ;
wire _5087_ ;
wire [15:0] \u_fir_pe4.mul  ;
wire _3993_ ;
wire _3573_ ;
wire _3153_ ;
wire [15:0] _4778_ ;
wire _4358_ ;
wire _57_ ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _2844_ ;
wire _2424_ ;
wire _2004_ ;
wire _3629_ ;
wire _3209_ ;
wire _3382_ ;
wire _4587_ ;
wire _4167_ ;
wire _606_ ;
wire _6313_ ;
wire _2653_ ;
wire _2233_ ;
wire _3858_ ;
wire _3438_ ;
wire _3018_ ;
wire _3191_ ;
wire _1924_ ;
wire _1504_ ;
wire _4396_ ;
wire _835_ ;
wire _415_ ;
wire _2709_ ;
wire _95_ ;
wire _6122_ ;
wire _2882_ ;
wire _2462_ ;
wire _2042_ ;
wire _3667_ ;
wire _3247_ ;
wire _5813_ ;
wire _1733_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _2938_ ;
wire _2518_ ;
wire _6351_ ;
wire _2691_ ;
wire _2271_ ;
wire _3896_ ;
wire _3476_ ;
wire _3056_ ;
wire _5622_ ;
wire _5202_ ;
wire _1962_ ;
wire _1542_ ;
wire _1122_ ;
wire _873_ ;
wire _453_ ;
wire _2747_ ;
wire _2327_ ;
wire _6160_ ;
wire [15:0] \u_fir_pe6.mul  ;
wire _2080_ ;
wire _3285_ ;
wire _5851_ ;
wire _5431_ ;
wire _5011_ ;
wire _929_ ;
wire _509_ ;
wire _6216_ ;
wire _1771_ ;
wire _1351_ ;
wire _682_ ;
wire _262_ ;
wire _2976_ ;
wire _2556_ ;
wire _2136_ ;
wire _4702_ ;
wire _5907_ ;
wire _3094_ ;
wire _1827_ ;
wire _1407_ ;
wire _4299_ ;
wire _5660_ ;
wire _5240_ ;
wire _738_ ;
wire _318_ ;
wire _6025_ ;
wire _1580_ ;
wire _1160_ ;
wire _491_ ;
wire _2785_ ;
wire _2365_ ;
wire _4931_ ;
wire _4511_ ;
wire _5716_ ;
wire _1636_ ;
wire _1216_ ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _6254_ ;
wire _2594_ ;
wire _2174_ ;
wire _3799_ ;
wire _3379_ ;
wire _4740_ ;
wire _4320_ ;
wire _5945_ ;
wire _5525_ ;
wire _5105_ ;
wire _1865_ ;
wire _1445_ ;
wire _1025_ ;
wire _776_ ;
wire _356_ ;
wire _6063_ ;
wire _3188_ ;
wire _5754_ ;
wire _5334_ ;
wire _6119_ ;
wire _1674_ ;
wire _1254_ ;
wire _585_ ;
wire _165_ ;
wire _2879_ ;
wire _2459_ ;
wire _2039_ ;
wire _3820_ ;
wire _3400_ ;
wire _6292_ ;
wire _4605_ ;
wire [15:0] \Y[4]  ;
wire _5983_ ;
wire _5563_ ;
wire _5143_ ;
wire _6348_ ;
wire _1483_ ;
wire _1063_ ;
wire _394_ ;
wire _2688_ ;
wire _2268_ ;
wire _4834_ ;
wire _4414_ ;
wire _5619_ ;
wire _1959_ ;
wire _1539_ ;
wire _1119_ ;
wire _2900_ ;
wire _5792_ ;
wire _5372_ ;
wire _6157_ ;
wire _1292_ ;
wire _2497_ ;
wire _2077_ ;
wire _4643_ ;
wire _4223_ ;
wire _5848_ ;
wire _5428_ ;
wire _5008_ ;
wire _1768_ ;
wire _1348_ ;
wire _5181_ ;
wire _679_ ;
wire _259_ ;
wire _3914_ ;
wire _4872_ ;
wire _4452_ ;
wire _4032_ ;
wire _5657_ ;
wire _5237_ ;
wire _1997_ ;
wire _1577_ ;
wire _1157_ ;
wire _488_ ;
wire _3723_ ;
wire _3303_ ;
wire _6195_ ;
wire _4928_ ;
wire _4508_ ;
wire _4681_ ;
wire _4261_ ;
wire _700_ ;
wire _5886_ ;
wire _5466_ ;
wire _5046_ ;
wire _1386_ ;
wire _297_ ;
wire _3952_ ;
wire _3532_ ;
wire _3112_ ;
wire _4737_ ;
wire _4317_ ;
wire _16_ ;
wire _4490_ ;
wire _4070_ ;
wire _2803_ ;
wire _5695_ ;
wire _5275_ ;
wire _1195_ ;
wire _3761_ ;
wire _3341_ ;
wire _4966_ ;
wire _4546_ ;
wire _4126_ ;
wire _2612_ ;
wire _5084_ ;
wire _3817_ ;
wire _6289_ ;
wire _3990_ ;
wire _3570_ ;
wire _3150_ ;
wire [15:0] _4775_ ;
wire _4355_ ;
wire _54_ ;
wire _2841_ ;
wire _2421_ ;
wire _2001_ ;
wire _3626_ ;
wire _3206_ ;
wire _6098_ ;
wire _4584_ ;
wire _4164_ ;
wire _603_ ;
wire _5789_ ;
wire _5369_ ;
wire _6310_ ;
wire _1289_ ;
wire _2650_ ;
wire _2230_ ;
wire _3855_ ;
wire _3435_ ;
wire _3015_ ;
wire _1921_ ;
wire _1501_ ;
wire _4393_ ;
wire _832_ ;
wire _412_ ;
wire _2706_ ;
wire _5598_ ;
wire _5178_ ;
wire _92_ ;
wire _1098_ ;
wire _3664_ ;
wire _3244_ ;
wire _4869_ ;
wire _4449_ ;
wire _4029_ ;
wire _5810_ ;
wire _1730_ ;
wire _1310_ ;
wire _641_ ;
wire _221_ ;
wire _2935_ ;
wire _2515_ ;
wire _3893_ ;
wire _3473_ ;
wire _3053_ ;
wire _4678_ ;
wire _4258_ ;
wire _870_ ;
wire _450_ ;
wire _2744_ ;
wire _2324_ ;
wire _3949_ ;
wire _3529_ ;
wire _3109_ ;
wire _3282_ ;
wire _4487_ ;
wire _4067_ ;
wire _926_ ;
wire _506_ ;
wire _6213_ ;
wire _2973_ ;
wire _2553_ ;
wire _2133_ ;
wire _3758_ ;
wire _3338_ ;
wire _5904_ ;
wire _3091_ ;
wire _1824_ ;
wire _1404_ ;
wire _4296_ ;
wire _735_ ;
wire _315_ ;
wire _2609_ ;
wire _6022_ ;
wire _2782_ ;
wire _2362_ ;
wire _3987_ ;
wire _3567_ ;
wire _3147_ ;
wire _5713_ ;
wire _1633_ ;
wire _1213_ ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire _2838_ ;
wire _2418_ ;
wire _6251_ ;
wire _2591_ ;
wire _2171_ ;
wire _3796_ ;
wire _3376_ ;
wire _5942_ ;
wire _5522_ ;
wire _5102_ ;
wire \X[6]_5_bF$buf1  ;
wire _6307_ ;
wire _1862_ ;
wire _1442_ ;
wire _1022_ ;
wire [15:0] \u_fir_pe4.rYin  ;
wire _773_ ;
wire _353_ ;
wire _2647_ ;
wire _2227_ ;
wire _6060_ ;
wire [15:0] _3185_ ;
wire _1918_ ;
wire _5751_ ;
wire _5331_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _6116_ ;
wire _1671_ ;
wire _1251_ ;
wire _582_ ;
wire _162_ ;
wire _2876_ ;
wire _2456_ ;
wire _2036_ ;
wire _4602_ ;
wire _5807_ ;
wire _1727_ ;
wire _1307_ ;
wire _4199_ ;
wire _5980_ ;
wire _5560_ ;
wire _5140_ ;
wire _638_ ;
wire _218_ ;
wire _6345_ ;
wire _1480_ ;
wire _1060_ ;
wire _391_ ;
wire _2685_ ;
wire _2265_ ;
wire _4831_ ;
wire _4411_ ;
wire _5616_ ;
wire _1956_ ;
wire _1536_ ;
wire _1116_ ;
wire _867_ ;
wire _447_ ;
wire _6154_ ;
wire _2494_ ;
wire _2074_ ;
wire _3699_ ;
wire _3279_ ;
wire _4640_ ;
wire _4220_ ;
wire _5845_ ;
wire _5425_ ;
wire _5005_ ;
wire _1765_ ;
wire _1345_ ;
wire _676_ ;
wire _256_ ;
wire _3911_ ;
wire _3088_ ;
wire _5654_ ;
wire _5234_ ;
wire _6019_ ;
wire _1994_ ;
wire _1574_ ;
wire _1154_ ;
wire _485_ ;
wire _2779_ ;
wire _2359_ ;
wire _3720_ ;
wire _3300_ ;
wire _6192_ ;
wire _4925_ ;
wire _4505_ ;
wire _5883_ ;
wire _5463_ ;
wire _5043_ ;
wire _6248_ ;
wire _1383_ ;
wire _294_ ;
wire _2588_ ;
wire _2168_ ;
wire _4734_ ;
wire _4314_ ;
wire _5939_ ;
wire _5519_ ;
wire _13_ ;
wire _1859_ ;
wire _1439_ ;
wire _1019_ ;
wire _2800_ ;
wire _5692_ ;
wire _5272_ ;
wire _6057_ ;
wire _1192_ ;
wire [7:0] \X[2]  ;
wire _2397_ ;
wire _4963_ ;
wire _4543_ ;
wire _4123_ ;
wire _5748_ ;
wire _5328_ ;
wire _1668_ ;
wire _1248_ ;
wire _5081_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire _3814_ ;
wire _6286_ ;
wire _4772_ ;
wire _4352_ ;
wire _5977_ ;
wire _5557_ ;
wire _5137_ ;
wire _51_ ;
wire _1897_ ;
wire _1477_ ;
wire _1057_ ;
wire _388_ ;
wire _3623_ ;
wire _3203_ ;
wire _6095_ ;
wire _4828_ ;
wire _4408_ ;
wire _4581_ ;
wire _4161_ ;
wire _600_ ;
wire _5786_ ;
wire _5366_ ;
wire _1286_ ;
wire _197_ ;
wire _3852_ ;
wire _3432_ ;
wire _3012_ ;
wire _4637_ ;
wire _4217_ ;
wire _4390_ ;
wire _2703_ ;
wire _5595_ ;
wire _5175_ ;
wire _3908_ ;
wire _1095_ ;
wire _3661_ ;
wire _3241_ ;
wire _4866_ ;
wire _4446_ ;
wire _4026_ ;
wire _2932_ ;
wire _2512_ ;
wire _3717_ ;
wire _6189_ ;
wire _3890_ ;
wire _3470_ ;
wire _3050_ ;
wire _4675_ ;
wire _4255_ ;
wire _2741_ ;
wire _2321_ ;
wire _3946_ ;
wire _3526_ ;
wire _3106_ ;
wire _7_ ;
wire _4484_ ;
wire _4064_ ;
wire _923_ ;
wire _503_ ;
wire _5689_ ;
wire _5269_ ;
wire _6210_ ;
wire _1189_ ;
wire _2970_ ;
wire _2550_ ;
wire _2130_ ;
wire _3755_ ;
wire _3335_ ;
wire _5901_ ;
wire _1821_ ;
wire _1401_ ;
wire _4293_ ;
wire _732_ ;
wire _312_ ;
wire _2606_ ;
wire _5498_ ;
wire _5078_ ;
wire [15:0] _3984_ ;
wire _3564_ ;
wire _3144_ ;
wire _4769_ ;
wire _4349_ ;
wire _5710_ ;
wire _48_ ;
wire _1630_ ;
wire _1210_ ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _2835_ ;
wire _2415_ ;
wire _3793_ ;
wire _3373_ ;
wire _4998_ ;
wire _4578_ ;
wire _4158_ ;
wire \X[5]_5_bF$buf3  ;
wire _6304_ ;
wire _770_ ;
wire _350_ ;
wire _2644_ ;
wire _2224_ ;
wire _3849_ ;
wire _3429_ ;
wire _3009_ ;
wire [15:0] _3182_ ;
wire _1915_ ;
wire _4387_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _6113_ ;
wire _2873_ ;
wire _2453_ ;
wire _2033_ ;
wire _3658_ ;
wire _3238_ ;
wire _5804_ ;
wire _1724_ ;
wire _1304_ ;
wire _4196_ ;
wire _635_ ;
wire _215_ ;
wire _2929_ ;
wire _2509_ ;
wire _6342_ ;
wire _2682_ ;
wire _2262_ ;
wire _3887_ ;
wire _3467_ ;
wire _3047_ ;
wire _5613_ ;
wire _1953_ ;
wire _1533_ ;
wire _1113_ ;
wire _864_ ;
wire _444_ ;
wire _2738_ ;
wire _2318_ ;
wire _6151_ ;
wire _2491_ ;
wire _2071_ ;
wire _3696_ ;
wire _3276_ ;
wire _5842_ ;
wire _5422_ ;
wire _5002_ ;
wire _6207_ ;
wire _1762_ ;
wire _1342_ ;
wire _673_ ;
wire _253_ ;
wire _2967_ ;
wire _2547_ ;
wire _2127_ ;
wire _3085_ ;
wire _1818_ ;
wire _5651_ ;
wire _5231_ ;
wire _729_ ;
wire _309_ ;
wire _6016_ ;
wire _1991_ ;
wire _1571_ ;
wire _1151_ ;
wire _482_ ;
wire _2776_ ;
wire _2356_ ;
wire _4922_ ;
wire _4502_ ;
wire _5707_ ;
wire _1627_ ;
wire _1207_ ;
wire _4099_ ;
wire _5880_ ;
wire _5460_ ;
wire _5040_ ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _6245_ ;
wire _1380_ ;
wire _291_ ;
wire _2585_ ;
wire _2165_ ;
wire _4731_ ;
wire _4311_ ;
wire _5936_ ;
wire _5516_ ;
wire _10_ ;
wire _1856_ ;
wire _1436_ ;
wire _1016_ ;
wire _767_ ;
wire _347_ ;
wire _6054_ ;
wire _2394_ ;
wire _3599_ ;
wire _3179_ ;
wire _4960_ ;
wire _4540_ ;
wire _4120_ ;
wire _5745_ ;
wire _5325_ ;
wire _1665_ ;
wire _1245_ ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire _3811_ ;
wire _6283_ ;
wire _5974_ ;
wire _5554_ ;
wire _5134_ ;
wire _6339_ ;
wire _1894_ ;
wire _1474_ ;
wire _1054_ ;
wire _385_ ;
wire _2679_ ;
wire _2259_ ;
wire _3620_ ;
wire _3200_ ;
wire _6092_ ;
wire _4825_ ;
wire _4405_ ;
wire _5783_ ;
wire _5363_ ;
wire _6148_ ;
wire _1283_ ;
wire _194_ ;
wire _2488_ ;
wire _2068_ ;
wire _4634_ ;
wire _4214_ ;
wire _5839_ ;
wire _5419_ ;
wire _1759_ ;
wire _1339_ ;
wire _2700_ ;
wire _5592_ ;
wire _5172_ ;
wire _3905_ ;
wire [15:0] _6377_ ;
wire _1092_ ;
wire _2297_ ;
wire _4863_ ;
wire _4443_ ;
wire _4023_ ;
wire _5648_ ;
wire _5228_ ;
wire _1988_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire _3714_ ;
wire _6186_ ;
wire _4919_ ;
wire _4672_ ;
wire _4252_ ;
wire _5877_ ;
wire _5457_ ;
wire _5037_ ;
wire _1797_ ;
wire _1377_ ;
wire _288_ ;
wire _3943_ ;
wire _3523_ ;
wire _3103_ ;
wire _4_ ;
wire _4728_ ;
wire _4308_ ;
wire _4481_ ;
wire _4061_ ;
wire _920_ ;
wire _500_ ;
wire _5686_ ;
wire _5266_ ;
wire _1186_ ;
wire _3752_ ;
wire _3332_ ;
wire _4957_ ;
wire _4537_ ;
wire _4117_ ;
wire _4290_ ;
wire _2603_ ;
wire _5495_ ;
wire _5075_ ;
wire _3808_ ;
wire [15:0] _3981_ ;
wire _3561_ ;
wire _3141_ ;
wire _4766_ ;
wire _4346_ ;
wire _45_ ;
wire _2832_ ;
wire _2412_ ;
wire _3617_ ;
wire _6089_ ;
wire [15:0] \u_fir_pe2.rYin  ;
wire _3790_ ;
wire _3370_ ;
wire _4995_ ;
wire _4575_ ;
wire _4155_ ;
wire \X[5]_5_bF$buf0  ;
wire _6301_ ;
wire _2641_ ;
wire _2221_ ;
wire _3846_ ;
wire _3426_ ;
wire _3006_ ;
wire _1912_ ;
wire _4384_ ;
wire _823_ ;
wire _403_ ;
wire _5589_ ;
wire _5169_ ;
wire _83_ ;
wire _6110_ ;
wire _1089_ ;
wire _2870_ ;
wire _2450_ ;
wire _2030_ ;
wire _3655_ ;
wire _3235_ ;
wire _5801_ ;
wire _1721_ ;
wire _1301_ ;
wire _4193_ ;
wire _632_ ;
wire _212_ ;
wire _2926_ ;
wire _2506_ ;
wire _5398_ ;
wire _3884_ ;
wire _3464_ ;
wire _3044_ ;
wire _4669_ ;
wire _4249_ ;
wire _5610_ ;
wire _1950_ ;
wire _1530_ ;
wire _1110_ ;
wire _861_ ;
wire _441_ ;
wire _2735_ ;
wire _2315_ ;
wire _3693_ ;
wire _3273_ ;
wire _4898_ ;
wire _4478_ ;
wire _4058_ ;
wire _917_ ;
wire _6204_ ;
wire _670_ ;
wire _250_ ;
wire _2964_ ;
wire _2544_ ;
wire _2124_ ;
wire _3749_ ;
wire _3329_ ;
wire _3082_ ;
wire _1815_ ;
wire _4287_ ;
wire _726_ ;
wire _306_ ;
wire _6013_ ;
wire _2773_ ;
wire _2353_ ;
wire [15:0] _3978_ ;
wire _3558_ ;
wire _3138_ ;
wire _5704_ ;
wire _1624_ ;
wire _1204_ ;
wire _4096_ ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _2829_ ;
wire _2409_ ;
wire _6242_ ;
wire _2582_ ;
wire _2162_ ;
wire _3787_ ;
wire _3367_ ;
wire _5933_ ;
wire _5513_ ;
wire _1853_ ;
wire _1433_ ;
wire _1013_ ;
wire _764_ ;
wire _344_ ;
wire _2638_ ;
wire _2218_ ;
wire _6051_ ;
wire _2391_ ;
wire _3596_ ;
wire _3176_ ;
wire _1909_ ;
wire _5742_ ;
wire _5322_ ;
wire _6107_ ;
wire _1662_ ;
wire _1242_ ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _2867_ ;
wire _2447_ ;
wire _2027_ ;
wire _6280_ ;
wire _1718_ ;
wire _5971_ ;
wire _5551_ ;
wire _5131_ ;
wire _629_ ;
wire _209_ ;
wire Xin_5_bF$buf0 ;
wire Xin_5_bF$buf1 ;
wire Xin_5_bF$buf2 ;
wire Xin_5_bF$buf3 ;
wire _6336_ ;
wire _1891_ ;
wire _1471_ ;
wire _1051_ ;
wire _382_ ;
wire _2676_ ;
wire _2256_ ;
wire clk_bF$buf50 ;
wire clk_bF$buf51 ;
wire clk_bF$buf52 ;
wire clk_bF$buf53 ;
wire clk_bF$buf54 ;
wire clk_bF$buf55 ;
wire clk_bF$buf56 ;
wire clk_bF$buf57 ;
wire _4822_ ;
wire _4402_ ;
wire _5607_ ;
wire _1947_ ;
wire _1527_ ;
wire _1107_ ;
wire _5780_ ;
wire _5360_ ;
wire _858_ ;
wire _438_ ;
wire _6145_ ;
wire _1280_ ;
wire _191_ ;
wire _2485_ ;
wire _2065_ ;
wire _4631_ ;
wire _4211_ ;
wire _5836_ ;
wire _5416_ ;
wire _1756_ ;
wire _1336_ ;
wire _667_ ;
wire _247_ ;
wire _3902_ ;
wire [15:0] _6374_ ;
wire _2294_ ;
wire _3499_ ;
wire _3079_ ;
wire _4860_ ;
wire _4440_ ;
wire _4020_ ;
wire _5645_ ;
wire _5225_ ;
wire _1985_ ;
wire _1565_ ;
wire _1145_ ;
wire _896_ ;
wire _476_ ;
wire _3711_ ;
wire _6183_ ;
wire _4916_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire clk_bF$buf8 ;
wire clk_bF$buf9 ;
wire _5874_ ;
wire _5454_ ;
wire _5034_ ;
wire _6239_ ;
wire _1794_ ;
wire _1374_ ;
wire _285_ ;
wire _2999_ ;
wire _2579_ ;
wire _2159_ ;
wire _3940_ ;
wire _3520_ ;
wire _3100_ ;
wire _1_ ;
wire _4725_ ;
wire _4305_ ;
wire _5683_ ;
wire _5263_ ;
wire _6048_ ;
wire _1183_ ;
wire [15:0] _2388_ ;
wire _4954_ ;
wire _4534_ ;
wire _4114_ ;
wire _5739_ ;
wire _5319_ ;
wire _1659_ ;
wire _1239_ ;
wire _2600_ ;
wire _5492_ ;
wire _5072_ ;
wire _3805_ ;
wire _6277_ ;
wire _2197_ ;
wire _4763_ ;
wire _4343_ ;
wire _5968_ ;
wire _5548_ ;
wire _5128_ ;
wire _42_ ;
wire _1888_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire _3614_ ;
wire _6086_ ;
wire _4819_ ;
wire _4992_ ;
wire _4572_ ;
wire _4152_ ;
wire _5777_ ;
wire _5357_ ;
wire \X[4]_5_bF$buf2  ;
wire _1697_ ;
wire _1277_ ;
wire _188_ ;
wire _3843_ ;
wire _3423_ ;
wire _3003_ ;
wire _4628_ ;
wire _4208_ ;
wire _4381_ ;
wire _820_ ;
wire _400_ ;
wire _5586_ ;
wire _5166_ ;
wire _80_ ;
wire _1086_ ;
wire _3652_ ;
wire _3232_ ;
wire _4857_ ;
wire _4437_ ;
wire _4017_ ;
wire _4190_ ;
wire [15:0] \u_fir_pe7.rYin  ;
wire _2923_ ;
wire _2503_ ;
wire _5395_ ;
wire _3708_ ;
wire _3881_ ;
wire _3461_ ;
wire _3041_ ;
wire _4666_ ;
wire _4246_ ;
wire _2732_ ;
wire _2312_ ;
wire _3937_ ;
wire _3517_ ;
wire _3690_ ;
wire _3270_ ;
wire _4895_ ;
wire _4475_ ;
wire _4055_ ;
wire _914_ ;
wire _6201_ ;
wire _2961_ ;
wire _2541_ ;
wire _2121_ ;
wire _3746_ ;
wire _3326_ ;
wire _1812_ ;
wire _4284_ ;
wire _723_ ;
wire _303_ ;
wire _5489_ ;
wire _5069_ ;
wire _6010_ ;
wire _2770_ ;
wire _2350_ ;
wire _3975_ ;
wire _3555_ ;
wire _3135_ ;
wire _5701_ ;
wire _39_ ;
wire _1621_ ;
wire _1201_ ;
wire _4093_ ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _2826_ ;
wire _2406_ ;
wire _5298_ ;
wire _3784_ ;
wire _3364_ ;
wire _4989_ ;
wire _4569_ ;
wire _4149_ ;
wire _5930_ ;
wire _5510_ ;
wire _1850_ ;
wire _1430_ ;
wire _1010_ ;
wire _761_ ;
wire _341_ ;
wire _2635_ ;
wire _2215_ ;
wire clk ;
wire _3593_ ;
wire _3173_ ;
wire _1906_ ;
wire _4798_ ;
wire _4378_ ;
wire _817_ ;
wire _77_ ;
wire _6104_ ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _2864_ ;
wire _2444_ ;
wire _2024_ ;
wire _3649_ ;
wire _3229_ ;
wire _1715_ ;
wire _4187_ ;
wire _626_ ;
wire _206_ ;
wire _6333_ ;
wire _2673_ ;
wire _2253_ ;
wire clk_bF$buf20 ;
wire clk_bF$buf21 ;
wire clk_bF$buf22 ;
wire clk_bF$buf23 ;
wire clk_bF$buf24 ;
wire clk_bF$buf25 ;
wire clk_bF$buf26 ;
wire clk_bF$buf27 ;
wire clk_bF$buf28 ;
wire clk_bF$buf29 ;
wire _3878_ ;
wire _3458_ ;
wire _3038_ ;
wire _5604_ ;
wire _1944_ ;
wire _1524_ ;
wire _1104_ ;
wire _855_ ;
wire _435_ ;
wire _2729_ ;
wire _2309_ ;
wire _6142_ ;
wire _2482_ ;
wire _2062_ ;
wire _3687_ ;
wire _3267_ ;
wire _5833_ ;
wire _5413_ ;
wire _1753_ ;
wire _1333_ ;
wire _664_ ;
wire _244_ ;
wire _2958_ ;
wire _2538_ ;
wire _2118_ ;
wire [15:0] _6371_ ;
wire _2291_ ;
wire _3496_ ;
wire _3076_ ;
wire _1809_ ;
wire _5642_ ;
wire _5222_ ;
wire _6007_ ;
wire _1982_ ;
wire _1562_ ;
wire _1142_ ;
wire _893_ ;
wire _473_ ;
wire _2767_ ;
wire _2347_ ;
wire _6180_ ;
wire _4913_ ;
wire _1618_ ;
wire _5871_ ;
wire _5451_ ;
wire _5031_ ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _6236_ ;
wire _1791_ ;
wire _1371_ ;
wire _282_ ;
wire _2996_ ;
wire _2576_ ;
wire _2156_ ;
wire _4722_ ;
wire _4302_ ;
wire _5927_ ;
wire _5507_ ;
wire _1847_ ;
wire _1427_ ;
wire _1007_ ;
wire _5680_ ;
wire _5260_ ;
wire _758_ ;
wire _338_ ;
wire _6045_ ;
wire _1180_ ;
wire [15:0] _2385_ ;
wire _4951_ ;
wire _4531_ ;
wire _4111_ ;
wire _5736_ ;
wire _5316_ ;
wire _1656_ ;
wire _1236_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _3802_ ;
wire _6274_ ;
wire _2194_ ;
wire _3399_ ;
wire _4760_ ;
wire _4340_ ;
wire _5965_ ;
wire _5545_ ;
wire _5125_ ;
wire _1885_ ;
wire _1465_ ;
wire _1045_ ;
wire [15:0] _796_ ;
wire _376_ ;
wire _3611_ ;
wire _6083_ ;
wire _4816_ ;
wire _5774_ ;
wire _5354_ ;
wire _6139_ ;
wire _1694_ ;
wire _1274_ ;
wire _185_ ;
wire _2899_ ;
wire _2479_ ;
wire _2059_ ;
wire _3840_ ;
wire _3420_ ;
wire _3000_ ;
wire _4625_ ;
wire _4205_ ;
wire [15:0] \Y[6]  ;
wire _5583_ ;
wire _5163_ ;
wire [15:0] _6368_ ;
wire _1083_ ;
wire _2288_ ;
wire _4854_ ;
wire _4434_ ;
wire _4014_ ;
wire _5639_ ;
wire _5219_ ;
wire _1979_ ;
wire _1559_ ;
wire _1139_ ;
wire _2920_ ;
wire _2500_ ;
wire _5392_ ;
wire _3705_ ;
wire _6177_ ;
wire _2097_ ;
wire _4663_ ;
wire _4243_ ;
wire _5868_ ;
wire _5448_ ;
wire _5028_ ;
wire _1788_ ;
wire _1368_ ;
wire _699_ ;
wire _279_ ;
wire _3934_ ;
wire _3514_ ;
wire _4719_ ;
wire _4892_ ;
wire _4472_ ;
wire _4052_ ;
wire _911_ ;
wire _5677_ ;
wire _5257_ ;
wire _1597_ ;
wire _1177_ ;
wire _3743_ ;
wire _3323_ ;
wire _4948_ ;
wire _4528_ ;
wire _4108_ ;
wire _4281_ ;
wire _720_ ;
wire _300_ ;
wire _5486_ ;
wire _5066_ ;
wire _3972_ ;
wire _3552_ ;
wire _3132_ ;
wire _4757_ ;
wire _4337_ ;
wire _36_ ;
wire _4090_ ;
wire _2823_ ;
wire _2403_ ;
wire _5295_ ;
wire _3608_ ;
wire _3781_ ;
wire _3361_ ;
wire _4986_ ;
wire _4566_ ;
wire _4146_ ;
wire _2632_ ;
wire _2212_ ;
wire _3837_ ;
wire _3417_ ;
wire _3590_ ;
wire _3170_ ;
wire _1903_ ;
wire _4795_ ;
wire _4375_ ;
wire _814_ ;
wire _74_ ;
wire _6101_ ;
wire _2861_ ;
wire _2441_ ;
wire _2021_ ;
wire _3646_ ;
wire _3226_ ;
wire _1712_ ;
wire _4184_ ;
wire _623_ ;
wire _203_ ;
wire _2917_ ;
wire _5389_ ;
wire _6330_ ;
wire _2670_ ;
wire _2250_ ;
wire _3875_ ;
wire _3455_ ;
wire _3035_ ;
wire _5601_ ;
wire _1941_ ;
wire _1521_ ;
wire _1101_ ;
wire _852_ ;
wire _432_ ;
wire _2726_ ;
wire _2306_ ;
wire _5198_ ;
wire _3684_ ;
wire _3264_ ;
wire _4889_ ;
wire _4469_ ;
wire _4049_ ;
wire _5830_ ;
wire _5410_ ;
wire _908_ ;
wire _1750_ ;
wire _1330_ ;
wire _661_ ;
wire _241_ ;
wire _2955_ ;
wire _2535_ ;
wire _2115_ ;
wire _3493_ ;
wire _3073_ ;
wire _1806_ ;
wire _4698_ ;
wire _4278_ ;
wire _717_ ;
wire _6004_ ;
wire _890_ ;
wire _470_ ;
wire _2764_ ;
wire _2344_ ;
wire _3969_ ;
wire _3549_ ;
wire _3129_ ;
wire _4910_ ;
wire _1615_ ;
wire _4087_ ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _6233_ ;
wire _2993_ ;
wire _2573_ ;
wire _2153_ ;
wire _3778_ ;
wire _3358_ ;
wire _5924_ ;
wire _5504_ ;
wire _1844_ ;
wire _1424_ ;
wire _1004_ ;
wire _755_ ;
wire _335_ ;
wire _2629_ ;
wire _2209_ ;
wire _6042_ ;
wire _2382_ ;
wire _3587_ ;
wire _3167_ ;
wire _5733_ ;
wire _5313_ ;
wire _1653_ ;
wire _1233_ ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _2858_ ;
wire _2438_ ;
wire _2018_ ;
wire _6271_ ;
wire _2191_ ;
wire _3396_ ;
wire _1709_ ;
wire _5962_ ;
wire _5542_ ;
wire _5122_ ;
wire _6327_ ;
wire _1882_ ;
wire _1462_ ;
wire _1042_ ;
wire [15:0] _793_ ;
wire _373_ ;
wire _2667_ ;
wire _2247_ ;
wire _6080_ ;
wire _4813_ ;
wire _1938_ ;
wire _1518_ ;
wire _5771_ ;
wire _5351_ ;
wire _849_ ;
wire _429_ ;
wire \X[3]_5_bF$buf1  ;
wire _6136_ ;
wire _1691_ ;
wire _1271_ ;
wire _182_ ;
wire _2896_ ;
wire _2476_ ;
wire _2056_ ;
wire _4622_ ;
wire _4202_ ;
wire _5827_ ;
wire _5407_ ;
wire _1747_ ;
wire _1327_ ;
wire _5580_ ;
wire _5160_ ;
wire _658_ ;
wire _238_ ;
wire _6365_ ;
wire _1080_ ;
wire [15:0] \u_fir_pe5.rYin  ;
wire _2285_ ;
wire _4851_ ;
wire _4431_ ;
wire _4011_ ;
wire _5636_ ;
wire _5216_ ;
wire _1976_ ;
wire _1556_ ;
wire _1136_ ;
wire _887_ ;
wire _467_ ;
wire _3702_ ;
wire _6174_ ;
wire _4907_ ;
wire _2094_ ;
wire _3299_ ;
wire _4660_ ;
wire _4240_ ;
wire _5865_ ;
wire _5445_ ;
wire _5025_ ;
wire _1785_ ;
wire _1365_ ;
wire _696_ ;
wire _276_ ;
wire _3931_ ;
wire _3511_ ;
wire _4716_ ;
wire _5674_ ;
wire _5254_ ;
wire _6039_ ;
wire _1594_ ;
wire _1174_ ;
wire _2799_ ;
wire _2379_ ;
wire _3740_ ;
wire _3320_ ;
wire _4945_ ;
wire _4525_ ;
wire _4105_ ;
wire _5483_ ;
wire _5063_ ;
wire _6268_ ;
wire _2188_ ;
wire _4754_ ;
wire _4334_ ;
wire _5959_ ;
wire _5539_ ;
wire _5119_ ;
wire _33_ ;
wire _1879_ ;
wire _1459_ ;
wire _1039_ ;
wire _2820_ ;
wire _2400_ ;
wire _5292_ ;
wire _3605_ ;
wire _6077_ ;
wire [7:0] \X[4]  ;
wire _4983_ ;
wire _4563_ ;
wire _4143_ ;
wire _5768_ ;
wire _5348_ ;
wire _1688_ ;
wire _1268_ ;
wire _599_ ;
wire _179_ ;
wire _3834_ ;
wire _3414_ ;
wire _4619_ ;
wire _1900_ ;
wire _4792_ ;
wire _4372_ ;
wire _811_ ;
wire _5997_ ;
wire [15:0] _5577_ ;
wire _5157_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire _3643_ ;
wire _3223_ ;
wire _4848_ ;
wire _4428_ ;
wire _4008_ ;
wire _4181_ ;
wire _620_ ;
wire _200_ ;
wire _2914_ ;
wire _5386_ ;
wire _3872_ ;
wire _3452_ ;
wire _3032_ ;
wire _4657_ ;
wire _4237_ ;
wire _2723_ ;
wire _2303_ ;
wire _5195_ ;
wire _3928_ ;
wire _3508_ ;
wire _3681_ ;
wire _3261_ ;
wire _4886_ ;
wire _4466_ ;
wire _4046_ ;
wire _905_ ;
wire _2952_ ;
wire _2532_ ;
wire _2112_ ;
wire _3737_ ;
wire _3317_ ;
wire _3490_ ;
wire _3070_ ;
wire _1803_ ;
wire _4695_ ;
wire _4275_ ;
wire _714_ ;
wire _6001_ ;
wire _2761_ ;
wire _2341_ ;
wire _3966_ ;
wire _3546_ ;
wire _3126_ ;
wire _1612_ ;
wire _4084_ ;
wire _943_ ;
wire _523_ ;
wire _103_ ;
wire _2817_ ;
wire _5289_ ;
wire _6230_ ;
wire _2990_ ;
wire _2570_ ;
wire _2150_ ;
wire _3775_ ;
wire _3355_ ;
wire _5921_ ;
wire _5501_ ;
wire _1841_ ;
wire _1421_ ;
wire _1001_ ;
wire _752_ ;
wire _332_ ;
wire _2626_ ;
wire _2206_ ;
wire _5098_ ;
wire _3584_ ;
wire _3164_ ;
wire _4789_ ;
wire _4369_ ;
wire _5730_ ;
wire _5310_ ;
wire _808_ ;
wire _68_ ;
wire _1650_ ;
wire _1230_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _2855_ ;
wire _2435_ ;
wire _2015_ ;
wire _3393_ ;
wire _1706_ ;
wire _4598_ ;
wire _4178_ ;
wire _617_ ;
wire _6324_ ;
wire [15:0] _790_ ;
wire _370_ ;
wire _2664_ ;
wire _2244_ ;
wire _3869_ ;
wire _3449_ ;
wire _3029_ ;
wire _4810_ ;
wire _1935_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire \X[2]_5_bF$buf3  ;
wire _6133_ ;
wire _2893_ ;
wire _2473_ ;
wire _2053_ ;
wire _3678_ ;
wire _3258_ ;
wire _5824_ ;
wire _5404_ ;
wire _1744_ ;
wire _1324_ ;
wire _655_ ;
wire _235_ ;
wire _2949_ ;
wire _2529_ ;
wire _2109_ ;
wire _6362_ ;
wire _2282_ ;
wire _3487_ ;
wire _3067_ ;
wire _5633_ ;
wire _5213_ ;
wire _1973_ ;
wire _1553_ ;
wire _1133_ ;
wire _884_ ;
wire _464_ ;
wire _2758_ ;
wire _2338_ ;
wire _6171_ ;
wire _4904_ ;
wire _2091_ ;
wire _3296_ ;
wire _1609_ ;
wire _5862_ ;
wire _5442_ ;
wire _5022_ ;
wire _6227_ ;
wire _1782_ ;
wire _1362_ ;
wire _693_ ;
wire _273_ ;
wire _2987_ ;
wire _2567_ ;
wire _2147_ ;
wire _4713_ ;
wire _5918_ ;
wire _1838_ ;
wire _1418_ ;
wire _5671_ ;
wire _5251_ ;
wire _749_ ;
wire _329_ ;
wire _6036_ ;
wire [15:0] _1591_ ;
wire _1171_ ;
wire _2796_ ;
wire _2376_ ;
wire _4942_ ;
wire _4522_ ;
wire _4102_ ;
wire _5727_ ;
wire _5307_ ;
wire _1647_ ;
wire _1227_ ;
wire _5480_ ;
wire _5060_ ;
wire _978_ ;
wire _558_ ;
wire _138_ ;
wire _6265_ ;
wire _2185_ ;
wire _4751_ ;
wire _4331_ ;
wire _5956_ ;
wire _5536_ ;
wire _5116_ ;
wire _30_ ;
wire _1876_ ;
wire _1456_ ;
wire _1036_ ;
wire _787_ ;
wire _367_ ;
wire _3602_ ;
wire _6074_ ;
wire _4807_ ;
wire _3199_ ;
wire _4980_ ;
wire _4560_ ;
wire _4140_ ;
wire _5765_ ;
wire _5345_ ;
wire _1685_ ;
wire _1265_ ;
wire _596_ ;
wire _176_ ;
wire _3831_ ;
wire _3411_ ;
wire _4616_ ;
wire _5994_ ;
wire [15:0] _5574_ ;
wire _5154_ ;
wire _6359_ ;
wire _1494_ ;
wire _1074_ ;
wire _2699_ ;
wire _2279_ ;
wire _3640_ ;
wire _3220_ ;
wire _4845_ ;
wire _4425_ ;
wire _4005_ ;
wire _2911_ ;
wire _5383_ ;
wire _6168_ ;
wire clk_hier0_bF$buf0 ;
wire clk_hier0_bF$buf1 ;
wire clk_hier0_bF$buf2 ;
wire clk_hier0_bF$buf3 ;
wire clk_hier0_bF$buf4 ;
wire clk_hier0_bF$buf5 ;
wire clk_hier0_bF$buf6 ;
wire _2088_ ;
wire _4654_ ;
wire _4234_ ;
wire _5859_ ;
wire _5439_ ;
wire _5019_ ;
wire _1779_ ;
wire _1359_ ;
wire _2720_ ;
wire _2300_ ;
wire _5192_ ;
wire _3925_ ;
wire _3505_ ;
wire _4883_ ;
wire _4463_ ;
wire _4043_ ;
wire _902_ ;
wire _5668_ ;
wire _5248_ ;
wire [15:0] _1588_ ;
wire _1168_ ;
wire _499_ ;
wire _3734_ ;
wire _3314_ ;
wire _4939_ ;
wire _4519_ ;
wire _1800_ ;
wire _4692_ ;
wire _4272_ ;
wire _711_ ;
wire _5897_ ;
wire _5477_ ;
wire _5057_ ;
wire _1397_ ;
wire _3963_ ;
wire _3543_ ;
wire _3123_ ;
wire _4748_ ;
wire _4328_ ;
wire _27_ ;
wire _4081_ ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire _2814_ ;
wire _5286_ ;
wire _3772_ ;
wire _3352_ ;
wire _4977_ ;
wire _4557_ ;
wire _4137_ ;
wire _2623_ ;
wire _2203_ ;
wire _5095_ ;
wire _3828_ ;
wire _3408_ ;
wire _3581_ ;
wire _3161_ ;
wire _4786_ ;
wire _4366_ ;
wire _805_ ;
wire _65_ ;
wire _2852_ ;
wire _2432_ ;
wire _2012_ ;
wire _3637_ ;
wire _3217_ ;
wire _3390_ ;
wire _1703_ ;
wire _4595_ ;
wire _4175_ ;
wire _614_ ;
wire _2908_ ;
wire _6321_ ;
wire _2661_ ;
wire _2241_ ;
wire _3866_ ;
wire _3446_ ;
wire _3026_ ;
wire _1932_ ;
wire _1512_ ;
wire _843_ ;
wire _423_ ;
wire _2717_ ;
wire _5189_ ;
wire \X[2]_5_bF$buf0  ;
wire _6130_ ;
wire _2890_ ;
wire _2470_ ;
wire _2050_ ;
wire _3675_ ;
wire _3255_ ;
wire _5821_ ;
wire _5401_ ;
wire _1741_ ;
wire _1321_ ;
wire _652_ ;
wire _232_ ;
wire _2946_ ;
wire _2526_ ;
wire _2106_ ;
wire _3484_ ;
wire _3064_ ;
wire _4689_ ;
wire _4269_ ;
wire _5630_ ;
wire _5210_ ;
wire _708_ ;
wire _1970_ ;
wire _1550_ ;
wire _1130_ ;
wire _881_ ;
wire _461_ ;
wire _2755_ ;
wire _2335_ ;
wire _4901_ ;
wire _3293_ ;
wire _1606_ ;
wire _4498_ ;
wire _4078_ ;
wire _937_ ;
wire _517_ ;
wire _6224_ ;
wire _690_ ;
wire _270_ ;
wire _2984_ ;
wire _2564_ ;
wire _2144_ ;
wire _3769_ ;
wire _3349_ ;
wire _4710_ ;
wire _5915_ ;
wire _1835_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _6033_ ;
wire _2793_ ;
wire _2373_ ;
wire _3998_ ;
wire _3578_ ;
wire _3158_ ;
wire _5724_ ;
wire _5304_ ;
wire _1644_ ;
wire _1224_ ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire _2849_ ;
wire _2429_ ;
wire _2009_ ;
wire _6262_ ;
wire _2182_ ;
wire [15:0] \Y[1]  ;
wire _3387_ ;
wire _5953_ ;
wire _5533_ ;
wire _5113_ ;
wire _6318_ ;
wire _1873_ ;
wire _1453_ ;
wire _1033_ ;
wire _784_ ;
wire _364_ ;
wire _2658_ ;
wire _2238_ ;
wire _6071_ ;
wire _4804_ ;
wire _3196_ ;
wire _1929_ ;
wire _1509_ ;
wire _5762_ ;
wire _5342_ ;
wire _6127_ ;
wire _1682_ ;
wire _1262_ ;
wire _593_ ;
wire _173_ ;
wire _2887_ ;
wire _2467_ ;
wire _2047_ ;
wire _4613_ ;
wire _5818_ ;
wire _1738_ ;
wire _1318_ ;
wire _5991_ ;
wire [15:0] _5571_ ;
wire _5151_ ;
wire _649_ ;
wire _229_ ;
wire _6356_ ;
wire _1491_ ;
wire _1071_ ;
wire _2696_ ;
wire _2276_ ;
wire _4842_ ;
wire _4422_ ;
wire _4002_ ;
wire _5627_ ;
wire _5207_ ;
wire _1967_ ;
wire _1547_ ;
wire _1127_ ;
wire _5380_ ;
wire _878_ ;
wire _458_ ;
wire _6165_ ;
wire _2085_ ;
wire _4651_ ;
wire _4231_ ;
wire _5856_ ;
wire _5436_ ;
wire _5016_ ;
wire _1776_ ;
wire _1356_ ;
wire _687_ ;
wire _267_ ;
wire _3922_ ;
wire _3502_ ;
wire _4707_ ;
wire _3099_ ;
wire _4880_ ;
wire _4460_ ;
wire _4040_ ;
wire _5665_ ;
wire _5245_ ;
wire _1585_ ;
wire _1165_ ;
wire _496_ ;
wire _3731_ ;
wire _3311_ ;
wire _4936_ ;
wire _4516_ ;
wire _5894_ ;
wire _5474_ ;
wire _5054_ ;
wire _6259_ ;
wire _1394_ ;
wire _2599_ ;
wire _2179_ ;
wire _3960_ ;
wire _3540_ ;
wire _3120_ ;
wire _4745_ ;
wire _4325_ ;
wire _24_ ;
wire _2811_ ;
wire _5283_ ;
wire _6068_ ;
wire _4974_ ;
wire _4554_ ;
wire _4134_ ;
wire _5759_ ;
wire _5339_ ;
wire _1679_ ;
wire _1259_ ;
wire _2620_ ;
wire _2200_ ;
wire _5092_ ;
wire _3825_ ;
wire _3405_ ;
wire _6297_ ;
wire _4783_ ;
wire _4363_ ;
wire _802_ ;
wire _5988_ ;
wire _5568_ ;
wire _5148_ ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire _399_ ;
wire _3634_ ;
wire _3214_ ;
wire _4839_ ;
wire _4419_ ;
wire _1700_ ;
wire _4592_ ;
wire _4172_ ;
wire _611_ ;
wire _2905_ ;
wire _5797_ ;
wire _5377_ ;
wire _1297_ ;
wire _3863_ ;
wire _3443_ ;
wire _3023_ ;
wire _4648_ ;
wire _4228_ ;
wire _840_ ;
wire _420_ ;
wire _2714_ ;
wire _5186_ ;
wire \X[1]_5_bF$buf2  ;
wire _3919_ ;
wire _3672_ ;
wire _3252_ ;
wire _4877_ ;
wire _4457_ ;
wire _4037_ ;
wire _2943_ ;
wire _2523_ ;
wire _2103_ ;
wire _3728_ ;
wire _3308_ ;
wire _3481_ ;
wire _3061_ ;
wire _4686_ ;
wire _4266_ ;
wire _705_ ;
wire _2752_ ;
wire _2332_ ;
wire _3957_ ;
wire _3537_ ;
wire _3117_ ;
wire _3290_ ;
wire _1603_ ;
wire _4495_ ;
wire _4075_ ;
wire _934_ ;
wire _514_ ;
wire _2808_ ;
wire _6221_ ;
wire _2981_ ;
wire _2561_ ;
wire _2141_ ;
wire _3766_ ;
wire _3346_ ;
wire _5912_ ;
wire _1832_ ;
wire _1412_ ;
wire _743_ ;
wire _323_ ;
wire _2617_ ;
wire _5089_ ;
wire _6030_ ;
wire _2790_ ;
wire _2370_ ;
wire _3995_ ;
wire _3575_ ;
wire _3155_ ;
wire _5721_ ;
wire _5301_ ;
wire _59_ ;
wire _1641_ ;
wire _1221_ ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _2846_ ;
wire _2426_ ;
wire _2006_ ;
wire _3384_ ;
wire _4589_ ;
wire _4169_ ;
wire _5950_ ;
wire _5530_ ;
wire _5110_ ;
wire _608_ ;
wire _6315_ ;
wire _1870_ ;
wire _1450_ ;
wire _1030_ ;
wire _781_ ;
wire _361_ ;
wire _2655_ ;
wire _2235_ ;
wire _4801_ ;
wire _3193_ ;
wire _1926_ ;
wire _1506_ ;
wire _4398_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _6124_ ;
wire _590_ ;
wire _170_ ;
wire _2884_ ;
wire _2464_ ;
wire _2044_ ;
wire _3669_ ;
wire _3249_ ;
wire _4610_ ;
wire _5815_ ;
wire _1735_ ;
wire _1315_ ;
wire _646_ ;
wire _226_ ;
wire _6353_ ;
wire _2693_ ;
wire _2273_ ;
wire _3898_ ;
wire _3478_ ;
wire _3058_ ;
wire _5624_ ;
wire _5204_ ;
wire _1964_ ;
wire _1544_ ;
wire _1124_ ;
wire _875_ ;
wire _455_ ;
wire _2749_ ;
wire _2329_ ;
wire _6162_ ;
wire _2082_ ;
wire _3287_ ;
wire _5853_ ;
wire _5433_ ;
wire _5013_ ;
wire _6218_ ;
wire _1773_ ;
wire _1353_ ;
wire _684_ ;
wire _264_ ;
wire _2978_ ;
wire _2558_ ;
wire _2138_ ;
wire _4704_ ;
wire _5909_ ;
wire _3096_ ;
wire _1829_ ;
wire _1409_ ;
wire _5662_ ;
wire _5242_ ;
wire _6027_ ;
wire _1582_ ;
wire _1162_ ;
wire _493_ ;
wire _2787_ ;
wire _2367_ ;
wire _4933_ ;
wire _4513_ ;
wire _5718_ ;
wire _1638_ ;
wire _1218_ ;
wire _5891_ ;
wire _5471_ ;
wire _5051_ ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire _6256_ ;
wire _1391_ ;
wire _2596_ ;
wire _2176_ ;
wire _4742_ ;
wire _4322_ ;
wire \X[7]_5_bF$buf1  ;
wire _5947_ ;
wire _5527_ ;
wire _5107_ ;
wire _21_ ;
wire _1867_ ;
wire _1447_ ;
wire _1027_ ;
wire _5280_ ;
wire _778_ ;
wire _358_ ;
wire _6065_ ;
wire _4971_ ;
wire _4551_ ;
wire _4131_ ;
wire _5756_ ;
wire _5336_ ;
wire _1676_ ;
wire _1256_ ;
wire _587_ ;
wire _167_ ;
wire _3822_ ;
wire _3402_ ;
wire _6294_ ;
wire _4607_ ;
wire [15:0] _4780_ ;
wire _4360_ ;
wire _5985_ ;
wire _5565_ ;
wire _5145_ ;
wire _1485_ ;
wire _1065_ ;
wire _396_ ;
wire _3631_ ;
wire _3211_ ;
wire _4836_ ;
wire _4416_ ;
wire _2902_ ;
wire _5794_ ;
wire _5374_ ;
wire _6159_ ;
wire _1294_ ;
wire _2499_ ;
wire _2079_ ;
wire _3860_ ;
wire _3440_ ;
wire _3020_ ;
wire _4645_ ;
wire _4225_ ;
wire _2711_ ;
wire _5183_ ;
wire _3916_ ;
wire _4874_ ;
wire _4454_ ;
wire _4034_ ;
wire _5659_ ;
wire _5239_ ;
wire _1999_ ;
wire _1579_ ;
wire _1159_ ;
wire _2940_ ;
wire _2520_ ;
wire _2100_ ;
wire _3725_ ;
wire _3305_ ;
wire _6197_ ;
wire _4683_ ;
wire _4263_ ;
wire _702_ ;
wire _5888_ ;
wire _5468_ ;
wire _5048_ ;
wire _1388_ ;
wire _299_ ;
wire _3954_ ;
wire _3534_ ;
wire _3114_ ;
wire _4739_ ;
wire _4319_ ;
wire _18_ ;
wire _1600_ ;
wire _4492_ ;
wire _4072_ ;
wire _931_ ;
wire _511_ ;
wire _2805_ ;
wire _5697_ ;
wire _5277_ ;
wire _1197_ ;
wire _3763_ ;
wire _3343_ ;
wire _4968_ ;
wire _4548_ ;
wire _4128_ ;
wire _740_ ;
wire _320_ ;
wire _2614_ ;
wire _5086_ ;
wire _3819_ ;
wire _3992_ ;
wire _3572_ ;
wire _3152_ ;
wire [15:0] _4777_ ;
wire _4357_ ;
wire _56_ ;
wire _2843_ ;
wire _2423_ ;
wire _2003_ ;
wire _3628_ ;
wire _3208_ ;
wire _3381_ ;
wire _4586_ ;
wire _4166_ ;
wire _605_ ;
wire _6312_ ;
wire _2652_ ;
wire _2232_ ;
wire _3857_ ;
wire _3437_ ;
wire _3017_ ;
wire _3190_ ;
wire _1923_ ;
wire _1503_ ;
wire _4395_ ;
wire _834_ ;
wire _414_ ;
wire _2708_ ;
wire _94_ ;
wire _6121_ ;
wire _2881_ ;
wire _2461_ ;
wire _2041_ ;
wire _3666_ ;
wire _3246_ ;
wire _5812_ ;
wire _1732_ ;
wire _1312_ ;
wire _643_ ;
wire _223_ ;
wire _2937_ ;
wire _2517_ ;
wire _6350_ ;
wire [15:0] \u_fir_pe5.mul  ;
wire _2690_ ;
wire _2270_ ;
wire _3895_ ;
wire _3475_ ;
wire _3055_ ;
wire _5621_ ;
wire _5201_ ;
wire _1961_ ;
wire _1541_ ;
wire _1121_ ;
wire _872_ ;
wire _452_ ;
wire _2746_ ;
wire _2326_ ;
wire _3284_ ;
wire _4489_ ;
wire _4069_ ;
wire _5850_ ;
wire _5430_ ;
wire _5010_ ;
wire _928_ ;
wire _508_ ;
wire _6215_ ;
wire _1770_ ;
wire _1350_ ;
wire _681_ ;
wire _261_ ;
wire _2975_ ;
wire _2555_ ;
wire _2135_ ;
wire _4701_ ;
wire _5906_ ;
wire _3093_ ;
wire _1826_ ;
wire _1406_ ;
wire _4298_ ;
wire _737_ ;
wire _317_ ;
wire _6024_ ;
wire _490_ ;
wire _2784_ ;
wire _2364_ ;
wire _3989_ ;
wire _3569_ ;
wire _3149_ ;
wire _4930_ ;
wire _4510_ ;
wire _5715_ ;
wire _1635_ ;
wire _1215_ ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire _6253_ ;
wire _2593_ ;
wire _2173_ ;
wire _3798_ ;
wire _3378_ ;
wire _5944_ ;
wire _5524_ ;
wire _5104_ ;
wire \X[6]_5_bF$buf3  ;
wire _6309_ ;
wire _1864_ ;
wire _1444_ ;
wire _1024_ ;
wire _775_ ;
wire _355_ ;
wire _2649_ ;
wire _2229_ ;
wire _6062_ ;
wire [15:0] \u_fir_pe7.mul  ;
wire [15:0] _3187_ ;
wire _5753_ ;
wire _5333_ ;
wire _6118_ ;
wire _1673_ ;
wire _1253_ ;
wire _584_ ;
wire _164_ ;
wire _2878_ ;
wire _2458_ ;
wire _2038_ ;
wire _6291_ ;
wire _4604_ ;
wire _5809_ ;
wire _1729_ ;
wire _1309_ ;
wire _5982_ ;
wire _5562_ ;
wire _5142_ ;
wire _6347_ ;
wire _1482_ ;
wire _1062_ ;
wire _393_ ;
wire _2687_ ;
wire _2267_ ;
wire _4833_ ;
wire _4413_ ;
wire _5618_ ;
wire _1958_ ;
wire _1538_ ;
wire _1118_ ;
wire _5791_ ;
wire _5371_ ;
wire _869_ ;
wire _449_ ;
wire _6156_ ;
wire _1291_ ;
wire _2496_ ;
wire _2076_ ;
wire _4642_ ;
wire _4222_ ;
wire _5847_ ;
wire _5427_ ;
wire _5007_ ;
wire _1767_ ;
wire _1347_ ;
wire _5180_ ;
wire _678_ ;
wire _258_ ;
wire _3913_ ;
wire _4871_ ;
wire _4451_ ;
wire _4031_ ;
wire _5656_ ;
wire _5236_ ;
wire _1996_ ;
wire _1576_ ;
wire _1156_ ;
wire _487_ ;
wire _3722_ ;
wire _3302_ ;
wire _6194_ ;
wire _4927_ ;
wire _4507_ ;
wire _4680_ ;
wire _4260_ ;
wire _5885_ ;
wire _5465_ ;
wire _5045_ ;
wire _1385_ ;
wire _296_ ;
wire _3951_ ;
wire _3531_ ;
wire _3111_ ;
wire _4736_ ;
wire _4316_ ;
wire _15_ ;
wire _2802_ ;
wire _5694_ ;
wire _5274_ ;
wire _6059_ ;
wire _1194_ ;
wire _2399_ ;
wire _3760_ ;
wire _3340_ ;
wire _4965_ ;
wire _4545_ ;
wire _4125_ ;
wire _2611_ ;
wire _5083_ ;
wire _3816_ ;
wire _6288_ ;
wire [15:0] _4774_ ;
wire _4354_ ;
wire _5979_ ;
wire _5559_ ;
wire _5139_ ;
wire _53_ ;
wire _1899_ ;
wire _1479_ ;
wire _1059_ ;
wire _2840_ ;
wire _2420_ ;
wire _2000_ ;
wire _3625_ ;
wire _3205_ ;
wire _6097_ ;
wire [7:0] \X[6]  ;
wire _4583_ ;
wire _4163_ ;
wire _602_ ;
wire _5788_ ;
wire _5368_ ;
wire _1288_ ;
wire _199_ ;
wire _3854_ ;
wire _3434_ ;
wire _3014_ ;
wire _4639_ ;
wire _4219_ ;
wire _1920_ ;
wire _1500_ ;
wire _4392_ ;
wire _831_ ;
wire _411_ ;
wire _2705_ ;
wire _5597_ ;
wire _5177_ ;
wire _91_ ;
wire _1097_ ;
wire _3663_ ;
wire _3243_ ;
wire _4868_ ;
wire _4448_ ;
wire _4028_ ;
wire _640_ ;
wire _220_ ;
wire _2934_ ;
wire _2514_ ;
wire _3719_ ;
wire _3892_ ;
wire _3472_ ;
wire _3052_ ;
wire _4677_ ;
wire _4257_ ;
wire _2743_ ;
wire _2323_ ;
wire _3948_ ;
wire _3528_ ;
wire _3108_ ;
wire _9_ ;
wire _3281_ ;
wire _4486_ ;
wire _4066_ ;
wire _925_ ;
wire _505_ ;
wire _6212_ ;
wire _2972_ ;
wire _2552_ ;
wire _2132_ ;
wire _3757_ ;
wire _3337_ ;
wire _5903_ ;
wire _3090_ ;
wire _1823_ ;
wire _1403_ ;
wire _4295_ ;
wire _734_ ;
wire _314_ ;
wire _2608_ ;
wire _6021_ ;
wire _2781_ ;
wire _2361_ ;
wire _3986_ ;
wire _3566_ ;
wire _3146_ ;
wire _5712_ ;
wire _1632_ ;
wire _1212_ ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _2837_ ;
wire _2417_ ;
wire _6250_ ;
wire _2590_ ;
wire _2170_ ;
wire _3795_ ;
wire _3375_ ;
wire _5941_ ;
wire _5521_ ;
wire _5101_ ;
wire \X[6]_5_bF$buf0  ;
wire _6306_ ;
wire _1861_ ;
wire _1441_ ;
wire _1021_ ;
wire _772_ ;
wire _352_ ;
wire _2646_ ;
wire _2226_ ;
wire [15:0] _3184_ ;
wire _1917_ ;
wire _4389_ ;
wire _5750_ ;
wire _5330_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _6115_ ;
wire _1670_ ;
wire _1250_ ;
wire _581_ ;
wire _161_ ;
wire _2875_ ;
wire _2455_ ;
wire _2035_ ;
wire _4601_ ;
wire _5806_ ;
wire _1726_ ;
wire _1306_ ;
wire _4198_ ;
wire _637_ ;
wire _217_ ;
wire _6344_ ;
wire _390_ ;
wire _2684_ ;
wire _2264_ ;
wire _3889_ ;
wire _3469_ ;
wire _3049_ ;
wire _4830_ ;
wire _4410_ ;
wire _5615_ ;
wire _1955_ ;
wire _1535_ ;
wire _1115_ ;
wire _866_ ;
wire _446_ ;
wire _6153_ ;
wire _2493_ ;
wire _2073_ ;
wire _3698_ ;
wire _3278_ ;
wire _5844_ ;
wire _5424_ ;
wire _5004_ ;
wire _6209_ ;
wire _1764_ ;
wire _1344_ ;
wire [15:0] Yin ;
wire _675_ ;
wire _255_ ;
wire _2969_ ;
wire _2549_ ;
wire _2129_ ;
wire _3910_ ;
wire _3087_ ;
wire _5653_ ;
wire _5233_ ;
wire _6018_ ;
wire _1993_ ;
wire _1573_ ;
wire _1153_ ;
wire _484_ ;
wire _2778_ ;
wire _2358_ ;
wire _6191_ ;
wire _4924_ ;
wire _4504_ ;
wire _5709_ ;
wire _1629_ ;
wire _1209_ ;
wire _5882_ ;
wire _5462_ ;
wire _5042_ ;
wire _6247_ ;
wire _1382_ ;
wire _293_ ;
wire _2587_ ;
wire _2167_ ;
wire _4733_ ;
wire _4313_ ;
wire _5938_ ;
wire _5518_ ;
wire _12_ ;
wire _1858_ ;
wire _1438_ ;
wire _1018_ ;
wire _5691_ ;
wire _5271_ ;
wire _769_ ;
wire _349_ ;
wire _6056_ ;
wire _1191_ ;
wire _2396_ ;
wire _4962_ ;
wire _4542_ ;
wire _4122_ ;
wire _5747_ ;
wire _5327_ ;
wire _1667_ ;
wire _1247_ ;
wire _5080_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _3813_ ;
wire _6285_ ;
wire _4771_ ;
wire _4351_ ;
wire _5976_ ;
wire _5556_ ;
wire _5136_ ;
wire _50_ ;
wire _1896_ ;
wire _1476_ ;
wire _1056_ ;
wire _387_ ;
wire _3622_ ;
wire _3202_ ;
wire _6094_ ;
wire _4827_ ;
wire _4407_ ;
wire _4580_ ;
wire _4160_ ;
wire _5785_ ;
wire _5365_ ;
wire _1285_ ;
wire _196_ ;
wire _3851_ ;
wire _3431_ ;
wire _3011_ ;
wire _4636_ ;
wire _4216_ ;
wire _2702_ ;
wire _5594_ ;
wire _5174_ ;
wire _3907_ ;
wire _1094_ ;
wire _2299_ ;
wire _3660_ ;
wire _3240_ ;
wire _4865_ ;
wire _4445_ ;
wire _4025_ ;
wire _2931_ ;
wire _2511_ ;
wire _3716_ ;
wire _6188_ ;
wire _4674_ ;
wire _4254_ ;
wire _5879_ ;
wire _5459_ ;
wire _5039_ ;
wire _1799_ ;
wire _1379_ ;
wire _2740_ ;
wire _2320_ ;
wire _3945_ ;
wire _3525_ ;
wire _3105_ ;
wire _6_ ;
wire _4483_ ;
wire _4063_ ;
wire _922_ ;
wire _502_ ;
wire _5688_ ;
wire _5268_ ;
wire _1188_ ;
wire _3754_ ;
wire _3334_ ;
wire _4959_ ;
wire _4539_ ;
wire _4119_ ;
wire _5900_ ;
wire _1820_ ;
wire _1400_ ;
wire _4292_ ;
wire _731_ ;
wire _311_ ;
wire _2605_ ;
wire _5497_ ;
wire _5077_ ;
wire [15:0] _3983_ ;
wire _3563_ ;
wire _3143_ ;
wire _4768_ ;
wire _4348_ ;
wire _47_ ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _2834_ ;
wire _2414_ ;
wire _3619_ ;
wire _3792_ ;
wire _3372_ ;
wire _4997_ ;
wire _4577_ ;
wire _4157_ ;
wire \X[5]_5_bF$buf2  ;
wire _6303_ ;
wire _2643_ ;
wire _2223_ ;
wire _3848_ ;
wire _3428_ ;
wire _3008_ ;
wire [15:0] _3181_ ;
wire _1914_ ;
wire _4386_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _6112_ ;
wire _2872_ ;
wire _2452_ ;
wire _2032_ ;
wire _3657_ ;
wire _3237_ ;
wire _5803_ ;
wire _1723_ ;
wire _1303_ ;
wire _4195_ ;
wire _634_ ;
wire _214_ ;
wire _2928_ ;
wire _2508_ ;
wire _6341_ ;
wire _2681_ ;
wire _2261_ ;
wire _3886_ ;
wire _3466_ ;
wire _3046_ ;
wire _5612_ ;
wire _1952_ ;
wire _1532_ ;
wire _1112_ ;
wire _863_ ;
wire _443_ ;
wire _2737_ ;
wire _2317_ ;
wire _6150_ ;
wire _2490_ ;
wire _2070_ ;
wire _3695_ ;
wire _3275_ ;
wire _5841_ ;
wire _5421_ ;
wire _5001_ ;
wire _919_ ;
wire _6206_ ;
wire _1761_ ;
wire _1341_ ;
wire _672_ ;
wire _252_ ;
wire _2966_ ;
wire _2546_ ;
wire _2126_ ;
wire _3084_ ;
wire _1817_ ;
wire _4289_ ;
wire _5650_ ;
wire _5230_ ;
wire _728_ ;
wire _308_ ;
wire _6015_ ;
wire _1990_ ;
wire _1570_ ;
wire _1150_ ;
wire _481_ ;
wire _2775_ ;
wire _2355_ ;
wire _4921_ ;
wire _4501_ ;
wire _5706_ ;
wire _1626_ ;
wire _1206_ ;
wire _4098_ ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire _6244_ ;
wire _290_ ;
wire _2584_ ;
wire _2164_ ;
wire _3789_ ;
wire _3369_ ;
wire _4730_ ;
wire _4310_ ;
wire _5935_ ;
wire _5515_ ;
wire _1855_ ;
wire _1435_ ;
wire _1015_ ;
wire _766_ ;
wire _346_ ;
wire _6053_ ;
wire _2393_ ;
wire _3598_ ;
wire _3178_ ;
wire _5744_ ;
wire _5324_ ;
wire _6109_ ;
wire _1664_ ;
wire _1244_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire _2869_ ;
wire _2449_ ;
wire _2029_ ;
wire _3810_ ;
wire _6282_ ;
wire [15:0] \Y[3]  ;
wire _5973_ ;
wire _5553_ ;
wire _5133_ ;
wire _6338_ ;
wire _1893_ ;
wire _1473_ ;
wire _1053_ ;
wire _384_ ;
wire _2678_ ;
wire _2258_ ;
wire _6091_ ;
wire _4824_ ;
wire _4404_ ;
wire _5609_ ;
wire _1949_ ;
wire _1529_ ;
wire _1109_ ;
wire _5782_ ;
wire _5362_ ;
wire _6147_ ;
wire _1282_ ;
wire _193_ ;
wire _2487_ ;
wire _2067_ ;
wire _4633_ ;
wire _4213_ ;
wire _5838_ ;
wire _5418_ ;
wire _1758_ ;
wire _1338_ ;
wire _5591_ ;
wire _5171_ ;
wire _669_ ;
wire _249_ ;
wire _3904_ ;
wire [7:0] _6376_ ;
wire _1091_ ;
wire _2296_ ;
wire _4862_ ;
wire _4442_ ;
wire _4022_ ;
wire _5647_ ;
wire _5227_ ;
wire _1987_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _3713_ ;
wire _6185_ ;
wire _4918_ ;
wire _4671_ ;
wire _4251_ ;
wire _5876_ ;
wire _5456_ ;
wire _5036_ ;
wire _1796_ ;
wire _1376_ ;
wire _287_ ;
wire _3942_ ;
wire _3522_ ;
wire _3102_ ;
wire _3_ ;
wire _4727_ ;
wire _4307_ ;
wire _4480_ ;
wire _4060_ ;
wire _5685_ ;
wire _5265_ ;
wire _1185_ ;
wire _3751_ ;
wire _3331_ ;
wire _4956_ ;
wire _4536_ ;
wire _4116_ ;
wire _2602_ ;
wire _5494_ ;
wire _5074_ ;
wire _3807_ ;
wire _6279_ ;
wire _2199_ ;
wire [15:0] _3980_ ;
wire _3560_ ;
wire _3140_ ;
wire _4765_ ;
wire _4345_ ;
wire _44_ ;
wire _2831_ ;
wire _2411_ ;
wire _3616_ ;
wire _6088_ ;
wire _4994_ ;
wire _4574_ ;
wire _4154_ ;
wire _5779_ ;
wire _5359_ ;
wire _6300_ ;
wire _1699_ ;
wire _1279_ ;
wire _2640_ ;
wire _2220_ ;
wire _3845_ ;
wire _3425_ ;
wire _3005_ ;
wire _1911_ ;
wire _4383_ ;
wire _822_ ;
wire _402_ ;
wire _5588_ ;
wire _5168_ ;
wire _82_ ;
wire _1088_ ;
wire _3654_ ;
wire _3234_ ;
wire _4859_ ;
wire _4439_ ;
wire _4019_ ;
wire _5800_ ;
wire _1720_ ;
wire _1300_ ;
wire _4192_ ;
wire _631_ ;
wire _211_ ;
wire _2925_ ;
wire _2505_ ;
wire _5397_ ;
wire _3883_ ;
wire _3463_ ;
wire _3043_ ;
wire _4668_ ;
wire _4248_ ;
wire _860_ ;
wire _440_ ;
wire _2734_ ;
wire _2314_ ;
wire _3939_ ;
wire _3519_ ;
wire _3692_ ;
wire _3272_ ;
wire _4897_ ;
wire _4477_ ;
wire _4057_ ;
wire _916_ ;
wire _6203_ ;
wire _2963_ ;
wire _2543_ ;
wire _2123_ ;
wire _3748_ ;
wire _3328_ ;
wire _3081_ ;
wire _1814_ ;
wire _4286_ ;
wire _725_ ;
wire _305_ ;
wire _6012_ ;
wire _2772_ ;
wire _2352_ ;
wire [15:0] _3977_ ;
wire _3557_ ;
wire _3137_ ;
wire _5703_ ;
wire _1623_ ;
wire _1203_ ;
wire _4095_ ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _2828_ ;
wire _2408_ ;
wire _6241_ ;
wire _2581_ ;
wire _2161_ ;
wire _3786_ ;
wire _3366_ ;
wire _5932_ ;
wire _5512_ ;
wire _1852_ ;
wire _1432_ ;
wire _1012_ ;
wire _763_ ;
wire _343_ ;
wire _2637_ ;
wire _2217_ ;
wire _6050_ ;
wire [15:0] _2390_ ;
wire _3595_ ;
wire _3175_ ;
wire _1908_ ;
wire _5741_ ;
wire _5321_ ;
wire _819_ ;
wire _79_ ;
wire _6106_ ;
wire _1661_ ;
wire _1241_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _2866_ ;
wire _2446_ ;
wire _2026_ ;
wire _1717_ ;
wire _4189_ ;
wire _5970_ ;
wire _5550_ ;
wire _5130_ ;
wire _628_ ;
wire _208_ ;
wire _6335_ ;
wire _1890_ ;
wire _1470_ ;
wire _1050_ ;
wire _381_ ;
wire _2675_ ;
wire _2255_ ;
wire clk_bF$buf40 ;
wire clk_bF$buf41 ;
wire clk_bF$buf42 ;
wire clk_bF$buf43 ;
wire clk_bF$buf44 ;
wire clk_bF$buf45 ;
wire clk_bF$buf46 ;
wire clk_bF$buf47 ;
wire clk_bF$buf48 ;
wire clk_bF$buf49 ;
wire _4821_ ;
wire _4401_ ;
wire _5606_ ;
wire _1946_ ;
wire _1526_ ;
wire _1106_ ;
wire _857_ ;
wire _437_ ;
wire _6144_ ;
wire _190_ ;
wire _2484_ ;
wire _2064_ ;
wire _3689_ ;
wire _3269_ ;
wire _4630_ ;
wire _4210_ ;
wire _5835_ ;
wire _5415_ ;
wire _1755_ ;
wire _1335_ ;
wire _666_ ;
wire _246_ ;
wire _3901_ ;
wire [15:0] _6373_ ;
wire _2293_ ;
wire _3498_ ;
wire _3078_ ;
wire _5644_ ;
wire _5224_ ;
wire _6009_ ;
wire _1984_ ;
wire _1564_ ;
wire _1144_ ;
wire _895_ ;
wire _475_ ;
wire _2769_ ;
wire _2349_ ;
wire _3710_ ;
wire _6182_ ;
wire _4915_ ;
wire [15:0] \u_fir_pe0.rYin  ;
wire _5873_ ;
wire _5453_ ;
wire _5033_ ;
wire _6238_ ;
wire _1793_ ;
wire _1373_ ;
wire _284_ ;
wire _2998_ ;
wire _2578_ ;
wire _2158_ ;
wire _0_ ;
wire _4724_ ;
wire _4304_ ;
wire _5929_ ;
wire _5509_ ;
wire _1849_ ;
wire _1429_ ;
wire _1009_ ;
wire _5682_ ;
wire _5262_ ;
wire _6047_ ;
wire _1182_ ;
wire [7:0] \X[1]  ;
wire [15:0] _2387_ ;
wire _4953_ ;
wire _4533_ ;
wire _4113_ ;
wire _5738_ ;
wire _5318_ ;
wire _1658_ ;
wire _1238_ ;
wire _5491_ ;
wire _5071_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire _3804_ ;
wire _6276_ ;
wire _2196_ ;
wire _4762_ ;
wire _4342_ ;
wire _5967_ ;
wire _5547_ ;
wire _5127_ ;
wire _41_ ;
wire _1887_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _3613_ ;
wire _6085_ ;
wire _4818_ ;
wire _4991_ ;
wire _4571_ ;
wire _4151_ ;
wire _5776_ ;
wire _5356_ ;
wire \X[4]_5_bF$buf1  ;
wire _1696_ ;
wire _1276_ ;
wire _187_ ;
wire _3842_ ;
wire _3422_ ;
wire _3002_ ;
wire _4627_ ;
wire _4207_ ;
wire _4380_ ;
wire _5585_ ;
wire _5165_ ;
wire _1085_ ;
wire _3651_ ;
wire _3231_ ;
wire _4856_ ;
wire _4436_ ;
wire _4016_ ;
wire _2922_ ;
wire _2502_ ;
wire _5394_ ;
wire _3707_ ;
wire _6179_ ;
wire _2099_ ;
wire _3880_ ;
wire _3460_ ;
wire _3040_ ;
wire _4665_ ;
wire _4245_ ;
wire _2731_ ;
wire _2311_ ;
wire [15:0] Yout ;
wire _3936_ ;
wire _3516_ ;
wire _4894_ ;
wire _4474_ ;
wire _4054_ ;
wire _913_ ;
wire _5679_ ;
wire _5259_ ;
wire _6200_ ;
wire _1599_ ;
wire _1179_ ;
wire _2960_ ;
wire _2540_ ;
wire _2120_ ;
wire _3745_ ;
wire _3325_ ;
wire _1811_ ;
wire _4283_ ;
wire _722_ ;
wire _302_ ;
wire _5488_ ;
wire _5068_ ;
wire _3974_ ;
wire _3554_ ;
wire _3134_ ;
wire _4759_ ;
wire _4339_ ;
wire _5700_ ;
wire _38_ ;
wire _1620_ ;
wire _1200_ ;
wire _4092_ ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _2825_ ;
wire _2405_ ;
wire _5297_ ;
wire _3783_ ;
wire _3363_ ;
wire _4988_ ;
wire _4568_ ;
wire _4148_ ;
wire _760_ ;
wire _340_ ;
wire _2634_ ;
wire _2214_ ;
wire _3839_ ;
wire _3419_ ;
wire _3592_ ;
wire _3172_ ;
wire _1905_ ;
wire _4797_ ;
wire _4377_ ;
wire _816_ ;
wire _76_ ;
wire _6103_ ;
wire _2863_ ;
wire _2443_ ;
wire _2023_ ;
wire _3648_ ;
wire _3228_ ;
wire _1714_ ;
wire _4186_ ;
wire _625_ ;
wire _205_ ;
wire _2919_ ;
wire _6332_ ;
wire _2672_ ;
wire _2252_ ;
wire clk_bF$buf10 ;
wire clk_bF$buf11 ;
wire clk_bF$buf12 ;
wire clk_bF$buf13 ;
wire clk_bF$buf14 ;
wire clk_bF$buf15 ;
wire clk_bF$buf16 ;
wire clk_bF$buf17 ;
wire clk_bF$buf18 ;
wire clk_bF$buf19 ;
wire _3877_ ;
wire _3457_ ;
wire _3037_ ;
wire _5603_ ;
wire _1943_ ;
wire _1523_ ;
wire _1103_ ;
wire _854_ ;
wire _434_ ;
wire _2728_ ;
wire _2308_ ;
wire _6141_ ;
wire _2481_ ;
wire _2061_ ;
wire _3686_ ;
wire _3266_ ;
wire _5832_ ;
wire _5412_ ;
wire _1752_ ;
wire _1332_ ;
wire _663_ ;
wire _243_ ;
wire _2957_ ;
wire _2537_ ;
wire _2117_ ;
wire [15:0] _6370_ ;
wire _2290_ ;
wire _3495_ ;
wire _3075_ ;
wire _1808_ ;
wire _5641_ ;
wire _5221_ ;
wire _719_ ;
wire _6006_ ;
wire _1981_ ;
wire _1561_ ;
wire _1141_ ;
wire _892_ ;
wire _472_ ;
wire _2766_ ;
wire _2346_ ;
wire _4912_ ;
wire _1617_ ;
wire _4089_ ;
wire _5870_ ;
wire _5450_ ;
wire _5030_ ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _6235_ ;
wire _1790_ ;
wire _1370_ ;
wire _281_ ;
wire _2995_ ;
wire _2575_ ;
wire _2155_ ;
wire _4721_ ;
wire _4301_ ;
wire _5926_ ;
wire _5506_ ;
wire _1846_ ;
wire _1426_ ;
wire _1006_ ;
wire _757_ ;
wire _337_ ;
wire _6044_ ;
wire [15:0] _2384_ ;
wire _3589_ ;
wire _3169_ ;
wire _4950_ ;
wire _4530_ ;
wire _4110_ ;
wire _5735_ ;
wire _5315_ ;
wire _1655_ ;
wire _1235_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire _3801_ ;
wire _6273_ ;
wire _2193_ ;
wire _3398_ ;
wire _5964_ ;
wire _5544_ ;
wire _5124_ ;
wire _6329_ ;
wire _1884_ ;
wire _1464_ ;
wire _1044_ ;
wire [15:0] _795_ ;
wire _375_ ;
wire _2669_ ;
wire _2249_ ;
wire _3610_ ;
wire _6082_ ;
wire _4815_ ;
wire _5773_ ;
wire _5353_ ;
wire \X[3]_5_bF$buf3  ;
wire _6138_ ;
wire _1693_ ;
wire _1273_ ;
wire _184_ ;
wire _2898_ ;
wire _2478_ ;
wire _2058_ ;
wire _4624_ ;
wire _4204_ ;
wire _5829_ ;
wire _5409_ ;
wire _1749_ ;
wire _1329_ ;
wire _5582_ ;
wire _5162_ ;
wire _6367_ ;
wire _1082_ ;
wire _2287_ ;
wire _4853_ ;
wire _4433_ ;
wire _4013_ ;
wire _5638_ ;
wire _5218_ ;
wire _1978_ ;
wire _1558_ ;
wire _1138_ ;
wire _5391_ ;
wire _889_ ;
wire _469_ ;
wire _3704_ ;
wire _6176_ ;
wire _4909_ ;
wire _2096_ ;
wire _4662_ ;
wire _4242_ ;
wire _5867_ ;
wire _5447_ ;
wire _5027_ ;
wire _1787_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _3933_ ;
wire _3513_ ;
wire _4718_ ;
wire _4891_ ;
wire _4471_ ;
wire _4051_ ;
wire _910_ ;
wire _5676_ ;
wire _5256_ ;
wire _1596_ ;
wire _1176_ ;
wire _3742_ ;
wire _3322_ ;
wire _4947_ ;
wire _4527_ ;
wire _4107_ ;
wire _4280_ ;
wire _5485_ ;
wire _5065_ ;
wire _3971_ ;
wire _3551_ ;
wire _3131_ ;
wire _4756_ ;
wire _4336_ ;
wire _35_ ;
wire _2822_ ;
wire _2402_ ;
wire _5294_ ;
wire _3607_ ;
wire _6079_ ;
wire _3780_ ;
wire _3360_ ;
wire _4985_ ;
wire _4565_ ;
wire _4145_ ;
wire _2631_ ;
wire _2211_ ;
wire [7:0] Xout ;
wire _3836_ ;
wire _3416_ ;
wire _1902_ ;
wire _4794_ ;
wire _4374_ ;
wire _813_ ;
wire _5999_ ;
wire _5579_ ;
wire _5159_ ;
wire _73_ ;
wire _6100_ ;
wire _1499_ ;
wire _1079_ ;
wire _2860_ ;
wire _2440_ ;
wire _2020_ ;
wire _3645_ ;
wire _3225_ ;
wire _1711_ ;
wire _4183_ ;
wire _622_ ;
wire _202_ ;
wire _2916_ ;
wire _5388_ ;
wire _3874_ ;
wire _3454_ ;
wire _3034_ ;
wire _4659_ ;
wire _4239_ ;
wire _5600_ ;
wire _1940_ ;
wire _1520_ ;
wire _1100_ ;
wire _851_ ;
wire _431_ ;
wire _2725_ ;
wire _2305_ ;
wire _5197_ ;
wire _3683_ ;
wire _3263_ ;
wire _4888_ ;
wire _4468_ ;
wire _4048_ ;
wire _907_ ;
wire _660_ ;
wire _240_ ;
wire _2954_ ;
wire _2534_ ;
wire _2114_ ;
wire _3739_ ;
wire _3319_ ;
wire _3492_ ;
wire _3072_ ;
wire _1805_ ;
wire _4697_ ;
wire _4277_ ;
wire _716_ ;
wire _6003_ ;
wire _2763_ ;
wire _2343_ ;
wire _3968_ ;
wire _3548_ ;
wire _3128_ ;
wire _1614_ ;
wire _4086_ ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _2819_ ;
wire _6232_ ;
wire _2992_ ;
wire _2572_ ;
wire _2152_ ;
wire _3777_ ;
wire _3357_ ;
wire _5923_ ;
wire _5503_ ;
wire _1843_ ;
wire _1423_ ;
wire _1003_ ;
wire _754_ ;
wire _334_ ;
wire _2628_ ;
wire _2208_ ;
wire _6041_ ;
wire _2381_ ;
wire _3586_ ;
wire _3166_ ;
wire _5732_ ;
wire _5312_ ;
wire _1652_ ;
wire _1232_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _2857_ ;
wire _2437_ ;
wire _2017_ ;
wire _6270_ ;
wire _2190_ ;
wire _3395_ ;
wire _1708_ ;
wire _5961_ ;
wire _5541_ ;
wire _5121_ ;
wire _619_ ;
wire _6326_ ;
wire _1881_ ;
wire _1461_ ;
wire _1041_ ;
wire [15:0] _792_ ;
wire _372_ ;
wire _2666_ ;
wire _2246_ ;
wire _4812_ ;
wire _1937_ ;
wire _1517_ ;
wire _5770_ ;
wire _5350_ ;
wire _848_ ;
wire _428_ ;
wire \X[3]_5_bF$buf0  ;
wire _6135_ ;
wire _1690_ ;
wire _1270_ ;
wire _181_ ;
wire _2895_ ;
wire _2475_ ;
wire _2055_ ;
wire _4621_ ;
wire _4201_ ;
wire _5826_ ;
wire _5406_ ;
wire _1746_ ;
wire _1326_ ;
wire _657_ ;
wire _237_ ;
wire _6364_ ;
wire _2284_ ;
wire _3489_ ;
wire _3069_ ;
wire _4850_ ;
wire _4430_ ;
wire _4010_ ;
wire _5635_ ;
wire _5215_ ;
wire _1975_ ;
wire _1555_ ;
wire _1135_ ;
wire _886_ ;
wire _466_ ;
wire _3701_ ;
wire _6173_ ;
wire _4906_ ;
wire _2093_ ;
wire _3298_ ;
wire _5864_ ;
wire _5444_ ;
wire _5024_ ;
wire _6229_ ;
wire _1784_ ;
wire _1364_ ;
wire _695_ ;
wire _275_ ;
wire _2989_ ;
wire _2569_ ;
wire _2149_ ;
wire _3930_ ;
wire _3510_ ;
wire _4715_ ;
wire _5673_ ;
wire _5253_ ;
wire _6038_ ;
wire [15:0] _1593_ ;
wire _1173_ ;
wire _2798_ ;
wire _2378_ ;
wire _4944_ ;
wire _4524_ ;
wire _4104_ ;
wire _5729_ ;
wire _5309_ ;
wire _1649_ ;
wire _1229_ ;
wire _5482_ ;
wire _5062_ ;
wire _6267_ ;
wire _2187_ ;
wire _4753_ ;
wire _4333_ ;
wire _5958_ ;
wire _5538_ ;
wire _5118_ ;
wire _32_ ;
wire _1878_ ;
wire _1458_ ;
wire _1038_ ;
wire _5291_ ;
wire [15:0] _789_ ;
wire _369_ ;
wire _3604_ ;
wire _6076_ ;
wire _4809_ ;
wire _4982_ ;
wire _4562_ ;
wire _4142_ ;
wire _5767_ ;
wire _5347_ ;
wire _1687_ ;
wire _1267_ ;
wire _598_ ;
wire _178_ ;
wire _3833_ ;
wire _3413_ ;
wire _4618_ ;
wire _4791_ ;
wire _4371_ ;
wire _810_ ;
wire _5996_ ;
wire [15:0] _5576_ ;
wire _5156_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _3642_ ;
wire _3222_ ;
wire _4847_ ;
wire _4427_ ;
wire _4007_ ;
wire _4180_ ;
wire _2913_ ;
wire _5385_ ;
wire _3871_ ;
wire _3451_ ;
wire _3031_ ;
wire _4656_ ;
wire _4236_ ;
wire _2722_ ;
wire _2302_ ;
wire _5194_ ;
wire _3927_ ;
wire _3507_ ;
wire _3680_ ;
wire _3260_ ;
wire _4885_ ;
wire _4465_ ;
wire _4045_ ;
wire _904_ ;
wire _2951_ ;
wire _2531_ ;
wire _2111_ ;
wire _3736_ ;
wire _3316_ ;
wire _1802_ ;
wire _4694_ ;
wire _4274_ ;
wire _713_ ;
wire _5899_ ;
wire _5479_ ;
wire _5059_ ;
wire _6000_ ;
wire _1399_ ;
wire _2760_ ;
wire _2340_ ;
wire _3965_ ;
wire _3545_ ;
wire _3125_ ;
wire _29_ ;
wire _1611_ ;
wire _4083_ ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _2816_ ;
wire _5288_ ;
wire _3774_ ;
wire _3354_ ;
wire _4979_ ;
wire _4559_ ;
wire _4139_ ;
wire _5920_ ;
wire _5500_ ;
wire _1840_ ;
wire _1420_ ;
wire _1000_ ;
wire _751_ ;
wire _331_ ;
wire _2625_ ;
wire _2205_ ;
wire _5097_ ;
wire _3583_ ;
wire _3163_ ;
wire _4788_ ;
wire _4368_ ;
wire [15:0] \u_fir_pe3.rYin  ;
wire _807_ ;
wire _67_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _2854_ ;
wire _2434_ ;
wire _2014_ ;
wire _3639_ ;
wire _3219_ ;
wire _3392_ ;
wire _1705_ ;
wire _4597_ ;
wire _4177_ ;
wire _616_ ;
wire _6323_ ;
wire _2663_ ;
wire _2243_ ;
wire _3868_ ;
wire _3448_ ;
wire _3028_ ;
wire _1934_ ;
wire _1514_ ;
wire _845_ ;
wire _425_ ;
wire _2719_ ;
wire \X[2]_5_bF$buf2  ;
wire _6132_ ;
wire _2892_ ;
wire _2472_ ;
wire _2052_ ;
wire _3677_ ;
wire _3257_ ;
wire _5823_ ;
wire _5403_ ;
wire _1743_ ;
wire _1323_ ;
wire _654_ ;
wire _234_ ;
wire _2948_ ;
wire _2528_ ;
wire _2108_ ;
wire _6361_ ;
wire _2281_ ;
wire _3486_ ;
wire _3066_ ;
wire _5632_ ;
wire _5212_ ;
wire _1972_ ;
wire _1552_ ;
wire _1132_ ;
wire _883_ ;
wire _463_ ;
wire _2757_ ;
wire _2337_ ;
wire _6170_ ;
wire _4903_ ;
wire _2090_ ;
wire _3295_ ;
wire _1608_ ;
wire _5861_ ;
wire _5441_ ;
wire _5021_ ;
wire _939_ ;
wire _519_ ;
wire _6226_ ;
wire _1781_ ;
wire _1361_ ;
wire _692_ ;
wire _272_ ;
wire _2986_ ;
wire _2566_ ;
wire _2146_ ;
wire _4712_ ;
wire _5917_ ;
wire _1837_ ;
wire _1417_ ;
wire _5670_ ;
wire _5250_ ;
wire _748_ ;
wire _328_ ;
wire _6035_ ;
wire [15:0] _1590_ ;
wire _1170_ ;
wire _2795_ ;
wire _2375_ ;
wire _4941_ ;
wire _4521_ ;
wire _4101_ ;
wire _5726_ ;
wire _5306_ ;
wire _1646_ ;
wire _1226_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire _6264_ ;
wire _2184_ ;
wire _3389_ ;
wire _4750_ ;
wire _4330_ ;
wire _5955_ ;
wire _5535_ ;
wire _5115_ ;
wire _1875_ ;
wire _1455_ ;
wire _1035_ ;
wire _786_ ;
wire _366_ ;
wire _3601_ ;
wire _6073_ ;
wire _4806_ ;
wire _3198_ ;
wire _5764_ ;
wire _5344_ ;
wire _6129_ ;
wire _1684_ ;
wire _1264_ ;
wire _595_ ;
wire _175_ ;
wire _2889_ ;
wire _2469_ ;
wire _2049_ ;
wire _3830_ ;
wire _3410_ ;
wire _4615_ ;
wire [15:0] \Y[5]  ;
wire _5993_ ;
wire [15:0] _5573_ ;
wire _5153_ ;
wire _6358_ ;
wire _1493_ ;
wire _1073_ ;
wire _2698_ ;
wire _2278_ ;
wire _4844_ ;
wire _4424_ ;
wire _4004_ ;
wire _5629_ ;
wire _5209_ ;
wire _1969_ ;
wire _1549_ ;
wire _1129_ ;
wire _2910_ ;
wire _5382_ ;
wire _6167_ ;
wire _2087_ ;
wire _4653_ ;
wire _4233_ ;
wire _5858_ ;
wire _5438_ ;
wire _5018_ ;
wire _1778_ ;
wire _1358_ ;
wire _5191_ ;
wire _689_ ;
wire _269_ ;
wire _3924_ ;
wire _3504_ ;
wire _4709_ ;
wire _4882_ ;
wire _4462_ ;
wire _4042_ ;
wire _901_ ;
wire _5667_ ;
wire _5247_ ;
wire [15:0] _1587_ ;
wire _1167_ ;
wire _498_ ;
wire _3733_ ;
wire _3313_ ;
wire _4938_ ;
wire _4518_ ;
wire _4691_ ;
wire _4271_ ;
wire _710_ ;
wire _5896_ ;
wire _5476_ ;
wire _5056_ ;
wire _1396_ ;
wire _3962_ ;
wire _3542_ ;
wire _3122_ ;
wire _4747_ ;
wire _4327_ ;
wire _26_ ;
wire _4080_ ;
wire _2813_ ;
wire _5285_ ;
wire _3771_ ;
wire _3351_ ;
wire _4976_ ;
wire _4556_ ;
wire _4136_ ;
wire _2622_ ;
wire _2202_ ;
wire _5094_ ;
wire _3827_ ;
wire _3407_ ;
wire _6299_ ;
wire _3580_ ;
wire _3160_ ;
wire _4785_ ;
wire _4365_ ;
wire _804_ ;
wire _64_ ;
wire _2851_ ;
wire _2431_ ;
wire _2011_ ;
wire _3636_ ;
wire _3216_ ;
wire _1702_ ;
wire _4594_ ;
wire _4174_ ;
wire _613_ ;
wire _2907_ ;
wire _5799_ ;
wire _5379_ ;
wire _6320_ ;
wire _1299_ ;
wire _2660_ ;
wire _2240_ ;
wire _3865_ ;
wire _3445_ ;
wire _3025_ ;
wire _1931_ ;
wire _1511_ ;
wire _842_ ;
wire _422_ ;
wire _2716_ ;
wire _5188_ ;
wire _3674_ ;
wire _3254_ ;
wire _4879_ ;
wire _4459_ ;
wire _4039_ ;
wire _5820_ ;
wire _5400_ ;
wire _1740_ ;
wire _1320_ ;
wire _651_ ;
wire _231_ ;
wire _2945_ ;
wire _2525_ ;
wire _2105_ ;
wire _3483_ ;
wire _3063_ ;
wire _4688_ ;
wire _4268_ ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _2754_ ;
wire _2334_ ;
wire _3959_ ;
wire _3539_ ;
wire _3119_ ;
wire _4900_ ;
wire _3292_ ;
wire _1605_ ;
wire _4497_ ;
wire _4077_ ;
wire _936_ ;
wire _516_ ;
wire _6223_ ;
wire _2983_ ;
wire _2563_ ;
wire _2143_ ;
wire _3768_ ;
wire _3348_ ;
wire _5914_ ;
wire _1834_ ;
wire _1414_ ;
wire _745_ ;
wire _325_ ;
wire _2619_ ;
wire _6032_ ;
wire _2792_ ;
wire _2372_ ;
wire _3997_ ;
wire _3577_ ;
wire _3157_ ;
wire _5723_ ;
wire _5303_ ;
wire _1643_ ;
wire _1223_ ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire _2848_ ;
wire _2428_ ;
wire _2008_ ;
wire _6261_ ;
wire _2181_ ;
wire _3386_ ;
wire _5952_ ;
wire _5532_ ;
wire _5112_ ;
wire _6317_ ;
wire _1872_ ;
wire _1452_ ;
wire _1032_ ;
wire _783_ ;
wire _363_ ;
wire _2657_ ;
wire _2237_ ;
wire _6070_ ;
wire _4803_ ;
wire _3195_ ;
wire _1928_ ;
wire _1508_ ;
wire _5761_ ;
wire _5341_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _6126_ ;
wire _1681_ ;
wire _1261_ ;
wire _592_ ;
wire _172_ ;
wire _2886_ ;
wire _2466_ ;
wire _2046_ ;
wire _4612_ ;
wire _5817_ ;
wire _1737_ ;
wire _1317_ ;
wire _5990_ ;
wire _5570_ ;
wire _5150_ ;
wire _648_ ;
wire _228_ ;
wire _6355_ ;
wire _1490_ ;
wire _1070_ ;
wire _2695_ ;
wire _2275_ ;
wire _4841_ ;
wire _4421_ ;
wire _4001_ ;
wire _5626_ ;
wire _5206_ ;
wire _1966_ ;
wire _1546_ ;
wire _1126_ ;
wire _877_ ;
wire _457_ ;
wire _6164_ ;
wire _2084_ ;
wire _3289_ ;
wire _4650_ ;
wire _4230_ ;
wire _5855_ ;
wire _5435_ ;
wire _5015_ ;
wire _1775_ ;
wire _1355_ ;
wire _686_ ;
wire _266_ ;
wire _3921_ ;
wire _3501_ ;
wire _4706_ ;
wire _3098_ ;
wire _5664_ ;
wire _5244_ ;
wire _6029_ ;
wire _1584_ ;
wire _1164_ ;
wire _495_ ;
wire _2789_ ;
wire _2369_ ;
wire _3730_ ;
wire _3310_ ;
wire _4935_ ;
wire _4515_ ;
wire _5893_ ;
wire _5473_ ;
wire _5053_ ;
wire [15:0] \u_fir_pe1.mul  ;
wire _6258_ ;
wire _1393_ ;
wire _2598_ ;
wire _2178_ ;
wire _4744_ ;
wire _4324_ ;
wire \X[7]_5_bF$buf3  ;
wire _5949_ ;
wire _5529_ ;
wire _5109_ ;
wire _23_ ;
wire _1869_ ;
wire _1449_ ;
wire _1029_ ;
wire _2810_ ;
wire _5282_ ;
wire _6067_ ;
wire [7:0] \X[3]  ;
wire _4973_ ;
wire _4553_ ;
wire _4133_ ;
wire _5758_ ;
wire _5338_ ;
wire _1678_ ;
wire _1258_ ;
wire _5091_ ;
wire _589_ ;
wire _169_ ;
wire _3824_ ;
wire _3404_ ;
wire _6296_ ;
wire _4609_ ;
wire _4782_ ;
wire _4362_ ;
wire _801_ ;
wire _5987_ ;
wire _5567_ ;
wire _5147_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _398_ ;
wire _3633_ ;
wire _3213_ ;
wire _4838_ ;
wire _4418_ ;
wire _4591_ ;
wire _4171_ ;
wire _610_ ;
wire _2904_ ;
wire _5796_ ;
wire _5376_ ;
wire _1296_ ;
wire _3862_ ;
wire _3442_ ;
wire _3022_ ;
wire _4647_ ;
wire _4227_ ;
wire _2713_ ;
wire _5185_ ;
wire [15:0] \u_fir_pe3.mul  ;
wire \X[1]_5_bF$buf1  ;
wire _3918_ ;
wire _3671_ ;
wire _3251_ ;
wire _4876_ ;
wire _4456_ ;
wire _4036_ ;
wire _2942_ ;
wire _2522_ ;
wire _2102_ ;
wire _3727_ ;
wire _3307_ ;
wire _6199_ ;
wire _3480_ ;
wire _3060_ ;
wire _4685_ ;
wire _4265_ ;
wire _704_ ;
wire _2751_ ;
wire _2331_ ;
wire _3956_ ;
wire _3536_ ;
wire _3116_ ;
wire _1602_ ;
wire _4494_ ;
wire _4074_ ;
wire _933_ ;
wire _513_ ;
wire _2807_ ;
wire _5699_ ;
wire _5279_ ;
wire _6220_ ;
wire _1199_ ;
wire _2980_ ;
wire _2560_ ;
wire _2140_ ;
wire _3765_ ;
wire _3345_ ;
wire _5911_ ;
wire _1831_ ;
wire _1411_ ;
wire _742_ ;
wire _322_ ;
wire _2616_ ;
wire _5088_ ;
wire _3994_ ;
wire _3574_ ;
wire _3154_ ;
wire [15:0] _4779_ ;
wire _4359_ ;
wire _5720_ ;
wire _5300_ ;
wire _58_ ;
wire _1640_ ;
wire _1220_ ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _2845_ ;
wire _2425_ ;
wire _2005_ ;
wire _3383_ ;
wire _4588_ ;
wire _4168_ ;
wire _607_ ;
wire _6314_ ;
wire _780_ ;
wire _360_ ;
wire _2654_ ;
wire _2234_ ;
wire _3859_ ;
wire _3439_ ;
wire _3019_ ;
wire _4800_ ;
wire _3192_ ;
wire _1925_ ;
wire _1505_ ;
wire _4397_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _6123_ ;
wire _2883_ ;
wire _2463_ ;
wire _2043_ ;
wire _3668_ ;
wire _3248_ ;
wire _5814_ ;
wire _1734_ ;
wire _1314_ ;
wire _645_ ;
wire _225_ ;
wire _2939_ ;
wire _2519_ ;
wire _6352_ ;
wire _2692_ ;
wire _2272_ ;
wire _3897_ ;
wire _3477_ ;
wire _3057_ ;
wire _5623_ ;
wire _5203_ ;
wire _1963_ ;
wire _1543_ ;
wire _1123_ ;
wire _874_ ;
wire _454_ ;
wire _2748_ ;
wire _2328_ ;
wire _6161_ ;
wire _2081_ ;
wire _3286_ ;
wire _5852_ ;
wire _5432_ ;
wire _5012_ ;
wire _6217_ ;
wire _1772_ ;
wire _1352_ ;
wire _683_ ;
wire _263_ ;
wire _2977_ ;
wire _2557_ ;
wire _2137_ ;
wire _4703_ ;
wire _5908_ ;
wire _3095_ ;
wire _1828_ ;
wire _1408_ ;
wire _5661_ ;
wire _5241_ ;
wire _739_ ;
wire _319_ ;
wire _6026_ ;
wire _1581_ ;
wire _1161_ ;
wire _492_ ;
wire _2786_ ;
wire _2366_ ;
wire _4932_ ;
wire _4512_ ;
wire _5717_ ;
wire _1637_ ;
wire _1217_ ;
wire _5890_ ;
wire _5470_ ;
wire _5050_ ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _6255_ ;
wire _1390_ ;
wire _2595_ ;
wire _2175_ ;
wire _4741_ ;
wire _4321_ ;
wire \X[7]_5_bF$buf0  ;
wire _5946_ ;
wire _5526_ ;
wire _5106_ ;
wire _20_ ;
wire _1866_ ;
wire _1446_ ;
wire _1026_ ;
wire _777_ ;
wire _357_ ;
wire _6064_ ;
wire _3189_ ;
wire _4970_ ;
wire _4550_ ;
wire _4130_ ;
wire _5755_ ;
wire _5335_ ;
wire _1675_ ;
wire _1255_ ;
wire _586_ ;
wire _166_ ;
wire _3821_ ;
wire _3401_ ;
wire _6293_ ;
wire _4606_ ;
wire _5984_ ;
wire _5564_ ;
wire _5144_ ;
wire _6349_ ;
wire _1484_ ;
wire _1064_ ;
wire _395_ ;
wire _2689_ ;
wire _2269_ ;
wire _3630_ ;
wire _3210_ ;
wire _4835_ ;
wire _4415_ ;
wire _2901_ ;
wire _5793_ ;
wire _5373_ ;
wire _6158_ ;
wire _1293_ ;
wire _2498_ ;
wire _2078_ ;
wire _4644_ ;
wire _4224_ ;
wire [15:0] \u_fir_pe6.rYin  ;
wire _5849_ ;
wire _5429_ ;
wire _5009_ ;
wire _1769_ ;
wire _1349_ ;
wire _2710_ ;
wire _5182_ ;
wire _3915_ ;
wire _4873_ ;
wire _4453_ ;
wire _4033_ ;
wire _5658_ ;
wire _5238_ ;
wire _1998_ ;
wire _1578_ ;
wire _1158_ ;
wire _489_ ;
wire _3724_ ;
wire _3304_ ;
wire _6196_ ;
wire _4929_ ;
wire _4509_ ;
wire _4682_ ;
wire _4262_ ;
wire _701_ ;
wire _5887_ ;
wire _5467_ ;
wire _5047_ ;
wire _1387_ ;
wire _298_ ;
wire _3953_ ;
wire _3533_ ;
wire _3113_ ;
wire _4738_ ;
wire _4318_ ;
wire _17_ ;
wire _4491_ ;
wire _4071_ ;
wire _930_ ;
wire _510_ ;
wire _2804_ ;
wire _5696_ ;
wire _5276_ ;
wire _1196_ ;
wire _3762_ ;
wire _3342_ ;
wire _4967_ ;
wire _4547_ ;
wire _4127_ ;
wire _2613_ ;
wire _5085_ ;
wire _3818_ ;
wire _3991_ ;
wire _3571_ ;
wire _3151_ ;
wire [15:0] _4776_ ;
wire _4356_ ;
wire _55_ ;
wire _2842_ ;
wire _2422_ ;
wire _2002_ ;
wire _3627_ ;
wire _3207_ ;
wire _6099_ ;
wire _3380_ ;
wire _4585_ ;
wire _4165_ ;
wire _604_ ;
wire _6311_ ;
wire _2651_ ;
wire _2231_ ;
wire _3856_ ;
wire _3436_ ;
wire _3016_ ;
wire _1922_ ;
wire _1502_ ;
wire _4394_ ;
wire _833_ ;
wire _413_ ;
wire _2707_ ;
wire _5599_ ;
wire _5179_ ;
wire _93_ ;
wire _6120_ ;
wire _1099_ ;
wire _2880_ ;
wire _2460_ ;
wire _2040_ ;
wire _3665_ ;
wire _3245_ ;
wire _5811_ ;
wire _1731_ ;
wire _1311_ ;
wire _642_ ;
wire _222_ ;
wire _2936_ ;
wire _2516_ ;
wire _3894_ ;
wire _3474_ ;
wire _3054_ ;
wire _4679_ ;
wire _4259_ ;
wire _5620_ ;
wire _5200_ ;
wire _1960_ ;
wire _1540_ ;
wire _1120_ ;
wire _871_ ;
wire _451_ ;
wire _2745_ ;
wire _2325_ ;
wire _3283_ ;
wire _4488_ ;
wire _4068_ ;
wire _927_ ;
wire _507_ ;
wire _6214_ ;
wire _680_ ;
wire _260_ ;
wire _2974_ ;
wire _2554_ ;
wire _2134_ ;
wire _3759_ ;
wire _3339_ ;
wire _4700_ ;
wire _5905_ ;
wire _3092_ ;
wire _1825_ ;
wire _1405_ ;
wire _4297_ ;
wire _736_ ;
wire _316_ ;
wire _6023_ ;
wire _2783_ ;
wire _2363_ ;
wire _3988_ ;
wire _3568_ ;
wire _3148_ ;
wire _5714_ ;
wire _1634_ ;
wire _1214_ ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _2839_ ;
wire _2419_ ;
wire _6252_ ;
wire _2592_ ;
wire _2172_ ;
wire _3797_ ;
wire _3377_ ;
wire _5943_ ;
wire _5523_ ;
wire _5103_ ;
wire \X[6]_5_bF$buf2  ;
wire _6308_ ;
wire _1863_ ;
wire _1443_ ;
wire _1023_ ;
wire _774_ ;
wire _354_ ;
wire _2648_ ;
wire _2228_ ;
wire _6061_ ;
wire [15:0] _3186_ ;
wire _1919_ ;
wire _5752_ ;
wire _5332_ ;
wire _6117_ ;
wire _1672_ ;
wire _1252_ ;
wire _583_ ;
wire _163_ ;
wire _2877_ ;
wire _2457_ ;
wire _2037_ ;
wire _6290_ ;
wire _4603_ ;
wire _5808_ ;
wire _1728_ ;
wire _1308_ ;
wire _5981_ ;
wire _5561_ ;
wire _5141_ ;
wire _639_ ;
wire _219_ ;
wire _6346_ ;
wire _1481_ ;
wire _1061_ ;
wire _392_ ;
wire _2686_ ;
wire _2266_ ;
wire _4832_ ;
wire _4412_ ;
wire _5617_ ;
wire _1957_ ;
wire _1537_ ;
wire _1117_ ;
wire _5790_ ;
wire _5370_ ;
wire _868_ ;
wire _448_ ;
wire _6155_ ;
wire _1290_ ;
wire _2495_ ;
wire _2075_ ;
wire _4641_ ;
wire _4221_ ;
wire _5846_ ;
wire _5426_ ;
wire _5006_ ;
wire _1766_ ;
wire _1346_ ;
wire _677_ ;
wire _257_ ;
wire _3912_ ;
wire _3089_ ;
wire _4870_ ;
wire _4450_ ;
wire _4030_ ;
wire _5655_ ;
wire _5235_ ;
wire _1995_ ;
wire _1575_ ;
wire _1155_ ;
wire _486_ ;
wire _3721_ ;
wire _3301_ ;
wire _6193_ ;
wire _4926_ ;
wire _4506_ ;
wire _5884_ ;
wire _5464_ ;
wire _5044_ ;
wire _6249_ ;
wire _1384_ ;
wire _295_ ;
wire _2589_ ;
wire _2169_ ;
wire _3950_ ;
wire _3530_ ;
wire _3110_ ;
wire _4735_ ;
wire _4315_ ;
wire _14_ ;
wire _2801_ ;
wire _5693_ ;
wire _5273_ ;
wire _6058_ ;
wire _1193_ ;
wire _2398_ ;
wire _4964_ ;
wire _4544_ ;
wire _4124_ ;
wire _5749_ ;
wire _5329_ ;
wire _1669_ ;
wire _1249_ ;
wire _2610_ ;
wire _5082_ ;
wire _3815_ ;
wire _6287_ ;
wire _4773_ ;
wire _4353_ ;
wire _5978_ ;
wire _5558_ ;
wire _5138_ ;
wire _52_ ;
wire _1898_ ;
wire _1478_ ;
wire _1058_ ;
wire _389_ ;
wire _3624_ ;
wire _3204_ ;
wire _6096_ ;
wire _4829_ ;
wire _4409_ ;
wire _4582_ ;
wire _4162_ ;
wire _601_ ;
wire _5787_ ;
wire _5367_ ;
wire _1287_ ;
wire _198_ ;
wire _3853_ ;
wire _3433_ ;
wire _3013_ ;
wire _4638_ ;
wire _4218_ ;
wire _4391_ ;
wire _830_ ;
wire _410_ ;
wire _2704_ ;
wire _5596_ ;
wire _5176_ ;
wire _90_ ;
wire _3909_ ;
wire _1096_ ;
wire _3662_ ;
wire _3242_ ;
wire _4867_ ;
wire _4447_ ;
wire _4027_ ;
wire _2933_ ;
wire _2513_ ;
wire _3718_ ;
wire _3891_ ;
wire _3471_ ;
wire _3051_ ;
wire _4676_ ;
wire _4256_ ;
wire _2742_ ;
wire _2322_ ;
wire _3947_ ;
wire _3527_ ;
wire _3107_ ;
wire _8_ ;
wire _3280_ ;
wire _4485_ ;
wire _4065_ ;
wire _924_ ;
wire _504_ ;
wire _6211_ ;
wire _2971_ ;
wire _2551_ ;
wire _2131_ ;
wire _3756_ ;
wire _3336_ ;
wire _5902_ ;
wire _1822_ ;
wire _1402_ ;
wire _4294_ ;
wire _733_ ;
wire _313_ ;
wire _2607_ ;
wire _5499_ ;
wire _5079_ ;
wire _6020_ ;
wire _2780_ ;
wire _2360_ ;
wire _3985_ ;
wire _3565_ ;
wire _3145_ ;
wire _5711_ ;
wire _49_ ;
wire _1631_ ;
wire _1211_ ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _2836_ ;
wire _2416_ ;
wire _3794_ ;
wire _3374_ ;
wire _4999_ ;
wire _4579_ ;
wire _4159_ ;
wire _5940_ ;
wire _5520_ ;
wire _5100_ ;
wire _6305_ ;
wire _1860_ ;
wire _1440_ ;
wire _1020_ ;
wire _771_ ;
wire _351_ ;
wire _2645_ ;
wire _2225_ ;
wire [15:0] _3183_ ;
wire _1916_ ;
wire _4388_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _6114_ ;
wire _580_ ;
wire _160_ ;
wire _2874_ ;
wire _2454_ ;
wire _2034_ ;
wire _3659_ ;
wire _3239_ ;
wire _4600_ ;
wire _5805_ ;
wire _1725_ ;
wire _1305_ ;
wire _4197_ ;
wire _636_ ;
wire _216_ ;
wire _6343_ ;
wire _2683_ ;
wire _2263_ ;
wire _3888_ ;
wire _3468_ ;
wire _3048_ ;
wire _5614_ ;
wire _1954_ ;
wire _1534_ ;
wire _1114_ ;
wire _865_ ;
wire _445_ ;
wire _2739_ ;
wire _2319_ ;
wire _6152_ ;
wire _2492_ ;
wire _2072_ ;
wire _3697_ ;
wire _3277_ ;
wire _5843_ ;
wire _5423_ ;
wire _5003_ ;
wire _6208_ ;
wire _1763_ ;
wire _1343_ ;
wire _674_ ;
wire _254_ ;
wire _2968_ ;
wire _2548_ ;
wire _2128_ ;
wire _3086_ ;
wire _1819_ ;
wire _5652_ ;
wire _5232_ ;
wire _6017_ ;
wire _1992_ ;
wire _1572_ ;
wire _1152_ ;
wire _483_ ;
wire _2777_ ;
wire _2357_ ;
wire _6190_ ;
wire _4923_ ;
wire _4503_ ;
wire _5708_ ;
wire _1628_ ;
wire _1208_ ;
wire _5881_ ;
wire _5461_ ;
wire _5041_ ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _6246_ ;
wire _1381_ ;
wire _292_ ;
wire _2586_ ;
wire _2166_ ;
wire _4732_ ;
wire _4312_ ;
wire _5937_ ;
wire _5517_ ;
wire _11_ ;
wire _1857_ ;
wire _1437_ ;
wire _1017_ ;
wire _5690_ ;
wire _5270_ ;
wire _768_ ;
wire _348_ ;
wire _6055_ ;
wire _1190_ ;
wire _2395_ ;
wire _4961_ ;
wire _4541_ ;
wire _4121_ ;
wire _5746_ ;
wire _5326_ ;
wire _1666_ ;
wire _1246_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _3812_ ;
wire _6284_ ;
wire _4770_ ;
wire _4350_ ;
wire _5975_ ;
wire _5555_ ;
wire _5135_ ;
wire _1895_ ;
wire _1475_ ;
wire _1055_ ;
wire _386_ ;
wire _3621_ ;
wire _3201_ ;
wire _6093_ ;
wire _4826_ ;
wire _4406_ ;
wire _5784_ ;
wire _5364_ ;
wire _6149_ ;
wire _1284_ ;
wire _195_ ;
wire _2489_ ;
wire _2069_ ;
wire _3850_ ;
wire _3430_ ;
wire _3010_ ;
wire _4635_ ;
wire _4215_ ;
wire [15:0] \Y[7]  ;
wire _2701_ ;
wire _5593_ ;
wire _5173_ ;
wire _3906_ ;
wire _1093_ ;
wire _2298_ ;
wire _4864_ ;
wire _4444_ ;
wire _4024_ ;
wire _5649_ ;
wire _5229_ ;
wire _1989_ ;
wire _1569_ ;
wire _1149_ ;
wire _2930_ ;
wire _2510_ ;
wire _3715_ ;
wire _6187_ ;
wire _4673_ ;
wire _4253_ ;
wire _5878_ ;
wire _5458_ ;
wire _5038_ ;
wire _1798_ ;
wire _1378_ ;
wire _289_ ;
wire _3944_ ;
wire _3524_ ;
wire _3104_ ;
wire _5_ ;
wire _4729_ ;
wire _4309_ ;
wire _4482_ ;
wire _4062_ ;
wire _921_ ;
wire _501_ ;
wire _5687_ ;
wire _5267_ ;
wire _1187_ ;
wire _3753_ ;
wire _3333_ ;
wire _4958_ ;
wire _4538_ ;
wire _4118_ ;
wire _4291_ ;
wire _730_ ;
wire _310_ ;
wire _2604_ ;
wire _5496_ ;
wire _5076_ ;
wire _3809_ ;
wire [15:0] _3982_ ;
wire _3562_ ;
wire _3142_ ;
wire _4767_ ;
wire _4347_ ;
wire _46_ ;
wire _2833_ ;
wire _2413_ ;
wire _3618_ ;
wire _3791_ ;
wire _3371_ ;
wire _4996_ ;
wire _4576_ ;
wire _4156_ ;
wire \X[5]_5_bF$buf1  ;
wire _6302_ ;
wire _2642_ ;
wire _2222_ ;
wire _3847_ ;
wire _3427_ ;
wire _3007_ ;
wire [15:0] _3180_ ;
wire _1913_ ;
wire _4385_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _6111_ ;
wire _2871_ ;
wire _2451_ ;
wire _2031_ ;
wire _3656_ ;
wire _3236_ ;
wire _5802_ ;
wire _1722_ ;
wire _1302_ ;
wire _4194_ ;
wire _633_ ;
wire _213_ ;
wire _2927_ ;
wire _2507_ ;
wire _5399_ ;
wire _6340_ ;
wire _2680_ ;
wire _2260_ ;
wire _3885_ ;
wire _3465_ ;
wire _3045_ ;
wire _5611_ ;
wire _1951_ ;
wire _1531_ ;
wire _1111_ ;
wire _862_ ;
wire _442_ ;
wire _2736_ ;
wire _2316_ ;
wire _3694_ ;
wire _3274_ ;
wire _4899_ ;
wire _4479_ ;
wire _4059_ ;
wire _5840_ ;
wire _5420_ ;
wire _5000_ ;
wire _918_ ;
wire _6205_ ;
wire _1760_ ;
wire _1340_ ;
wire _671_ ;
wire _251_ ;
wire _2965_ ;
wire _2545_ ;
wire _2125_ ;
wire _3083_ ;
wire _1816_ ;
wire _4288_ ;
wire _727_ ;
wire _307_ ;
wire _6014_ ;
wire _480_ ;
wire _2774_ ;
wire _2354_ ;
wire [15:0] _3979_ ;
wire _3559_ ;
wire _3139_ ;
wire _4920_ ;
wire _4500_ ;
wire _5705_ ;
wire _1625_ ;
wire _1205_ ;
wire _4097_ ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _6243_ ;
wire _2583_ ;
wire _2163_ ;
wire _3788_ ;
wire _3368_ ;
wire _5934_ ;
wire _5514_ ;
wire _1854_ ;
wire _1434_ ;
wire _1014_ ;
wire _765_ ;
wire _345_ ;
wire _2639_ ;
wire _2219_ ;
wire _6052_ ;
wire _2392_ ;
wire _3597_ ;
wire _3177_ ;
wire _5743_ ;
wire _5323_ ;
wire _6108_ ;
wire _1663_ ;
wire _1243_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _2868_ ;
wire _2448_ ;
wire _2028_ ;
wire _6281_ ;
wire _1719_ ;
wire _5972_ ;
wire _5552_ ;
wire _5132_ ;
wire _6337_ ;
wire _1892_ ;
wire _1472_ ;
wire _1052_ ;
wire _383_ ;
wire _2677_ ;
wire _2257_ ;
wire _6090_ ;
wire _4823_ ;
wire _4403_ ;
wire _5608_ ;
wire _1948_ ;
wire _1528_ ;
wire _1108_ ;
wire _5781_ ;
wire _5361_ ;
wire _859_ ;
wire _439_ ;
wire _6146_ ;
wire _1281_ ;
wire _192_ ;
wire _2486_ ;
wire _2066_ ;
wire _4632_ ;
wire _4212_ ;
wire _5837_ ;
wire _5417_ ;
wire _1757_ ;
wire _1337_ ;
wire _5590_ ;
wire _5170_ ;
wire _668_ ;
wire _248_ ;
wire _3903_ ;
wire [15:0] _6375_ ;
wire _1090_ ;
wire _2295_ ;
wire _4861_ ;
wire _4441_ ;
wire _4021_ ;
wire _5646_ ;
wire _5226_ ;
wire _1986_ ;
wire _1566_ ;
wire _1146_ ;
wire _897_ ;
wire _477_ ;
wire _3712_ ;
wire _6184_ ;
wire _4917_ ;
wire _4670_ ;
wire _4250_ ;
wire _5875_ ;
wire _5455_ ;
wire _5035_ ;
wire _1795_ ;
wire _1375_ ;
wire _286_ ;
wire _3941_ ;
wire _3521_ ;
wire _3101_ ;
wire _2_ ;
wire _4726_ ;
wire _4306_ ;
wire _5684_ ;
wire _5264_ ;
wire _6049_ ;
wire _1184_ ;
wire [15:0] _2389_ ;
wire _3750_ ;
wire _3330_ ;
wire _4955_ ;
wire _4535_ ;
wire _4115_ ;
wire _2601_ ;
wire _5493_ ;
wire _5073_ ;
wire _3806_ ;
wire _6278_ ;
wire _2198_ ;
wire _4764_ ;
wire _4344_ ;
wire _5969_ ;
wire _5549_ ;
wire _5129_ ;
wire _43_ ;
wire _1889_ ;
wire _1469_ ;
wire _1049_ ;
wire _2830_ ;
wire _2410_ ;
wire _3615_ ;
wire _6087_ ;
wire [7:0] \X[5]  ;
wire _4993_ ;
wire _4573_ ;
wire _4153_ ;
wire _5778_ ;
wire _5358_ ;
wire \X[4]_5_bF$buf3  ;
wire _1698_ ;
wire _1278_ ;
wire _189_ ;
wire _3844_ ;
wire _3424_ ;
wire _3004_ ;
wire _4629_ ;
wire _4209_ ;
wire _1910_ ;
wire _4382_ ;
wire _821_ ;
wire _401_ ;
wire _5587_ ;
wire _5167_ ;
wire _81_ ;
wire _1087_ ;
wire _3653_ ;
wire _3233_ ;
wire _4858_ ;
wire _4438_ ;
wire _4018_ ;
wire _4191_ ;
wire _630_ ;
wire _210_ ;
wire _2924_ ;
wire _2504_ ;
wire _5396_ ;
wire _3709_ ;
wire _3882_ ;
wire _3462_ ;
wire _3042_ ;
wire _4667_ ;
wire _4247_ ;
wire _2733_ ;
wire _2313_ ;
wire _3938_ ;
wire _3518_ ;
wire _3691_ ;
wire _3271_ ;
wire _4896_ ;
wire _4476_ ;
wire _4056_ ;
wire _915_ ;
wire _6202_ ;
wire _2962_ ;
wire _2542_ ;
wire _2122_ ;
wire _3747_ ;
wire _3327_ ;
wire _3080_ ;
wire _1813_ ;
wire _4285_ ;
wire _724_ ;
wire _304_ ;
wire _6011_ ;
wire _2771_ ;
wire _2351_ ;
wire _3976_ ;
wire _3556_ ;
wire _3136_ ;
wire _5702_ ;
wire _1622_ ;
wire _1202_ ;
wire _4094_ ;
wire _953_ ;
wire _533_ ;
wire _113_ ;
wire _2827_ ;
wire _2407_ ;
wire _5299_ ;
wire _6240_ ;
wire _2580_ ;
wire _2160_ ;
wire _3785_ ;
wire _3365_ ;
wire _5931_ ;
wire _5511_ ;
wire _1851_ ;
wire _1431_ ;
wire _1011_ ;
wire _762_ ;
wire _342_ ;
wire _2636_ ;
wire _2216_ ;
wire _3594_ ;
wire _3174_ ;
wire _1907_ ;
wire _4799_ ;
wire _4379_ ;
wire _5740_ ;
wire _5320_ ;
wire _818_ ;
wire _78_ ;
wire _6105_ ;
wire _1660_ ;
wire _1240_ ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _2865_ ;
wire _2445_ ;
wire _2025_ ;
wire _1716_ ;
wire _4188_ ;
wire _627_ ;
wire _207_ ;
wire _6334_ ;
wire _380_ ;
wire _2674_ ;
wire _2254_ ;
wire clk_bF$buf30 ;
wire clk_bF$buf31 ;
wire clk_bF$buf32 ;
wire clk_bF$buf33 ;
wire clk_bF$buf34 ;
wire clk_bF$buf35 ;
wire clk_bF$buf36 ;
wire clk_bF$buf37 ;
wire clk_bF$buf38 ;
wire clk_bF$buf39 ;
wire _3879_ ;
wire _3459_ ;
wire _3039_ ;
wire _4820_ ;
wire _4400_ ;
wire _5605_ ;
wire _1945_ ;
wire _1525_ ;
wire _1105_ ;
wire _856_ ;
wire _436_ ;
wire _6143_ ;
wire _2483_ ;
wire _2063_ ;
wire _3688_ ;
wire _3268_ ;
wire _5834_ ;
wire _5414_ ;
wire _1754_ ;
wire _1334_ ;
wire [7:0] Xin ;
wire _665_ ;
wire _245_ ;
wire _2959_ ;
wire _2539_ ;
wire _2119_ ;
wire _3900_ ;
wire [15:0] _6372_ ;
wire _2292_ ;
wire _3497_ ;
wire _3077_ ;
wire _5643_ ;
wire _5223_ ;
wire _6008_ ;
wire _1983_ ;
wire _1563_ ;
wire _1143_ ;
wire _894_ ;
wire _474_ ;
wire _2768_ ;
wire _2348_ ;
wire _6181_ ;
wire _4914_ ;
wire _1619_ ;
wire _5872_ ;
wire _5452_ ;
wire _5032_ ;
wire _6237_ ;
wire _1792_ ;
wire _1372_ ;
wire _283_ ;
wire _2997_ ;
wire _2577_ ;
wire _2157_ ;
wire _4723_ ;
wire _4303_ ;
wire _5928_ ;
wire _5508_ ;
wire _1848_ ;
wire _1428_ ;
wire _1008_ ;
wire _5681_ ;
wire _5261_ ;
wire _759_ ;
wire _339_ ;
wire _6046_ ;
wire _1181_ ;
wire [15:0] _2386_ ;
wire _4952_ ;
wire _4532_ ;
wire _4112_ ;
wire _5737_ ;
wire _5317_ ;
wire _1657_ ;
wire _1237_ ;
wire _5490_ ;
wire _5070_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _3803_ ;
wire _6275_ ;
wire _2195_ ;
wire _4761_ ;
wire _4341_ ;
wire _5966_ ;
wire _5546_ ;
wire _5126_ ;
wire _40_ ;
wire _1886_ ;
wire _1466_ ;
wire _1046_ ;
wire _797_ ;
wire _377_ ;
wire _3612_ ;
wire _6084_ ;
wire _4817_ ;
wire _4990_ ;
wire _4570_ ;
wire _4150_ ;
wire _5775_ ;
wire _5355_ ;
wire \X[4]_5_bF$buf0  ;
wire _1695_ ;
wire _1275_ ;
wire _186_ ;
wire _3841_ ;
wire _3421_ ;
wire _3001_ ;
wire _4626_ ;
wire _4206_ ;
wire _5584_ ;
wire _5164_ ;
wire [15:0] _6369_ ;
wire _1084_ ;
wire _2289_ ;
wire _3650_ ;
wire _3230_ ;
wire _4855_ ;
wire _4435_ ;
wire _4015_ ;
wire _2921_ ;
wire _2501_ ;
wire _5393_ ;
wire _3706_ ;
wire _6178_ ;
wire _2098_ ;
wire _4664_ ;
wire _4244_ ;
wire _5869_ ;
wire _5449_ ;
wire _5029_ ;
wire _1789_ ;
wire _1369_ ;
wire _2730_ ;
wire _2310_ ;
wire _3935_ ;
wire _3515_ ;
wire _4893_ ;
wire _4473_ ;
wire _4053_ ;
wire _912_ ;
wire _5678_ ;
wire _5258_ ;
wire _1598_ ;
wire _1178_ ;
wire _3744_ ;
wire _3324_ ;
wire _4949_ ;
wire _4529_ ;
wire _4109_ ;
wire _1810_ ;
wire _4282_ ;
wire _721_ ;
wire _301_ ;
wire _5487_ ;
wire _5067_ ;
wire _3973_ ;
wire _3553_ ;
wire _3133_ ;
wire _4758_ ;
wire _4338_ ;
wire _37_ ;
wire _4091_ ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _2824_ ;
wire _2404_ ;
wire _5296_ ;
wire _3609_ ;
wire _3782_ ;
wire _3362_ ;
wire _4987_ ;
wire _4567_ ;
wire _4147_ ;
wire _2633_ ;
wire _2213_ ;
wire _3838_ ;
wire _3418_ ;
wire _3591_ ;
wire _3171_ ;
wire _1904_ ;
wire _4796_ ;
wire _4376_ ;
wire _815_ ;
wire _75_ ;
wire _6102_ ;
wire _2862_ ;
wire _2442_ ;
wire _2022_ ;
wire _3647_ ;
wire _3227_ ;
wire _1713_ ;
wire _4185_ ;
wire _624_ ;
wire _204_ ;
wire _2918_ ;
wire _6331_ ;
wire _2671_ ;
wire _2251_ ;
wire _3876_ ;
wire _3456_ ;
wire _3036_ ;
wire _5602_ ;
wire _1942_ ;
wire _1522_ ;
wire _1102_ ;
wire _853_ ;
wire _433_ ;
wire _2727_ ;
wire _2307_ ;
wire _5199_ ;
wire _6140_ ;
wire _2480_ ;
wire _2060_ ;
wire _3685_ ;
wire _3265_ ;
wire _5831_ ;
wire _5411_ ;
wire _909_ ;
wire _1751_ ;
wire _1331_ ;
wire _662_ ;
wire _242_ ;
wire _2956_ ;
wire _2536_ ;
wire _2116_ ;
wire _3494_ ;
wire _3074_ ;
wire _1807_ ;
wire _4699_ ;
wire _4279_ ;
wire _5640_ ;
wire _5220_ ;
wire _718_ ;
wire _6005_ ;
wire _1980_ ;
wire _1560_ ;
wire _1140_ ;
wire _891_ ;
wire _471_ ;
wire _2765_ ;
wire _2345_ ;
wire _4911_ ;
wire _1616_ ;
wire _4088_ ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _6234_ ;
wire _280_ ;
wire _2994_ ;
wire _2574_ ;
wire _2154_ ;
wire _3779_ ;
wire _3359_ ;
wire _4720_ ;
wire _4300_ ;
wire _5925_ ;
wire _5505_ ;
wire _1845_ ;
wire _1425_ ;
wire _1005_ ;
wire _756_ ;
wire _336_ ;
wire _6043_ ;
wire [15:0] _2383_ ;
wire _3588_ ;
wire _3168_ ;
wire _5734_ ;
wire _5314_ ;
wire _1654_ ;
wire _1234_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _2859_ ;
wire _2439_ ;
wire _2019_ ;
wire _3800_ ;
wire _6272_ ;
wire _2192_ ;
wire [15:0] \Y[2]  ;
wire _3397_ ;
wire _5963_ ;
wire _5543_ ;
wire _5123_ ;
wire _6328_ ;
wire _1883_ ;
wire _1463_ ;
wire _1043_ ;
wire [15:0] _794_ ;
wire _374_ ;
wire _2668_ ;
wire _2248_ ;
wire _6081_ ;
wire _4814_ ;
wire _1939_ ;
wire _1519_ ;
wire _5772_ ;
wire _5352_ ;
wire \X[3]_5_bF$buf2  ;
wire _6137_ ;
wire _1692_ ;
wire _1272_ ;
wire _183_ ;
wire _2897_ ;
wire _2477_ ;
wire _2057_ ;
wire _4623_ ;
wire _4203_ ;
wire _5828_ ;
wire _5408_ ;
wire _1748_ ;
wire _1328_ ;
wire _5581_ ;
wire _5161_ ;
wire _659_ ;
wire _239_ ;
wire _6366_ ;
wire _1081_ ;
wire _2286_ ;
wire _4852_ ;
wire _4432_ ;
wire _4012_ ;
wire _5637_ ;
wire _5217_ ;
wire _1977_ ;
wire _1557_ ;
wire _1137_ ;
wire _5390_ ;
wire _888_ ;
wire _468_ ;
wire _3703_ ;
wire _6175_ ;
wire _4908_ ;
wire _2095_ ;
wire _4661_ ;
wire _4241_ ;
wire _5866_ ;
wire _5446_ ;
wire _5026_ ;
wire _1786_ ;
wire _1366_ ;
wire _697_ ;
wire _277_ ;
wire _3932_ ;
wire _3512_ ;
wire _4717_ ;
wire _4890_ ;
wire _4470_ ;
wire _4050_ ;
wire _5675_ ;
wire _5255_ ;
wire _1595_ ;
wire _1175_ ;
wire _3741_ ;
wire _3321_ ;
wire _4946_ ;
wire _4526_ ;
wire _4106_ ;
wire _5484_ ;
wire _5064_ ;
wire _6269_ ;
wire _2189_ ;
wire _3970_ ;
wire _3550_ ;
wire _3130_ ;
wire _4755_ ;
wire _4335_ ;
wire _34_ ;
wire _2821_ ;
wire _2401_ ;
wire _5293_ ;
wire _3606_ ;
wire _6078_ ;
wire _4984_ ;
wire _4564_ ;
wire _4144_ ;
wire _5769_ ;
wire _5349_ ;
wire _1689_ ;
wire _1269_ ;
wire _2630_ ;
wire _2210_ ;
wire _3835_ ;
wire _3415_ ;
wire _1901_ ;
wire _4793_ ;
wire _4373_ ;
wire _812_ ;
wire _5998_ ;
wire [15:0] _5578_ ;
wire _5158_ ;
wire _72_ ;
wire _1498_ ;
wire _1078_ ;
wire _3644_ ;
wire _3224_ ;
wire _4849_ ;
wire _4429_ ;
wire _4009_ ;
wire _1710_ ;
wire _4182_ ;
wire _621_ ;
wire _201_ ;
wire _2915_ ;
wire _5387_ ;
wire _3873_ ;
wire _3453_ ;
wire _3033_ ;
wire _4658_ ;
wire _4238_ ;
wire _850_ ;
wire _430_ ;
wire _2724_ ;
wire _2304_ ;
wire _5196_ ;
wire _3929_ ;
wire _3509_ ;
wire _3682_ ;
wire _3262_ ;
wire _4887_ ;
wire _4467_ ;
wire _4047_ ;
wire _906_ ;
wire _2953_ ;
wire _2533_ ;
wire _2113_ ;
wire _3738_ ;
wire _3318_ ;
wire _3491_ ;
wire _3071_ ;
wire _1804_ ;
wire _4696_ ;
wire _4276_ ;
wire _715_ ;
wire _6002_ ;
wire _2762_ ;
wire _2342_ ;
wire _3967_ ;
wire _3547_ ;
wire _3127_ ;
wire _1613_ ;
wire _4085_ ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire _2818_ ;
wire _6231_ ;
wire _2991_ ;
wire _2571_ ;
wire _2151_ ;
wire _3776_ ;
wire _3356_ ;
wire _5922_ ;
wire _5502_ ;
wire _1842_ ;
wire _1422_ ;
wire _1002_ ;
wire _753_ ;
wire _333_ ;
wire _2627_ ;
wire _2207_ ;
wire _5099_ ;
wire _6040_ ;
wire _2380_ ;
wire _3585_ ;
wire _3165_ ;
wire _5731_ ;
wire _5311_ ;
wire _809_ ;
wire _69_ ;
wire _1651_ ;
wire _1231_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _2856_ ;
wire _2436_ ;
wire _2016_ ;
wire _3394_ ;
wire _1707_ ;
wire _4599_ ;
wire _4179_ ;
wire _5960_ ;
wire _5540_ ;
wire _5120_ ;
wire _618_ ;
wire _6325_ ;
wire _1880_ ;
wire _1460_ ;
wire _1040_ ;
wire [15:0] _791_ ;
wire _371_ ;
wire _2665_ ;
wire _2245_ ;
wire _4811_ ;
wire _1936_ ;
wire _1516_ ;
wire _847_ ;
wire _427_ ;
wire _6134_ ;
wire _180_ ;
wire _2894_ ;
wire _2474_ ;
wire _2054_ ;
wire _3679_ ;
wire _3259_ ;
wire _4620_ ;
wire _4200_ ;
wire _5825_ ;
wire _5405_ ;
wire _1745_ ;
wire _1325_ ;
wire _656_ ;
wire _236_ ;
wire _6363_ ;
wire _2283_ ;
wire _3488_ ;
wire _3068_ ;
wire _5634_ ;
wire _5214_ ;
wire _1974_ ;
wire _1554_ ;
wire _1134_ ;
wire _885_ ;
wire _465_ ;
wire _2759_ ;
wire _2339_ ;
wire _3700_ ;
wire _6172_ ;
wire _4905_ ;
wire _2092_ ;
wire _3297_ ;
wire _5863_ ;
wire _5443_ ;
wire _5023_ ;
wire _6228_ ;
wire _1783_ ;
wire _1363_ ;
wire _694_ ;
wire _274_ ;
wire _2988_ ;
wire _2568_ ;
wire _2148_ ;
wire _4714_ ;
wire _5919_ ;
wire _1839_ ;
wire _1419_ ;
wire _5672_ ;
wire _5252_ ;
wire _6037_ ;
wire [15:0] _1592_ ;
wire _1172_ ;
wire _2797_ ;
wire _2377_ ;
wire _4943_ ;
wire _4523_ ;
wire _4103_ ;
wire _5728_ ;
wire _5308_ ;
wire _1648_ ;
wire _1228_ ;
wire _5481_ ;
wire _5061_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _6266_ ;
wire _2186_ ;
wire _4752_ ;
wire _4332_ ;
wire _5957_ ;
wire _5537_ ;
wire _5117_ ;
wire _31_ ;
wire _1877_ ;
wire _1457_ ;
wire _1037_ ;
wire _5290_ ;
wire _788_ ;
wire _368_ ;
wire _3603_ ;
wire _6075_ ;
wire _4808_ ;
wire _4981_ ;
wire _4561_ ;
wire _4141_ ;
wire _5766_ ;
wire _5346_ ;
wire _1686_ ;
wire _1266_ ;
wire _597_ ;
wire _177_ ;
wire _3832_ ;
wire _3412_ ;
wire _4617_ ;
wire _4790_ ;
wire _4370_ ;
wire _5995_ ;
wire [15:0] _5575_ ;
wire _5155_ ;
wire _1495_ ;
wire _1075_ ;
wire _3641_ ;
wire _3221_ ;
wire _4846_ ;
wire _4426_ ;
wire _4006_ ;
wire _2912_ ;
wire _5384_ ;
wire _6169_ ;
wire _2089_ ;
wire _3870_ ;
wire _3450_ ;
wire _3030_ ;
wire _4655_ ;
wire _4235_ ;
wire _2721_ ;
wire _2301_ ;
wire _5193_ ;
wire _3926_ ;
wire _3506_ ;
wire _4884_ ;
wire _4464_ ;
wire _4044_ ;
wire _903_ ;
wire _5669_ ;
wire _5249_ ;
wire [15:0] _1589_ ;
wire _1169_ ;
wire _2950_ ;
wire _2530_ ;
wire _2110_ ;
wire _3735_ ;
wire _3315_ ;
wire _1801_ ;
wire _4693_ ;
wire _4273_ ;
wire _712_ ;
wire _5898_ ;
wire _5478_ ;
wire _5058_ ;
wire _1398_ ;
wire _3964_ ;
wire _3544_ ;
wire _3124_ ;
wire _4749_ ;
wire _4329_ ;
wire _28_ ;
wire _1610_ ;
wire _4082_ ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _2815_ ;
wire _5287_ ;
wire _3773_ ;
wire _3353_ ;
wire _4978_ ;
wire _4558_ ;
wire _4138_ ;
wire _750_ ;
wire _330_ ;
wire _2624_ ;
wire _2204_ ;
wire _5096_ ;
wire _3829_ ;
wire _3409_ ;
wire _3582_ ;
wire _3162_ ;
wire _4787_ ;
wire _4367_ ;
wire _806_ ;
wire _66_ ;
wire _2853_ ;
wire _2433_ ;
wire _2013_ ;
wire _3638_ ;
wire _3218_ ;
wire _3391_ ;
wire _1704_ ;
wire _4596_ ;
wire _4176_ ;
wire _615_ ;
wire _2909_ ;
wire _6322_ ;
wire _2662_ ;
wire _2242_ ;
wire _3867_ ;
wire _3447_ ;
wire _3027_ ;
wire _1933_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire _2718_ ;
wire \X[2]_5_bF$buf1  ;
wire _6131_ ;
wire _2891_ ;
wire _2471_ ;
wire _2051_ ;
wire _3676_ ;
wire _3256_ ;
wire _5822_ ;
wire _5402_ ;
wire _1742_ ;
wire _1322_ ;
wire _653_ ;
wire _233_ ;
wire _2947_ ;
wire _2527_ ;
wire _2107_ ;
wire _6360_ ;
wire _2280_ ;
wire _3485_ ;
wire _3065_ ;
wire _5631_ ;
wire _5211_ ;
wire _709_ ;
wire _1971_ ;
wire _1551_ ;
wire _1131_ ;
wire _882_ ;
wire _462_ ;
wire _2756_ ;
wire _2336_ ;
wire _4902_ ;
wire _3294_ ;
wire _1607_ ;
wire _4499_ ;
wire _4079_ ;
wire _5860_ ;
wire _5440_ ;
wire _5020_ ;
wire _938_ ;
wire _518_ ;
wire _6225_ ;
wire _1780_ ;
wire _1360_ ;
wire _691_ ;
wire _271_ ;
wire _2985_ ;
wire _2565_ ;
wire _2145_ ;
wire _4711_ ;
wire _5916_ ;
wire _1836_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _6034_ ;
wire _2794_ ;
wire _2374_ ;
wire _3999_ ;
wire _3579_ ;
wire _3159_ ;
wire _4940_ ;
wire _4520_ ;
wire _4100_ ;
wire _5725_ ;
wire _5305_ ;
wire _1645_ ;
wire _1225_ ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire _6263_ ;
wire _2183_ ;
wire _3388_ ;
wire _5954_ ;
wire _5534_ ;
wire _5114_ ;
wire _6319_ ;
wire _1874_ ;
wire _1454_ ;
wire _1034_ ;
wire _785_ ;
wire _365_ ;
wire _2659_ ;
wire _2239_ ;
wire _3600_ ;
wire _6072_ ;
wire _4805_ ;
wire _3197_ ;
wire _5763_ ;
wire _5343_ ;
wire _6128_ ;
wire _1683_ ;
wire _1263_ ;
wire _594_ ;
wire _174_ ;
wire _2888_ ;
wire _2468_ ;
wire _2048_ ;
wire _4614_ ;
wire _5819_ ;
wire _1739_ ;
wire _1319_ ;
wire _5992_ ;
wire [15:0] _5572_ ;
wire _5152_ ;
wire _6357_ ;
wire _1492_ ;
wire _1072_ ;
wire _2697_ ;
wire _2277_ ;
wire _4843_ ;
wire _4423_ ;
wire _4003_ ;
wire _5628_ ;
wire _5208_ ;
wire _1968_ ;
wire _1548_ ;
wire _1128_ ;
wire _5381_ ;
wire _879_ ;
wire _459_ ;
wire _6166_ ;
wire _2086_ ;
wire _4652_ ;
wire _4232_ ;
wire _5857_ ;
wire _5437_ ;
wire _5017_ ;
wire _1777_ ;
wire _1357_ ;
wire _5190_ ;
wire _688_ ;
wire _268_ ;
wire _3923_ ;
wire _3503_ ;
wire _4708_ ;
wire _4881_ ;
wire _4461_ ;
wire _4041_ ;
wire _900_ ;
wire _5666_ ;
wire _5246_ ;
wire [15:0] _1586_ ;
wire _1166_ ;
wire [15:0] \u_fir_pe1.rYin  ;
wire _497_ ;
wire _3732_ ;
wire _3312_ ;
wire _4937_ ;
wire _4517_ ;
wire _4690_ ;
wire _4270_ ;
wire _5895_ ;
wire _5475_ ;
wire _5055_ ;
wire _1395_ ;
wire _3961_ ;
wire _3541_ ;
wire _3121_ ;
wire _4746_ ;
wire _4326_ ;
wire _25_ ;
wire _2812_ ;
wire _5284_ ;
wire _6069_ ;
wire _3770_ ;
wire _3350_ ;
wire _4975_ ;
wire _4555_ ;
wire _4135_ ;
wire _2621_ ;
wire _2201_ ;
wire _5093_ ;
wire _3826_ ;
wire _3406_ ;
wire _6298_ ;
wire _4784_ ;
wire _4364_ ;
wire _803_ ;
wire _5989_ ;
wire _5569_ ;
wire _5149_ ;
wire _63_ ;
wire _1489_ ;
wire _1069_ ;
wire _2850_ ;
wire _2430_ ;
wire _2010_ ;
wire _3635_ ;
wire _3215_ ;
wire [7:0] \X[7]  ;
wire _1701_ ;
wire _4593_ ;
wire _4173_ ;
wire _612_ ;
wire _2906_ ;
wire _5798_ ;
wire _5378_ ;
wire _1298_ ;
wire _3864_ ;
wire _3444_ ;
wire _3024_ ;
wire _4649_ ;
wire _4229_ ;
wire _1930_ ;
wire _1510_ ;
wire _841_ ;
wire _421_ ;
wire _2715_ ;
wire _5187_ ;
wire \X[1]_5_bF$buf3  ;
wire _3673_ ;
wire _3253_ ;
wire _4878_ ;
wire _4458_ ;
wire _4038_ ;
wire _650_ ;
wire _230_ ;
wire _2944_ ;
wire _2524_ ;
wire _2104_ ;
wire _3729_ ;
wire _3309_ ;
wire _3482_ ;
wire _3062_ ;
wire _4687_ ;
wire _4267_ ;
wire _706_ ;
wire _2753_ ;
wire _2333_ ;
wire _3958_ ;
wire _3538_ ;
wire _3118_ ;
wire _3291_ ;
wire _1604_ ;
wire _4496_ ;
wire _4076_ ;
wire _935_ ;
wire _515_ ;
wire _2809_ ;
wire _6222_ ;
wire _2982_ ;
wire _2562_ ;
wire _2142_ ;
wire _3767_ ;
wire _3347_ ;
wire _5913_ ;
wire _1833_ ;
wire _1413_ ;
wire _744_ ;
wire _324_ ;
wire _2618_ ;
wire _6031_ ;
wire _2791_ ;
wire _2371_ ;
wire _3996_ ;
wire _3576_ ;
wire _3156_ ;
wire _5722_ ;
wire _5302_ ;
wire _1642_ ;
wire _1222_ ;
wire _973_ ;
wire _553_ ;
wire _133_ ;
wire _2847_ ;
wire _2427_ ;
wire _2007_ ;
wire _6260_ ;
wire _2180_ ;
wire _3385_ ;
wire _5951_ ;
wire _5531_ ;
wire _5111_ ;
wire _609_ ;
wire _6316_ ;
wire _1871_ ;
wire _1451_ ;
wire _1031_ ;
wire _782_ ;
wire _362_ ;
wire _2656_ ;
wire _2236_ ;
wire _4802_ ;
wire _3194_ ;
wire _1927_ ;
wire _1507_ ;
wire _4399_ ;
wire _5760_ ;
wire _5340_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _6125_ ;
wire _1680_ ;
wire _1260_ ;
wire _591_ ;
wire _171_ ;
wire _2885_ ;
wire _2465_ ;
wire _2045_ ;
wire _4611_ ;
wire _5816_ ;
wire _1736_ ;
wire _1316_ ;
wire _647_ ;
wire _227_ ;
wire _6354_ ;
wire _2694_ ;
wire _2274_ ;
wire _3899_ ;
wire _3479_ ;
wire _3059_ ;
wire _4840_ ;
wire _4420_ ;
wire _4000_ ;
wire _5625_ ;
wire _5205_ ;
wire _1965_ ;
wire _1545_ ;
wire _1125_ ;
wire _876_ ;
wire _456_ ;
wire _6163_ ;
wire _2083_ ;
wire _3288_ ;
wire _5854_ ;
wire _5434_ ;
wire _5014_ ;
wire _6219_ ;
wire _1774_ ;
wire _1354_ ;
wire _685_ ;
wire _265_ ;
wire _2979_ ;
wire _2559_ ;
wire _2139_ ;
wire _3920_ ;
wire _3500_ ;
wire _4705_ ;
wire _3097_ ;
wire _5663_ ;
wire _5243_ ;
wire [15:0] \u_fir_pe0.mul  ;
wire _6028_ ;
wire _1583_ ;
wire _1163_ ;
wire _494_ ;
wire _2788_ ;
wire _2368_ ;
wire _4934_ ;
wire _4514_ ;
wire _5719_ ;
wire _1639_ ;
wire _1219_ ;
wire _5892_ ;
wire _5472_ ;
wire _5052_ ;
wire _6257_ ;
wire _1392_ ;
wire _2597_ ;
wire _2177_ ;
wire _4743_ ;
wire _4323_ ;
wire \X[7]_5_bF$buf2  ;
wire _5948_ ;
wire _5528_ ;
wire _5108_ ;
wire _22_ ;
wire _1868_ ;
wire _1448_ ;
wire _1028_ ;
wire _5281_ ;
wire _779_ ;
wire _359_ ;
wire _6066_ ;

CLKBUF1 CLKBUF1_insert96 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_hier0_bF$buf0)
);

CLKBUF1 CLKBUF1_insert95 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_hier0_bF$buf1)
);

CLKBUF1 CLKBUF1_insert94 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_hier0_bF$buf2)
);

CLKBUF1 CLKBUF1_insert93 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_hier0_bF$buf3)
);

CLKBUF1 CLKBUF1_insert92 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_hier0_bF$buf4)
);

CLKBUF1 CLKBUF1_insert91 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_hier0_bF$buf5)
);

CLKBUF1 CLKBUF1_insert90 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_hier0_bF$buf6)
);

BUFX2 BUFX2_insert89 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [5]),
    .Y(\X[7]_5_bF$buf0 )
);

BUFX2 BUFX2_insert88 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [5]),
    .Y(\X[7]_5_bF$buf1 )
);

BUFX2 BUFX2_insert87 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [5]),
    .Y(\X[7]_5_bF$buf2 )
);

BUFX2 BUFX2_insert86 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [5]),
    .Y(\X[7]_5_bF$buf3 )
);

BUFX2 BUFX2_insert85 (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[5]),
    .Y(Xin_5_bF$buf0)
);

BUFX2 BUFX2_insert84 (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[5]),
    .Y(Xin_5_bF$buf1)
);

BUFX2 BUFX2_insert83 (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[5]),
    .Y(Xin_5_bF$buf2)
);

BUFX2 BUFX2_insert82 (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[5]),
    .Y(Xin_5_bF$buf3)
);

BUFX2 BUFX2_insert81 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [5]),
    .Y(\X[6]_5_bF$buf0 )
);

BUFX2 BUFX2_insert80 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [5]),
    .Y(\X[6]_5_bF$buf1 )
);

BUFX2 BUFX2_insert79 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [5]),
    .Y(\X[6]_5_bF$buf2 )
);

BUFX2 BUFX2_insert78 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [5]),
    .Y(\X[6]_5_bF$buf3 )
);

BUFX2 BUFX2_insert77 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [5]),
    .Y(\X[4]_5_bF$buf0 )
);

BUFX2 BUFX2_insert76 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [5]),
    .Y(\X[4]_5_bF$buf1 )
);

BUFX2 BUFX2_insert75 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [5]),
    .Y(\X[4]_5_bF$buf2 )
);

BUFX2 BUFX2_insert74 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [5]),
    .Y(\X[4]_5_bF$buf3 )
);

BUFX2 BUFX2_insert73 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [5]),
    .Y(\X[2]_5_bF$buf0 )
);

BUFX2 BUFX2_insert72 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [5]),
    .Y(\X[2]_5_bF$buf1 )
);

BUFX2 BUFX2_insert71 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [5]),
    .Y(\X[2]_5_bF$buf2 )
);

BUFX2 BUFX2_insert70 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [5]),
    .Y(\X[2]_5_bF$buf3 )
);

CLKBUF1 CLKBUF1_insert69 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert68 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert67 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert66 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert65 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert64 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert63 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert62 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert61 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf8)
);

CLKBUF1 CLKBUF1_insert60 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf9)
);

CLKBUF1 CLKBUF1_insert59 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf10)
);

CLKBUF1 CLKBUF1_insert58 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf11)
);

CLKBUF1 CLKBUF1_insert57 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf12)
);

CLKBUF1 CLKBUF1_insert56 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf13)
);

CLKBUF1 CLKBUF1_insert55 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf14)
);

CLKBUF1 CLKBUF1_insert54 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf15)
);

CLKBUF1 CLKBUF1_insert53 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf16)
);

CLKBUF1 CLKBUF1_insert52 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf17)
);

CLKBUF1 CLKBUF1_insert51 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf18)
);

CLKBUF1 CLKBUF1_insert50 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf19)
);

CLKBUF1 CLKBUF1_insert49 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf20)
);

CLKBUF1 CLKBUF1_insert48 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf21)
);

CLKBUF1 CLKBUF1_insert47 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf22)
);

CLKBUF1 CLKBUF1_insert46 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf23)
);

CLKBUF1 CLKBUF1_insert45 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf24)
);

CLKBUF1 CLKBUF1_insert44 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf25)
);

CLKBUF1 CLKBUF1_insert43 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf26)
);

CLKBUF1 CLKBUF1_insert42 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf27)
);

CLKBUF1 CLKBUF1_insert41 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf28)
);

CLKBUF1 CLKBUF1_insert40 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf29)
);

CLKBUF1 CLKBUF1_insert39 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf30)
);

CLKBUF1 CLKBUF1_insert38 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf31)
);

CLKBUF1 CLKBUF1_insert37 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf32)
);

CLKBUF1 CLKBUF1_insert36 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf33)
);

CLKBUF1 CLKBUF1_insert35 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf34)
);

CLKBUF1 CLKBUF1_insert34 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf35)
);

CLKBUF1 CLKBUF1_insert33 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf36)
);

CLKBUF1 CLKBUF1_insert32 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf37)
);

CLKBUF1 CLKBUF1_insert31 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf38)
);

CLKBUF1 CLKBUF1_insert30 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf39)
);

CLKBUF1 CLKBUF1_insert29 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf40)
);

CLKBUF1 CLKBUF1_insert28 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf41)
);

CLKBUF1 CLKBUF1_insert27 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf42)
);

CLKBUF1 CLKBUF1_insert26 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf43)
);

CLKBUF1 CLKBUF1_insert25 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf44)
);

CLKBUF1 CLKBUF1_insert24 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf45)
);

CLKBUF1 CLKBUF1_insert23 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf46)
);

CLKBUF1 CLKBUF1_insert22 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf47)
);

CLKBUF1 CLKBUF1_insert21 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf48)
);

CLKBUF1 CLKBUF1_insert20 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf49)
);

CLKBUF1 CLKBUF1_insert19 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf50)
);

CLKBUF1 CLKBUF1_insert18 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf51)
);

CLKBUF1 CLKBUF1_insert17 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf52)
);

CLKBUF1 CLKBUF1_insert16 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf53)
);

CLKBUF1 CLKBUF1_insert15 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf54)
);

CLKBUF1 CLKBUF1_insert14 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf55)
);

CLKBUF1 CLKBUF1_insert13 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf56)
);

CLKBUF1 CLKBUF1_insert12 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf57)
);

BUFX2 BUFX2_insert11 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [5]),
    .Y(\X[5]_5_bF$buf0 )
);

BUFX2 BUFX2_insert10 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [5]),
    .Y(\X[5]_5_bF$buf1 )
);

BUFX2 BUFX2_insert9 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [5]),
    .Y(\X[5]_5_bF$buf2 )
);

BUFX2 BUFX2_insert8 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [5]),
    .Y(\X[5]_5_bF$buf3 )
);

BUFX2 BUFX2_insert7 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [5]),
    .Y(\X[3]_5_bF$buf0 )
);

BUFX2 BUFX2_insert6 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [5]),
    .Y(\X[3]_5_bF$buf1 )
);

BUFX2 BUFX2_insert5 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [5]),
    .Y(\X[3]_5_bF$buf2 )
);

BUFX2 BUFX2_insert4 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [5]),
    .Y(\X[3]_5_bF$buf3 )
);

BUFX2 BUFX2_insert3 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [5]),
    .Y(\X[1]_5_bF$buf0 )
);

BUFX2 BUFX2_insert2 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [5]),
    .Y(\X[1]_5_bF$buf1 )
);

BUFX2 BUFX2_insert1 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [5]),
    .Y(\X[1]_5_bF$buf2 )
);

BUFX2 BUFX2_insert0 (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [5]),
    .Y(\X[1]_5_bF$buf3 )
);

NAND2X1 _10000_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [3]),
    .Y(_3281_)
);

NAND3X1 _10001_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [2]),
    .C(_3281_),
    .Y(_3282_)
);

NAND3X1 _10002_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3273_),
    .B(_3280_),
    .C(_3282_),
    .Y(_3283_)
);

NAND3X1 _10003_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3272_),
    .B(_3283_),
    .C(_3279_),
    .Y(_3284_)
);

INVX1 _10004_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3272_),
    .Y(_3285_)
);

AOI21X1 _10005_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3280_),
    .B(_3282_),
    .C(_3273_),
    .Y(_3286_)
);

AOI22X1 _10006_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[4] [4]),
    .C(_3276_),
    .D(_3278_),
    .Y(_3287_)
);

OAI21X1 _10007_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3286_),
    .B(_3287_),
    .C(_3285_),
    .Y(_3288_)
);

NAND3X1 _10008_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3284_),
    .B(_3270_),
    .C(_3288_),
    .Y(_3289_)
);

NAND2X1 _10009_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3269_),
    .B(_3265_),
    .Y(_3290_)
);

OAI21X1 _10010_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3286_),
    .B(_3287_),
    .C(_3272_),
    .Y(_3291_)
);

NAND3X1 _10011_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3283_),
    .B(_3279_),
    .C(_3285_),
    .Y(_3292_)
);

NAND3X1 _10012_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3290_),
    .B(_3292_),
    .C(_3291_),
    .Y(_3293_)
);

NAND3X1 _10013_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3289_),
    .B(_3293_),
    .C(_3257_),
    .Y(_3294_)
);

AOI21X1 _10014_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3216_),
    .B(_3236_),
    .C(_3250_),
    .Y(_3295_)
);

AOI21X1 _10015_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3291_),
    .B(_3292_),
    .C(_3290_),
    .Y(_3296_)
);

AOI21X1 _10016_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3288_),
    .B(_3284_),
    .C(_3270_),
    .Y(_3297_)
);

OAI21X1 _10017_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3296_),
    .B(_3297_),
    .C(_3295_),
    .Y(_3298_)
);

NAND3X1 _10018_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3214_),
    .B(_3294_),
    .C(_3298_),
    .Y(_3299_)
);

INVX1 _10019_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3214_),
    .Y(_3300_)
);

OAI21X1 _10020_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3296_),
    .B(_3297_),
    .C(_3257_),
    .Y(_3301_)
);

NAND3X1 _10021_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3289_),
    .B(_3293_),
    .C(_3295_),
    .Y(_3302_)
);

NAND3X1 _10022_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3300_),
    .B(_3301_),
    .C(_3302_),
    .Y(_3303_)
);

NAND3X1 _10023_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3241_),
    .B(_3299_),
    .C(_3303_),
    .Y(_3304_)
);

NAND3X1 _10024_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3300_),
    .B(_3294_),
    .C(_3298_),
    .Y(_3305_)
);

NAND3X1 _10025_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3214_),
    .B(_3301_),
    .C(_3302_),
    .Y(_3306_)
);

NAND3X1 _10026_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3242_),
    .B(_3305_),
    .C(_3306_),
    .Y(_3307_)
);

NAND3X1 _10027_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3304_),
    .B(_3307_),
    .C(_3256_),
    .Y(_3308_)
);

INVX1 _10028_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3208_),
    .Y(_3309_)
);

NAND3X1 _10029_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3309_),
    .B(_3242_),
    .C(_3245_),
    .Y(_3310_)
);

NAND3X1 _10030_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3242_),
    .B(_3299_),
    .C(_3303_),
    .Y(_3311_)
);

NAND3X1 _10031_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3241_),
    .B(_3305_),
    .C(_3306_),
    .Y(_3312_)
);

NAND3X1 _10032_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3311_),
    .B(_3312_),
    .C(_3310_),
    .Y(_3313_)
);

NAND3X1 _10033_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3308_),
    .B(_3313_),
    .C(_3255_),
    .Y(_3314_)
);

INVX1 _10034_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3255_),
    .Y(_3315_)
);

INVX1 _10035_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3308_),
    .Y(_3316_)
);

INVX1 _10036_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3313_),
    .Y(_3317_)
);

OAI21X1 _10037_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3316_),
    .B(_3317_),
    .C(_3315_),
    .Y(_3318_)
);

AND2X2 _10038_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3318_),
    .B(_3314_),
    .Y(_3984_[5])
);

AND2X2 _10039_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [0]),
    .B(gnd),
    .Y(_3319_)
);

NAND2X1 _10040_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4]_5_bF$buf3 ),
    .Y(_3320_)
);

OAI21X1 _10041_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3898_),
    .B(_3320_),
    .C(_3265_),
    .Y(_3321_)
);

OR2X2 _10042_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3321_),
    .B(_3319_),
    .Y(_3322_)
);

NAND2X1 _10043_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3319_),
    .B(_3321_),
    .Y(_3323_)
);

NAND2X1 _10044_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3323_),
    .B(_3322_),
    .Y(_3324_)
);

AOI21X1 _10045_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3279_),
    .B(_3283_),
    .C(_3272_),
    .Y(_3325_)
);

OAI21X1 _10046_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3290_),
    .B(_3325_),
    .C(_3284_),
    .Y(_3326_)
);

NAND2X1 _10047_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [1]),
    .B(vdd),
    .Y(_3327_)
);

INVX1 _10048_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3327_),
    .Y(_3328_)
);

AND2X2 _10049_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [2]),
    .B(gnd),
    .Y(_3329_)
);

AND2X2 _10050_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [6]),
    .Y(_3330_)
);

NAND2X1 _10051_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3329_),
    .B(_3330_),
    .Y(_3331_)
);

INVX2 _10052_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [6]),
    .Y(_3332_)
);

NAND2X1 _10053_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [2]),
    .B(gnd),
    .Y(_3333_)
);

OAI21X1 _10054_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3966_),
    .B(_3332_),
    .C(_3333_),
    .Y(_3334_)
);

NAND3X1 _10055_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3334_),
    .B(_3328_),
    .C(_3331_),
    .Y(_3335_)
);

NAND3X1 _10056_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [6]),
    .C(_3333_),
    .Y(_3336_)
);

NAND2X1 _10057_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [6]),
    .Y(_3337_)
);

NAND2X1 _10058_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3337_),
    .B(_3329_),
    .Y(_3338_)
);

NAND3X1 _10059_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3327_),
    .B(_3336_),
    .C(_3338_),
    .Y(_3339_)
);

AND2X2 _10060_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3335_),
    .B(_3339_),
    .Y(_3340_)
);

NAND2X1 _10061_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [3]),
    .Y(_3341_)
);

AOI22X1 _10062_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [2]),
    .C(gnd),
    .D(\X[4] [3]),
    .Y(_3342_)
);

OAI22X1 _10063_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3230_),
    .B(_3341_),
    .C(_3273_),
    .D(_3342_),
    .Y(_3343_)
);

NAND2X1 _10064_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[4]_5_bF$buf2 ),
    .Y(_3344_)
);

INVX1 _10065_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3344_),
    .Y(_3345_)
);

AND2X2 _10066_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [4]),
    .Y(_3346_)
);

NAND2X1 _10067_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3275_),
    .B(_3346_),
    .Y(_3347_)
);

AOI22X1 _10068_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [3]),
    .C(gnd),
    .D(\X[4] [4]),
    .Y(_3348_)
);

INVX1 _10069_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3348_),
    .Y(_3349_)
);

NAND3X1 _10070_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3345_),
    .B(_3349_),
    .C(_3347_),
    .Y(_3350_)
);

NAND3X1 _10071_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [4]),
    .C(_3341_),
    .Y(_3351_)
);

NAND2X1 _10072_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [4]),
    .Y(_3352_)
);

NAND3X1 _10073_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [3]),
    .C(_3352_),
    .Y(_3353_)
);

NAND3X1 _10074_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3344_),
    .B(_3351_),
    .C(_3353_),
    .Y(_3354_)
);

NAND3X1 _10075_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3343_),
    .B(_3354_),
    .C(_3350_),
    .Y(_3355_)
);

INVX1 _10076_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3343_),
    .Y(_3356_)
);

AOI21X1 _10077_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3351_),
    .B(_3353_),
    .C(_3344_),
    .Y(_3357_)
);

AOI22X1 _10078_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[4]_5_bF$buf1 ),
    .C(_3347_),
    .D(_3349_),
    .Y(_3358_)
);

OAI21X1 _10079_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3357_),
    .B(_3358_),
    .C(_3356_),
    .Y(_3359_)
);

NAND3X1 _10080_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3355_),
    .B(_3340_),
    .C(_3359_),
    .Y(_3360_)
);

NAND2X1 _10081_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3339_),
    .B(_3335_),
    .Y(_3361_)
);

OAI21X1 _10082_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3357_),
    .B(_3358_),
    .C(_3343_),
    .Y(_3362_)
);

NAND3X1 _10083_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3350_),
    .B(_3354_),
    .C(_3356_),
    .Y(_3363_)
);

NAND3X1 _10084_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3361_),
    .B(_3363_),
    .C(_3362_),
    .Y(_3364_)
);

NAND3X1 _10085_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3360_),
    .B(_3326_),
    .C(_3364_),
    .Y(_3365_)
);

INVX1 _10086_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3284_),
    .Y(_3366_)
);

AOI21X1 _10087_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3270_),
    .B(_3288_),
    .C(_3366_),
    .Y(_3367_)
);

AOI21X1 _10088_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3362_),
    .B(_3363_),
    .C(_3361_),
    .Y(_3368_)
);

AOI21X1 _10089_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3359_),
    .B(_3355_),
    .C(_3340_),
    .Y(_3369_)
);

OAI21X1 _10090_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3368_),
    .B(_3369_),
    .C(_3367_),
    .Y(_3370_)
);

NAND3X1 _10091_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3324_),
    .B(_3365_),
    .C(_3370_),
    .Y(_3371_)
);

AND2X2 _10092_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3322_),
    .B(_3323_),
    .Y(_3372_)
);

OAI21X1 _10093_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3368_),
    .B(_3369_),
    .C(_3326_),
    .Y(_3373_)
);

NAND3X1 _10094_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3360_),
    .B(_3364_),
    .C(_3367_),
    .Y(_3374_)
);

NAND3X1 _10095_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3372_),
    .B(_3373_),
    .C(_3374_),
    .Y(_3375_)
);

AOI22X1 _10096_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3299_),
    .B(_3294_),
    .C(_3371_),
    .D(_3375_),
    .Y(_3376_)
);

AOI21X1 _10097_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3289_),
    .B(_3293_),
    .C(_3257_),
    .Y(_3377_)
);

OAI21X1 _10098_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3300_),
    .B(_3377_),
    .C(_3294_),
    .Y(_3378_)
);

NAND3X1 _10099_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3372_),
    .B(_3365_),
    .C(_3370_),
    .Y(_3379_)
);

NAND3X1 _10100_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3324_),
    .B(_3373_),
    .C(_3374_),
    .Y(_3380_)
);

AOI21X1 _10101_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3380_),
    .B(_3379_),
    .C(_3378_),
    .Y(_3381_)
);

OAI21X1 _10102_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3381_),
    .B(_3376_),
    .C(_3304_),
    .Y(_3382_)
);

AOI21X1 _10103_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3306_),
    .B(_3305_),
    .C(_3242_),
    .Y(_3383_)
);

NAND3X1 _10104_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3378_),
    .B(_3379_),
    .C(_3380_),
    .Y(_3384_)
);

INVX1 _10105_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3294_),
    .Y(_3385_)
);

AOI21X1 _10106_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3214_),
    .B(_3298_),
    .C(_3385_),
    .Y(_3386_)
);

AOI21X1 _10107_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3374_),
    .B(_3373_),
    .C(_3324_),
    .Y(_3387_)
);

AOI21X1 _10108_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3370_),
    .B(_3365_),
    .C(_3372_),
    .Y(_3388_)
);

OAI21X1 _10109_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3387_),
    .B(_3388_),
    .C(_3386_),
    .Y(_3389_)
);

NAND3X1 _10110_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3383_),
    .B(_3384_),
    .C(_3389_),
    .Y(_3390_)
);

NAND2X1 _10111_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3390_),
    .B(_3382_),
    .Y(_3391_)
);

AOI21X1 _10112_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3308_),
    .B(_3314_),
    .C(_3391_),
    .Y(_3392_)
);

OAI21X1 _10113_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3317_),
    .B(_3315_),
    .C(_3308_),
    .Y(_3393_)
);

AOI21X1 _10114_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3382_),
    .B(_3390_),
    .C(_3393_),
    .Y(_3394_)
);

NOR2X1 _10115_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3392_),
    .B(_3394_),
    .Y(_3984_[6])
);

INVX1 _10116_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3390_),
    .Y(_3395_)
);

AOI21X1 _10117_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3360_),
    .B(_3364_),
    .C(_3326_),
    .Y(_3396_)
);

OAI21X1 _10118_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3324_),
    .B(_3396_),
    .C(_3365_),
    .Y(_3397_)
);

NAND2X1 _10119_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [0]),
    .B(gnd),
    .Y(_3398_)
);

INVX1 _10120_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3398_),
    .Y(_3399_)
);

NAND2X1 _10121_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [1]),
    .B(gnd),
    .Y(_3400_)
);

INVX1 _10122_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3400_),
    .Y(_3401_)
);

AND2X2 _10123_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3333_),
    .B(_3337_),
    .Y(_3402_)
);

OAI21X1 _10124_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3327_),
    .B(_3402_),
    .C(_3331_),
    .Y(_3403_)
);

NAND2X1 _10125_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3401_),
    .B(_3403_),
    .Y(_3404_)
);

NAND3X1 _10126_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3331_),
    .B(_3400_),
    .C(_3335_),
    .Y(_3405_)
);

NAND3X1 _10127_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3399_),
    .B(_3405_),
    .C(_3404_),
    .Y(_3406_)
);

AOI21X1 _10128_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3335_),
    .B(_3331_),
    .C(_3400_),
    .Y(_3407_)
);

NOR2X1 _10129_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3401_),
    .B(_3403_),
    .Y(_3408_)
);

OAI21X1 _10130_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3407_),
    .B(_3408_),
    .C(_3398_),
    .Y(_3409_)
);

NAND2X1 _10131_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3406_),
    .B(_3409_),
    .Y(_3410_)
);

AOI21X1 _10132_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3350_),
    .B(_3354_),
    .C(_3343_),
    .Y(_3411_)
);

OAI21X1 _10133_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3361_),
    .B(_3411_),
    .C(_3355_),
    .Y(_3412_)
);

NAND2X1 _10134_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [2]),
    .B(vdd),
    .Y(_3413_)
);

INVX1 _10135_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3413_),
    .Y(_3414_)
);

AND2X2 _10136_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [3]),
    .B(gnd),
    .Y(_3415_)
);

AND2X2 _10137_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [7]),
    .Y(_3416_)
);

NAND2X1 _10138_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3415_),
    .B(_3416_),
    .Y(_3417_)
);

AOI22X1 _10139_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [7]),
    .C(\X[4] [3]),
    .D(gnd),
    .Y(_3418_)
);

INVX1 _10140_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3418_),
    .Y(_3419_)
);

NAND3X1 _10141_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3414_),
    .B(_3419_),
    .C(_3417_),
    .Y(_3420_)
);

INVX1 _10142_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_3421_)
);

OAI21X1 _10143_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3203_),
    .B(_3421_),
    .C(_3416_),
    .Y(_3422_)
);

INVX1 _10144_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [7]),
    .Y(_3423_)
);

OAI21X1 _10145_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3966_),
    .B(_3423_),
    .C(_3415_),
    .Y(_3424_)
);

NAND3X1 _10146_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3413_),
    .B(_3422_),
    .C(_3424_),
    .Y(_3425_)
);

NAND2X1 _10147_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3420_),
    .B(_3425_),
    .Y(_3426_)
);

OAI21X1 _10148_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3344_),
    .B(_3348_),
    .C(_3347_),
    .Y(_3427_)
);

NAND2X1 _10149_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[4] [6]),
    .Y(_3428_)
);

NAND2X1 _10150_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [4]),
    .Y(_3429_)
);

AND2X2 _10151_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4]_5_bF$buf0 ),
    .Y(_3430_)
);

NAND2X1 _10152_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3429_),
    .B(_3430_),
    .Y(_3431_)
);

OAI21X1 _10153_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3277_),
    .B(_3262_),
    .C(_3346_),
    .Y(_3432_)
);

AOI21X1 _10154_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3432_),
    .B(_3431_),
    .C(_3428_),
    .Y(_3433_)
);

INVX1 _10155_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3428_),
    .Y(_3434_)
);

NAND2X1 _10156_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3346_),
    .B(_3430_),
    .Y(_3435_)
);

AOI22X1 _10157_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [4]),
    .C(gnd),
    .D(\X[4]_5_bF$buf3 ),
    .Y(_3436_)
);

INVX1 _10158_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3436_),
    .Y(_3437_)
);

AOI21X1 _10159_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3435_),
    .B(_3437_),
    .C(_3434_),
    .Y(_3438_)
);

OAI21X1 _10160_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3438_),
    .B(_3433_),
    .C(_3427_),
    .Y(_3439_)
);

AOI22X1 _10161_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3275_),
    .B(_3346_),
    .C(_3349_),
    .D(_3345_),
    .Y(_3440_)
);

NAND3X1 _10162_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3434_),
    .B(_3437_),
    .C(_3435_),
    .Y(_3441_)
);

NAND2X1 _10163_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4]_5_bF$buf2 ),
    .Y(_3442_)
);

NOR2X1 _10164_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3429_),
    .B(_3442_),
    .Y(_3443_)
);

OAI21X1 _10165_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3436_),
    .B(_3443_),
    .C(_3428_),
    .Y(_3444_)
);

NAND3X1 _10166_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3441_),
    .B(_3440_),
    .C(_3444_),
    .Y(_3445_)
);

AOI21X1 _10167_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3439_),
    .B(_3445_),
    .C(_3426_),
    .Y(_3446_)
);

AND2X2 _10168_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3425_),
    .B(_3420_),
    .Y(_3447_)
);

NAND3X1 _10169_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3427_),
    .B(_3441_),
    .C(_3444_),
    .Y(_3448_)
);

OAI21X1 _10170_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3438_),
    .B(_3433_),
    .C(_3440_),
    .Y(_3449_)
);

AOI21X1 _10171_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3449_),
    .B(_3448_),
    .C(_3447_),
    .Y(_3450_)
);

OAI21X1 _10172_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3446_),
    .B(_3450_),
    .C(_3412_),
    .Y(_3451_)
);

INVX1 _10173_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3355_),
    .Y(_3452_)
);

AOI21X1 _10174_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3340_),
    .B(_3359_),
    .C(_3452_),
    .Y(_3453_)
);

NAND3X1 _10175_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3448_),
    .B(_3447_),
    .C(_3449_),
    .Y(_3454_)
);

NAND3X1 _10176_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3426_),
    .B(_3445_),
    .C(_3439_),
    .Y(_3455_)
);

NAND3X1 _10177_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3454_),
    .B(_3455_),
    .C(_3453_),
    .Y(_3456_)
);

AOI21X1 _10178_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3456_),
    .B(_3451_),
    .C(_3410_),
    .Y(_3457_)
);

AND2X2 _10179_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3409_),
    .B(_3406_),
    .Y(_3458_)
);

NAND3X1 _10180_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3412_),
    .B(_3454_),
    .C(_3455_),
    .Y(_3459_)
);

OAI21X1 _10181_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3446_),
    .B(_3450_),
    .C(_3453_),
    .Y(_3460_)
);

AOI21X1 _10182_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3460_),
    .B(_3459_),
    .C(_3458_),
    .Y(_3461_)
);

OAI21X1 _10183_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3461_),
    .B(_3457_),
    .C(_3397_),
    .Y(_3462_)
);

INVX1 _10184_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3365_),
    .Y(_3463_)
);

AOI21X1 _10185_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3372_),
    .B(_3370_),
    .C(_3463_),
    .Y(_3464_)
);

NAND3X1 _10186_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3459_),
    .B(_3458_),
    .C(_3460_),
    .Y(_3465_)
);

NAND3X1 _10187_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3410_),
    .B(_3451_),
    .C(_3456_),
    .Y(_3466_)
);

NAND3X1 _10188_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3465_),
    .B(_3466_),
    .C(_3464_),
    .Y(_3467_)
);

AOI21X1 _10189_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3467_),
    .B(_3462_),
    .C(_3323_),
    .Y(_3468_)
);

INVX1 _10190_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3323_),
    .Y(_3469_)
);

NAND3X1 _10191_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3397_),
    .B(_3465_),
    .C(_3466_),
    .Y(_3470_)
);

OAI21X1 _10192_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3457_),
    .B(_3461_),
    .C(_3464_),
    .Y(_3471_)
);

AOI21X1 _10193_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3471_),
    .B(_3470_),
    .C(_3469_),
    .Y(_3472_)
);

OAI21X1 _10194_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3472_),
    .B(_3468_),
    .C(_3384_),
    .Y(_3473_)
);

NAND3X1 _10195_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3469_),
    .B(_3470_),
    .C(_3471_),
    .Y(_3474_)
);

NAND3X1 _10196_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3323_),
    .B(_3462_),
    .C(_3467_),
    .Y(_3475_)
);

NAND3X1 _10197_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3376_),
    .B(_3474_),
    .C(_3475_),
    .Y(_3476_)
);

AND2X2 _10198_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3473_),
    .B(_3476_),
    .Y(_3477_)
);

OAI21X1 _10199_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3395_),
    .B(_3392_),
    .C(_3477_),
    .Y(_3478_)
);

NOR2X1 _10200_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3395_),
    .B(_3392_),
    .Y(_3479_)
);

AOI21X1 _10201_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3475_),
    .B(_3474_),
    .C(_3376_),
    .Y(_3480_)
);

INVX1 _10202_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3476_),
    .Y(_3481_)
);

OAI21X1 _10203_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3480_),
    .B(_3481_),
    .C(_3479_),
    .Y(_3482_)
);

AND2X2 _10204_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3482_),
    .B(_3478_),
    .Y(_3984_[7])
);

NAND3X1 _10205_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3473_),
    .B(_3476_),
    .C(_3392_),
    .Y(_3483_)
);

AOI21X1 _10206_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3395_),
    .B(_3473_),
    .C(_3481_),
    .Y(_3484_)
);

NAND2X1 _10207_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3484_),
    .B(_3483_),
    .Y(_3485_)
);

INVX1 _10208_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3470_),
    .Y(_3486_)
);

AOI21X1 _10209_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3469_),
    .B(_3471_),
    .C(_3486_),
    .Y(_3487_)
);

OAI21X1 _10210_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3398_),
    .B(_3408_),
    .C(_3404_),
    .Y(_3488_)
);

INVX1 _10211_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3488_),
    .Y(_3489_)
);

AOI21X1 _10212_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3454_),
    .B(_3455_),
    .C(_3412_),
    .Y(_3490_)
);

OAI21X1 _10213_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3410_),
    .B(_3490_),
    .C(_3459_),
    .Y(_3491_)
);

NAND2X1 _10214_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [1]),
    .B(gnd),
    .Y(_3492_)
);

INVX2 _10215_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_3493_)
);

NOR2X1 _10216_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3958_),
    .B(_3493_),
    .Y(_3494_)
);

OAI21X1 _10217_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3413_),
    .B(_3418_),
    .C(_3417_),
    .Y(_3495_)
);

NOR2X1 _10218_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3494_),
    .B(_3495_),
    .Y(_3496_)
);

AND2X2 _10219_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3495_),
    .B(_3494_),
    .Y(_3497_)
);

OAI21X1 _10220_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3496_),
    .B(_3497_),
    .C(_3492_),
    .Y(_3498_)
);

INVX1 _10221_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3492_),
    .Y(_3499_)
);

OR2X2 _10222_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3495_),
    .B(_3494_),
    .Y(_3500_)
);

NAND2X1 _10223_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3494_),
    .B(_3495_),
    .Y(_3501_)
);

NAND3X1 _10224_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3499_),
    .B(_3501_),
    .C(_3500_),
    .Y(_3502_)
);

NAND2X1 _10225_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3498_),
    .B(_3502_),
    .Y(_3503_)
);

AOI21X1 _10226_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3444_),
    .B(_3441_),
    .C(_3427_),
    .Y(_3504_)
);

OAI21X1 _10227_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3426_),
    .B(_3504_),
    .C(_3448_),
    .Y(_3505_)
);

NAND2X1 _10228_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [3]),
    .B(gnd),
    .Y(_3506_)
);

INVX1 _10229_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .Y(_3507_)
);

OAI21X1 _10230_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3203_),
    .B(_3507_),
    .C(_3213_),
    .Y(_3508_)
);

NAND2X1 _10231_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [4]),
    .B(vdd),
    .Y(_3509_)
);

OAI21X1 _10232_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3506_),
    .B(_3509_),
    .C(_3508_),
    .Y(_3510_)
);

OAI21X1 _10233_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3428_),
    .B(_3436_),
    .C(_3435_),
    .Y(_3511_)
);

NAND2X1 _10234_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[4] [7]),
    .Y(_3512_)
);

NAND2X1 _10235_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4]_5_bF$buf1 ),
    .Y(_3513_)
);

NAND3X1 _10236_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [6]),
    .C(_3513_),
    .Y(_3514_)
);

AND2X2 _10237_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4]_5_bF$buf0 ),
    .Y(_3515_)
);

OAI21X1 _10238_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3277_),
    .B(_3332_),
    .C(_3515_),
    .Y(_3516_)
);

AOI21X1 _10239_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3516_),
    .B(_3514_),
    .C(_3512_),
    .Y(_3517_)
);

INVX1 _10240_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3512_),
    .Y(_3518_)
);

AND2X2 _10241_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [6]),
    .Y(_3519_)
);

NAND2X1 _10242_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3515_),
    .B(_3519_),
    .Y(_3520_)
);

NAND2X1 _10243_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [6]),
    .Y(_3521_)
);

NAND2X1 _10244_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3513_),
    .B(_3521_),
    .Y(_3522_)
);

AOI21X1 _10245_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3520_),
    .B(_3522_),
    .C(_3518_),
    .Y(_3523_)
);

OAI21X1 _10246_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3523_),
    .B(_3517_),
    .C(_3511_),
    .Y(_3524_)
);

AOI21X1 _10247_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3434_),
    .B(_3437_),
    .C(_3443_),
    .Y(_3525_)
);

NAND3X1 _10248_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3518_),
    .B(_3522_),
    .C(_3520_),
    .Y(_3526_)
);

NAND3X1 _10249_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3512_),
    .B(_3514_),
    .C(_3516_),
    .Y(_3527_)
);

NAND3X1 _10250_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3526_),
    .B(_3527_),
    .C(_3525_),
    .Y(_3528_)
);

AOI21X1 _10251_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3524_),
    .B(_3528_),
    .C(_3510_),
    .Y(_3529_)
);

INVX1 _10252_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3510_),
    .Y(_3530_)
);

NAND3X1 _10253_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3511_),
    .B(_3526_),
    .C(_3527_),
    .Y(_3531_)
);

OAI21X1 _10254_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3523_),
    .B(_3517_),
    .C(_3525_),
    .Y(_3532_)
);

AOI21X1 _10255_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3532_),
    .B(_3531_),
    .C(_3530_),
    .Y(_3533_)
);

OAI21X1 _10256_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3529_),
    .B(_3533_),
    .C(_3505_),
    .Y(_3534_)
);

INVX1 _10257_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3448_),
    .Y(_3535_)
);

AOI21X1 _10258_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3447_),
    .B(_3449_),
    .C(_3535_),
    .Y(_3536_)
);

NAND3X1 _10259_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3530_),
    .B(_3531_),
    .C(_3532_),
    .Y(_3537_)
);

NAND3X1 _10260_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3510_),
    .B(_3528_),
    .C(_3524_),
    .Y(_3538_)
);

NAND3X1 _10261_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3537_),
    .B(_3538_),
    .C(_3536_),
    .Y(_3539_)
);

AOI21X1 _10262_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3539_),
    .B(_3534_),
    .C(_3503_),
    .Y(_3540_)
);

AND2X2 _10263_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3502_),
    .B(_3498_),
    .Y(_3541_)
);

NAND3X1 _10264_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3537_),
    .B(_3538_),
    .C(_3505_),
    .Y(_3542_)
);

OAI21X1 _10265_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3529_),
    .B(_3533_),
    .C(_3536_),
    .Y(_3543_)
);

AOI21X1 _10266_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3543_),
    .B(_3542_),
    .C(_3541_),
    .Y(_3544_)
);

OAI21X1 _10267_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3544_),
    .B(_3540_),
    .C(_3491_),
    .Y(_3545_)
);

INVX1 _10268_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3459_),
    .Y(_3546_)
);

AOI21X1 _10269_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3458_),
    .B(_3460_),
    .C(_3546_),
    .Y(_3547_)
);

NAND3X1 _10270_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3541_),
    .B(_3542_),
    .C(_3543_),
    .Y(_3548_)
);

NAND3X1 _10271_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3503_),
    .B(_3534_),
    .C(_3539_),
    .Y(_3549_)
);

NAND3X1 _10272_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3548_),
    .B(_3549_),
    .C(_3547_),
    .Y(_3550_)
);

AOI21X1 _10273_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3545_),
    .B(_3550_),
    .C(_3489_),
    .Y(_3551_)
);

NAND3X1 _10274_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3491_),
    .B(_3548_),
    .C(_3549_),
    .Y(_3552_)
);

OAI21X1 _10275_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3544_),
    .B(_3540_),
    .C(_3547_),
    .Y(_3553_)
);

AOI21X1 _10276_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3553_),
    .B(_3552_),
    .C(_3488_),
    .Y(_3554_)
);

OAI21X1 _10277_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3554_),
    .B(_3551_),
    .C(_3487_),
    .Y(_3555_)
);

AOI21X1 _10278_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3466_),
    .B(_3465_),
    .C(_3397_),
    .Y(_3556_)
);

OAI21X1 _10279_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3323_),
    .B(_3556_),
    .C(_3470_),
    .Y(_3557_)
);

NAND3X1 _10280_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3488_),
    .B(_3552_),
    .C(_3553_),
    .Y(_3558_)
);

NAND3X1 _10281_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3489_),
    .B(_3550_),
    .C(_3545_),
    .Y(_3559_)
);

NAND3X1 _10282_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3557_),
    .B(_3558_),
    .C(_3559_),
    .Y(_3560_)
);

NAND2X1 _10283_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3560_),
    .B(_3555_),
    .Y(_3561_)
);

NAND2X1 _10284_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3561_),
    .B(_3485_),
    .Y(_3562_)
);

OAI21X1 _10285_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3390_),
    .B(_3480_),
    .C(_3476_),
    .Y(_3563_)
);

AOI21X1 _10286_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3477_),
    .B(_3392_),
    .C(_3563_),
    .Y(_3564_)
);

AND2X2 _10287_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3555_),
    .B(_3560_),
    .Y(_3565_)
);

NAND2X1 _10288_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3565_),
    .B(_3564_),
    .Y(_3566_)
);

NAND2X1 _10289_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3562_),
    .B(_3566_),
    .Y(_3984_[8])
);

INVX1 _10290_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3560_),
    .Y(_3567_)
);

AOI21X1 _10291_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3485_),
    .B(_3555_),
    .C(_3567_),
    .Y(_3568_)
);

AOI21X1 _10292_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3549_),
    .B(_3548_),
    .C(_3491_),
    .Y(_3569_)
);

OAI21X1 _10293_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3489_),
    .B(_3569_),
    .C(_3552_),
    .Y(_3570_)
);

OAI21X1 _10294_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3492_),
    .B(_3496_),
    .C(_3501_),
    .Y(_3571_)
);

AOI21X1 _10295_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3537_),
    .B(_3538_),
    .C(_3505_),
    .Y(_3572_)
);

OAI21X1 _10296_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3503_),
    .B(_3572_),
    .C(_3542_),
    .Y(_3573_)
);

NAND2X1 _10297_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [2]),
    .B(gnd),
    .Y(_3574_)
);

NOR2X1 _10298_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3506_),
    .B(_3509_),
    .Y(_3575_)
);

NAND2X1 _10299_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_3575_),
    .Y(_3576_)
);

INVX1 _10300_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3576_),
    .Y(_3577_)
);

AOI21X1 _10301_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [3]),
    .B(gnd),
    .C(_3575_),
    .Y(_3578_)
);

OAI21X1 _10302_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3578_),
    .B(_3577_),
    .C(_3574_),
    .Y(_3579_)
);

INVX1 _10303_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3574_),
    .Y(_3580_)
);

INVX1 _10304_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3578_),
    .Y(_3581_)
);

NAND3X1 _10305_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3580_),
    .B(_3576_),
    .C(_3581_),
    .Y(_3582_)
);

AND2X2 _10306_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3582_),
    .B(_3579_),
    .Y(_3583_)
);

AOI21X1 _10307_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3527_),
    .B(_3526_),
    .C(_3511_),
    .Y(_3584_)
);

OAI21X1 _10308_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3510_),
    .B(_3584_),
    .C(_3531_),
    .Y(_3585_)
);

NOR2X1 _10309_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3320_),
    .B(_3509_),
    .Y(_3586_)
);

AND2X2 _10310_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3320_),
    .B(_3509_),
    .Y(_3587_)
);

NOR2X1 _10311_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3586_),
    .B(_3587_),
    .Y(_3588_)
);

NAND2X1 _10312_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [6]),
    .Y(_3589_)
);

AOI22X1 _10313_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4]_5_bF$buf3 ),
    .C(gnd),
    .D(\X[4] [6]),
    .Y(_3590_)
);

OAI22X1 _10314_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3442_),
    .B(_3589_),
    .C(_3512_),
    .D(_3590_),
    .Y(_3591_)
);

AOI22X1 _10315_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [6]),
    .C(gnd),
    .D(\X[4] [7]),
    .Y(_3592_)
);

AND2X2 _10316_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [7]),
    .Y(_3593_)
);

AOI21X1 _10317_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3519_),
    .B(_3593_),
    .C(_3592_),
    .Y(_3594_)
);

NAND2X1 _10318_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3594_),
    .B(_3591_),
    .Y(_3595_)
);

AND2X2 _10319_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [6]),
    .Y(_3596_)
);

AOI22X1 _10320_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3430_),
    .B(_3596_),
    .C(_3522_),
    .D(_3518_),
    .Y(_3597_)
);

NAND2X1 _10321_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [7]),
    .Y(_3598_)
);

NAND2X1 _10322_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3589_),
    .B(_3598_),
    .Y(_3599_)
);

NAND2X1 _10323_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [7]),
    .Y(_3600_)
);

OAI21X1 _10324_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3521_),
    .B(_3600_),
    .C(_3599_),
    .Y(_3601_)
);

NAND2X1 _10325_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3601_),
    .B(_3597_),
    .Y(_3602_)
);

NAND3X1 _10326_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3588_),
    .B(_3595_),
    .C(_3602_),
    .Y(_3603_)
);

NAND2X1 _10327_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4]_5_bF$buf2 ),
    .B(vdd),
    .Y(_3604_)
);

INVX1 _10328_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [4]),
    .Y(_3605_)
);

OAI21X1 _10329_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3605_),
    .B(_3507_),
    .C(_3320_),
    .Y(_3606_)
);

OAI21X1 _10330_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3213_),
    .B(_3604_),
    .C(_3606_),
    .Y(_3607_)
);

NAND2X1 _10331_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3591_),
    .B(_3601_),
    .Y(_3608_)
);

NAND2X1 _10332_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3594_),
    .B(_3597_),
    .Y(_3609_)
);

NAND3X1 _10333_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3607_),
    .B(_3608_),
    .C(_3609_),
    .Y(_3610_)
);

NAND3X1 _10334_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3603_),
    .B(_3610_),
    .C(_3585_),
    .Y(_3611_)
);

NAND2X1 _10335_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3603_),
    .B(_3610_),
    .Y(_3612_)
);

NAND3X1 _10336_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3531_),
    .B(_3537_),
    .C(_3612_),
    .Y(_3613_)
);

NAND3X1 _10337_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3583_),
    .B(_3611_),
    .C(_3613_),
    .Y(_3614_)
);

NAND2X1 _10338_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3579_),
    .B(_3582_),
    .Y(_3615_)
);

AOI21X1 _10339_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3531_),
    .B(_3537_),
    .C(_3612_),
    .Y(_3616_)
);

AOI21X1 _10340_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3603_),
    .B(_3610_),
    .C(_3585_),
    .Y(_3617_)
);

OAI21X1 _10341_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3617_),
    .B(_3616_),
    .C(_3615_),
    .Y(_3618_)
);

NAND3X1 _10342_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3614_),
    .B(_3618_),
    .C(_3573_),
    .Y(_3619_)
);

INVX1 _10343_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3542_),
    .Y(_3620_)
);

AOI21X1 _10344_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3541_),
    .B(_3543_),
    .C(_3620_),
    .Y(_3621_)
);

INVX1 _10345_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3614_),
    .Y(_3622_)
);

AOI21X1 _10346_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3613_),
    .B(_3611_),
    .C(_3583_),
    .Y(_3623_)
);

OAI21X1 _10347_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3623_),
    .B(_3622_),
    .C(_3621_),
    .Y(_3624_)
);

NAND3X1 _10348_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3571_),
    .B(_3619_),
    .C(_3624_),
    .Y(_3625_)
);

INVX1 _10349_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3571_),
    .Y(_3626_)
);

INVX1 _10350_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3619_),
    .Y(_3627_)
);

AOI21X1 _10351_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3618_),
    .B(_3614_),
    .C(_3573_),
    .Y(_3628_)
);

OAI21X1 _10352_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3628_),
    .B(_3627_),
    .C(_3626_),
    .Y(_3629_)
);

NAND3X1 _10353_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3570_),
    .B(_3625_),
    .C(_3629_),
    .Y(_3630_)
);

INVX1 _10354_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3552_),
    .Y(_3631_)
);

AOI21X1 _10355_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3488_),
    .B(_3553_),
    .C(_3631_),
    .Y(_3632_)
);

OAI21X1 _10356_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3623_),
    .B(_3622_),
    .C(_3573_),
    .Y(_3633_)
);

NAND3X1 _10357_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3614_),
    .B(_3618_),
    .C(_3621_),
    .Y(_3634_)
);

AOI21X1 _10358_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3634_),
    .B(_3633_),
    .C(_3626_),
    .Y(_3635_)
);

AOI21X1 _10359_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3624_),
    .B(_3619_),
    .C(_3571_),
    .Y(_3636_)
);

OAI21X1 _10360_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3635_),
    .B(_3636_),
    .C(_3632_),
    .Y(_3637_)
);

AND2X2 _10361_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3637_),
    .B(_3630_),
    .Y(_3638_)
);

OR2X2 _10362_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3568_),
    .B(_3638_),
    .Y(_3639_)
);

NAND2X1 _10363_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3638_),
    .B(_3568_),
    .Y(_3640_)
);

NAND2X1 _10364_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3640_),
    .B(_3639_),
    .Y(_3984_[9])
);

NAND2X1 _10365_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3630_),
    .B(_3637_),
    .Y(_3641_)
);

NOR2X1 _10366_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3561_),
    .B(_3641_),
    .Y(_3642_)
);

NAND2X1 _10367_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3642_),
    .B(_3485_),
    .Y(_3643_)
);

AOI21X1 _10368_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3629_),
    .B(_3625_),
    .C(_3570_),
    .Y(_3644_)
);

AOI21X1 _10369_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3560_),
    .B(_3630_),
    .C(_3644_),
    .Y(_3645_)
);

INVX1 _10370_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3645_),
    .Y(_3646_)
);

OAI21X1 _10371_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3626_),
    .B(_3628_),
    .C(_3619_),
    .Y(_3647_)
);

OAI21X1 _10372_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3574_),
    .B(_3578_),
    .C(_3576_),
    .Y(_3648_)
);

OAI21X1 _10373_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3615_),
    .B(_3617_),
    .C(_3611_),
    .Y(_3649_)
);

INVX2 _10374_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_3650_)
);

NOR3X1 _10375_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3493_),
    .B(_3320_),
    .C(_3509_),
    .Y(_3651_)
);

OAI22X1 _10376_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3605_),
    .B(_3493_),
    .C(_3213_),
    .D(_3604_),
    .Y(_3652_)
);

INVX1 _10377_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3652_),
    .Y(_3653_)
);

OAI22X1 _10378_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3203_),
    .B(_3650_),
    .C(_3651_),
    .D(_3653_),
    .Y(_3654_)
);

NOR2X1 _10379_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3203_),
    .B(_3650_),
    .Y(_3655_)
);

NAND2X1 _10380_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_3586_),
    .Y(_3656_)
);

NAND3X1 _10381_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3655_),
    .B(_3652_),
    .C(_3656_),
    .Y(_3657_)
);

AND2X2 _10382_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3654_),
    .B(_3657_),
    .Y(_3658_)
);

NOR2X1 _10383_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3594_),
    .B(_3591_),
    .Y(_3659_)
);

OAI21X1 _10384_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3607_),
    .B(_3659_),
    .C(_3595_),
    .Y(_3660_)
);

NAND2X1 _10385_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [6]),
    .Y(_3661_)
);

NOR2X1 _10386_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3661_),
    .B(_3604_),
    .Y(_3662_)
);

AND2X2 _10387_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3661_),
    .B(_3604_),
    .Y(_3663_)
);

OAI22X1 _10388_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3519_),
    .B(_3600_),
    .C(_3662_),
    .D(_3663_),
    .Y(_3664_)
);

AND2X2 _10389_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [6]),
    .Y(_3665_)
);

AND2X2 _10390_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4]_5_bF$buf1 ),
    .B(vdd),
    .Y(_3666_)
);

NAND2X1 _10391_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3665_),
    .B(_3666_),
    .Y(_3667_)
);

OAI21X1 _10392_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3262_),
    .B(_3507_),
    .C(_3661_),
    .Y(_3668_)
);

AOI21X1 _10393_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [6]),
    .C(_3600_),
    .Y(_3669_)
);

NAND3X1 _10394_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3668_),
    .B(_3669_),
    .C(_3667_),
    .Y(_3670_)
);

AND2X2 _10395_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3664_),
    .B(_3670_),
    .Y(_3671_)
);

NAND2X1 _10396_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3671_),
    .B(_3660_),
    .Y(_3672_)
);

NAND2X1 _10397_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3670_),
    .B(_3664_),
    .Y(_3673_)
);

NAND3X1 _10398_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3595_),
    .B(_3673_),
    .C(_3603_),
    .Y(_3674_)
);

NAND3X1 _10399_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3658_),
    .B(_3674_),
    .C(_3672_),
    .Y(_3675_)
);

NAND2X1 _10400_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3657_),
    .B(_3654_),
    .Y(_3676_)
);

NAND2X1 _10401_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3673_),
    .B(_3660_),
    .Y(_3677_)
);

NAND3X1 _10402_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3595_),
    .B(_3671_),
    .C(_3603_),
    .Y(_3678_)
);

NAND3X1 _10403_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3676_),
    .B(_3678_),
    .C(_3677_),
    .Y(_3679_)
);

NAND3X1 _10404_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3675_),
    .B(_3679_),
    .C(_3649_),
    .Y(_3680_)
);

NAND2X1 _10405_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3679_),
    .B(_3675_),
    .Y(_3681_)
);

NAND3X1 _10406_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3611_),
    .B(_3614_),
    .C(_3681_),
    .Y(_3682_)
);

NAND3X1 _10407_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3648_),
    .B(_3682_),
    .C(_3680_),
    .Y(_3683_)
);

INVX1 _10408_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3648_),
    .Y(_3684_)
);

NAND2X1 _10409_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3681_),
    .B(_3649_),
    .Y(_3685_)
);

AOI21X1 _10410_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3583_),
    .B(_3613_),
    .C(_3616_),
    .Y(_3686_)
);

AND2X2 _10411_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3675_),
    .B(_3679_),
    .Y(_3687_)
);

NAND2X1 _10412_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3686_),
    .B(_3687_),
    .Y(_3688_)
);

NAND3X1 _10413_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3684_),
    .B(_3685_),
    .C(_3688_),
    .Y(_3689_)
);

AOI21X1 _10414_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3683_),
    .B(_3689_),
    .C(_3647_),
    .Y(_3690_)
);

NAND2X1 _10415_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3683_),
    .B(_3689_),
    .Y(_3691_)
);

AOI21X1 _10416_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3619_),
    .B(_3625_),
    .C(_3691_),
    .Y(_3692_)
);

NOR2X1 _10417_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3690_),
    .B(_3692_),
    .Y(_3693_)
);

INVX1 _10418_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3693_),
    .Y(_3694_)
);

AOI21X1 _10419_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3643_),
    .B(_3646_),
    .C(_3694_),
    .Y(_3695_)
);

NAND2X1 _10420_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3565_),
    .B(_3638_),
    .Y(_3696_)
);

OAI21X1 _10421_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3696_),
    .B(_3564_),
    .C(_3646_),
    .Y(_3697_)
);

NOR2X1 _10422_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3693_),
    .B(_3697_),
    .Y(_3698_)
);

NOR2X1 _10423_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3695_),
    .B(_3698_),
    .Y(_3984_[10])
);

NAND3X1 _10424_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3683_),
    .B(_3689_),
    .C(_3647_),
    .Y(_3699_)
);

NAND2X1 _10425_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3693_),
    .B(_3697_),
    .Y(_3700_)
);

NOR2X1 _10426_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3681_),
    .B(_3686_),
    .Y(_3701_)
);

AOI21X1 _10427_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3648_),
    .B(_3682_),
    .C(_3701_),
    .Y(_3702_)
);

NAND2X1 _10428_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3656_),
    .B(_3657_),
    .Y(_3703_)
);

NAND2X1 _10429_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3672_),
    .B(_3675_),
    .Y(_3704_)
);

NOR3X1 _10430_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3493_),
    .B(_3661_),
    .C(_3604_),
    .Y(_3705_)
);

AOI22X1 _10431_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4]_5_bF$buf0 ),
    .B(gnd),
    .C(_3665_),
    .D(_3666_),
    .Y(_3706_)
);

OAI22X1 _10432_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3605_),
    .B(_3650_),
    .C(_3706_),
    .D(_3705_),
    .Y(_3707_)
);

NOR2X1 _10433_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3605_),
    .B(_3650_),
    .Y(_3708_)
);

NAND2X1 _10434_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_3662_),
    .Y(_3709_)
);

OAI21X1 _10435_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3262_),
    .B(_3493_),
    .C(_3667_),
    .Y(_3710_)
);

NAND3X1 _10436_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3708_),
    .B(_3709_),
    .C(_3710_),
    .Y(_3711_)
);

NAND2X1 _10437_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3707_),
    .B(_3711_),
    .Y(_3712_)
);

NAND2X1 _10438_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3519_),
    .B(_3593_),
    .Y(_3713_)
);

NAND2X1 _10439_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[4] [7]),
    .Y(_3714_)
);

OAI22X1 _10440_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3421_),
    .B(_3423_),
    .C(_3507_),
    .D(_3332_),
    .Y(_3715_)
);

OAI21X1 _10441_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3661_),
    .B(_3714_),
    .C(_3715_),
    .Y(_3716_)
);

NAND3X1 _10442_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3713_),
    .B(_3716_),
    .C(_3670_),
    .Y(_3717_)
);

INVX1 _10443_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3717_),
    .Y(_3718_)
);

AOI21X1 _10444_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3670_),
    .B(_3713_),
    .C(_3716_),
    .Y(_3719_)
);

OAI21X1 _10445_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3719_),
    .B(_3718_),
    .C(_3712_),
    .Y(_3720_)
);

AND2X2 _10446_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3711_),
    .B(_3707_),
    .Y(_3721_)
);

INVX1 _10447_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3719_),
    .Y(_3722_)
);

NAND3X1 _10448_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3717_),
    .B(_3722_),
    .C(_3721_),
    .Y(_3723_)
);

AND2X2 _10449_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3723_),
    .B(_3720_),
    .Y(_3724_)
);

NAND2X1 _10450_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3724_),
    .B(_3704_),
    .Y(_3725_)
);

AOI21X1 _10451_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3603_),
    .B(_3595_),
    .C(_3673_),
    .Y(_3726_)
);

AOI21X1 _10452_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3658_),
    .B(_3674_),
    .C(_3726_),
    .Y(_3727_)
);

NAND2X1 _10453_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3720_),
    .B(_3723_),
    .Y(_3728_)
);

NAND2X1 _10454_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3728_),
    .B(_3727_),
    .Y(_3729_)
);

NAND3X1 _10455_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3703_),
    .B(_3729_),
    .C(_3725_),
    .Y(_3730_)
);

INVX1 _10456_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3703_),
    .Y(_3731_)
);

NAND2X1 _10457_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3728_),
    .B(_3704_),
    .Y(_3732_)
);

NAND2X1 _10458_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3727_),
    .B(_3724_),
    .Y(_3733_)
);

NAND3X1 _10459_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3731_),
    .B(_3733_),
    .C(_3732_),
    .Y(_3734_)
);

NAND2X1 _10460_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3730_),
    .B(_3734_),
    .Y(_3735_)
);

NAND2X1 _10461_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3735_),
    .B(_3702_),
    .Y(_3736_)
);

AOI21X1 _10462_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3675_),
    .B(_3679_),
    .C(_3649_),
    .Y(_3737_)
);

OAI21X1 _10463_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3684_),
    .B(_3737_),
    .C(_3680_),
    .Y(_3738_)
);

NAND3X1 _10464_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3730_),
    .B(_3734_),
    .C(_3738_),
    .Y(_3739_)
);

NAND2X1 _10465_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3736_),
    .B(_3739_),
    .Y(_3740_)
);

INVX1 _10466_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3740_),
    .Y(_3741_)
);

NAND3X1 _10467_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3699_),
    .B(_3741_),
    .C(_3700_),
    .Y(_3742_)
);

OAI21X1 _10468_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3692_),
    .B(_3695_),
    .C(_3740_),
    .Y(_3743_)
);

NAND2X1 _10469_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3742_),
    .B(_3743_),
    .Y(_3984_[11])
);

NOR3X1 _10470_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3690_),
    .B(_3692_),
    .C(_3740_),
    .Y(_3744_)
);

NAND3X1 _10471_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3642_),
    .B(_3744_),
    .C(_3485_),
    .Y(_3745_)
);

OAI21X1 _10472_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3699_),
    .B(_3740_),
    .C(_3739_),
    .Y(_3746_)
);

AOI21X1 _10473_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3744_),
    .B(_3645_),
    .C(_3746_),
    .Y(_3747_)
);

AND2X2 _10474_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3730_),
    .B(_3725_),
    .Y(_3748_)
);

OAI21X1 _10475_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3493_),
    .B(_3667_),
    .C(_3711_),
    .Y(_3749_)
);

OAI21X1 _10476_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3718_),
    .B(_3712_),
    .C(_3722_),
    .Y(_3750_)
);

INVX1 _10477_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3750_),
    .Y(_3751_)
);

INVX1 _10478_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3714_),
    .Y(_3752_)
);

NOR2X1 _10479_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3262_),
    .B(_3650_),
    .Y(_3753_)
);

NOR2X1 _10480_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3661_),
    .B(_3714_),
    .Y(_3754_)
);

NOR2X1 _10481_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3332_),
    .B(_3493_),
    .Y(_3755_)
);

NOR2X1 _10482_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3755_),
    .B(_3754_),
    .Y(_3756_)
);

AOI21X1 _10483_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_3754_),
    .C(_3756_),
    .Y(_3757_)
);

OR2X2 _10484_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3757_),
    .B(_3753_),
    .Y(_3758_)
);

NAND2X1 _10485_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3753_),
    .B(_3757_),
    .Y(_3759_)
);

NAND3X1 _10486_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3752_),
    .B(_3759_),
    .C(_3758_),
    .Y(_3760_)
);

NOR2X1 _10487_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3753_),
    .B(_3757_),
    .Y(_3761_)
);

INVX1 _10488_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3759_),
    .Y(_3762_)
);

OAI21X1 _10489_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3761_),
    .B(_3762_),
    .C(_3714_),
    .Y(_3763_)
);

NAND2X1 _10490_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3760_),
    .B(_3763_),
    .Y(_3764_)
);

NAND2X1 _10491_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3751_),
    .B(_3764_),
    .Y(_3765_)
);

NAND3X1 _10492_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3750_),
    .B(_3760_),
    .C(_3763_),
    .Y(_3766_)
);

AOI21X1 _10493_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3765_),
    .B(_3766_),
    .C(_3749_),
    .Y(_3767_)
);

NAND3X1 _10494_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3749_),
    .B(_3766_),
    .C(_3765_),
    .Y(_3768_)
);

INVX1 _10495_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3768_),
    .Y(_3769_)
);

OAI21X1 _10496_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3767_),
    .B(_3769_),
    .C(_3748_),
    .Y(_3770_)
);

OR2X2 _10497_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3769_),
    .B(_3767_),
    .Y(_3771_)
);

OR2X2 _10498_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3771_),
    .B(_3748_),
    .Y(_3772_)
);

NAND2X1 _10499_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3770_),
    .B(_3772_),
    .Y(_3773_)
);

AOI21X1 _10500_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3745_),
    .B(_3747_),
    .C(_3773_),
    .Y(_3774_)
);

NAND3X1 _10501_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3565_),
    .B(_3638_),
    .C(_3744_),
    .Y(_3775_)
);

OAI21X1 _10502_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3564_),
    .B(_3775_),
    .C(_3747_),
    .Y(_3776_)
);

INVX1 _10503_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3773_),
    .Y(_3777_)
);

NOR2X1 _10504_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3777_),
    .B(_3776_),
    .Y(_3778_)
);

NOR2X1 _10505_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3774_),
    .B(_3778_),
    .Y(_3984_[12])
);

NOR2X1 _10506_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3748_),
    .B(_3771_),
    .Y(_3779_)
);

INVX1 _10507_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3754_),
    .Y(_3780_)
);

OAI21X1 _10508_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3493_),
    .B(_3780_),
    .C(_3759_),
    .Y(_3781_)
);

INVX1 _10509_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3781_),
    .Y(_3782_)
);

NOR2X1 _10510_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3423_),
    .B(_3650_),
    .Y(_3783_)
);

NAND2X1 _10511_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3755_),
    .B(_3783_),
    .Y(_3784_)
);

OAI22X1 _10512_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3332_),
    .B(_3650_),
    .C(_3493_),
    .D(_3423_),
    .Y(_3785_)
);

NAND2X1 _10513_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3785_),
    .B(_3784_),
    .Y(_3786_)
);

NAND2X1 _10514_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3786_),
    .B(_3760_),
    .Y(_3787_)
);

OR2X2 _10515_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3760_),
    .B(_3786_),
    .Y(_3788_)
);

NAND2X1 _10516_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3787_),
    .B(_3788_),
    .Y(_3789_)
);

NAND2X1 _10517_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3782_),
    .B(_3789_),
    .Y(_3790_)
);

OR2X2 _10518_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3789_),
    .B(_3782_),
    .Y(_3791_)
);

NAND2X1 _10519_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3790_),
    .B(_3791_),
    .Y(_3792_)
);

NAND3X1 _10520_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3766_),
    .B(_3768_),
    .C(_3792_),
    .Y(_3793_)
);

OAI21X1 _10521_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3751_),
    .B(_3764_),
    .C(_3768_),
    .Y(_3794_)
);

AND2X2 _10522_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3791_),
    .B(_3790_),
    .Y(_3795_)
);

NAND2X1 _10523_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3794_),
    .B(_3795_),
    .Y(_3796_)
);

NAND2X1 _10524_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3793_),
    .B(_3796_),
    .Y(_3797_)
);

OAI21X1 _10525_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3779_),
    .B(_3774_),
    .C(_3797_),
    .Y(_3798_)
);

NAND2X1 _10526_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3777_),
    .B(_3776_),
    .Y(_3799_)
);

AND2X2 _10527_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3796_),
    .B(_3793_),
    .Y(_3800_)
);

NAND3X1 _10528_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3772_),
    .B(_3800_),
    .C(_3799_),
    .Y(_3801_)
);

NAND2X1 _10529_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3801_),
    .B(_3798_),
    .Y(_3984_[13])
);

NAND3X1 _10530_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3770_),
    .B(_3772_),
    .C(_3800_),
    .Y(_3802_)
);

AOI21X1 _10531_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3745_),
    .B(_3747_),
    .C(_3802_),
    .Y(_3803_)
);

OAI21X1 _10532_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3772_),
    .B(_3797_),
    .C(_3796_),
    .Y(_3804_)
);

OAI21X1 _10533_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3782_),
    .B(_3789_),
    .C(_3788_),
    .Y(_3805_)
);

AND2X2 _10534_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3784_),
    .B(_3783_),
    .Y(_3806_)
);

OR2X2 _10535_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3805_),
    .B(_3806_),
    .Y(_3807_)
);

NAND2X1 _10536_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3806_),
    .B(_3805_),
    .Y(_3808_)
);

NAND2X1 _10537_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3808_),
    .B(_3807_),
    .Y(_3809_)
);

OAI21X1 _10538_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3804_),
    .B(_3803_),
    .C(_3809_),
    .Y(_3810_)
);

INVX1 _10539_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3770_),
    .Y(_3811_)
);

NOR3X1 _10540_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3811_),
    .B(_3779_),
    .C(_3797_),
    .Y(_3812_)
);

NAND2X1 _10541_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3812_),
    .B(_3776_),
    .Y(_3813_)
);

INVX1 _10542_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3804_),
    .Y(_3814_)
);

INVX1 _10543_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3809_),
    .Y(_3815_)
);

NAND3X1 _10544_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3814_),
    .B(_3815_),
    .C(_3813_),
    .Y(_3816_)
);

NAND2X1 _10545_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3816_),
    .B(_3810_),
    .Y(_3984_[14])
);

OAI21X1 _10546_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3804_),
    .B(_3803_),
    .C(_3815_),
    .Y(_3817_)
);

OAI21X1 _10547_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3755_),
    .B(_3805_),
    .C(_3783_),
    .Y(_3818_)
);

NAND2X1 _10548_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3818_),
    .B(_3817_),
    .Y(_3984_[15])
);

INVX1 _10549_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3212_),
    .Y(_3979_[0])
);

AND2X2 _10550_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [0]),
    .B(\u_fir_pe4.mul [0]),
    .Y(_3819_)
);

INVX1 _10551_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [1]),
    .Y(_3820_)
);

INVX1 _10552_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.mul [1]),
    .Y(_3821_)
);

NOR2X1 _10553_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3820_),
    .B(_3821_),
    .Y(_3822_)
);

NOR2X1 _10554_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [1]),
    .B(\u_fir_pe4.mul [1]),
    .Y(_3823_)
);

NOR2X1 _10555_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3823_),
    .B(_3822_),
    .Y(_3824_)
);

NAND2X1 _10556_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3819_),
    .B(_3824_),
    .Y(_3825_)
);

INVX1 _10557_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3825_),
    .Y(_3826_)
);

NOR2X1 _10558_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3819_),
    .B(_3824_),
    .Y(_3827_)
);

NOR2X1 _10559_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3827_),
    .B(_3826_),
    .Y(_3978_[1])
);

OAI21X1 _10560_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3820_),
    .B(_3821_),
    .C(_3825_),
    .Y(_3828_)
);

AND2X2 _10561_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [2]),
    .B(\u_fir_pe4.mul [2]),
    .Y(_3829_)
);

NOR2X1 _10562_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [2]),
    .B(\u_fir_pe4.mul [2]),
    .Y(_3830_)
);

OAI21X1 _10563_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3829_),
    .B(_3830_),
    .C(_3828_),
    .Y(_3831_)
);

INVX1 _10564_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3828_),
    .Y(_3832_)
);

NOR2X1 _10565_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3830_),
    .B(_3829_),
    .Y(_3833_)
);

NAND2X1 _10566_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3833_),
    .B(_3832_),
    .Y(_3834_)
);

NAND2X1 _10567_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3831_),
    .B(_3834_),
    .Y(_3978_[2])
);

AOI21X1 _10568_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3828_),
    .B(_3833_),
    .C(_3829_),
    .Y(_3835_)
);

INVX1 _10569_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [3]),
    .Y(_3836_)
);

INVX1 _10570_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.mul [3]),
    .Y(_3837_)
);

NOR2X1 _10571_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3836_),
    .B(_3837_),
    .Y(_3838_)
);

NOR2X1 _10572_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [3]),
    .B(\u_fir_pe4.mul [3]),
    .Y(_3839_)
);

NOR2X1 _10573_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3839_),
    .B(_3838_),
    .Y(_3840_)
);

NAND2X1 _10574_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3840_),
    .B(_3835_),
    .Y(_3841_)
);

OR2X2 _10575_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3835_),
    .B(_3840_),
    .Y(_3842_)
);

NAND2X1 _10576_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3841_),
    .B(_3842_),
    .Y(_3978_[3])
);

INVX1 _10577_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [4]),
    .Y(_3843_)
);

INVX1 _10578_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.mul [4]),
    .Y(_3844_)
);

NOR2X1 _10579_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3843_),
    .B(_3844_),
    .Y(_3845_)
);

NOR2X1 _10580_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [4]),
    .B(\u_fir_pe4.mul [4]),
    .Y(_3846_)
);

NOR2X1 _10581_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3846_),
    .B(_3845_),
    .Y(_3847_)
);

INVX1 _10582_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3838_),
    .Y(_3848_)
);

OAI21X1 _10583_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3839_),
    .B(_3835_),
    .C(_3848_),
    .Y(_3849_)
);

NAND2X1 _10584_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3847_),
    .B(_3849_),
    .Y(_3850_)
);

OR2X2 _10585_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3849_),
    .B(_3847_),
    .Y(_3851_)
);

AND2X2 _10586_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3851_),
    .B(_3850_),
    .Y(_3978_[4])
);

OAI21X1 _10587_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3843_),
    .B(_3844_),
    .C(_3850_),
    .Y(_3852_)
);

INVX1 _10588_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [5]),
    .Y(_3853_)
);

INVX1 _10589_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.mul [5]),
    .Y(_3854_)
);

NOR2X1 _10590_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3853_),
    .B(_3854_),
    .Y(_3855_)
);

NOR2X1 _10591_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [5]),
    .B(\u_fir_pe4.mul [5]),
    .Y(_3856_)
);

NOR2X1 _10592_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3856_),
    .B(_3855_),
    .Y(_3857_)
);

NAND2X1 _10593_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3857_),
    .B(_3852_),
    .Y(_3858_)
);

OR2X2 _10594_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3852_),
    .B(_3857_),
    .Y(_3859_)
);

AND2X2 _10595_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3859_),
    .B(_3858_),
    .Y(_3978_[5])
);

OAI21X1 _10596_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3853_),
    .B(_3854_),
    .C(_3858_),
    .Y(_3860_)
);

INVX1 _10597_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [6]),
    .Y(_3861_)
);

INVX1 _10598_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.mul [6]),
    .Y(_3862_)
);

NOR2X1 _10599_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3861_),
    .B(_3862_),
    .Y(_3863_)
);

NOR2X1 _10600_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [6]),
    .B(\u_fir_pe4.mul [6]),
    .Y(_3864_)
);

NOR2X1 _10601_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3864_),
    .B(_3863_),
    .Y(_3865_)
);

NAND2X1 _10602_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3865_),
    .B(_3860_),
    .Y(_3866_)
);

OR2X2 _10603_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3860_),
    .B(_3865_),
    .Y(_3867_)
);

AND2X2 _10604_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3867_),
    .B(_3866_),
    .Y(_3978_[6])
);

OAI21X1 _10605_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3861_),
    .B(_3862_),
    .C(_3866_),
    .Y(_3868_)
);

INVX1 _10606_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [7]),
    .Y(_3869_)
);

INVX1 _10607_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.mul [7]),
    .Y(_3870_)
);

NOR2X1 _10608_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3869_),
    .B(_3870_),
    .Y(_3871_)
);

NOR2X1 _10609_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [7]),
    .B(\u_fir_pe4.mul [7]),
    .Y(_3872_)
);

OAI21X1 _10610_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3871_),
    .B(_3872_),
    .C(_3868_),
    .Y(_3873_)
);

INVX1 _10611_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3868_),
    .Y(_3874_)
);

NOR2X1 _10612_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3872_),
    .B(_3871_),
    .Y(_3875_)
);

NAND2X1 _10613_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3875_),
    .B(_3874_),
    .Y(_3876_)
);

NAND2X1 _10614_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3873_),
    .B(_3876_),
    .Y(_3978_[7])
);

INVX1 _10615_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [8]),
    .Y(_3878_)
);

INVX1 _10616_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.mul [8]),
    .Y(_3879_)
);

NOR2X1 _10617_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3878_),
    .B(_3879_),
    .Y(_3880_)
);

NOR2X1 _10618_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [8]),
    .B(\u_fir_pe4.mul [8]),
    .Y(_3881_)
);

NAND2X1 _10619_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3845_),
    .B(_3857_),
    .Y(_3882_)
);

OAI21X1 _10620_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3853_),
    .B(_3854_),
    .C(_3882_),
    .Y(_3883_)
);

NAND2X1 _10621_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3863_),
    .B(_3875_),
    .Y(_3884_)
);

OAI21X1 _10622_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3869_),
    .B(_3870_),
    .C(_3884_),
    .Y(_3885_)
);

AND2X2 _10623_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3865_),
    .B(_3875_),
    .Y(_3886_)
);

AOI21X1 _10624_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3883_),
    .B(_3886_),
    .C(_3885_),
    .Y(_3887_)
);

AND2X2 _10625_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3847_),
    .B(_3857_),
    .Y(_3889_)
);

NAND3X1 _10626_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3889_),
    .B(_3886_),
    .C(_3849_),
    .Y(_3890_)
);

NAND2X1 _10627_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3887_),
    .B(_3890_),
    .Y(_3891_)
);

OAI21X1 _10628_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3880_),
    .B(_3881_),
    .C(_3891_),
    .Y(_3892_)
);

NOR2X1 _10629_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3881_),
    .B(_3880_),
    .Y(_3893_)
);

INVX1 _10630_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3891_),
    .Y(_3894_)
);

NAND2X1 _10631_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3893_),
    .B(_3894_),
    .Y(_3895_)
);

NAND2X1 _10632_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3892_),
    .B(_3895_),
    .Y(_3978_[8])
);

INVX1 _10633_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3880_),
    .Y(_3896_)
);

INVX1 _10634_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3893_),
    .Y(_3897_)
);

OAI21X1 _10635_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3897_),
    .B(_3894_),
    .C(_3896_),
    .Y(_3899_)
);

AND2X2 _10636_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [9]),
    .B(\u_fir_pe4.mul [9]),
    .Y(_3900_)
);

NOR2X1 _10637_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [9]),
    .B(\u_fir_pe4.mul [9]),
    .Y(_3901_)
);

NOR2X1 _10638_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3901_),
    .B(_3900_),
    .Y(_3902_)
);

INVX1 _10639_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3902_),
    .Y(_3903_)
);

OR2X2 _10640_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3899_),
    .B(_3903_),
    .Y(_3904_)
);

OAI21X1 _10641_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3900_),
    .B(_3901_),
    .C(_3899_),
    .Y(_3905_)
);

NAND2X1 _10642_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3905_),
    .B(_3904_),
    .Y(_3978_[9])
);

NOR2X1 _10643_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3903_),
    .B(_3897_),
    .Y(_3906_)
);

AOI21X1 _10644_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3902_),
    .B(_3880_),
    .C(_3900_),
    .Y(_3907_)
);

INVX1 _10645_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3907_),
    .Y(_3909_)
);

AOI21X1 _10646_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3891_),
    .B(_3906_),
    .C(_3909_),
    .Y(_3910_)
);

INVX1 _10647_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3910_),
    .Y(_3911_)
);

INVX1 _10648_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [10]),
    .Y(_3912_)
);

INVX1 _10649_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.mul [10]),
    .Y(_3913_)
);

NOR2X1 _10650_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3912_),
    .B(_3913_),
    .Y(_3914_)
);

NOR2X1 _10651_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [10]),
    .B(\u_fir_pe4.mul [10]),
    .Y(_3915_)
);

NOR2X1 _10652_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3915_),
    .B(_3914_),
    .Y(_3916_)
);

NAND2X1 _10653_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3916_),
    .B(_3911_),
    .Y(_3917_)
);

OAI21X1 _10654_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3914_),
    .B(_3915_),
    .C(_3910_),
    .Y(_3918_)
);

AND2X2 _10655_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3917_),
    .B(_3918_),
    .Y(_3978_[10])
);

OAI21X1 _10656_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3912_),
    .B(_3913_),
    .C(_3917_),
    .Y(_3920_)
);

AND2X2 _10657_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [11]),
    .B(\u_fir_pe4.mul [11]),
    .Y(_3921_)
);

NOR2X1 _10658_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [11]),
    .B(\u_fir_pe4.mul [11]),
    .Y(_3922_)
);

NOR2X1 _10659_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3922_),
    .B(_3921_),
    .Y(_3923_)
);

NOR2X1 _10660_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3923_),
    .B(_3920_),
    .Y(_3924_)
);

AND2X2 _10661_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3920_),
    .B(_3923_),
    .Y(_3925_)
);

NOR2X1 _10662_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3924_),
    .B(_3925_),
    .Y(_3978_[11])
);

AOI21X1 _10663_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3923_),
    .B(_3914_),
    .C(_3921_),
    .Y(_3926_)
);

NAND2X1 _10664_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3923_),
    .B(_3916_),
    .Y(_3927_)
);

OAI21X1 _10665_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3927_),
    .B(_3910_),
    .C(_3926_),
    .Y(_3929_)
);

INVX1 _10666_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [12]),
    .Y(_3930_)
);

INVX1 _10667_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.mul [12]),
    .Y(_3931_)
);

NOR2X1 _10668_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3930_),
    .B(_3931_),
    .Y(_3932_)
);

NOR2X1 _10669_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [12]),
    .B(\u_fir_pe4.mul [12]),
    .Y(_3933_)
);

NOR2X1 _10670_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3933_),
    .B(_3932_),
    .Y(_3934_)
);

NAND2X1 _10671_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3934_),
    .B(_3929_),
    .Y(_3935_)
);

OR2X2 _10672_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3929_),
    .B(_3934_),
    .Y(_3936_)
);

AND2X2 _10673_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3936_),
    .B(_3935_),
    .Y(_3978_[12])
);

OAI21X1 _10674_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3930_),
    .B(_3931_),
    .C(_3935_),
    .Y(_3937_)
);

INVX1 _10675_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [13]),
    .Y(_3939_)
);

INVX1 _10676_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.mul [13]),
    .Y(_3940_)
);

NOR2X1 _10677_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3939_),
    .B(_3940_),
    .Y(_3941_)
);

NOR2X1 _10678_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [13]),
    .B(\u_fir_pe4.mul [13]),
    .Y(_3942_)
);

NOR2X1 _10679_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3942_),
    .B(_3941_),
    .Y(_3943_)
);

NAND2X1 _10680_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3943_),
    .B(_3937_),
    .Y(_3944_)
);

OR2X2 _10681_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3937_),
    .B(_3943_),
    .Y(_3945_)
);

AND2X2 _10682_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3945_),
    .B(_3944_),
    .Y(_3978_[13])
);

OAI21X1 _10683_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3939_),
    .B(_3940_),
    .C(_3944_),
    .Y(_3946_)
);

INVX1 _10684_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [14]),
    .Y(_3947_)
);

INVX1 _10685_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.mul [14]),
    .Y(_3949_)
);

NOR2X1 _10686_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3947_),
    .B(_3949_),
    .Y(_3950_)
);

NOR2X1 _10687_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [14]),
    .B(\u_fir_pe4.mul [14]),
    .Y(_3951_)
);

NOR2X1 _10688_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3951_),
    .B(_3950_),
    .Y(_3952_)
);

AND2X2 _10689_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3946_),
    .B(_3952_),
    .Y(_3953_)
);

NOR2X1 _10690_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3952_),
    .B(_3946_),
    .Y(_3954_)
);

NOR2X1 _10691_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3954_),
    .B(_3953_),
    .Y(_3978_[14])
);

INVX1 _10692_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3950_),
    .Y(_3955_)
);

NAND2X1 _10693_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3952_),
    .B(_3946_),
    .Y(_3956_)
);

NAND2X1 _10694_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [15]),
    .B(\u_fir_pe4.mul [15]),
    .Y(_3957_)
);

OR2X2 _10695_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [15]),
    .B(\u_fir_pe4.mul [15]),
    .Y(_3959_)
);

NAND2X1 _10696_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3957_),
    .B(_3959_),
    .Y(_3960_)
);

INVX1 _10697_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3960_),
    .Y(_3961_)
);

NAND3X1 _10698_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3955_),
    .B(_3961_),
    .C(_3956_),
    .Y(_3962_)
);

OAI21X1 _10699_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3950_),
    .B(_3953_),
    .C(_3960_),
    .Y(_3963_)
);

NAND2X1 _10700_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3962_),
    .B(_3963_),
    .Y(_3978_[15])
);

NOR2X1 _10701_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe4.rYin [0]),
    .B(\u_fir_pe4.mul [0]),
    .Y(_3964_)
);

NOR2X1 _10702_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3964_),
    .B(_3819_),
    .Y(_3977_[0])
);

AOI21X1 _10703_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [0]),
    .B(vdd),
    .C(_3888_),
    .Y(_3965_)
);

NOR2X1 _10704_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3965_),
    .B(_3908_),
    .Y(_3980_[1])
);

NOR2X1 _10705_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3908_),
    .B(_3972_),
    .Y(_3967_)
);

NOR2X1 _10706_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3967_),
    .B(_3974_),
    .Y(_3981_[2])
);

DFFPOSX1 _10707_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf57),
    .D(_3977_[0]),
    .Q(\Y[5] [0])
);

DFFPOSX1 _10708_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf56),
    .D(_3978_[1]),
    .Q(\Y[5] [1])
);

DFFPOSX1 _10709_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf55),
    .D(_3978_[2]),
    .Q(\Y[5] [2])
);

DFFPOSX1 _10710_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf54),
    .D(_3978_[3]),
    .Q(\Y[5] [3])
);

DFFPOSX1 _10711_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf53),
    .D(_3978_[4]),
    .Q(\Y[5] [4])
);

DFFPOSX1 _10712_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf52),
    .D(_3978_[5]),
    .Q(\Y[5] [5])
);

DFFPOSX1 _10713_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf51),
    .D(_3978_[6]),
    .Q(\Y[5] [6])
);

DFFPOSX1 _10714_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf50),
    .D(_3978_[7]),
    .Q(\Y[5] [7])
);

DFFPOSX1 _10715_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf49),
    .D(_3978_[8]),
    .Q(\Y[5] [8])
);

DFFPOSX1 _10716_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf48),
    .D(_3978_[9]),
    .Q(\Y[5] [9])
);

DFFPOSX1 _10717_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf47),
    .D(_3978_[10]),
    .Q(\Y[5] [10])
);

DFFPOSX1 _10718_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf46),
    .D(_3978_[11]),
    .Q(\Y[5] [11])
);

DFFPOSX1 _10719_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf45),
    .D(_3978_[12]),
    .Q(\Y[5] [12])
);

DFFPOSX1 _10720_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf44),
    .D(_3978_[13]),
    .Q(\Y[5] [13])
);

DFFPOSX1 _10721_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf43),
    .D(_3978_[14]),
    .Q(\Y[5] [14])
);

DFFPOSX1 _10722_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf42),
    .D(_3978_[15]),
    .Q(\Y[5] [15])
);

DFFPOSX1 _10723_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf41),
    .D(\X[4] [0]),
    .Q(\X[5] [0])
);

DFFPOSX1 _10724_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf40),
    .D(\X[4] [1]),
    .Q(\X[5] [1])
);

DFFPOSX1 _10725_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf39),
    .D(\X[4] [2]),
    .Q(\X[5] [2])
);

DFFPOSX1 _10726_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf38),
    .D(\X[4] [3]),
    .Q(\X[5] [3])
);

DFFPOSX1 _10727_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf37),
    .D(\X[4] [4]),
    .Q(\X[5] [4])
);

DFFPOSX1 _10728_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf36),
    .D(\X[4]_5_bF$buf3 ),
    .Q(\X[5] [5])
);

DFFPOSX1 _10729_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf35),
    .D(\X[4] [6]),
    .Q(\X[5] [6])
);

DFFPOSX1 _10730_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf34),
    .D(\X[4] [7]),
    .Q(\X[5] [7])
);

DFFPOSX1 _10731_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf33),
    .D(\Y[4] [0]),
    .Q(\u_fir_pe4.rYin [0])
);

DFFPOSX1 _10732_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf32),
    .D(\Y[4] [1]),
    .Q(\u_fir_pe4.rYin [1])
);

DFFPOSX1 _10733_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf31),
    .D(\Y[4] [2]),
    .Q(\u_fir_pe4.rYin [2])
);

DFFPOSX1 _10734_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf30),
    .D(\Y[4] [3]),
    .Q(\u_fir_pe4.rYin [3])
);

DFFPOSX1 _10735_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf29),
    .D(\Y[4] [4]),
    .Q(\u_fir_pe4.rYin [4])
);

DFFPOSX1 _10736_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf28),
    .D(\Y[4] [5]),
    .Q(\u_fir_pe4.rYin [5])
);

DFFPOSX1 _10737_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf27),
    .D(\Y[4] [6]),
    .Q(\u_fir_pe4.rYin [6])
);

DFFPOSX1 _10738_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf26),
    .D(\Y[4] [7]),
    .Q(\u_fir_pe4.rYin [7])
);

DFFPOSX1 _10739_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf25),
    .D(\Y[4] [8]),
    .Q(\u_fir_pe4.rYin [8])
);

DFFPOSX1 _10740_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf24),
    .D(\Y[4] [9]),
    .Q(\u_fir_pe4.rYin [9])
);

DFFPOSX1 _10741_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf23),
    .D(\Y[4] [10]),
    .Q(\u_fir_pe4.rYin [10])
);

DFFPOSX1 _10742_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf22),
    .D(\Y[4] [11]),
    .Q(\u_fir_pe4.rYin [11])
);

DFFPOSX1 _10743_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf21),
    .D(\Y[4] [12]),
    .Q(\u_fir_pe4.rYin [12])
);

DFFPOSX1 _10744_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf20),
    .D(\Y[4] [13]),
    .Q(\u_fir_pe4.rYin [13])
);

DFFPOSX1 _10745_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf19),
    .D(\Y[4] [14]),
    .Q(\u_fir_pe4.rYin [14])
);

DFFPOSX1 _10746_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf18),
    .D(\Y[4] [15]),
    .Q(\u_fir_pe4.rYin [15])
);

DFFPOSX1 _10747_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf17),
    .D(_3979_[0]),
    .Q(\u_fir_pe4.mul [0])
);

DFFPOSX1 _10748_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf16),
    .D(_3980_[1]),
    .Q(\u_fir_pe4.mul [1])
);

DFFPOSX1 _10749_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf15),
    .D(_3981_[2]),
    .Q(\u_fir_pe4.mul [2])
);

DFFPOSX1 _10750_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf14),
    .D(_3982_[3]),
    .Q(\u_fir_pe4.mul [3])
);

DFFPOSX1 _10751_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf13),
    .D(_3983_[4]),
    .Q(\u_fir_pe4.mul [4])
);

DFFPOSX1 _10752_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf12),
    .D(_3984_[5]),
    .Q(\u_fir_pe4.mul [5])
);

DFFPOSX1 _10753_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf11),
    .D(_3984_[6]),
    .Q(\u_fir_pe4.mul [6])
);

DFFPOSX1 _10754_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf10),
    .D(_3984_[7]),
    .Q(\u_fir_pe4.mul [7])
);

DFFPOSX1 _10755_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf9),
    .D(_3984_[8]),
    .Q(\u_fir_pe4.mul [8])
);

DFFPOSX1 _10756_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf8),
    .D(_3984_[9]),
    .Q(\u_fir_pe4.mul [9])
);

DFFPOSX1 _10757_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf7),
    .D(_3984_[10]),
    .Q(\u_fir_pe4.mul [10])
);

DFFPOSX1 _10758_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_3984_[11]),
    .Q(\u_fir_pe4.mul [11])
);

DFFPOSX1 _10759_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_3984_[12]),
    .Q(\u_fir_pe4.mul [12])
);

DFFPOSX1 _10760_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_3984_[13]),
    .Q(\u_fir_pe4.mul [13])
);

DFFPOSX1 _10761_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_3984_[14]),
    .Q(\u_fir_pe4.mul [14])
);

DFFPOSX1 _10762_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_3984_[15]),
    .Q(\u_fir_pe4.mul [15])
);

NAND2X1 _10763_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [0]),
    .B(gnd),
    .Y(_4674_)
);

AND2X2 _10764_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [1]),
    .B(vdd),
    .Y(_4685_)
);

INVX1 _10765_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4685_),
    .Y(_4695_)
);

NOR2X1 _10766_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4674_),
    .B(_4695_),
    .Y(_4705_)
);

NAND2X1 _10767_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [1]),
    .Y(_4716_)
);

NOR2X1 _10768_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4674_),
    .B(_4716_),
    .Y(_4725_)
);

AOI22X1 _10769_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [0]),
    .B(gnd),
    .C(\X[5] [1]),
    .D(gnd),
    .Y(_4735_)
);

NOR2X1 _10770_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4735_),
    .B(_4725_),
    .Y(_4745_)
);

INVX1 _10771_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [2]),
    .Y(_4755_)
);

INVX2 _10772_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .Y(_4763_)
);

NOR2X1 _10773_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4755_),
    .B(_4763_),
    .Y(_4765_)
);

NAND2X1 _10774_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4765_),
    .B(_4745_),
    .Y(_4766_)
);

INVX1 _10775_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4766_),
    .Y(_4767_)
);

NOR2X1 _10776_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4765_),
    .B(_4745_),
    .Y(_4768_)
);

NOR2X1 _10777_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4768_),
    .B(_4767_),
    .Y(_4769_)
);

NAND2X1 _10778_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4705_),
    .B(_4769_),
    .Y(_4770_)
);

INVX1 _10779_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4770_),
    .Y(_4771_)
);

NAND2X1 _10780_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [3]),
    .Y(_4772_)
);

INVX1 _10781_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4772_),
    .Y(_4773_)
);

NAND2X1 _10782_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [2]),
    .Y(_3985_)
);

INVX1 _10783_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3985_),
    .Y(_3986_)
);

NAND2X1 _10784_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [0]),
    .Y(_3987_)
);

OR2X2 _10785_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4716_),
    .B(_3987_),
    .Y(_3988_)
);

AOI22X1 _10786_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [0]),
    .C(gnd),
    .D(\X[5] [1]),
    .Y(_3989_)
);

INVX1 _10787_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3989_),
    .Y(_3990_)
);

NAND3X1 _10788_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3986_),
    .B(_3990_),
    .C(_3988_),
    .Y(_3991_)
);

NOR2X1 _10789_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4716_),
    .B(_3987_),
    .Y(_3992_)
);

OAI21X1 _10790_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3989_),
    .B(_3992_),
    .C(_3985_),
    .Y(_3993_)
);

NAND3X1 _10791_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4725_),
    .B(_3993_),
    .C(_3991_),
    .Y(_3994_)
);

INVX1 _10792_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4725_),
    .Y(_3995_)
);

NAND3X1 _10793_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3985_),
    .B(_3990_),
    .C(_3988_),
    .Y(_3996_)
);

OAI21X1 _10794_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3989_),
    .B(_3992_),
    .C(_3986_),
    .Y(_3997_)
);

NAND3X1 _10795_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3995_),
    .B(_3997_),
    .C(_3996_),
    .Y(_3998_)
);

NAND3X1 _10796_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4773_),
    .B(_3998_),
    .C(_3994_),
    .Y(_3999_)
);

INVX2 _10797_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [3]),
    .Y(_4000_)
);

NAND2X1 _10798_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3998_),
    .B(_3994_),
    .Y(_4001_)
);

OAI21X1 _10799_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4763_),
    .B(_4000_),
    .C(_4001_),
    .Y(_4002_)
);

NAND2X1 _10800_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3999_),
    .B(_4002_),
    .Y(_4003_)
);

NAND2X1 _10801_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4766_),
    .B(_4003_),
    .Y(_4004_)
);

NAND3X1 _10802_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4767_),
    .B(_3999_),
    .C(_4002_),
    .Y(_4005_)
);

NAND3X1 _10803_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4005_),
    .B(_4771_),
    .C(_4004_),
    .Y(_4006_)
);

INVX1 _10804_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4006_),
    .Y(_4007_)
);

AOI21X1 _10805_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4004_),
    .B(_4005_),
    .C(_4771_),
    .Y(_4008_)
);

NOR2X1 _10806_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4008_),
    .B(_4007_),
    .Y(_4779_[3])
);

NAND2X1 _10807_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [0]),
    .B(vdd),
    .Y(_4009_)
);

NAND2X1 _10808_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [4]),
    .B(vdd),
    .Y(_4010_)
);

NOR2X1 _10809_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4009_),
    .B(_4010_),
    .Y(_4011_)
);

AOI22X1 _10810_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [0]),
    .B(vdd),
    .C(vdd),
    .D(\X[5] [4]),
    .Y(_4012_)
);

NOR2X1 _10811_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4012_),
    .B(_4011_),
    .Y(_4013_)
);

INVX1 _10812_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4013_),
    .Y(_4014_)
);

NAND2X1 _10813_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [0]),
    .B(gnd),
    .Y(_4015_)
);

NAND2X1 _10814_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [1]),
    .Y(_4016_)
);

OAI22X1 _10815_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4015_),
    .B(_4016_),
    .C(_3985_),
    .D(_3989_),
    .Y(_4017_)
);

NAND2X1 _10816_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [3]),
    .Y(_4018_)
);

INVX1 _10817_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4018_),
    .Y(_4019_)
);

AND2X2 _10818_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [1]),
    .Y(_4020_)
);

AND2X2 _10819_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [2]),
    .Y(_4021_)
);

NAND2X1 _10820_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4020_),
    .B(_4021_),
    .Y(_4022_)
);

AOI22X1 _10821_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [1]),
    .C(gnd),
    .D(\X[5] [2]),
    .Y(_4023_)
);

INVX1 _10822_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4023_),
    .Y(_4024_)
);

NAND3X1 _10823_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4019_),
    .B(_4024_),
    .C(_4022_),
    .Y(_4025_)
);

NAND3X1 _10824_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [2]),
    .C(_4016_),
    .Y(_4026_)
);

NAND2X1 _10825_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [2]),
    .Y(_4027_)
);

NAND3X1 _10826_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [1]),
    .C(_4027_),
    .Y(_4028_)
);

NAND3X1 _10827_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4018_),
    .B(_4026_),
    .C(_4028_),
    .Y(_4029_)
);

NAND3X1 _10828_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4017_),
    .B(_4029_),
    .C(_4025_),
    .Y(_4030_)
);

INVX1 _10829_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4017_),
    .Y(_4031_)
);

NAND2X1 _10830_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4029_),
    .B(_4025_),
    .Y(_4032_)
);

NAND2X1 _10831_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4031_),
    .B(_4032_),
    .Y(_4033_)
);

NAND3X1 _10832_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4014_),
    .B(_4030_),
    .C(_4033_),
    .Y(_4034_)
);

NAND2X1 _10833_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4017_),
    .B(_4032_),
    .Y(_4035_)
);

NAND3X1 _10834_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4025_),
    .B(_4029_),
    .C(_4031_),
    .Y(_4036_)
);

NAND3X1 _10835_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4013_),
    .B(_4036_),
    .C(_4035_),
    .Y(_4037_)
);

AOI22X1 _10836_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3994_),
    .B(_3999_),
    .C(_4034_),
    .D(_4037_),
    .Y(_4038_)
);

INVX1 _10837_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4038_),
    .Y(_4039_)
);

NAND2X1 _10838_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3994_),
    .B(_3999_),
    .Y(_4040_)
);

NAND2X1 _10839_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4034_),
    .B(_4037_),
    .Y(_4041_)
);

OR2X2 _10840_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4041_),
    .B(_4040_),
    .Y(_4042_)
);

NAND2X1 _10841_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4039_),
    .B(_4042_),
    .Y(_4043_)
);

OAI21X1 _10842_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4766_),
    .B(_4003_),
    .C(_4006_),
    .Y(_4044_)
);

OR2X2 _10843_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4044_),
    .B(_4043_),
    .Y(_4045_)
);

NAND3X1 _10844_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4013_),
    .B(_4030_),
    .C(_4033_),
    .Y(_4046_)
);

INVX1 _10845_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4030_),
    .Y(_4047_)
);

AOI21X1 _10846_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4025_),
    .B(_4029_),
    .C(_4017_),
    .Y(_4048_)
);

OAI21X1 _10847_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4048_),
    .B(_4047_),
    .C(_4014_),
    .Y(_4049_)
);

AOI21X1 _10848_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4046_),
    .B(_4049_),
    .C(_4040_),
    .Y(_4050_)
);

OAI21X1 _10849_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4038_),
    .B(_4050_),
    .C(_4044_),
    .Y(_4051_)
);

NAND2X1 _10850_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4051_),
    .B(_4045_),
    .Y(_4780_[4])
);

NOR2X1 _10851_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4006_),
    .B(_4043_),
    .Y(_4052_)
);

NOR3X1 _10852_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4038_),
    .B(_4005_),
    .C(_4050_),
    .Y(_4053_)
);

OAI21X1 _10853_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4014_),
    .B(_4048_),
    .C(_4030_),
    .Y(_4054_)
);

NAND2X1 _10854_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [0]),
    .B(gnd),
    .Y(_4055_)
);

INVX1 _10855_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4055_),
    .Y(_4056_)
);

AND2X2 _10856_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5]_5_bF$buf3 ),
    .Y(_4057_)
);

NAND2X1 _10857_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4685_),
    .B(_4057_),
    .Y(_4058_)
);

INVX2 _10858_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5]_5_bF$buf2 ),
    .Y(_4059_)
);

NAND2X1 _10859_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [1]),
    .B(vdd),
    .Y(_4060_)
);

OAI21X1 _10860_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4763_),
    .B(_4059_),
    .C(_4060_),
    .Y(_4061_)
);

NAND3X1 _10861_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4061_),
    .B(_4056_),
    .C(_4058_),
    .Y(_4062_)
);

NAND3X1 _10862_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5]_5_bF$buf1 ),
    .C(_4060_),
    .Y(_4063_)
);

NAND2X1 _10863_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5]_5_bF$buf0 ),
    .Y(_4064_)
);

NAND3X1 _10864_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [1]),
    .B(vdd),
    .C(_4064_),
    .Y(_4065_)
);

NAND3X1 _10865_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4055_),
    .B(_4063_),
    .C(_4065_),
    .Y(_4066_)
);

AND2X2 _10866_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4062_),
    .B(_4066_),
    .Y(_4067_)
);

NAND2X1 _10867_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [2]),
    .Y(_4068_)
);

OAI22X1 _10868_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4716_),
    .B(_4068_),
    .C(_4018_),
    .D(_4023_),
    .Y(_4069_)
);

NAND2X1 _10869_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [4]),
    .Y(_4070_)
);

INVX1 _10870_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4070_),
    .Y(_4071_)
);

AND2X2 _10871_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [3]),
    .Y(_4072_)
);

NAND2X1 _10872_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4021_),
    .B(_4072_),
    .Y(_4073_)
);

INVX1 _10873_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_4074_)
);

OAI21X1 _10874_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4074_),
    .B(_4000_),
    .C(_4068_),
    .Y(_4075_)
);

NAND3X1 _10875_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4071_),
    .B(_4075_),
    .C(_4073_),
    .Y(_4076_)
);

NAND3X1 _10876_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [3]),
    .C(_4068_),
    .Y(_4077_)
);

NAND2X1 _10877_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [3]),
    .Y(_4078_)
);

NAND3X1 _10878_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [2]),
    .C(_4078_),
    .Y(_4079_)
);

NAND3X1 _10879_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4070_),
    .B(_4077_),
    .C(_4079_),
    .Y(_4080_)
);

NAND3X1 _10880_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4069_),
    .B(_4080_),
    .C(_4076_),
    .Y(_4081_)
);

INVX1 _10881_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4069_),
    .Y(_4082_)
);

AOI21X1 _10882_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4077_),
    .B(_4079_),
    .C(_4070_),
    .Y(_4083_)
);

AOI22X1 _10883_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [4]),
    .C(_4073_),
    .D(_4075_),
    .Y(_4084_)
);

OAI21X1 _10884_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4083_),
    .B(_4084_),
    .C(_4082_),
    .Y(_4085_)
);

NAND3X1 _10885_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4081_),
    .B(_4067_),
    .C(_4085_),
    .Y(_4086_)
);

NAND2X1 _10886_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4066_),
    .B(_4062_),
    .Y(_4087_)
);

OAI21X1 _10887_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4083_),
    .B(_4084_),
    .C(_4069_),
    .Y(_4088_)
);

NAND3X1 _10888_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4080_),
    .B(_4076_),
    .C(_4082_),
    .Y(_4089_)
);

NAND3X1 _10889_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4087_),
    .B(_4089_),
    .C(_4088_),
    .Y(_4090_)
);

NAND3X1 _10890_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4086_),
    .B(_4090_),
    .C(_4054_),
    .Y(_4091_)
);

AOI21X1 _10891_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4013_),
    .B(_4033_),
    .C(_4047_),
    .Y(_4092_)
);

AOI21X1 _10892_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4088_),
    .B(_4089_),
    .C(_4087_),
    .Y(_4093_)
);

AOI21X1 _10893_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4085_),
    .B(_4081_),
    .C(_4067_),
    .Y(_4094_)
);

OAI21X1 _10894_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4093_),
    .B(_4094_),
    .C(_4092_),
    .Y(_4095_)
);

NAND3X1 _10895_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4011_),
    .B(_4091_),
    .C(_4095_),
    .Y(_4096_)
);

INVX1 _10896_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4011_),
    .Y(_4097_)
);

OAI21X1 _10897_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4093_),
    .B(_4094_),
    .C(_4054_),
    .Y(_4098_)
);

NAND3X1 _10898_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4086_),
    .B(_4090_),
    .C(_4092_),
    .Y(_4099_)
);

NAND3X1 _10899_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4097_),
    .B(_4098_),
    .C(_4099_),
    .Y(_4100_)
);

NAND3X1 _10900_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4038_),
    .B(_4096_),
    .C(_4100_),
    .Y(_4101_)
);

NAND3X1 _10901_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4097_),
    .B(_4091_),
    .C(_4095_),
    .Y(_4102_)
);

NAND3X1 _10902_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4011_),
    .B(_4098_),
    .C(_4099_),
    .Y(_4103_)
);

NAND3X1 _10903_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4039_),
    .B(_4102_),
    .C(_4103_),
    .Y(_4104_)
);

NAND3X1 _10904_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4101_),
    .B(_4104_),
    .C(_4053_),
    .Y(_4105_)
);

INVX1 _10905_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4005_),
    .Y(_4106_)
);

NAND3X1 _10906_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4106_),
    .B(_4039_),
    .C(_4042_),
    .Y(_4107_)
);

NAND3X1 _10907_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4039_),
    .B(_4096_),
    .C(_4100_),
    .Y(_4108_)
);

NAND3X1 _10908_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4038_),
    .B(_4102_),
    .C(_4103_),
    .Y(_4109_)
);

NAND3X1 _10909_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4108_),
    .B(_4109_),
    .C(_4107_),
    .Y(_4110_)
);

NAND3X1 _10910_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4105_),
    .B(_4110_),
    .C(_4052_),
    .Y(_4111_)
);

INVX1 _10911_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4052_),
    .Y(_4112_)
);

INVX1 _10912_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4105_),
    .Y(_4113_)
);

INVX1 _10913_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4110_),
    .Y(_4114_)
);

OAI21X1 _10914_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4113_),
    .B(_4114_),
    .C(_4112_),
    .Y(_4115_)
);

AND2X2 _10915_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4115_),
    .B(_4111_),
    .Y(_4781_[5])
);

AND2X2 _10916_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [0]),
    .B(gnd),
    .Y(_4116_)
);

NAND2X1 _10917_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5]_5_bF$buf3 ),
    .Y(_4117_)
);

OAI21X1 _10918_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4695_),
    .B(_4117_),
    .C(_4062_),
    .Y(_4118_)
);

OR2X2 _10919_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4118_),
    .B(_4116_),
    .Y(_4119_)
);

NAND2X1 _10920_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4116_),
    .B(_4118_),
    .Y(_4120_)
);

NAND2X1 _10921_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4120_),
    .B(_4119_),
    .Y(_4121_)
);

AOI21X1 _10922_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4076_),
    .B(_4080_),
    .C(_4069_),
    .Y(_4122_)
);

OAI21X1 _10923_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4087_),
    .B(_4122_),
    .C(_4081_),
    .Y(_4123_)
);

NAND2X1 _10924_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [1]),
    .B(gnd),
    .Y(_4124_)
);

INVX1 _10925_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4124_),
    .Y(_4125_)
);

AND2X2 _10926_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [2]),
    .B(vdd),
    .Y(_4126_)
);

AND2X2 _10927_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [6]),
    .Y(_4127_)
);

NAND2X1 _10928_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4126_),
    .B(_4127_),
    .Y(_4128_)
);

INVX2 _10929_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [6]),
    .Y(_4129_)
);

NAND2X1 _10930_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [2]),
    .B(vdd),
    .Y(_4130_)
);

OAI21X1 _10931_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4763_),
    .B(_4129_),
    .C(_4130_),
    .Y(_4131_)
);

NAND3X1 _10932_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4131_),
    .B(_4125_),
    .C(_4128_),
    .Y(_4132_)
);

NAND3X1 _10933_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [6]),
    .C(_4130_),
    .Y(_4133_)
);

NAND2X1 _10934_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [6]),
    .Y(_4134_)
);

NAND2X1 _10935_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4134_),
    .B(_4126_),
    .Y(_4135_)
);

NAND3X1 _10936_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4124_),
    .B(_4133_),
    .C(_4135_),
    .Y(_4136_)
);

AND2X2 _10937_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4132_),
    .B(_4136_),
    .Y(_4137_)
);

NAND2X1 _10938_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [3]),
    .Y(_4138_)
);

AOI22X1 _10939_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [2]),
    .C(gnd),
    .D(\X[5] [3]),
    .Y(_4139_)
);

OAI22X1 _10940_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4027_),
    .B(_4138_),
    .C(_4070_),
    .D(_4139_),
    .Y(_4140_)
);

NAND2X1 _10941_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5]_5_bF$buf2 ),
    .Y(_4141_)
);

INVX1 _10942_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4141_),
    .Y(_4142_)
);

AND2X2 _10943_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [4]),
    .Y(_4143_)
);

NAND2X1 _10944_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4072_),
    .B(_4143_),
    .Y(_4144_)
);

AOI22X1 _10945_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [3]),
    .C(gnd),
    .D(\X[5] [4]),
    .Y(_4145_)
);

INVX1 _10946_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4145_),
    .Y(_4146_)
);

NAND3X1 _10947_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4142_),
    .B(_4146_),
    .C(_4144_),
    .Y(_4147_)
);

NAND3X1 _10948_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [4]),
    .C(_4138_),
    .Y(_4148_)
);

NAND2X1 _10949_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [4]),
    .Y(_4149_)
);

NAND3X1 _10950_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [3]),
    .C(_4149_),
    .Y(_4150_)
);

NAND3X1 _10951_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4141_),
    .B(_4148_),
    .C(_4150_),
    .Y(_4151_)
);

NAND3X1 _10952_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4140_),
    .B(_4151_),
    .C(_4147_),
    .Y(_4152_)
);

INVX1 _10953_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4140_),
    .Y(_4153_)
);

AOI21X1 _10954_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4148_),
    .B(_4150_),
    .C(_4141_),
    .Y(_4154_)
);

AOI22X1 _10955_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5]_5_bF$buf1 ),
    .C(_4144_),
    .D(_4146_),
    .Y(_4155_)
);

OAI21X1 _10956_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4154_),
    .B(_4155_),
    .C(_4153_),
    .Y(_4156_)
);

NAND3X1 _10957_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4152_),
    .B(_4137_),
    .C(_4156_),
    .Y(_4157_)
);

NAND2X1 _10958_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4136_),
    .B(_4132_),
    .Y(_4158_)
);

OAI21X1 _10959_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4154_),
    .B(_4155_),
    .C(_4140_),
    .Y(_4159_)
);

NAND3X1 _10960_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4147_),
    .B(_4151_),
    .C(_4153_),
    .Y(_4160_)
);

NAND3X1 _10961_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4158_),
    .B(_4160_),
    .C(_4159_),
    .Y(_4161_)
);

NAND3X1 _10962_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4157_),
    .B(_4123_),
    .C(_4161_),
    .Y(_4162_)
);

INVX1 _10963_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4081_),
    .Y(_4163_)
);

AOI21X1 _10964_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4067_),
    .B(_4085_),
    .C(_4163_),
    .Y(_4164_)
);

AOI21X1 _10965_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4159_),
    .B(_4160_),
    .C(_4158_),
    .Y(_4165_)
);

AOI21X1 _10966_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4156_),
    .B(_4152_),
    .C(_4137_),
    .Y(_4166_)
);

OAI21X1 _10967_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4165_),
    .B(_4166_),
    .C(_4164_),
    .Y(_4167_)
);

NAND3X1 _10968_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4121_),
    .B(_4162_),
    .C(_4167_),
    .Y(_4168_)
);

AND2X2 _10969_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4119_),
    .B(_4120_),
    .Y(_4169_)
);

OAI21X1 _10970_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4165_),
    .B(_4166_),
    .C(_4123_),
    .Y(_4170_)
);

NAND3X1 _10971_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4157_),
    .B(_4161_),
    .C(_4164_),
    .Y(_4171_)
);

NAND3X1 _10972_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4169_),
    .B(_4170_),
    .C(_4171_),
    .Y(_4172_)
);

AOI22X1 _10973_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4096_),
    .B(_4091_),
    .C(_4168_),
    .D(_4172_),
    .Y(_4173_)
);

AOI21X1 _10974_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4086_),
    .B(_4090_),
    .C(_4054_),
    .Y(_4174_)
);

OAI21X1 _10975_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4097_),
    .B(_4174_),
    .C(_4091_),
    .Y(_4175_)
);

NAND3X1 _10976_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4169_),
    .B(_4162_),
    .C(_4167_),
    .Y(_4176_)
);

NAND3X1 _10977_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4121_),
    .B(_4170_),
    .C(_4171_),
    .Y(_4177_)
);

AOI21X1 _10978_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4177_),
    .B(_4176_),
    .C(_4175_),
    .Y(_4178_)
);

OAI21X1 _10979_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4178_),
    .B(_4173_),
    .C(_4101_),
    .Y(_4179_)
);

AOI21X1 _10980_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4103_),
    .B(_4102_),
    .C(_4039_),
    .Y(_4180_)
);

NAND3X1 _10981_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4175_),
    .B(_4176_),
    .C(_4177_),
    .Y(_4181_)
);

INVX1 _10982_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4091_),
    .Y(_4182_)
);

AOI21X1 _10983_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4011_),
    .B(_4095_),
    .C(_4182_),
    .Y(_4183_)
);

AOI21X1 _10984_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4171_),
    .B(_4170_),
    .C(_4121_),
    .Y(_4184_)
);

AOI21X1 _10985_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4167_),
    .B(_4162_),
    .C(_4169_),
    .Y(_4185_)
);

OAI21X1 _10986_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4184_),
    .B(_4185_),
    .C(_4183_),
    .Y(_4186_)
);

NAND3X1 _10987_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4180_),
    .B(_4181_),
    .C(_4186_),
    .Y(_4187_)
);

NAND2X1 _10988_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4187_),
    .B(_4179_),
    .Y(_4188_)
);

AOI21X1 _10989_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4105_),
    .B(_4111_),
    .C(_4188_),
    .Y(_4189_)
);

OAI21X1 _10990_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4114_),
    .B(_4112_),
    .C(_4105_),
    .Y(_4190_)
);

AOI21X1 _10991_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4179_),
    .B(_4187_),
    .C(_4190_),
    .Y(_4191_)
);

NOR2X1 _10992_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4189_),
    .B(_4191_),
    .Y(_4781_[6])
);

INVX1 _10993_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4187_),
    .Y(_4192_)
);

AOI21X1 _10994_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4157_),
    .B(_4161_),
    .C(_4123_),
    .Y(_4193_)
);

OAI21X1 _10995_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4121_),
    .B(_4193_),
    .C(_4162_),
    .Y(_4194_)
);

NAND2X1 _10996_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [0]),
    .B(gnd),
    .Y(_4195_)
);

INVX1 _10997_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4195_),
    .Y(_4196_)
);

NAND2X1 _10998_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [1]),
    .B(gnd),
    .Y(_4197_)
);

INVX1 _10999_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4197_),
    .Y(_4198_)
);

AND2X2 _11000_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4130_),
    .B(_4134_),
    .Y(_4199_)
);

OAI21X1 _11001_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4124_),
    .B(_4199_),
    .C(_4128_),
    .Y(_4200_)
);

NAND2X1 _11002_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4198_),
    .B(_4200_),
    .Y(_4201_)
);

NAND3X1 _11003_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4128_),
    .B(_4197_),
    .C(_4132_),
    .Y(_4202_)
);

NAND3X1 _11004_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4196_),
    .B(_4202_),
    .C(_4201_),
    .Y(_4203_)
);

AOI21X1 _11005_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4132_),
    .B(_4128_),
    .C(_4197_),
    .Y(_4204_)
);

NOR2X1 _11006_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4198_),
    .B(_4200_),
    .Y(_4205_)
);

OAI21X1 _11007_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4204_),
    .B(_4205_),
    .C(_4195_),
    .Y(_4206_)
);

NAND2X1 _11008_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4203_),
    .B(_4206_),
    .Y(_4207_)
);

AOI21X1 _11009_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4147_),
    .B(_4151_),
    .C(_4140_),
    .Y(_4208_)
);

OAI21X1 _11010_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4158_),
    .B(_4208_),
    .C(_4152_),
    .Y(_4209_)
);

NAND2X1 _11011_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [2]),
    .B(gnd),
    .Y(_4210_)
);

INVX1 _11012_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4210_),
    .Y(_4211_)
);

AND2X2 _11013_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [3]),
    .B(vdd),
    .Y(_4212_)
);

AND2X2 _11014_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [7]),
    .Y(_4213_)
);

NAND2X1 _11015_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4212_),
    .B(_4213_),
    .Y(_4214_)
);

AOI22X1 _11016_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [7]),
    .C(\X[5] [3]),
    .D(vdd),
    .Y(_4215_)
);

INVX1 _11017_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4215_),
    .Y(_4216_)
);

NAND3X1 _11018_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4211_),
    .B(_4216_),
    .C(_4214_),
    .Y(_4217_)
);

INVX1 _11019_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .Y(_4218_)
);

OAI21X1 _11020_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4000_),
    .B(_4218_),
    .C(_4213_),
    .Y(_4219_)
);

INVX1 _11021_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [7]),
    .Y(_4220_)
);

OAI21X1 _11022_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4763_),
    .B(_4220_),
    .C(_4212_),
    .Y(_4221_)
);

NAND3X1 _11023_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4210_),
    .B(_4219_),
    .C(_4221_),
    .Y(_4222_)
);

NAND2X1 _11024_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4217_),
    .B(_4222_),
    .Y(_4223_)
);

OAI21X1 _11025_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4141_),
    .B(_4145_),
    .C(_4144_),
    .Y(_4224_)
);

NAND2X1 _11026_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [6]),
    .Y(_4225_)
);

NAND2X1 _11027_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [4]),
    .Y(_4226_)
);

AND2X2 _11028_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5]_5_bF$buf0 ),
    .Y(_4227_)
);

NAND2X1 _11029_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4226_),
    .B(_4227_),
    .Y(_4228_)
);

OAI21X1 _11030_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4074_),
    .B(_4059_),
    .C(_4143_),
    .Y(_4229_)
);

AOI21X1 _11031_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4229_),
    .B(_4228_),
    .C(_4225_),
    .Y(_4230_)
);

INVX1 _11032_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4225_),
    .Y(_4231_)
);

NAND2X1 _11033_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4143_),
    .B(_4227_),
    .Y(_4232_)
);

AOI22X1 _11034_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [4]),
    .C(gnd),
    .D(\X[5]_5_bF$buf3 ),
    .Y(_4233_)
);

INVX1 _11035_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4233_),
    .Y(_4234_)
);

AOI21X1 _11036_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4232_),
    .B(_4234_),
    .C(_4231_),
    .Y(_4235_)
);

OAI21X1 _11037_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4235_),
    .B(_4230_),
    .C(_4224_),
    .Y(_4236_)
);

AOI22X1 _11038_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4072_),
    .B(_4143_),
    .C(_4146_),
    .D(_4142_),
    .Y(_4237_)
);

NAND3X1 _11039_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4231_),
    .B(_4234_),
    .C(_4232_),
    .Y(_4238_)
);

NAND2X1 _11040_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5]_5_bF$buf2 ),
    .Y(_4239_)
);

NOR2X1 _11041_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4226_),
    .B(_4239_),
    .Y(_4240_)
);

OAI21X1 _11042_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4233_),
    .B(_4240_),
    .C(_4225_),
    .Y(_4241_)
);

NAND3X1 _11043_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4238_),
    .B(_4237_),
    .C(_4241_),
    .Y(_4242_)
);

AOI21X1 _11044_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4236_),
    .B(_4242_),
    .C(_4223_),
    .Y(_4243_)
);

AND2X2 _11045_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4222_),
    .B(_4217_),
    .Y(_4244_)
);

NAND3X1 _11046_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4224_),
    .B(_4238_),
    .C(_4241_),
    .Y(_4245_)
);

OAI21X1 _11047_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4235_),
    .B(_4230_),
    .C(_4237_),
    .Y(_4246_)
);

AOI21X1 _11048_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4246_),
    .B(_4245_),
    .C(_4244_),
    .Y(_4247_)
);

OAI21X1 _11049_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4243_),
    .B(_4247_),
    .C(_4209_),
    .Y(_4248_)
);

INVX1 _11050_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4152_),
    .Y(_4249_)
);

AOI21X1 _11051_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4137_),
    .B(_4156_),
    .C(_4249_),
    .Y(_4250_)
);

NAND3X1 _11052_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4245_),
    .B(_4244_),
    .C(_4246_),
    .Y(_4251_)
);

NAND3X1 _11053_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4223_),
    .B(_4242_),
    .C(_4236_),
    .Y(_4252_)
);

NAND3X1 _11054_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4251_),
    .B(_4252_),
    .C(_4250_),
    .Y(_4253_)
);

AOI21X1 _11055_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4253_),
    .B(_4248_),
    .C(_4207_),
    .Y(_4254_)
);

AND2X2 _11056_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4206_),
    .B(_4203_),
    .Y(_4255_)
);

NAND3X1 _11057_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4209_),
    .B(_4251_),
    .C(_4252_),
    .Y(_4256_)
);

OAI21X1 _11058_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4243_),
    .B(_4247_),
    .C(_4250_),
    .Y(_4257_)
);

AOI21X1 _11059_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4257_),
    .B(_4256_),
    .C(_4255_),
    .Y(_4258_)
);

OAI21X1 _11060_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4258_),
    .B(_4254_),
    .C(_4194_),
    .Y(_4259_)
);

INVX1 _11061_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4162_),
    .Y(_4260_)
);

AOI21X1 _11062_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4169_),
    .B(_4167_),
    .C(_4260_),
    .Y(_4261_)
);

NAND3X1 _11063_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4256_),
    .B(_4255_),
    .C(_4257_),
    .Y(_4262_)
);

NAND3X1 _11064_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4207_),
    .B(_4248_),
    .C(_4253_),
    .Y(_4263_)
);

NAND3X1 _11065_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4262_),
    .B(_4263_),
    .C(_4261_),
    .Y(_4264_)
);

AOI21X1 _11066_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4264_),
    .B(_4259_),
    .C(_4120_),
    .Y(_4265_)
);

INVX1 _11067_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4120_),
    .Y(_4266_)
);

NAND3X1 _11068_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4194_),
    .B(_4262_),
    .C(_4263_),
    .Y(_4267_)
);

OAI21X1 _11069_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4254_),
    .B(_4258_),
    .C(_4261_),
    .Y(_4268_)
);

AOI21X1 _11070_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4268_),
    .B(_4267_),
    .C(_4266_),
    .Y(_4269_)
);

OAI21X1 _11071_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4269_),
    .B(_4265_),
    .C(_4181_),
    .Y(_4270_)
);

NAND3X1 _11072_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4266_),
    .B(_4267_),
    .C(_4268_),
    .Y(_4271_)
);

NAND3X1 _11073_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4120_),
    .B(_4259_),
    .C(_4264_),
    .Y(_4272_)
);

NAND3X1 _11074_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4173_),
    .B(_4271_),
    .C(_4272_),
    .Y(_4273_)
);

AND2X2 _11075_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4270_),
    .B(_4273_),
    .Y(_4274_)
);

OAI21X1 _11076_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4192_),
    .B(_4189_),
    .C(_4274_),
    .Y(_4275_)
);

NOR2X1 _11077_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4192_),
    .B(_4189_),
    .Y(_4276_)
);

AOI21X1 _11078_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4272_),
    .B(_4271_),
    .C(_4173_),
    .Y(_4277_)
);

INVX1 _11079_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4273_),
    .Y(_4278_)
);

OAI21X1 _11080_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4277_),
    .B(_4278_),
    .C(_4276_),
    .Y(_4279_)
);

AND2X2 _11081_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4279_),
    .B(_4275_),
    .Y(_4781_[7])
);

NAND3X1 _11082_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4270_),
    .B(_4273_),
    .C(_4189_),
    .Y(_4280_)
);

AOI21X1 _11083_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4192_),
    .B(_4270_),
    .C(_4278_),
    .Y(_4281_)
);

NAND2X1 _11084_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4281_),
    .B(_4280_),
    .Y(_4282_)
);

INVX1 _11085_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4267_),
    .Y(_4283_)
);

AOI21X1 _11086_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4266_),
    .B(_4268_),
    .C(_4283_),
    .Y(_4284_)
);

OAI21X1 _11087_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4195_),
    .B(_4205_),
    .C(_4201_),
    .Y(_4285_)
);

INVX1 _11088_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4285_),
    .Y(_4286_)
);

AOI21X1 _11089_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4251_),
    .B(_4252_),
    .C(_4209_),
    .Y(_4287_)
);

OAI21X1 _11090_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4207_),
    .B(_4287_),
    .C(_4256_),
    .Y(_4288_)
);

NAND2X1 _11091_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [1]),
    .B(gnd),
    .Y(_4289_)
);

INVX2 _11092_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_4290_)
);

NOR2X1 _11093_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4755_),
    .B(_4290_),
    .Y(_4291_)
);

OAI21X1 _11094_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4210_),
    .B(_4215_),
    .C(_4214_),
    .Y(_4292_)
);

NOR2X1 _11095_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4291_),
    .B(_4292_),
    .Y(_4293_)
);

AND2X2 _11096_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4292_),
    .B(_4291_),
    .Y(_4294_)
);

OAI21X1 _11097_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4293_),
    .B(_4294_),
    .C(_4289_),
    .Y(_4295_)
);

INVX1 _11098_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4289_),
    .Y(_4296_)
);

OR2X2 _11099_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4292_),
    .B(_4291_),
    .Y(_4297_)
);

NAND2X1 _11100_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4291_),
    .B(_4292_),
    .Y(_4298_)
);

NAND3X1 _11101_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4296_),
    .B(_4298_),
    .C(_4297_),
    .Y(_4299_)
);

NAND2X1 _11102_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4295_),
    .B(_4299_),
    .Y(_4300_)
);

AOI21X1 _11103_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4241_),
    .B(_4238_),
    .C(_4224_),
    .Y(_4301_)
);

OAI21X1 _11104_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4223_),
    .B(_4301_),
    .C(_4245_),
    .Y(_4302_)
);

NAND2X1 _11105_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [3]),
    .B(vdd),
    .Y(_4303_)
);

INVX1 _11106_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_4304_)
);

OAI21X1 _11107_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4000_),
    .B(_4304_),
    .C(_4010_),
    .Y(_4305_)
);

NAND2X1 _11108_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [4]),
    .B(gnd),
    .Y(_4306_)
);

OAI21X1 _11109_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4303_),
    .B(_4306_),
    .C(_4305_),
    .Y(_4307_)
);

OAI21X1 _11110_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4225_),
    .B(_4233_),
    .C(_4232_),
    .Y(_4308_)
);

NAND2X1 _11111_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [7]),
    .Y(_4309_)
);

NAND2X1 _11112_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5]_5_bF$buf1 ),
    .Y(_4310_)
);

NAND3X1 _11113_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [6]),
    .C(_4310_),
    .Y(_4311_)
);

AND2X2 _11114_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5]_5_bF$buf0 ),
    .Y(_4312_)
);

OAI21X1 _11115_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4074_),
    .B(_4129_),
    .C(_4312_),
    .Y(_4313_)
);

AOI21X1 _11116_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4313_),
    .B(_4311_),
    .C(_4309_),
    .Y(_4314_)
);

INVX1 _11117_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4309_),
    .Y(_4315_)
);

AND2X2 _11118_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [6]),
    .Y(_4316_)
);

NAND2X1 _11119_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4312_),
    .B(_4316_),
    .Y(_4317_)
);

NAND2X1 _11120_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [6]),
    .Y(_4318_)
);

NAND2X1 _11121_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4310_),
    .B(_4318_),
    .Y(_4319_)
);

AOI21X1 _11122_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4317_),
    .B(_4319_),
    .C(_4315_),
    .Y(_4320_)
);

OAI21X1 _11123_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4320_),
    .B(_4314_),
    .C(_4308_),
    .Y(_4321_)
);

AOI21X1 _11124_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4231_),
    .B(_4234_),
    .C(_4240_),
    .Y(_4322_)
);

NAND3X1 _11125_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4315_),
    .B(_4319_),
    .C(_4317_),
    .Y(_4323_)
);

NAND3X1 _11126_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4309_),
    .B(_4311_),
    .C(_4313_),
    .Y(_4324_)
);

NAND3X1 _11127_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4323_),
    .B(_4324_),
    .C(_4322_),
    .Y(_4325_)
);

AOI21X1 _11128_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4321_),
    .B(_4325_),
    .C(_4307_),
    .Y(_4326_)
);

INVX1 _11129_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4307_),
    .Y(_4327_)
);

NAND3X1 _11130_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4308_),
    .B(_4323_),
    .C(_4324_),
    .Y(_4328_)
);

OAI21X1 _11131_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4320_),
    .B(_4314_),
    .C(_4322_),
    .Y(_4329_)
);

AOI21X1 _11132_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4329_),
    .B(_4328_),
    .C(_4327_),
    .Y(_4330_)
);

OAI21X1 _11133_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4326_),
    .B(_4330_),
    .C(_4302_),
    .Y(_4331_)
);

INVX1 _11134_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4245_),
    .Y(_4332_)
);

AOI21X1 _11135_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4244_),
    .B(_4246_),
    .C(_4332_),
    .Y(_4333_)
);

NAND3X1 _11136_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4327_),
    .B(_4328_),
    .C(_4329_),
    .Y(_4334_)
);

NAND3X1 _11137_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4307_),
    .B(_4325_),
    .C(_4321_),
    .Y(_4335_)
);

NAND3X1 _11138_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4334_),
    .B(_4335_),
    .C(_4333_),
    .Y(_4336_)
);

AOI21X1 _11139_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4336_),
    .B(_4331_),
    .C(_4300_),
    .Y(_4337_)
);

AND2X2 _11140_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4299_),
    .B(_4295_),
    .Y(_4338_)
);

NAND3X1 _11141_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4334_),
    .B(_4335_),
    .C(_4302_),
    .Y(_4339_)
);

OAI21X1 _11142_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4326_),
    .B(_4330_),
    .C(_4333_),
    .Y(_4340_)
);

AOI21X1 _11143_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4340_),
    .B(_4339_),
    .C(_4338_),
    .Y(_4341_)
);

OAI21X1 _11144_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4341_),
    .B(_4337_),
    .C(_4288_),
    .Y(_4342_)
);

INVX1 _11145_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4256_),
    .Y(_4343_)
);

AOI21X1 _11146_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4255_),
    .B(_4257_),
    .C(_4343_),
    .Y(_4344_)
);

NAND3X1 _11147_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4338_),
    .B(_4339_),
    .C(_4340_),
    .Y(_4345_)
);

NAND3X1 _11148_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4300_),
    .B(_4331_),
    .C(_4336_),
    .Y(_4346_)
);

NAND3X1 _11149_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4345_),
    .B(_4346_),
    .C(_4344_),
    .Y(_4347_)
);

AOI21X1 _11150_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4342_),
    .B(_4347_),
    .C(_4286_),
    .Y(_4348_)
);

NAND3X1 _11151_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4288_),
    .B(_4345_),
    .C(_4346_),
    .Y(_4349_)
);

OAI21X1 _11152_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4341_),
    .B(_4337_),
    .C(_4344_),
    .Y(_4350_)
);

AOI21X1 _11153_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4350_),
    .B(_4349_),
    .C(_4285_),
    .Y(_4351_)
);

OAI21X1 _11154_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4351_),
    .B(_4348_),
    .C(_4284_),
    .Y(_4352_)
);

AOI21X1 _11155_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4263_),
    .B(_4262_),
    .C(_4194_),
    .Y(_4353_)
);

OAI21X1 _11156_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4120_),
    .B(_4353_),
    .C(_4267_),
    .Y(_4354_)
);

NAND3X1 _11157_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4285_),
    .B(_4349_),
    .C(_4350_),
    .Y(_4355_)
);

NAND3X1 _11158_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4286_),
    .B(_4347_),
    .C(_4342_),
    .Y(_4356_)
);

NAND3X1 _11159_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4354_),
    .B(_4355_),
    .C(_4356_),
    .Y(_4357_)
);

NAND2X1 _11160_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4357_),
    .B(_4352_),
    .Y(_4358_)
);

NAND2X1 _11161_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4358_),
    .B(_4282_),
    .Y(_4359_)
);

OAI21X1 _11162_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4187_),
    .B(_4277_),
    .C(_4273_),
    .Y(_4360_)
);

AOI21X1 _11163_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4274_),
    .B(_4189_),
    .C(_4360_),
    .Y(_4361_)
);

AND2X2 _11164_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4352_),
    .B(_4357_),
    .Y(_4362_)
);

NAND2X1 _11165_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4362_),
    .B(_4361_),
    .Y(_4363_)
);

NAND2X1 _11166_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4359_),
    .B(_4363_),
    .Y(_4781_[8])
);

INVX1 _11167_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4357_),
    .Y(_4364_)
);

AOI21X1 _11168_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4282_),
    .B(_4352_),
    .C(_4364_),
    .Y(_4365_)
);

AOI21X1 _11169_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4346_),
    .B(_4345_),
    .C(_4288_),
    .Y(_4366_)
);

OAI21X1 _11170_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4286_),
    .B(_4366_),
    .C(_4349_),
    .Y(_4367_)
);

OAI21X1 _11171_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4289_),
    .B(_4293_),
    .C(_4298_),
    .Y(_4368_)
);

AOI21X1 _11172_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4334_),
    .B(_4335_),
    .C(_4302_),
    .Y(_4369_)
);

OAI21X1 _11173_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4300_),
    .B(_4369_),
    .C(_4339_),
    .Y(_4370_)
);

NAND2X1 _11174_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [2]),
    .B(gnd),
    .Y(_4371_)
);

NOR2X1 _11175_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4303_),
    .B(_4306_),
    .Y(_4372_)
);

NAND2X1 _11176_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_4372_),
    .Y(_4373_)
);

INVX1 _11177_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4373_),
    .Y(_4374_)
);

AOI21X1 _11178_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [3]),
    .B(gnd),
    .C(_4372_),
    .Y(_4375_)
);

OAI21X1 _11179_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4375_),
    .B(_4374_),
    .C(_4371_),
    .Y(_4376_)
);

INVX1 _11180_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4371_),
    .Y(_4377_)
);

INVX1 _11181_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4375_),
    .Y(_4378_)
);

NAND3X1 _11182_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4377_),
    .B(_4373_),
    .C(_4378_),
    .Y(_4379_)
);

AND2X2 _11183_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4379_),
    .B(_4376_),
    .Y(_4380_)
);

AOI21X1 _11184_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4324_),
    .B(_4323_),
    .C(_4308_),
    .Y(_4381_)
);

OAI21X1 _11185_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4307_),
    .B(_4381_),
    .C(_4328_),
    .Y(_4382_)
);

NOR2X1 _11186_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4117_),
    .B(_4306_),
    .Y(_4383_)
);

AND2X2 _11187_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4117_),
    .B(_4306_),
    .Y(_4384_)
);

NOR2X1 _11188_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4383_),
    .B(_4384_),
    .Y(_4385_)
);

NAND2X1 _11189_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [6]),
    .Y(_4386_)
);

AOI22X1 _11190_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5]_5_bF$buf3 ),
    .C(gnd),
    .D(\X[5] [6]),
    .Y(_4387_)
);

OAI22X1 _11191_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4239_),
    .B(_4386_),
    .C(_4309_),
    .D(_4387_),
    .Y(_4388_)
);

AOI22X1 _11192_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [6]),
    .C(gnd),
    .D(\X[5] [7]),
    .Y(_4389_)
);

AND2X2 _11193_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [7]),
    .Y(_4390_)
);

AOI21X1 _11194_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4316_),
    .B(_4390_),
    .C(_4389_),
    .Y(_4391_)
);

NAND2X1 _11195_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4391_),
    .B(_4388_),
    .Y(_4392_)
);

AND2X2 _11196_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [6]),
    .Y(_4393_)
);

AOI22X1 _11197_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4227_),
    .B(_4393_),
    .C(_4319_),
    .D(_4315_),
    .Y(_4394_)
);

NAND2X1 _11198_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [7]),
    .Y(_4395_)
);

NAND2X1 _11199_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4386_),
    .B(_4395_),
    .Y(_4396_)
);

NAND2X1 _11200_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [7]),
    .Y(_4397_)
);

OAI21X1 _11201_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4318_),
    .B(_4397_),
    .C(_4396_),
    .Y(_4398_)
);

NAND2X1 _11202_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4398_),
    .B(_4394_),
    .Y(_4399_)
);

NAND3X1 _11203_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4385_),
    .B(_4392_),
    .C(_4399_),
    .Y(_4400_)
);

NAND2X1 _11204_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5]_5_bF$buf2 ),
    .B(gnd),
    .Y(_4401_)
);

INVX1 _11205_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [4]),
    .Y(_4402_)
);

OAI21X1 _11206_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4402_),
    .B(_4304_),
    .C(_4117_),
    .Y(_4403_)
);

OAI21X1 _11207_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4010_),
    .B(_4401_),
    .C(_4403_),
    .Y(_4404_)
);

NAND2X1 _11208_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4388_),
    .B(_4398_),
    .Y(_4405_)
);

NAND2X1 _11209_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4391_),
    .B(_4394_),
    .Y(_4406_)
);

NAND3X1 _11210_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4404_),
    .B(_4405_),
    .C(_4406_),
    .Y(_4407_)
);

NAND3X1 _11211_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4400_),
    .B(_4407_),
    .C(_4382_),
    .Y(_4408_)
);

NAND2X1 _11212_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4400_),
    .B(_4407_),
    .Y(_4409_)
);

NAND3X1 _11213_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4328_),
    .B(_4334_),
    .C(_4409_),
    .Y(_4410_)
);

NAND3X1 _11214_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4380_),
    .B(_4408_),
    .C(_4410_),
    .Y(_4411_)
);

NAND2X1 _11215_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4376_),
    .B(_4379_),
    .Y(_4412_)
);

AOI21X1 _11216_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4328_),
    .B(_4334_),
    .C(_4409_),
    .Y(_4413_)
);

AOI21X1 _11217_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4400_),
    .B(_4407_),
    .C(_4382_),
    .Y(_4414_)
);

OAI21X1 _11218_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4414_),
    .B(_4413_),
    .C(_4412_),
    .Y(_4415_)
);

NAND3X1 _11219_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4411_),
    .B(_4415_),
    .C(_4370_),
    .Y(_4416_)
);

INVX1 _11220_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4339_),
    .Y(_4417_)
);

AOI21X1 _11221_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4338_),
    .B(_4340_),
    .C(_4417_),
    .Y(_4418_)
);

INVX1 _11222_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4411_),
    .Y(_4419_)
);

AOI21X1 _11223_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4410_),
    .B(_4408_),
    .C(_4380_),
    .Y(_4420_)
);

OAI21X1 _11224_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4420_),
    .B(_4419_),
    .C(_4418_),
    .Y(_4421_)
);

NAND3X1 _11225_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4368_),
    .B(_4416_),
    .C(_4421_),
    .Y(_4422_)
);

INVX1 _11226_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4368_),
    .Y(_4423_)
);

INVX1 _11227_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4416_),
    .Y(_4424_)
);

AOI21X1 _11228_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4415_),
    .B(_4411_),
    .C(_4370_),
    .Y(_4425_)
);

OAI21X1 _11229_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4425_),
    .B(_4424_),
    .C(_4423_),
    .Y(_4426_)
);

NAND3X1 _11230_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4367_),
    .B(_4422_),
    .C(_4426_),
    .Y(_4427_)
);

INVX1 _11231_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4349_),
    .Y(_4428_)
);

AOI21X1 _11232_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4285_),
    .B(_4350_),
    .C(_4428_),
    .Y(_4429_)
);

OAI21X1 _11233_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4420_),
    .B(_4419_),
    .C(_4370_),
    .Y(_4430_)
);

NAND3X1 _11234_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4411_),
    .B(_4415_),
    .C(_4418_),
    .Y(_4431_)
);

AOI21X1 _11235_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4431_),
    .B(_4430_),
    .C(_4423_),
    .Y(_4432_)
);

AOI21X1 _11236_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4421_),
    .B(_4416_),
    .C(_4368_),
    .Y(_4433_)
);

OAI21X1 _11237_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4432_),
    .B(_4433_),
    .C(_4429_),
    .Y(_4434_)
);

AND2X2 _11238_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4434_),
    .B(_4427_),
    .Y(_4435_)
);

OR2X2 _11239_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4365_),
    .B(_4435_),
    .Y(_4436_)
);

NAND2X1 _11240_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4435_),
    .B(_4365_),
    .Y(_4437_)
);

NAND2X1 _11241_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4437_),
    .B(_4436_),
    .Y(_4781_[9])
);

NAND2X1 _11242_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4427_),
    .B(_4434_),
    .Y(_4438_)
);

NOR2X1 _11243_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4358_),
    .B(_4438_),
    .Y(_4439_)
);

NAND2X1 _11244_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4439_),
    .B(_4282_),
    .Y(_4440_)
);

AOI21X1 _11245_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4426_),
    .B(_4422_),
    .C(_4367_),
    .Y(_4441_)
);

AOI21X1 _11246_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4357_),
    .B(_4427_),
    .C(_4441_),
    .Y(_4442_)
);

INVX1 _11247_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4442_),
    .Y(_4443_)
);

OAI21X1 _11248_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4423_),
    .B(_4425_),
    .C(_4416_),
    .Y(_4444_)
);

OAI21X1 _11249_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4371_),
    .B(_4375_),
    .C(_4373_),
    .Y(_4445_)
);

OAI21X1 _11250_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4412_),
    .B(_4414_),
    .C(_4408_),
    .Y(_4446_)
);

INVX2 _11251_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_4447_)
);

NOR3X1 _11252_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4290_),
    .B(_4117_),
    .C(_4306_),
    .Y(_4448_)
);

OAI22X1 _11253_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4402_),
    .B(_4290_),
    .C(_4010_),
    .D(_4401_),
    .Y(_4449_)
);

INVX1 _11254_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4449_),
    .Y(_4450_)
);

OAI22X1 _11255_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4000_),
    .B(_4447_),
    .C(_4448_),
    .D(_4450_),
    .Y(_4451_)
);

NOR2X1 _11256_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4000_),
    .B(_4447_),
    .Y(_4452_)
);

NAND2X1 _11257_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_4383_),
    .Y(_4453_)
);

NAND3X1 _11258_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4452_),
    .B(_4449_),
    .C(_4453_),
    .Y(_4454_)
);

AND2X2 _11259_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4451_),
    .B(_4454_),
    .Y(_4455_)
);

NOR2X1 _11260_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4391_),
    .B(_4388_),
    .Y(_4456_)
);

OAI21X1 _11261_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4404_),
    .B(_4456_),
    .C(_4392_),
    .Y(_4457_)
);

NAND2X1 _11262_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [6]),
    .Y(_4458_)
);

NOR2X1 _11263_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4458_),
    .B(_4401_),
    .Y(_4459_)
);

AND2X2 _11264_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4458_),
    .B(_4401_),
    .Y(_4460_)
);

OAI22X1 _11265_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4316_),
    .B(_4397_),
    .C(_4459_),
    .D(_4460_),
    .Y(_4461_)
);

AND2X2 _11266_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[5] [6]),
    .Y(_4462_)
);

AND2X2 _11267_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5]_5_bF$buf1 ),
    .B(gnd),
    .Y(_4463_)
);

NAND2X1 _11268_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4462_),
    .B(_4463_),
    .Y(_4464_)
);

OAI21X1 _11269_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4059_),
    .B(_4304_),
    .C(_4458_),
    .Y(_4465_)
);

AOI21X1 _11270_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [6]),
    .C(_4397_),
    .Y(_4466_)
);

NAND3X1 _11271_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4465_),
    .B(_4466_),
    .C(_4464_),
    .Y(_4467_)
);

AND2X2 _11272_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4461_),
    .B(_4467_),
    .Y(_4468_)
);

NAND2X1 _11273_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4468_),
    .B(_4457_),
    .Y(_4469_)
);

NAND2X1 _11274_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4467_),
    .B(_4461_),
    .Y(_4470_)
);

NAND3X1 _11275_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4392_),
    .B(_4470_),
    .C(_4400_),
    .Y(_4471_)
);

NAND3X1 _11276_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4455_),
    .B(_4471_),
    .C(_4469_),
    .Y(_4472_)
);

NAND2X1 _11277_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4454_),
    .B(_4451_),
    .Y(_4473_)
);

NAND2X1 _11278_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4470_),
    .B(_4457_),
    .Y(_4474_)
);

NAND3X1 _11279_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4392_),
    .B(_4468_),
    .C(_4400_),
    .Y(_4475_)
);

NAND3X1 _11280_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4473_),
    .B(_4475_),
    .C(_4474_),
    .Y(_4476_)
);

NAND3X1 _11281_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4472_),
    .B(_4476_),
    .C(_4446_),
    .Y(_4477_)
);

NAND2X1 _11282_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4476_),
    .B(_4472_),
    .Y(_4478_)
);

NAND3X1 _11283_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4408_),
    .B(_4411_),
    .C(_4478_),
    .Y(_4479_)
);

NAND3X1 _11284_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4445_),
    .B(_4479_),
    .C(_4477_),
    .Y(_4480_)
);

INVX1 _11285_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4445_),
    .Y(_4481_)
);

NAND2X1 _11286_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4478_),
    .B(_4446_),
    .Y(_4482_)
);

AOI21X1 _11287_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4380_),
    .B(_4410_),
    .C(_4413_),
    .Y(_4483_)
);

AND2X2 _11288_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4472_),
    .B(_4476_),
    .Y(_4484_)
);

NAND2X1 _11289_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4483_),
    .B(_4484_),
    .Y(_4485_)
);

NAND3X1 _11290_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4481_),
    .B(_4482_),
    .C(_4485_),
    .Y(_4486_)
);

AOI21X1 _11291_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4480_),
    .B(_4486_),
    .C(_4444_),
    .Y(_4487_)
);

NAND2X1 _11292_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4480_),
    .B(_4486_),
    .Y(_4488_)
);

AOI21X1 _11293_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4416_),
    .B(_4422_),
    .C(_4488_),
    .Y(_4489_)
);

NOR2X1 _11294_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4487_),
    .B(_4489_),
    .Y(_4490_)
);

INVX1 _11295_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4490_),
    .Y(_4491_)
);

AOI21X1 _11296_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4440_),
    .B(_4443_),
    .C(_4491_),
    .Y(_4492_)
);

NAND2X1 _11297_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4362_),
    .B(_4435_),
    .Y(_4493_)
);

OAI21X1 _11298_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4493_),
    .B(_4361_),
    .C(_4443_),
    .Y(_4494_)
);

NOR2X1 _11299_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4490_),
    .B(_4494_),
    .Y(_4495_)
);

NOR2X1 _11300_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4492_),
    .B(_4495_),
    .Y(_4781_[10])
);

NAND3X1 _11301_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4480_),
    .B(_4486_),
    .C(_4444_),
    .Y(_4496_)
);

NAND2X1 _11302_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4490_),
    .B(_4494_),
    .Y(_4497_)
);

NOR2X1 _11303_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4478_),
    .B(_4483_),
    .Y(_4498_)
);

AOI21X1 _11304_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4445_),
    .B(_4479_),
    .C(_4498_),
    .Y(_4499_)
);

NAND2X1 _11305_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4453_),
    .B(_4454_),
    .Y(_4500_)
);

NAND2X1 _11306_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4469_),
    .B(_4472_),
    .Y(_4501_)
);

NOR3X1 _11307_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4290_),
    .B(_4458_),
    .C(_4401_),
    .Y(_4502_)
);

AOI22X1 _11308_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5]_5_bF$buf0 ),
    .B(gnd),
    .C(_4462_),
    .D(_4463_),
    .Y(_4503_)
);

OAI22X1 _11309_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4402_),
    .B(_4447_),
    .C(_4503_),
    .D(_4502_),
    .Y(_4504_)
);

NOR2X1 _11310_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4402_),
    .B(_4447_),
    .Y(_4505_)
);

NAND2X1 _11311_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_4459_),
    .Y(_4506_)
);

OAI21X1 _11312_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4059_),
    .B(_4290_),
    .C(_4464_),
    .Y(_4507_)
);

NAND3X1 _11313_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4505_),
    .B(_4506_),
    .C(_4507_),
    .Y(_4508_)
);

NAND2X1 _11314_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4504_),
    .B(_4508_),
    .Y(_4509_)
);

NAND2X1 _11315_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4316_),
    .B(_4390_),
    .Y(_4510_)
);

NAND2X1 _11316_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[5] [7]),
    .Y(_4511_)
);

OAI22X1 _11317_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4218_),
    .B(_4220_),
    .C(_4304_),
    .D(_4129_),
    .Y(_4512_)
);

OAI21X1 _11318_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4458_),
    .B(_4511_),
    .C(_4512_),
    .Y(_4513_)
);

NAND3X1 _11319_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4510_),
    .B(_4513_),
    .C(_4467_),
    .Y(_4514_)
);

INVX1 _11320_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4514_),
    .Y(_4515_)
);

AOI21X1 _11321_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4467_),
    .B(_4510_),
    .C(_4513_),
    .Y(_4516_)
);

OAI21X1 _11322_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4516_),
    .B(_4515_),
    .C(_4509_),
    .Y(_4517_)
);

AND2X2 _11323_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4508_),
    .B(_4504_),
    .Y(_4518_)
);

INVX1 _11324_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4516_),
    .Y(_4519_)
);

NAND3X1 _11325_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4514_),
    .B(_4519_),
    .C(_4518_),
    .Y(_4520_)
);

AND2X2 _11326_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4520_),
    .B(_4517_),
    .Y(_4521_)
);

NAND2X1 _11327_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4521_),
    .B(_4501_),
    .Y(_4522_)
);

AOI21X1 _11328_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4400_),
    .B(_4392_),
    .C(_4470_),
    .Y(_4523_)
);

AOI21X1 _11329_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4455_),
    .B(_4471_),
    .C(_4523_),
    .Y(_4524_)
);

NAND2X1 _11330_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4517_),
    .B(_4520_),
    .Y(_4525_)
);

NAND2X1 _11331_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4525_),
    .B(_4524_),
    .Y(_4526_)
);

NAND3X1 _11332_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4500_),
    .B(_4526_),
    .C(_4522_),
    .Y(_4527_)
);

INVX1 _11333_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4500_),
    .Y(_4528_)
);

NAND2X1 _11334_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4525_),
    .B(_4501_),
    .Y(_4529_)
);

NAND2X1 _11335_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4524_),
    .B(_4521_),
    .Y(_4530_)
);

NAND3X1 _11336_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4528_),
    .B(_4530_),
    .C(_4529_),
    .Y(_4531_)
);

NAND2X1 _11337_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4527_),
    .B(_4531_),
    .Y(_4532_)
);

NAND2X1 _11338_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4532_),
    .B(_4499_),
    .Y(_4533_)
);

AOI21X1 _11339_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4472_),
    .B(_4476_),
    .C(_4446_),
    .Y(_4534_)
);

OAI21X1 _11340_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4481_),
    .B(_4534_),
    .C(_4477_),
    .Y(_4535_)
);

NAND3X1 _11341_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4527_),
    .B(_4531_),
    .C(_4535_),
    .Y(_4536_)
);

NAND2X1 _11342_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4533_),
    .B(_4536_),
    .Y(_4537_)
);

INVX1 _11343_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4537_),
    .Y(_4538_)
);

NAND3X1 _11344_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4496_),
    .B(_4538_),
    .C(_4497_),
    .Y(_4539_)
);

OAI21X1 _11345_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4489_),
    .B(_4492_),
    .C(_4537_),
    .Y(_4540_)
);

NAND2X1 _11346_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4539_),
    .B(_4540_),
    .Y(_4781_[11])
);

NOR3X1 _11347_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4487_),
    .B(_4489_),
    .C(_4537_),
    .Y(_4541_)
);

NAND3X1 _11348_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4439_),
    .B(_4541_),
    .C(_4282_),
    .Y(_4542_)
);

OAI21X1 _11349_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4496_),
    .B(_4537_),
    .C(_4536_),
    .Y(_4543_)
);

AOI21X1 _11350_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4541_),
    .B(_4442_),
    .C(_4543_),
    .Y(_4544_)
);

AND2X2 _11351_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4527_),
    .B(_4522_),
    .Y(_4545_)
);

OAI21X1 _11352_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4290_),
    .B(_4464_),
    .C(_4508_),
    .Y(_4546_)
);

OAI21X1 _11353_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4515_),
    .B(_4509_),
    .C(_4519_),
    .Y(_4547_)
);

INVX1 _11354_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4547_),
    .Y(_4548_)
);

INVX1 _11355_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4511_),
    .Y(_4549_)
);

NOR2X1 _11356_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4059_),
    .B(_4447_),
    .Y(_4550_)
);

NOR2X1 _11357_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4458_),
    .B(_4511_),
    .Y(_4551_)
);

NOR2X1 _11358_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4129_),
    .B(_4290_),
    .Y(_4552_)
);

NOR2X1 _11359_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4552_),
    .B(_4551_),
    .Y(_4553_)
);

AOI21X1 _11360_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_4551_),
    .C(_4553_),
    .Y(_4554_)
);

OR2X2 _11361_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4554_),
    .B(_4550_),
    .Y(_4555_)
);

NAND2X1 _11362_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4550_),
    .B(_4554_),
    .Y(_4556_)
);

NAND3X1 _11363_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4549_),
    .B(_4556_),
    .C(_4555_),
    .Y(_4557_)
);

NOR2X1 _11364_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4550_),
    .B(_4554_),
    .Y(_4558_)
);

INVX1 _11365_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4556_),
    .Y(_4559_)
);

OAI21X1 _11366_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4558_),
    .B(_4559_),
    .C(_4511_),
    .Y(_4560_)
);

NAND2X1 _11367_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4557_),
    .B(_4560_),
    .Y(_4561_)
);

NAND2X1 _11368_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4548_),
    .B(_4561_),
    .Y(_4562_)
);

NAND3X1 _11369_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4547_),
    .B(_4557_),
    .C(_4560_),
    .Y(_4563_)
);

AOI21X1 _11370_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4562_),
    .B(_4563_),
    .C(_4546_),
    .Y(_4564_)
);

NAND3X1 _11371_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4546_),
    .B(_4563_),
    .C(_4562_),
    .Y(_4565_)
);

INVX1 _11372_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4565_),
    .Y(_4566_)
);

OAI21X1 _11373_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4564_),
    .B(_4566_),
    .C(_4545_),
    .Y(_4567_)
);

OR2X2 _11374_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4566_),
    .B(_4564_),
    .Y(_4568_)
);

OR2X2 _11375_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4568_),
    .B(_4545_),
    .Y(_4569_)
);

NAND2X1 _11376_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4567_),
    .B(_4569_),
    .Y(_4570_)
);

AOI21X1 _11377_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4542_),
    .B(_4544_),
    .C(_4570_),
    .Y(_4571_)
);

NAND3X1 _11378_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4362_),
    .B(_4435_),
    .C(_4541_),
    .Y(_4572_)
);

OAI21X1 _11379_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4361_),
    .B(_4572_),
    .C(_4544_),
    .Y(_4573_)
);

INVX1 _11380_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4570_),
    .Y(_4574_)
);

NOR2X1 _11381_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4574_),
    .B(_4573_),
    .Y(_4575_)
);

NOR2X1 _11382_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4571_),
    .B(_4575_),
    .Y(_4781_[12])
);

NOR2X1 _11383_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4545_),
    .B(_4568_),
    .Y(_4576_)
);

INVX1 _11384_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4551_),
    .Y(_4577_)
);

OAI21X1 _11385_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4290_),
    .B(_4577_),
    .C(_4556_),
    .Y(_4578_)
);

INVX1 _11386_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4578_),
    .Y(_4579_)
);

NOR2X1 _11387_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4220_),
    .B(_4447_),
    .Y(_4580_)
);

NAND2X1 _11388_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4552_),
    .B(_4580_),
    .Y(_4581_)
);

OAI22X1 _11389_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4129_),
    .B(_4447_),
    .C(_4290_),
    .D(_4220_),
    .Y(_4582_)
);

NAND2X1 _11390_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4582_),
    .B(_4581_),
    .Y(_4583_)
);

NAND2X1 _11391_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4583_),
    .B(_4557_),
    .Y(_4584_)
);

OR2X2 _11392_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4557_),
    .B(_4583_),
    .Y(_4585_)
);

NAND2X1 _11393_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4584_),
    .B(_4585_),
    .Y(_4586_)
);

NAND2X1 _11394_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4579_),
    .B(_4586_),
    .Y(_4587_)
);

OR2X2 _11395_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4586_),
    .B(_4579_),
    .Y(_4588_)
);

NAND2X1 _11396_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4587_),
    .B(_4588_),
    .Y(_4589_)
);

NAND3X1 _11397_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4563_),
    .B(_4565_),
    .C(_4589_),
    .Y(_4590_)
);

OAI21X1 _11398_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4548_),
    .B(_4561_),
    .C(_4565_),
    .Y(_4591_)
);

AND2X2 _11399_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4588_),
    .B(_4587_),
    .Y(_4592_)
);

NAND2X1 _11400_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4591_),
    .B(_4592_),
    .Y(_4593_)
);

NAND2X1 _11401_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4590_),
    .B(_4593_),
    .Y(_4594_)
);

OAI21X1 _11402_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4576_),
    .B(_4571_),
    .C(_4594_),
    .Y(_4595_)
);

NAND2X1 _11403_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4574_),
    .B(_4573_),
    .Y(_4596_)
);

AND2X2 _11404_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4593_),
    .B(_4590_),
    .Y(_4597_)
);

NAND3X1 _11405_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4569_),
    .B(_4597_),
    .C(_4596_),
    .Y(_4598_)
);

NAND2X1 _11406_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4598_),
    .B(_4595_),
    .Y(_4781_[13])
);

NAND3X1 _11407_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4567_),
    .B(_4569_),
    .C(_4597_),
    .Y(_4599_)
);

AOI21X1 _11408_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4542_),
    .B(_4544_),
    .C(_4599_),
    .Y(_4600_)
);

OAI21X1 _11409_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4569_),
    .B(_4594_),
    .C(_4593_),
    .Y(_4601_)
);

OAI21X1 _11410_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4579_),
    .B(_4586_),
    .C(_4585_),
    .Y(_4602_)
);

AND2X2 _11411_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4581_),
    .B(_4580_),
    .Y(_4603_)
);

OR2X2 _11412_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4602_),
    .B(_4603_),
    .Y(_4604_)
);

NAND2X1 _11413_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4603_),
    .B(_4602_),
    .Y(_4605_)
);

NAND2X1 _11414_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4605_),
    .B(_4604_),
    .Y(_4606_)
);

OAI21X1 _11415_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4601_),
    .B(_4600_),
    .C(_4606_),
    .Y(_4607_)
);

INVX1 _11416_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4567_),
    .Y(_4608_)
);

NOR3X1 _11417_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4608_),
    .B(_4576_),
    .C(_4594_),
    .Y(_4609_)
);

NAND2X1 _11418_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4609_),
    .B(_4573_),
    .Y(_4610_)
);

INVX1 _11419_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4601_),
    .Y(_4611_)
);

INVX1 _11420_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4606_),
    .Y(_4612_)
);

NAND3X1 _11421_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4611_),
    .B(_4612_),
    .C(_4610_),
    .Y(_4613_)
);

NAND2X1 _11422_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4613_),
    .B(_4607_),
    .Y(_4781_[14])
);

OAI21X1 _11423_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4601_),
    .B(_4600_),
    .C(_4612_),
    .Y(_4614_)
);

OAI21X1 _11424_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4552_),
    .B(_4602_),
    .C(_4580_),
    .Y(_4615_)
);

NAND2X1 _11425_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4615_),
    .B(_4614_),
    .Y(_4781_[15])
);

INVX1 _11426_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4009_),
    .Y(_4776_[0])
);

AND2X2 _11427_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [0]),
    .B(\u_fir_pe5.mul [0]),
    .Y(_4616_)
);

INVX1 _11428_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [1]),
    .Y(_4617_)
);

INVX1 _11429_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.mul [1]),
    .Y(_4618_)
);

NOR2X1 _11430_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4617_),
    .B(_4618_),
    .Y(_4619_)
);

NOR2X1 _11431_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [1]),
    .B(\u_fir_pe5.mul [1]),
    .Y(_4620_)
);

NOR2X1 _11432_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4620_),
    .B(_4619_),
    .Y(_4621_)
);

NAND2X1 _11433_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4616_),
    .B(_4621_),
    .Y(_4622_)
);

INVX1 _11434_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4622_),
    .Y(_4623_)
);

NOR2X1 _11435_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4616_),
    .B(_4621_),
    .Y(_4624_)
);

NOR2X1 _11436_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4624_),
    .B(_4623_),
    .Y(_4775_[1])
);

OAI21X1 _11437_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4617_),
    .B(_4618_),
    .C(_4622_),
    .Y(_4625_)
);

AND2X2 _11438_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [2]),
    .B(\u_fir_pe5.mul [2]),
    .Y(_4626_)
);

NOR2X1 _11439_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [2]),
    .B(\u_fir_pe5.mul [2]),
    .Y(_4627_)
);

OAI21X1 _11440_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4626_),
    .B(_4627_),
    .C(_4625_),
    .Y(_4628_)
);

INVX1 _11441_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4625_),
    .Y(_4629_)
);

NOR2X1 _11442_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4627_),
    .B(_4626_),
    .Y(_4630_)
);

NAND2X1 _11443_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4630_),
    .B(_4629_),
    .Y(_4631_)
);

NAND2X1 _11444_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4628_),
    .B(_4631_),
    .Y(_4775_[2])
);

AOI21X1 _11445_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4625_),
    .B(_4630_),
    .C(_4626_),
    .Y(_4632_)
);

INVX1 _11446_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [3]),
    .Y(_4633_)
);

INVX1 _11447_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.mul [3]),
    .Y(_4634_)
);

NOR2X1 _11448_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4633_),
    .B(_4634_),
    .Y(_4635_)
);

NOR2X1 _11449_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [3]),
    .B(\u_fir_pe5.mul [3]),
    .Y(_4636_)
);

NOR2X1 _11450_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4636_),
    .B(_4635_),
    .Y(_4637_)
);

NAND2X1 _11451_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4637_),
    .B(_4632_),
    .Y(_4638_)
);

OR2X2 _11452_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4632_),
    .B(_4637_),
    .Y(_4639_)
);

NAND2X1 _11453_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4638_),
    .B(_4639_),
    .Y(_4775_[3])
);

INVX1 _11454_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [4]),
    .Y(_4640_)
);

INVX1 _11455_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.mul [4]),
    .Y(_4641_)
);

NOR2X1 _11456_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4640_),
    .B(_4641_),
    .Y(_4642_)
);

NOR2X1 _11457_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [4]),
    .B(\u_fir_pe5.mul [4]),
    .Y(_4643_)
);

NOR2X1 _11458_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4643_),
    .B(_4642_),
    .Y(_4644_)
);

INVX1 _11459_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4635_),
    .Y(_4645_)
);

OAI21X1 _11460_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4636_),
    .B(_4632_),
    .C(_4645_),
    .Y(_4646_)
);

NAND2X1 _11461_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4644_),
    .B(_4646_),
    .Y(_4647_)
);

OR2X2 _11462_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4646_),
    .B(_4644_),
    .Y(_4648_)
);

AND2X2 _11463_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4648_),
    .B(_4647_),
    .Y(_4775_[4])
);

OAI21X1 _11464_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4640_),
    .B(_4641_),
    .C(_4647_),
    .Y(_4649_)
);

INVX1 _11465_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [5]),
    .Y(_4650_)
);

INVX1 _11466_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.mul [5]),
    .Y(_4651_)
);

NOR2X1 _11467_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4650_),
    .B(_4651_),
    .Y(_4652_)
);

NOR2X1 _11468_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [5]),
    .B(\u_fir_pe5.mul [5]),
    .Y(_4653_)
);

NOR2X1 _11469_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4653_),
    .B(_4652_),
    .Y(_4654_)
);

NAND2X1 _11470_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4654_),
    .B(_4649_),
    .Y(_4655_)
);

OR2X2 _11471_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4649_),
    .B(_4654_),
    .Y(_4656_)
);

AND2X2 _11472_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4656_),
    .B(_4655_),
    .Y(_4775_[5])
);

OAI21X1 _11473_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4650_),
    .B(_4651_),
    .C(_4655_),
    .Y(_4657_)
);

INVX1 _11474_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [6]),
    .Y(_4658_)
);

INVX1 _11475_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.mul [6]),
    .Y(_4659_)
);

NOR2X1 _11476_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4658_),
    .B(_4659_),
    .Y(_4660_)
);

NOR2X1 _11477_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [6]),
    .B(\u_fir_pe5.mul [6]),
    .Y(_4661_)
);

NOR2X1 _11478_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4661_),
    .B(_4660_),
    .Y(_4662_)
);

NAND2X1 _11479_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4662_),
    .B(_4657_),
    .Y(_4663_)
);

OR2X2 _11480_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4657_),
    .B(_4662_),
    .Y(_4664_)
);

AND2X2 _11481_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4664_),
    .B(_4663_),
    .Y(_4775_[6])
);

OAI21X1 _11482_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4658_),
    .B(_4659_),
    .C(_4663_),
    .Y(_4665_)
);

INVX1 _11483_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [7]),
    .Y(_4666_)
);

INVX1 _11484_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.mul [7]),
    .Y(_4667_)
);

NOR2X1 _11485_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4666_),
    .B(_4667_),
    .Y(_4668_)
);

NOR2X1 _11486_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [7]),
    .B(\u_fir_pe5.mul [7]),
    .Y(_4669_)
);

OAI21X1 _11487_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4668_),
    .B(_4669_),
    .C(_4665_),
    .Y(_4670_)
);

INVX1 _11488_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4665_),
    .Y(_4671_)
);

NOR2X1 _11489_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4669_),
    .B(_4668_),
    .Y(_4672_)
);

NAND2X1 _11490_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4672_),
    .B(_4671_),
    .Y(_4673_)
);

NAND2X1 _11491_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4670_),
    .B(_4673_),
    .Y(_4775_[7])
);

INVX1 _11492_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [8]),
    .Y(_4675_)
);

INVX1 _11493_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.mul [8]),
    .Y(_4676_)
);

NOR2X1 _11494_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4675_),
    .B(_4676_),
    .Y(_4677_)
);

NOR2X1 _11495_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [8]),
    .B(\u_fir_pe5.mul [8]),
    .Y(_4678_)
);

NAND2X1 _11496_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4642_),
    .B(_4654_),
    .Y(_4679_)
);

OAI21X1 _11497_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4650_),
    .B(_4651_),
    .C(_4679_),
    .Y(_4680_)
);

NAND2X1 _11498_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4660_),
    .B(_4672_),
    .Y(_4681_)
);

OAI21X1 _11499_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4666_),
    .B(_4667_),
    .C(_4681_),
    .Y(_4682_)
);

AND2X2 _11500_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4662_),
    .B(_4672_),
    .Y(_4683_)
);

AOI21X1 _11501_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4680_),
    .B(_4683_),
    .C(_4682_),
    .Y(_4684_)
);

AND2X2 _11502_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4644_),
    .B(_4654_),
    .Y(_4686_)
);

NAND3X1 _11503_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4686_),
    .B(_4683_),
    .C(_4646_),
    .Y(_4687_)
);

NAND2X1 _11504_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4684_),
    .B(_4687_),
    .Y(_4688_)
);

OAI21X1 _11505_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4677_),
    .B(_4678_),
    .C(_4688_),
    .Y(_4689_)
);

NOR2X1 _11506_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4678_),
    .B(_4677_),
    .Y(_4690_)
);

INVX1 _11507_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4688_),
    .Y(_4691_)
);

NAND2X1 _11508_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4690_),
    .B(_4691_),
    .Y(_4692_)
);

NAND2X1 _11509_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4689_),
    .B(_4692_),
    .Y(_4775_[8])
);

INVX1 _11510_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4677_),
    .Y(_4693_)
);

INVX1 _11511_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4690_),
    .Y(_4694_)
);

OAI21X1 _11512_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4694_),
    .B(_4691_),
    .C(_4693_),
    .Y(_4696_)
);

AND2X2 _11513_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [9]),
    .B(\u_fir_pe5.mul [9]),
    .Y(_4697_)
);

NOR2X1 _11514_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [9]),
    .B(\u_fir_pe5.mul [9]),
    .Y(_4698_)
);

NOR2X1 _11515_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4698_),
    .B(_4697_),
    .Y(_4699_)
);

INVX1 _11516_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4699_),
    .Y(_4700_)
);

OR2X2 _11517_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4696_),
    .B(_4700_),
    .Y(_4701_)
);

OAI21X1 _11518_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4697_),
    .B(_4698_),
    .C(_4696_),
    .Y(_4702_)
);

NAND2X1 _11519_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4702_),
    .B(_4701_),
    .Y(_4775_[9])
);

NOR2X1 _11520_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4700_),
    .B(_4694_),
    .Y(_4703_)
);

AOI21X1 _11521_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4699_),
    .B(_4677_),
    .C(_4697_),
    .Y(_4704_)
);

INVX1 _11522_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4704_),
    .Y(_4706_)
);

AOI21X1 _11523_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4688_),
    .B(_4703_),
    .C(_4706_),
    .Y(_4707_)
);

INVX1 _11524_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4707_),
    .Y(_4708_)
);

INVX1 _11525_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [10]),
    .Y(_4709_)
);

INVX1 _11526_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.mul [10]),
    .Y(_4710_)
);

NOR2X1 _11527_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4709_),
    .B(_4710_),
    .Y(_4711_)
);

NOR2X1 _11528_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [10]),
    .B(\u_fir_pe5.mul [10]),
    .Y(_4712_)
);

NOR2X1 _11529_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4712_),
    .B(_4711_),
    .Y(_4713_)
);

NAND2X1 _11530_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4713_),
    .B(_4708_),
    .Y(_4714_)
);

OAI21X1 _11531_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4711_),
    .B(_4712_),
    .C(_4707_),
    .Y(_4715_)
);

AND2X2 _11532_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4714_),
    .B(_4715_),
    .Y(_4775_[10])
);

OAI21X1 _11533_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4709_),
    .B(_4710_),
    .C(_4714_),
    .Y(_4717_)
);

AND2X2 _11534_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [11]),
    .B(\u_fir_pe5.mul [11]),
    .Y(_4718_)
);

NOR2X1 _11535_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [11]),
    .B(\u_fir_pe5.mul [11]),
    .Y(_4719_)
);

NOR2X1 _11536_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4719_),
    .B(_4718_),
    .Y(_4720_)
);

NOR2X1 _11537_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4720_),
    .B(_4717_),
    .Y(_4721_)
);

AND2X2 _11538_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4717_),
    .B(_4720_),
    .Y(_4722_)
);

NOR2X1 _11539_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4721_),
    .B(_4722_),
    .Y(_4775_[11])
);

AOI21X1 _11540_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4720_),
    .B(_4711_),
    .C(_4718_),
    .Y(_4723_)
);

NAND2X1 _11541_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4720_),
    .B(_4713_),
    .Y(_4724_)
);

OAI21X1 _11542_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4724_),
    .B(_4707_),
    .C(_4723_),
    .Y(_4726_)
);

INVX1 _11543_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [12]),
    .Y(_4727_)
);

INVX1 _11544_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.mul [12]),
    .Y(_4728_)
);

NOR2X1 _11545_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4727_),
    .B(_4728_),
    .Y(_4729_)
);

NOR2X1 _11546_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [12]),
    .B(\u_fir_pe5.mul [12]),
    .Y(_4730_)
);

NOR2X1 _11547_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4730_),
    .B(_4729_),
    .Y(_4731_)
);

NAND2X1 _11548_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4731_),
    .B(_4726_),
    .Y(_4732_)
);

OR2X2 _11549_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4726_),
    .B(_4731_),
    .Y(_4733_)
);

AND2X2 _11550_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4733_),
    .B(_4732_),
    .Y(_4775_[12])
);

OAI21X1 _11551_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4727_),
    .B(_4728_),
    .C(_4732_),
    .Y(_4734_)
);

INVX1 _11552_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [13]),
    .Y(_4736_)
);

INVX1 _11553_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.mul [13]),
    .Y(_4737_)
);

NOR2X1 _11554_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4736_),
    .B(_4737_),
    .Y(_4738_)
);

NOR2X1 _11555_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [13]),
    .B(\u_fir_pe5.mul [13]),
    .Y(_4739_)
);

NOR2X1 _11556_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4739_),
    .B(_4738_),
    .Y(_4740_)
);

NAND2X1 _11557_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4740_),
    .B(_4734_),
    .Y(_4741_)
);

OR2X2 _11558_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4734_),
    .B(_4740_),
    .Y(_4742_)
);

AND2X2 _11559_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4742_),
    .B(_4741_),
    .Y(_4775_[13])
);

OAI21X1 _11560_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4736_),
    .B(_4737_),
    .C(_4741_),
    .Y(_4743_)
);

INVX1 _11561_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [14]),
    .Y(_4744_)
);

INVX1 _11562_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.mul [14]),
    .Y(_4746_)
);

NOR2X1 _11563_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4744_),
    .B(_4746_),
    .Y(_4747_)
);

NOR2X1 _11564_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [14]),
    .B(\u_fir_pe5.mul [14]),
    .Y(_4748_)
);

NOR2X1 _11565_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4748_),
    .B(_4747_),
    .Y(_4749_)
);

AND2X2 _11566_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4743_),
    .B(_4749_),
    .Y(_4750_)
);

NOR2X1 _11567_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4749_),
    .B(_4743_),
    .Y(_4751_)
);

NOR2X1 _11568_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4751_),
    .B(_4750_),
    .Y(_4775_[14])
);

INVX1 _11569_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4747_),
    .Y(_4752_)
);

NAND2X1 _11570_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4749_),
    .B(_4743_),
    .Y(_4753_)
);

NAND2X1 _11571_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [15]),
    .B(\u_fir_pe5.mul [15]),
    .Y(_4754_)
);

OR2X2 _11572_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [15]),
    .B(\u_fir_pe5.mul [15]),
    .Y(_4756_)
);

NAND2X1 _11573_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4754_),
    .B(_4756_),
    .Y(_4757_)
);

INVX1 _11574_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4757_),
    .Y(_4758_)
);

NAND3X1 _11575_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4752_),
    .B(_4758_),
    .C(_4753_),
    .Y(_4759_)
);

OAI21X1 _11576_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4747_),
    .B(_4750_),
    .C(_4757_),
    .Y(_4760_)
);

NAND2X1 _11577_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4759_),
    .B(_4760_),
    .Y(_4775_[15])
);

NOR2X1 _11578_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe5.rYin [0]),
    .B(\u_fir_pe5.mul [0]),
    .Y(_4761_)
);

NOR2X1 _11579_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4761_),
    .B(_4616_),
    .Y(_4774_[0])
);

AOI21X1 _11580_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[5] [0]),
    .B(gnd),
    .C(_4685_),
    .Y(_4762_)
);

NOR2X1 _11581_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4762_),
    .B(_4705_),
    .Y(_4777_[1])
);

NOR2X1 _11582_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4705_),
    .B(_4769_),
    .Y(_4764_)
);

NOR2X1 _11583_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4764_),
    .B(_4771_),
    .Y(_4778_[2])
);

DFFPOSX1 _11584_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_4774_[0]),
    .Q(\Y[6] [0])
);

DFFPOSX1 _11585_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_4775_[1]),
    .Q(\Y[6] [1])
);

DFFPOSX1 _11586_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf57),
    .D(_4775_[2]),
    .Q(\Y[6] [2])
);

DFFPOSX1 _11587_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf56),
    .D(_4775_[3]),
    .Q(\Y[6] [3])
);

DFFPOSX1 _11588_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf55),
    .D(_4775_[4]),
    .Q(\Y[6] [4])
);

DFFPOSX1 _11589_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf54),
    .D(_4775_[5]),
    .Q(\Y[6] [5])
);

DFFPOSX1 _11590_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf53),
    .D(_4775_[6]),
    .Q(\Y[6] [6])
);

DFFPOSX1 _11591_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf52),
    .D(_4775_[7]),
    .Q(\Y[6] [7])
);

DFFPOSX1 _11592_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf51),
    .D(_4775_[8]),
    .Q(\Y[6] [8])
);

DFFPOSX1 _11593_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf50),
    .D(_4775_[9]),
    .Q(\Y[6] [9])
);

DFFPOSX1 _11594_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf49),
    .D(_4775_[10]),
    .Q(\Y[6] [10])
);

DFFPOSX1 _11595_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf48),
    .D(_4775_[11]),
    .Q(\Y[6] [11])
);

DFFPOSX1 _11596_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf47),
    .D(_4775_[12]),
    .Q(\Y[6] [12])
);

DFFPOSX1 _11597_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf46),
    .D(_4775_[13]),
    .Q(\Y[6] [13])
);

DFFPOSX1 _11598_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf45),
    .D(_4775_[14]),
    .Q(\Y[6] [14])
);

DFFPOSX1 _11599_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf44),
    .D(_4775_[15]),
    .Q(\Y[6] [15])
);

DFFPOSX1 _11600_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf43),
    .D(\X[5] [0]),
    .Q(\X[6] [0])
);

DFFPOSX1 _11601_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf42),
    .D(\X[5] [1]),
    .Q(\X[6] [1])
);

DFFPOSX1 _11602_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf41),
    .D(\X[5] [2]),
    .Q(\X[6] [2])
);

DFFPOSX1 _11603_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf40),
    .D(\X[5] [3]),
    .Q(\X[6] [3])
);

DFFPOSX1 _11604_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf39),
    .D(\X[5] [4]),
    .Q(\X[6] [4])
);

DFFPOSX1 _11605_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf38),
    .D(\X[5]_5_bF$buf3 ),
    .Q(\X[6] [5])
);

DFFPOSX1 _11606_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf37),
    .D(\X[5] [6]),
    .Q(\X[6] [6])
);

DFFPOSX1 _11607_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf36),
    .D(\X[5] [7]),
    .Q(\X[6] [7])
);

DFFPOSX1 _11608_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf35),
    .D(\Y[5] [0]),
    .Q(\u_fir_pe5.rYin [0])
);

DFFPOSX1 _11609_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf34),
    .D(\Y[5] [1]),
    .Q(\u_fir_pe5.rYin [1])
);

DFFPOSX1 _11610_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf33),
    .D(\Y[5] [2]),
    .Q(\u_fir_pe5.rYin [2])
);

DFFPOSX1 _11611_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf32),
    .D(\Y[5] [3]),
    .Q(\u_fir_pe5.rYin [3])
);

DFFPOSX1 _11612_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf31),
    .D(\Y[5] [4]),
    .Q(\u_fir_pe5.rYin [4])
);

DFFPOSX1 _11613_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf30),
    .D(\Y[5] [5]),
    .Q(\u_fir_pe5.rYin [5])
);

DFFPOSX1 _11614_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf29),
    .D(\Y[5] [6]),
    .Q(\u_fir_pe5.rYin [6])
);

DFFPOSX1 _11615_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf28),
    .D(\Y[5] [7]),
    .Q(\u_fir_pe5.rYin [7])
);

DFFPOSX1 _11616_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf27),
    .D(\Y[5] [8]),
    .Q(\u_fir_pe5.rYin [8])
);

DFFPOSX1 _11617_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf26),
    .D(\Y[5] [9]),
    .Q(\u_fir_pe5.rYin [9])
);

DFFPOSX1 _11618_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf25),
    .D(\Y[5] [10]),
    .Q(\u_fir_pe5.rYin [10])
);

DFFPOSX1 _11619_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf24),
    .D(\Y[5] [11]),
    .Q(\u_fir_pe5.rYin [11])
);

DFFPOSX1 _11620_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf23),
    .D(\Y[5] [12]),
    .Q(\u_fir_pe5.rYin [12])
);

DFFPOSX1 _11621_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf22),
    .D(\Y[5] [13]),
    .Q(\u_fir_pe5.rYin [13])
);

DFFPOSX1 _11622_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf21),
    .D(\Y[5] [14]),
    .Q(\u_fir_pe5.rYin [14])
);

DFFPOSX1 _11623_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf20),
    .D(\Y[5] [15]),
    .Q(\u_fir_pe5.rYin [15])
);

DFFPOSX1 _11624_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf19),
    .D(_4776_[0]),
    .Q(\u_fir_pe5.mul [0])
);

DFFPOSX1 _11625_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf18),
    .D(_4777_[1]),
    .Q(\u_fir_pe5.mul [1])
);

DFFPOSX1 _11626_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf17),
    .D(_4778_[2]),
    .Q(\u_fir_pe5.mul [2])
);

DFFPOSX1 _11627_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf16),
    .D(_4779_[3]),
    .Q(\u_fir_pe5.mul [3])
);

DFFPOSX1 _11628_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf15),
    .D(_4780_[4]),
    .Q(\u_fir_pe5.mul [4])
);

DFFPOSX1 _11629_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf14),
    .D(_4781_[5]),
    .Q(\u_fir_pe5.mul [5])
);

DFFPOSX1 _11630_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf13),
    .D(_4781_[6]),
    .Q(\u_fir_pe5.mul [6])
);

DFFPOSX1 _11631_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf12),
    .D(_4781_[7]),
    .Q(\u_fir_pe5.mul [7])
);

DFFPOSX1 _11632_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf11),
    .D(_4781_[8]),
    .Q(\u_fir_pe5.mul [8])
);

DFFPOSX1 _11633_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf10),
    .D(_4781_[9]),
    .Q(\u_fir_pe5.mul [9])
);

DFFPOSX1 _11634_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf9),
    .D(_4781_[10]),
    .Q(\u_fir_pe5.mul [10])
);

DFFPOSX1 _11635_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf8),
    .D(_4781_[11]),
    .Q(\u_fir_pe5.mul [11])
);

DFFPOSX1 _11636_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf7),
    .D(_4781_[12]),
    .Q(\u_fir_pe5.mul [12])
);

DFFPOSX1 _11637_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_4781_[13]),
    .Q(\u_fir_pe5.mul [13])
);

DFFPOSX1 _11638_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_4781_[14]),
    .Q(\u_fir_pe5.mul [14])
);

DFFPOSX1 _11639_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_4781_[15]),
    .Q(\u_fir_pe5.mul [15])
);

NAND2X1 _11640_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [0]),
    .B(gnd),
    .Y(_5471_)
);

AND2X2 _11641_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [1]),
    .B(gnd),
    .Y(_5482_)
);

INVX1 _11642_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5482_),
    .Y(_5492_)
);

NOR2X1 _11643_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5471_),
    .B(_5492_),
    .Y(_5502_)
);

NAND2X1 _11644_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[7] [1]),
    .Y(_5513_)
);

NOR2X1 _11645_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5471_),
    .B(_5513_),
    .Y(_5522_)
);

AOI22X1 _11646_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [0]),
    .B(vdd),
    .C(\X[7] [1]),
    .D(gnd),
    .Y(_5532_)
);

NOR2X1 _11647_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5532_),
    .B(_5522_),
    .Y(_5542_)
);

INVX1 _11648_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [2]),
    .Y(_5552_)
);

INVX2 _11649_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_5560_)
);

NOR2X1 _11650_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5552_),
    .B(_5560_),
    .Y(_5562_)
);

NAND2X1 _11651_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5562_),
    .B(_5542_),
    .Y(_5563_)
);

INVX1 _11652_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5563_),
    .Y(_5564_)
);

NOR2X1 _11653_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5562_),
    .B(_5542_),
    .Y(_5565_)
);

NOR2X1 _11654_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5565_),
    .B(_5564_),
    .Y(_5566_)
);

NAND2X1 _11655_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5502_),
    .B(_5566_),
    .Y(_5567_)
);

INVX1 _11656_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5567_),
    .Y(_5568_)
);

NAND2X1 _11657_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [3]),
    .Y(_5569_)
);

INVX1 _11658_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5569_),
    .Y(_5570_)
);

NAND2X1 _11659_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [2]),
    .Y(_4782_)
);

INVX1 _11660_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4782_),
    .Y(_4783_)
);

NAND2X1 _11661_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [0]),
    .Y(_4784_)
);

OR2X2 _11662_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5513_),
    .B(_4784_),
    .Y(_4785_)
);

AOI22X1 _11663_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [0]),
    .C(vdd),
    .D(\X[7] [1]),
    .Y(_4786_)
);

INVX1 _11664_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4786_),
    .Y(_4787_)
);

NAND3X1 _11665_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4783_),
    .B(_4787_),
    .C(_4785_),
    .Y(_4788_)
);

NOR2X1 _11666_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5513_),
    .B(_4784_),
    .Y(_4789_)
);

OAI21X1 _11667_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4786_),
    .B(_4789_),
    .C(_4782_),
    .Y(_4790_)
);

NAND3X1 _11668_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5522_),
    .B(_4790_),
    .C(_4788_),
    .Y(_4791_)
);

INVX1 _11669_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5522_),
    .Y(_4792_)
);

NAND3X1 _11670_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4782_),
    .B(_4787_),
    .C(_4785_),
    .Y(_4793_)
);

OAI21X1 _11671_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4786_),
    .B(_4789_),
    .C(_4783_),
    .Y(_4794_)
);

NAND3X1 _11672_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4792_),
    .B(_4794_),
    .C(_4793_),
    .Y(_4795_)
);

NAND3X1 _11673_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5570_),
    .B(_4795_),
    .C(_4791_),
    .Y(_4796_)
);

INVX2 _11674_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [3]),
    .Y(_4797_)
);

NAND2X1 _11675_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4795_),
    .B(_4791_),
    .Y(_4798_)
);

OAI21X1 _11676_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5560_),
    .B(_4797_),
    .C(_4798_),
    .Y(_4799_)
);

NAND2X1 _11677_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4796_),
    .B(_4799_),
    .Y(_4800_)
);

NAND2X1 _11678_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5563_),
    .B(_4800_),
    .Y(_4801_)
);

NAND3X1 _11679_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5564_),
    .B(_4796_),
    .C(_4799_),
    .Y(_4802_)
);

NAND3X1 _11680_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4802_),
    .B(_5568_),
    .C(_4801_),
    .Y(_4803_)
);

INVX1 _11681_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4803_),
    .Y(_4804_)
);

AOI21X1 _11682_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4801_),
    .B(_4802_),
    .C(_5568_),
    .Y(_4805_)
);

NOR2X1 _11683_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4805_),
    .B(_4804_),
    .Y(_5576_[3])
);

NAND2X1 _11684_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [0]),
    .B(gnd),
    .Y(_4806_)
);

NAND2X1 _11685_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [4]),
    .B(gnd),
    .Y(_4807_)
);

NOR2X1 _11686_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4806_),
    .B(_4807_),
    .Y(_4808_)
);

AOI22X1 _11687_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [0]),
    .B(gnd),
    .C(gnd),
    .D(\X[7] [4]),
    .Y(_4809_)
);

NOR2X1 _11688_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4809_),
    .B(_4808_),
    .Y(_4810_)
);

INVX1 _11689_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4810_),
    .Y(_4811_)
);

NAND2X1 _11690_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [0]),
    .B(vdd),
    .Y(_4812_)
);

NAND2X1 _11691_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [1]),
    .Y(_4813_)
);

OAI22X1 _11692_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4812_),
    .B(_4813_),
    .C(_4782_),
    .D(_4786_),
    .Y(_4814_)
);

NAND2X1 _11693_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [3]),
    .Y(_4815_)
);

INVX1 _11694_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4815_),
    .Y(_4816_)
);

AND2X2 _11695_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[7] [1]),
    .Y(_4817_)
);

AND2X2 _11696_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [2]),
    .Y(_4818_)
);

NAND2X1 _11697_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4817_),
    .B(_4818_),
    .Y(_4819_)
);

AOI22X1 _11698_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [1]),
    .C(vdd),
    .D(\X[7] [2]),
    .Y(_4820_)
);

INVX1 _11699_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4820_),
    .Y(_4821_)
);

NAND3X1 _11700_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4816_),
    .B(_4821_),
    .C(_4819_),
    .Y(_4822_)
);

NAND3X1 _11701_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[7] [2]),
    .C(_4813_),
    .Y(_4823_)
);

NAND2X1 _11702_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[7] [2]),
    .Y(_4824_)
);

NAND3X1 _11703_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [1]),
    .C(_4824_),
    .Y(_4825_)
);

NAND3X1 _11704_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4815_),
    .B(_4823_),
    .C(_4825_),
    .Y(_4826_)
);

NAND3X1 _11705_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4814_),
    .B(_4826_),
    .C(_4822_),
    .Y(_4827_)
);

INVX1 _11706_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4814_),
    .Y(_4828_)
);

NAND2X1 _11707_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4826_),
    .B(_4822_),
    .Y(_4829_)
);

NAND2X1 _11708_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4828_),
    .B(_4829_),
    .Y(_4830_)
);

NAND3X1 _11709_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4811_),
    .B(_4827_),
    .C(_4830_),
    .Y(_4831_)
);

NAND2X1 _11710_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4814_),
    .B(_4829_),
    .Y(_4832_)
);

NAND3X1 _11711_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4822_),
    .B(_4826_),
    .C(_4828_),
    .Y(_4833_)
);

NAND3X1 _11712_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4810_),
    .B(_4833_),
    .C(_4832_),
    .Y(_4834_)
);

AOI22X1 _11713_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4791_),
    .B(_4796_),
    .C(_4831_),
    .D(_4834_),
    .Y(_4835_)
);

INVX1 _11714_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4835_),
    .Y(_4836_)
);

NAND2X1 _11715_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4791_),
    .B(_4796_),
    .Y(_4837_)
);

NAND2X1 _11716_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4831_),
    .B(_4834_),
    .Y(_4838_)
);

OR2X2 _11717_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4838_),
    .B(_4837_),
    .Y(_4839_)
);

NAND2X1 _11718_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4836_),
    .B(_4839_),
    .Y(_4840_)
);

OAI21X1 _11719_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5563_),
    .B(_4800_),
    .C(_4803_),
    .Y(_4841_)
);

OR2X2 _11720_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4841_),
    .B(_4840_),
    .Y(_4842_)
);

NAND3X1 _11721_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4810_),
    .B(_4827_),
    .C(_4830_),
    .Y(_4843_)
);

INVX1 _11722_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4827_),
    .Y(_4844_)
);

AOI21X1 _11723_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4822_),
    .B(_4826_),
    .C(_4814_),
    .Y(_4845_)
);

OAI21X1 _11724_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4845_),
    .B(_4844_),
    .C(_4811_),
    .Y(_4846_)
);

AOI21X1 _11725_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4843_),
    .B(_4846_),
    .C(_4837_),
    .Y(_4847_)
);

OAI21X1 _11726_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4835_),
    .B(_4847_),
    .C(_4841_),
    .Y(_4848_)
);

NAND2X1 _11727_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4848_),
    .B(_4842_),
    .Y(_5577_[4])
);

NOR2X1 _11728_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4803_),
    .B(_4840_),
    .Y(_4849_)
);

NOR3X1 _11729_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4835_),
    .B(_4802_),
    .C(_4847_),
    .Y(_4850_)
);

OAI21X1 _11730_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4811_),
    .B(_4845_),
    .C(_4827_),
    .Y(_4851_)
);

NAND2X1 _11731_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [0]),
    .B(gnd),
    .Y(_4852_)
);

INVX1 _11732_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4852_),
    .Y(_4853_)
);

AND2X2 _11733_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7]_5_bF$buf3 ),
    .Y(_4854_)
);

NAND2X1 _11734_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5482_),
    .B(_4854_),
    .Y(_4855_)
);

INVX2 _11735_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7]_5_bF$buf2 ),
    .Y(_4856_)
);

NAND2X1 _11736_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [1]),
    .B(gnd),
    .Y(_4857_)
);

OAI21X1 _11737_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5560_),
    .B(_4856_),
    .C(_4857_),
    .Y(_4858_)
);

NAND3X1 _11738_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4858_),
    .B(_4853_),
    .C(_4855_),
    .Y(_4859_)
);

NAND3X1 _11739_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7]_5_bF$buf1 ),
    .C(_4857_),
    .Y(_4860_)
);

NAND2X1 _11740_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7]_5_bF$buf0 ),
    .Y(_4861_)
);

NAND3X1 _11741_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [1]),
    .B(gnd),
    .C(_4861_),
    .Y(_4862_)
);

NAND3X1 _11742_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4852_),
    .B(_4860_),
    .C(_4862_),
    .Y(_4863_)
);

AND2X2 _11743_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4859_),
    .B(_4863_),
    .Y(_4864_)
);

NAND2X1 _11744_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [2]),
    .Y(_4865_)
);

OAI22X1 _11745_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5513_),
    .B(_4865_),
    .C(_4815_),
    .D(_4820_),
    .Y(_4866_)
);

NAND2X1 _11746_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [4]),
    .Y(_4867_)
);

INVX1 _11747_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4867_),
    .Y(_4868_)
);

AND2X2 _11748_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[7] [3]),
    .Y(_4869_)
);

NAND2X1 _11749_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4818_),
    .B(_4869_),
    .Y(_4870_)
);

INVX1 _11750_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .Y(_4871_)
);

OAI21X1 _11751_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4871_),
    .B(_4797_),
    .C(_4865_),
    .Y(_4872_)
);

NAND3X1 _11752_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4868_),
    .B(_4872_),
    .C(_4870_),
    .Y(_4873_)
);

NAND3X1 _11753_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[7] [3]),
    .C(_4865_),
    .Y(_4874_)
);

NAND2X1 _11754_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[7] [3]),
    .Y(_4875_)
);

NAND3X1 _11755_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [2]),
    .C(_4875_),
    .Y(_4876_)
);

NAND3X1 _11756_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4867_),
    .B(_4874_),
    .C(_4876_),
    .Y(_4877_)
);

NAND3X1 _11757_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4866_),
    .B(_4877_),
    .C(_4873_),
    .Y(_4878_)
);

INVX1 _11758_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4866_),
    .Y(_4879_)
);

AOI21X1 _11759_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4874_),
    .B(_4876_),
    .C(_4867_),
    .Y(_4880_)
);

AOI22X1 _11760_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [4]),
    .C(_4870_),
    .D(_4872_),
    .Y(_4881_)
);

OAI21X1 _11761_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4880_),
    .B(_4881_),
    .C(_4879_),
    .Y(_4882_)
);

NAND3X1 _11762_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4878_),
    .B(_4864_),
    .C(_4882_),
    .Y(_4883_)
);

NAND2X1 _11763_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4863_),
    .B(_4859_),
    .Y(_4884_)
);

OAI21X1 _11764_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4880_),
    .B(_4881_),
    .C(_4866_),
    .Y(_4885_)
);

NAND3X1 _11765_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4877_),
    .B(_4873_),
    .C(_4879_),
    .Y(_4886_)
);

NAND3X1 _11766_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4884_),
    .B(_4886_),
    .C(_4885_),
    .Y(_4887_)
);

NAND3X1 _11767_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4883_),
    .B(_4887_),
    .C(_4851_),
    .Y(_4888_)
);

AOI21X1 _11768_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4810_),
    .B(_4830_),
    .C(_4844_),
    .Y(_4889_)
);

AOI21X1 _11769_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4885_),
    .B(_4886_),
    .C(_4884_),
    .Y(_4890_)
);

AOI21X1 _11770_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4882_),
    .B(_4878_),
    .C(_4864_),
    .Y(_4891_)
);

OAI21X1 _11771_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4890_),
    .B(_4891_),
    .C(_4889_),
    .Y(_4892_)
);

NAND3X1 _11772_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4808_),
    .B(_4888_),
    .C(_4892_),
    .Y(_4893_)
);

INVX1 _11773_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4808_),
    .Y(_4894_)
);

OAI21X1 _11774_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4890_),
    .B(_4891_),
    .C(_4851_),
    .Y(_4895_)
);

NAND3X1 _11775_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4883_),
    .B(_4887_),
    .C(_4889_),
    .Y(_4896_)
);

NAND3X1 _11776_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4894_),
    .B(_4895_),
    .C(_4896_),
    .Y(_4897_)
);

NAND3X1 _11777_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4835_),
    .B(_4893_),
    .C(_4897_),
    .Y(_4898_)
);

NAND3X1 _11778_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4894_),
    .B(_4888_),
    .C(_4892_),
    .Y(_4899_)
);

NAND3X1 _11779_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4808_),
    .B(_4895_),
    .C(_4896_),
    .Y(_4900_)
);

NAND3X1 _11780_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4836_),
    .B(_4899_),
    .C(_4900_),
    .Y(_4901_)
);

NAND3X1 _11781_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4898_),
    .B(_4901_),
    .C(_4850_),
    .Y(_4902_)
);

INVX1 _11782_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4802_),
    .Y(_4903_)
);

NAND3X1 _11783_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4903_),
    .B(_4836_),
    .C(_4839_),
    .Y(_4904_)
);

NAND3X1 _11784_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4836_),
    .B(_4893_),
    .C(_4897_),
    .Y(_4905_)
);

NAND3X1 _11785_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4835_),
    .B(_4899_),
    .C(_4900_),
    .Y(_4906_)
);

NAND3X1 _11786_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4905_),
    .B(_4906_),
    .C(_4904_),
    .Y(_4907_)
);

NAND3X1 _11787_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4902_),
    .B(_4907_),
    .C(_4849_),
    .Y(_4908_)
);

INVX1 _11788_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4849_),
    .Y(_4909_)
);

INVX1 _11789_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4902_),
    .Y(_4910_)
);

INVX1 _11790_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4907_),
    .Y(_4911_)
);

OAI21X1 _11791_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4910_),
    .B(_4911_),
    .C(_4909_),
    .Y(_4912_)
);

AND2X2 _11792_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4912_),
    .B(_4908_),
    .Y(_5578_[5])
);

AND2X2 _11793_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [0]),
    .B(gnd),
    .Y(_4913_)
);

NAND2X1 _11794_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7]_5_bF$buf3 ),
    .Y(_4914_)
);

OAI21X1 _11795_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5492_),
    .B(_4914_),
    .C(_4859_),
    .Y(_4915_)
);

OR2X2 _11796_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4915_),
    .B(_4913_),
    .Y(_4916_)
);

NAND2X1 _11797_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4913_),
    .B(_4915_),
    .Y(_4917_)
);

NAND2X1 _11798_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4917_),
    .B(_4916_),
    .Y(_4918_)
);

AOI21X1 _11799_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4873_),
    .B(_4877_),
    .C(_4866_),
    .Y(_4919_)
);

OAI21X1 _11800_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4884_),
    .B(_4919_),
    .C(_4878_),
    .Y(_4920_)
);

NAND2X1 _11801_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [1]),
    .B(gnd),
    .Y(_4921_)
);

INVX1 _11802_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4921_),
    .Y(_4922_)
);

AND2X2 _11803_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [2]),
    .B(gnd),
    .Y(_4923_)
);

AND2X2 _11804_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [6]),
    .Y(_4924_)
);

NAND2X1 _11805_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4923_),
    .B(_4924_),
    .Y(_4925_)
);

INVX2 _11806_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [6]),
    .Y(_4926_)
);

NAND2X1 _11807_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [2]),
    .B(gnd),
    .Y(_4927_)
);

OAI21X1 _11808_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5560_),
    .B(_4926_),
    .C(_4927_),
    .Y(_4928_)
);

NAND3X1 _11809_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4928_),
    .B(_4922_),
    .C(_4925_),
    .Y(_4929_)
);

NAND3X1 _11810_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [6]),
    .C(_4927_),
    .Y(_4930_)
);

NAND2X1 _11811_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [6]),
    .Y(_4931_)
);

NAND2X1 _11812_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4931_),
    .B(_4923_),
    .Y(_4932_)
);

NAND3X1 _11813_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4921_),
    .B(_4930_),
    .C(_4932_),
    .Y(_4933_)
);

AND2X2 _11814_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4929_),
    .B(_4933_),
    .Y(_4934_)
);

NAND2X1 _11815_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [3]),
    .Y(_4935_)
);

AOI22X1 _11816_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [2]),
    .C(vdd),
    .D(\X[7] [3]),
    .Y(_4936_)
);

OAI22X1 _11817_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4824_),
    .B(_4935_),
    .C(_4867_),
    .D(_4936_),
    .Y(_4937_)
);

NAND2X1 _11818_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7]_5_bF$buf2 ),
    .Y(_4938_)
);

INVX1 _11819_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4938_),
    .Y(_4939_)
);

AND2X2 _11820_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [4]),
    .Y(_4940_)
);

NAND2X1 _11821_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4869_),
    .B(_4940_),
    .Y(_4941_)
);

AOI22X1 _11822_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [3]),
    .C(vdd),
    .D(\X[7] [4]),
    .Y(_4942_)
);

INVX1 _11823_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4942_),
    .Y(_4943_)
);

NAND3X1 _11824_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4939_),
    .B(_4943_),
    .C(_4941_),
    .Y(_4944_)
);

NAND3X1 _11825_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[7] [4]),
    .C(_4935_),
    .Y(_4945_)
);

NAND2X1 _11826_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[7] [4]),
    .Y(_4946_)
);

NAND3X1 _11827_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [3]),
    .C(_4946_),
    .Y(_4947_)
);

NAND3X1 _11828_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4938_),
    .B(_4945_),
    .C(_4947_),
    .Y(_4948_)
);

NAND3X1 _11829_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4937_),
    .B(_4948_),
    .C(_4944_),
    .Y(_4949_)
);

INVX1 _11830_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4937_),
    .Y(_4950_)
);

AOI21X1 _11831_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4945_),
    .B(_4947_),
    .C(_4938_),
    .Y(_4951_)
);

AOI22X1 _11832_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7]_5_bF$buf1 ),
    .C(_4941_),
    .D(_4943_),
    .Y(_4952_)
);

OAI21X1 _11833_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4951_),
    .B(_4952_),
    .C(_4950_),
    .Y(_4953_)
);

NAND3X1 _11834_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4949_),
    .B(_4934_),
    .C(_4953_),
    .Y(_4954_)
);

NAND2X1 _11835_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4933_),
    .B(_4929_),
    .Y(_4955_)
);

OAI21X1 _11836_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4951_),
    .B(_4952_),
    .C(_4937_),
    .Y(_4956_)
);

NAND3X1 _11837_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4944_),
    .B(_4948_),
    .C(_4950_),
    .Y(_4957_)
);

NAND3X1 _11838_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4955_),
    .B(_4957_),
    .C(_4956_),
    .Y(_4958_)
);

NAND3X1 _11839_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4954_),
    .B(_4920_),
    .C(_4958_),
    .Y(_4959_)
);

INVX1 _11840_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4878_),
    .Y(_4960_)
);

AOI21X1 _11841_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4864_),
    .B(_4882_),
    .C(_4960_),
    .Y(_4961_)
);

AOI21X1 _11842_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4956_),
    .B(_4957_),
    .C(_4955_),
    .Y(_4962_)
);

AOI21X1 _11843_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4953_),
    .B(_4949_),
    .C(_4934_),
    .Y(_4963_)
);

OAI21X1 _11844_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4962_),
    .B(_4963_),
    .C(_4961_),
    .Y(_4964_)
);

NAND3X1 _11845_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4918_),
    .B(_4959_),
    .C(_4964_),
    .Y(_4965_)
);

AND2X2 _11846_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4916_),
    .B(_4917_),
    .Y(_4966_)
);

OAI21X1 _11847_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4962_),
    .B(_4963_),
    .C(_4920_),
    .Y(_4967_)
);

NAND3X1 _11848_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4954_),
    .B(_4958_),
    .C(_4961_),
    .Y(_4968_)
);

NAND3X1 _11849_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4966_),
    .B(_4967_),
    .C(_4968_),
    .Y(_4969_)
);

AOI22X1 _11850_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4893_),
    .B(_4888_),
    .C(_4965_),
    .D(_4969_),
    .Y(_4970_)
);

AOI21X1 _11851_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4883_),
    .B(_4887_),
    .C(_4851_),
    .Y(_4971_)
);

OAI21X1 _11852_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4894_),
    .B(_4971_),
    .C(_4888_),
    .Y(_4972_)
);

NAND3X1 _11853_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4966_),
    .B(_4959_),
    .C(_4964_),
    .Y(_4973_)
);

NAND3X1 _11854_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4918_),
    .B(_4967_),
    .C(_4968_),
    .Y(_4974_)
);

AOI21X1 _11855_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4974_),
    .B(_4973_),
    .C(_4972_),
    .Y(_4975_)
);

OAI21X1 _11856_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4975_),
    .B(_4970_),
    .C(_4898_),
    .Y(_4976_)
);

AOI21X1 _11857_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4900_),
    .B(_4899_),
    .C(_4836_),
    .Y(_4977_)
);

NAND3X1 _11858_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4972_),
    .B(_4973_),
    .C(_4974_),
    .Y(_4978_)
);

INVX1 _11859_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4888_),
    .Y(_4979_)
);

AOI21X1 _11860_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4808_),
    .B(_4892_),
    .C(_4979_),
    .Y(_4980_)
);

AOI21X1 _11861_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4968_),
    .B(_4967_),
    .C(_4918_),
    .Y(_4981_)
);

AOI21X1 _11862_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4964_),
    .B(_4959_),
    .C(_4966_),
    .Y(_4982_)
);

OAI21X1 _11863_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4981_),
    .B(_4982_),
    .C(_4980_),
    .Y(_4983_)
);

NAND3X1 _11864_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4977_),
    .B(_4978_),
    .C(_4983_),
    .Y(_4984_)
);

NAND2X1 _11865_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4984_),
    .B(_4976_),
    .Y(_4985_)
);

AOI21X1 _11866_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4902_),
    .B(_4908_),
    .C(_4985_),
    .Y(_4986_)
);

OAI21X1 _11867_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4911_),
    .B(_4909_),
    .C(_4902_),
    .Y(_4987_)
);

AOI21X1 _11868_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4976_),
    .B(_4984_),
    .C(_4987_),
    .Y(_4988_)
);

NOR2X1 _11869_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4986_),
    .B(_4988_),
    .Y(_5578_[6])
);

INVX1 _11870_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4984_),
    .Y(_4989_)
);

AOI21X1 _11871_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4954_),
    .B(_4958_),
    .C(_4920_),
    .Y(_4990_)
);

OAI21X1 _11872_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4918_),
    .B(_4990_),
    .C(_4959_),
    .Y(_4991_)
);

NAND2X1 _11873_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [0]),
    .B(gnd),
    .Y(_4992_)
);

INVX1 _11874_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4992_),
    .Y(_4993_)
);

NAND2X1 _11875_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [1]),
    .B(gnd),
    .Y(_4994_)
);

INVX1 _11876_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4994_),
    .Y(_4995_)
);

AND2X2 _11877_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4927_),
    .B(_4931_),
    .Y(_4996_)
);

OAI21X1 _11878_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4921_),
    .B(_4996_),
    .C(_4925_),
    .Y(_4997_)
);

NAND2X1 _11879_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4995_),
    .B(_4997_),
    .Y(_4998_)
);

NAND3X1 _11880_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4925_),
    .B(_4994_),
    .C(_4929_),
    .Y(_4999_)
);

NAND3X1 _11881_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4993_),
    .B(_4999_),
    .C(_4998_),
    .Y(_5000_)
);

AOI21X1 _11882_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4929_),
    .B(_4925_),
    .C(_4994_),
    .Y(_5001_)
);

NOR2X1 _11883_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4995_),
    .B(_4997_),
    .Y(_5002_)
);

OAI21X1 _11884_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5001_),
    .B(_5002_),
    .C(_4992_),
    .Y(_5003_)
);

NAND2X1 _11885_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5000_),
    .B(_5003_),
    .Y(_5004_)
);

AOI21X1 _11886_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4944_),
    .B(_4948_),
    .C(_4937_),
    .Y(_5005_)
);

OAI21X1 _11887_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4955_),
    .B(_5005_),
    .C(_4949_),
    .Y(_5006_)
);

NAND2X1 _11888_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [2]),
    .B(gnd),
    .Y(_5007_)
);

INVX1 _11889_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5007_),
    .Y(_5008_)
);

AND2X2 _11890_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [3]),
    .B(gnd),
    .Y(_5009_)
);

AND2X2 _11891_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [7]),
    .Y(_5010_)
);

NAND2X1 _11892_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5009_),
    .B(_5010_),
    .Y(_5011_)
);

AOI22X1 _11893_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [7]),
    .C(\X[7] [3]),
    .D(gnd),
    .Y(_5012_)
);

INVX1 _11894_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5012_),
    .Y(_5013_)
);

NAND3X1 _11895_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5008_),
    .B(_5013_),
    .C(_5011_),
    .Y(_5014_)
);

INVX1 _11896_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_5015_)
);

OAI21X1 _11897_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4797_),
    .B(_5015_),
    .C(_5010_),
    .Y(_5016_)
);

INVX1 _11898_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [7]),
    .Y(_5017_)
);

OAI21X1 _11899_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5560_),
    .B(_5017_),
    .C(_5009_),
    .Y(_5018_)
);

NAND3X1 _11900_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5007_),
    .B(_5016_),
    .C(_5018_),
    .Y(_5019_)
);

NAND2X1 _11901_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5014_),
    .B(_5019_),
    .Y(_5020_)
);

OAI21X1 _11902_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4938_),
    .B(_4942_),
    .C(_4941_),
    .Y(_5021_)
);

NAND2X1 _11903_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [6]),
    .Y(_5022_)
);

NAND2X1 _11904_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [4]),
    .Y(_5023_)
);

AND2X2 _11905_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[7]_5_bF$buf0 ),
    .Y(_5024_)
);

NAND2X1 _11906_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5023_),
    .B(_5024_),
    .Y(_5025_)
);

OAI21X1 _11907_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4871_),
    .B(_4856_),
    .C(_4940_),
    .Y(_5026_)
);

AOI21X1 _11908_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5026_),
    .B(_5025_),
    .C(_5022_),
    .Y(_5027_)
);

INVX1 _11909_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5022_),
    .Y(_5028_)
);

NAND2X1 _11910_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4940_),
    .B(_5024_),
    .Y(_5029_)
);

AOI22X1 _11911_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [4]),
    .C(vdd),
    .D(\X[7]_5_bF$buf3 ),
    .Y(_5030_)
);

INVX1 _11912_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5030_),
    .Y(_5031_)
);

AOI21X1 _11913_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5029_),
    .B(_5031_),
    .C(_5028_),
    .Y(_5032_)
);

OAI21X1 _11914_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5032_),
    .B(_5027_),
    .C(_5021_),
    .Y(_5033_)
);

AOI22X1 _11915_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4869_),
    .B(_4940_),
    .C(_4943_),
    .D(_4939_),
    .Y(_5034_)
);

NAND3X1 _11916_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5028_),
    .B(_5031_),
    .C(_5029_),
    .Y(_5035_)
);

NAND2X1 _11917_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[7]_5_bF$buf2 ),
    .Y(_5036_)
);

NOR2X1 _11918_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5023_),
    .B(_5036_),
    .Y(_5037_)
);

OAI21X1 _11919_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5030_),
    .B(_5037_),
    .C(_5022_),
    .Y(_5038_)
);

NAND3X1 _11920_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5035_),
    .B(_5034_),
    .C(_5038_),
    .Y(_5039_)
);

AOI21X1 _11921_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5033_),
    .B(_5039_),
    .C(_5020_),
    .Y(_5040_)
);

AND2X2 _11922_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5019_),
    .B(_5014_),
    .Y(_5041_)
);

NAND3X1 _11923_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5021_),
    .B(_5035_),
    .C(_5038_),
    .Y(_5042_)
);

OAI21X1 _11924_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5032_),
    .B(_5027_),
    .C(_5034_),
    .Y(_5043_)
);

AOI21X1 _11925_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5043_),
    .B(_5042_),
    .C(_5041_),
    .Y(_5044_)
);

OAI21X1 _11926_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5040_),
    .B(_5044_),
    .C(_5006_),
    .Y(_5045_)
);

INVX1 _11927_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4949_),
    .Y(_5046_)
);

AOI21X1 _11928_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4934_),
    .B(_4953_),
    .C(_5046_),
    .Y(_5047_)
);

NAND3X1 _11929_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5042_),
    .B(_5041_),
    .C(_5043_),
    .Y(_5048_)
);

NAND3X1 _11930_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5020_),
    .B(_5039_),
    .C(_5033_),
    .Y(_5049_)
);

NAND3X1 _11931_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5048_),
    .B(_5049_),
    .C(_5047_),
    .Y(_5050_)
);

AOI21X1 _11932_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5050_),
    .B(_5045_),
    .C(_5004_),
    .Y(_5051_)
);

AND2X2 _11933_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5003_),
    .B(_5000_),
    .Y(_5052_)
);

NAND3X1 _11934_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5006_),
    .B(_5048_),
    .C(_5049_),
    .Y(_5053_)
);

OAI21X1 _11935_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5040_),
    .B(_5044_),
    .C(_5047_),
    .Y(_5054_)
);

AOI21X1 _11936_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5054_),
    .B(_5053_),
    .C(_5052_),
    .Y(_5055_)
);

OAI21X1 _11937_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5055_),
    .B(_5051_),
    .C(_4991_),
    .Y(_5056_)
);

INVX1 _11938_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4959_),
    .Y(_5057_)
);

AOI21X1 _11939_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4966_),
    .B(_4964_),
    .C(_5057_),
    .Y(_5058_)
);

NAND3X1 _11940_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5053_),
    .B(_5052_),
    .C(_5054_),
    .Y(_5059_)
);

NAND3X1 _11941_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5004_),
    .B(_5045_),
    .C(_5050_),
    .Y(_5060_)
);

NAND3X1 _11942_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5059_),
    .B(_5060_),
    .C(_5058_),
    .Y(_5061_)
);

AOI21X1 _11943_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5061_),
    .B(_5056_),
    .C(_4917_),
    .Y(_5062_)
);

INVX1 _11944_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4917_),
    .Y(_5063_)
);

NAND3X1 _11945_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4991_),
    .B(_5059_),
    .C(_5060_),
    .Y(_5064_)
);

OAI21X1 _11946_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5051_),
    .B(_5055_),
    .C(_5058_),
    .Y(_5065_)
);

AOI21X1 _11947_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5065_),
    .B(_5064_),
    .C(_5063_),
    .Y(_5066_)
);

OAI21X1 _11948_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5066_),
    .B(_5062_),
    .C(_4978_),
    .Y(_5067_)
);

NAND3X1 _11949_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5063_),
    .B(_5064_),
    .C(_5065_),
    .Y(_5068_)
);

NAND3X1 _11950_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4917_),
    .B(_5056_),
    .C(_5061_),
    .Y(_5069_)
);

NAND3X1 _11951_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4970_),
    .B(_5068_),
    .C(_5069_),
    .Y(_5070_)
);

AND2X2 _11952_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5067_),
    .B(_5070_),
    .Y(_5071_)
);

OAI21X1 _11953_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4989_),
    .B(_4986_),
    .C(_5071_),
    .Y(_5072_)
);

NOR2X1 _11954_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4989_),
    .B(_4986_),
    .Y(_5073_)
);

AOI21X1 _11955_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5069_),
    .B(_5068_),
    .C(_4970_),
    .Y(_5074_)
);

INVX1 _11956_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5070_),
    .Y(_5075_)
);

OAI21X1 _11957_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5074_),
    .B(_5075_),
    .C(_5073_),
    .Y(_5076_)
);

AND2X2 _11958_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5076_),
    .B(_5072_),
    .Y(_5578_[7])
);

NAND3X1 _11959_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5067_),
    .B(_5070_),
    .C(_4986_),
    .Y(_5077_)
);

AOI21X1 _11960_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4989_),
    .B(_5067_),
    .C(_5075_),
    .Y(_5078_)
);

NAND2X1 _11961_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5078_),
    .B(_5077_),
    .Y(_5079_)
);

INVX1 _11962_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5064_),
    .Y(_5080_)
);

AOI21X1 _11963_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5063_),
    .B(_5065_),
    .C(_5080_),
    .Y(_5081_)
);

OAI21X1 _11964_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4992_),
    .B(_5002_),
    .C(_4998_),
    .Y(_5082_)
);

INVX1 _11965_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5082_),
    .Y(_5083_)
);

AOI21X1 _11966_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5048_),
    .B(_5049_),
    .C(_5006_),
    .Y(_5084_)
);

OAI21X1 _11967_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5004_),
    .B(_5084_),
    .C(_5053_),
    .Y(_5085_)
);

NAND2X1 _11968_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [1]),
    .B(gnd),
    .Y(_5086_)
);

INVX2 _11969_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_5087_)
);

NOR2X1 _11970_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5552_),
    .B(_5087_),
    .Y(_5088_)
);

OAI21X1 _11971_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5007_),
    .B(_5012_),
    .C(_5011_),
    .Y(_5089_)
);

NOR2X1 _11972_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5088_),
    .B(_5089_),
    .Y(_5090_)
);

AND2X2 _11973_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5089_),
    .B(_5088_),
    .Y(_5091_)
);

OAI21X1 _11974_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5090_),
    .B(_5091_),
    .C(_5086_),
    .Y(_5092_)
);

INVX1 _11975_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5086_),
    .Y(_5093_)
);

OR2X2 _11976_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5089_),
    .B(_5088_),
    .Y(_5094_)
);

NAND2X1 _11977_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5088_),
    .B(_5089_),
    .Y(_5095_)
);

NAND3X1 _11978_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5093_),
    .B(_5095_),
    .C(_5094_),
    .Y(_5096_)
);

NAND2X1 _11979_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5092_),
    .B(_5096_),
    .Y(_5097_)
);

AOI21X1 _11980_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5038_),
    .B(_5035_),
    .C(_5021_),
    .Y(_5098_)
);

OAI21X1 _11981_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5020_),
    .B(_5098_),
    .C(_5042_),
    .Y(_5099_)
);

NAND2X1 _11982_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [3]),
    .B(gnd),
    .Y(_5100_)
);

INVX1 _11983_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_5101_)
);

OAI21X1 _11984_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4797_),
    .B(_5101_),
    .C(_4807_),
    .Y(_5102_)
);

NAND2X1 _11985_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [4]),
    .B(gnd),
    .Y(_5103_)
);

OAI21X1 _11986_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5100_),
    .B(_5103_),
    .C(_5102_),
    .Y(_5104_)
);

OAI21X1 _11987_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5022_),
    .B(_5030_),
    .C(_5029_),
    .Y(_5105_)
);

NAND2X1 _11988_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [7]),
    .Y(_5106_)
);

NAND2X1 _11989_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7]_5_bF$buf1 ),
    .Y(_5107_)
);

NAND3X1 _11990_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[7] [6]),
    .C(_5107_),
    .Y(_5108_)
);

AND2X2 _11991_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7]_5_bF$buf0 ),
    .Y(_5109_)
);

OAI21X1 _11992_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4871_),
    .B(_4926_),
    .C(_5109_),
    .Y(_5110_)
);

AOI21X1 _11993_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5110_),
    .B(_5108_),
    .C(_5106_),
    .Y(_5111_)
);

INVX1 _11994_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5106_),
    .Y(_5112_)
);

AND2X2 _11995_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[7] [6]),
    .Y(_5113_)
);

NAND2X1 _11996_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5109_),
    .B(_5113_),
    .Y(_5114_)
);

NAND2X1 _11997_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[7] [6]),
    .Y(_5115_)
);

NAND2X1 _11998_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5107_),
    .B(_5115_),
    .Y(_5116_)
);

AOI21X1 _11999_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5114_),
    .B(_5116_),
    .C(_5112_),
    .Y(_5117_)
);

OAI21X1 _12000_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5117_),
    .B(_5111_),
    .C(_5105_),
    .Y(_5118_)
);

AOI21X1 _12001_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5028_),
    .B(_5031_),
    .C(_5037_),
    .Y(_5119_)
);

NAND3X1 _12002_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5112_),
    .B(_5116_),
    .C(_5114_),
    .Y(_5120_)
);

NAND3X1 _12003_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5106_),
    .B(_5108_),
    .C(_5110_),
    .Y(_5121_)
);

NAND3X1 _12004_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5120_),
    .B(_5121_),
    .C(_5119_),
    .Y(_5122_)
);

AOI21X1 _12005_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5118_),
    .B(_5122_),
    .C(_5104_),
    .Y(_5123_)
);

INVX1 _12006_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5104_),
    .Y(_5124_)
);

NAND3X1 _12007_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5105_),
    .B(_5120_),
    .C(_5121_),
    .Y(_5125_)
);

OAI21X1 _12008_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5117_),
    .B(_5111_),
    .C(_5119_),
    .Y(_5126_)
);

AOI21X1 _12009_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5126_),
    .B(_5125_),
    .C(_5124_),
    .Y(_5127_)
);

OAI21X1 _12010_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5123_),
    .B(_5127_),
    .C(_5099_),
    .Y(_5128_)
);

INVX1 _12011_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5042_),
    .Y(_5129_)
);

AOI21X1 _12012_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5041_),
    .B(_5043_),
    .C(_5129_),
    .Y(_5130_)
);

NAND3X1 _12013_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5124_),
    .B(_5125_),
    .C(_5126_),
    .Y(_5131_)
);

NAND3X1 _12014_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5104_),
    .B(_5122_),
    .C(_5118_),
    .Y(_5132_)
);

NAND3X1 _12015_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5131_),
    .B(_5132_),
    .C(_5130_),
    .Y(_5133_)
);

AOI21X1 _12016_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5133_),
    .B(_5128_),
    .C(_5097_),
    .Y(_5134_)
);

AND2X2 _12017_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5096_),
    .B(_5092_),
    .Y(_5135_)
);

NAND3X1 _12018_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5131_),
    .B(_5132_),
    .C(_5099_),
    .Y(_5136_)
);

OAI21X1 _12019_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5123_),
    .B(_5127_),
    .C(_5130_),
    .Y(_5137_)
);

AOI21X1 _12020_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5137_),
    .B(_5136_),
    .C(_5135_),
    .Y(_5138_)
);

OAI21X1 _12021_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5138_),
    .B(_5134_),
    .C(_5085_),
    .Y(_5139_)
);

INVX1 _12022_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5053_),
    .Y(_5140_)
);

AOI21X1 _12023_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5052_),
    .B(_5054_),
    .C(_5140_),
    .Y(_5141_)
);

NAND3X1 _12024_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5135_),
    .B(_5136_),
    .C(_5137_),
    .Y(_5142_)
);

NAND3X1 _12025_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5097_),
    .B(_5128_),
    .C(_5133_),
    .Y(_5143_)
);

NAND3X1 _12026_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5142_),
    .B(_5143_),
    .C(_5141_),
    .Y(_5144_)
);

AOI21X1 _12027_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5139_),
    .B(_5144_),
    .C(_5083_),
    .Y(_5145_)
);

NAND3X1 _12028_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5085_),
    .B(_5142_),
    .C(_5143_),
    .Y(_5146_)
);

OAI21X1 _12029_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5138_),
    .B(_5134_),
    .C(_5141_),
    .Y(_5147_)
);

AOI21X1 _12030_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5147_),
    .B(_5146_),
    .C(_5082_),
    .Y(_5148_)
);

OAI21X1 _12031_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5148_),
    .B(_5145_),
    .C(_5081_),
    .Y(_5149_)
);

AOI21X1 _12032_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5060_),
    .B(_5059_),
    .C(_4991_),
    .Y(_5150_)
);

OAI21X1 _12033_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4917_),
    .B(_5150_),
    .C(_5064_),
    .Y(_5151_)
);

NAND3X1 _12034_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5082_),
    .B(_5146_),
    .C(_5147_),
    .Y(_5152_)
);

NAND3X1 _12035_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5083_),
    .B(_5144_),
    .C(_5139_),
    .Y(_5153_)
);

NAND3X1 _12036_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5151_),
    .B(_5152_),
    .C(_5153_),
    .Y(_5154_)
);

NAND2X1 _12037_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5154_),
    .B(_5149_),
    .Y(_5155_)
);

NAND2X1 _12038_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5155_),
    .B(_5079_),
    .Y(_5156_)
);

OAI21X1 _12039_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4984_),
    .B(_5074_),
    .C(_5070_),
    .Y(_5157_)
);

AOI21X1 _12040_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5071_),
    .B(_4986_),
    .C(_5157_),
    .Y(_5158_)
);

AND2X2 _12041_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5149_),
    .B(_5154_),
    .Y(_5159_)
);

NAND2X1 _12042_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5159_),
    .B(_5158_),
    .Y(_5160_)
);

NAND2X1 _12043_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5156_),
    .B(_5160_),
    .Y(_5578_[8])
);

INVX1 _12044_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5154_),
    .Y(_5161_)
);

AOI21X1 _12045_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5079_),
    .B(_5149_),
    .C(_5161_),
    .Y(_5162_)
);

AOI21X1 _12046_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5143_),
    .B(_5142_),
    .C(_5085_),
    .Y(_5163_)
);

OAI21X1 _12047_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5083_),
    .B(_5163_),
    .C(_5146_),
    .Y(_5164_)
);

OAI21X1 _12048_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5086_),
    .B(_5090_),
    .C(_5095_),
    .Y(_5165_)
);

AOI21X1 _12049_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5131_),
    .B(_5132_),
    .C(_5099_),
    .Y(_5166_)
);

OAI21X1 _12050_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5097_),
    .B(_5166_),
    .C(_5136_),
    .Y(_5167_)
);

NAND2X1 _12051_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [2]),
    .B(gnd),
    .Y(_5168_)
);

NOR2X1 _12052_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5100_),
    .B(_5103_),
    .Y(_5169_)
);

NAND2X1 _12053_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_5169_),
    .Y(_5170_)
);

INVX1 _12054_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5170_),
    .Y(_5171_)
);

AOI21X1 _12055_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [3]),
    .B(gnd),
    .C(_5169_),
    .Y(_5172_)
);

OAI21X1 _12056_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5172_),
    .B(_5171_),
    .C(_5168_),
    .Y(_5173_)
);

INVX1 _12057_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5168_),
    .Y(_5174_)
);

INVX1 _12058_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5172_),
    .Y(_5175_)
);

NAND3X1 _12059_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5174_),
    .B(_5170_),
    .C(_5175_),
    .Y(_5176_)
);

AND2X2 _12060_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5176_),
    .B(_5173_),
    .Y(_5177_)
);

AOI21X1 _12061_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5121_),
    .B(_5120_),
    .C(_5105_),
    .Y(_5178_)
);

OAI21X1 _12062_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5104_),
    .B(_5178_),
    .C(_5125_),
    .Y(_5179_)
);

NOR2X1 _12063_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4914_),
    .B(_5103_),
    .Y(_5180_)
);

AND2X2 _12064_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4914_),
    .B(_5103_),
    .Y(_5181_)
);

NOR2X1 _12065_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5180_),
    .B(_5181_),
    .Y(_5182_)
);

NAND2X1 _12066_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [6]),
    .Y(_5183_)
);

AOI22X1 _12067_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7]_5_bF$buf3 ),
    .C(vdd),
    .D(\X[7] [6]),
    .Y(_5184_)
);

OAI22X1 _12068_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5036_),
    .B(_5183_),
    .C(_5106_),
    .D(_5184_),
    .Y(_5185_)
);

AOI22X1 _12069_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [6]),
    .C(vdd),
    .D(\X[7] [7]),
    .Y(_5186_)
);

AND2X2 _12070_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [7]),
    .Y(_5187_)
);

AOI21X1 _12071_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5113_),
    .B(_5187_),
    .C(_5186_),
    .Y(_5188_)
);

NAND2X1 _12072_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5188_),
    .B(_5185_),
    .Y(_5189_)
);

AND2X2 _12073_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [6]),
    .Y(_5190_)
);

AOI22X1 _12074_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5024_),
    .B(_5190_),
    .C(_5116_),
    .D(_5112_),
    .Y(_5191_)
);

NAND2X1 _12075_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[7] [7]),
    .Y(_5192_)
);

NAND2X1 _12076_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5183_),
    .B(_5192_),
    .Y(_5193_)
);

NAND2X1 _12077_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [7]),
    .Y(_5194_)
);

OAI21X1 _12078_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5115_),
    .B(_5194_),
    .C(_5193_),
    .Y(_5195_)
);

NAND2X1 _12079_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5195_),
    .B(_5191_),
    .Y(_5196_)
);

NAND3X1 _12080_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5182_),
    .B(_5189_),
    .C(_5196_),
    .Y(_5197_)
);

NAND2X1 _12081_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7]_5_bF$buf2 ),
    .B(gnd),
    .Y(_5198_)
);

INVX1 _12082_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [4]),
    .Y(_5199_)
);

OAI21X1 _12083_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5199_),
    .B(_5101_),
    .C(_4914_),
    .Y(_5200_)
);

OAI21X1 _12084_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4807_),
    .B(_5198_),
    .C(_5200_),
    .Y(_5201_)
);

NAND2X1 _12085_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5185_),
    .B(_5195_),
    .Y(_5202_)
);

NAND2X1 _12086_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5188_),
    .B(_5191_),
    .Y(_5203_)
);

NAND3X1 _12087_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5201_),
    .B(_5202_),
    .C(_5203_),
    .Y(_5204_)
);

NAND3X1 _12088_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5197_),
    .B(_5204_),
    .C(_5179_),
    .Y(_5205_)
);

NAND2X1 _12089_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5197_),
    .B(_5204_),
    .Y(_5206_)
);

NAND3X1 _12090_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5125_),
    .B(_5131_),
    .C(_5206_),
    .Y(_5207_)
);

NAND3X1 _12091_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5177_),
    .B(_5205_),
    .C(_5207_),
    .Y(_5208_)
);

NAND2X1 _12092_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5173_),
    .B(_5176_),
    .Y(_5209_)
);

AOI21X1 _12093_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5125_),
    .B(_5131_),
    .C(_5206_),
    .Y(_5210_)
);

AOI21X1 _12094_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5197_),
    .B(_5204_),
    .C(_5179_),
    .Y(_5211_)
);

OAI21X1 _12095_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5211_),
    .B(_5210_),
    .C(_5209_),
    .Y(_5212_)
);

NAND3X1 _12096_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5208_),
    .B(_5212_),
    .C(_5167_),
    .Y(_5213_)
);

INVX1 _12097_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5136_),
    .Y(_5214_)
);

AOI21X1 _12098_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5135_),
    .B(_5137_),
    .C(_5214_),
    .Y(_5215_)
);

INVX1 _12099_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5208_),
    .Y(_5216_)
);

AOI21X1 _12100_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5207_),
    .B(_5205_),
    .C(_5177_),
    .Y(_5217_)
);

OAI21X1 _12101_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5217_),
    .B(_5216_),
    .C(_5215_),
    .Y(_5218_)
);

NAND3X1 _12102_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5165_),
    .B(_5213_),
    .C(_5218_),
    .Y(_5219_)
);

INVX1 _12103_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5165_),
    .Y(_5220_)
);

INVX1 _12104_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5213_),
    .Y(_5221_)
);

AOI21X1 _12105_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5212_),
    .B(_5208_),
    .C(_5167_),
    .Y(_5222_)
);

OAI21X1 _12106_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5222_),
    .B(_5221_),
    .C(_5220_),
    .Y(_5223_)
);

NAND3X1 _12107_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5164_),
    .B(_5219_),
    .C(_5223_),
    .Y(_5224_)
);

INVX1 _12108_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5146_),
    .Y(_5225_)
);

AOI21X1 _12109_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5082_),
    .B(_5147_),
    .C(_5225_),
    .Y(_5226_)
);

OAI21X1 _12110_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5217_),
    .B(_5216_),
    .C(_5167_),
    .Y(_5227_)
);

NAND3X1 _12111_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5208_),
    .B(_5212_),
    .C(_5215_),
    .Y(_5228_)
);

AOI21X1 _12112_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5228_),
    .B(_5227_),
    .C(_5220_),
    .Y(_5229_)
);

AOI21X1 _12113_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5218_),
    .B(_5213_),
    .C(_5165_),
    .Y(_5230_)
);

OAI21X1 _12114_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5229_),
    .B(_5230_),
    .C(_5226_),
    .Y(_5231_)
);

AND2X2 _12115_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5231_),
    .B(_5224_),
    .Y(_5232_)
);

OR2X2 _12116_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5162_),
    .B(_5232_),
    .Y(_5233_)
);

NAND2X1 _12117_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5232_),
    .B(_5162_),
    .Y(_5234_)
);

NAND2X1 _12118_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5234_),
    .B(_5233_),
    .Y(_5578_[9])
);

NAND2X1 _12119_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5224_),
    .B(_5231_),
    .Y(_5235_)
);

NOR2X1 _12120_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5155_),
    .B(_5235_),
    .Y(_5236_)
);

NAND2X1 _12121_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5236_),
    .B(_5079_),
    .Y(_5237_)
);

AOI21X1 _12122_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5223_),
    .B(_5219_),
    .C(_5164_),
    .Y(_5238_)
);

AOI21X1 _12123_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5154_),
    .B(_5224_),
    .C(_5238_),
    .Y(_5239_)
);

INVX1 _12124_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5239_),
    .Y(_5240_)
);

OAI21X1 _12125_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5220_),
    .B(_5222_),
    .C(_5213_),
    .Y(_5241_)
);

OAI21X1 _12126_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5168_),
    .B(_5172_),
    .C(_5170_),
    .Y(_5242_)
);

OAI21X1 _12127_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5209_),
    .B(_5211_),
    .C(_5205_),
    .Y(_5243_)
);

INVX2 _12128_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_5244_)
);

NOR3X1 _12129_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5087_),
    .B(_4914_),
    .C(_5103_),
    .Y(_5245_)
);

OAI22X1 _12130_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5199_),
    .B(_5087_),
    .C(_4807_),
    .D(_5198_),
    .Y(_5246_)
);

INVX1 _12131_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5246_),
    .Y(_5247_)
);

OAI22X1 _12132_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4797_),
    .B(_5244_),
    .C(_5245_),
    .D(_5247_),
    .Y(_5248_)
);

NOR2X1 _12133_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4797_),
    .B(_5244_),
    .Y(_5249_)
);

NAND2X1 _12134_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_5180_),
    .Y(_5250_)
);

NAND3X1 _12135_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5249_),
    .B(_5246_),
    .C(_5250_),
    .Y(_5251_)
);

AND2X2 _12136_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5248_),
    .B(_5251_),
    .Y(_5252_)
);

NOR2X1 _12137_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5188_),
    .B(_5185_),
    .Y(_5253_)
);

OAI21X1 _12138_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5201_),
    .B(_5253_),
    .C(_5189_),
    .Y(_5254_)
);

NAND2X1 _12139_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [6]),
    .Y(_5255_)
);

NOR2X1 _12140_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5255_),
    .B(_5198_),
    .Y(_5256_)
);

AND2X2 _12141_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5255_),
    .B(_5198_),
    .Y(_5257_)
);

OAI22X1 _12142_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5113_),
    .B(_5194_),
    .C(_5256_),
    .D(_5257_),
    .Y(_5258_)
);

AND2X2 _12143_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [6]),
    .Y(_5259_)
);

AND2X2 _12144_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7]_5_bF$buf1 ),
    .B(gnd),
    .Y(_5260_)
);

NAND2X1 _12145_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5259_),
    .B(_5260_),
    .Y(_5261_)
);

OAI21X1 _12146_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4856_),
    .B(_5101_),
    .C(_5255_),
    .Y(_5262_)
);

AOI21X1 _12147_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[7] [6]),
    .C(_5194_),
    .Y(_5263_)
);

NAND3X1 _12148_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5262_),
    .B(_5263_),
    .C(_5261_),
    .Y(_5264_)
);

AND2X2 _12149_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5258_),
    .B(_5264_),
    .Y(_5265_)
);

NAND2X1 _12150_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5265_),
    .B(_5254_),
    .Y(_5266_)
);

NAND2X1 _12151_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5264_),
    .B(_5258_),
    .Y(_5267_)
);

NAND3X1 _12152_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5189_),
    .B(_5267_),
    .C(_5197_),
    .Y(_5268_)
);

NAND3X1 _12153_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5252_),
    .B(_5268_),
    .C(_5266_),
    .Y(_5269_)
);

NAND2X1 _12154_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5251_),
    .B(_5248_),
    .Y(_5270_)
);

NAND2X1 _12155_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5267_),
    .B(_5254_),
    .Y(_5271_)
);

NAND3X1 _12156_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5189_),
    .B(_5265_),
    .C(_5197_),
    .Y(_5272_)
);

NAND3X1 _12157_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5270_),
    .B(_5272_),
    .C(_5271_),
    .Y(_5273_)
);

NAND3X1 _12158_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5269_),
    .B(_5273_),
    .C(_5243_),
    .Y(_5274_)
);

NAND2X1 _12159_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5273_),
    .B(_5269_),
    .Y(_5275_)
);

NAND3X1 _12160_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5205_),
    .B(_5208_),
    .C(_5275_),
    .Y(_5276_)
);

NAND3X1 _12161_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5242_),
    .B(_5276_),
    .C(_5274_),
    .Y(_5277_)
);

INVX1 _12162_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5242_),
    .Y(_5278_)
);

NAND2X1 _12163_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5275_),
    .B(_5243_),
    .Y(_5279_)
);

AOI21X1 _12164_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5177_),
    .B(_5207_),
    .C(_5210_),
    .Y(_5280_)
);

AND2X2 _12165_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5269_),
    .B(_5273_),
    .Y(_5281_)
);

NAND2X1 _12166_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5280_),
    .B(_5281_),
    .Y(_5282_)
);

NAND3X1 _12167_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5278_),
    .B(_5279_),
    .C(_5282_),
    .Y(_5283_)
);

AOI21X1 _12168_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5277_),
    .B(_5283_),
    .C(_5241_),
    .Y(_5284_)
);

NAND2X1 _12169_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5277_),
    .B(_5283_),
    .Y(_5285_)
);

AOI21X1 _12170_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5213_),
    .B(_5219_),
    .C(_5285_),
    .Y(_5286_)
);

NOR2X1 _12171_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5284_),
    .B(_5286_),
    .Y(_5287_)
);

INVX1 _12172_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5287_),
    .Y(_5288_)
);

AOI21X1 _12173_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5237_),
    .B(_5240_),
    .C(_5288_),
    .Y(_5289_)
);

NAND2X1 _12174_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5159_),
    .B(_5232_),
    .Y(_5290_)
);

OAI21X1 _12175_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5290_),
    .B(_5158_),
    .C(_5240_),
    .Y(_5291_)
);

NOR2X1 _12176_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5287_),
    .B(_5291_),
    .Y(_5292_)
);

NOR2X1 _12177_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5289_),
    .B(_5292_),
    .Y(_5578_[10])
);

NAND3X1 _12178_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5277_),
    .B(_5283_),
    .C(_5241_),
    .Y(_5293_)
);

NAND2X1 _12179_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5287_),
    .B(_5291_),
    .Y(_5294_)
);

NOR2X1 _12180_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5275_),
    .B(_5280_),
    .Y(_5295_)
);

AOI21X1 _12181_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5242_),
    .B(_5276_),
    .C(_5295_),
    .Y(_5296_)
);

NAND2X1 _12182_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5250_),
    .B(_5251_),
    .Y(_5297_)
);

NAND2X1 _12183_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5266_),
    .B(_5269_),
    .Y(_5298_)
);

NOR3X1 _12184_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5087_),
    .B(_5255_),
    .C(_5198_),
    .Y(_5299_)
);

AOI22X1 _12185_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7]_5_bF$buf0 ),
    .B(gnd),
    .C(_5259_),
    .D(_5260_),
    .Y(_5300_)
);

OAI22X1 _12186_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5199_),
    .B(_5244_),
    .C(_5300_),
    .D(_5299_),
    .Y(_5301_)
);

NOR2X1 _12187_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5199_),
    .B(_5244_),
    .Y(_5302_)
);

NAND2X1 _12188_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_5256_),
    .Y(_5303_)
);

OAI21X1 _12189_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4856_),
    .B(_5087_),
    .C(_5261_),
    .Y(_5304_)
);

NAND3X1 _12190_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5302_),
    .B(_5303_),
    .C(_5304_),
    .Y(_5305_)
);

NAND2X1 _12191_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5301_),
    .B(_5305_),
    .Y(_5306_)
);

NAND2X1 _12192_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5113_),
    .B(_5187_),
    .Y(_5307_)
);

NAND2X1 _12193_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[7] [7]),
    .Y(_5308_)
);

OAI22X1 _12194_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5015_),
    .B(_5017_),
    .C(_5101_),
    .D(_4926_),
    .Y(_5309_)
);

OAI21X1 _12195_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5255_),
    .B(_5308_),
    .C(_5309_),
    .Y(_5310_)
);

NAND3X1 _12196_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5307_),
    .B(_5310_),
    .C(_5264_),
    .Y(_5311_)
);

INVX1 _12197_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5311_),
    .Y(_5312_)
);

AOI21X1 _12198_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5264_),
    .B(_5307_),
    .C(_5310_),
    .Y(_5313_)
);

OAI21X1 _12199_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5313_),
    .B(_5312_),
    .C(_5306_),
    .Y(_5314_)
);

AND2X2 _12200_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5305_),
    .B(_5301_),
    .Y(_5315_)
);

INVX1 _12201_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5313_),
    .Y(_5316_)
);

NAND3X1 _12202_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5311_),
    .B(_5316_),
    .C(_5315_),
    .Y(_5317_)
);

AND2X2 _12203_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5317_),
    .B(_5314_),
    .Y(_5318_)
);

NAND2X1 _12204_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5318_),
    .B(_5298_),
    .Y(_5319_)
);

AOI21X1 _12205_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5197_),
    .B(_5189_),
    .C(_5267_),
    .Y(_5320_)
);

AOI21X1 _12206_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5252_),
    .B(_5268_),
    .C(_5320_),
    .Y(_5321_)
);

NAND2X1 _12207_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5314_),
    .B(_5317_),
    .Y(_5322_)
);

NAND2X1 _12208_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5322_),
    .B(_5321_),
    .Y(_5323_)
);

NAND3X1 _12209_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5297_),
    .B(_5323_),
    .C(_5319_),
    .Y(_5324_)
);

INVX1 _12210_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5297_),
    .Y(_5325_)
);

NAND2X1 _12211_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5322_),
    .B(_5298_),
    .Y(_5326_)
);

NAND2X1 _12212_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5321_),
    .B(_5318_),
    .Y(_5327_)
);

NAND3X1 _12213_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5325_),
    .B(_5327_),
    .C(_5326_),
    .Y(_5328_)
);

NAND2X1 _12214_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5324_),
    .B(_5328_),
    .Y(_5329_)
);

NAND2X1 _12215_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5329_),
    .B(_5296_),
    .Y(_5330_)
);

AOI21X1 _12216_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5269_),
    .B(_5273_),
    .C(_5243_),
    .Y(_5331_)
);

OAI21X1 _12217_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5278_),
    .B(_5331_),
    .C(_5274_),
    .Y(_5332_)
);

NAND3X1 _12218_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5324_),
    .B(_5328_),
    .C(_5332_),
    .Y(_5333_)
);

NAND2X1 _12219_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5330_),
    .B(_5333_),
    .Y(_5334_)
);

INVX1 _12220_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5334_),
    .Y(_5335_)
);

NAND3X1 _12221_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5293_),
    .B(_5335_),
    .C(_5294_),
    .Y(_5336_)
);

OAI21X1 _12222_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5286_),
    .B(_5289_),
    .C(_5334_),
    .Y(_5337_)
);

NAND2X1 _12223_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5336_),
    .B(_5337_),
    .Y(_5578_[11])
);

NOR3X1 _12224_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5284_),
    .B(_5286_),
    .C(_5334_),
    .Y(_5338_)
);

NAND3X1 _12225_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5236_),
    .B(_5338_),
    .C(_5079_),
    .Y(_5339_)
);

OAI21X1 _12226_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5293_),
    .B(_5334_),
    .C(_5333_),
    .Y(_5340_)
);

AOI21X1 _12227_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5338_),
    .B(_5239_),
    .C(_5340_),
    .Y(_5341_)
);

AND2X2 _12228_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5324_),
    .B(_5319_),
    .Y(_5342_)
);

OAI21X1 _12229_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5087_),
    .B(_5261_),
    .C(_5305_),
    .Y(_5343_)
);

OAI21X1 _12230_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5312_),
    .B(_5306_),
    .C(_5316_),
    .Y(_5344_)
);

INVX1 _12231_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5344_),
    .Y(_5345_)
);

INVX1 _12232_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5308_),
    .Y(_5346_)
);

NOR2X1 _12233_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4856_),
    .B(_5244_),
    .Y(_5347_)
);

NOR2X1 _12234_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5255_),
    .B(_5308_),
    .Y(_5348_)
);

NOR2X1 _12235_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4926_),
    .B(_5087_),
    .Y(_5349_)
);

NOR2X1 _12236_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5349_),
    .B(_5348_),
    .Y(_5350_)
);

AOI21X1 _12237_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_5348_),
    .C(_5350_),
    .Y(_5351_)
);

OR2X2 _12238_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5351_),
    .B(_5347_),
    .Y(_5352_)
);

NAND2X1 _12239_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5347_),
    .B(_5351_),
    .Y(_5353_)
);

NAND3X1 _12240_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5346_),
    .B(_5353_),
    .C(_5352_),
    .Y(_5354_)
);

NOR2X1 _12241_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5347_),
    .B(_5351_),
    .Y(_5355_)
);

INVX1 _12242_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5353_),
    .Y(_5356_)
);

OAI21X1 _12243_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5355_),
    .B(_5356_),
    .C(_5308_),
    .Y(_5357_)
);

NAND2X1 _12244_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5354_),
    .B(_5357_),
    .Y(_5358_)
);

NAND2X1 _12245_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5345_),
    .B(_5358_),
    .Y(_5359_)
);

NAND3X1 _12246_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5344_),
    .B(_5354_),
    .C(_5357_),
    .Y(_5360_)
);

AOI21X1 _12247_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5359_),
    .B(_5360_),
    .C(_5343_),
    .Y(_5361_)
);

NAND3X1 _12248_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5343_),
    .B(_5360_),
    .C(_5359_),
    .Y(_5362_)
);

INVX1 _12249_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5362_),
    .Y(_5363_)
);

OAI21X1 _12250_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5361_),
    .B(_5363_),
    .C(_5342_),
    .Y(_5364_)
);

OR2X2 _12251_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5363_),
    .B(_5361_),
    .Y(_5365_)
);

OR2X2 _12252_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5365_),
    .B(_5342_),
    .Y(_5366_)
);

NAND2X1 _12253_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5364_),
    .B(_5366_),
    .Y(_5367_)
);

AOI21X1 _12254_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5339_),
    .B(_5341_),
    .C(_5367_),
    .Y(_5368_)
);

NAND3X1 _12255_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5159_),
    .B(_5232_),
    .C(_5338_),
    .Y(_5369_)
);

OAI21X1 _12256_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5158_),
    .B(_5369_),
    .C(_5341_),
    .Y(_5370_)
);

INVX1 _12257_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5367_),
    .Y(_5371_)
);

NOR2X1 _12258_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5371_),
    .B(_5370_),
    .Y(_5372_)
);

NOR2X1 _12259_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5368_),
    .B(_5372_),
    .Y(_5578_[12])
);

NOR2X1 _12260_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5342_),
    .B(_5365_),
    .Y(_5373_)
);

INVX1 _12261_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5348_),
    .Y(_5374_)
);

OAI21X1 _12262_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5087_),
    .B(_5374_),
    .C(_5353_),
    .Y(_5375_)
);

INVX1 _12263_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5375_),
    .Y(_5376_)
);

NOR2X1 _12264_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5017_),
    .B(_5244_),
    .Y(_5377_)
);

NAND2X1 _12265_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5349_),
    .B(_5377_),
    .Y(_5378_)
);

OAI22X1 _12266_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4926_),
    .B(_5244_),
    .C(_5087_),
    .D(_5017_),
    .Y(_5379_)
);

NAND2X1 _12267_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5379_),
    .B(_5378_),
    .Y(_5380_)
);

NAND2X1 _12268_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5380_),
    .B(_5354_),
    .Y(_5381_)
);

OR2X2 _12269_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5354_),
    .B(_5380_),
    .Y(_5382_)
);

NAND2X1 _12270_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5381_),
    .B(_5382_),
    .Y(_5383_)
);

NAND2X1 _12271_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5376_),
    .B(_5383_),
    .Y(_5384_)
);

OR2X2 _12272_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5383_),
    .B(_5376_),
    .Y(_5385_)
);

NAND2X1 _12273_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5384_),
    .B(_5385_),
    .Y(_5386_)
);

NAND3X1 _12274_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5360_),
    .B(_5362_),
    .C(_5386_),
    .Y(_5387_)
);

OAI21X1 _12275_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5345_),
    .B(_5358_),
    .C(_5362_),
    .Y(_5388_)
);

AND2X2 _12276_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5385_),
    .B(_5384_),
    .Y(_5389_)
);

NAND2X1 _12277_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5388_),
    .B(_5389_),
    .Y(_5390_)
);

NAND2X1 _12278_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5387_),
    .B(_5390_),
    .Y(_5391_)
);

OAI21X1 _12279_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5373_),
    .B(_5368_),
    .C(_5391_),
    .Y(_5392_)
);

NAND2X1 _12280_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5371_),
    .B(_5370_),
    .Y(_5393_)
);

AND2X2 _12281_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5390_),
    .B(_5387_),
    .Y(_5394_)
);

NAND3X1 _12282_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5366_),
    .B(_5394_),
    .C(_5393_),
    .Y(_5395_)
);

NAND2X1 _12283_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5395_),
    .B(_5392_),
    .Y(_5578_[13])
);

NAND3X1 _12284_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5364_),
    .B(_5366_),
    .C(_5394_),
    .Y(_5396_)
);

AOI21X1 _12285_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5339_),
    .B(_5341_),
    .C(_5396_),
    .Y(_5397_)
);

OAI21X1 _12286_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5366_),
    .B(_5391_),
    .C(_5390_),
    .Y(_5398_)
);

OAI21X1 _12287_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5376_),
    .B(_5383_),
    .C(_5382_),
    .Y(_5399_)
);

AND2X2 _12288_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5378_),
    .B(_5377_),
    .Y(_5400_)
);

OR2X2 _12289_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5399_),
    .B(_5400_),
    .Y(_5401_)
);

NAND2X1 _12290_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5400_),
    .B(_5399_),
    .Y(_5402_)
);

NAND2X1 _12291_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5402_),
    .B(_5401_),
    .Y(_5403_)
);

OAI21X1 _12292_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5398_),
    .B(_5397_),
    .C(_5403_),
    .Y(_5404_)
);

INVX1 _12293_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5364_),
    .Y(_5405_)
);

NOR3X1 _12294_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5405_),
    .B(_5373_),
    .C(_5391_),
    .Y(_5406_)
);

NAND2X1 _12295_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5406_),
    .B(_5370_),
    .Y(_5407_)
);

INVX1 _12296_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5398_),
    .Y(_5408_)
);

INVX1 _12297_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5403_),
    .Y(_5409_)
);

NAND3X1 _12298_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5408_),
    .B(_5409_),
    .C(_5407_),
    .Y(_5410_)
);

NAND2X1 _12299_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5410_),
    .B(_5404_),
    .Y(_5578_[14])
);

OAI21X1 _12300_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5398_),
    .B(_5397_),
    .C(_5409_),
    .Y(_5411_)
);

OAI21X1 _12301_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5349_),
    .B(_5399_),
    .C(_5377_),
    .Y(_5412_)
);

NAND2X1 _12302_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5412_),
    .B(_5411_),
    .Y(_5578_[15])
);

INVX1 _12303_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4806_),
    .Y(_5573_[0])
);

AND2X2 _12304_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [0]),
    .B(\u_fir_pe6.mul [0]),
    .Y(_5413_)
);

INVX1 _12305_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [1]),
    .Y(_5414_)
);

INVX1 _12306_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.mul [1]),
    .Y(_5415_)
);

NOR2X1 _12307_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5414_),
    .B(_5415_),
    .Y(_5416_)
);

NOR2X1 _12308_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [1]),
    .B(\u_fir_pe6.mul [1]),
    .Y(_5417_)
);

NOR2X1 _12309_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5417_),
    .B(_5416_),
    .Y(_5418_)
);

NAND2X1 _12310_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5413_),
    .B(_5418_),
    .Y(_5419_)
);

INVX1 _12311_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5419_),
    .Y(_5420_)
);

NOR2X1 _12312_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5413_),
    .B(_5418_),
    .Y(_5421_)
);

NOR2X1 _12313_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5421_),
    .B(_5420_),
    .Y(_5572_[1])
);

OAI21X1 _12314_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5414_),
    .B(_5415_),
    .C(_5419_),
    .Y(_5422_)
);

AND2X2 _12315_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [2]),
    .B(\u_fir_pe6.mul [2]),
    .Y(_5423_)
);

NOR2X1 _12316_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [2]),
    .B(\u_fir_pe6.mul [2]),
    .Y(_5424_)
);

OAI21X1 _12317_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5423_),
    .B(_5424_),
    .C(_5422_),
    .Y(_5425_)
);

INVX1 _12318_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5422_),
    .Y(_5426_)
);

NOR2X1 _12319_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5424_),
    .B(_5423_),
    .Y(_5427_)
);

NAND2X1 _12320_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5427_),
    .B(_5426_),
    .Y(_5428_)
);

NAND2X1 _12321_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5425_),
    .B(_5428_),
    .Y(_5572_[2])
);

AOI21X1 _12322_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5422_),
    .B(_5427_),
    .C(_5423_),
    .Y(_5429_)
);

INVX1 _12323_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [3]),
    .Y(_5430_)
);

INVX1 _12324_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.mul [3]),
    .Y(_5431_)
);

NOR2X1 _12325_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5430_),
    .B(_5431_),
    .Y(_5432_)
);

NOR2X1 _12326_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [3]),
    .B(\u_fir_pe6.mul [3]),
    .Y(_5433_)
);

NOR2X1 _12327_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5433_),
    .B(_5432_),
    .Y(_5434_)
);

NAND2X1 _12328_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5434_),
    .B(_5429_),
    .Y(_5435_)
);

OR2X2 _12329_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5429_),
    .B(_5434_),
    .Y(_5436_)
);

NAND2X1 _12330_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5435_),
    .B(_5436_),
    .Y(_5572_[3])
);

INVX1 _12331_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [4]),
    .Y(_5437_)
);

INVX1 _12332_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.mul [4]),
    .Y(_5438_)
);

NOR2X1 _12333_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5437_),
    .B(_5438_),
    .Y(_5439_)
);

NOR2X1 _12334_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [4]),
    .B(\u_fir_pe6.mul [4]),
    .Y(_5440_)
);

NOR2X1 _12335_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5440_),
    .B(_5439_),
    .Y(_5441_)
);

INVX1 _12336_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5432_),
    .Y(_5442_)
);

OAI21X1 _12337_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5433_),
    .B(_5429_),
    .C(_5442_),
    .Y(_5443_)
);

NAND2X1 _12338_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5441_),
    .B(_5443_),
    .Y(_5444_)
);

OR2X2 _12339_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5443_),
    .B(_5441_),
    .Y(_5445_)
);

AND2X2 _12340_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5445_),
    .B(_5444_),
    .Y(_5572_[4])
);

OAI21X1 _12341_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5437_),
    .B(_5438_),
    .C(_5444_),
    .Y(_5446_)
);

INVX1 _12342_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [5]),
    .Y(_5447_)
);

INVX1 _12343_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.mul [5]),
    .Y(_5448_)
);

NOR2X1 _12344_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5447_),
    .B(_5448_),
    .Y(_5449_)
);

NOR2X1 _12345_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [5]),
    .B(\u_fir_pe6.mul [5]),
    .Y(_5450_)
);

NOR2X1 _12346_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5450_),
    .B(_5449_),
    .Y(_5451_)
);

NAND2X1 _12347_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5451_),
    .B(_5446_),
    .Y(_5452_)
);

OR2X2 _12348_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5446_),
    .B(_5451_),
    .Y(_5453_)
);

AND2X2 _12349_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5453_),
    .B(_5452_),
    .Y(_5572_[5])
);

OAI21X1 _12350_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5447_),
    .B(_5448_),
    .C(_5452_),
    .Y(_5454_)
);

INVX1 _12351_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [6]),
    .Y(_5455_)
);

INVX1 _12352_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.mul [6]),
    .Y(_5456_)
);

NOR2X1 _12353_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5455_),
    .B(_5456_),
    .Y(_5457_)
);

NOR2X1 _12354_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [6]),
    .B(\u_fir_pe6.mul [6]),
    .Y(_5458_)
);

NOR2X1 _12355_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5458_),
    .B(_5457_),
    .Y(_5459_)
);

NAND2X1 _12356_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5459_),
    .B(_5454_),
    .Y(_5460_)
);

OR2X2 _12357_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5454_),
    .B(_5459_),
    .Y(_5461_)
);

AND2X2 _12358_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5461_),
    .B(_5460_),
    .Y(_5572_[6])
);

OAI21X1 _12359_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5455_),
    .B(_5456_),
    .C(_5460_),
    .Y(_5462_)
);

INVX1 _12360_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [7]),
    .Y(_5463_)
);

INVX1 _12361_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.mul [7]),
    .Y(_5464_)
);

NOR2X1 _12362_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5463_),
    .B(_5464_),
    .Y(_5465_)
);

NOR2X1 _12363_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [7]),
    .B(\u_fir_pe6.mul [7]),
    .Y(_5466_)
);

OAI21X1 _12364_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5465_),
    .B(_5466_),
    .C(_5462_),
    .Y(_5467_)
);

INVX1 _12365_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5462_),
    .Y(_5468_)
);

NOR2X1 _12366_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5466_),
    .B(_5465_),
    .Y(_5469_)
);

NAND2X1 _12367_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5469_),
    .B(_5468_),
    .Y(_5470_)
);

NAND2X1 _12368_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5467_),
    .B(_5470_),
    .Y(_5572_[7])
);

INVX1 _12369_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [8]),
    .Y(_5472_)
);

INVX1 _12370_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.mul [8]),
    .Y(_5473_)
);

NOR2X1 _12371_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5472_),
    .B(_5473_),
    .Y(_5474_)
);

NOR2X1 _12372_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [8]),
    .B(\u_fir_pe6.mul [8]),
    .Y(_5475_)
);

NAND2X1 _12373_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5439_),
    .B(_5451_),
    .Y(_5476_)
);

OAI21X1 _12374_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5447_),
    .B(_5448_),
    .C(_5476_),
    .Y(_5477_)
);

NAND2X1 _12375_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5457_),
    .B(_5469_),
    .Y(_5478_)
);

OAI21X1 _12376_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5463_),
    .B(_5464_),
    .C(_5478_),
    .Y(_5479_)
);

AND2X2 _12377_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5459_),
    .B(_5469_),
    .Y(_5480_)
);

AOI21X1 _12378_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5477_),
    .B(_5480_),
    .C(_5479_),
    .Y(_5481_)
);

AND2X2 _12379_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5441_),
    .B(_5451_),
    .Y(_5483_)
);

NAND3X1 _12380_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5483_),
    .B(_5480_),
    .C(_5443_),
    .Y(_5484_)
);

NAND2X1 _12381_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5481_),
    .B(_5484_),
    .Y(_5485_)
);

OAI21X1 _12382_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5474_),
    .B(_5475_),
    .C(_5485_),
    .Y(_5486_)
);

NOR2X1 _12383_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5475_),
    .B(_5474_),
    .Y(_5487_)
);

INVX1 _12384_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5485_),
    .Y(_5488_)
);

NAND2X1 _12385_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5487_),
    .B(_5488_),
    .Y(_5489_)
);

NAND2X1 _12386_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5486_),
    .B(_5489_),
    .Y(_5572_[8])
);

INVX1 _12387_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5474_),
    .Y(_5490_)
);

INVX1 _12388_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5487_),
    .Y(_5491_)
);

OAI21X1 _12389_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5491_),
    .B(_5488_),
    .C(_5490_),
    .Y(_5493_)
);

AND2X2 _12390_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [9]),
    .B(\u_fir_pe6.mul [9]),
    .Y(_5494_)
);

NOR2X1 _12391_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [9]),
    .B(\u_fir_pe6.mul [9]),
    .Y(_5495_)
);

NOR2X1 _12392_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5495_),
    .B(_5494_),
    .Y(_5496_)
);

INVX1 _12393_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5496_),
    .Y(_5497_)
);

OR2X2 _12394_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5493_),
    .B(_5497_),
    .Y(_5498_)
);

OAI21X1 _12395_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5494_),
    .B(_5495_),
    .C(_5493_),
    .Y(_5499_)
);

NAND2X1 _12396_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5499_),
    .B(_5498_),
    .Y(_5572_[9])
);

NOR2X1 _12397_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5497_),
    .B(_5491_),
    .Y(_5500_)
);

AOI21X1 _12398_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5496_),
    .B(_5474_),
    .C(_5494_),
    .Y(_5501_)
);

INVX1 _12399_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5501_),
    .Y(_5503_)
);

AOI21X1 _12400_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5485_),
    .B(_5500_),
    .C(_5503_),
    .Y(_5504_)
);

INVX1 _12401_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5504_),
    .Y(_5505_)
);

INVX1 _12402_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [10]),
    .Y(_5506_)
);

INVX1 _12403_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.mul [10]),
    .Y(_5507_)
);

NOR2X1 _12404_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5506_),
    .B(_5507_),
    .Y(_5508_)
);

NOR2X1 _12405_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [10]),
    .B(\u_fir_pe6.mul [10]),
    .Y(_5509_)
);

NOR2X1 _12406_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5509_),
    .B(_5508_),
    .Y(_5510_)
);

NAND2X1 _12407_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5510_),
    .B(_5505_),
    .Y(_5511_)
);

OAI21X1 _12408_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5508_),
    .B(_5509_),
    .C(_5504_),
    .Y(_5512_)
);

AND2X2 _12409_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5511_),
    .B(_5512_),
    .Y(_5572_[10])
);

OAI21X1 _12410_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5506_),
    .B(_5507_),
    .C(_5511_),
    .Y(_5514_)
);

AND2X2 _12411_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [11]),
    .B(\u_fir_pe6.mul [11]),
    .Y(_5515_)
);

NOR2X1 _12412_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [11]),
    .B(\u_fir_pe6.mul [11]),
    .Y(_5516_)
);

NOR2X1 _12413_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5516_),
    .B(_5515_),
    .Y(_5517_)
);

NOR2X1 _12414_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5517_),
    .B(_5514_),
    .Y(_5518_)
);

AND2X2 _12415_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5514_),
    .B(_5517_),
    .Y(_5519_)
);

NOR2X1 _12416_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5518_),
    .B(_5519_),
    .Y(_5572_[11])
);

AOI21X1 _12417_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5517_),
    .B(_5508_),
    .C(_5515_),
    .Y(_5520_)
);

NAND2X1 _12418_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5517_),
    .B(_5510_),
    .Y(_5521_)
);

OAI21X1 _12419_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5521_),
    .B(_5504_),
    .C(_5520_),
    .Y(_5523_)
);

INVX1 _12420_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [12]),
    .Y(_5524_)
);

INVX1 _12421_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.mul [12]),
    .Y(_5525_)
);

NOR2X1 _12422_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5524_),
    .B(_5525_),
    .Y(_5526_)
);

NOR2X1 _12423_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [12]),
    .B(\u_fir_pe6.mul [12]),
    .Y(_5527_)
);

NOR2X1 _12424_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5527_),
    .B(_5526_),
    .Y(_5528_)
);

NAND2X1 _12425_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5528_),
    .B(_5523_),
    .Y(_5529_)
);

OR2X2 _12426_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5523_),
    .B(_5528_),
    .Y(_5530_)
);

AND2X2 _12427_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5530_),
    .B(_5529_),
    .Y(_5572_[12])
);

OAI21X1 _12428_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5524_),
    .B(_5525_),
    .C(_5529_),
    .Y(_5531_)
);

INVX1 _12429_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [13]),
    .Y(_5533_)
);

INVX1 _12430_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.mul [13]),
    .Y(_5534_)
);

NOR2X1 _12431_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5533_),
    .B(_5534_),
    .Y(_5535_)
);

NOR2X1 _12432_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [13]),
    .B(\u_fir_pe6.mul [13]),
    .Y(_5536_)
);

NOR2X1 _12433_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5536_),
    .B(_5535_),
    .Y(_5537_)
);

NAND2X1 _12434_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5537_),
    .B(_5531_),
    .Y(_5538_)
);

OR2X2 _12435_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5531_),
    .B(_5537_),
    .Y(_5539_)
);

AND2X2 _12436_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5539_),
    .B(_5538_),
    .Y(_5572_[13])
);

OAI21X1 _12437_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5533_),
    .B(_5534_),
    .C(_5538_),
    .Y(_5540_)
);

INVX1 _12438_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [14]),
    .Y(_5541_)
);

INVX1 _12439_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.mul [14]),
    .Y(_5543_)
);

NOR2X1 _12440_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5541_),
    .B(_5543_),
    .Y(_5544_)
);

NOR2X1 _12441_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [14]),
    .B(\u_fir_pe6.mul [14]),
    .Y(_5545_)
);

NOR2X1 _12442_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5545_),
    .B(_5544_),
    .Y(_5546_)
);

AND2X2 _12443_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5540_),
    .B(_5546_),
    .Y(_5547_)
);

NOR2X1 _12444_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5546_),
    .B(_5540_),
    .Y(_5548_)
);

NOR2X1 _12445_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5548_),
    .B(_5547_),
    .Y(_5572_[14])
);

INVX1 _12446_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5544_),
    .Y(_5549_)
);

NAND2X1 _12447_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5546_),
    .B(_5540_),
    .Y(_5550_)
);

NAND2X1 _12448_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [15]),
    .B(\u_fir_pe6.mul [15]),
    .Y(_5551_)
);

OR2X2 _12449_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [15]),
    .B(\u_fir_pe6.mul [15]),
    .Y(_5553_)
);

NAND2X1 _12450_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5551_),
    .B(_5553_),
    .Y(_5554_)
);

INVX1 _12451_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5554_),
    .Y(_5555_)
);

NAND3X1 _12452_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5549_),
    .B(_5555_),
    .C(_5550_),
    .Y(_5556_)
);

OAI21X1 _12453_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5544_),
    .B(_5547_),
    .C(_5554_),
    .Y(_5557_)
);

NAND2X1 _12454_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5556_),
    .B(_5557_),
    .Y(_5572_[15])
);

NOR2X1 _12455_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe6.rYin [0]),
    .B(\u_fir_pe6.mul [0]),
    .Y(_5558_)
);

NOR2X1 _12456_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5558_),
    .B(_5413_),
    .Y(_5571_[0])
);

AOI21X1 _12457_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[7] [0]),
    .B(gnd),
    .C(_5482_),
    .Y(_5559_)
);

NOR2X1 _12458_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5559_),
    .B(_5502_),
    .Y(_5574_[1])
);

NOR2X1 _12459_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5502_),
    .B(_5566_),
    .Y(_5561_)
);

NOR2X1 _12460_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5561_),
    .B(_5568_),
    .Y(_5575_[2])
);

DFFPOSX1 _12461_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_5571_[0]),
    .Q(_6377_[0])
);

DFFPOSX1 _12462_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_5572_[1]),
    .Q(_6377_[1])
);

DFFPOSX1 _12463_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_5572_[2]),
    .Q(_6377_[2])
);

DFFPOSX1 _12464_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_5572_[3]),
    .Q(_6377_[3])
);

DFFPOSX1 _12465_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf57),
    .D(_5572_[4]),
    .Q(_6377_[4])
);

DFFPOSX1 _12466_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf56),
    .D(_5572_[5]),
    .Q(_6377_[5])
);

DFFPOSX1 _12467_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf55),
    .D(_5572_[6]),
    .Q(_6377_[6])
);

DFFPOSX1 _12468_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf54),
    .D(_5572_[7]),
    .Q(_6377_[7])
);

DFFPOSX1 _12469_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf53),
    .D(_5572_[8]),
    .Q(_6377_[8])
);

DFFPOSX1 _12470_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf52),
    .D(_5572_[9]),
    .Q(_6377_[9])
);

DFFPOSX1 _12471_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf51),
    .D(_5572_[10]),
    .Q(_6377_[10])
);

DFFPOSX1 _12472_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf50),
    .D(_5572_[11]),
    .Q(_6377_[11])
);

DFFPOSX1 _12473_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf49),
    .D(_5572_[12]),
    .Q(_6377_[12])
);

DFFPOSX1 _12474_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf48),
    .D(_5572_[13]),
    .Q(_6377_[13])
);

DFFPOSX1 _12475_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf47),
    .D(_5572_[14]),
    .Q(_6377_[14])
);

DFFPOSX1 _12476_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf46),
    .D(_5572_[15]),
    .Q(_6377_[15])
);

DFFPOSX1 _12477_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf45),
    .D(\X[7] [0]),
    .Q(_6376_[0])
);

DFFPOSX1 _12478_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf44),
    .D(\X[7] [1]),
    .Q(_6376_[1])
);

DFFPOSX1 _12479_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf43),
    .D(\X[7] [2]),
    .Q(_6376_[2])
);

DFFPOSX1 _12480_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf42),
    .D(\X[7] [3]),
    .Q(_6376_[3])
);

DFFPOSX1 _12481_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf41),
    .D(\X[7] [4]),
    .Q(_6376_[4])
);

DFFPOSX1 _12482_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf40),
    .D(\X[7]_5_bF$buf3 ),
    .Q(_6376_[5])
);

DFFPOSX1 _12483_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf39),
    .D(\X[7] [6]),
    .Q(_6376_[6])
);

DFFPOSX1 _12484_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf38),
    .D(\X[7] [7]),
    .Q(_6376_[7])
);

DFFPOSX1 _12485_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf37),
    .D(\Y[7] [0]),
    .Q(\u_fir_pe6.rYin [0])
);

DFFPOSX1 _12486_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf36),
    .D(\Y[7] [1]),
    .Q(\u_fir_pe6.rYin [1])
);

DFFPOSX1 _12487_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf35),
    .D(\Y[7] [2]),
    .Q(\u_fir_pe6.rYin [2])
);

DFFPOSX1 _12488_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf34),
    .D(\Y[7] [3]),
    .Q(\u_fir_pe6.rYin [3])
);

DFFPOSX1 _12489_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf33),
    .D(\Y[7] [4]),
    .Q(\u_fir_pe6.rYin [4])
);

DFFPOSX1 _12490_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf32),
    .D(\Y[7] [5]),
    .Q(\u_fir_pe6.rYin [5])
);

DFFPOSX1 _12491_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf31),
    .D(\Y[7] [6]),
    .Q(\u_fir_pe6.rYin [6])
);

DFFPOSX1 _12492_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf30),
    .D(\Y[7] [7]),
    .Q(\u_fir_pe6.rYin [7])
);

DFFPOSX1 _12493_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf29),
    .D(\Y[7] [8]),
    .Q(\u_fir_pe6.rYin [8])
);

DFFPOSX1 _12494_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf28),
    .D(\Y[7] [9]),
    .Q(\u_fir_pe6.rYin [9])
);

DFFPOSX1 _12495_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf27),
    .D(\Y[7] [10]),
    .Q(\u_fir_pe6.rYin [10])
);

DFFPOSX1 _12496_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf26),
    .D(\Y[7] [11]),
    .Q(\u_fir_pe6.rYin [11])
);

DFFPOSX1 _12497_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf25),
    .D(\Y[7] [12]),
    .Q(\u_fir_pe6.rYin [12])
);

DFFPOSX1 _12498_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf24),
    .D(\Y[7] [13]),
    .Q(\u_fir_pe6.rYin [13])
);

DFFPOSX1 _12499_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf23),
    .D(\Y[7] [14]),
    .Q(\u_fir_pe6.rYin [14])
);

DFFPOSX1 _12500_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf22),
    .D(\Y[7] [15]),
    .Q(\u_fir_pe6.rYin [15])
);

DFFPOSX1 _12501_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf21),
    .D(_5573_[0]),
    .Q(\u_fir_pe6.mul [0])
);

DFFPOSX1 _12502_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf20),
    .D(_5574_[1]),
    .Q(\u_fir_pe6.mul [1])
);

DFFPOSX1 _12503_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf19),
    .D(_5575_[2]),
    .Q(\u_fir_pe6.mul [2])
);

DFFPOSX1 _12504_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf18),
    .D(_5576_[3]),
    .Q(\u_fir_pe6.mul [3])
);

DFFPOSX1 _12505_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf17),
    .D(_5577_[4]),
    .Q(\u_fir_pe6.mul [4])
);

DFFPOSX1 _12506_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf16),
    .D(_5578_[5]),
    .Q(\u_fir_pe6.mul [5])
);

DFFPOSX1 _12507_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf15),
    .D(_5578_[6]),
    .Q(\u_fir_pe6.mul [6])
);

DFFPOSX1 _12508_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf14),
    .D(_5578_[7]),
    .Q(\u_fir_pe6.mul [7])
);

DFFPOSX1 _12509_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf13),
    .D(_5578_[8]),
    .Q(\u_fir_pe6.mul [8])
);

DFFPOSX1 _12510_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf12),
    .D(_5578_[9]),
    .Q(\u_fir_pe6.mul [9])
);

DFFPOSX1 _12511_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf11),
    .D(_5578_[10]),
    .Q(\u_fir_pe6.mul [10])
);

DFFPOSX1 _12512_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf10),
    .D(_5578_[11]),
    .Q(\u_fir_pe6.mul [11])
);

DFFPOSX1 _12513_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf9),
    .D(_5578_[12]),
    .Q(\u_fir_pe6.mul [12])
);

DFFPOSX1 _12514_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf8),
    .D(_5578_[13]),
    .Q(\u_fir_pe6.mul [13])
);

DFFPOSX1 _12515_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf7),
    .D(_5578_[14]),
    .Q(\u_fir_pe6.mul [14])
);

DFFPOSX1 _12516_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_5578_[15]),
    .Q(\u_fir_pe6.mul [15])
);

NAND2X1 _12517_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [0]),
    .B(gnd),
    .Y(_6268_)
);

AND2X2 _12518_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [1]),
    .B(gnd),
    .Y(_6279_)
);

INVX1 _12519_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6279_),
    .Y(_6289_)
);

NOR2X1 _12520_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6268_),
    .B(_6289_),
    .Y(_6299_)
);

NAND2X1 _12521_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [1]),
    .Y(_6310_)
);

NOR2X1 _12522_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6268_),
    .B(_6310_),
    .Y(_6319_)
);

AOI22X1 _12523_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [0]),
    .B(vdd),
    .C(\X[6] [1]),
    .D(gnd),
    .Y(_6329_)
);

NOR2X1 _12524_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6329_),
    .B(_6319_),
    .Y(_6339_)
);

INVX1 _12525_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [2]),
    .Y(_6349_)
);

INVX2 _12526_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_6357_)
);

NOR2X1 _12527_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6349_),
    .B(_6357_),
    .Y(_6359_)
);

NAND2X1 _12528_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6359_),
    .B(_6339_),
    .Y(_6360_)
);

INVX1 _12529_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6360_),
    .Y(_6361_)
);

NOR2X1 _12530_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6359_),
    .B(_6339_),
    .Y(_6362_)
);

NOR2X1 _12531_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6362_),
    .B(_6361_),
    .Y(_6363_)
);

NAND2X1 _12532_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6299_),
    .B(_6363_),
    .Y(_6364_)
);

INVX1 _12533_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6364_),
    .Y(_6365_)
);

NAND2X1 _12534_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6] [3]),
    .Y(_6366_)
);

INVX1 _12535_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6366_),
    .Y(_6367_)
);

NAND2X1 _12536_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6] [2]),
    .Y(_5579_)
);

INVX1 _12537_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5579_),
    .Y(_5580_)
);

NAND2X1 _12538_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [0]),
    .Y(_5581_)
);

OR2X2 _12539_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6310_),
    .B(_5581_),
    .Y(_5582_)
);

AOI22X1 _12540_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [0]),
    .C(vdd),
    .D(\X[6] [1]),
    .Y(_5583_)
);

INVX1 _12541_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5583_),
    .Y(_5584_)
);

NAND3X1 _12542_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5580_),
    .B(_5584_),
    .C(_5582_),
    .Y(_5585_)
);

NOR2X1 _12543_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6310_),
    .B(_5581_),
    .Y(_5586_)
);

OAI21X1 _12544_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5583_),
    .B(_5586_),
    .C(_5579_),
    .Y(_5587_)
);

NAND3X1 _12545_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6319_),
    .B(_5587_),
    .C(_5585_),
    .Y(_5588_)
);

INVX1 _12546_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6319_),
    .Y(_5589_)
);

NAND3X1 _12547_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5579_),
    .B(_5584_),
    .C(_5582_),
    .Y(_5590_)
);

OAI21X1 _12548_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5583_),
    .B(_5586_),
    .C(_5580_),
    .Y(_5591_)
);

NAND3X1 _12549_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5589_),
    .B(_5591_),
    .C(_5590_),
    .Y(_5592_)
);

NAND3X1 _12550_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6367_),
    .B(_5592_),
    .C(_5588_),
    .Y(_5593_)
);

INVX2 _12551_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [3]),
    .Y(_5594_)
);

NAND2X1 _12552_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5592_),
    .B(_5588_),
    .Y(_5595_)
);

OAI21X1 _12553_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6357_),
    .B(_5594_),
    .C(_5595_),
    .Y(_5596_)
);

NAND2X1 _12554_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5593_),
    .B(_5596_),
    .Y(_5597_)
);

NAND2X1 _12555_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6360_),
    .B(_5597_),
    .Y(_5598_)
);

NAND3X1 _12556_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6361_),
    .B(_5593_),
    .C(_5596_),
    .Y(_5599_)
);

NAND3X1 _12557_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5599_),
    .B(_6365_),
    .C(_5598_),
    .Y(_5600_)
);

INVX1 _12558_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5600_),
    .Y(_5601_)
);

AOI21X1 _12559_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5598_),
    .B(_5599_),
    .C(_6365_),
    .Y(_5602_)
);

NOR2X1 _12560_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5602_),
    .B(_5601_),
    .Y(_6373_[3])
);

NAND2X1 _12561_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [0]),
    .B(gnd),
    .Y(_5603_)
);

NAND2X1 _12562_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [4]),
    .B(gnd),
    .Y(_5604_)
);

NOR2X1 _12563_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5603_),
    .B(_5604_),
    .Y(_5605_)
);

AOI22X1 _12564_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [0]),
    .B(gnd),
    .C(gnd),
    .D(\X[6] [4]),
    .Y(_5606_)
);

NOR2X1 _12565_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5606_),
    .B(_5605_),
    .Y(_5607_)
);

INVX1 _12566_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5607_),
    .Y(_5608_)
);

NAND2X1 _12567_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [0]),
    .B(vdd),
    .Y(_5609_)
);

NAND2X1 _12568_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [1]),
    .Y(_5610_)
);

OAI22X1 _12569_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5609_),
    .B(_5610_),
    .C(_5579_),
    .D(_5583_),
    .Y(_5611_)
);

NAND2X1 _12570_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6] [3]),
    .Y(_5612_)
);

INVX1 _12571_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5612_),
    .Y(_5613_)
);

AND2X2 _12572_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [1]),
    .Y(_5614_)
);

AND2X2 _12573_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [2]),
    .Y(_5615_)
);

NAND2X1 _12574_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5614_),
    .B(_5615_),
    .Y(_5616_)
);

AOI22X1 _12575_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [1]),
    .C(vdd),
    .D(\X[6] [2]),
    .Y(_5617_)
);

INVX1 _12576_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5617_),
    .Y(_5618_)
);

NAND3X1 _12577_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5613_),
    .B(_5618_),
    .C(_5616_),
    .Y(_5619_)
);

NAND3X1 _12578_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [2]),
    .C(_5610_),
    .Y(_5620_)
);

NAND2X1 _12579_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [2]),
    .Y(_5621_)
);

NAND3X1 _12580_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [1]),
    .C(_5621_),
    .Y(_5622_)
);

NAND3X1 _12581_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5612_),
    .B(_5620_),
    .C(_5622_),
    .Y(_5623_)
);

NAND3X1 _12582_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5611_),
    .B(_5623_),
    .C(_5619_),
    .Y(_5624_)
);

INVX1 _12583_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5611_),
    .Y(_5625_)
);

NAND2X1 _12584_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5623_),
    .B(_5619_),
    .Y(_5626_)
);

NAND2X1 _12585_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5625_),
    .B(_5626_),
    .Y(_5627_)
);

NAND3X1 _12586_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5608_),
    .B(_5624_),
    .C(_5627_),
    .Y(_5628_)
);

NAND2X1 _12587_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5611_),
    .B(_5626_),
    .Y(_5629_)
);

NAND3X1 _12588_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5619_),
    .B(_5623_),
    .C(_5625_),
    .Y(_5630_)
);

NAND3X1 _12589_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5607_),
    .B(_5630_),
    .C(_5629_),
    .Y(_5631_)
);

AOI22X1 _12590_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5588_),
    .B(_5593_),
    .C(_5628_),
    .D(_5631_),
    .Y(_5632_)
);

INVX1 _12591_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5632_),
    .Y(_5633_)
);

NAND2X1 _12592_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5588_),
    .B(_5593_),
    .Y(_5634_)
);

NAND2X1 _12593_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5628_),
    .B(_5631_),
    .Y(_5635_)
);

OR2X2 _12594_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5635_),
    .B(_5634_),
    .Y(_5636_)
);

NAND2X1 _12595_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5633_),
    .B(_5636_),
    .Y(_5637_)
);

OAI21X1 _12596_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6360_),
    .B(_5597_),
    .C(_5600_),
    .Y(_5638_)
);

OR2X2 _12597_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5638_),
    .B(_5637_),
    .Y(_5639_)
);

NAND3X1 _12598_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5607_),
    .B(_5624_),
    .C(_5627_),
    .Y(_5640_)
);

INVX1 _12599_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5624_),
    .Y(_5641_)
);

AOI21X1 _12600_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5619_),
    .B(_5623_),
    .C(_5611_),
    .Y(_5642_)
);

OAI21X1 _12601_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5642_),
    .B(_5641_),
    .C(_5608_),
    .Y(_5643_)
);

AOI21X1 _12602_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5640_),
    .B(_5643_),
    .C(_5634_),
    .Y(_5644_)
);

OAI21X1 _12603_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5632_),
    .B(_5644_),
    .C(_5638_),
    .Y(_5645_)
);

NAND2X1 _12604_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5645_),
    .B(_5639_),
    .Y(_6374_[4])
);

NOR2X1 _12605_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5600_),
    .B(_5637_),
    .Y(_5646_)
);

NOR3X1 _12606_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5632_),
    .B(_5599_),
    .C(_5644_),
    .Y(_5647_)
);

OAI21X1 _12607_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5608_),
    .B(_5642_),
    .C(_5624_),
    .Y(_5648_)
);

NAND2X1 _12608_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [0]),
    .B(gnd),
    .Y(_5649_)
);

INVX1 _12609_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5649_),
    .Y(_5650_)
);

AND2X2 _12610_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6]_5_bF$buf3 ),
    .Y(_5651_)
);

NAND2X1 _12611_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6279_),
    .B(_5651_),
    .Y(_5652_)
);

INVX2 _12612_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6]_5_bF$buf2 ),
    .Y(_5653_)
);

NAND2X1 _12613_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [1]),
    .B(gnd),
    .Y(_5654_)
);

OAI21X1 _12614_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6357_),
    .B(_5653_),
    .C(_5654_),
    .Y(_5655_)
);

NAND3X1 _12615_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5655_),
    .B(_5650_),
    .C(_5652_),
    .Y(_5656_)
);

NAND3X1 _12616_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6]_5_bF$buf1 ),
    .C(_5654_),
    .Y(_5657_)
);

NAND2X1 _12617_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6]_5_bF$buf0 ),
    .Y(_5658_)
);

NAND3X1 _12618_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [1]),
    .B(gnd),
    .C(_5658_),
    .Y(_5659_)
);

NAND3X1 _12619_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5649_),
    .B(_5657_),
    .C(_5659_),
    .Y(_5660_)
);

AND2X2 _12620_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5656_),
    .B(_5660_),
    .Y(_5661_)
);

NAND2X1 _12621_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [2]),
    .Y(_5662_)
);

OAI22X1 _12622_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6310_),
    .B(_5662_),
    .C(_5612_),
    .D(_5617_),
    .Y(_5663_)
);

NAND2X1 _12623_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6] [4]),
    .Y(_5664_)
);

INVX1 _12624_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5664_),
    .Y(_5665_)
);

AND2X2 _12625_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [3]),
    .Y(_5666_)
);

NAND2X1 _12626_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5615_),
    .B(_5666_),
    .Y(_5667_)
);

INVX1 _12627_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .Y(_5668_)
);

OAI21X1 _12628_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5668_),
    .B(_5594_),
    .C(_5662_),
    .Y(_5669_)
);

NAND3X1 _12629_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5665_),
    .B(_5669_),
    .C(_5667_),
    .Y(_5670_)
);

NAND3X1 _12630_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [3]),
    .C(_5662_),
    .Y(_5671_)
);

NAND2X1 _12631_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [3]),
    .Y(_5672_)
);

NAND3X1 _12632_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [2]),
    .C(_5672_),
    .Y(_5673_)
);

NAND3X1 _12633_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5664_),
    .B(_5671_),
    .C(_5673_),
    .Y(_5674_)
);

NAND3X1 _12634_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5663_),
    .B(_5674_),
    .C(_5670_),
    .Y(_5675_)
);

INVX1 _12635_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5663_),
    .Y(_5676_)
);

AOI21X1 _12636_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5671_),
    .B(_5673_),
    .C(_5664_),
    .Y(_5677_)
);

AOI22X1 _12637_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6] [4]),
    .C(_5667_),
    .D(_5669_),
    .Y(_5678_)
);

OAI21X1 _12638_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5677_),
    .B(_5678_),
    .C(_5676_),
    .Y(_5679_)
);

NAND3X1 _12639_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5675_),
    .B(_5661_),
    .C(_5679_),
    .Y(_5680_)
);

NAND2X1 _12640_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5660_),
    .B(_5656_),
    .Y(_5681_)
);

OAI21X1 _12641_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5677_),
    .B(_5678_),
    .C(_5663_),
    .Y(_5682_)
);

NAND3X1 _12642_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5674_),
    .B(_5670_),
    .C(_5676_),
    .Y(_5683_)
);

NAND3X1 _12643_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5681_),
    .B(_5683_),
    .C(_5682_),
    .Y(_5684_)
);

NAND3X1 _12644_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5680_),
    .B(_5684_),
    .C(_5648_),
    .Y(_5685_)
);

AOI21X1 _12645_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5607_),
    .B(_5627_),
    .C(_5641_),
    .Y(_5686_)
);

AOI21X1 _12646_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5682_),
    .B(_5683_),
    .C(_5681_),
    .Y(_5687_)
);

AOI21X1 _12647_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5679_),
    .B(_5675_),
    .C(_5661_),
    .Y(_5688_)
);

OAI21X1 _12648_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5687_),
    .B(_5688_),
    .C(_5686_),
    .Y(_5689_)
);

NAND3X1 _12649_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5605_),
    .B(_5685_),
    .C(_5689_),
    .Y(_5690_)
);

INVX1 _12650_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5605_),
    .Y(_5691_)
);

OAI21X1 _12651_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5687_),
    .B(_5688_),
    .C(_5648_),
    .Y(_5692_)
);

NAND3X1 _12652_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5680_),
    .B(_5684_),
    .C(_5686_),
    .Y(_5693_)
);

NAND3X1 _12653_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5691_),
    .B(_5692_),
    .C(_5693_),
    .Y(_5694_)
);

NAND3X1 _12654_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5632_),
    .B(_5690_),
    .C(_5694_),
    .Y(_5695_)
);

NAND3X1 _12655_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5691_),
    .B(_5685_),
    .C(_5689_),
    .Y(_5696_)
);

NAND3X1 _12656_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5605_),
    .B(_5692_),
    .C(_5693_),
    .Y(_5697_)
);

NAND3X1 _12657_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5633_),
    .B(_5696_),
    .C(_5697_),
    .Y(_5698_)
);

NAND3X1 _12658_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5695_),
    .B(_5698_),
    .C(_5647_),
    .Y(_5699_)
);

INVX1 _12659_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5599_),
    .Y(_5700_)
);

NAND3X1 _12660_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5700_),
    .B(_5633_),
    .C(_5636_),
    .Y(_5701_)
);

NAND3X1 _12661_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5633_),
    .B(_5690_),
    .C(_5694_),
    .Y(_5702_)
);

NAND3X1 _12662_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5632_),
    .B(_5696_),
    .C(_5697_),
    .Y(_5703_)
);

NAND3X1 _12663_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5702_),
    .B(_5703_),
    .C(_5701_),
    .Y(_5704_)
);

NAND3X1 _12664_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5699_),
    .B(_5704_),
    .C(_5646_),
    .Y(_5705_)
);

INVX1 _12665_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5646_),
    .Y(_5706_)
);

INVX1 _12666_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5699_),
    .Y(_5707_)
);

INVX1 _12667_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5704_),
    .Y(_5708_)
);

OAI21X1 _12668_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5707_),
    .B(_5708_),
    .C(_5706_),
    .Y(_5709_)
);

AND2X2 _12669_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5709_),
    .B(_5705_),
    .Y(_6375_[5])
);

AND2X2 _12670_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [0]),
    .B(gnd),
    .Y(_5710_)
);

NAND2X1 _12671_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6]_5_bF$buf3 ),
    .Y(_5711_)
);

OAI21X1 _12672_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6289_),
    .B(_5711_),
    .C(_5656_),
    .Y(_5712_)
);

OR2X2 _12673_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5712_),
    .B(_5710_),
    .Y(_5713_)
);

NAND2X1 _12674_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5710_),
    .B(_5712_),
    .Y(_5714_)
);

NAND2X1 _12675_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5714_),
    .B(_5713_),
    .Y(_5715_)
);

AOI21X1 _12676_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5670_),
    .B(_5674_),
    .C(_5663_),
    .Y(_5716_)
);

OAI21X1 _12677_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5681_),
    .B(_5716_),
    .C(_5675_),
    .Y(_5717_)
);

NAND2X1 _12678_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [1]),
    .B(gnd),
    .Y(_5718_)
);

INVX1 _12679_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5718_),
    .Y(_5719_)
);

AND2X2 _12680_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [2]),
    .B(gnd),
    .Y(_5720_)
);

AND2X2 _12681_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6] [6]),
    .Y(_5721_)
);

NAND2X1 _12682_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5720_),
    .B(_5721_),
    .Y(_5722_)
);

INVX2 _12683_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [6]),
    .Y(_5723_)
);

NAND2X1 _12684_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [2]),
    .B(gnd),
    .Y(_5724_)
);

OAI21X1 _12685_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6357_),
    .B(_5723_),
    .C(_5724_),
    .Y(_5725_)
);

NAND3X1 _12686_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5725_),
    .B(_5719_),
    .C(_5722_),
    .Y(_5726_)
);

NAND3X1 _12687_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6] [6]),
    .C(_5724_),
    .Y(_5727_)
);

NAND2X1 _12688_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6] [6]),
    .Y(_5728_)
);

NAND2X1 _12689_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5728_),
    .B(_5720_),
    .Y(_5729_)
);

NAND3X1 _12690_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5718_),
    .B(_5727_),
    .C(_5729_),
    .Y(_5730_)
);

AND2X2 _12691_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5726_),
    .B(_5730_),
    .Y(_5731_)
);

NAND2X1 _12692_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [3]),
    .Y(_5732_)
);

AOI22X1 _12693_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [2]),
    .C(vdd),
    .D(\X[6] [3]),
    .Y(_5733_)
);

OAI22X1 _12694_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5621_),
    .B(_5732_),
    .C(_5664_),
    .D(_5733_),
    .Y(_5734_)
);

NAND2X1 _12695_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6]_5_bF$buf2 ),
    .Y(_5735_)
);

INVX1 _12696_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5735_),
    .Y(_5736_)
);

AND2X2 _12697_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [4]),
    .Y(_5737_)
);

NAND2X1 _12698_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5666_),
    .B(_5737_),
    .Y(_5738_)
);

AOI22X1 _12699_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [3]),
    .C(vdd),
    .D(\X[6] [4]),
    .Y(_5739_)
);

INVX1 _12700_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5739_),
    .Y(_5740_)
);

NAND3X1 _12701_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5736_),
    .B(_5740_),
    .C(_5738_),
    .Y(_5741_)
);

NAND3X1 _12702_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [4]),
    .C(_5732_),
    .Y(_5742_)
);

NAND2X1 _12703_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [4]),
    .Y(_5743_)
);

NAND3X1 _12704_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [3]),
    .C(_5743_),
    .Y(_5744_)
);

NAND3X1 _12705_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5735_),
    .B(_5742_),
    .C(_5744_),
    .Y(_5745_)
);

NAND3X1 _12706_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5734_),
    .B(_5745_),
    .C(_5741_),
    .Y(_5746_)
);

INVX1 _12707_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5734_),
    .Y(_5747_)
);

AOI21X1 _12708_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5742_),
    .B(_5744_),
    .C(_5735_),
    .Y(_5748_)
);

AOI22X1 _12709_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6]_5_bF$buf1 ),
    .C(_5738_),
    .D(_5740_),
    .Y(_5749_)
);

OAI21X1 _12710_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5748_),
    .B(_5749_),
    .C(_5747_),
    .Y(_5750_)
);

NAND3X1 _12711_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5746_),
    .B(_5731_),
    .C(_5750_),
    .Y(_5751_)
);

NAND2X1 _12712_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5730_),
    .B(_5726_),
    .Y(_5752_)
);

OAI21X1 _12713_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5748_),
    .B(_5749_),
    .C(_5734_),
    .Y(_5753_)
);

NAND3X1 _12714_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5741_),
    .B(_5745_),
    .C(_5747_),
    .Y(_5754_)
);

NAND3X1 _12715_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5752_),
    .B(_5754_),
    .C(_5753_),
    .Y(_5755_)
);

NAND3X1 _12716_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5751_),
    .B(_5717_),
    .C(_5755_),
    .Y(_5756_)
);

INVX1 _12717_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5675_),
    .Y(_5757_)
);

AOI21X1 _12718_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5661_),
    .B(_5679_),
    .C(_5757_),
    .Y(_5758_)
);

AOI21X1 _12719_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5753_),
    .B(_5754_),
    .C(_5752_),
    .Y(_5759_)
);

AOI21X1 _12720_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5750_),
    .B(_5746_),
    .C(_5731_),
    .Y(_5760_)
);

OAI21X1 _12721_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5759_),
    .B(_5760_),
    .C(_5758_),
    .Y(_5761_)
);

NAND3X1 _12722_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5715_),
    .B(_5756_),
    .C(_5761_),
    .Y(_5762_)
);

AND2X2 _12723_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5713_),
    .B(_5714_),
    .Y(_5763_)
);

OAI21X1 _12724_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5759_),
    .B(_5760_),
    .C(_5717_),
    .Y(_5764_)
);

NAND3X1 _12725_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5751_),
    .B(_5755_),
    .C(_5758_),
    .Y(_5765_)
);

NAND3X1 _12726_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5763_),
    .B(_5764_),
    .C(_5765_),
    .Y(_5766_)
);

AOI22X1 _12727_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5690_),
    .B(_5685_),
    .C(_5762_),
    .D(_5766_),
    .Y(_5767_)
);

AOI21X1 _12728_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5680_),
    .B(_5684_),
    .C(_5648_),
    .Y(_5768_)
);

OAI21X1 _12729_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5691_),
    .B(_5768_),
    .C(_5685_),
    .Y(_5769_)
);

NAND3X1 _12730_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5763_),
    .B(_5756_),
    .C(_5761_),
    .Y(_5770_)
);

NAND3X1 _12731_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5715_),
    .B(_5764_),
    .C(_5765_),
    .Y(_5771_)
);

AOI21X1 _12732_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5771_),
    .B(_5770_),
    .C(_5769_),
    .Y(_5772_)
);

OAI21X1 _12733_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5772_),
    .B(_5767_),
    .C(_5695_),
    .Y(_5773_)
);

AOI21X1 _12734_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5697_),
    .B(_5696_),
    .C(_5633_),
    .Y(_5774_)
);

NAND3X1 _12735_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5769_),
    .B(_5770_),
    .C(_5771_),
    .Y(_5775_)
);

INVX1 _12736_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5685_),
    .Y(_5776_)
);

AOI21X1 _12737_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5605_),
    .B(_5689_),
    .C(_5776_),
    .Y(_5777_)
);

AOI21X1 _12738_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5765_),
    .B(_5764_),
    .C(_5715_),
    .Y(_5778_)
);

AOI21X1 _12739_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5761_),
    .B(_5756_),
    .C(_5763_),
    .Y(_5779_)
);

OAI21X1 _12740_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5778_),
    .B(_5779_),
    .C(_5777_),
    .Y(_5780_)
);

NAND3X1 _12741_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5774_),
    .B(_5775_),
    .C(_5780_),
    .Y(_5781_)
);

NAND2X1 _12742_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5781_),
    .B(_5773_),
    .Y(_5782_)
);

AOI21X1 _12743_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5699_),
    .B(_5705_),
    .C(_5782_),
    .Y(_5783_)
);

OAI21X1 _12744_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5708_),
    .B(_5706_),
    .C(_5699_),
    .Y(_5784_)
);

AOI21X1 _12745_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5773_),
    .B(_5781_),
    .C(_5784_),
    .Y(_5785_)
);

NOR2X1 _12746_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5783_),
    .B(_5785_),
    .Y(_6375_[6])
);

INVX1 _12747_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5781_),
    .Y(_5786_)
);

AOI21X1 _12748_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5751_),
    .B(_5755_),
    .C(_5717_),
    .Y(_5787_)
);

OAI21X1 _12749_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5715_),
    .B(_5787_),
    .C(_5756_),
    .Y(_5788_)
);

NAND2X1 _12750_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [0]),
    .B(gnd),
    .Y(_5789_)
);

INVX1 _12751_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5789_),
    .Y(_5790_)
);

NAND2X1 _12752_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [1]),
    .B(gnd),
    .Y(_5791_)
);

INVX1 _12753_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5791_),
    .Y(_5792_)
);

AND2X2 _12754_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5724_),
    .B(_5728_),
    .Y(_5793_)
);

OAI21X1 _12755_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5718_),
    .B(_5793_),
    .C(_5722_),
    .Y(_5794_)
);

NAND2X1 _12756_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5792_),
    .B(_5794_),
    .Y(_5795_)
);

NAND3X1 _12757_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5722_),
    .B(_5791_),
    .C(_5726_),
    .Y(_5796_)
);

NAND3X1 _12758_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5790_),
    .B(_5796_),
    .C(_5795_),
    .Y(_5797_)
);

AOI21X1 _12759_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5726_),
    .B(_5722_),
    .C(_5791_),
    .Y(_5798_)
);

NOR2X1 _12760_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5792_),
    .B(_5794_),
    .Y(_5799_)
);

OAI21X1 _12761_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5798_),
    .B(_5799_),
    .C(_5789_),
    .Y(_5800_)
);

NAND2X1 _12762_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5797_),
    .B(_5800_),
    .Y(_5801_)
);

AOI21X1 _12763_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5741_),
    .B(_5745_),
    .C(_5734_),
    .Y(_5802_)
);

OAI21X1 _12764_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5752_),
    .B(_5802_),
    .C(_5746_),
    .Y(_5803_)
);

NAND2X1 _12765_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [2]),
    .B(gnd),
    .Y(_5804_)
);

INVX1 _12766_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5804_),
    .Y(_5805_)
);

AND2X2 _12767_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [3]),
    .B(gnd),
    .Y(_5806_)
);

AND2X2 _12768_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6] [7]),
    .Y(_5807_)
);

NAND2X1 _12769_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5806_),
    .B(_5807_),
    .Y(_5808_)
);

AOI22X1 _12770_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6] [7]),
    .C(\X[6] [3]),
    .D(gnd),
    .Y(_5809_)
);

INVX1 _12771_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5809_),
    .Y(_5810_)
);

NAND3X1 _12772_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5805_),
    .B(_5810_),
    .C(_5808_),
    .Y(_5811_)
);

INVX1 _12773_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_5812_)
);

OAI21X1 _12774_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5594_),
    .B(_5812_),
    .C(_5807_),
    .Y(_5813_)
);

INVX1 _12775_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [7]),
    .Y(_5814_)
);

OAI21X1 _12776_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6357_),
    .B(_5814_),
    .C(_5806_),
    .Y(_5815_)
);

NAND3X1 _12777_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5804_),
    .B(_5813_),
    .C(_5815_),
    .Y(_5816_)
);

NAND2X1 _12778_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5811_),
    .B(_5816_),
    .Y(_5817_)
);

OAI21X1 _12779_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5735_),
    .B(_5739_),
    .C(_5738_),
    .Y(_5818_)
);

NAND2X1 _12780_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6] [6]),
    .Y(_5819_)
);

NAND2X1 _12781_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [4]),
    .Y(_5820_)
);

AND2X2 _12782_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6]_5_bF$buf0 ),
    .Y(_5821_)
);

NAND2X1 _12783_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5820_),
    .B(_5821_),
    .Y(_5822_)
);

OAI21X1 _12784_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5668_),
    .B(_5653_),
    .C(_5737_),
    .Y(_5823_)
);

AOI21X1 _12785_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5823_),
    .B(_5822_),
    .C(_5819_),
    .Y(_5824_)
);

INVX1 _12786_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5819_),
    .Y(_5825_)
);

NAND2X1 _12787_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5737_),
    .B(_5821_),
    .Y(_5826_)
);

AOI22X1 _12788_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [4]),
    .C(vdd),
    .D(\X[6]_5_bF$buf3 ),
    .Y(_5827_)
);

INVX1 _12789_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5827_),
    .Y(_5828_)
);

AOI21X1 _12790_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5826_),
    .B(_5828_),
    .C(_5825_),
    .Y(_5829_)
);

OAI21X1 _12791_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5829_),
    .B(_5824_),
    .C(_5818_),
    .Y(_5830_)
);

AOI22X1 _12792_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5666_),
    .B(_5737_),
    .C(_5740_),
    .D(_5736_),
    .Y(_5831_)
);

NAND3X1 _12793_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5825_),
    .B(_5828_),
    .C(_5826_),
    .Y(_5832_)
);

NAND2X1 _12794_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6]_5_bF$buf2 ),
    .Y(_5833_)
);

NOR2X1 _12795_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5820_),
    .B(_5833_),
    .Y(_5834_)
);

OAI21X1 _12796_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5827_),
    .B(_5834_),
    .C(_5819_),
    .Y(_5835_)
);

NAND3X1 _12797_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5832_),
    .B(_5831_),
    .C(_5835_),
    .Y(_5836_)
);

AOI21X1 _12798_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5830_),
    .B(_5836_),
    .C(_5817_),
    .Y(_5837_)
);

AND2X2 _12799_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5816_),
    .B(_5811_),
    .Y(_5838_)
);

NAND3X1 _12800_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5818_),
    .B(_5832_),
    .C(_5835_),
    .Y(_5839_)
);

OAI21X1 _12801_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5829_),
    .B(_5824_),
    .C(_5831_),
    .Y(_5840_)
);

AOI21X1 _12802_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5840_),
    .B(_5839_),
    .C(_5838_),
    .Y(_5841_)
);

OAI21X1 _12803_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5837_),
    .B(_5841_),
    .C(_5803_),
    .Y(_5842_)
);

INVX1 _12804_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5746_),
    .Y(_5843_)
);

AOI21X1 _12805_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5731_),
    .B(_5750_),
    .C(_5843_),
    .Y(_5844_)
);

NAND3X1 _12806_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5839_),
    .B(_5838_),
    .C(_5840_),
    .Y(_5845_)
);

NAND3X1 _12807_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5817_),
    .B(_5836_),
    .C(_5830_),
    .Y(_5846_)
);

NAND3X1 _12808_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5845_),
    .B(_5846_),
    .C(_5844_),
    .Y(_5847_)
);

AOI21X1 _12809_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5847_),
    .B(_5842_),
    .C(_5801_),
    .Y(_5848_)
);

AND2X2 _12810_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5800_),
    .B(_5797_),
    .Y(_5849_)
);

NAND3X1 _12811_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5803_),
    .B(_5845_),
    .C(_5846_),
    .Y(_5850_)
);

OAI21X1 _12812_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5837_),
    .B(_5841_),
    .C(_5844_),
    .Y(_5851_)
);

AOI21X1 _12813_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5851_),
    .B(_5850_),
    .C(_5849_),
    .Y(_5852_)
);

OAI21X1 _12814_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5852_),
    .B(_5848_),
    .C(_5788_),
    .Y(_5853_)
);

INVX1 _12815_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5756_),
    .Y(_5854_)
);

AOI21X1 _12816_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5763_),
    .B(_5761_),
    .C(_5854_),
    .Y(_5855_)
);

NAND3X1 _12817_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5850_),
    .B(_5849_),
    .C(_5851_),
    .Y(_5856_)
);

NAND3X1 _12818_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5801_),
    .B(_5842_),
    .C(_5847_),
    .Y(_5857_)
);

NAND3X1 _12819_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5856_),
    .B(_5857_),
    .C(_5855_),
    .Y(_5858_)
);

AOI21X1 _12820_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5858_),
    .B(_5853_),
    .C(_5714_),
    .Y(_5859_)
);

INVX1 _12821_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5714_),
    .Y(_5860_)
);

NAND3X1 _12822_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5788_),
    .B(_5856_),
    .C(_5857_),
    .Y(_5861_)
);

OAI21X1 _12823_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5848_),
    .B(_5852_),
    .C(_5855_),
    .Y(_5862_)
);

AOI21X1 _12824_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5862_),
    .B(_5861_),
    .C(_5860_),
    .Y(_5863_)
);

OAI21X1 _12825_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5863_),
    .B(_5859_),
    .C(_5775_),
    .Y(_5864_)
);

NAND3X1 _12826_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5860_),
    .B(_5861_),
    .C(_5862_),
    .Y(_5865_)
);

NAND3X1 _12827_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5714_),
    .B(_5853_),
    .C(_5858_),
    .Y(_5866_)
);

NAND3X1 _12828_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5767_),
    .B(_5865_),
    .C(_5866_),
    .Y(_5867_)
);

AND2X2 _12829_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5864_),
    .B(_5867_),
    .Y(_5868_)
);

OAI21X1 _12830_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5786_),
    .B(_5783_),
    .C(_5868_),
    .Y(_5869_)
);

NOR2X1 _12831_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5786_),
    .B(_5783_),
    .Y(_5870_)
);

AOI21X1 _12832_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5866_),
    .B(_5865_),
    .C(_5767_),
    .Y(_5871_)
);

INVX1 _12833_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5867_),
    .Y(_5872_)
);

OAI21X1 _12834_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5871_),
    .B(_5872_),
    .C(_5870_),
    .Y(_5873_)
);

AND2X2 _12835_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5873_),
    .B(_5869_),
    .Y(_6375_[7])
);

NAND3X1 _12836_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5864_),
    .B(_5867_),
    .C(_5783_),
    .Y(_5874_)
);

AOI21X1 _12837_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5786_),
    .B(_5864_),
    .C(_5872_),
    .Y(_5875_)
);

NAND2X1 _12838_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5875_),
    .B(_5874_),
    .Y(_5876_)
);

INVX1 _12839_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5861_),
    .Y(_5877_)
);

AOI21X1 _12840_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5860_),
    .B(_5862_),
    .C(_5877_),
    .Y(_5878_)
);

OAI21X1 _12841_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5789_),
    .B(_5799_),
    .C(_5795_),
    .Y(_5879_)
);

INVX1 _12842_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5879_),
    .Y(_5880_)
);

AOI21X1 _12843_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5845_),
    .B(_5846_),
    .C(_5803_),
    .Y(_5881_)
);

OAI21X1 _12844_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5801_),
    .B(_5881_),
    .C(_5850_),
    .Y(_5882_)
);

NAND2X1 _12845_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [1]),
    .B(gnd),
    .Y(_5883_)
);

INVX2 _12846_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_5884_)
);

NOR2X1 _12847_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6349_),
    .B(_5884_),
    .Y(_5885_)
);

OAI21X1 _12848_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5804_),
    .B(_5809_),
    .C(_5808_),
    .Y(_5886_)
);

NOR2X1 _12849_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5885_),
    .B(_5886_),
    .Y(_5887_)
);

AND2X2 _12850_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5886_),
    .B(_5885_),
    .Y(_5888_)
);

OAI21X1 _12851_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5887_),
    .B(_5888_),
    .C(_5883_),
    .Y(_5889_)
);

INVX1 _12852_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5883_),
    .Y(_5890_)
);

OR2X2 _12853_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5886_),
    .B(_5885_),
    .Y(_5891_)
);

NAND2X1 _12854_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5885_),
    .B(_5886_),
    .Y(_5892_)
);

NAND3X1 _12855_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5890_),
    .B(_5892_),
    .C(_5891_),
    .Y(_5893_)
);

NAND2X1 _12856_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5889_),
    .B(_5893_),
    .Y(_5894_)
);

AOI21X1 _12857_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5835_),
    .B(_5832_),
    .C(_5818_),
    .Y(_5895_)
);

OAI21X1 _12858_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5817_),
    .B(_5895_),
    .C(_5839_),
    .Y(_5896_)
);

NAND2X1 _12859_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [3]),
    .B(gnd),
    .Y(_5897_)
);

INVX1 _12860_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_5898_)
);

OAI21X1 _12861_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5594_),
    .B(_5898_),
    .C(_5604_),
    .Y(_5899_)
);

NAND2X1 _12862_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [4]),
    .B(gnd),
    .Y(_5900_)
);

OAI21X1 _12863_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5897_),
    .B(_5900_),
    .C(_5899_),
    .Y(_5901_)
);

OAI21X1 _12864_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5819_),
    .B(_5827_),
    .C(_5826_),
    .Y(_5902_)
);

NAND2X1 _12865_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6] [7]),
    .Y(_5903_)
);

NAND2X1 _12866_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6]_5_bF$buf1 ),
    .Y(_5904_)
);

NAND3X1 _12867_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [6]),
    .C(_5904_),
    .Y(_5905_)
);

AND2X2 _12868_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6]_5_bF$buf0 ),
    .Y(_5906_)
);

OAI21X1 _12869_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5668_),
    .B(_5723_),
    .C(_5906_),
    .Y(_5907_)
);

AOI21X1 _12870_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5907_),
    .B(_5905_),
    .C(_5903_),
    .Y(_5908_)
);

INVX1 _12871_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5903_),
    .Y(_5909_)
);

AND2X2 _12872_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [6]),
    .Y(_5910_)
);

NAND2X1 _12873_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5906_),
    .B(_5910_),
    .Y(_5911_)
);

NAND2X1 _12874_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [6]),
    .Y(_5912_)
);

NAND2X1 _12875_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5904_),
    .B(_5912_),
    .Y(_5913_)
);

AOI21X1 _12876_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5911_),
    .B(_5913_),
    .C(_5909_),
    .Y(_5914_)
);

OAI21X1 _12877_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5914_),
    .B(_5908_),
    .C(_5902_),
    .Y(_5915_)
);

AOI21X1 _12878_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5825_),
    .B(_5828_),
    .C(_5834_),
    .Y(_5916_)
);

NAND3X1 _12879_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5909_),
    .B(_5913_),
    .C(_5911_),
    .Y(_5917_)
);

NAND3X1 _12880_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5903_),
    .B(_5905_),
    .C(_5907_),
    .Y(_5918_)
);

NAND3X1 _12881_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5917_),
    .B(_5918_),
    .C(_5916_),
    .Y(_5919_)
);

AOI21X1 _12882_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5915_),
    .B(_5919_),
    .C(_5901_),
    .Y(_5920_)
);

INVX1 _12883_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5901_),
    .Y(_5921_)
);

NAND3X1 _12884_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5902_),
    .B(_5917_),
    .C(_5918_),
    .Y(_5922_)
);

OAI21X1 _12885_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5914_),
    .B(_5908_),
    .C(_5916_),
    .Y(_5923_)
);

AOI21X1 _12886_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5923_),
    .B(_5922_),
    .C(_5921_),
    .Y(_5924_)
);

OAI21X1 _12887_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5920_),
    .B(_5924_),
    .C(_5896_),
    .Y(_5925_)
);

INVX1 _12888_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5839_),
    .Y(_5926_)
);

AOI21X1 _12889_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5838_),
    .B(_5840_),
    .C(_5926_),
    .Y(_5927_)
);

NAND3X1 _12890_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5921_),
    .B(_5922_),
    .C(_5923_),
    .Y(_5928_)
);

NAND3X1 _12891_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5901_),
    .B(_5919_),
    .C(_5915_),
    .Y(_5929_)
);

NAND3X1 _12892_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5928_),
    .B(_5929_),
    .C(_5927_),
    .Y(_5930_)
);

AOI21X1 _12893_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5930_),
    .B(_5925_),
    .C(_5894_),
    .Y(_5931_)
);

AND2X2 _12894_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5893_),
    .B(_5889_),
    .Y(_5932_)
);

NAND3X1 _12895_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5928_),
    .B(_5929_),
    .C(_5896_),
    .Y(_5933_)
);

OAI21X1 _12896_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5920_),
    .B(_5924_),
    .C(_5927_),
    .Y(_5934_)
);

AOI21X1 _12897_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5934_),
    .B(_5933_),
    .C(_5932_),
    .Y(_5935_)
);

OAI21X1 _12898_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5935_),
    .B(_5931_),
    .C(_5882_),
    .Y(_5936_)
);

INVX1 _12899_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5850_),
    .Y(_5937_)
);

AOI21X1 _12900_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5849_),
    .B(_5851_),
    .C(_5937_),
    .Y(_5938_)
);

NAND3X1 _12901_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5932_),
    .B(_5933_),
    .C(_5934_),
    .Y(_5939_)
);

NAND3X1 _12902_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5894_),
    .B(_5925_),
    .C(_5930_),
    .Y(_5940_)
);

NAND3X1 _12903_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5939_),
    .B(_5940_),
    .C(_5938_),
    .Y(_5941_)
);

AOI21X1 _12904_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5936_),
    .B(_5941_),
    .C(_5880_),
    .Y(_5942_)
);

NAND3X1 _12905_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5882_),
    .B(_5939_),
    .C(_5940_),
    .Y(_5943_)
);

OAI21X1 _12906_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5935_),
    .B(_5931_),
    .C(_5938_),
    .Y(_5944_)
);

AOI21X1 _12907_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5944_),
    .B(_5943_),
    .C(_5879_),
    .Y(_5945_)
);

OAI21X1 _12908_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5945_),
    .B(_5942_),
    .C(_5878_),
    .Y(_5946_)
);

AOI21X1 _12909_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5857_),
    .B(_5856_),
    .C(_5788_),
    .Y(_5947_)
);

OAI21X1 _12910_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5714_),
    .B(_5947_),
    .C(_5861_),
    .Y(_5948_)
);

NAND3X1 _12911_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5879_),
    .B(_5943_),
    .C(_5944_),
    .Y(_5949_)
);

NAND3X1 _12912_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5880_),
    .B(_5941_),
    .C(_5936_),
    .Y(_5950_)
);

NAND3X1 _12913_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5948_),
    .B(_5949_),
    .C(_5950_),
    .Y(_5951_)
);

NAND2X1 _12914_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5951_),
    .B(_5946_),
    .Y(_5952_)
);

NAND2X1 _12915_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5952_),
    .B(_5876_),
    .Y(_5953_)
);

OAI21X1 _12916_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5781_),
    .B(_5871_),
    .C(_5867_),
    .Y(_5954_)
);

AOI21X1 _12917_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5868_),
    .B(_5783_),
    .C(_5954_),
    .Y(_5955_)
);

AND2X2 _12918_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5946_),
    .B(_5951_),
    .Y(_5956_)
);

NAND2X1 _12919_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5956_),
    .B(_5955_),
    .Y(_5957_)
);

NAND2X1 _12920_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5953_),
    .B(_5957_),
    .Y(_6375_[8])
);

INVX1 _12921_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5951_),
    .Y(_5958_)
);

AOI21X1 _12922_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5876_),
    .B(_5946_),
    .C(_5958_),
    .Y(_5959_)
);

AOI21X1 _12923_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5940_),
    .B(_5939_),
    .C(_5882_),
    .Y(_5960_)
);

OAI21X1 _12924_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5880_),
    .B(_5960_),
    .C(_5943_),
    .Y(_5961_)
);

OAI21X1 _12925_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5883_),
    .B(_5887_),
    .C(_5892_),
    .Y(_5962_)
);

AOI21X1 _12926_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5928_),
    .B(_5929_),
    .C(_5896_),
    .Y(_5963_)
);

OAI21X1 _12927_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5894_),
    .B(_5963_),
    .C(_5933_),
    .Y(_5964_)
);

NAND2X1 _12928_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [2]),
    .B(gnd),
    .Y(_5965_)
);

NOR2X1 _12929_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5897_),
    .B(_5900_),
    .Y(_5966_)
);

NAND2X1 _12930_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_5966_),
    .Y(_5967_)
);

INVX1 _12931_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5967_),
    .Y(_5968_)
);

AOI21X1 _12932_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [3]),
    .B(gnd),
    .C(_5966_),
    .Y(_5969_)
);

OAI21X1 _12933_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5969_),
    .B(_5968_),
    .C(_5965_),
    .Y(_5970_)
);

INVX1 _12934_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5965_),
    .Y(_5971_)
);

INVX1 _12935_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5969_),
    .Y(_5972_)
);

NAND3X1 _12936_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5971_),
    .B(_5967_),
    .C(_5972_),
    .Y(_5973_)
);

AND2X2 _12937_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5973_),
    .B(_5970_),
    .Y(_5974_)
);

AOI21X1 _12938_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5918_),
    .B(_5917_),
    .C(_5902_),
    .Y(_5975_)
);

OAI21X1 _12939_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5901_),
    .B(_5975_),
    .C(_5922_),
    .Y(_5976_)
);

NOR2X1 _12940_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5711_),
    .B(_5900_),
    .Y(_5977_)
);

AND2X2 _12941_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5711_),
    .B(_5900_),
    .Y(_5978_)
);

NOR2X1 _12942_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5977_),
    .B(_5978_),
    .Y(_5979_)
);

NAND2X1 _12943_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [6]),
    .Y(_5980_)
);

AOI22X1 _12944_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6]_5_bF$buf3 ),
    .C(vdd),
    .D(\X[6] [6]),
    .Y(_5981_)
);

OAI22X1 _12945_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5833_),
    .B(_5980_),
    .C(_5903_),
    .D(_5981_),
    .Y(_5982_)
);

AOI22X1 _12946_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [6]),
    .C(vdd),
    .D(\X[6] [7]),
    .Y(_5983_)
);

AND2X2 _12947_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [7]),
    .Y(_5984_)
);

AOI21X1 _12948_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5910_),
    .B(_5984_),
    .C(_5983_),
    .Y(_5985_)
);

NAND2X1 _12949_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5985_),
    .B(_5982_),
    .Y(_5986_)
);

AND2X2 _12950_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [6]),
    .Y(_5987_)
);

AOI22X1 _12951_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5821_),
    .B(_5987_),
    .C(_5913_),
    .D(_5909_),
    .Y(_5988_)
);

NAND2X1 _12952_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [7]),
    .Y(_5989_)
);

NAND2X1 _12953_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5980_),
    .B(_5989_),
    .Y(_5990_)
);

NAND2X1 _12954_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [7]),
    .Y(_5991_)
);

OAI21X1 _12955_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5912_),
    .B(_5991_),
    .C(_5990_),
    .Y(_5992_)
);

NAND2X1 _12956_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5992_),
    .B(_5988_),
    .Y(_5993_)
);

NAND3X1 _12957_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5979_),
    .B(_5986_),
    .C(_5993_),
    .Y(_5994_)
);

NAND2X1 _12958_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6]_5_bF$buf2 ),
    .B(gnd),
    .Y(_5995_)
);

INVX1 _12959_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [4]),
    .Y(_5996_)
);

OAI21X1 _12960_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5996_),
    .B(_5898_),
    .C(_5711_),
    .Y(_5997_)
);

OAI21X1 _12961_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5604_),
    .B(_5995_),
    .C(_5997_),
    .Y(_5998_)
);

NAND2X1 _12962_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5982_),
    .B(_5992_),
    .Y(_5999_)
);

NAND2X1 _12963_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5985_),
    .B(_5988_),
    .Y(_6000_)
);

NAND3X1 _12964_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5998_),
    .B(_5999_),
    .C(_6000_),
    .Y(_6001_)
);

NAND3X1 _12965_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5994_),
    .B(_6001_),
    .C(_5976_),
    .Y(_6002_)
);

NAND2X1 _12966_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5994_),
    .B(_6001_),
    .Y(_6003_)
);

NAND3X1 _12967_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5922_),
    .B(_5928_),
    .C(_6003_),
    .Y(_6004_)
);

NAND3X1 _12968_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5974_),
    .B(_6002_),
    .C(_6004_),
    .Y(_6005_)
);

NAND2X1 _12969_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5970_),
    .B(_5973_),
    .Y(_6006_)
);

AOI21X1 _12970_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5922_),
    .B(_5928_),
    .C(_6003_),
    .Y(_6007_)
);

AOI21X1 _12971_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5994_),
    .B(_6001_),
    .C(_5976_),
    .Y(_6008_)
);

OAI21X1 _12972_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6008_),
    .B(_6007_),
    .C(_6006_),
    .Y(_6009_)
);

NAND3X1 _12973_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6005_),
    .B(_6009_),
    .C(_5964_),
    .Y(_6010_)
);

INVX1 _12974_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5933_),
    .Y(_6011_)
);

AOI21X1 _12975_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5932_),
    .B(_5934_),
    .C(_6011_),
    .Y(_6012_)
);

INVX1 _12976_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6005_),
    .Y(_6013_)
);

AOI21X1 _12977_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6004_),
    .B(_6002_),
    .C(_5974_),
    .Y(_6014_)
);

OAI21X1 _12978_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6014_),
    .B(_6013_),
    .C(_6012_),
    .Y(_6015_)
);

NAND3X1 _12979_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5962_),
    .B(_6010_),
    .C(_6015_),
    .Y(_6016_)
);

INVX1 _12980_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5962_),
    .Y(_6017_)
);

INVX1 _12981_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6010_),
    .Y(_6018_)
);

AOI21X1 _12982_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6009_),
    .B(_6005_),
    .C(_5964_),
    .Y(_6019_)
);

OAI21X1 _12983_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6019_),
    .B(_6018_),
    .C(_6017_),
    .Y(_6020_)
);

NAND3X1 _12984_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5961_),
    .B(_6016_),
    .C(_6020_),
    .Y(_6021_)
);

INVX1 _12985_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5943_),
    .Y(_6022_)
);

AOI21X1 _12986_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5879_),
    .B(_5944_),
    .C(_6022_),
    .Y(_6023_)
);

OAI21X1 _12987_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6014_),
    .B(_6013_),
    .C(_5964_),
    .Y(_6024_)
);

NAND3X1 _12988_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6005_),
    .B(_6009_),
    .C(_6012_),
    .Y(_6025_)
);

AOI21X1 _12989_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6025_),
    .B(_6024_),
    .C(_6017_),
    .Y(_6026_)
);

AOI21X1 _12990_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6015_),
    .B(_6010_),
    .C(_5962_),
    .Y(_6027_)
);

OAI21X1 _12991_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6026_),
    .B(_6027_),
    .C(_6023_),
    .Y(_6028_)
);

AND2X2 _12992_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6028_),
    .B(_6021_),
    .Y(_6029_)
);

OR2X2 _12993_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5959_),
    .B(_6029_),
    .Y(_6030_)
);

NAND2X1 _12994_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6029_),
    .B(_5959_),
    .Y(_6031_)
);

NAND2X1 _12995_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6031_),
    .B(_6030_),
    .Y(_6375_[9])
);

NAND2X1 _12996_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6021_),
    .B(_6028_),
    .Y(_6032_)
);

NOR2X1 _12997_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5952_),
    .B(_6032_),
    .Y(_6033_)
);

NAND2X1 _12998_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6033_),
    .B(_5876_),
    .Y(_6034_)
);

AOI21X1 _12999_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6020_),
    .B(_6016_),
    .C(_5961_),
    .Y(_6035_)
);

AOI21X1 _13000_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5951_),
    .B(_6021_),
    .C(_6035_),
    .Y(_6036_)
);

INVX1 _13001_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6036_),
    .Y(_6037_)
);

OAI21X1 _13002_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6017_),
    .B(_6019_),
    .C(_6010_),
    .Y(_6038_)
);

OAI21X1 _13003_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5965_),
    .B(_5969_),
    .C(_5967_),
    .Y(_6039_)
);

OAI21X1 _13004_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6006_),
    .B(_6008_),
    .C(_6002_),
    .Y(_6040_)
);

INVX2 _13005_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_6041_)
);

NOR3X1 _13006_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5884_),
    .B(_5711_),
    .C(_5900_),
    .Y(_6042_)
);

OAI22X1 _13007_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5996_),
    .B(_5884_),
    .C(_5604_),
    .D(_5995_),
    .Y(_6043_)
);

INVX1 _13008_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6043_),
    .Y(_6044_)
);

OAI22X1 _13009_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5594_),
    .B(_6041_),
    .C(_6042_),
    .D(_6044_),
    .Y(_6045_)
);

NOR2X1 _13010_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5594_),
    .B(_6041_),
    .Y(_6046_)
);

NAND2X1 _13011_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_5977_),
    .Y(_6047_)
);

NAND3X1 _13012_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6046_),
    .B(_6043_),
    .C(_6047_),
    .Y(_6048_)
);

AND2X2 _13013_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6045_),
    .B(_6048_),
    .Y(_6049_)
);

NOR2X1 _13014_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5985_),
    .B(_5982_),
    .Y(_6050_)
);

OAI21X1 _13015_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5998_),
    .B(_6050_),
    .C(_5986_),
    .Y(_6051_)
);

NAND2X1 _13016_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6] [6]),
    .Y(_6052_)
);

NOR2X1 _13017_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6052_),
    .B(_5995_),
    .Y(_6053_)
);

AND2X2 _13018_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6052_),
    .B(_5995_),
    .Y(_6054_)
);

OAI22X1 _13019_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5910_),
    .B(_5991_),
    .C(_6053_),
    .D(_6054_),
    .Y(_6055_)
);

AND2X2 _13020_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6] [6]),
    .Y(_6056_)
);

AND2X2 _13021_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6]_5_bF$buf1 ),
    .B(gnd),
    .Y(_6057_)
);

NAND2X1 _13022_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6056_),
    .B(_6057_),
    .Y(_6058_)
);

OAI21X1 _13023_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5653_),
    .B(_5898_),
    .C(_6052_),
    .Y(_6059_)
);

AOI21X1 _13024_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[6] [6]),
    .C(_5991_),
    .Y(_6060_)
);

NAND3X1 _13025_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6059_),
    .B(_6060_),
    .C(_6058_),
    .Y(_6061_)
);

AND2X2 _13026_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6055_),
    .B(_6061_),
    .Y(_6062_)
);

NAND2X1 _13027_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6062_),
    .B(_6051_),
    .Y(_6063_)
);

NAND2X1 _13028_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6061_),
    .B(_6055_),
    .Y(_6064_)
);

NAND3X1 _13029_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5986_),
    .B(_6064_),
    .C(_5994_),
    .Y(_6065_)
);

NAND3X1 _13030_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6049_),
    .B(_6065_),
    .C(_6063_),
    .Y(_6066_)
);

NAND2X1 _13031_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6048_),
    .B(_6045_),
    .Y(_6067_)
);

NAND2X1 _13032_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6064_),
    .B(_6051_),
    .Y(_6068_)
);

NAND3X1 _13033_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5986_),
    .B(_6062_),
    .C(_5994_),
    .Y(_6069_)
);

NAND3X1 _13034_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6067_),
    .B(_6069_),
    .C(_6068_),
    .Y(_6070_)
);

NAND3X1 _13035_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6066_),
    .B(_6070_),
    .C(_6040_),
    .Y(_6071_)
);

NAND2X1 _13036_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6070_),
    .B(_6066_),
    .Y(_6072_)
);

NAND3X1 _13037_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6002_),
    .B(_6005_),
    .C(_6072_),
    .Y(_6073_)
);

NAND3X1 _13038_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6039_),
    .B(_6073_),
    .C(_6071_),
    .Y(_6074_)
);

INVX1 _13039_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6039_),
    .Y(_6075_)
);

NAND2X1 _13040_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6072_),
    .B(_6040_),
    .Y(_6076_)
);

AOI21X1 _13041_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5974_),
    .B(_6004_),
    .C(_6007_),
    .Y(_6077_)
);

AND2X2 _13042_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6066_),
    .B(_6070_),
    .Y(_6078_)
);

NAND2X1 _13043_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6077_),
    .B(_6078_),
    .Y(_6079_)
);

NAND3X1 _13044_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6075_),
    .B(_6076_),
    .C(_6079_),
    .Y(_6080_)
);

AOI21X1 _13045_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6074_),
    .B(_6080_),
    .C(_6038_),
    .Y(_6081_)
);

NAND2X1 _13046_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6074_),
    .B(_6080_),
    .Y(_6082_)
);

AOI21X1 _13047_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6010_),
    .B(_6016_),
    .C(_6082_),
    .Y(_6083_)
);

NOR2X1 _13048_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6081_),
    .B(_6083_),
    .Y(_6084_)
);

INVX1 _13049_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6084_),
    .Y(_6085_)
);

AOI21X1 _13050_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6034_),
    .B(_6037_),
    .C(_6085_),
    .Y(_6086_)
);

NAND2X1 _13051_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5956_),
    .B(_6029_),
    .Y(_6087_)
);

OAI21X1 _13052_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6087_),
    .B(_5955_),
    .C(_6037_),
    .Y(_6088_)
);

NOR2X1 _13053_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6084_),
    .B(_6088_),
    .Y(_6089_)
);

NOR2X1 _13054_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6086_),
    .B(_6089_),
    .Y(_6375_[10])
);

NAND3X1 _13055_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6074_),
    .B(_6080_),
    .C(_6038_),
    .Y(_6090_)
);

NAND2X1 _13056_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6084_),
    .B(_6088_),
    .Y(_6091_)
);

NOR2X1 _13057_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6072_),
    .B(_6077_),
    .Y(_6092_)
);

AOI21X1 _13058_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6039_),
    .B(_6073_),
    .C(_6092_),
    .Y(_6093_)
);

NAND2X1 _13059_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6047_),
    .B(_6048_),
    .Y(_6094_)
);

NAND2X1 _13060_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6063_),
    .B(_6066_),
    .Y(_6095_)
);

NOR3X1 _13061_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5884_),
    .B(_6052_),
    .C(_5995_),
    .Y(_6096_)
);

AOI22X1 _13062_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6]_5_bF$buf0 ),
    .B(gnd),
    .C(_6056_),
    .D(_6057_),
    .Y(_6097_)
);

OAI22X1 _13063_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5996_),
    .B(_6041_),
    .C(_6097_),
    .D(_6096_),
    .Y(_6098_)
);

NOR2X1 _13064_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5996_),
    .B(_6041_),
    .Y(_6099_)
);

NAND2X1 _13065_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_6053_),
    .Y(_6100_)
);

OAI21X1 _13066_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5653_),
    .B(_5884_),
    .C(_6058_),
    .Y(_6101_)
);

NAND3X1 _13067_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6099_),
    .B(_6100_),
    .C(_6101_),
    .Y(_6102_)
);

NAND2X1 _13068_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6098_),
    .B(_6102_),
    .Y(_6103_)
);

NAND2X1 _13069_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5910_),
    .B(_5984_),
    .Y(_6104_)
);

NAND2X1 _13070_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[6] [7]),
    .Y(_6105_)
);

OAI22X1 _13071_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5812_),
    .B(_5814_),
    .C(_5898_),
    .D(_5723_),
    .Y(_6106_)
);

OAI21X1 _13072_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6052_),
    .B(_6105_),
    .C(_6106_),
    .Y(_6107_)
);

NAND3X1 _13073_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6104_),
    .B(_6107_),
    .C(_6061_),
    .Y(_6108_)
);

INVX1 _13074_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6108_),
    .Y(_6109_)
);

AOI21X1 _13075_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6061_),
    .B(_6104_),
    .C(_6107_),
    .Y(_6110_)
);

OAI21X1 _13076_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6110_),
    .B(_6109_),
    .C(_6103_),
    .Y(_6111_)
);

AND2X2 _13077_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6102_),
    .B(_6098_),
    .Y(_6112_)
);

INVX1 _13078_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6110_),
    .Y(_6113_)
);

NAND3X1 _13079_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6108_),
    .B(_6113_),
    .C(_6112_),
    .Y(_6114_)
);

AND2X2 _13080_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6114_),
    .B(_6111_),
    .Y(_6115_)
);

NAND2X1 _13081_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6115_),
    .B(_6095_),
    .Y(_6116_)
);

AOI21X1 _13082_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5994_),
    .B(_5986_),
    .C(_6064_),
    .Y(_6117_)
);

AOI21X1 _13083_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6049_),
    .B(_6065_),
    .C(_6117_),
    .Y(_6118_)
);

NAND2X1 _13084_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6111_),
    .B(_6114_),
    .Y(_6119_)
);

NAND2X1 _13085_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6119_),
    .B(_6118_),
    .Y(_6120_)
);

NAND3X1 _13086_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6094_),
    .B(_6120_),
    .C(_6116_),
    .Y(_6121_)
);

INVX1 _13087_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6094_),
    .Y(_6122_)
);

NAND2X1 _13088_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6119_),
    .B(_6095_),
    .Y(_6123_)
);

NAND2X1 _13089_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6118_),
    .B(_6115_),
    .Y(_6124_)
);

NAND3X1 _13090_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6122_),
    .B(_6124_),
    .C(_6123_),
    .Y(_6125_)
);

NAND2X1 _13091_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6121_),
    .B(_6125_),
    .Y(_6126_)
);

NAND2X1 _13092_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6126_),
    .B(_6093_),
    .Y(_6127_)
);

AOI21X1 _13093_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6066_),
    .B(_6070_),
    .C(_6040_),
    .Y(_6128_)
);

OAI21X1 _13094_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6075_),
    .B(_6128_),
    .C(_6071_),
    .Y(_6129_)
);

NAND3X1 _13095_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6121_),
    .B(_6125_),
    .C(_6129_),
    .Y(_6130_)
);

NAND2X1 _13096_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6127_),
    .B(_6130_),
    .Y(_6131_)
);

INVX1 _13097_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6131_),
    .Y(_6132_)
);

NAND3X1 _13098_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6090_),
    .B(_6132_),
    .C(_6091_),
    .Y(_6133_)
);

OAI21X1 _13099_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6083_),
    .B(_6086_),
    .C(_6131_),
    .Y(_6134_)
);

NAND2X1 _13100_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6133_),
    .B(_6134_),
    .Y(_6375_[11])
);

NOR3X1 _13101_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6081_),
    .B(_6083_),
    .C(_6131_),
    .Y(_6135_)
);

NAND3X1 _13102_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6033_),
    .B(_6135_),
    .C(_5876_),
    .Y(_6136_)
);

OAI21X1 _13103_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6090_),
    .B(_6131_),
    .C(_6130_),
    .Y(_6137_)
);

AOI21X1 _13104_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6135_),
    .B(_6036_),
    .C(_6137_),
    .Y(_6138_)
);

AND2X2 _13105_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6121_),
    .B(_6116_),
    .Y(_6139_)
);

OAI21X1 _13106_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5884_),
    .B(_6058_),
    .C(_6102_),
    .Y(_6140_)
);

OAI21X1 _13107_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6109_),
    .B(_6103_),
    .C(_6113_),
    .Y(_6141_)
);

INVX1 _13108_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6141_),
    .Y(_6142_)
);

INVX1 _13109_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6105_),
    .Y(_6143_)
);

NOR2X1 _13110_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5653_),
    .B(_6041_),
    .Y(_6144_)
);

NOR2X1 _13111_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6052_),
    .B(_6105_),
    .Y(_6145_)
);

NOR2X1 _13112_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5723_),
    .B(_5884_),
    .Y(_6146_)
);

NOR2X1 _13113_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6146_),
    .B(_6145_),
    .Y(_6147_)
);

AOI21X1 _13114_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_6145_),
    .C(_6147_),
    .Y(_6148_)
);

OR2X2 _13115_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6148_),
    .B(_6144_),
    .Y(_6149_)
);

NAND2X1 _13116_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6144_),
    .B(_6148_),
    .Y(_6150_)
);

NAND3X1 _13117_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6143_),
    .B(_6150_),
    .C(_6149_),
    .Y(_6151_)
);

NOR2X1 _13118_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6144_),
    .B(_6148_),
    .Y(_6152_)
);

INVX1 _13119_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6150_),
    .Y(_6153_)
);

OAI21X1 _13120_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6152_),
    .B(_6153_),
    .C(_6105_),
    .Y(_6154_)
);

NAND2X1 _13121_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6151_),
    .B(_6154_),
    .Y(_6155_)
);

NAND2X1 _13122_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6142_),
    .B(_6155_),
    .Y(_6156_)
);

NAND3X1 _13123_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6141_),
    .B(_6151_),
    .C(_6154_),
    .Y(_6157_)
);

AOI21X1 _13124_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6156_),
    .B(_6157_),
    .C(_6140_),
    .Y(_6158_)
);

NAND3X1 _13125_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6140_),
    .B(_6157_),
    .C(_6156_),
    .Y(_6159_)
);

INVX1 _13126_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6159_),
    .Y(_6160_)
);

OAI21X1 _13127_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6158_),
    .B(_6160_),
    .C(_6139_),
    .Y(_6161_)
);

OR2X2 _13128_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6160_),
    .B(_6158_),
    .Y(_6162_)
);

OR2X2 _13129_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6162_),
    .B(_6139_),
    .Y(_6163_)
);

NAND2X1 _13130_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6161_),
    .B(_6163_),
    .Y(_6164_)
);

AOI21X1 _13131_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6136_),
    .B(_6138_),
    .C(_6164_),
    .Y(_6165_)
);

NAND3X1 _13132_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5956_),
    .B(_6029_),
    .C(_6135_),
    .Y(_6166_)
);

OAI21X1 _13133_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5955_),
    .B(_6166_),
    .C(_6138_),
    .Y(_6167_)
);

INVX1 _13134_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6164_),
    .Y(_6168_)
);

NOR2X1 _13135_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6168_),
    .B(_6167_),
    .Y(_6169_)
);

NOR2X1 _13136_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6165_),
    .B(_6169_),
    .Y(_6375_[12])
);

NOR2X1 _13137_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6139_),
    .B(_6162_),
    .Y(_6170_)
);

INVX1 _13138_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6145_),
    .Y(_6171_)
);

OAI21X1 _13139_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5884_),
    .B(_6171_),
    .C(_6150_),
    .Y(_6172_)
);

INVX1 _13140_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6172_),
    .Y(_6173_)
);

NOR2X1 _13141_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5814_),
    .B(_6041_),
    .Y(_6174_)
);

NAND2X1 _13142_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6146_),
    .B(_6174_),
    .Y(_6175_)
);

OAI22X1 _13143_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5723_),
    .B(_6041_),
    .C(_5884_),
    .D(_5814_),
    .Y(_6176_)
);

NAND2X1 _13144_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6176_),
    .B(_6175_),
    .Y(_6177_)
);

NAND2X1 _13145_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6177_),
    .B(_6151_),
    .Y(_6178_)
);

OR2X2 _13146_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6151_),
    .B(_6177_),
    .Y(_6179_)
);

NAND2X1 _13147_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6178_),
    .B(_6179_),
    .Y(_6180_)
);

NAND2X1 _13148_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6173_),
    .B(_6180_),
    .Y(_6181_)
);

OR2X2 _13149_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6180_),
    .B(_6173_),
    .Y(_6182_)
);

NAND2X1 _13150_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6181_),
    .B(_6182_),
    .Y(_6183_)
);

NAND3X1 _13151_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6157_),
    .B(_6159_),
    .C(_6183_),
    .Y(_6184_)
);

OAI21X1 _13152_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6142_),
    .B(_6155_),
    .C(_6159_),
    .Y(_6185_)
);

AND2X2 _13153_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6182_),
    .B(_6181_),
    .Y(_6186_)
);

NAND2X1 _13154_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6185_),
    .B(_6186_),
    .Y(_6187_)
);

NAND2X1 _13155_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6184_),
    .B(_6187_),
    .Y(_6188_)
);

OAI21X1 _13156_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6170_),
    .B(_6165_),
    .C(_6188_),
    .Y(_6189_)
);

NAND2X1 _13157_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6168_),
    .B(_6167_),
    .Y(_6190_)
);

AND2X2 _13158_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6187_),
    .B(_6184_),
    .Y(_6191_)
);

NAND3X1 _13159_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6163_),
    .B(_6191_),
    .C(_6190_),
    .Y(_6192_)
);

NAND2X1 _13160_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6192_),
    .B(_6189_),
    .Y(_6375_[13])
);

NAND3X1 _13161_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6161_),
    .B(_6163_),
    .C(_6191_),
    .Y(_6193_)
);

AOI21X1 _13162_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6136_),
    .B(_6138_),
    .C(_6193_),
    .Y(_6194_)
);

OAI21X1 _13163_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6163_),
    .B(_6188_),
    .C(_6187_),
    .Y(_6195_)
);

OAI21X1 _13164_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6173_),
    .B(_6180_),
    .C(_6179_),
    .Y(_6196_)
);

AND2X2 _13165_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6175_),
    .B(_6174_),
    .Y(_6197_)
);

OR2X2 _13166_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6196_),
    .B(_6197_),
    .Y(_6198_)
);

NAND2X1 _13167_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6197_),
    .B(_6196_),
    .Y(_6199_)
);

NAND2X1 _13168_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6199_),
    .B(_6198_),
    .Y(_6200_)
);

OAI21X1 _13169_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6195_),
    .B(_6194_),
    .C(_6200_),
    .Y(_6201_)
);

INVX1 _13170_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6161_),
    .Y(_6202_)
);

NOR3X1 _13171_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6202_),
    .B(_6170_),
    .C(_6188_),
    .Y(_6203_)
);

NAND2X1 _13172_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6203_),
    .B(_6167_),
    .Y(_6204_)
);

INVX1 _13173_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6195_),
    .Y(_6205_)
);

INVX1 _13174_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6200_),
    .Y(_6206_)
);

NAND3X1 _13175_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6205_),
    .B(_6206_),
    .C(_6204_),
    .Y(_6207_)
);

NAND2X1 _13176_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6207_),
    .B(_6201_),
    .Y(_6375_[14])
);

OAI21X1 _13177_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6195_),
    .B(_6194_),
    .C(_6206_),
    .Y(_6208_)
);

OAI21X1 _13178_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6146_),
    .B(_6196_),
    .C(_6174_),
    .Y(_6209_)
);

NAND2X1 _13179_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6209_),
    .B(_6208_),
    .Y(_6375_[15])
);

INVX1 _13180_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_5603_),
    .Y(_6370_[0])
);

AND2X2 _13181_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [0]),
    .B(\u_fir_pe7.mul [0]),
    .Y(_6210_)
);

INVX1 _13182_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [1]),
    .Y(_6211_)
);

INVX1 _13183_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.mul [1]),
    .Y(_6212_)
);

NOR2X1 _13184_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6211_),
    .B(_6212_),
    .Y(_6213_)
);

NOR2X1 _13185_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [1]),
    .B(\u_fir_pe7.mul [1]),
    .Y(_6214_)
);

NOR2X1 _13186_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6214_),
    .B(_6213_),
    .Y(_6215_)
);

NAND2X1 _13187_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6210_),
    .B(_6215_),
    .Y(_6216_)
);

INVX1 _13188_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6216_),
    .Y(_6217_)
);

NOR2X1 _13189_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6210_),
    .B(_6215_),
    .Y(_6218_)
);

NOR2X1 _13190_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6218_),
    .B(_6217_),
    .Y(_6369_[1])
);

OAI21X1 _13191_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6211_),
    .B(_6212_),
    .C(_6216_),
    .Y(_6219_)
);

AND2X2 _13192_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [2]),
    .B(\u_fir_pe7.mul [2]),
    .Y(_6220_)
);

NOR2X1 _13193_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [2]),
    .B(\u_fir_pe7.mul [2]),
    .Y(_6221_)
);

OAI21X1 _13194_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6220_),
    .B(_6221_),
    .C(_6219_),
    .Y(_6222_)
);

INVX1 _13195_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6219_),
    .Y(_6223_)
);

NOR2X1 _13196_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6221_),
    .B(_6220_),
    .Y(_6224_)
);

NAND2X1 _13197_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6224_),
    .B(_6223_),
    .Y(_6225_)
);

NAND2X1 _13198_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6222_),
    .B(_6225_),
    .Y(_6369_[2])
);

AOI21X1 _13199_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6219_),
    .B(_6224_),
    .C(_6220_),
    .Y(_6226_)
);

INVX1 _13200_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [3]),
    .Y(_6227_)
);

INVX1 _13201_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.mul [3]),
    .Y(_6228_)
);

NOR2X1 _13202_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6227_),
    .B(_6228_),
    .Y(_6229_)
);

NOR2X1 _13203_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [3]),
    .B(\u_fir_pe7.mul [3]),
    .Y(_6230_)
);

NOR2X1 _13204_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6230_),
    .B(_6229_),
    .Y(_6231_)
);

NAND2X1 _13205_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6231_),
    .B(_6226_),
    .Y(_6232_)
);

OR2X2 _13206_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6226_),
    .B(_6231_),
    .Y(_6233_)
);

NAND2X1 _13207_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6232_),
    .B(_6233_),
    .Y(_6369_[3])
);

INVX1 _13208_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [4]),
    .Y(_6234_)
);

INVX1 _13209_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.mul [4]),
    .Y(_6235_)
);

NOR2X1 _13210_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6234_),
    .B(_6235_),
    .Y(_6236_)
);

NOR2X1 _13211_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [4]),
    .B(\u_fir_pe7.mul [4]),
    .Y(_6237_)
);

NOR2X1 _13212_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6237_),
    .B(_6236_),
    .Y(_6238_)
);

INVX1 _13213_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6229_),
    .Y(_6239_)
);

OAI21X1 _13214_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6230_),
    .B(_6226_),
    .C(_6239_),
    .Y(_6240_)
);

NAND2X1 _13215_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6238_),
    .B(_6240_),
    .Y(_6241_)
);

OR2X2 _13216_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6240_),
    .B(_6238_),
    .Y(_6242_)
);

AND2X2 _13217_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6242_),
    .B(_6241_),
    .Y(_6369_[4])
);

OAI21X1 _13218_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6234_),
    .B(_6235_),
    .C(_6241_),
    .Y(_6243_)
);

INVX1 _13219_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [5]),
    .Y(_6244_)
);

INVX1 _13220_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.mul [5]),
    .Y(_6245_)
);

NOR2X1 _13221_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6244_),
    .B(_6245_),
    .Y(_6246_)
);

NOR2X1 _13222_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [5]),
    .B(\u_fir_pe7.mul [5]),
    .Y(_6247_)
);

NOR2X1 _13223_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6247_),
    .B(_6246_),
    .Y(_6248_)
);

NAND2X1 _13224_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6248_),
    .B(_6243_),
    .Y(_6249_)
);

OR2X2 _13225_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6243_),
    .B(_6248_),
    .Y(_6250_)
);

AND2X2 _13226_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6250_),
    .B(_6249_),
    .Y(_6369_[5])
);

OAI21X1 _13227_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6244_),
    .B(_6245_),
    .C(_6249_),
    .Y(_6251_)
);

INVX1 _13228_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [6]),
    .Y(_6252_)
);

INVX1 _13229_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.mul [6]),
    .Y(_6253_)
);

NOR2X1 _13230_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6252_),
    .B(_6253_),
    .Y(_6254_)
);

NOR2X1 _13231_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [6]),
    .B(\u_fir_pe7.mul [6]),
    .Y(_6255_)
);

NOR2X1 _13232_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6255_),
    .B(_6254_),
    .Y(_6256_)
);

NAND2X1 _13233_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6256_),
    .B(_6251_),
    .Y(_6257_)
);

OR2X2 _13234_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6251_),
    .B(_6256_),
    .Y(_6258_)
);

AND2X2 _13235_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6258_),
    .B(_6257_),
    .Y(_6369_[6])
);

OAI21X1 _13236_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6252_),
    .B(_6253_),
    .C(_6257_),
    .Y(_6259_)
);

INVX1 _13237_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [7]),
    .Y(_6260_)
);

INVX1 _13238_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.mul [7]),
    .Y(_6261_)
);

NOR2X1 _13239_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6260_),
    .B(_6261_),
    .Y(_6262_)
);

NOR2X1 _13240_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [7]),
    .B(\u_fir_pe7.mul [7]),
    .Y(_6263_)
);

OAI21X1 _13241_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6262_),
    .B(_6263_),
    .C(_6259_),
    .Y(_6264_)
);

INVX1 _13242_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6259_),
    .Y(_6265_)
);

NOR2X1 _13243_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6263_),
    .B(_6262_),
    .Y(_6266_)
);

NAND2X1 _13244_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6266_),
    .B(_6265_),
    .Y(_6267_)
);

NAND2X1 _13245_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6264_),
    .B(_6267_),
    .Y(_6369_[7])
);

INVX1 _13246_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [8]),
    .Y(_6269_)
);

INVX1 _13247_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.mul [8]),
    .Y(_6270_)
);

NOR2X1 _13248_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6269_),
    .B(_6270_),
    .Y(_6271_)
);

NOR2X1 _13249_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [8]),
    .B(\u_fir_pe7.mul [8]),
    .Y(_6272_)
);

NAND2X1 _13250_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6236_),
    .B(_6248_),
    .Y(_6273_)
);

OAI21X1 _13251_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6244_),
    .B(_6245_),
    .C(_6273_),
    .Y(_6274_)
);

NAND2X1 _13252_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6254_),
    .B(_6266_),
    .Y(_6275_)
);

OAI21X1 _13253_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6260_),
    .B(_6261_),
    .C(_6275_),
    .Y(_6276_)
);

AND2X2 _13254_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6256_),
    .B(_6266_),
    .Y(_6277_)
);

AOI21X1 _13255_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6274_),
    .B(_6277_),
    .C(_6276_),
    .Y(_6278_)
);

AND2X2 _13256_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6238_),
    .B(_6248_),
    .Y(_6280_)
);

NAND3X1 _13257_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6280_),
    .B(_6277_),
    .C(_6240_),
    .Y(_6281_)
);

NAND2X1 _13258_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6278_),
    .B(_6281_),
    .Y(_6282_)
);

OAI21X1 _13259_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6271_),
    .B(_6272_),
    .C(_6282_),
    .Y(_6283_)
);

NOR2X1 _13260_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6272_),
    .B(_6271_),
    .Y(_6284_)
);

INVX1 _13261_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6282_),
    .Y(_6285_)
);

NAND2X1 _13262_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6284_),
    .B(_6285_),
    .Y(_6286_)
);

NAND2X1 _13263_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6283_),
    .B(_6286_),
    .Y(_6369_[8])
);

INVX1 _13264_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6271_),
    .Y(_6287_)
);

INVX1 _13265_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6284_),
    .Y(_6288_)
);

OAI21X1 _13266_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6288_),
    .B(_6285_),
    .C(_6287_),
    .Y(_6290_)
);

AND2X2 _13267_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [9]),
    .B(\u_fir_pe7.mul [9]),
    .Y(_6291_)
);

NOR2X1 _13268_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [9]),
    .B(\u_fir_pe7.mul [9]),
    .Y(_6292_)
);

NOR2X1 _13269_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6292_),
    .B(_6291_),
    .Y(_6293_)
);

INVX1 _13270_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6293_),
    .Y(_6294_)
);

OR2X2 _13271_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6290_),
    .B(_6294_),
    .Y(_6295_)
);

OAI21X1 _13272_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6291_),
    .B(_6292_),
    .C(_6290_),
    .Y(_6296_)
);

NAND2X1 _13273_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6296_),
    .B(_6295_),
    .Y(_6369_[9])
);

NOR2X1 _13274_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6294_),
    .B(_6288_),
    .Y(_6297_)
);

AOI21X1 _13275_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6293_),
    .B(_6271_),
    .C(_6291_),
    .Y(_6298_)
);

INVX1 _13276_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6298_),
    .Y(_6300_)
);

AOI21X1 _13277_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6282_),
    .B(_6297_),
    .C(_6300_),
    .Y(_6301_)
);

INVX1 _13278_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6301_),
    .Y(_6302_)
);

INVX1 _13279_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [10]),
    .Y(_6303_)
);

INVX1 _13280_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.mul [10]),
    .Y(_6304_)
);

NOR2X1 _13281_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6303_),
    .B(_6304_),
    .Y(_6305_)
);

NOR2X1 _13282_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [10]),
    .B(\u_fir_pe7.mul [10]),
    .Y(_6306_)
);

NOR2X1 _13283_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6306_),
    .B(_6305_),
    .Y(_6307_)
);

NAND2X1 _13284_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6307_),
    .B(_6302_),
    .Y(_6308_)
);

OAI21X1 _13285_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6305_),
    .B(_6306_),
    .C(_6301_),
    .Y(_6309_)
);

AND2X2 _13286_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6308_),
    .B(_6309_),
    .Y(_6369_[10])
);

OAI21X1 _13287_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6303_),
    .B(_6304_),
    .C(_6308_),
    .Y(_6311_)
);

AND2X2 _13288_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [11]),
    .B(\u_fir_pe7.mul [11]),
    .Y(_6312_)
);

NOR2X1 _13289_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [11]),
    .B(\u_fir_pe7.mul [11]),
    .Y(_6313_)
);

NOR2X1 _13290_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6313_),
    .B(_6312_),
    .Y(_6314_)
);

NOR2X1 _13291_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6314_),
    .B(_6311_),
    .Y(_6315_)
);

AND2X2 _13292_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6311_),
    .B(_6314_),
    .Y(_6316_)
);

NOR2X1 _13293_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6315_),
    .B(_6316_),
    .Y(_6369_[11])
);

AOI21X1 _13294_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6314_),
    .B(_6305_),
    .C(_6312_),
    .Y(_6317_)
);

NAND2X1 _13295_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6314_),
    .B(_6307_),
    .Y(_6318_)
);

OAI21X1 _13296_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6318_),
    .B(_6301_),
    .C(_6317_),
    .Y(_6320_)
);

INVX1 _13297_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [12]),
    .Y(_6321_)
);

INVX1 _13298_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.mul [12]),
    .Y(_6322_)
);

NOR2X1 _13299_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6321_),
    .B(_6322_),
    .Y(_6323_)
);

NOR2X1 _13300_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [12]),
    .B(\u_fir_pe7.mul [12]),
    .Y(_6324_)
);

NOR2X1 _13301_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6324_),
    .B(_6323_),
    .Y(_6325_)
);

NAND2X1 _13302_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6325_),
    .B(_6320_),
    .Y(_6326_)
);

OR2X2 _13303_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6320_),
    .B(_6325_),
    .Y(_6327_)
);

AND2X2 _13304_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6327_),
    .B(_6326_),
    .Y(_6369_[12])
);

OAI21X1 _13305_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6321_),
    .B(_6322_),
    .C(_6326_),
    .Y(_6328_)
);

INVX1 _13306_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [13]),
    .Y(_6330_)
);

INVX1 _13307_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.mul [13]),
    .Y(_6331_)
);

NOR2X1 _13308_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6330_),
    .B(_6331_),
    .Y(_6332_)
);

NOR2X1 _13309_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [13]),
    .B(\u_fir_pe7.mul [13]),
    .Y(_6333_)
);

NOR2X1 _13310_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6333_),
    .B(_6332_),
    .Y(_6334_)
);

NAND2X1 _13311_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6334_),
    .B(_6328_),
    .Y(_6335_)
);

OR2X2 _13312_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6328_),
    .B(_6334_),
    .Y(_6336_)
);

AND2X2 _13313_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6336_),
    .B(_6335_),
    .Y(_6369_[13])
);

OAI21X1 _13314_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6330_),
    .B(_6331_),
    .C(_6335_),
    .Y(_6337_)
);

INVX1 _13315_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [14]),
    .Y(_6338_)
);

INVX1 _13316_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.mul [14]),
    .Y(_6340_)
);

NOR2X1 _13317_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6338_),
    .B(_6340_),
    .Y(_6341_)
);

NOR2X1 _13318_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [14]),
    .B(\u_fir_pe7.mul [14]),
    .Y(_6342_)
);

NOR2X1 _13319_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6342_),
    .B(_6341_),
    .Y(_6343_)
);

AND2X2 _13320_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6337_),
    .B(_6343_),
    .Y(_6344_)
);

NOR2X1 _13321_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6343_),
    .B(_6337_),
    .Y(_6345_)
);

NOR2X1 _13322_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6345_),
    .B(_6344_),
    .Y(_6369_[14])
);

INVX1 _13323_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6341_),
    .Y(_6346_)
);

NAND2X1 _13324_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6343_),
    .B(_6337_),
    .Y(_6347_)
);

NAND2X1 _13325_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [15]),
    .B(\u_fir_pe7.mul [15]),
    .Y(_6348_)
);

OR2X2 _13326_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [15]),
    .B(\u_fir_pe7.mul [15]),
    .Y(_6350_)
);

NAND2X1 _13327_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6348_),
    .B(_6350_),
    .Y(_6351_)
);

INVX1 _13328_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6351_),
    .Y(_6352_)
);

NAND3X1 _13329_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6346_),
    .B(_6352_),
    .C(_6347_),
    .Y(_6353_)
);

OAI21X1 _13330_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6341_),
    .B(_6344_),
    .C(_6351_),
    .Y(_6354_)
);

NAND2X1 _13331_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6353_),
    .B(_6354_),
    .Y(_6369_[15])
);

NOR2X1 _13332_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe7.rYin [0]),
    .B(\u_fir_pe7.mul [0]),
    .Y(_6355_)
);

NOR2X1 _13333_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6355_),
    .B(_6210_),
    .Y(_6368_[0])
);

AOI21X1 _13334_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[6] [0]),
    .B(gnd),
    .C(_6279_),
    .Y(_6356_)
);

NOR2X1 _13335_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6356_),
    .B(_6299_),
    .Y(_6371_[1])
);

NOR2X1 _13336_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6299_),
    .B(_6363_),
    .Y(_6358_)
);

NOR2X1 _13337_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6358_),
    .B(_6365_),
    .Y(_6372_[2])
);

DFFPOSX1 _13338_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_6368_[0]),
    .Q(\Y[7] [0])
);

DFFPOSX1 _13339_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_6369_[1]),
    .Q(\Y[7] [1])
);

DFFPOSX1 _13340_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_6369_[2]),
    .Q(\Y[7] [2])
);

DFFPOSX1 _13341_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_6369_[3]),
    .Q(\Y[7] [3])
);

DFFPOSX1 _13342_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_6369_[4]),
    .Q(\Y[7] [4])
);

DFFPOSX1 _13343_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_6369_[5]),
    .Q(\Y[7] [5])
);

DFFPOSX1 _13344_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf57),
    .D(_6369_[6]),
    .Q(\Y[7] [6])
);

DFFPOSX1 _13345_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf56),
    .D(_6369_[7]),
    .Q(\Y[7] [7])
);

DFFPOSX1 _13346_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf55),
    .D(_6369_[8]),
    .Q(\Y[7] [8])
);

DFFPOSX1 _13347_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf54),
    .D(_6369_[9]),
    .Q(\Y[7] [9])
);

DFFPOSX1 _13348_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf53),
    .D(_6369_[10]),
    .Q(\Y[7] [10])
);

DFFPOSX1 _13349_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf52),
    .D(_6369_[11]),
    .Q(\Y[7] [11])
);

DFFPOSX1 _13350_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf51),
    .D(_6369_[12]),
    .Q(\Y[7] [12])
);

DFFPOSX1 _13351_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf50),
    .D(_6369_[13]),
    .Q(\Y[7] [13])
);

DFFPOSX1 _13352_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf49),
    .D(_6369_[14]),
    .Q(\Y[7] [14])
);

DFFPOSX1 _13353_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf48),
    .D(_6369_[15]),
    .Q(\Y[7] [15])
);

DFFPOSX1 _13354_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf47),
    .D(\X[6] [0]),
    .Q(\X[7] [0])
);

DFFPOSX1 _13355_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf46),
    .D(\X[6] [1]),
    .Q(\X[7] [1])
);

DFFPOSX1 _13356_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf45),
    .D(\X[6] [2]),
    .Q(\X[7] [2])
);

DFFPOSX1 _13357_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf44),
    .D(\X[6] [3]),
    .Q(\X[7] [3])
);

DFFPOSX1 _13358_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf43),
    .D(\X[6] [4]),
    .Q(\X[7] [4])
);

DFFPOSX1 _13359_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf42),
    .D(\X[6]_5_bF$buf3 ),
    .Q(\X[7] [5])
);

DFFPOSX1 _13360_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf41),
    .D(\X[6] [6]),
    .Q(\X[7] [6])
);

DFFPOSX1 _13361_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf40),
    .D(\X[6] [7]),
    .Q(\X[7] [7])
);

DFFPOSX1 _13362_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf39),
    .D(\Y[6] [0]),
    .Q(\u_fir_pe7.rYin [0])
);

DFFPOSX1 _13363_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf38),
    .D(\Y[6] [1]),
    .Q(\u_fir_pe7.rYin [1])
);

DFFPOSX1 _13364_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf37),
    .D(\Y[6] [2]),
    .Q(\u_fir_pe7.rYin [2])
);

DFFPOSX1 _13365_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf36),
    .D(\Y[6] [3]),
    .Q(\u_fir_pe7.rYin [3])
);

DFFPOSX1 _13366_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf35),
    .D(\Y[6] [4]),
    .Q(\u_fir_pe7.rYin [4])
);

DFFPOSX1 _13367_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf34),
    .D(\Y[6] [5]),
    .Q(\u_fir_pe7.rYin [5])
);

DFFPOSX1 _13368_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf33),
    .D(\Y[6] [6]),
    .Q(\u_fir_pe7.rYin [6])
);

DFFPOSX1 _13369_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf32),
    .D(\Y[6] [7]),
    .Q(\u_fir_pe7.rYin [7])
);

DFFPOSX1 _13370_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf31),
    .D(\Y[6] [8]),
    .Q(\u_fir_pe7.rYin [8])
);

DFFPOSX1 _13371_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf30),
    .D(\Y[6] [9]),
    .Q(\u_fir_pe7.rYin [9])
);

DFFPOSX1 _13372_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf29),
    .D(\Y[6] [10]),
    .Q(\u_fir_pe7.rYin [10])
);

DFFPOSX1 _13373_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf28),
    .D(\Y[6] [11]),
    .Q(\u_fir_pe7.rYin [11])
);

DFFPOSX1 _13374_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf27),
    .D(\Y[6] [12]),
    .Q(\u_fir_pe7.rYin [12])
);

DFFPOSX1 _13375_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf26),
    .D(\Y[6] [13]),
    .Q(\u_fir_pe7.rYin [13])
);

DFFPOSX1 _13376_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf25),
    .D(\Y[6] [14]),
    .Q(\u_fir_pe7.rYin [14])
);

DFFPOSX1 _13377_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf24),
    .D(\Y[6] [15]),
    .Q(\u_fir_pe7.rYin [15])
);

DFFPOSX1 _13378_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf23),
    .D(_6370_[0]),
    .Q(\u_fir_pe7.mul [0])
);

DFFPOSX1 _13379_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf22),
    .D(_6371_[1]),
    .Q(\u_fir_pe7.mul [1])
);

DFFPOSX1 _13380_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf21),
    .D(_6372_[2]),
    .Q(\u_fir_pe7.mul [2])
);

DFFPOSX1 _13381_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf20),
    .D(_6373_[3]),
    .Q(\u_fir_pe7.mul [3])
);

DFFPOSX1 _13382_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf19),
    .D(_6374_[4]),
    .Q(\u_fir_pe7.mul [4])
);

DFFPOSX1 _13383_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf18),
    .D(_6375_[5]),
    .Q(\u_fir_pe7.mul [5])
);

DFFPOSX1 _13384_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf17),
    .D(_6375_[6]),
    .Q(\u_fir_pe7.mul [6])
);

DFFPOSX1 _13385_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf16),
    .D(_6375_[7]),
    .Q(\u_fir_pe7.mul [7])
);

DFFPOSX1 _13386_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf15),
    .D(_6375_[8]),
    .Q(\u_fir_pe7.mul [8])
);

DFFPOSX1 _13387_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf14),
    .D(_6375_[9]),
    .Q(\u_fir_pe7.mul [9])
);

DFFPOSX1 _13388_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf13),
    .D(_6375_[10]),
    .Q(\u_fir_pe7.mul [10])
);

DFFPOSX1 _13389_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf12),
    .D(_6375_[11]),
    .Q(\u_fir_pe7.mul [11])
);

DFFPOSX1 _13390_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf11),
    .D(_6375_[12]),
    .Q(\u_fir_pe7.mul [12])
);

DFFPOSX1 _13391_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf10),
    .D(_6375_[13]),
    .Q(\u_fir_pe7.mul [13])
);

DFFPOSX1 _13392_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf9),
    .D(_6375_[14]),
    .Q(\u_fir_pe7.mul [14])
);

DFFPOSX1 _13393_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf8),
    .D(_6375_[15]),
    .Q(\u_fir_pe7.mul [15])
);

BUFX2 _13394_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6376_[0]),
    .Y(Xout[0])
);

BUFX2 _13395_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6376_[1]),
    .Y(Xout[1])
);

BUFX2 _13396_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6376_[2]),
    .Y(Xout[2])
);

BUFX2 _13397_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6376_[3]),
    .Y(Xout[3])
);

BUFX2 _13398_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6376_[4]),
    .Y(Xout[4])
);

BUFX2 _13399_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6376_[5]),
    .Y(Xout[5])
);

BUFX2 _13400_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6376_[6]),
    .Y(Xout[6])
);

BUFX2 _13401_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6376_[7]),
    .Y(Xout[7])
);

BUFX2 _13402_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6377_[0]),
    .Y(Yout[0])
);

BUFX2 _13403_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6377_[1]),
    .Y(Yout[1])
);

BUFX2 _13404_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6377_[10]),
    .Y(Yout[10])
);

BUFX2 _13405_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6377_[11]),
    .Y(Yout[11])
);

BUFX2 _13406_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6377_[12]),
    .Y(Yout[12])
);

BUFX2 _13407_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6377_[13]),
    .Y(Yout[13])
);

BUFX2 _13408_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6377_[14]),
    .Y(Yout[14])
);

BUFX2 _13409_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6377_[15]),
    .Y(Yout[15])
);

BUFX2 _13410_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6377_[2]),
    .Y(Yout[2])
);

BUFX2 _13411_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6377_[3]),
    .Y(Yout[3])
);

BUFX2 _13412_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6377_[4]),
    .Y(Yout[4])
);

BUFX2 _13413_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6377_[5]),
    .Y(Yout[5])
);

BUFX2 _13414_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6377_[6]),
    .Y(Yout[6])
);

BUFX2 _13415_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6377_[7]),
    .Y(Yout[7])
);

BUFX2 _13416_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6377_[8]),
    .Y(Yout[8])
);

BUFX2 _13417_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_6377_[9]),
    .Y(Yout[9])
);

NAND2X1 _6378_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[0]),
    .B(gnd),
    .Y(_689_)
);

AND2X2 _6379_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[1]),
    .B(gnd),
    .Y(_700_)
);

INVX1 _6380_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_700_),
    .Y(_710_)
);

NOR2X1 _6381_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_689_),
    .B(_710_),
    .Y(_720_)
);

NAND2X1 _6382_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(Xin[1]),
    .Y(_731_)
);

NOR2X1 _6383_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_689_),
    .B(_731_),
    .Y(_740_)
);

AOI22X1 _6384_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[0]),
    .B(vdd),
    .C(Xin[1]),
    .D(gnd),
    .Y(_750_)
);

NOR2X1 _6385_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_750_),
    .B(_740_),
    .Y(_760_)
);

INVX1 _6386_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[2]),
    .Y(_770_)
);

INVX2 _6387_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_778_)
);

NOR2X1 _6388_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_770_),
    .B(_778_),
    .Y(_780_)
);

NAND2X1 _6389_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_780_),
    .B(_760_),
    .Y(_781_)
);

INVX1 _6390_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_781_),
    .Y(_782_)
);

NOR2X1 _6391_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_780_),
    .B(_760_),
    .Y(_783_)
);

NOR2X1 _6392_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_783_),
    .B(_782_),
    .Y(_784_)
);

NAND2X1 _6393_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720_),
    .B(_784_),
    .Y(_785_)
);

INVX1 _6394_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_785_),
    .Y(_786_)
);

NAND2X1 _6395_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[3]),
    .Y(_787_)
);

INVX1 _6396_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_787_),
    .Y(_788_)
);

NAND2X1 _6397_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[2]),
    .Y(_0_)
);

INVX1 _6398_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_0_),
    .Y(_1_)
);

NAND2X1 _6399_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[0]),
    .Y(_2_)
);

OR2X2 _6400_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_731_),
    .B(_2_),
    .Y(_3_)
);

AOI22X1 _6401_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[0]),
    .C(vdd),
    .D(Xin[1]),
    .Y(_4_)
);

INVX1 _6402_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4_),
    .Y(_5_)
);

NAND3X1 _6403_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1_),
    .B(_5_),
    .C(_3_),
    .Y(_6_)
);

NOR2X1 _6404_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_731_),
    .B(_2_),
    .Y(_7_)
);

OAI21X1 _6405_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4_),
    .B(_7_),
    .C(_0_),
    .Y(_8_)
);

NAND3X1 _6406_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_740_),
    .B(_8_),
    .C(_6_),
    .Y(_9_)
);

INVX1 _6407_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_740_),
    .Y(_10_)
);

NAND3X1 _6408_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_0_),
    .B(_5_),
    .C(_3_),
    .Y(_11_)
);

OAI21X1 _6409_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_4_),
    .B(_7_),
    .C(_1_),
    .Y(_12_)
);

NAND3X1 _6410_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_10_),
    .B(_12_),
    .C(_11_),
    .Y(_13_)
);

NAND3X1 _6411_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_788_),
    .B(_13_),
    .C(_9_),
    .Y(_14_)
);

INVX2 _6412_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[3]),
    .Y(_15_)
);

NAND2X1 _6413_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_13_),
    .B(_9_),
    .Y(_16_)
);

OAI21X1 _6414_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_778_),
    .B(_15_),
    .C(_16_),
    .Y(_17_)
);

NAND2X1 _6415_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_14_),
    .B(_17_),
    .Y(_18_)
);

NAND2X1 _6416_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_781_),
    .B(_18_),
    .Y(_19_)
);

NAND3X1 _6417_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_782_),
    .B(_14_),
    .C(_17_),
    .Y(_20_)
);

NAND3X1 _6418_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_20_),
    .B(_786_),
    .C(_19_),
    .Y(_21_)
);

INVX1 _6419_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_21_),
    .Y(_22_)
);

AOI21X1 _6420_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_19_),
    .B(_20_),
    .C(_786_),
    .Y(_23_)
);

NOR2X1 _6421_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_23_),
    .B(_22_),
    .Y(_794_[3])
);

NAND2X1 _6422_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[0]),
    .B(gnd),
    .Y(_24_)
);

NAND2X1 _6423_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[4]),
    .B(gnd),
    .Y(_25_)
);

NOR2X1 _6424_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_24_),
    .B(_25_),
    .Y(_26_)
);

AOI22X1 _6425_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[0]),
    .B(gnd),
    .C(gnd),
    .D(Xin[4]),
    .Y(_27_)
);

NOR2X1 _6426_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_27_),
    .B(_26_),
    .Y(_28_)
);

INVX1 _6427_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_28_),
    .Y(_29_)
);

NAND2X1 _6428_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[0]),
    .B(vdd),
    .Y(_30_)
);

NAND2X1 _6429_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[1]),
    .Y(_31_)
);

OAI22X1 _6430_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_30_),
    .B(_31_),
    .C(_0_),
    .D(_4_),
    .Y(_32_)
);

NAND2X1 _6431_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[3]),
    .Y(_33_)
);

INVX1 _6432_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_33_),
    .Y(_34_)
);

AND2X2 _6433_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(Xin[1]),
    .Y(_35_)
);

AND2X2 _6434_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[2]),
    .Y(_36_)
);

NAND2X1 _6435_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_35_),
    .B(_36_),
    .Y(_37_)
);

AOI22X1 _6436_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[1]),
    .C(vdd),
    .D(Xin[2]),
    .Y(_38_)
);

INVX1 _6437_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_38_),
    .Y(_39_)
);

NAND3X1 _6438_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_34_),
    .B(_39_),
    .C(_37_),
    .Y(_40_)
);

NAND3X1 _6439_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(Xin[2]),
    .C(_31_),
    .Y(_41_)
);

NAND2X1 _6440_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(Xin[2]),
    .Y(_42_)
);

NAND3X1 _6441_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[1]),
    .C(_42_),
    .Y(_43_)
);

NAND3X1 _6442_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_33_),
    .B(_41_),
    .C(_43_),
    .Y(_44_)
);

NAND3X1 _6443_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_32_),
    .B(_44_),
    .C(_40_),
    .Y(_45_)
);

INVX1 _6444_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_32_),
    .Y(_46_)
);

NAND2X1 _6445_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_44_),
    .B(_40_),
    .Y(_47_)
);

NAND2X1 _6446_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_46_),
    .B(_47_),
    .Y(_48_)
);

NAND3X1 _6447_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_29_),
    .B(_45_),
    .C(_48_),
    .Y(_49_)
);

NAND2X1 _6448_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_32_),
    .B(_47_),
    .Y(_50_)
);

NAND3X1 _6449_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_40_),
    .B(_44_),
    .C(_46_),
    .Y(_51_)
);

NAND3X1 _6450_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_28_),
    .B(_51_),
    .C(_50_),
    .Y(_52_)
);

AOI22X1 _6451_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_9_),
    .B(_14_),
    .C(_49_),
    .D(_52_),
    .Y(_53_)
);

INVX1 _6452_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_53_),
    .Y(_54_)
);

NAND2X1 _6453_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_9_),
    .B(_14_),
    .Y(_55_)
);

NAND2X1 _6454_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_49_),
    .B(_52_),
    .Y(_56_)
);

OR2X2 _6455_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_56_),
    .B(_55_),
    .Y(_57_)
);

NAND2X1 _6456_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_54_),
    .B(_57_),
    .Y(_58_)
);

OAI21X1 _6457_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_781_),
    .B(_18_),
    .C(_21_),
    .Y(_59_)
);

OR2X2 _6458_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_59_),
    .B(_58_),
    .Y(_60_)
);

NAND3X1 _6459_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_28_),
    .B(_45_),
    .C(_48_),
    .Y(_61_)
);

INVX1 _6460_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_45_),
    .Y(_62_)
);

AOI21X1 _6461_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_40_),
    .B(_44_),
    .C(_32_),
    .Y(_63_)
);

OAI21X1 _6462_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_63_),
    .B(_62_),
    .C(_29_),
    .Y(_64_)
);

AOI21X1 _6463_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_61_),
    .B(_64_),
    .C(_55_),
    .Y(_65_)
);

OAI21X1 _6464_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_53_),
    .B(_65_),
    .C(_59_),
    .Y(_66_)
);

NAND2X1 _6465_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_66_),
    .B(_60_),
    .Y(_795_[4])
);

NOR2X1 _6466_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_21_),
    .B(_58_),
    .Y(_67_)
);

NOR3X1 _6467_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_53_),
    .B(_20_),
    .C(_65_),
    .Y(_68_)
);

OAI21X1 _6468_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_29_),
    .B(_63_),
    .C(_45_),
    .Y(_69_)
);

NAND2X1 _6469_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[0]),
    .B(gnd),
    .Y(_70_)
);

INVX1 _6470_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_70_),
    .Y(_71_)
);

AND2X2 _6471_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin_5_bF$buf3),
    .Y(_72_)
);

NAND2X1 _6472_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_700_),
    .B(_72_),
    .Y(_73_)
);

INVX2 _6473_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin_5_bF$buf2),
    .Y(_74_)
);

NAND2X1 _6474_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[1]),
    .B(gnd),
    .Y(_75_)
);

OAI21X1 _6475_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_778_),
    .B(_74_),
    .C(_75_),
    .Y(_76_)
);

NAND3X1 _6476_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_76_),
    .B(_71_),
    .C(_73_),
    .Y(_77_)
);

NAND3X1 _6477_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin_5_bF$buf1),
    .C(_75_),
    .Y(_78_)
);

NAND2X1 _6478_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin_5_bF$buf0),
    .Y(_79_)
);

NAND3X1 _6479_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[1]),
    .B(gnd),
    .C(_79_),
    .Y(_80_)
);

NAND3X1 _6480_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_70_),
    .B(_78_),
    .C(_80_),
    .Y(_81_)
);

AND2X2 _6481_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_77_),
    .B(_81_),
    .Y(_82_)
);

NAND2X1 _6482_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[2]),
    .Y(_83_)
);

OAI22X1 _6483_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_731_),
    .B(_83_),
    .C(_33_),
    .D(_38_),
    .Y(_84_)
);

NAND2X1 _6484_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[4]),
    .Y(_85_)
);

INVX1 _6485_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_85_),
    .Y(_86_)
);

AND2X2 _6486_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(Xin[3]),
    .Y(_87_)
);

NAND2X1 _6487_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_36_),
    .B(_87_),
    .Y(_88_)
);

INVX1 _6488_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .Y(_89_)
);

OAI21X1 _6489_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_89_),
    .B(_15_),
    .C(_83_),
    .Y(_90_)
);

NAND3X1 _6490_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_86_),
    .B(_90_),
    .C(_88_),
    .Y(_91_)
);

NAND3X1 _6491_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(Xin[3]),
    .C(_83_),
    .Y(_92_)
);

NAND2X1 _6492_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(Xin[3]),
    .Y(_93_)
);

NAND3X1 _6493_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[2]),
    .C(_93_),
    .Y(_94_)
);

NAND3X1 _6494_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_85_),
    .B(_92_),
    .C(_94_),
    .Y(_95_)
);

NAND3X1 _6495_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_84_),
    .B(_95_),
    .C(_91_),
    .Y(_96_)
);

INVX1 _6496_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_84_),
    .Y(_97_)
);

AOI21X1 _6497_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_92_),
    .B(_94_),
    .C(_85_),
    .Y(_98_)
);

AOI22X1 _6498_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[4]),
    .C(_88_),
    .D(_90_),
    .Y(_99_)
);

OAI21X1 _6499_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_98_),
    .B(_99_),
    .C(_97_),
    .Y(_100_)
);

NAND3X1 _6500_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_96_),
    .B(_82_),
    .C(_100_),
    .Y(_101_)
);

NAND2X1 _6501_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_81_),
    .B(_77_),
    .Y(_102_)
);

OAI21X1 _6502_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_98_),
    .B(_99_),
    .C(_84_),
    .Y(_103_)
);

NAND3X1 _6503_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_95_),
    .B(_91_),
    .C(_97_),
    .Y(_104_)
);

NAND3X1 _6504_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_102_),
    .B(_104_),
    .C(_103_),
    .Y(_105_)
);

NAND3X1 _6505_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_101_),
    .B(_105_),
    .C(_69_),
    .Y(_106_)
);

AOI21X1 _6506_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_28_),
    .B(_48_),
    .C(_62_),
    .Y(_107_)
);

AOI21X1 _6507_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_103_),
    .B(_104_),
    .C(_102_),
    .Y(_108_)
);

AOI21X1 _6508_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_100_),
    .B(_96_),
    .C(_82_),
    .Y(_109_)
);

OAI21X1 _6509_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_108_),
    .B(_109_),
    .C(_107_),
    .Y(_110_)
);

NAND3X1 _6510_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_26_),
    .B(_106_),
    .C(_110_),
    .Y(_111_)
);

INVX1 _6511_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_26_),
    .Y(_112_)
);

OAI21X1 _6512_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_108_),
    .B(_109_),
    .C(_69_),
    .Y(_113_)
);

NAND3X1 _6513_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_101_),
    .B(_105_),
    .C(_107_),
    .Y(_114_)
);

NAND3X1 _6514_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_112_),
    .B(_113_),
    .C(_114_),
    .Y(_115_)
);

NAND3X1 _6515_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_53_),
    .B(_111_),
    .C(_115_),
    .Y(_116_)
);

NAND3X1 _6516_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_112_),
    .B(_106_),
    .C(_110_),
    .Y(_117_)
);

NAND3X1 _6517_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_26_),
    .B(_113_),
    .C(_114_),
    .Y(_118_)
);

NAND3X1 _6518_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_54_),
    .B(_117_),
    .C(_118_),
    .Y(_119_)
);

NAND3X1 _6519_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_116_),
    .B(_119_),
    .C(_68_),
    .Y(_120_)
);

INVX1 _6520_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_20_),
    .Y(_121_)
);

NAND3X1 _6521_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_121_),
    .B(_54_),
    .C(_57_),
    .Y(_122_)
);

NAND3X1 _6522_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_54_),
    .B(_111_),
    .C(_115_),
    .Y(_123_)
);

NAND3X1 _6523_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_53_),
    .B(_117_),
    .C(_118_),
    .Y(_124_)
);

NAND3X1 _6524_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_123_),
    .B(_124_),
    .C(_122_),
    .Y(_125_)
);

NAND3X1 _6525_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_120_),
    .B(_125_),
    .C(_67_),
    .Y(_126_)
);

INVX1 _6526_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_67_),
    .Y(_127_)
);

INVX1 _6527_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_120_),
    .Y(_128_)
);

INVX1 _6528_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_125_),
    .Y(_129_)
);

OAI21X1 _6529_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_128_),
    .B(_129_),
    .C(_127_),
    .Y(_130_)
);

AND2X2 _6530_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_130_),
    .B(_126_),
    .Y(_796_[5])
);

AND2X2 _6531_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[0]),
    .B(gnd),
    .Y(_131_)
);

NAND2X1 _6532_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin_5_bF$buf3),
    .Y(_132_)
);

OAI21X1 _6533_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_710_),
    .B(_132_),
    .C(_77_),
    .Y(_133_)
);

OR2X2 _6534_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_133_),
    .B(_131_),
    .Y(_134_)
);

NAND2X1 _6535_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_131_),
    .B(_133_),
    .Y(_135_)
);

NAND2X1 _6536_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_135_),
    .B(_134_),
    .Y(_136_)
);

AOI21X1 _6537_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_91_),
    .B(_95_),
    .C(_84_),
    .Y(_137_)
);

OAI21X1 _6538_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_102_),
    .B(_137_),
    .C(_96_),
    .Y(_138_)
);

NAND2X1 _6539_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[1]),
    .B(gnd),
    .Y(_139_)
);

INVX1 _6540_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_139_),
    .Y(_140_)
);

AND2X2 _6541_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[2]),
    .B(gnd),
    .Y(_141_)
);

AND2X2 _6542_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[6]),
    .Y(_142_)
);

NAND2X1 _6543_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_141_),
    .B(_142_),
    .Y(_143_)
);

INVX2 _6544_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[6]),
    .Y(_144_)
);

NAND2X1 _6545_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[2]),
    .B(gnd),
    .Y(_145_)
);

OAI21X1 _6546_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_778_),
    .B(_144_),
    .C(_145_),
    .Y(_146_)
);

NAND3X1 _6547_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_146_),
    .B(_140_),
    .C(_143_),
    .Y(_147_)
);

NAND3X1 _6548_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[6]),
    .C(_145_),
    .Y(_148_)
);

NAND2X1 _6549_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[6]),
    .Y(_149_)
);

NAND2X1 _6550_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_149_),
    .B(_141_),
    .Y(_150_)
);

NAND3X1 _6551_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_139_),
    .B(_148_),
    .C(_150_),
    .Y(_151_)
);

AND2X2 _6552_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_147_),
    .B(_151_),
    .Y(_152_)
);

NAND2X1 _6553_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[3]),
    .Y(_153_)
);

AOI22X1 _6554_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[2]),
    .C(vdd),
    .D(Xin[3]),
    .Y(_154_)
);

OAI22X1 _6555_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_42_),
    .B(_153_),
    .C(_85_),
    .D(_154_),
    .Y(_155_)
);

NAND2X1 _6556_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin_5_bF$buf2),
    .Y(_156_)
);

INVX1 _6557_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_156_),
    .Y(_157_)
);

AND2X2 _6558_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[4]),
    .Y(_158_)
);

NAND2X1 _6559_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_87_),
    .B(_158_),
    .Y(_159_)
);

AOI22X1 _6560_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[3]),
    .C(vdd),
    .D(Xin[4]),
    .Y(_160_)
);

INVX1 _6561_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_160_),
    .Y(_161_)
);

NAND3X1 _6562_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_157_),
    .B(_161_),
    .C(_159_),
    .Y(_162_)
);

NAND3X1 _6563_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(Xin[4]),
    .C(_153_),
    .Y(_163_)
);

NAND2X1 _6564_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(Xin[4]),
    .Y(_164_)
);

NAND3X1 _6565_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[3]),
    .C(_164_),
    .Y(_165_)
);

NAND3X1 _6566_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_156_),
    .B(_163_),
    .C(_165_),
    .Y(_166_)
);

NAND3X1 _6567_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_155_),
    .B(_166_),
    .C(_162_),
    .Y(_167_)
);

INVX1 _6568_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_155_),
    .Y(_168_)
);

AOI21X1 _6569_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_163_),
    .B(_165_),
    .C(_156_),
    .Y(_169_)
);

AOI22X1 _6570_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin_5_bF$buf1),
    .C(_159_),
    .D(_161_),
    .Y(_170_)
);

OAI21X1 _6571_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_169_),
    .B(_170_),
    .C(_168_),
    .Y(_171_)
);

NAND3X1 _6572_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_167_),
    .B(_152_),
    .C(_171_),
    .Y(_172_)
);

NAND2X1 _6573_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_151_),
    .B(_147_),
    .Y(_173_)
);

OAI21X1 _6574_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_169_),
    .B(_170_),
    .C(_155_),
    .Y(_174_)
);

NAND3X1 _6575_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_162_),
    .B(_166_),
    .C(_168_),
    .Y(_175_)
);

NAND3X1 _6576_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_173_),
    .B(_175_),
    .C(_174_),
    .Y(_176_)
);

NAND3X1 _6577_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_172_),
    .B(_138_),
    .C(_176_),
    .Y(_177_)
);

INVX1 _6578_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_96_),
    .Y(_178_)
);

AOI21X1 _6579_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_82_),
    .B(_100_),
    .C(_178_),
    .Y(_179_)
);

AOI21X1 _6580_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_174_),
    .B(_175_),
    .C(_173_),
    .Y(_180_)
);

AOI21X1 _6581_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_171_),
    .B(_167_),
    .C(_152_),
    .Y(_181_)
);

OAI21X1 _6582_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_180_),
    .B(_181_),
    .C(_179_),
    .Y(_182_)
);

NAND3X1 _6583_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_136_),
    .B(_177_),
    .C(_182_),
    .Y(_183_)
);

AND2X2 _6584_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_134_),
    .B(_135_),
    .Y(_184_)
);

OAI21X1 _6585_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_180_),
    .B(_181_),
    .C(_138_),
    .Y(_185_)
);

NAND3X1 _6586_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_172_),
    .B(_176_),
    .C(_179_),
    .Y(_186_)
);

NAND3X1 _6587_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_184_),
    .B(_185_),
    .C(_186_),
    .Y(_187_)
);

AOI22X1 _6588_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_111_),
    .B(_106_),
    .C(_183_),
    .D(_187_),
    .Y(_188_)
);

AOI21X1 _6589_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_101_),
    .B(_105_),
    .C(_69_),
    .Y(_189_)
);

OAI21X1 _6590_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_112_),
    .B(_189_),
    .C(_106_),
    .Y(_190_)
);

NAND3X1 _6591_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_184_),
    .B(_177_),
    .C(_182_),
    .Y(_191_)
);

NAND3X1 _6592_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_136_),
    .B(_185_),
    .C(_186_),
    .Y(_192_)
);

AOI21X1 _6593_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_192_),
    .B(_191_),
    .C(_190_),
    .Y(_193_)
);

OAI21X1 _6594_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_193_),
    .B(_188_),
    .C(_116_),
    .Y(_194_)
);

AOI21X1 _6595_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_118_),
    .B(_117_),
    .C(_54_),
    .Y(_195_)
);

NAND3X1 _6596_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_190_),
    .B(_191_),
    .C(_192_),
    .Y(_196_)
);

INVX1 _6597_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_106_),
    .Y(_197_)
);

AOI21X1 _6598_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_26_),
    .B(_110_),
    .C(_197_),
    .Y(_198_)
);

AOI21X1 _6599_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_186_),
    .B(_185_),
    .C(_136_),
    .Y(_199_)
);

AOI21X1 _6600_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_182_),
    .B(_177_),
    .C(_184_),
    .Y(_200_)
);

OAI21X1 _6601_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_199_),
    .B(_200_),
    .C(_198_),
    .Y(_201_)
);

NAND3X1 _6602_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_195_),
    .B(_196_),
    .C(_201_),
    .Y(_202_)
);

NAND2X1 _6603_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_202_),
    .B(_194_),
    .Y(_203_)
);

AOI21X1 _6604_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_120_),
    .B(_126_),
    .C(_203_),
    .Y(_204_)
);

OAI21X1 _6605_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_129_),
    .B(_127_),
    .C(_120_),
    .Y(_205_)
);

AOI21X1 _6606_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_194_),
    .B(_202_),
    .C(_205_),
    .Y(_206_)
);

NOR2X1 _6607_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_204_),
    .B(_206_),
    .Y(_796_[6])
);

INVX1 _6608_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_202_),
    .Y(_207_)
);

AOI21X1 _6609_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_172_),
    .B(_176_),
    .C(_138_),
    .Y(_208_)
);

OAI21X1 _6610_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_136_),
    .B(_208_),
    .C(_177_),
    .Y(_209_)
);

NAND2X1 _6611_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[0]),
    .B(gnd),
    .Y(_210_)
);

INVX1 _6612_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_210_),
    .Y(_211_)
);

NAND2X1 _6613_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[1]),
    .B(gnd),
    .Y(_212_)
);

INVX1 _6614_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_212_),
    .Y(_213_)
);

AND2X2 _6615_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_145_),
    .B(_149_),
    .Y(_214_)
);

OAI21X1 _6616_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_139_),
    .B(_214_),
    .C(_143_),
    .Y(_215_)
);

NAND2X1 _6617_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_213_),
    .B(_215_),
    .Y(_216_)
);

NAND3X1 _6618_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_143_),
    .B(_212_),
    .C(_147_),
    .Y(_217_)
);

NAND3X1 _6619_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_211_),
    .B(_217_),
    .C(_216_),
    .Y(_218_)
);

AOI21X1 _6620_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_147_),
    .B(_143_),
    .C(_212_),
    .Y(_219_)
);

NOR2X1 _6621_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_213_),
    .B(_215_),
    .Y(_220_)
);

OAI21X1 _6622_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_219_),
    .B(_220_),
    .C(_210_),
    .Y(_221_)
);

NAND2X1 _6623_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_218_),
    .B(_221_),
    .Y(_222_)
);

AOI21X1 _6624_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_162_),
    .B(_166_),
    .C(_155_),
    .Y(_223_)
);

OAI21X1 _6625_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_173_),
    .B(_223_),
    .C(_167_),
    .Y(_224_)
);

NAND2X1 _6626_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[2]),
    .B(gnd),
    .Y(_225_)
);

INVX1 _6627_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_225_),
    .Y(_226_)
);

AND2X2 _6628_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[3]),
    .B(gnd),
    .Y(_227_)
);

AND2X2 _6629_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[7]),
    .Y(_228_)
);

NAND2X1 _6630_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_227_),
    .B(_228_),
    .Y(_229_)
);

AOI22X1 _6631_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[7]),
    .C(Xin[3]),
    .D(gnd),
    .Y(_230_)
);

INVX1 _6632_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_230_),
    .Y(_231_)
);

NAND3X1 _6633_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_226_),
    .B(_231_),
    .C(_229_),
    .Y(_232_)
);

INVX1 _6634_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_233_)
);

OAI21X1 _6635_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_15_),
    .B(_233_),
    .C(_228_),
    .Y(_234_)
);

INVX1 _6636_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[7]),
    .Y(_235_)
);

OAI21X1 _6637_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_778_),
    .B(_235_),
    .C(_227_),
    .Y(_236_)
);

NAND3X1 _6638_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_225_),
    .B(_234_),
    .C(_236_),
    .Y(_237_)
);

NAND2X1 _6639_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_232_),
    .B(_237_),
    .Y(_238_)
);

OAI21X1 _6640_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_156_),
    .B(_160_),
    .C(_159_),
    .Y(_239_)
);

NAND2X1 _6641_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[6]),
    .Y(_240_)
);

NAND2X1 _6642_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[4]),
    .Y(_241_)
);

AND2X2 _6643_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(Xin_5_bF$buf0),
    .Y(_242_)
);

NAND2X1 _6644_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_241_),
    .B(_242_),
    .Y(_243_)
);

OAI21X1 _6645_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_89_),
    .B(_74_),
    .C(_158_),
    .Y(_244_)
);

AOI21X1 _6646_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_244_),
    .B(_243_),
    .C(_240_),
    .Y(_245_)
);

INVX1 _6647_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_240_),
    .Y(_246_)
);

NAND2X1 _6648_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_158_),
    .B(_242_),
    .Y(_247_)
);

AOI22X1 _6649_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[4]),
    .C(vdd),
    .D(Xin_5_bF$buf3),
    .Y(_248_)
);

INVX1 _6650_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_248_),
    .Y(_249_)
);

AOI21X1 _6651_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_247_),
    .B(_249_),
    .C(_246_),
    .Y(_250_)
);

OAI21X1 _6652_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_250_),
    .B(_245_),
    .C(_239_),
    .Y(_251_)
);

AOI22X1 _6653_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_87_),
    .B(_158_),
    .C(_161_),
    .D(_157_),
    .Y(_252_)
);

NAND3X1 _6654_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_246_),
    .B(_249_),
    .C(_247_),
    .Y(_253_)
);

NAND2X1 _6655_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(Xin_5_bF$buf2),
    .Y(_254_)
);

NOR2X1 _6656_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_241_),
    .B(_254_),
    .Y(_255_)
);

OAI21X1 _6657_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_248_),
    .B(_255_),
    .C(_240_),
    .Y(_256_)
);

NAND3X1 _6658_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_253_),
    .B(_252_),
    .C(_256_),
    .Y(_257_)
);

AOI21X1 _6659_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_251_),
    .B(_257_),
    .C(_238_),
    .Y(_258_)
);

AND2X2 _6660_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_237_),
    .B(_232_),
    .Y(_259_)
);

NAND3X1 _6661_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_239_),
    .B(_253_),
    .C(_256_),
    .Y(_260_)
);

OAI21X1 _6662_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_250_),
    .B(_245_),
    .C(_252_),
    .Y(_261_)
);

AOI21X1 _6663_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_261_),
    .B(_260_),
    .C(_259_),
    .Y(_262_)
);

OAI21X1 _6664_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_258_),
    .B(_262_),
    .C(_224_),
    .Y(_263_)
);

INVX1 _6665_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_167_),
    .Y(_264_)
);

AOI21X1 _6666_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_152_),
    .B(_171_),
    .C(_264_),
    .Y(_265_)
);

NAND3X1 _6667_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_260_),
    .B(_259_),
    .C(_261_),
    .Y(_266_)
);

NAND3X1 _6668_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_238_),
    .B(_257_),
    .C(_251_),
    .Y(_267_)
);

NAND3X1 _6669_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_266_),
    .B(_267_),
    .C(_265_),
    .Y(_268_)
);

AOI21X1 _6670_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_268_),
    .B(_263_),
    .C(_222_),
    .Y(_269_)
);

AND2X2 _6671_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_221_),
    .B(_218_),
    .Y(_270_)
);

NAND3X1 _6672_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_224_),
    .B(_266_),
    .C(_267_),
    .Y(_271_)
);

OAI21X1 _6673_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_258_),
    .B(_262_),
    .C(_265_),
    .Y(_272_)
);

AOI21X1 _6674_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_272_),
    .B(_271_),
    .C(_270_),
    .Y(_273_)
);

OAI21X1 _6675_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_273_),
    .B(_269_),
    .C(_209_),
    .Y(_274_)
);

INVX1 _6676_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_177_),
    .Y(_275_)
);

AOI21X1 _6677_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_184_),
    .B(_182_),
    .C(_275_),
    .Y(_276_)
);

NAND3X1 _6678_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_271_),
    .B(_270_),
    .C(_272_),
    .Y(_277_)
);

NAND3X1 _6679_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_222_),
    .B(_263_),
    .C(_268_),
    .Y(_278_)
);

NAND3X1 _6680_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_277_),
    .B(_278_),
    .C(_276_),
    .Y(_279_)
);

AOI21X1 _6681_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_279_),
    .B(_274_),
    .C(_135_),
    .Y(_280_)
);

INVX1 _6682_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_135_),
    .Y(_281_)
);

NAND3X1 _6683_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_209_),
    .B(_277_),
    .C(_278_),
    .Y(_282_)
);

OAI21X1 _6684_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_269_),
    .B(_273_),
    .C(_276_),
    .Y(_283_)
);

AOI21X1 _6685_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_283_),
    .B(_282_),
    .C(_281_),
    .Y(_284_)
);

OAI21X1 _6686_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_284_),
    .B(_280_),
    .C(_196_),
    .Y(_285_)
);

NAND3X1 _6687_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_281_),
    .B(_282_),
    .C(_283_),
    .Y(_286_)
);

NAND3X1 _6688_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_135_),
    .B(_274_),
    .C(_279_),
    .Y(_287_)
);

NAND3X1 _6689_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_188_),
    .B(_286_),
    .C(_287_),
    .Y(_288_)
);

AND2X2 _6690_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_285_),
    .B(_288_),
    .Y(_289_)
);

OAI21X1 _6691_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_207_),
    .B(_204_),
    .C(_289_),
    .Y(_290_)
);

NOR2X1 _6692_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_207_),
    .B(_204_),
    .Y(_291_)
);

AOI21X1 _6693_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_287_),
    .B(_286_),
    .C(_188_),
    .Y(_292_)
);

INVX1 _6694_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_288_),
    .Y(_293_)
);

OAI21X1 _6695_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_292_),
    .B(_293_),
    .C(_291_),
    .Y(_294_)
);

AND2X2 _6696_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_294_),
    .B(_290_),
    .Y(_796_[7])
);

NAND3X1 _6697_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_285_),
    .B(_288_),
    .C(_204_),
    .Y(_295_)
);

AOI21X1 _6698_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_207_),
    .B(_285_),
    .C(_293_),
    .Y(_296_)
);

NAND2X1 _6699_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_296_),
    .B(_295_),
    .Y(_297_)
);

INVX1 _6700_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_282_),
    .Y(_298_)
);

AOI21X1 _6701_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_281_),
    .B(_283_),
    .C(_298_),
    .Y(_299_)
);

OAI21X1 _6702_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_210_),
    .B(_220_),
    .C(_216_),
    .Y(_300_)
);

INVX1 _6703_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_300_),
    .Y(_301_)
);

AOI21X1 _6704_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_266_),
    .B(_267_),
    .C(_224_),
    .Y(_302_)
);

OAI21X1 _6705_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_222_),
    .B(_302_),
    .C(_271_),
    .Y(_303_)
);

NAND2X1 _6706_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[1]),
    .B(gnd),
    .Y(_304_)
);

INVX2 _6707_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_305_)
);

NOR2X1 _6708_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_770_),
    .B(_305_),
    .Y(_306_)
);

OAI21X1 _6709_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_225_),
    .B(_230_),
    .C(_229_),
    .Y(_307_)
);

NOR2X1 _6710_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_306_),
    .B(_307_),
    .Y(_308_)
);

AND2X2 _6711_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_307_),
    .B(_306_),
    .Y(_309_)
);

OAI21X1 _6712_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_308_),
    .B(_309_),
    .C(_304_),
    .Y(_310_)
);

INVX1 _6713_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_304_),
    .Y(_311_)
);

OR2X2 _6714_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_307_),
    .B(_306_),
    .Y(_312_)
);

NAND2X1 _6715_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_306_),
    .B(_307_),
    .Y(_313_)
);

NAND3X1 _6716_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_311_),
    .B(_313_),
    .C(_312_),
    .Y(_314_)
);

NAND2X1 _6717_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_310_),
    .B(_314_),
    .Y(_315_)
);

AOI21X1 _6718_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_256_),
    .B(_253_),
    .C(_239_),
    .Y(_316_)
);

OAI21X1 _6719_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_238_),
    .B(_316_),
    .C(_260_),
    .Y(_317_)
);

NAND2X1 _6720_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[3]),
    .B(gnd),
    .Y(_318_)
);

INVX1 _6721_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_319_)
);

OAI21X1 _6722_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_15_),
    .B(_319_),
    .C(_25_),
    .Y(_320_)
);

NAND2X1 _6723_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[4]),
    .B(gnd),
    .Y(_321_)
);

OAI21X1 _6724_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_318_),
    .B(_321_),
    .C(_320_),
    .Y(_322_)
);

OAI21X1 _6725_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_240_),
    .B(_248_),
    .C(_247_),
    .Y(_323_)
);

NAND2X1 _6726_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[7]),
    .Y(_324_)
);

NAND2X1 _6727_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin_5_bF$buf1),
    .Y(_325_)
);

NAND3X1 _6728_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(Xin[6]),
    .C(_325_),
    .Y(_326_)
);

AND2X2 _6729_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin_5_bF$buf0),
    .Y(_327_)
);

OAI21X1 _6730_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_89_),
    .B(_144_),
    .C(_327_),
    .Y(_328_)
);

AOI21X1 _6731_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_328_),
    .B(_326_),
    .C(_324_),
    .Y(_329_)
);

INVX1 _6732_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_324_),
    .Y(_330_)
);

AND2X2 _6733_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(Xin[6]),
    .Y(_331_)
);

NAND2X1 _6734_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_327_),
    .B(_331_),
    .Y(_332_)
);

NAND2X1 _6735_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(Xin[6]),
    .Y(_333_)
);

NAND2X1 _6736_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_325_),
    .B(_333_),
    .Y(_334_)
);

AOI21X1 _6737_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_332_),
    .B(_334_),
    .C(_330_),
    .Y(_335_)
);

OAI21X1 _6738_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_335_),
    .B(_329_),
    .C(_323_),
    .Y(_336_)
);

AOI21X1 _6739_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_246_),
    .B(_249_),
    .C(_255_),
    .Y(_337_)
);

NAND3X1 _6740_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_330_),
    .B(_334_),
    .C(_332_),
    .Y(_338_)
);

NAND3X1 _6741_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_324_),
    .B(_326_),
    .C(_328_),
    .Y(_339_)
);

NAND3X1 _6742_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_338_),
    .B(_339_),
    .C(_337_),
    .Y(_340_)
);

AOI21X1 _6743_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_336_),
    .B(_340_),
    .C(_322_),
    .Y(_341_)
);

INVX1 _6744_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_322_),
    .Y(_342_)
);

NAND3X1 _6745_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_323_),
    .B(_338_),
    .C(_339_),
    .Y(_343_)
);

OAI21X1 _6746_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_335_),
    .B(_329_),
    .C(_337_),
    .Y(_344_)
);

AOI21X1 _6747_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_344_),
    .B(_343_),
    .C(_342_),
    .Y(_345_)
);

OAI21X1 _6748_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_341_),
    .B(_345_),
    .C(_317_),
    .Y(_346_)
);

INVX1 _6749_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_260_),
    .Y(_347_)
);

AOI21X1 _6750_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_259_),
    .B(_261_),
    .C(_347_),
    .Y(_348_)
);

NAND3X1 _6751_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_342_),
    .B(_343_),
    .C(_344_),
    .Y(_349_)
);

NAND3X1 _6752_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_322_),
    .B(_340_),
    .C(_336_),
    .Y(_350_)
);

NAND3X1 _6753_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_349_),
    .B(_350_),
    .C(_348_),
    .Y(_351_)
);

AOI21X1 _6754_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_351_),
    .B(_346_),
    .C(_315_),
    .Y(_352_)
);

AND2X2 _6755_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_314_),
    .B(_310_),
    .Y(_353_)
);

NAND3X1 _6756_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_349_),
    .B(_350_),
    .C(_317_),
    .Y(_354_)
);

OAI21X1 _6757_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_341_),
    .B(_345_),
    .C(_348_),
    .Y(_355_)
);

AOI21X1 _6758_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_355_),
    .B(_354_),
    .C(_353_),
    .Y(_356_)
);

OAI21X1 _6759_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_356_),
    .B(_352_),
    .C(_303_),
    .Y(_357_)
);

INVX1 _6760_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_271_),
    .Y(_358_)
);

AOI21X1 _6761_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_270_),
    .B(_272_),
    .C(_358_),
    .Y(_359_)
);

NAND3X1 _6762_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_353_),
    .B(_354_),
    .C(_355_),
    .Y(_360_)
);

NAND3X1 _6763_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_315_),
    .B(_346_),
    .C(_351_),
    .Y(_361_)
);

NAND3X1 _6764_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_360_),
    .B(_361_),
    .C(_359_),
    .Y(_362_)
);

AOI21X1 _6765_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_357_),
    .B(_362_),
    .C(_301_),
    .Y(_363_)
);

NAND3X1 _6766_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_303_),
    .B(_360_),
    .C(_361_),
    .Y(_364_)
);

OAI21X1 _6767_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_356_),
    .B(_352_),
    .C(_359_),
    .Y(_365_)
);

AOI21X1 _6768_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_365_),
    .B(_364_),
    .C(_300_),
    .Y(_366_)
);

OAI21X1 _6769_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_366_),
    .B(_363_),
    .C(_299_),
    .Y(_367_)
);

AOI21X1 _6770_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_278_),
    .B(_277_),
    .C(_209_),
    .Y(_368_)
);

OAI21X1 _6771_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_135_),
    .B(_368_),
    .C(_282_),
    .Y(_369_)
);

NAND3X1 _6772_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_300_),
    .B(_364_),
    .C(_365_),
    .Y(_370_)
);

NAND3X1 _6773_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_301_),
    .B(_362_),
    .C(_357_),
    .Y(_371_)
);

NAND3X1 _6774_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_369_),
    .B(_370_),
    .C(_371_),
    .Y(_372_)
);

NAND2X1 _6775_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_372_),
    .B(_367_),
    .Y(_373_)
);

NAND2X1 _6776_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_373_),
    .B(_297_),
    .Y(_374_)
);

OAI21X1 _6777_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_202_),
    .B(_292_),
    .C(_288_),
    .Y(_375_)
);

AOI21X1 _6778_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_289_),
    .B(_204_),
    .C(_375_),
    .Y(_376_)
);

AND2X2 _6779_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_367_),
    .B(_372_),
    .Y(_377_)
);

NAND2X1 _6780_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_377_),
    .B(_376_),
    .Y(_378_)
);

NAND2X1 _6781_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_374_),
    .B(_378_),
    .Y(_796_[8])
);

INVX1 _6782_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_372_),
    .Y(_379_)
);

AOI21X1 _6783_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_297_),
    .B(_367_),
    .C(_379_),
    .Y(_380_)
);

AOI21X1 _6784_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_361_),
    .B(_360_),
    .C(_303_),
    .Y(_381_)
);

OAI21X1 _6785_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_301_),
    .B(_381_),
    .C(_364_),
    .Y(_382_)
);

OAI21X1 _6786_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_304_),
    .B(_308_),
    .C(_313_),
    .Y(_383_)
);

AOI21X1 _6787_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_349_),
    .B(_350_),
    .C(_317_),
    .Y(_384_)
);

OAI21X1 _6788_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_315_),
    .B(_384_),
    .C(_354_),
    .Y(_385_)
);

NAND2X1 _6789_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[2]),
    .B(gnd),
    .Y(_386_)
);

NOR2X1 _6790_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_318_),
    .B(_321_),
    .Y(_387_)
);

NAND2X1 _6791_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_387_),
    .Y(_388_)
);

INVX1 _6792_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_388_),
    .Y(_389_)
);

AOI21X1 _6793_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[3]),
    .B(gnd),
    .C(_387_),
    .Y(_390_)
);

OAI21X1 _6794_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_390_),
    .B(_389_),
    .C(_386_),
    .Y(_391_)
);

INVX1 _6795_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_386_),
    .Y(_392_)
);

INVX1 _6796_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_390_),
    .Y(_393_)
);

NAND3X1 _6797_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_392_),
    .B(_388_),
    .C(_393_),
    .Y(_394_)
);

AND2X2 _6798_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_394_),
    .B(_391_),
    .Y(_395_)
);

AOI21X1 _6799_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_339_),
    .B(_338_),
    .C(_323_),
    .Y(_396_)
);

OAI21X1 _6800_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_322_),
    .B(_396_),
    .C(_343_),
    .Y(_397_)
);

NOR2X1 _6801_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_132_),
    .B(_321_),
    .Y(_398_)
);

AND2X2 _6802_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_132_),
    .B(_321_),
    .Y(_399_)
);

NOR2X1 _6803_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_398_),
    .B(_399_),
    .Y(_400_)
);

NAND2X1 _6804_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[6]),
    .Y(_401_)
);

AOI22X1 _6805_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin_5_bF$buf3),
    .C(vdd),
    .D(Xin[6]),
    .Y(_402_)
);

OAI22X1 _6806_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_254_),
    .B(_401_),
    .C(_324_),
    .D(_402_),
    .Y(_403_)
);

AOI22X1 _6807_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[6]),
    .C(vdd),
    .D(Xin[7]),
    .Y(_404_)
);

AND2X2 _6808_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[7]),
    .Y(_405_)
);

AOI21X1 _6809_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_331_),
    .B(_405_),
    .C(_404_),
    .Y(_406_)
);

NAND2X1 _6810_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_406_),
    .B(_403_),
    .Y(_407_)
);

AND2X2 _6811_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[6]),
    .Y(_408_)
);

AOI22X1 _6812_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_242_),
    .B(_408_),
    .C(_334_),
    .D(_330_),
    .Y(_409_)
);

NAND2X1 _6813_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(Xin[7]),
    .Y(_410_)
);

NAND2X1 _6814_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_401_),
    .B(_410_),
    .Y(_411_)
);

NAND2X1 _6815_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[7]),
    .Y(_412_)
);

OAI21X1 _6816_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_333_),
    .B(_412_),
    .C(_411_),
    .Y(_413_)
);

NAND2X1 _6817_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_413_),
    .B(_409_),
    .Y(_414_)
);

NAND3X1 _6818_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_400_),
    .B(_407_),
    .C(_414_),
    .Y(_415_)
);

NAND2X1 _6819_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin_5_bF$buf2),
    .B(gnd),
    .Y(_416_)
);

INVX1 _6820_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[4]),
    .Y(_417_)
);

OAI21X1 _6821_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_417_),
    .B(_319_),
    .C(_132_),
    .Y(_418_)
);

OAI21X1 _6822_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_25_),
    .B(_416_),
    .C(_418_),
    .Y(_419_)
);

NAND2X1 _6823_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_403_),
    .B(_413_),
    .Y(_420_)
);

NAND2X1 _6824_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_406_),
    .B(_409_),
    .Y(_421_)
);

NAND3X1 _6825_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_419_),
    .B(_420_),
    .C(_421_),
    .Y(_422_)
);

NAND3X1 _6826_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_415_),
    .B(_422_),
    .C(_397_),
    .Y(_423_)
);

NAND2X1 _6827_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_415_),
    .B(_422_),
    .Y(_424_)
);

NAND3X1 _6828_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_343_),
    .B(_349_),
    .C(_424_),
    .Y(_425_)
);

NAND3X1 _6829_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_395_),
    .B(_423_),
    .C(_425_),
    .Y(_426_)
);

NAND2X1 _6830_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_391_),
    .B(_394_),
    .Y(_427_)
);

AOI21X1 _6831_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_343_),
    .B(_349_),
    .C(_424_),
    .Y(_428_)
);

AOI21X1 _6832_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_415_),
    .B(_422_),
    .C(_397_),
    .Y(_429_)
);

OAI21X1 _6833_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_429_),
    .B(_428_),
    .C(_427_),
    .Y(_430_)
);

NAND3X1 _6834_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_426_),
    .B(_430_),
    .C(_385_),
    .Y(_431_)
);

INVX1 _6835_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_354_),
    .Y(_432_)
);

AOI21X1 _6836_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_353_),
    .B(_355_),
    .C(_432_),
    .Y(_433_)
);

INVX1 _6837_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_426_),
    .Y(_434_)
);

AOI21X1 _6838_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_425_),
    .B(_423_),
    .C(_395_),
    .Y(_435_)
);

OAI21X1 _6839_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_435_),
    .B(_434_),
    .C(_433_),
    .Y(_436_)
);

NAND3X1 _6840_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_383_),
    .B(_431_),
    .C(_436_),
    .Y(_437_)
);

INVX1 _6841_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_383_),
    .Y(_438_)
);

INVX1 _6842_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_431_),
    .Y(_439_)
);

AOI21X1 _6843_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_430_),
    .B(_426_),
    .C(_385_),
    .Y(_440_)
);

OAI21X1 _6844_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_440_),
    .B(_439_),
    .C(_438_),
    .Y(_441_)
);

NAND3X1 _6845_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_382_),
    .B(_437_),
    .C(_441_),
    .Y(_442_)
);

INVX1 _6846_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_364_),
    .Y(_443_)
);

AOI21X1 _6847_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_300_),
    .B(_365_),
    .C(_443_),
    .Y(_444_)
);

OAI21X1 _6848_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_435_),
    .B(_434_),
    .C(_385_),
    .Y(_445_)
);

NAND3X1 _6849_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_426_),
    .B(_430_),
    .C(_433_),
    .Y(_446_)
);

AOI21X1 _6850_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_446_),
    .B(_445_),
    .C(_438_),
    .Y(_447_)
);

AOI21X1 _6851_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_436_),
    .B(_431_),
    .C(_383_),
    .Y(_448_)
);

OAI21X1 _6852_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_447_),
    .B(_448_),
    .C(_444_),
    .Y(_449_)
);

AND2X2 _6853_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_449_),
    .B(_442_),
    .Y(_450_)
);

OR2X2 _6854_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_380_),
    .B(_450_),
    .Y(_451_)
);

NAND2X1 _6855_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_450_),
    .B(_380_),
    .Y(_452_)
);

NAND2X1 _6856_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_452_),
    .B(_451_),
    .Y(_796_[9])
);

NAND2X1 _6857_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_442_),
    .B(_449_),
    .Y(_453_)
);

NOR2X1 _6858_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_373_),
    .B(_453_),
    .Y(_454_)
);

NAND2X1 _6859_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_454_),
    .B(_297_),
    .Y(_455_)
);

AOI21X1 _6860_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_441_),
    .B(_437_),
    .C(_382_),
    .Y(_456_)
);

AOI21X1 _6861_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_372_),
    .B(_442_),
    .C(_456_),
    .Y(_457_)
);

INVX1 _6862_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_457_),
    .Y(_458_)
);

OAI21X1 _6863_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_438_),
    .B(_440_),
    .C(_431_),
    .Y(_459_)
);

OAI21X1 _6864_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_386_),
    .B(_390_),
    .C(_388_),
    .Y(_460_)
);

OAI21X1 _6865_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_427_),
    .B(_429_),
    .C(_423_),
    .Y(_461_)
);

INVX2 _6866_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_462_)
);

NOR3X1 _6867_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_305_),
    .B(_132_),
    .C(_321_),
    .Y(_463_)
);

OAI22X1 _6868_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_417_),
    .B(_305_),
    .C(_25_),
    .D(_416_),
    .Y(_464_)
);

INVX1 _6869_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_464_),
    .Y(_465_)
);

OAI22X1 _6870_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_15_),
    .B(_462_),
    .C(_463_),
    .D(_465_),
    .Y(_466_)
);

NOR2X1 _6871_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_15_),
    .B(_462_),
    .Y(_467_)
);

NAND2X1 _6872_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_398_),
    .Y(_468_)
);

NAND3X1 _6873_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_467_),
    .B(_464_),
    .C(_468_),
    .Y(_469_)
);

AND2X2 _6874_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_466_),
    .B(_469_),
    .Y(_470_)
);

NOR2X1 _6875_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_406_),
    .B(_403_),
    .Y(_471_)
);

OAI21X1 _6876_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_419_),
    .B(_471_),
    .C(_407_),
    .Y(_472_)
);

NAND2X1 _6877_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[6]),
    .Y(_473_)
);

NOR2X1 _6878_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_473_),
    .B(_416_),
    .Y(_474_)
);

AND2X2 _6879_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_473_),
    .B(_416_),
    .Y(_475_)
);

OAI22X1 _6880_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_331_),
    .B(_412_),
    .C(_474_),
    .D(_475_),
    .Y(_476_)
);

AND2X2 _6881_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[6]),
    .Y(_477_)
);

AND2X2 _6882_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin_5_bF$buf1),
    .B(gnd),
    .Y(_478_)
);

NAND2X1 _6883_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_477_),
    .B(_478_),
    .Y(_479_)
);

OAI21X1 _6884_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_74_),
    .B(_319_),
    .C(_473_),
    .Y(_480_)
);

AOI21X1 _6885_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(Xin[6]),
    .C(_412_),
    .Y(_481_)
);

NAND3X1 _6886_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_480_),
    .B(_481_),
    .C(_479_),
    .Y(_482_)
);

AND2X2 _6887_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_476_),
    .B(_482_),
    .Y(_483_)
);

NAND2X1 _6888_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_483_),
    .B(_472_),
    .Y(_484_)
);

NAND2X1 _6889_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_482_),
    .B(_476_),
    .Y(_485_)
);

NAND3X1 _6890_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_407_),
    .B(_485_),
    .C(_415_),
    .Y(_486_)
);

NAND3X1 _6891_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_470_),
    .B(_486_),
    .C(_484_),
    .Y(_487_)
);

NAND2X1 _6892_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_469_),
    .B(_466_),
    .Y(_488_)
);

NAND2X1 _6893_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_485_),
    .B(_472_),
    .Y(_489_)
);

NAND3X1 _6894_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_407_),
    .B(_483_),
    .C(_415_),
    .Y(_490_)
);

NAND3X1 _6895_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_488_),
    .B(_490_),
    .C(_489_),
    .Y(_491_)
);

NAND3X1 _6896_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_487_),
    .B(_491_),
    .C(_461_),
    .Y(_492_)
);

NAND2X1 _6897_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_491_),
    .B(_487_),
    .Y(_493_)
);

NAND3X1 _6898_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_423_),
    .B(_426_),
    .C(_493_),
    .Y(_494_)
);

NAND3X1 _6899_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_460_),
    .B(_494_),
    .C(_492_),
    .Y(_495_)
);

INVX1 _6900_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_460_),
    .Y(_496_)
);

NAND2X1 _6901_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_493_),
    .B(_461_),
    .Y(_497_)
);

AOI21X1 _6902_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_395_),
    .B(_425_),
    .C(_428_),
    .Y(_498_)
);

AND2X2 _6903_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_487_),
    .B(_491_),
    .Y(_499_)
);

NAND2X1 _6904_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_498_),
    .B(_499_),
    .Y(_500_)
);

NAND3X1 _6905_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_496_),
    .B(_497_),
    .C(_500_),
    .Y(_501_)
);

AOI21X1 _6906_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_495_),
    .B(_501_),
    .C(_459_),
    .Y(_502_)
);

NAND2X1 _6907_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_495_),
    .B(_501_),
    .Y(_503_)
);

AOI21X1 _6908_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_431_),
    .B(_437_),
    .C(_503_),
    .Y(_504_)
);

NOR2X1 _6909_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_502_),
    .B(_504_),
    .Y(_505_)
);

INVX1 _6910_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_505_),
    .Y(_506_)
);

AOI21X1 _6911_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_455_),
    .B(_458_),
    .C(_506_),
    .Y(_507_)
);

NAND2X1 _6912_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_377_),
    .B(_450_),
    .Y(_508_)
);

OAI21X1 _6913_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_508_),
    .B(_376_),
    .C(_458_),
    .Y(_509_)
);

NOR2X1 _6914_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_505_),
    .B(_509_),
    .Y(_510_)
);

NOR2X1 _6915_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_507_),
    .B(_510_),
    .Y(_796_[10])
);

NAND3X1 _6916_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_495_),
    .B(_501_),
    .C(_459_),
    .Y(_511_)
);

NAND2X1 _6917_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_505_),
    .B(_509_),
    .Y(_512_)
);

NOR2X1 _6918_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_493_),
    .B(_498_),
    .Y(_513_)
);

AOI21X1 _6919_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_460_),
    .B(_494_),
    .C(_513_),
    .Y(_514_)
);

NAND2X1 _6920_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_468_),
    .B(_469_),
    .Y(_515_)
);

NAND2X1 _6921_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_484_),
    .B(_487_),
    .Y(_516_)
);

NOR3X1 _6922_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_305_),
    .B(_473_),
    .C(_416_),
    .Y(_517_)
);

AOI22X1 _6923_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin_5_bF$buf0),
    .B(gnd),
    .C(_477_),
    .D(_478_),
    .Y(_518_)
);

OAI22X1 _6924_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_417_),
    .B(_462_),
    .C(_518_),
    .D(_517_),
    .Y(_519_)
);

NOR2X1 _6925_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_417_),
    .B(_462_),
    .Y(_520_)
);

NAND2X1 _6926_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_474_),
    .Y(_521_)
);

OAI21X1 _6927_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_74_),
    .B(_305_),
    .C(_479_),
    .Y(_522_)
);

NAND3X1 _6928_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_520_),
    .B(_521_),
    .C(_522_),
    .Y(_523_)
);

NAND2X1 _6929_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_519_),
    .B(_523_),
    .Y(_524_)
);

NAND2X1 _6930_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_331_),
    .B(_405_),
    .Y(_525_)
);

NAND2X1 _6931_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(Xin[7]),
    .Y(_526_)
);

OAI22X1 _6932_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_233_),
    .B(_235_),
    .C(_319_),
    .D(_144_),
    .Y(_527_)
);

OAI21X1 _6933_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_473_),
    .B(_526_),
    .C(_527_),
    .Y(_528_)
);

NAND3X1 _6934_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_525_),
    .B(_528_),
    .C(_482_),
    .Y(_529_)
);

INVX1 _6935_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_529_),
    .Y(_530_)
);

AOI21X1 _6936_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_482_),
    .B(_525_),
    .C(_528_),
    .Y(_531_)
);

OAI21X1 _6937_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_531_),
    .B(_530_),
    .C(_524_),
    .Y(_532_)
);

AND2X2 _6938_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_523_),
    .B(_519_),
    .Y(_533_)
);

INVX1 _6939_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_531_),
    .Y(_534_)
);

NAND3X1 _6940_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_529_),
    .B(_534_),
    .C(_533_),
    .Y(_535_)
);

AND2X2 _6941_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_535_),
    .B(_532_),
    .Y(_536_)
);

NAND2X1 _6942_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_536_),
    .B(_516_),
    .Y(_537_)
);

AOI21X1 _6943_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_415_),
    .B(_407_),
    .C(_485_),
    .Y(_538_)
);

AOI21X1 _6944_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_470_),
    .B(_486_),
    .C(_538_),
    .Y(_539_)
);

NAND2X1 _6945_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_532_),
    .B(_535_),
    .Y(_540_)
);

NAND2X1 _6946_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_540_),
    .B(_539_),
    .Y(_541_)
);

NAND3X1 _6947_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_515_),
    .B(_541_),
    .C(_537_),
    .Y(_542_)
);

INVX1 _6948_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_515_),
    .Y(_543_)
);

NAND2X1 _6949_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_540_),
    .B(_516_),
    .Y(_544_)
);

NAND2X1 _6950_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_539_),
    .B(_536_),
    .Y(_545_)
);

NAND3X1 _6951_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_543_),
    .B(_545_),
    .C(_544_),
    .Y(_546_)
);

NAND2X1 _6952_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_542_),
    .B(_546_),
    .Y(_547_)
);

NAND2X1 _6953_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_547_),
    .B(_514_),
    .Y(_548_)
);

AOI21X1 _6954_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_487_),
    .B(_491_),
    .C(_461_),
    .Y(_549_)
);

OAI21X1 _6955_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_496_),
    .B(_549_),
    .C(_492_),
    .Y(_550_)
);

NAND3X1 _6956_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_542_),
    .B(_546_),
    .C(_550_),
    .Y(_551_)
);

NAND2X1 _6957_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_548_),
    .B(_551_),
    .Y(_552_)
);

INVX1 _6958_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_552_),
    .Y(_553_)
);

NAND3X1 _6959_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_511_),
    .B(_553_),
    .C(_512_),
    .Y(_554_)
);

OAI21X1 _6960_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_504_),
    .B(_507_),
    .C(_552_),
    .Y(_555_)
);

NAND2X1 _6961_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_554_),
    .B(_555_),
    .Y(_796_[11])
);

NOR3X1 _6962_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_502_),
    .B(_504_),
    .C(_552_),
    .Y(_556_)
);

NAND3X1 _6963_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_454_),
    .B(_556_),
    .C(_297_),
    .Y(_557_)
);

OAI21X1 _6964_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_511_),
    .B(_552_),
    .C(_551_),
    .Y(_558_)
);

AOI21X1 _6965_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_556_),
    .B(_457_),
    .C(_558_),
    .Y(_559_)
);

AND2X2 _6966_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_542_),
    .B(_537_),
    .Y(_560_)
);

OAI21X1 _6967_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_305_),
    .B(_479_),
    .C(_523_),
    .Y(_561_)
);

OAI21X1 _6968_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_530_),
    .B(_524_),
    .C(_534_),
    .Y(_562_)
);

INVX1 _6969_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_562_),
    .Y(_563_)
);

INVX1 _6970_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_526_),
    .Y(_564_)
);

NOR2X1 _6971_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_74_),
    .B(_462_),
    .Y(_565_)
);

NOR2X1 _6972_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_473_),
    .B(_526_),
    .Y(_566_)
);

NOR2X1 _6973_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_144_),
    .B(_305_),
    .Y(_567_)
);

NOR2X1 _6974_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_567_),
    .B(_566_),
    .Y(_568_)
);

AOI21X1 _6975_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_566_),
    .C(_568_),
    .Y(_569_)
);

OR2X2 _6976_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_569_),
    .B(_565_),
    .Y(_570_)
);

NAND2X1 _6977_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_565_),
    .B(_569_),
    .Y(_571_)
);

NAND3X1 _6978_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_564_),
    .B(_571_),
    .C(_570_),
    .Y(_572_)
);

NOR2X1 _6979_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_565_),
    .B(_569_),
    .Y(_573_)
);

INVX1 _6980_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_571_),
    .Y(_574_)
);

OAI21X1 _6981_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_573_),
    .B(_574_),
    .C(_526_),
    .Y(_575_)
);

NAND2X1 _6982_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_572_),
    .B(_575_),
    .Y(_576_)
);

NAND2X1 _6983_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_563_),
    .B(_576_),
    .Y(_577_)
);

NAND3X1 _6984_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_562_),
    .B(_572_),
    .C(_575_),
    .Y(_578_)
);

AOI21X1 _6985_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_577_),
    .B(_578_),
    .C(_561_),
    .Y(_579_)
);

NAND3X1 _6986_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_561_),
    .B(_578_),
    .C(_577_),
    .Y(_580_)
);

INVX1 _6987_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_580_),
    .Y(_581_)
);

OAI21X1 _6988_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_579_),
    .B(_581_),
    .C(_560_),
    .Y(_582_)
);

OR2X2 _6989_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_581_),
    .B(_579_),
    .Y(_583_)
);

OR2X2 _6990_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_583_),
    .B(_560_),
    .Y(_584_)
);

NAND2X1 _6991_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_582_),
    .B(_584_),
    .Y(_585_)
);

AOI21X1 _6992_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_557_),
    .B(_559_),
    .C(_585_),
    .Y(_586_)
);

NAND3X1 _6993_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_377_),
    .B(_450_),
    .C(_556_),
    .Y(_587_)
);

OAI21X1 _6994_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_376_),
    .B(_587_),
    .C(_559_),
    .Y(_588_)
);

INVX1 _6995_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_585_),
    .Y(_589_)
);

NOR2X1 _6996_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_589_),
    .B(_588_),
    .Y(_590_)
);

NOR2X1 _6997_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_586_),
    .B(_590_),
    .Y(_796_[12])
);

NOR2X1 _6998_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_560_),
    .B(_583_),
    .Y(_591_)
);

INVX1 _6999_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_566_),
    .Y(_592_)
);

OAI21X1 _7000_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_305_),
    .B(_592_),
    .C(_571_),
    .Y(_593_)
);

INVX1 _7001_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_593_),
    .Y(_594_)
);

NOR2X1 _7002_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_235_),
    .B(_462_),
    .Y(_595_)
);

NAND2X1 _7003_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_567_),
    .B(_595_),
    .Y(_596_)
);

OAI22X1 _7004_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_144_),
    .B(_462_),
    .C(_305_),
    .D(_235_),
    .Y(_597_)
);

NAND2X1 _7005_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_597_),
    .B(_596_),
    .Y(_598_)
);

NAND2X1 _7006_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_598_),
    .B(_572_),
    .Y(_599_)
);

OR2X2 _7007_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_572_),
    .B(_598_),
    .Y(_600_)
);

NAND2X1 _7008_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_599_),
    .B(_600_),
    .Y(_601_)
);

NAND2X1 _7009_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_594_),
    .B(_601_),
    .Y(_602_)
);

OR2X2 _7010_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_601_),
    .B(_594_),
    .Y(_603_)
);

NAND2X1 _7011_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_602_),
    .B(_603_),
    .Y(_604_)
);

NAND3X1 _7012_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_578_),
    .B(_580_),
    .C(_604_),
    .Y(_605_)
);

OAI21X1 _7013_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_563_),
    .B(_576_),
    .C(_580_),
    .Y(_606_)
);

AND2X2 _7014_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_603_),
    .B(_602_),
    .Y(_607_)
);

NAND2X1 _7015_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_606_),
    .B(_607_),
    .Y(_608_)
);

NAND2X1 _7016_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_605_),
    .B(_608_),
    .Y(_609_)
);

OAI21X1 _7017_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_591_),
    .B(_586_),
    .C(_609_),
    .Y(_610_)
);

NAND2X1 _7018_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_589_),
    .B(_588_),
    .Y(_611_)
);

AND2X2 _7019_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_608_),
    .B(_605_),
    .Y(_612_)
);

NAND3X1 _7020_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_584_),
    .B(_612_),
    .C(_611_),
    .Y(_613_)
);

NAND2X1 _7021_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_613_),
    .B(_610_),
    .Y(_796_[13])
);

NAND3X1 _7022_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_582_),
    .B(_584_),
    .C(_612_),
    .Y(_614_)
);

AOI21X1 _7023_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_557_),
    .B(_559_),
    .C(_614_),
    .Y(_615_)
);

OAI21X1 _7024_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_584_),
    .B(_609_),
    .C(_608_),
    .Y(_616_)
);

OAI21X1 _7025_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_594_),
    .B(_601_),
    .C(_600_),
    .Y(_617_)
);

AND2X2 _7026_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_596_),
    .B(_595_),
    .Y(_618_)
);

OR2X2 _7027_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_617_),
    .B(_618_),
    .Y(_619_)
);

NAND2X1 _7028_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_618_),
    .B(_617_),
    .Y(_620_)
);

NAND2X1 _7029_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_620_),
    .B(_619_),
    .Y(_621_)
);

OAI21X1 _7030_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_616_),
    .B(_615_),
    .C(_621_),
    .Y(_622_)
);

INVX1 _7031_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_582_),
    .Y(_623_)
);

NOR3X1 _7032_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_623_),
    .B(_591_),
    .C(_609_),
    .Y(_624_)
);

NAND2X1 _7033_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_624_),
    .B(_588_),
    .Y(_625_)
);

INVX1 _7034_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_616_),
    .Y(_626_)
);

INVX1 _7035_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_621_),
    .Y(_627_)
);

NAND3X1 _7036_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_626_),
    .B(_627_),
    .C(_625_),
    .Y(_628_)
);

NAND2X1 _7037_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_628_),
    .B(_622_),
    .Y(_796_[14])
);

OAI21X1 _7038_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_616_),
    .B(_615_),
    .C(_627_),
    .Y(_629_)
);

OAI21X1 _7039_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_567_),
    .B(_617_),
    .C(_595_),
    .Y(_630_)
);

NAND2X1 _7040_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_630_),
    .B(_629_),
    .Y(_796_[15])
);

INVX1 _7041_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_24_),
    .Y(_791_[0])
);

AND2X2 _7042_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [0]),
    .B(\u_fir_pe0.mul [0]),
    .Y(_631_)
);

INVX1 _7043_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [1]),
    .Y(_632_)
);

INVX1 _7044_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.mul [1]),
    .Y(_633_)
);

NOR2X1 _7045_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_632_),
    .B(_633_),
    .Y(_634_)
);

NOR2X1 _7046_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [1]),
    .B(\u_fir_pe0.mul [1]),
    .Y(_635_)
);

NOR2X1 _7047_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_635_),
    .B(_634_),
    .Y(_636_)
);

NAND2X1 _7048_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_631_),
    .B(_636_),
    .Y(_637_)
);

INVX1 _7049_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_637_),
    .Y(_638_)
);

NOR2X1 _7050_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_631_),
    .B(_636_),
    .Y(_639_)
);

NOR2X1 _7051_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_639_),
    .B(_638_),
    .Y(_790_[1])
);

OAI21X1 _7052_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_632_),
    .B(_633_),
    .C(_637_),
    .Y(_640_)
);

AND2X2 _7053_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [2]),
    .B(\u_fir_pe0.mul [2]),
    .Y(_641_)
);

NOR2X1 _7054_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [2]),
    .B(\u_fir_pe0.mul [2]),
    .Y(_642_)
);

OAI21X1 _7055_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_641_),
    .B(_642_),
    .C(_640_),
    .Y(_643_)
);

INVX1 _7056_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_640_),
    .Y(_644_)
);

NOR2X1 _7057_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_642_),
    .B(_641_),
    .Y(_645_)
);

NAND2X1 _7058_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_645_),
    .B(_644_),
    .Y(_646_)
);

NAND2X1 _7059_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_643_),
    .B(_646_),
    .Y(_790_[2])
);

AOI21X1 _7060_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_640_),
    .B(_645_),
    .C(_641_),
    .Y(_647_)
);

INVX1 _7061_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [3]),
    .Y(_648_)
);

INVX1 _7062_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.mul [3]),
    .Y(_649_)
);

NOR2X1 _7063_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_648_),
    .B(_649_),
    .Y(_650_)
);

NOR2X1 _7064_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [3]),
    .B(\u_fir_pe0.mul [3]),
    .Y(_651_)
);

NOR2X1 _7065_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_651_),
    .B(_650_),
    .Y(_652_)
);

NAND2X1 _7066_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_652_),
    .B(_647_),
    .Y(_653_)
);

OR2X2 _7067_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_647_),
    .B(_652_),
    .Y(_654_)
);

NAND2X1 _7068_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_653_),
    .B(_654_),
    .Y(_790_[3])
);

INVX1 _7069_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [4]),
    .Y(_655_)
);

INVX1 _7070_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.mul [4]),
    .Y(_656_)
);

NOR2X1 _7071_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_655_),
    .B(_656_),
    .Y(_657_)
);

NOR2X1 _7072_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [4]),
    .B(\u_fir_pe0.mul [4]),
    .Y(_658_)
);

NOR2X1 _7073_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_658_),
    .B(_657_),
    .Y(_659_)
);

INVX1 _7074_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_650_),
    .Y(_660_)
);

OAI21X1 _7075_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_651_),
    .B(_647_),
    .C(_660_),
    .Y(_661_)
);

NAND2X1 _7076_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_659_),
    .B(_661_),
    .Y(_662_)
);

OR2X2 _7077_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_661_),
    .B(_659_),
    .Y(_663_)
);

AND2X2 _7078_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_663_),
    .B(_662_),
    .Y(_790_[4])
);

OAI21X1 _7079_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_655_),
    .B(_656_),
    .C(_662_),
    .Y(_664_)
);

INVX1 _7080_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [5]),
    .Y(_665_)
);

INVX1 _7081_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.mul [5]),
    .Y(_666_)
);

NOR2X1 _7082_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_665_),
    .B(_666_),
    .Y(_667_)
);

NOR2X1 _7083_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [5]),
    .B(\u_fir_pe0.mul [5]),
    .Y(_668_)
);

NOR2X1 _7084_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_668_),
    .B(_667_),
    .Y(_669_)
);

NAND2X1 _7085_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_669_),
    .B(_664_),
    .Y(_670_)
);

OR2X2 _7086_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_664_),
    .B(_669_),
    .Y(_671_)
);

AND2X2 _7087_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_671_),
    .B(_670_),
    .Y(_790_[5])
);

OAI21X1 _7088_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_665_),
    .B(_666_),
    .C(_670_),
    .Y(_672_)
);

INVX1 _7089_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [6]),
    .Y(_673_)
);

INVX1 _7090_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.mul [6]),
    .Y(_674_)
);

NOR2X1 _7091_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_673_),
    .B(_674_),
    .Y(_675_)
);

NOR2X1 _7092_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [6]),
    .B(\u_fir_pe0.mul [6]),
    .Y(_676_)
);

NOR2X1 _7093_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_676_),
    .B(_675_),
    .Y(_677_)
);

NAND2X1 _7094_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_677_),
    .B(_672_),
    .Y(_678_)
);

OR2X2 _7095_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_672_),
    .B(_677_),
    .Y(_679_)
);

AND2X2 _7096_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_679_),
    .B(_678_),
    .Y(_790_[6])
);

OAI21X1 _7097_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_673_),
    .B(_674_),
    .C(_678_),
    .Y(_680_)
);

INVX1 _7098_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [7]),
    .Y(_681_)
);

INVX1 _7099_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.mul [7]),
    .Y(_682_)
);

NOR2X1 _7100_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_681_),
    .B(_682_),
    .Y(_683_)
);

NOR2X1 _7101_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [7]),
    .B(\u_fir_pe0.mul [7]),
    .Y(_684_)
);

OAI21X1 _7102_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_683_),
    .B(_684_),
    .C(_680_),
    .Y(_685_)
);

INVX1 _7103_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_680_),
    .Y(_686_)
);

NOR2X1 _7104_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_684_),
    .B(_683_),
    .Y(_687_)
);

NAND2X1 _7105_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_687_),
    .B(_686_),
    .Y(_688_)
);

NAND2X1 _7106_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_685_),
    .B(_688_),
    .Y(_790_[7])
);

INVX1 _7107_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [8]),
    .Y(_690_)
);

INVX1 _7108_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.mul [8]),
    .Y(_691_)
);

NOR2X1 _7109_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_690_),
    .B(_691_),
    .Y(_692_)
);

NOR2X1 _7110_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [8]),
    .B(\u_fir_pe0.mul [8]),
    .Y(_693_)
);

NAND2X1 _7111_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_657_),
    .B(_669_),
    .Y(_694_)
);

OAI21X1 _7112_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_665_),
    .B(_666_),
    .C(_694_),
    .Y(_695_)
);

NAND2X1 _7113_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_675_),
    .B(_687_),
    .Y(_696_)
);

OAI21X1 _7114_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_681_),
    .B(_682_),
    .C(_696_),
    .Y(_697_)
);

AND2X2 _7115_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_677_),
    .B(_687_),
    .Y(_698_)
);

AOI21X1 _7116_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_695_),
    .B(_698_),
    .C(_697_),
    .Y(_699_)
);

AND2X2 _7117_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_659_),
    .B(_669_),
    .Y(_701_)
);

NAND3X1 _7118_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_701_),
    .B(_698_),
    .C(_661_),
    .Y(_702_)
);

NAND2X1 _7119_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_699_),
    .B(_702_),
    .Y(_703_)
);

OAI21X1 _7120_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_692_),
    .B(_693_),
    .C(_703_),
    .Y(_704_)
);

NOR2X1 _7121_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_693_),
    .B(_692_),
    .Y(_705_)
);

INVX1 _7122_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_703_),
    .Y(_706_)
);

NAND2X1 _7123_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_705_),
    .B(_706_),
    .Y(_707_)
);

NAND2X1 _7124_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_704_),
    .B(_707_),
    .Y(_790_[8])
);

INVX1 _7125_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_692_),
    .Y(_708_)
);

INVX1 _7126_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_705_),
    .Y(_709_)
);

OAI21X1 _7127_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_709_),
    .B(_706_),
    .C(_708_),
    .Y(_711_)
);

AND2X2 _7128_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [9]),
    .B(\u_fir_pe0.mul [9]),
    .Y(_712_)
);

NOR2X1 _7129_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [9]),
    .B(\u_fir_pe0.mul [9]),
    .Y(_713_)
);

NOR2X1 _7130_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_713_),
    .B(_712_),
    .Y(_714_)
);

INVX1 _7131_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_714_),
    .Y(_715_)
);

OR2X2 _7132_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_711_),
    .B(_715_),
    .Y(_716_)
);

OAI21X1 _7133_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_712_),
    .B(_713_),
    .C(_711_),
    .Y(_717_)
);

NAND2X1 _7134_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_717_),
    .B(_716_),
    .Y(_790_[9])
);

NOR2X1 _7135_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_715_),
    .B(_709_),
    .Y(_718_)
);

AOI21X1 _7136_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_714_),
    .B(_692_),
    .C(_712_),
    .Y(_719_)
);

INVX1 _7137_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_719_),
    .Y(_721_)
);

AOI21X1 _7138_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_703_),
    .B(_718_),
    .C(_721_),
    .Y(_722_)
);

INVX1 _7139_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_722_),
    .Y(_723_)
);

INVX1 _7140_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [10]),
    .Y(_724_)
);

INVX1 _7141_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.mul [10]),
    .Y(_725_)
);

NOR2X1 _7142_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_724_),
    .B(_725_),
    .Y(_726_)
);

NOR2X1 _7143_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [10]),
    .B(\u_fir_pe0.mul [10]),
    .Y(_727_)
);

NOR2X1 _7144_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_727_),
    .B(_726_),
    .Y(_728_)
);

NAND2X1 _7145_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_728_),
    .B(_723_),
    .Y(_729_)
);

OAI21X1 _7146_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_726_),
    .B(_727_),
    .C(_722_),
    .Y(_730_)
);

AND2X2 _7147_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_729_),
    .B(_730_),
    .Y(_790_[10])
);

OAI21X1 _7148_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_724_),
    .B(_725_),
    .C(_729_),
    .Y(_732_)
);

AND2X2 _7149_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [11]),
    .B(\u_fir_pe0.mul [11]),
    .Y(_733_)
);

NOR2X1 _7150_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [11]),
    .B(\u_fir_pe0.mul [11]),
    .Y(_734_)
);

NOR2X1 _7151_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_734_),
    .B(_733_),
    .Y(_735_)
);

NOR2X1 _7152_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_735_),
    .B(_732_),
    .Y(_736_)
);

AND2X2 _7153_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_732_),
    .B(_735_),
    .Y(_737_)
);

NOR2X1 _7154_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_736_),
    .B(_737_),
    .Y(_790_[11])
);

AOI21X1 _7155_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_735_),
    .B(_726_),
    .C(_733_),
    .Y(_738_)
);

NAND2X1 _7156_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_735_),
    .B(_728_),
    .Y(_739_)
);

OAI21X1 _7157_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_739_),
    .B(_722_),
    .C(_738_),
    .Y(_741_)
);

INVX1 _7158_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [12]),
    .Y(_742_)
);

INVX1 _7159_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.mul [12]),
    .Y(_743_)
);

NOR2X1 _7160_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_742_),
    .B(_743_),
    .Y(_744_)
);

NOR2X1 _7161_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [12]),
    .B(\u_fir_pe0.mul [12]),
    .Y(_745_)
);

NOR2X1 _7162_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_745_),
    .B(_744_),
    .Y(_746_)
);

NAND2X1 _7163_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_746_),
    .B(_741_),
    .Y(_747_)
);

OR2X2 _7164_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_741_),
    .B(_746_),
    .Y(_748_)
);

AND2X2 _7165_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_748_),
    .B(_747_),
    .Y(_790_[12])
);

OAI21X1 _7166_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_742_),
    .B(_743_),
    .C(_747_),
    .Y(_749_)
);

INVX1 _7167_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [13]),
    .Y(_751_)
);

INVX1 _7168_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.mul [13]),
    .Y(_752_)
);

NOR2X1 _7169_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_751_),
    .B(_752_),
    .Y(_753_)
);

NOR2X1 _7170_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [13]),
    .B(\u_fir_pe0.mul [13]),
    .Y(_754_)
);

NOR2X1 _7171_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_754_),
    .B(_753_),
    .Y(_755_)
);

NAND2X1 _7172_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_755_),
    .B(_749_),
    .Y(_756_)
);

OR2X2 _7173_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_749_),
    .B(_755_),
    .Y(_757_)
);

AND2X2 _7174_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_757_),
    .B(_756_),
    .Y(_790_[13])
);

OAI21X1 _7175_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_751_),
    .B(_752_),
    .C(_756_),
    .Y(_758_)
);

INVX1 _7176_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [14]),
    .Y(_759_)
);

INVX1 _7177_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.mul [14]),
    .Y(_761_)
);

NOR2X1 _7178_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_759_),
    .B(_761_),
    .Y(_762_)
);

NOR2X1 _7179_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [14]),
    .B(\u_fir_pe0.mul [14]),
    .Y(_763_)
);

NOR2X1 _7180_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_763_),
    .B(_762_),
    .Y(_764_)
);

AND2X2 _7181_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_758_),
    .B(_764_),
    .Y(_765_)
);

NOR2X1 _7182_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_764_),
    .B(_758_),
    .Y(_766_)
);

NOR2X1 _7183_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_766_),
    .B(_765_),
    .Y(_790_[14])
);

INVX1 _7184_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_762_),
    .Y(_767_)
);

NAND2X1 _7185_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_764_),
    .B(_758_),
    .Y(_768_)
);

NAND2X1 _7186_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [15]),
    .B(\u_fir_pe0.mul [15]),
    .Y(_769_)
);

OR2X2 _7187_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [15]),
    .B(\u_fir_pe0.mul [15]),
    .Y(_771_)
);

NAND2X1 _7188_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_769_),
    .B(_771_),
    .Y(_772_)
);

INVX1 _7189_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_772_),
    .Y(_773_)
);

NAND3X1 _7190_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_767_),
    .B(_773_),
    .C(_768_),
    .Y(_774_)
);

OAI21X1 _7191_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_762_),
    .B(_765_),
    .C(_772_),
    .Y(_775_)
);

NAND2X1 _7192_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_774_),
    .B(_775_),
    .Y(_790_[15])
);

NOR2X1 _7193_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe0.rYin [0]),
    .B(\u_fir_pe0.mul [0]),
    .Y(_776_)
);

NOR2X1 _7194_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_776_),
    .B(_631_),
    .Y(_789_[0])
);

AOI21X1 _7195_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[0]),
    .B(gnd),
    .C(_700_),
    .Y(_777_)
);

NOR2X1 _7196_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_777_),
    .B(_720_),
    .Y(_792_[1])
);

NOR2X1 _7197_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720_),
    .B(_784_),
    .Y(_779_)
);

NOR2X1 _7198_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_779_),
    .B(_786_),
    .Y(_793_[2])
);

DFFPOSX1 _7199_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf7),
    .D(_789_[0]),
    .Q(\Y[1] [0])
);

DFFPOSX1 _7200_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_790_[1]),
    .Q(\Y[1] [1])
);

DFFPOSX1 _7201_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_790_[2]),
    .Q(\Y[1] [2])
);

DFFPOSX1 _7202_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_790_[3]),
    .Q(\Y[1] [3])
);

DFFPOSX1 _7203_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_790_[4]),
    .Q(\Y[1] [4])
);

DFFPOSX1 _7204_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_790_[5]),
    .Q(\Y[1] [5])
);

DFFPOSX1 _7205_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_790_[6]),
    .Q(\Y[1] [6])
);

DFFPOSX1 _7206_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_790_[7]),
    .Q(\Y[1] [7])
);

DFFPOSX1 _7207_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf57),
    .D(_790_[8]),
    .Q(\Y[1] [8])
);

DFFPOSX1 _7208_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf56),
    .D(_790_[9]),
    .Q(\Y[1] [9])
);

DFFPOSX1 _7209_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf55),
    .D(_790_[10]),
    .Q(\Y[1] [10])
);

DFFPOSX1 _7210_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf54),
    .D(_790_[11]),
    .Q(\Y[1] [11])
);

DFFPOSX1 _7211_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf53),
    .D(_790_[12]),
    .Q(\Y[1] [12])
);

DFFPOSX1 _7212_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf52),
    .D(_790_[13]),
    .Q(\Y[1] [13])
);

DFFPOSX1 _7213_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf51),
    .D(_790_[14]),
    .Q(\Y[1] [14])
);

DFFPOSX1 _7214_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf50),
    .D(_790_[15]),
    .Q(\Y[1] [15])
);

DFFPOSX1 _7215_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf49),
    .D(Xin[0]),
    .Q(\X[1] [0])
);

DFFPOSX1 _7216_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf48),
    .D(Xin[1]),
    .Q(\X[1] [1])
);

DFFPOSX1 _7217_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf47),
    .D(Xin[2]),
    .Q(\X[1] [2])
);

DFFPOSX1 _7218_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf46),
    .D(Xin[3]),
    .Q(\X[1] [3])
);

DFFPOSX1 _7219_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf45),
    .D(Xin[4]),
    .Q(\X[1] [4])
);

DFFPOSX1 _7220_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf44),
    .D(Xin_5_bF$buf3),
    .Q(\X[1] [5])
);

DFFPOSX1 _7221_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf43),
    .D(Xin[6]),
    .Q(\X[1] [6])
);

DFFPOSX1 _7222_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf42),
    .D(Xin[7]),
    .Q(\X[1] [7])
);

DFFPOSX1 _7223_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf41),
    .D(Yin[0]),
    .Q(\u_fir_pe0.rYin [0])
);

DFFPOSX1 _7224_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf40),
    .D(Yin[1]),
    .Q(\u_fir_pe0.rYin [1])
);

DFFPOSX1 _7225_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf39),
    .D(Yin[2]),
    .Q(\u_fir_pe0.rYin [2])
);

DFFPOSX1 _7226_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf38),
    .D(Yin[3]),
    .Q(\u_fir_pe0.rYin [3])
);

DFFPOSX1 _7227_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf37),
    .D(Yin[4]),
    .Q(\u_fir_pe0.rYin [4])
);

DFFPOSX1 _7228_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf36),
    .D(Yin[5]),
    .Q(\u_fir_pe0.rYin [5])
);

DFFPOSX1 _7229_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf35),
    .D(Yin[6]),
    .Q(\u_fir_pe0.rYin [6])
);

DFFPOSX1 _7230_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf34),
    .D(Yin[7]),
    .Q(\u_fir_pe0.rYin [7])
);

DFFPOSX1 _7231_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf33),
    .D(Yin[8]),
    .Q(\u_fir_pe0.rYin [8])
);

DFFPOSX1 _7232_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf32),
    .D(Yin[9]),
    .Q(\u_fir_pe0.rYin [9])
);

DFFPOSX1 _7233_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf31),
    .D(Yin[10]),
    .Q(\u_fir_pe0.rYin [10])
);

DFFPOSX1 _7234_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf30),
    .D(Yin[11]),
    .Q(\u_fir_pe0.rYin [11])
);

DFFPOSX1 _7235_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf29),
    .D(Yin[12]),
    .Q(\u_fir_pe0.rYin [12])
);

DFFPOSX1 _7236_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf28),
    .D(Yin[13]),
    .Q(\u_fir_pe0.rYin [13])
);

DFFPOSX1 _7237_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf27),
    .D(Yin[14]),
    .Q(\u_fir_pe0.rYin [14])
);

DFFPOSX1 _7238_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf26),
    .D(Yin[15]),
    .Q(\u_fir_pe0.rYin [15])
);

DFFPOSX1 _7239_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf25),
    .D(_791_[0]),
    .Q(\u_fir_pe0.mul [0])
);

DFFPOSX1 _7240_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf24),
    .D(_792_[1]),
    .Q(\u_fir_pe0.mul [1])
);

DFFPOSX1 _7241_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf23),
    .D(_793_[2]),
    .Q(\u_fir_pe0.mul [2])
);

DFFPOSX1 _7242_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf22),
    .D(_794_[3]),
    .Q(\u_fir_pe0.mul [3])
);

DFFPOSX1 _7243_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf21),
    .D(_795_[4]),
    .Q(\u_fir_pe0.mul [4])
);

DFFPOSX1 _7244_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf20),
    .D(_796_[5]),
    .Q(\u_fir_pe0.mul [5])
);

DFFPOSX1 _7245_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf19),
    .D(_796_[6]),
    .Q(\u_fir_pe0.mul [6])
);

DFFPOSX1 _7246_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf18),
    .D(_796_[7]),
    .Q(\u_fir_pe0.mul [7])
);

DFFPOSX1 _7247_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf17),
    .D(_796_[8]),
    .Q(\u_fir_pe0.mul [8])
);

DFFPOSX1 _7248_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf16),
    .D(_796_[9]),
    .Q(\u_fir_pe0.mul [9])
);

DFFPOSX1 _7249_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf15),
    .D(_796_[10]),
    .Q(\u_fir_pe0.mul [10])
);

DFFPOSX1 _7250_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf14),
    .D(_796_[11]),
    .Q(\u_fir_pe0.mul [11])
);

DFFPOSX1 _7251_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf13),
    .D(_796_[12]),
    .Q(\u_fir_pe0.mul [12])
);

DFFPOSX1 _7252_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf12),
    .D(_796_[13]),
    .Q(\u_fir_pe0.mul [13])
);

DFFPOSX1 _7253_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf11),
    .D(_796_[14]),
    .Q(\u_fir_pe0.mul [14])
);

DFFPOSX1 _7254_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf10),
    .D(_796_[15]),
    .Q(\u_fir_pe0.mul [15])
);

NAND2X1 _7255_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [0]),
    .B(gnd),
    .Y(_1486_)
);

AND2X2 _7256_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [1]),
    .B(gnd),
    .Y(_1497_)
);

INVX1 _7257_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1497_),
    .Y(_1507_)
);

NOR2X1 _7258_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1486_),
    .B(_1507_),
    .Y(_1517_)
);

NAND2X1 _7259_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [1]),
    .Y(_1528_)
);

NOR2X1 _7260_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1486_),
    .B(_1528_),
    .Y(_1537_)
);

AOI22X1 _7261_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [0]),
    .B(vdd),
    .C(\X[1] [1]),
    .D(gnd),
    .Y(_1547_)
);

NOR2X1 _7262_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1547_),
    .B(_1537_),
    .Y(_1557_)
);

INVX1 _7263_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [2]),
    .Y(_1567_)
);

INVX2 _7264_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_1575_)
);

NOR2X1 _7265_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1567_),
    .B(_1575_),
    .Y(_1577_)
);

NAND2X1 _7266_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1577_),
    .B(_1557_),
    .Y(_1578_)
);

INVX1 _7267_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1578_),
    .Y(_1579_)
);

NOR2X1 _7268_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1577_),
    .B(_1557_),
    .Y(_1580_)
);

NOR2X1 _7269_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1580_),
    .B(_1579_),
    .Y(_1581_)
);

NAND2X1 _7270_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1517_),
    .B(_1581_),
    .Y(_1582_)
);

INVX1 _7271_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1582_),
    .Y(_1583_)
);

NAND2X1 _7272_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1] [3]),
    .Y(_1584_)
);

INVX1 _7273_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1584_),
    .Y(_1585_)
);

NAND2X1 _7274_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1] [2]),
    .Y(_797_)
);

INVX1 _7275_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_797_),
    .Y(_798_)
);

NAND2X1 _7276_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [0]),
    .Y(_799_)
);

OR2X2 _7277_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1528_),
    .B(_799_),
    .Y(_800_)
);

AOI22X1 _7278_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [0]),
    .C(vdd),
    .D(\X[1] [1]),
    .Y(_801_)
);

INVX1 _7279_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_801_),
    .Y(_802_)
);

NAND3X1 _7280_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_798_),
    .B(_802_),
    .C(_800_),
    .Y(_803_)
);

NOR2X1 _7281_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1528_),
    .B(_799_),
    .Y(_804_)
);

OAI21X1 _7282_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_801_),
    .B(_804_),
    .C(_797_),
    .Y(_805_)
);

NAND3X1 _7283_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1537_),
    .B(_805_),
    .C(_803_),
    .Y(_806_)
);

INVX1 _7284_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1537_),
    .Y(_807_)
);

NAND3X1 _7285_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_797_),
    .B(_802_),
    .C(_800_),
    .Y(_808_)
);

OAI21X1 _7286_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_801_),
    .B(_804_),
    .C(_798_),
    .Y(_809_)
);

NAND3X1 _7287_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_807_),
    .B(_809_),
    .C(_808_),
    .Y(_810_)
);

NAND3X1 _7288_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1585_),
    .B(_810_),
    .C(_806_),
    .Y(_811_)
);

INVX2 _7289_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [3]),
    .Y(_812_)
);

NAND2X1 _7290_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_810_),
    .B(_806_),
    .Y(_813_)
);

OAI21X1 _7291_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1575_),
    .B(_812_),
    .C(_813_),
    .Y(_814_)
);

NAND2X1 _7292_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_811_),
    .B(_814_),
    .Y(_815_)
);

NAND2X1 _7293_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1578_),
    .B(_815_),
    .Y(_816_)
);

NAND3X1 _7294_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1579_),
    .B(_811_),
    .C(_814_),
    .Y(_817_)
);

NAND3X1 _7295_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_817_),
    .B(_1583_),
    .C(_816_),
    .Y(_818_)
);

INVX1 _7296_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_818_),
    .Y(_819_)
);

AOI21X1 _7297_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_816_),
    .B(_817_),
    .C(_1583_),
    .Y(_820_)
);

NOR2X1 _7298_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_820_),
    .B(_819_),
    .Y(_1591_[3])
);

NAND2X1 _7299_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [0]),
    .B(gnd),
    .Y(_821_)
);

NAND2X1 _7300_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [4]),
    .B(gnd),
    .Y(_822_)
);

NOR2X1 _7301_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_821_),
    .B(_822_),
    .Y(_823_)
);

AOI22X1 _7302_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [0]),
    .B(gnd),
    .C(gnd),
    .D(\X[1] [4]),
    .Y(_824_)
);

NOR2X1 _7303_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_824_),
    .B(_823_),
    .Y(_825_)
);

INVX1 _7304_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_825_),
    .Y(_826_)
);

NAND2X1 _7305_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [0]),
    .B(vdd),
    .Y(_827_)
);

NAND2X1 _7306_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [1]),
    .Y(_828_)
);

OAI22X1 _7307_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_827_),
    .B(_828_),
    .C(_797_),
    .D(_801_),
    .Y(_829_)
);

NAND2X1 _7308_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1] [3]),
    .Y(_830_)
);

INVX1 _7309_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_830_),
    .Y(_831_)
);

AND2X2 _7310_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [1]),
    .Y(_832_)
);

AND2X2 _7311_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [2]),
    .Y(_833_)
);

NAND2X1 _7312_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_832_),
    .B(_833_),
    .Y(_834_)
);

AOI22X1 _7313_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [1]),
    .C(vdd),
    .D(\X[1] [2]),
    .Y(_835_)
);

INVX1 _7314_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_835_),
    .Y(_836_)
);

NAND3X1 _7315_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_831_),
    .B(_836_),
    .C(_834_),
    .Y(_837_)
);

NAND3X1 _7316_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [2]),
    .C(_828_),
    .Y(_838_)
);

NAND2X1 _7317_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [2]),
    .Y(_839_)
);

NAND3X1 _7318_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [1]),
    .C(_839_),
    .Y(_840_)
);

NAND3X1 _7319_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_830_),
    .B(_838_),
    .C(_840_),
    .Y(_841_)
);

NAND3X1 _7320_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_829_),
    .B(_841_),
    .C(_837_),
    .Y(_842_)
);

INVX1 _7321_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_829_),
    .Y(_843_)
);

NAND2X1 _7322_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_841_),
    .B(_837_),
    .Y(_844_)
);

NAND2X1 _7323_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_843_),
    .B(_844_),
    .Y(_845_)
);

NAND3X1 _7324_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_826_),
    .B(_842_),
    .C(_845_),
    .Y(_846_)
);

NAND2X1 _7325_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_829_),
    .B(_844_),
    .Y(_847_)
);

NAND3X1 _7326_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_837_),
    .B(_841_),
    .C(_843_),
    .Y(_848_)
);

NAND3X1 _7327_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_825_),
    .B(_848_),
    .C(_847_),
    .Y(_849_)
);

AOI22X1 _7328_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_806_),
    .B(_811_),
    .C(_846_),
    .D(_849_),
    .Y(_850_)
);

INVX1 _7329_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_850_),
    .Y(_851_)
);

NAND2X1 _7330_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_806_),
    .B(_811_),
    .Y(_852_)
);

NAND2X1 _7331_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_846_),
    .B(_849_),
    .Y(_853_)
);

OR2X2 _7332_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_853_),
    .B(_852_),
    .Y(_854_)
);

NAND2X1 _7333_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_851_),
    .B(_854_),
    .Y(_855_)
);

OAI21X1 _7334_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1578_),
    .B(_815_),
    .C(_818_),
    .Y(_856_)
);

OR2X2 _7335_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_856_),
    .B(_855_),
    .Y(_857_)
);

NAND3X1 _7336_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_825_),
    .B(_842_),
    .C(_845_),
    .Y(_858_)
);

INVX1 _7337_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_842_),
    .Y(_859_)
);

AOI21X1 _7338_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_837_),
    .B(_841_),
    .C(_829_),
    .Y(_860_)
);

OAI21X1 _7339_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_860_),
    .B(_859_),
    .C(_826_),
    .Y(_861_)
);

AOI21X1 _7340_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_858_),
    .B(_861_),
    .C(_852_),
    .Y(_862_)
);

OAI21X1 _7341_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_850_),
    .B(_862_),
    .C(_856_),
    .Y(_863_)
);

NAND2X1 _7342_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_863_),
    .B(_857_),
    .Y(_1592_[4])
);

NOR2X1 _7343_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_818_),
    .B(_855_),
    .Y(_864_)
);

NOR3X1 _7344_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_850_),
    .B(_817_),
    .C(_862_),
    .Y(_865_)
);

OAI21X1 _7345_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_826_),
    .B(_860_),
    .C(_842_),
    .Y(_866_)
);

NAND2X1 _7346_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [0]),
    .B(gnd),
    .Y(_867_)
);

INVX1 _7347_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_867_),
    .Y(_868_)
);

AND2X2 _7348_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1]_5_bF$buf3 ),
    .Y(_869_)
);

NAND2X1 _7349_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1497_),
    .B(_869_),
    .Y(_870_)
);

INVX2 _7350_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1]_5_bF$buf2 ),
    .Y(_871_)
);

NAND2X1 _7351_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [1]),
    .B(gnd),
    .Y(_872_)
);

OAI21X1 _7352_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1575_),
    .B(_871_),
    .C(_872_),
    .Y(_873_)
);

NAND3X1 _7353_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_873_),
    .B(_868_),
    .C(_870_),
    .Y(_874_)
);

NAND3X1 _7354_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1]_5_bF$buf1 ),
    .C(_872_),
    .Y(_875_)
);

NAND2X1 _7355_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1]_5_bF$buf0 ),
    .Y(_876_)
);

NAND3X1 _7356_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [1]),
    .B(gnd),
    .C(_876_),
    .Y(_877_)
);

NAND3X1 _7357_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_867_),
    .B(_875_),
    .C(_877_),
    .Y(_878_)
);

AND2X2 _7358_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_874_),
    .B(_878_),
    .Y(_879_)
);

NAND2X1 _7359_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [2]),
    .Y(_880_)
);

OAI22X1 _7360_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1528_),
    .B(_880_),
    .C(_830_),
    .D(_835_),
    .Y(_881_)
);

NAND2X1 _7361_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1] [4]),
    .Y(_882_)
);

INVX1 _7362_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_882_),
    .Y(_883_)
);

AND2X2 _7363_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [3]),
    .Y(_884_)
);

NAND2X1 _7364_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_833_),
    .B(_884_),
    .Y(_885_)
);

INVX1 _7365_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .Y(_886_)
);

OAI21X1 _7366_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886_),
    .B(_812_),
    .C(_880_),
    .Y(_887_)
);

NAND3X1 _7367_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_883_),
    .B(_887_),
    .C(_885_),
    .Y(_888_)
);

NAND3X1 _7368_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [3]),
    .C(_880_),
    .Y(_889_)
);

NAND2X1 _7369_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [3]),
    .Y(_890_)
);

NAND3X1 _7370_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [2]),
    .C(_890_),
    .Y(_891_)
);

NAND3X1 _7371_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_882_),
    .B(_889_),
    .C(_891_),
    .Y(_892_)
);

NAND3X1 _7372_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_881_),
    .B(_892_),
    .C(_888_),
    .Y(_893_)
);

INVX1 _7373_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_881_),
    .Y(_894_)
);

AOI21X1 _7374_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_889_),
    .B(_891_),
    .C(_882_),
    .Y(_895_)
);

AOI22X1 _7375_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1] [4]),
    .C(_885_),
    .D(_887_),
    .Y(_896_)
);

OAI21X1 _7376_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_895_),
    .B(_896_),
    .C(_894_),
    .Y(_897_)
);

NAND3X1 _7377_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_893_),
    .B(_879_),
    .C(_897_),
    .Y(_898_)
);

NAND2X1 _7378_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_878_),
    .B(_874_),
    .Y(_899_)
);

OAI21X1 _7379_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_895_),
    .B(_896_),
    .C(_881_),
    .Y(_900_)
);

NAND3X1 _7380_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_892_),
    .B(_888_),
    .C(_894_),
    .Y(_901_)
);

NAND3X1 _7381_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_899_),
    .B(_901_),
    .C(_900_),
    .Y(_902_)
);

NAND3X1 _7382_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_898_),
    .B(_902_),
    .C(_866_),
    .Y(_903_)
);

AOI21X1 _7383_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_825_),
    .B(_845_),
    .C(_859_),
    .Y(_904_)
);

AOI21X1 _7384_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_900_),
    .B(_901_),
    .C(_899_),
    .Y(_905_)
);

AOI21X1 _7385_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_897_),
    .B(_893_),
    .C(_879_),
    .Y(_906_)
);

OAI21X1 _7386_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_905_),
    .B(_906_),
    .C(_904_),
    .Y(_907_)
);

NAND3X1 _7387_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_823_),
    .B(_903_),
    .C(_907_),
    .Y(_908_)
);

INVX1 _7388_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_823_),
    .Y(_909_)
);

OAI21X1 _7389_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_905_),
    .B(_906_),
    .C(_866_),
    .Y(_910_)
);

NAND3X1 _7390_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_898_),
    .B(_902_),
    .C(_904_),
    .Y(_911_)
);

NAND3X1 _7391_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_909_),
    .B(_910_),
    .C(_911_),
    .Y(_912_)
);

NAND3X1 _7392_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_850_),
    .B(_908_),
    .C(_912_),
    .Y(_913_)
);

NAND3X1 _7393_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_909_),
    .B(_903_),
    .C(_907_),
    .Y(_914_)
);

NAND3X1 _7394_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_823_),
    .B(_910_),
    .C(_911_),
    .Y(_915_)
);

NAND3X1 _7395_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_851_),
    .B(_914_),
    .C(_915_),
    .Y(_916_)
);

NAND3X1 _7396_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_913_),
    .B(_916_),
    .C(_865_),
    .Y(_917_)
);

INVX1 _7397_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_817_),
    .Y(_918_)
);

NAND3X1 _7398_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_918_),
    .B(_851_),
    .C(_854_),
    .Y(_919_)
);

NAND3X1 _7399_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_851_),
    .B(_908_),
    .C(_912_),
    .Y(_920_)
);

NAND3X1 _7400_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_850_),
    .B(_914_),
    .C(_915_),
    .Y(_921_)
);

NAND3X1 _7401_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_920_),
    .B(_921_),
    .C(_919_),
    .Y(_922_)
);

NAND3X1 _7402_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_917_),
    .B(_922_),
    .C(_864_),
    .Y(_923_)
);

INVX1 _7403_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_864_),
    .Y(_924_)
);

INVX1 _7404_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_917_),
    .Y(_925_)
);

INVX1 _7405_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_922_),
    .Y(_926_)
);

OAI21X1 _7406_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_925_),
    .B(_926_),
    .C(_924_),
    .Y(_927_)
);

AND2X2 _7407_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_927_),
    .B(_923_),
    .Y(_1593_[5])
);

AND2X2 _7408_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [0]),
    .B(gnd),
    .Y(_928_)
);

NAND2X1 _7409_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1]_5_bF$buf3 ),
    .Y(_929_)
);

OAI21X1 _7410_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1507_),
    .B(_929_),
    .C(_874_),
    .Y(_930_)
);

OR2X2 _7411_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_930_),
    .B(_928_),
    .Y(_931_)
);

NAND2X1 _7412_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_928_),
    .B(_930_),
    .Y(_932_)
);

NAND2X1 _7413_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_932_),
    .B(_931_),
    .Y(_933_)
);

AOI21X1 _7414_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_888_),
    .B(_892_),
    .C(_881_),
    .Y(_934_)
);

OAI21X1 _7415_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_899_),
    .B(_934_),
    .C(_893_),
    .Y(_935_)
);

NAND2X1 _7416_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [1]),
    .B(gnd),
    .Y(_936_)
);

INVX1 _7417_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_936_),
    .Y(_937_)
);

AND2X2 _7418_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [2]),
    .B(gnd),
    .Y(_938_)
);

AND2X2 _7419_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1] [6]),
    .Y(_939_)
);

NAND2X1 _7420_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_938_),
    .B(_939_),
    .Y(_940_)
);

INVX2 _7421_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [6]),
    .Y(_941_)
);

NAND2X1 _7422_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [2]),
    .B(gnd),
    .Y(_942_)
);

OAI21X1 _7423_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1575_),
    .B(_941_),
    .C(_942_),
    .Y(_943_)
);

NAND3X1 _7424_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_943_),
    .B(_937_),
    .C(_940_),
    .Y(_944_)
);

NAND3X1 _7425_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1] [6]),
    .C(_942_),
    .Y(_945_)
);

NAND2X1 _7426_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1] [6]),
    .Y(_946_)
);

NAND2X1 _7427_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_946_),
    .B(_938_),
    .Y(_947_)
);

NAND3X1 _7428_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_936_),
    .B(_945_),
    .C(_947_),
    .Y(_948_)
);

AND2X2 _7429_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_944_),
    .B(_948_),
    .Y(_949_)
);

NAND2X1 _7430_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [3]),
    .Y(_950_)
);

AOI22X1 _7431_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [2]),
    .C(vdd),
    .D(\X[1] [3]),
    .Y(_951_)
);

OAI22X1 _7432_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_839_),
    .B(_950_),
    .C(_882_),
    .D(_951_),
    .Y(_952_)
);

NAND2X1 _7433_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1]_5_bF$buf2 ),
    .Y(_953_)
);

INVX1 _7434_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_953_),
    .Y(_954_)
);

AND2X2 _7435_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [4]),
    .Y(_955_)
);

NAND2X1 _7436_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_884_),
    .B(_955_),
    .Y(_956_)
);

AOI22X1 _7437_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [3]),
    .C(vdd),
    .D(\X[1] [4]),
    .Y(_957_)
);

INVX1 _7438_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_957_),
    .Y(_958_)
);

NAND3X1 _7439_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_954_),
    .B(_958_),
    .C(_956_),
    .Y(_959_)
);

NAND3X1 _7440_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [4]),
    .C(_950_),
    .Y(_960_)
);

NAND2X1 _7441_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [4]),
    .Y(_961_)
);

NAND3X1 _7442_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [3]),
    .C(_961_),
    .Y(_962_)
);

NAND3X1 _7443_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_953_),
    .B(_960_),
    .C(_962_),
    .Y(_963_)
);

NAND3X1 _7444_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_952_),
    .B(_963_),
    .C(_959_),
    .Y(_964_)
);

INVX1 _7445_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_952_),
    .Y(_965_)
);

AOI21X1 _7446_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_960_),
    .B(_962_),
    .C(_953_),
    .Y(_966_)
);

AOI22X1 _7447_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1]_5_bF$buf1 ),
    .C(_956_),
    .D(_958_),
    .Y(_967_)
);

OAI21X1 _7448_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_966_),
    .B(_967_),
    .C(_965_),
    .Y(_968_)
);

NAND3X1 _7449_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_964_),
    .B(_949_),
    .C(_968_),
    .Y(_969_)
);

NAND2X1 _7450_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_948_),
    .B(_944_),
    .Y(_970_)
);

OAI21X1 _7451_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_966_),
    .B(_967_),
    .C(_952_),
    .Y(_971_)
);

NAND3X1 _7452_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_959_),
    .B(_963_),
    .C(_965_),
    .Y(_972_)
);

NAND3X1 _7453_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_970_),
    .B(_972_),
    .C(_971_),
    .Y(_973_)
);

NAND3X1 _7454_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_969_),
    .B(_935_),
    .C(_973_),
    .Y(_974_)
);

INVX1 _7455_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_893_),
    .Y(_975_)
);

AOI21X1 _7456_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_879_),
    .B(_897_),
    .C(_975_),
    .Y(_976_)
);

AOI21X1 _7457_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_971_),
    .B(_972_),
    .C(_970_),
    .Y(_977_)
);

AOI21X1 _7458_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_968_),
    .B(_964_),
    .C(_949_),
    .Y(_978_)
);

OAI21X1 _7459_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_977_),
    .B(_978_),
    .C(_976_),
    .Y(_979_)
);

NAND3X1 _7460_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_933_),
    .B(_974_),
    .C(_979_),
    .Y(_980_)
);

AND2X2 _7461_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931_),
    .B(_932_),
    .Y(_981_)
);

OAI21X1 _7462_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_977_),
    .B(_978_),
    .C(_935_),
    .Y(_982_)
);

NAND3X1 _7463_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_969_),
    .B(_973_),
    .C(_976_),
    .Y(_983_)
);

NAND3X1 _7464_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_981_),
    .B(_982_),
    .C(_983_),
    .Y(_984_)
);

AOI22X1 _7465_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_908_),
    .B(_903_),
    .C(_980_),
    .D(_984_),
    .Y(_985_)
);

AOI21X1 _7466_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_898_),
    .B(_902_),
    .C(_866_),
    .Y(_986_)
);

OAI21X1 _7467_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_909_),
    .B(_986_),
    .C(_903_),
    .Y(_987_)
);

NAND3X1 _7468_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_981_),
    .B(_974_),
    .C(_979_),
    .Y(_988_)
);

NAND3X1 _7469_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_933_),
    .B(_982_),
    .C(_983_),
    .Y(_989_)
);

AOI21X1 _7470_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_989_),
    .B(_988_),
    .C(_987_),
    .Y(_990_)
);

OAI21X1 _7471_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_990_),
    .B(_985_),
    .C(_913_),
    .Y(_991_)
);

AOI21X1 _7472_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_915_),
    .B(_914_),
    .C(_851_),
    .Y(_992_)
);

NAND3X1 _7473_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_987_),
    .B(_988_),
    .C(_989_),
    .Y(_993_)
);

INVX1 _7474_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_903_),
    .Y(_994_)
);

AOI21X1 _7475_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_823_),
    .B(_907_),
    .C(_994_),
    .Y(_995_)
);

AOI21X1 _7476_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_983_),
    .B(_982_),
    .C(_933_),
    .Y(_996_)
);

AOI21X1 _7477_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_979_),
    .B(_974_),
    .C(_981_),
    .Y(_997_)
);

OAI21X1 _7478_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_996_),
    .B(_997_),
    .C(_995_),
    .Y(_998_)
);

NAND3X1 _7479_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_992_),
    .B(_993_),
    .C(_998_),
    .Y(_999_)
);

NAND2X1 _7480_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_999_),
    .B(_991_),
    .Y(_1000_)
);

AOI21X1 _7481_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_917_),
    .B(_923_),
    .C(_1000_),
    .Y(_1001_)
);

OAI21X1 _7482_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_926_),
    .B(_924_),
    .C(_917_),
    .Y(_1002_)
);

AOI21X1 _7483_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_991_),
    .B(_999_),
    .C(_1002_),
    .Y(_1003_)
);

NOR2X1 _7484_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1001_),
    .B(_1003_),
    .Y(_1593_[6])
);

INVX1 _7485_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_999_),
    .Y(_1004_)
);

AOI21X1 _7486_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_969_),
    .B(_973_),
    .C(_935_),
    .Y(_1005_)
);

OAI21X1 _7487_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_933_),
    .B(_1005_),
    .C(_974_),
    .Y(_1006_)
);

NAND2X1 _7488_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [0]),
    .B(gnd),
    .Y(_1007_)
);

INVX1 _7489_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1007_),
    .Y(_1008_)
);

NAND2X1 _7490_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [1]),
    .B(gnd),
    .Y(_1009_)
);

INVX1 _7491_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1009_),
    .Y(_1010_)
);

AND2X2 _7492_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_942_),
    .B(_946_),
    .Y(_1011_)
);

OAI21X1 _7493_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_936_),
    .B(_1011_),
    .C(_940_),
    .Y(_1012_)
);

NAND2X1 _7494_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1010_),
    .B(_1012_),
    .Y(_1013_)
);

NAND3X1 _7495_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_940_),
    .B(_1009_),
    .C(_944_),
    .Y(_1014_)
);

NAND3X1 _7496_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1008_),
    .B(_1014_),
    .C(_1013_),
    .Y(_1015_)
);

AOI21X1 _7497_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_944_),
    .B(_940_),
    .C(_1009_),
    .Y(_1016_)
);

NOR2X1 _7498_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1010_),
    .B(_1012_),
    .Y(_1017_)
);

OAI21X1 _7499_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1016_),
    .B(_1017_),
    .C(_1007_),
    .Y(_1018_)
);

NAND2X1 _7500_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1015_),
    .B(_1018_),
    .Y(_1019_)
);

AOI21X1 _7501_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_959_),
    .B(_963_),
    .C(_952_),
    .Y(_1020_)
);

OAI21X1 _7502_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_970_),
    .B(_1020_),
    .C(_964_),
    .Y(_1021_)
);

NAND2X1 _7503_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [2]),
    .B(gnd),
    .Y(_1022_)
);

INVX1 _7504_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1022_),
    .Y(_1023_)
);

AND2X2 _7505_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [3]),
    .B(gnd),
    .Y(_1024_)
);

AND2X2 _7506_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1] [7]),
    .Y(_1025_)
);

NAND2X1 _7507_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1024_),
    .B(_1025_),
    .Y(_1026_)
);

AOI22X1 _7508_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1] [7]),
    .C(\X[1] [3]),
    .D(gnd),
    .Y(_1027_)
);

INVX1 _7509_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1027_),
    .Y(_1028_)
);

NAND3X1 _7510_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1023_),
    .B(_1028_),
    .C(_1026_),
    .Y(_1029_)
);

INVX1 _7511_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_1030_)
);

OAI21X1 _7512_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_812_),
    .B(_1030_),
    .C(_1025_),
    .Y(_1031_)
);

INVX1 _7513_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [7]),
    .Y(_1032_)
);

OAI21X1 _7514_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1575_),
    .B(_1032_),
    .C(_1024_),
    .Y(_1033_)
);

NAND3X1 _7515_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1022_),
    .B(_1031_),
    .C(_1033_),
    .Y(_1034_)
);

NAND2X1 _7516_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1029_),
    .B(_1034_),
    .Y(_1035_)
);

OAI21X1 _7517_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_953_),
    .B(_957_),
    .C(_956_),
    .Y(_1036_)
);

NAND2X1 _7518_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1] [6]),
    .Y(_1037_)
);

NAND2X1 _7519_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [4]),
    .Y(_1038_)
);

AND2X2 _7520_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1]_5_bF$buf0 ),
    .Y(_1039_)
);

NAND2X1 _7521_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1038_),
    .B(_1039_),
    .Y(_1040_)
);

OAI21X1 _7522_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886_),
    .B(_871_),
    .C(_955_),
    .Y(_1041_)
);

AOI21X1 _7523_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1041_),
    .B(_1040_),
    .C(_1037_),
    .Y(_1042_)
);

INVX1 _7524_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1037_),
    .Y(_1043_)
);

NAND2X1 _7525_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_955_),
    .B(_1039_),
    .Y(_1044_)
);

AOI22X1 _7526_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [4]),
    .C(vdd),
    .D(\X[1]_5_bF$buf3 ),
    .Y(_1045_)
);

INVX1 _7527_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1045_),
    .Y(_1046_)
);

AOI21X1 _7528_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1044_),
    .B(_1046_),
    .C(_1043_),
    .Y(_1047_)
);

OAI21X1 _7529_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1047_),
    .B(_1042_),
    .C(_1036_),
    .Y(_1048_)
);

AOI22X1 _7530_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_884_),
    .B(_955_),
    .C(_958_),
    .D(_954_),
    .Y(_1049_)
);

NAND3X1 _7531_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1043_),
    .B(_1046_),
    .C(_1044_),
    .Y(_1050_)
);

NAND2X1 _7532_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1]_5_bF$buf2 ),
    .Y(_1051_)
);

NOR2X1 _7533_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1038_),
    .B(_1051_),
    .Y(_1052_)
);

OAI21X1 _7534_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1045_),
    .B(_1052_),
    .C(_1037_),
    .Y(_1053_)
);

NAND3X1 _7535_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1050_),
    .B(_1049_),
    .C(_1053_),
    .Y(_1054_)
);

AOI21X1 _7536_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1048_),
    .B(_1054_),
    .C(_1035_),
    .Y(_1055_)
);

AND2X2 _7537_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1034_),
    .B(_1029_),
    .Y(_1056_)
);

NAND3X1 _7538_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1036_),
    .B(_1050_),
    .C(_1053_),
    .Y(_1057_)
);

OAI21X1 _7539_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1047_),
    .B(_1042_),
    .C(_1049_),
    .Y(_1058_)
);

AOI21X1 _7540_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1058_),
    .B(_1057_),
    .C(_1056_),
    .Y(_1059_)
);

OAI21X1 _7541_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1055_),
    .B(_1059_),
    .C(_1021_),
    .Y(_1060_)
);

INVX1 _7542_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_964_),
    .Y(_1061_)
);

AOI21X1 _7543_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_949_),
    .B(_968_),
    .C(_1061_),
    .Y(_1062_)
);

NAND3X1 _7544_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1057_),
    .B(_1056_),
    .C(_1058_),
    .Y(_1063_)
);

NAND3X1 _7545_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1035_),
    .B(_1054_),
    .C(_1048_),
    .Y(_1064_)
);

NAND3X1 _7546_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1063_),
    .B(_1064_),
    .C(_1062_),
    .Y(_1065_)
);

AOI21X1 _7547_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1065_),
    .B(_1060_),
    .C(_1019_),
    .Y(_1066_)
);

AND2X2 _7548_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1018_),
    .B(_1015_),
    .Y(_1067_)
);

NAND3X1 _7549_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1021_),
    .B(_1063_),
    .C(_1064_),
    .Y(_1068_)
);

OAI21X1 _7550_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1055_),
    .B(_1059_),
    .C(_1062_),
    .Y(_1069_)
);

AOI21X1 _7551_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1069_),
    .B(_1068_),
    .C(_1067_),
    .Y(_1070_)
);

OAI21X1 _7552_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1070_),
    .B(_1066_),
    .C(_1006_),
    .Y(_1071_)
);

INVX1 _7553_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_974_),
    .Y(_1072_)
);

AOI21X1 _7554_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_981_),
    .B(_979_),
    .C(_1072_),
    .Y(_1073_)
);

NAND3X1 _7555_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1068_),
    .B(_1067_),
    .C(_1069_),
    .Y(_1074_)
);

NAND3X1 _7556_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1019_),
    .B(_1060_),
    .C(_1065_),
    .Y(_1075_)
);

NAND3X1 _7557_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1074_),
    .B(_1075_),
    .C(_1073_),
    .Y(_1076_)
);

AOI21X1 _7558_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1076_),
    .B(_1071_),
    .C(_932_),
    .Y(_1077_)
);

INVX1 _7559_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_932_),
    .Y(_1078_)
);

NAND3X1 _7560_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1006_),
    .B(_1074_),
    .C(_1075_),
    .Y(_1079_)
);

OAI21X1 _7561_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1066_),
    .B(_1070_),
    .C(_1073_),
    .Y(_1080_)
);

AOI21X1 _7562_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1080_),
    .B(_1079_),
    .C(_1078_),
    .Y(_1081_)
);

OAI21X1 _7563_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1081_),
    .B(_1077_),
    .C(_993_),
    .Y(_1082_)
);

NAND3X1 _7564_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1078_),
    .B(_1079_),
    .C(_1080_),
    .Y(_1083_)
);

NAND3X1 _7565_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_932_),
    .B(_1071_),
    .C(_1076_),
    .Y(_1084_)
);

NAND3X1 _7566_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_985_),
    .B(_1083_),
    .C(_1084_),
    .Y(_1085_)
);

AND2X2 _7567_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1082_),
    .B(_1085_),
    .Y(_1086_)
);

OAI21X1 _7568_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1004_),
    .B(_1001_),
    .C(_1086_),
    .Y(_1087_)
);

NOR2X1 _7569_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1004_),
    .B(_1001_),
    .Y(_1088_)
);

AOI21X1 _7570_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1084_),
    .B(_1083_),
    .C(_985_),
    .Y(_1089_)
);

INVX1 _7571_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1085_),
    .Y(_1090_)
);

OAI21X1 _7572_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1089_),
    .B(_1090_),
    .C(_1088_),
    .Y(_1091_)
);

AND2X2 _7573_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1091_),
    .B(_1087_),
    .Y(_1593_[7])
);

NAND3X1 _7574_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1082_),
    .B(_1085_),
    .C(_1001_),
    .Y(_1092_)
);

AOI21X1 _7575_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1004_),
    .B(_1082_),
    .C(_1090_),
    .Y(_1093_)
);

NAND2X1 _7576_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1093_),
    .B(_1092_),
    .Y(_1094_)
);

INVX1 _7577_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1079_),
    .Y(_1095_)
);

AOI21X1 _7578_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1078_),
    .B(_1080_),
    .C(_1095_),
    .Y(_1096_)
);

OAI21X1 _7579_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1007_),
    .B(_1017_),
    .C(_1013_),
    .Y(_1097_)
);

INVX1 _7580_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1097_),
    .Y(_1098_)
);

AOI21X1 _7581_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1063_),
    .B(_1064_),
    .C(_1021_),
    .Y(_1099_)
);

OAI21X1 _7582_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1019_),
    .B(_1099_),
    .C(_1068_),
    .Y(_1100_)
);

NAND2X1 _7583_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [1]),
    .B(gnd),
    .Y(_1101_)
);

INVX2 _7584_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_1102_)
);

NOR2X1 _7585_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1567_),
    .B(_1102_),
    .Y(_1103_)
);

OAI21X1 _7586_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1022_),
    .B(_1027_),
    .C(_1026_),
    .Y(_1104_)
);

NOR2X1 _7587_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1103_),
    .B(_1104_),
    .Y(_1105_)
);

AND2X2 _7588_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1104_),
    .B(_1103_),
    .Y(_1106_)
);

OAI21X1 _7589_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1105_),
    .B(_1106_),
    .C(_1101_),
    .Y(_1107_)
);

INVX1 _7590_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1101_),
    .Y(_1108_)
);

OR2X2 _7591_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1104_),
    .B(_1103_),
    .Y(_1109_)
);

NAND2X1 _7592_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1103_),
    .B(_1104_),
    .Y(_1110_)
);

NAND3X1 _7593_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1108_),
    .B(_1110_),
    .C(_1109_),
    .Y(_1111_)
);

NAND2X1 _7594_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1107_),
    .B(_1111_),
    .Y(_1112_)
);

AOI21X1 _7595_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1053_),
    .B(_1050_),
    .C(_1036_),
    .Y(_1113_)
);

OAI21X1 _7596_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1035_),
    .B(_1113_),
    .C(_1057_),
    .Y(_1114_)
);

NAND2X1 _7597_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [3]),
    .B(gnd),
    .Y(_1115_)
);

INVX1 _7598_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_1116_)
);

OAI21X1 _7599_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_812_),
    .B(_1116_),
    .C(_822_),
    .Y(_1117_)
);

NAND2X1 _7600_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [4]),
    .B(gnd),
    .Y(_1118_)
);

OAI21X1 _7601_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1115_),
    .B(_1118_),
    .C(_1117_),
    .Y(_1119_)
);

OAI21X1 _7602_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1037_),
    .B(_1045_),
    .C(_1044_),
    .Y(_1120_)
);

NAND2X1 _7603_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1] [7]),
    .Y(_1121_)
);

NAND2X1 _7604_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1]_5_bF$buf1 ),
    .Y(_1122_)
);

NAND3X1 _7605_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [6]),
    .C(_1122_),
    .Y(_1123_)
);

AND2X2 _7606_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1]_5_bF$buf0 ),
    .Y(_1124_)
);

OAI21X1 _7607_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886_),
    .B(_941_),
    .C(_1124_),
    .Y(_1125_)
);

AOI21X1 _7608_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1125_),
    .B(_1123_),
    .C(_1121_),
    .Y(_1126_)
);

INVX1 _7609_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1121_),
    .Y(_1127_)
);

AND2X2 _7610_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [6]),
    .Y(_1128_)
);

NAND2X1 _7611_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1124_),
    .B(_1128_),
    .Y(_1129_)
);

NAND2X1 _7612_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [6]),
    .Y(_1130_)
);

NAND2X1 _7613_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1122_),
    .B(_1130_),
    .Y(_1131_)
);

AOI21X1 _7614_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1129_),
    .B(_1131_),
    .C(_1127_),
    .Y(_1132_)
);

OAI21X1 _7615_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1132_),
    .B(_1126_),
    .C(_1120_),
    .Y(_1133_)
);

AOI21X1 _7616_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1043_),
    .B(_1046_),
    .C(_1052_),
    .Y(_1134_)
);

NAND3X1 _7617_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1127_),
    .B(_1131_),
    .C(_1129_),
    .Y(_1135_)
);

NAND3X1 _7618_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1121_),
    .B(_1123_),
    .C(_1125_),
    .Y(_1136_)
);

NAND3X1 _7619_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1135_),
    .B(_1136_),
    .C(_1134_),
    .Y(_1137_)
);

AOI21X1 _7620_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1133_),
    .B(_1137_),
    .C(_1119_),
    .Y(_1138_)
);

INVX1 _7621_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1119_),
    .Y(_1139_)
);

NAND3X1 _7622_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1120_),
    .B(_1135_),
    .C(_1136_),
    .Y(_1140_)
);

OAI21X1 _7623_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1132_),
    .B(_1126_),
    .C(_1134_),
    .Y(_1141_)
);

AOI21X1 _7624_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1141_),
    .B(_1140_),
    .C(_1139_),
    .Y(_1142_)
);

OAI21X1 _7625_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1138_),
    .B(_1142_),
    .C(_1114_),
    .Y(_1143_)
);

INVX1 _7626_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1057_),
    .Y(_1144_)
);

AOI21X1 _7627_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1056_),
    .B(_1058_),
    .C(_1144_),
    .Y(_1145_)
);

NAND3X1 _7628_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1139_),
    .B(_1140_),
    .C(_1141_),
    .Y(_1146_)
);

NAND3X1 _7629_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1119_),
    .B(_1137_),
    .C(_1133_),
    .Y(_1147_)
);

NAND3X1 _7630_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1146_),
    .B(_1147_),
    .C(_1145_),
    .Y(_1148_)
);

AOI21X1 _7631_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1148_),
    .B(_1143_),
    .C(_1112_),
    .Y(_1149_)
);

AND2X2 _7632_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1111_),
    .B(_1107_),
    .Y(_1150_)
);

NAND3X1 _7633_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1146_),
    .B(_1147_),
    .C(_1114_),
    .Y(_1151_)
);

OAI21X1 _7634_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1138_),
    .B(_1142_),
    .C(_1145_),
    .Y(_1152_)
);

AOI21X1 _7635_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1152_),
    .B(_1151_),
    .C(_1150_),
    .Y(_1153_)
);

OAI21X1 _7636_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1153_),
    .B(_1149_),
    .C(_1100_),
    .Y(_1154_)
);

INVX1 _7637_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1068_),
    .Y(_1155_)
);

AOI21X1 _7638_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1067_),
    .B(_1069_),
    .C(_1155_),
    .Y(_1156_)
);

NAND3X1 _7639_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1150_),
    .B(_1151_),
    .C(_1152_),
    .Y(_1157_)
);

NAND3X1 _7640_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1112_),
    .B(_1143_),
    .C(_1148_),
    .Y(_1158_)
);

NAND3X1 _7641_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1157_),
    .B(_1158_),
    .C(_1156_),
    .Y(_1159_)
);

AOI21X1 _7642_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1154_),
    .B(_1159_),
    .C(_1098_),
    .Y(_1160_)
);

NAND3X1 _7643_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1100_),
    .B(_1157_),
    .C(_1158_),
    .Y(_1161_)
);

OAI21X1 _7644_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1153_),
    .B(_1149_),
    .C(_1156_),
    .Y(_1162_)
);

AOI21X1 _7645_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1162_),
    .B(_1161_),
    .C(_1097_),
    .Y(_1163_)
);

OAI21X1 _7646_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1163_),
    .B(_1160_),
    .C(_1096_),
    .Y(_1164_)
);

AOI21X1 _7647_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1075_),
    .B(_1074_),
    .C(_1006_),
    .Y(_1165_)
);

OAI21X1 _7648_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_932_),
    .B(_1165_),
    .C(_1079_),
    .Y(_1166_)
);

NAND3X1 _7649_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1097_),
    .B(_1161_),
    .C(_1162_),
    .Y(_1167_)
);

NAND3X1 _7650_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1098_),
    .B(_1159_),
    .C(_1154_),
    .Y(_1168_)
);

NAND3X1 _7651_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1166_),
    .B(_1167_),
    .C(_1168_),
    .Y(_1169_)
);

NAND2X1 _7652_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1169_),
    .B(_1164_),
    .Y(_1170_)
);

NAND2X1 _7653_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1170_),
    .B(_1094_),
    .Y(_1171_)
);

OAI21X1 _7654_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_999_),
    .B(_1089_),
    .C(_1085_),
    .Y(_1172_)
);

AOI21X1 _7655_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1086_),
    .B(_1001_),
    .C(_1172_),
    .Y(_1173_)
);

AND2X2 _7656_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1164_),
    .B(_1169_),
    .Y(_1174_)
);

NAND2X1 _7657_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1174_),
    .B(_1173_),
    .Y(_1175_)
);

NAND2X1 _7658_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1171_),
    .B(_1175_),
    .Y(_1593_[8])
);

INVX1 _7659_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1169_),
    .Y(_1176_)
);

AOI21X1 _7660_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1094_),
    .B(_1164_),
    .C(_1176_),
    .Y(_1177_)
);

AOI21X1 _7661_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1158_),
    .B(_1157_),
    .C(_1100_),
    .Y(_1178_)
);

OAI21X1 _7662_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1098_),
    .B(_1178_),
    .C(_1161_),
    .Y(_1179_)
);

OAI21X1 _7663_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1101_),
    .B(_1105_),
    .C(_1110_),
    .Y(_1180_)
);

AOI21X1 _7664_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1146_),
    .B(_1147_),
    .C(_1114_),
    .Y(_1181_)
);

OAI21X1 _7665_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1112_),
    .B(_1181_),
    .C(_1151_),
    .Y(_1182_)
);

NAND2X1 _7666_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [2]),
    .B(gnd),
    .Y(_1183_)
);

NOR2X1 _7667_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1115_),
    .B(_1118_),
    .Y(_1184_)
);

NAND2X1 _7668_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_1184_),
    .Y(_1185_)
);

INVX1 _7669_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1185_),
    .Y(_1186_)
);

AOI21X1 _7670_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [3]),
    .B(gnd),
    .C(_1184_),
    .Y(_1187_)
);

OAI21X1 _7671_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1187_),
    .B(_1186_),
    .C(_1183_),
    .Y(_1188_)
);

INVX1 _7672_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1183_),
    .Y(_1189_)
);

INVX1 _7673_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1187_),
    .Y(_1190_)
);

NAND3X1 _7674_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1189_),
    .B(_1185_),
    .C(_1190_),
    .Y(_1191_)
);

AND2X2 _7675_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1191_),
    .B(_1188_),
    .Y(_1192_)
);

AOI21X1 _7676_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1136_),
    .B(_1135_),
    .C(_1120_),
    .Y(_1193_)
);

OAI21X1 _7677_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1119_),
    .B(_1193_),
    .C(_1140_),
    .Y(_1194_)
);

NOR2X1 _7678_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_929_),
    .B(_1118_),
    .Y(_1195_)
);

AND2X2 _7679_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_929_),
    .B(_1118_),
    .Y(_1196_)
);

NOR2X1 _7680_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1195_),
    .B(_1196_),
    .Y(_1197_)
);

NAND2X1 _7681_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [6]),
    .Y(_1198_)
);

AOI22X1 _7682_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1]_5_bF$buf3 ),
    .C(vdd),
    .D(\X[1] [6]),
    .Y(_1199_)
);

OAI22X1 _7683_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1051_),
    .B(_1198_),
    .C(_1121_),
    .D(_1199_),
    .Y(_1200_)
);

AOI22X1 _7684_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [6]),
    .C(vdd),
    .D(\X[1] [7]),
    .Y(_1201_)
);

AND2X2 _7685_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [7]),
    .Y(_1202_)
);

AOI21X1 _7686_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1128_),
    .B(_1202_),
    .C(_1201_),
    .Y(_1203_)
);

NAND2X1 _7687_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1203_),
    .B(_1200_),
    .Y(_1204_)
);

AND2X2 _7688_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [6]),
    .Y(_1205_)
);

AOI22X1 _7689_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1039_),
    .B(_1205_),
    .C(_1131_),
    .D(_1127_),
    .Y(_1206_)
);

NAND2X1 _7690_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [7]),
    .Y(_1207_)
);

NAND2X1 _7691_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1198_),
    .B(_1207_),
    .Y(_1208_)
);

NAND2X1 _7692_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [7]),
    .Y(_1209_)
);

OAI21X1 _7693_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1130_),
    .B(_1209_),
    .C(_1208_),
    .Y(_1210_)
);

NAND2X1 _7694_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1210_),
    .B(_1206_),
    .Y(_1211_)
);

NAND3X1 _7695_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1197_),
    .B(_1204_),
    .C(_1211_),
    .Y(_1212_)
);

NAND2X1 _7696_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1]_5_bF$buf2 ),
    .B(gnd),
    .Y(_1213_)
);

INVX1 _7697_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [4]),
    .Y(_1214_)
);

OAI21X1 _7698_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1214_),
    .B(_1116_),
    .C(_929_),
    .Y(_1215_)
);

OAI21X1 _7699_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_822_),
    .B(_1213_),
    .C(_1215_),
    .Y(_1216_)
);

NAND2X1 _7700_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1200_),
    .B(_1210_),
    .Y(_1217_)
);

NAND2X1 _7701_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1203_),
    .B(_1206_),
    .Y(_1218_)
);

NAND3X1 _7702_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1216_),
    .B(_1217_),
    .C(_1218_),
    .Y(_1219_)
);

NAND3X1 _7703_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1212_),
    .B(_1219_),
    .C(_1194_),
    .Y(_1220_)
);

NAND2X1 _7704_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1212_),
    .B(_1219_),
    .Y(_1221_)
);

NAND3X1 _7705_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1140_),
    .B(_1146_),
    .C(_1221_),
    .Y(_1222_)
);

NAND3X1 _7706_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1192_),
    .B(_1220_),
    .C(_1222_),
    .Y(_1223_)
);

NAND2X1 _7707_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1188_),
    .B(_1191_),
    .Y(_1224_)
);

AOI21X1 _7708_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1140_),
    .B(_1146_),
    .C(_1221_),
    .Y(_1225_)
);

AOI21X1 _7709_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1212_),
    .B(_1219_),
    .C(_1194_),
    .Y(_1226_)
);

OAI21X1 _7710_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1226_),
    .B(_1225_),
    .C(_1224_),
    .Y(_1227_)
);

NAND3X1 _7711_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1223_),
    .B(_1227_),
    .C(_1182_),
    .Y(_1228_)
);

INVX1 _7712_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1151_),
    .Y(_1229_)
);

AOI21X1 _7713_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1150_),
    .B(_1152_),
    .C(_1229_),
    .Y(_1230_)
);

INVX1 _7714_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1223_),
    .Y(_1231_)
);

AOI21X1 _7715_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1222_),
    .B(_1220_),
    .C(_1192_),
    .Y(_1232_)
);

OAI21X1 _7716_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1232_),
    .B(_1231_),
    .C(_1230_),
    .Y(_1233_)
);

NAND3X1 _7717_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1180_),
    .B(_1228_),
    .C(_1233_),
    .Y(_1234_)
);

INVX1 _7718_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1180_),
    .Y(_1235_)
);

INVX1 _7719_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1228_),
    .Y(_1236_)
);

AOI21X1 _7720_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1227_),
    .B(_1223_),
    .C(_1182_),
    .Y(_1237_)
);

OAI21X1 _7721_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1237_),
    .B(_1236_),
    .C(_1235_),
    .Y(_1238_)
);

NAND3X1 _7722_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1179_),
    .B(_1234_),
    .C(_1238_),
    .Y(_1239_)
);

INVX1 _7723_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1161_),
    .Y(_1240_)
);

AOI21X1 _7724_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1097_),
    .B(_1162_),
    .C(_1240_),
    .Y(_1241_)
);

OAI21X1 _7725_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1232_),
    .B(_1231_),
    .C(_1182_),
    .Y(_1242_)
);

NAND3X1 _7726_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1223_),
    .B(_1227_),
    .C(_1230_),
    .Y(_1243_)
);

AOI21X1 _7727_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1243_),
    .B(_1242_),
    .C(_1235_),
    .Y(_1244_)
);

AOI21X1 _7728_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1233_),
    .B(_1228_),
    .C(_1180_),
    .Y(_1245_)
);

OAI21X1 _7729_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1244_),
    .B(_1245_),
    .C(_1241_),
    .Y(_1246_)
);

AND2X2 _7730_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1246_),
    .B(_1239_),
    .Y(_1247_)
);

OR2X2 _7731_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1177_),
    .B(_1247_),
    .Y(_1248_)
);

NAND2X1 _7732_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1247_),
    .B(_1177_),
    .Y(_1249_)
);

NAND2X1 _7733_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1249_),
    .B(_1248_),
    .Y(_1593_[9])
);

NAND2X1 _7734_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1239_),
    .B(_1246_),
    .Y(_1250_)
);

NOR2X1 _7735_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1170_),
    .B(_1250_),
    .Y(_1251_)
);

NAND2X1 _7736_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1251_),
    .B(_1094_),
    .Y(_1252_)
);

AOI21X1 _7737_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1238_),
    .B(_1234_),
    .C(_1179_),
    .Y(_1253_)
);

AOI21X1 _7738_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1169_),
    .B(_1239_),
    .C(_1253_),
    .Y(_1254_)
);

INVX1 _7739_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1254_),
    .Y(_1255_)
);

OAI21X1 _7740_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1235_),
    .B(_1237_),
    .C(_1228_),
    .Y(_1256_)
);

OAI21X1 _7741_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1183_),
    .B(_1187_),
    .C(_1185_),
    .Y(_1257_)
);

OAI21X1 _7742_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1224_),
    .B(_1226_),
    .C(_1220_),
    .Y(_1258_)
);

INVX2 _7743_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_1259_)
);

NOR3X1 _7744_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1102_),
    .B(_929_),
    .C(_1118_),
    .Y(_1260_)
);

OAI22X1 _7745_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1214_),
    .B(_1102_),
    .C(_822_),
    .D(_1213_),
    .Y(_1261_)
);

INVX1 _7746_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1261_),
    .Y(_1262_)
);

OAI22X1 _7747_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_812_),
    .B(_1259_),
    .C(_1260_),
    .D(_1262_),
    .Y(_1263_)
);

NOR2X1 _7748_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_812_),
    .B(_1259_),
    .Y(_1264_)
);

NAND2X1 _7749_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_1195_),
    .Y(_1265_)
);

NAND3X1 _7750_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1264_),
    .B(_1261_),
    .C(_1265_),
    .Y(_1266_)
);

AND2X2 _7751_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1263_),
    .B(_1266_),
    .Y(_1267_)
);

NOR2X1 _7752_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1203_),
    .B(_1200_),
    .Y(_1268_)
);

OAI21X1 _7753_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1216_),
    .B(_1268_),
    .C(_1204_),
    .Y(_1269_)
);

NAND2X1 _7754_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1] [6]),
    .Y(_1270_)
);

NOR2X1 _7755_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1270_),
    .B(_1213_),
    .Y(_1271_)
);

AND2X2 _7756_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1270_),
    .B(_1213_),
    .Y(_1272_)
);

OAI22X1 _7757_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1128_),
    .B(_1209_),
    .C(_1271_),
    .D(_1272_),
    .Y(_1273_)
);

AND2X2 _7758_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1] [6]),
    .Y(_1274_)
);

AND2X2 _7759_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1]_5_bF$buf1 ),
    .B(gnd),
    .Y(_1275_)
);

NAND2X1 _7760_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1274_),
    .B(_1275_),
    .Y(_1276_)
);

OAI21X1 _7761_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_871_),
    .B(_1116_),
    .C(_1270_),
    .Y(_1277_)
);

AOI21X1 _7762_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[1] [6]),
    .C(_1209_),
    .Y(_1278_)
);

NAND3X1 _7763_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1277_),
    .B(_1278_),
    .C(_1276_),
    .Y(_1279_)
);

AND2X2 _7764_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1273_),
    .B(_1279_),
    .Y(_1280_)
);

NAND2X1 _7765_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1280_),
    .B(_1269_),
    .Y(_1281_)
);

NAND2X1 _7766_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1279_),
    .B(_1273_),
    .Y(_1282_)
);

NAND3X1 _7767_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1204_),
    .B(_1282_),
    .C(_1212_),
    .Y(_1283_)
);

NAND3X1 _7768_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1267_),
    .B(_1283_),
    .C(_1281_),
    .Y(_1284_)
);

NAND2X1 _7769_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1266_),
    .B(_1263_),
    .Y(_1285_)
);

NAND2X1 _7770_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1282_),
    .B(_1269_),
    .Y(_1286_)
);

NAND3X1 _7771_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1204_),
    .B(_1280_),
    .C(_1212_),
    .Y(_1287_)
);

NAND3X1 _7772_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1285_),
    .B(_1287_),
    .C(_1286_),
    .Y(_1288_)
);

NAND3X1 _7773_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1284_),
    .B(_1288_),
    .C(_1258_),
    .Y(_1289_)
);

NAND2X1 _7774_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1288_),
    .B(_1284_),
    .Y(_1290_)
);

NAND3X1 _7775_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1220_),
    .B(_1223_),
    .C(_1290_),
    .Y(_1291_)
);

NAND3X1 _7776_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1257_),
    .B(_1291_),
    .C(_1289_),
    .Y(_1292_)
);

INVX1 _7777_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1257_),
    .Y(_1293_)
);

NAND2X1 _7778_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1290_),
    .B(_1258_),
    .Y(_1294_)
);

AOI21X1 _7779_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1192_),
    .B(_1222_),
    .C(_1225_),
    .Y(_1295_)
);

AND2X2 _7780_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1284_),
    .B(_1288_),
    .Y(_1296_)
);

NAND2X1 _7781_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1295_),
    .B(_1296_),
    .Y(_1297_)
);

NAND3X1 _7782_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1293_),
    .B(_1294_),
    .C(_1297_),
    .Y(_1298_)
);

AOI21X1 _7783_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1292_),
    .B(_1298_),
    .C(_1256_),
    .Y(_1299_)
);

NAND2X1 _7784_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1292_),
    .B(_1298_),
    .Y(_1300_)
);

AOI21X1 _7785_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1228_),
    .B(_1234_),
    .C(_1300_),
    .Y(_1301_)
);

NOR2X1 _7786_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1299_),
    .B(_1301_),
    .Y(_1302_)
);

INVX1 _7787_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1302_),
    .Y(_1303_)
);

AOI21X1 _7788_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1252_),
    .B(_1255_),
    .C(_1303_),
    .Y(_1304_)
);

NAND2X1 _7789_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1174_),
    .B(_1247_),
    .Y(_1305_)
);

OAI21X1 _7790_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1305_),
    .B(_1173_),
    .C(_1255_),
    .Y(_1306_)
);

NOR2X1 _7791_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1302_),
    .B(_1306_),
    .Y(_1307_)
);

NOR2X1 _7792_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1304_),
    .B(_1307_),
    .Y(_1593_[10])
);

NAND3X1 _7793_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1292_),
    .B(_1298_),
    .C(_1256_),
    .Y(_1308_)
);

NAND2X1 _7794_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1302_),
    .B(_1306_),
    .Y(_1309_)
);

NOR2X1 _7795_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1290_),
    .B(_1295_),
    .Y(_1310_)
);

AOI21X1 _7796_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1257_),
    .B(_1291_),
    .C(_1310_),
    .Y(_1311_)
);

NAND2X1 _7797_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1265_),
    .B(_1266_),
    .Y(_1312_)
);

NAND2X1 _7798_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1281_),
    .B(_1284_),
    .Y(_1313_)
);

NOR3X1 _7799_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1102_),
    .B(_1270_),
    .C(_1213_),
    .Y(_1314_)
);

AOI22X1 _7800_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1]_5_bF$buf0 ),
    .B(gnd),
    .C(_1274_),
    .D(_1275_),
    .Y(_1315_)
);

OAI22X1 _7801_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1214_),
    .B(_1259_),
    .C(_1315_),
    .D(_1314_),
    .Y(_1316_)
);

NOR2X1 _7802_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1214_),
    .B(_1259_),
    .Y(_1317_)
);

NAND2X1 _7803_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_1271_),
    .Y(_1318_)
);

OAI21X1 _7804_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_871_),
    .B(_1102_),
    .C(_1276_),
    .Y(_1319_)
);

NAND3X1 _7805_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1317_),
    .B(_1318_),
    .C(_1319_),
    .Y(_1320_)
);

NAND2X1 _7806_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1316_),
    .B(_1320_),
    .Y(_1321_)
);

NAND2X1 _7807_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1128_),
    .B(_1202_),
    .Y(_1322_)
);

NAND2X1 _7808_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[1] [7]),
    .Y(_1323_)
);

OAI22X1 _7809_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1030_),
    .B(_1032_),
    .C(_1116_),
    .D(_941_),
    .Y(_1324_)
);

OAI21X1 _7810_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1270_),
    .B(_1323_),
    .C(_1324_),
    .Y(_1325_)
);

NAND3X1 _7811_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1322_),
    .B(_1325_),
    .C(_1279_),
    .Y(_1326_)
);

INVX1 _7812_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1326_),
    .Y(_1327_)
);

AOI21X1 _7813_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1279_),
    .B(_1322_),
    .C(_1325_),
    .Y(_1328_)
);

OAI21X1 _7814_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1328_),
    .B(_1327_),
    .C(_1321_),
    .Y(_1329_)
);

AND2X2 _7815_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1320_),
    .B(_1316_),
    .Y(_1330_)
);

INVX1 _7816_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1328_),
    .Y(_1331_)
);

NAND3X1 _7817_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1326_),
    .B(_1331_),
    .C(_1330_),
    .Y(_1332_)
);

AND2X2 _7818_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1332_),
    .B(_1329_),
    .Y(_1333_)
);

NAND2X1 _7819_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1333_),
    .B(_1313_),
    .Y(_1334_)
);

AOI21X1 _7820_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1212_),
    .B(_1204_),
    .C(_1282_),
    .Y(_1335_)
);

AOI21X1 _7821_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1267_),
    .B(_1283_),
    .C(_1335_),
    .Y(_1336_)
);

NAND2X1 _7822_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1329_),
    .B(_1332_),
    .Y(_1337_)
);

NAND2X1 _7823_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1337_),
    .B(_1336_),
    .Y(_1338_)
);

NAND3X1 _7824_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1312_),
    .B(_1338_),
    .C(_1334_),
    .Y(_1339_)
);

INVX1 _7825_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1312_),
    .Y(_1340_)
);

NAND2X1 _7826_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1337_),
    .B(_1313_),
    .Y(_1341_)
);

NAND2X1 _7827_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1336_),
    .B(_1333_),
    .Y(_1342_)
);

NAND3X1 _7828_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1340_),
    .B(_1342_),
    .C(_1341_),
    .Y(_1343_)
);

NAND2X1 _7829_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1339_),
    .B(_1343_),
    .Y(_1344_)
);

NAND2X1 _7830_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1344_),
    .B(_1311_),
    .Y(_1345_)
);

AOI21X1 _7831_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1284_),
    .B(_1288_),
    .C(_1258_),
    .Y(_1346_)
);

OAI21X1 _7832_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1293_),
    .B(_1346_),
    .C(_1289_),
    .Y(_1347_)
);

NAND3X1 _7833_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1339_),
    .B(_1343_),
    .C(_1347_),
    .Y(_1348_)
);

NAND2X1 _7834_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1345_),
    .B(_1348_),
    .Y(_1349_)
);

INVX1 _7835_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1349_),
    .Y(_1350_)
);

NAND3X1 _7836_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1308_),
    .B(_1350_),
    .C(_1309_),
    .Y(_1351_)
);

OAI21X1 _7837_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1301_),
    .B(_1304_),
    .C(_1349_),
    .Y(_1352_)
);

NAND2X1 _7838_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1351_),
    .B(_1352_),
    .Y(_1593_[11])
);

NOR3X1 _7839_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1299_),
    .B(_1301_),
    .C(_1349_),
    .Y(_1353_)
);

NAND3X1 _7840_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1251_),
    .B(_1353_),
    .C(_1094_),
    .Y(_1354_)
);

OAI21X1 _7841_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1308_),
    .B(_1349_),
    .C(_1348_),
    .Y(_1355_)
);

AOI21X1 _7842_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1353_),
    .B(_1254_),
    .C(_1355_),
    .Y(_1356_)
);

AND2X2 _7843_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1339_),
    .B(_1334_),
    .Y(_1357_)
);

OAI21X1 _7844_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1102_),
    .B(_1276_),
    .C(_1320_),
    .Y(_1358_)
);

OAI21X1 _7845_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1327_),
    .B(_1321_),
    .C(_1331_),
    .Y(_1359_)
);

INVX1 _7846_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1359_),
    .Y(_1360_)
);

INVX1 _7847_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1323_),
    .Y(_1361_)
);

NOR2X1 _7848_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_871_),
    .B(_1259_),
    .Y(_1362_)
);

NOR2X1 _7849_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1270_),
    .B(_1323_),
    .Y(_1363_)
);

NOR2X1 _7850_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_941_),
    .B(_1102_),
    .Y(_1364_)
);

NOR2X1 _7851_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1364_),
    .B(_1363_),
    .Y(_1365_)
);

AOI21X1 _7852_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_1363_),
    .C(_1365_),
    .Y(_1366_)
);

OR2X2 _7853_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1366_),
    .B(_1362_),
    .Y(_1367_)
);

NAND2X1 _7854_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1362_),
    .B(_1366_),
    .Y(_1368_)
);

NAND3X1 _7855_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1361_),
    .B(_1368_),
    .C(_1367_),
    .Y(_1369_)
);

NOR2X1 _7856_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1362_),
    .B(_1366_),
    .Y(_1370_)
);

INVX1 _7857_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1368_),
    .Y(_1371_)
);

OAI21X1 _7858_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1370_),
    .B(_1371_),
    .C(_1323_),
    .Y(_1372_)
);

NAND2X1 _7859_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1369_),
    .B(_1372_),
    .Y(_1373_)
);

NAND2X1 _7860_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1360_),
    .B(_1373_),
    .Y(_1374_)
);

NAND3X1 _7861_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1359_),
    .B(_1369_),
    .C(_1372_),
    .Y(_1375_)
);

AOI21X1 _7862_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1374_),
    .B(_1375_),
    .C(_1358_),
    .Y(_1376_)
);

NAND3X1 _7863_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1358_),
    .B(_1375_),
    .C(_1374_),
    .Y(_1377_)
);

INVX1 _7864_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1377_),
    .Y(_1378_)
);

OAI21X1 _7865_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1376_),
    .B(_1378_),
    .C(_1357_),
    .Y(_1379_)
);

OR2X2 _7866_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1378_),
    .B(_1376_),
    .Y(_1380_)
);

OR2X2 _7867_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1380_),
    .B(_1357_),
    .Y(_1381_)
);

NAND2X1 _7868_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1379_),
    .B(_1381_),
    .Y(_1382_)
);

AOI21X1 _7869_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1354_),
    .B(_1356_),
    .C(_1382_),
    .Y(_1383_)
);

NAND3X1 _7870_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1174_),
    .B(_1247_),
    .C(_1353_),
    .Y(_1384_)
);

OAI21X1 _7871_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1173_),
    .B(_1384_),
    .C(_1356_),
    .Y(_1385_)
);

INVX1 _7872_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1382_),
    .Y(_1386_)
);

NOR2X1 _7873_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1386_),
    .B(_1385_),
    .Y(_1387_)
);

NOR2X1 _7874_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1383_),
    .B(_1387_),
    .Y(_1593_[12])
);

NOR2X1 _7875_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1357_),
    .B(_1380_),
    .Y(_1388_)
);

INVX1 _7876_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1363_),
    .Y(_1389_)
);

OAI21X1 _7877_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1102_),
    .B(_1389_),
    .C(_1368_),
    .Y(_1390_)
);

INVX1 _7878_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1390_),
    .Y(_1391_)
);

NOR2X1 _7879_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1032_),
    .B(_1259_),
    .Y(_1392_)
);

NAND2X1 _7880_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1364_),
    .B(_1392_),
    .Y(_1393_)
);

OAI22X1 _7881_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_941_),
    .B(_1259_),
    .C(_1102_),
    .D(_1032_),
    .Y(_1394_)
);

NAND2X1 _7882_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1394_),
    .B(_1393_),
    .Y(_1395_)
);

NAND2X1 _7883_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1395_),
    .B(_1369_),
    .Y(_1396_)
);

OR2X2 _7884_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1369_),
    .B(_1395_),
    .Y(_1397_)
);

NAND2X1 _7885_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1396_),
    .B(_1397_),
    .Y(_1398_)
);

NAND2X1 _7886_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1391_),
    .B(_1398_),
    .Y(_1399_)
);

OR2X2 _7887_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1398_),
    .B(_1391_),
    .Y(_1400_)
);

NAND2X1 _7888_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1399_),
    .B(_1400_),
    .Y(_1401_)
);

NAND3X1 _7889_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1375_),
    .B(_1377_),
    .C(_1401_),
    .Y(_1402_)
);

OAI21X1 _7890_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1360_),
    .B(_1373_),
    .C(_1377_),
    .Y(_1403_)
);

AND2X2 _7891_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1400_),
    .B(_1399_),
    .Y(_1404_)
);

NAND2X1 _7892_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1403_),
    .B(_1404_),
    .Y(_1405_)
);

NAND2X1 _7893_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1402_),
    .B(_1405_),
    .Y(_1406_)
);

OAI21X1 _7894_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1388_),
    .B(_1383_),
    .C(_1406_),
    .Y(_1407_)
);

NAND2X1 _7895_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1386_),
    .B(_1385_),
    .Y(_1408_)
);

AND2X2 _7896_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1405_),
    .B(_1402_),
    .Y(_1409_)
);

NAND3X1 _7897_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1381_),
    .B(_1409_),
    .C(_1408_),
    .Y(_1410_)
);

NAND2X1 _7898_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1410_),
    .B(_1407_),
    .Y(_1593_[13])
);

NAND3X1 _7899_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1379_),
    .B(_1381_),
    .C(_1409_),
    .Y(_1411_)
);

AOI21X1 _7900_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1354_),
    .B(_1356_),
    .C(_1411_),
    .Y(_1412_)
);

OAI21X1 _7901_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1381_),
    .B(_1406_),
    .C(_1405_),
    .Y(_1413_)
);

OAI21X1 _7902_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1391_),
    .B(_1398_),
    .C(_1397_),
    .Y(_1414_)
);

AND2X2 _7903_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1393_),
    .B(_1392_),
    .Y(_1415_)
);

OR2X2 _7904_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1414_),
    .B(_1415_),
    .Y(_1416_)
);

NAND2X1 _7905_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1415_),
    .B(_1414_),
    .Y(_1417_)
);

NAND2X1 _7906_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1417_),
    .B(_1416_),
    .Y(_1418_)
);

OAI21X1 _7907_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1413_),
    .B(_1412_),
    .C(_1418_),
    .Y(_1419_)
);

INVX1 _7908_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1379_),
    .Y(_1420_)
);

NOR3X1 _7909_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1420_),
    .B(_1388_),
    .C(_1406_),
    .Y(_1421_)
);

NAND2X1 _7910_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1421_),
    .B(_1385_),
    .Y(_1422_)
);

INVX1 _7911_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1413_),
    .Y(_1423_)
);

INVX1 _7912_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1418_),
    .Y(_1424_)
);

NAND3X1 _7913_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1423_),
    .B(_1424_),
    .C(_1422_),
    .Y(_1425_)
);

NAND2X1 _7914_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1425_),
    .B(_1419_),
    .Y(_1593_[14])
);

OAI21X1 _7915_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1413_),
    .B(_1412_),
    .C(_1424_),
    .Y(_1426_)
);

OAI21X1 _7916_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1364_),
    .B(_1414_),
    .C(_1392_),
    .Y(_1427_)
);

NAND2X1 _7917_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1427_),
    .B(_1426_),
    .Y(_1593_[15])
);

INVX1 _7918_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_821_),
    .Y(_1588_[0])
);

AND2X2 _7919_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [0]),
    .B(\u_fir_pe1.mul [0]),
    .Y(_1428_)
);

INVX1 _7920_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [1]),
    .Y(_1429_)
);

INVX1 _7921_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.mul [1]),
    .Y(_1430_)
);

NOR2X1 _7922_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1429_),
    .B(_1430_),
    .Y(_1431_)
);

NOR2X1 _7923_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [1]),
    .B(\u_fir_pe1.mul [1]),
    .Y(_1432_)
);

NOR2X1 _7924_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1432_),
    .B(_1431_),
    .Y(_1433_)
);

NAND2X1 _7925_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1428_),
    .B(_1433_),
    .Y(_1434_)
);

INVX1 _7926_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1434_),
    .Y(_1435_)
);

NOR2X1 _7927_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1428_),
    .B(_1433_),
    .Y(_1436_)
);

NOR2X1 _7928_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1436_),
    .B(_1435_),
    .Y(_1587_[1])
);

OAI21X1 _7929_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1429_),
    .B(_1430_),
    .C(_1434_),
    .Y(_1437_)
);

AND2X2 _7930_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [2]),
    .B(\u_fir_pe1.mul [2]),
    .Y(_1438_)
);

NOR2X1 _7931_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [2]),
    .B(\u_fir_pe1.mul [2]),
    .Y(_1439_)
);

OAI21X1 _7932_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1438_),
    .B(_1439_),
    .C(_1437_),
    .Y(_1440_)
);

INVX1 _7933_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1437_),
    .Y(_1441_)
);

NOR2X1 _7934_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1439_),
    .B(_1438_),
    .Y(_1442_)
);

NAND2X1 _7935_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1442_),
    .B(_1441_),
    .Y(_1443_)
);

NAND2X1 _7936_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1440_),
    .B(_1443_),
    .Y(_1587_[2])
);

AOI21X1 _7937_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1437_),
    .B(_1442_),
    .C(_1438_),
    .Y(_1444_)
);

INVX1 _7938_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [3]),
    .Y(_1445_)
);

INVX1 _7939_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.mul [3]),
    .Y(_1446_)
);

NOR2X1 _7940_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1445_),
    .B(_1446_),
    .Y(_1447_)
);

NOR2X1 _7941_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [3]),
    .B(\u_fir_pe1.mul [3]),
    .Y(_1448_)
);

NOR2X1 _7942_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1448_),
    .B(_1447_),
    .Y(_1449_)
);

NAND2X1 _7943_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1449_),
    .B(_1444_),
    .Y(_1450_)
);

OR2X2 _7944_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1444_),
    .B(_1449_),
    .Y(_1451_)
);

NAND2X1 _7945_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1450_),
    .B(_1451_),
    .Y(_1587_[3])
);

INVX1 _7946_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [4]),
    .Y(_1452_)
);

INVX1 _7947_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.mul [4]),
    .Y(_1453_)
);

NOR2X1 _7948_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1452_),
    .B(_1453_),
    .Y(_1454_)
);

NOR2X1 _7949_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [4]),
    .B(\u_fir_pe1.mul [4]),
    .Y(_1455_)
);

NOR2X1 _7950_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1455_),
    .B(_1454_),
    .Y(_1456_)
);

INVX1 _7951_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1447_),
    .Y(_1457_)
);

OAI21X1 _7952_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1448_),
    .B(_1444_),
    .C(_1457_),
    .Y(_1458_)
);

NAND2X1 _7953_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1456_),
    .B(_1458_),
    .Y(_1459_)
);

OR2X2 _7954_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1458_),
    .B(_1456_),
    .Y(_1460_)
);

AND2X2 _7955_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1460_),
    .B(_1459_),
    .Y(_1587_[4])
);

OAI21X1 _7956_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1452_),
    .B(_1453_),
    .C(_1459_),
    .Y(_1461_)
);

INVX1 _7957_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [5]),
    .Y(_1462_)
);

INVX1 _7958_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.mul [5]),
    .Y(_1463_)
);

NOR2X1 _7959_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1462_),
    .B(_1463_),
    .Y(_1464_)
);

NOR2X1 _7960_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [5]),
    .B(\u_fir_pe1.mul [5]),
    .Y(_1465_)
);

NOR2X1 _7961_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1465_),
    .B(_1464_),
    .Y(_1466_)
);

NAND2X1 _7962_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1466_),
    .B(_1461_),
    .Y(_1467_)
);

OR2X2 _7963_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1461_),
    .B(_1466_),
    .Y(_1468_)
);

AND2X2 _7964_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1468_),
    .B(_1467_),
    .Y(_1587_[5])
);

OAI21X1 _7965_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1462_),
    .B(_1463_),
    .C(_1467_),
    .Y(_1469_)
);

INVX1 _7966_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [6]),
    .Y(_1470_)
);

INVX1 _7967_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.mul [6]),
    .Y(_1471_)
);

NOR2X1 _7968_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1470_),
    .B(_1471_),
    .Y(_1472_)
);

NOR2X1 _7969_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [6]),
    .B(\u_fir_pe1.mul [6]),
    .Y(_1473_)
);

NOR2X1 _7970_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1473_),
    .B(_1472_),
    .Y(_1474_)
);

NAND2X1 _7971_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1474_),
    .B(_1469_),
    .Y(_1475_)
);

OR2X2 _7972_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1469_),
    .B(_1474_),
    .Y(_1476_)
);

AND2X2 _7973_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1476_),
    .B(_1475_),
    .Y(_1587_[6])
);

OAI21X1 _7974_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1470_),
    .B(_1471_),
    .C(_1475_),
    .Y(_1477_)
);

INVX1 _7975_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [7]),
    .Y(_1478_)
);

INVX1 _7976_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.mul [7]),
    .Y(_1479_)
);

NOR2X1 _7977_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1478_),
    .B(_1479_),
    .Y(_1480_)
);

NOR2X1 _7978_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [7]),
    .B(\u_fir_pe1.mul [7]),
    .Y(_1481_)
);

OAI21X1 _7979_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1480_),
    .B(_1481_),
    .C(_1477_),
    .Y(_1482_)
);

INVX1 _7980_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1477_),
    .Y(_1483_)
);

NOR2X1 _7981_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1481_),
    .B(_1480_),
    .Y(_1484_)
);

NAND2X1 _7982_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1484_),
    .B(_1483_),
    .Y(_1485_)
);

NAND2X1 _7983_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1482_),
    .B(_1485_),
    .Y(_1587_[7])
);

INVX1 _7984_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [8]),
    .Y(_1487_)
);

INVX1 _7985_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.mul [8]),
    .Y(_1488_)
);

NOR2X1 _7986_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1487_),
    .B(_1488_),
    .Y(_1489_)
);

NOR2X1 _7987_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [8]),
    .B(\u_fir_pe1.mul [8]),
    .Y(_1490_)
);

NAND2X1 _7988_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1454_),
    .B(_1466_),
    .Y(_1491_)
);

OAI21X1 _7989_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1462_),
    .B(_1463_),
    .C(_1491_),
    .Y(_1492_)
);

NAND2X1 _7990_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1472_),
    .B(_1484_),
    .Y(_1493_)
);

OAI21X1 _7991_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1478_),
    .B(_1479_),
    .C(_1493_),
    .Y(_1494_)
);

AND2X2 _7992_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1474_),
    .B(_1484_),
    .Y(_1495_)
);

AOI21X1 _7993_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1492_),
    .B(_1495_),
    .C(_1494_),
    .Y(_1496_)
);

AND2X2 _7994_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1456_),
    .B(_1466_),
    .Y(_1498_)
);

NAND3X1 _7995_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1498_),
    .B(_1495_),
    .C(_1458_),
    .Y(_1499_)
);

NAND2X1 _7996_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1496_),
    .B(_1499_),
    .Y(_1500_)
);

OAI21X1 _7997_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1489_),
    .B(_1490_),
    .C(_1500_),
    .Y(_1501_)
);

NOR2X1 _7998_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1490_),
    .B(_1489_),
    .Y(_1502_)
);

INVX1 _7999_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1500_),
    .Y(_1503_)
);

NAND2X1 _8000_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1502_),
    .B(_1503_),
    .Y(_1504_)
);

NAND2X1 _8001_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1501_),
    .B(_1504_),
    .Y(_1587_[8])
);

INVX1 _8002_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1489_),
    .Y(_1505_)
);

INVX1 _8003_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1502_),
    .Y(_1506_)
);

OAI21X1 _8004_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1506_),
    .B(_1503_),
    .C(_1505_),
    .Y(_1508_)
);

AND2X2 _8005_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [9]),
    .B(\u_fir_pe1.mul [9]),
    .Y(_1509_)
);

NOR2X1 _8006_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [9]),
    .B(\u_fir_pe1.mul [9]),
    .Y(_1510_)
);

NOR2X1 _8007_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1510_),
    .B(_1509_),
    .Y(_1511_)
);

INVX1 _8008_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1511_),
    .Y(_1512_)
);

OR2X2 _8009_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1508_),
    .B(_1512_),
    .Y(_1513_)
);

OAI21X1 _8010_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1509_),
    .B(_1510_),
    .C(_1508_),
    .Y(_1514_)
);

NAND2X1 _8011_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1514_),
    .B(_1513_),
    .Y(_1587_[9])
);

NOR2X1 _8012_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1512_),
    .B(_1506_),
    .Y(_1515_)
);

AOI21X1 _8013_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1511_),
    .B(_1489_),
    .C(_1509_),
    .Y(_1516_)
);

INVX1 _8014_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1516_),
    .Y(_1518_)
);

AOI21X1 _8015_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1500_),
    .B(_1515_),
    .C(_1518_),
    .Y(_1519_)
);

INVX1 _8016_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1519_),
    .Y(_1520_)
);

INVX1 _8017_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [10]),
    .Y(_1521_)
);

INVX1 _8018_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.mul [10]),
    .Y(_1522_)
);

NOR2X1 _8019_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1521_),
    .B(_1522_),
    .Y(_1523_)
);

NOR2X1 _8020_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [10]),
    .B(\u_fir_pe1.mul [10]),
    .Y(_1524_)
);

NOR2X1 _8021_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1524_),
    .B(_1523_),
    .Y(_1525_)
);

NAND2X1 _8022_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1525_),
    .B(_1520_),
    .Y(_1526_)
);

OAI21X1 _8023_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1523_),
    .B(_1524_),
    .C(_1519_),
    .Y(_1527_)
);

AND2X2 _8024_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1526_),
    .B(_1527_),
    .Y(_1587_[10])
);

OAI21X1 _8025_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1521_),
    .B(_1522_),
    .C(_1526_),
    .Y(_1529_)
);

AND2X2 _8026_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [11]),
    .B(\u_fir_pe1.mul [11]),
    .Y(_1530_)
);

NOR2X1 _8027_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [11]),
    .B(\u_fir_pe1.mul [11]),
    .Y(_1531_)
);

NOR2X1 _8028_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1531_),
    .B(_1530_),
    .Y(_1532_)
);

NOR2X1 _8029_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1532_),
    .B(_1529_),
    .Y(_1533_)
);

AND2X2 _8030_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1529_),
    .B(_1532_),
    .Y(_1534_)
);

NOR2X1 _8031_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1533_),
    .B(_1534_),
    .Y(_1587_[11])
);

AOI21X1 _8032_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1532_),
    .B(_1523_),
    .C(_1530_),
    .Y(_1535_)
);

NAND2X1 _8033_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1532_),
    .B(_1525_),
    .Y(_1536_)
);

OAI21X1 _8034_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1536_),
    .B(_1519_),
    .C(_1535_),
    .Y(_1538_)
);

INVX1 _8035_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [12]),
    .Y(_1539_)
);

INVX1 _8036_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.mul [12]),
    .Y(_1540_)
);

NOR2X1 _8037_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1539_),
    .B(_1540_),
    .Y(_1541_)
);

NOR2X1 _8038_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [12]),
    .B(\u_fir_pe1.mul [12]),
    .Y(_1542_)
);

NOR2X1 _8039_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1542_),
    .B(_1541_),
    .Y(_1543_)
);

NAND2X1 _8040_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1543_),
    .B(_1538_),
    .Y(_1544_)
);

OR2X2 _8041_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1538_),
    .B(_1543_),
    .Y(_1545_)
);

AND2X2 _8042_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1545_),
    .B(_1544_),
    .Y(_1587_[12])
);

OAI21X1 _8043_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1539_),
    .B(_1540_),
    .C(_1544_),
    .Y(_1546_)
);

INVX1 _8044_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [13]),
    .Y(_1548_)
);

INVX1 _8045_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.mul [13]),
    .Y(_1549_)
);

NOR2X1 _8046_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1548_),
    .B(_1549_),
    .Y(_1550_)
);

NOR2X1 _8047_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [13]),
    .B(\u_fir_pe1.mul [13]),
    .Y(_1551_)
);

NOR2X1 _8048_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1551_),
    .B(_1550_),
    .Y(_1552_)
);

NAND2X1 _8049_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1552_),
    .B(_1546_),
    .Y(_1553_)
);

OR2X2 _8050_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1546_),
    .B(_1552_),
    .Y(_1554_)
);

AND2X2 _8051_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1554_),
    .B(_1553_),
    .Y(_1587_[13])
);

OAI21X1 _8052_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1548_),
    .B(_1549_),
    .C(_1553_),
    .Y(_1555_)
);

INVX1 _8053_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [14]),
    .Y(_1556_)
);

INVX1 _8054_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.mul [14]),
    .Y(_1558_)
);

NOR2X1 _8055_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1556_),
    .B(_1558_),
    .Y(_1559_)
);

NOR2X1 _8056_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [14]),
    .B(\u_fir_pe1.mul [14]),
    .Y(_1560_)
);

NOR2X1 _8057_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1560_),
    .B(_1559_),
    .Y(_1561_)
);

AND2X2 _8058_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1555_),
    .B(_1561_),
    .Y(_1562_)
);

NOR2X1 _8059_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1561_),
    .B(_1555_),
    .Y(_1563_)
);

NOR2X1 _8060_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1563_),
    .B(_1562_),
    .Y(_1587_[14])
);

INVX1 _8061_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1559_),
    .Y(_1564_)
);

NAND2X1 _8062_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1561_),
    .B(_1555_),
    .Y(_1565_)
);

NAND2X1 _8063_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [15]),
    .B(\u_fir_pe1.mul [15]),
    .Y(_1566_)
);

OR2X2 _8064_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [15]),
    .B(\u_fir_pe1.mul [15]),
    .Y(_1568_)
);

NAND2X1 _8065_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1566_),
    .B(_1568_),
    .Y(_1569_)
);

INVX1 _8066_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1569_),
    .Y(_1570_)
);

NAND3X1 _8067_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1564_),
    .B(_1570_),
    .C(_1565_),
    .Y(_1571_)
);

OAI21X1 _8068_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1559_),
    .B(_1562_),
    .C(_1569_),
    .Y(_1572_)
);

NAND2X1 _8069_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1571_),
    .B(_1572_),
    .Y(_1587_[15])
);

NOR2X1 _8070_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe1.rYin [0]),
    .B(\u_fir_pe1.mul [0]),
    .Y(_1573_)
);

NOR2X1 _8071_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1573_),
    .B(_1428_),
    .Y(_1586_[0])
);

AOI21X1 _8072_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[1] [0]),
    .B(gnd),
    .C(_1497_),
    .Y(_1574_)
);

NOR2X1 _8073_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1574_),
    .B(_1517_),
    .Y(_1589_[1])
);

NOR2X1 _8074_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1517_),
    .B(_1581_),
    .Y(_1576_)
);

NOR2X1 _8075_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1576_),
    .B(_1583_),
    .Y(_1590_[2])
);

DFFPOSX1 _8076_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf9),
    .D(_1586_[0]),
    .Q(\Y[2] [0])
);

DFFPOSX1 _8077_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf8),
    .D(_1587_[1]),
    .Q(\Y[2] [1])
);

DFFPOSX1 _8078_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf7),
    .D(_1587_[2]),
    .Q(\Y[2] [2])
);

DFFPOSX1 _8079_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_1587_[3]),
    .Q(\Y[2] [3])
);

DFFPOSX1 _8080_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_1587_[4]),
    .Q(\Y[2] [4])
);

DFFPOSX1 _8081_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_1587_[5]),
    .Q(\Y[2] [5])
);

DFFPOSX1 _8082_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_1587_[6]),
    .Q(\Y[2] [6])
);

DFFPOSX1 _8083_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_1587_[7]),
    .Q(\Y[2] [7])
);

DFFPOSX1 _8084_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_1587_[8]),
    .Q(\Y[2] [8])
);

DFFPOSX1 _8085_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_1587_[9]),
    .Q(\Y[2] [9])
);

DFFPOSX1 _8086_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf57),
    .D(_1587_[10]),
    .Q(\Y[2] [10])
);

DFFPOSX1 _8087_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf56),
    .D(_1587_[11]),
    .Q(\Y[2] [11])
);

DFFPOSX1 _8088_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf55),
    .D(_1587_[12]),
    .Q(\Y[2] [12])
);

DFFPOSX1 _8089_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf54),
    .D(_1587_[13]),
    .Q(\Y[2] [13])
);

DFFPOSX1 _8090_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf53),
    .D(_1587_[14]),
    .Q(\Y[2] [14])
);

DFFPOSX1 _8091_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf52),
    .D(_1587_[15]),
    .Q(\Y[2] [15])
);

DFFPOSX1 _8092_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf51),
    .D(\X[1] [0]),
    .Q(\X[2] [0])
);

DFFPOSX1 _8093_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf50),
    .D(\X[1] [1]),
    .Q(\X[2] [1])
);

DFFPOSX1 _8094_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf49),
    .D(\X[1] [2]),
    .Q(\X[2] [2])
);

DFFPOSX1 _8095_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf48),
    .D(\X[1] [3]),
    .Q(\X[2] [3])
);

DFFPOSX1 _8096_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf47),
    .D(\X[1] [4]),
    .Q(\X[2] [4])
);

DFFPOSX1 _8097_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf46),
    .D(\X[1]_5_bF$buf3 ),
    .Q(\X[2] [5])
);

DFFPOSX1 _8098_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf45),
    .D(\X[1] [6]),
    .Q(\X[2] [6])
);

DFFPOSX1 _8099_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf44),
    .D(\X[1] [7]),
    .Q(\X[2] [7])
);

DFFPOSX1 _8100_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf43),
    .D(\Y[1] [0]),
    .Q(\u_fir_pe1.rYin [0])
);

DFFPOSX1 _8101_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf42),
    .D(\Y[1] [1]),
    .Q(\u_fir_pe1.rYin [1])
);

DFFPOSX1 _8102_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf41),
    .D(\Y[1] [2]),
    .Q(\u_fir_pe1.rYin [2])
);

DFFPOSX1 _8103_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf40),
    .D(\Y[1] [3]),
    .Q(\u_fir_pe1.rYin [3])
);

DFFPOSX1 _8104_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf39),
    .D(\Y[1] [4]),
    .Q(\u_fir_pe1.rYin [4])
);

DFFPOSX1 _8105_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf38),
    .D(\Y[1] [5]),
    .Q(\u_fir_pe1.rYin [5])
);

DFFPOSX1 _8106_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf37),
    .D(\Y[1] [6]),
    .Q(\u_fir_pe1.rYin [6])
);

DFFPOSX1 _8107_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf36),
    .D(\Y[1] [7]),
    .Q(\u_fir_pe1.rYin [7])
);

DFFPOSX1 _8108_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf35),
    .D(\Y[1] [8]),
    .Q(\u_fir_pe1.rYin [8])
);

DFFPOSX1 _8109_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf34),
    .D(\Y[1] [9]),
    .Q(\u_fir_pe1.rYin [9])
);

DFFPOSX1 _8110_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf33),
    .D(\Y[1] [10]),
    .Q(\u_fir_pe1.rYin [10])
);

DFFPOSX1 _8111_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf32),
    .D(\Y[1] [11]),
    .Q(\u_fir_pe1.rYin [11])
);

DFFPOSX1 _8112_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf31),
    .D(\Y[1] [12]),
    .Q(\u_fir_pe1.rYin [12])
);

DFFPOSX1 _8113_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf30),
    .D(\Y[1] [13]),
    .Q(\u_fir_pe1.rYin [13])
);

DFFPOSX1 _8114_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf29),
    .D(\Y[1] [14]),
    .Q(\u_fir_pe1.rYin [14])
);

DFFPOSX1 _8115_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf28),
    .D(\Y[1] [15]),
    .Q(\u_fir_pe1.rYin [15])
);

DFFPOSX1 _8116_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf27),
    .D(_1588_[0]),
    .Q(\u_fir_pe1.mul [0])
);

DFFPOSX1 _8117_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf26),
    .D(_1589_[1]),
    .Q(\u_fir_pe1.mul [1])
);

DFFPOSX1 _8118_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf25),
    .D(_1590_[2]),
    .Q(\u_fir_pe1.mul [2])
);

DFFPOSX1 _8119_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf24),
    .D(_1591_[3]),
    .Q(\u_fir_pe1.mul [3])
);

DFFPOSX1 _8120_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf23),
    .D(_1592_[4]),
    .Q(\u_fir_pe1.mul [4])
);

DFFPOSX1 _8121_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf22),
    .D(_1593_[5]),
    .Q(\u_fir_pe1.mul [5])
);

DFFPOSX1 _8122_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf21),
    .D(_1593_[6]),
    .Q(\u_fir_pe1.mul [6])
);

DFFPOSX1 _8123_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf20),
    .D(_1593_[7]),
    .Q(\u_fir_pe1.mul [7])
);

DFFPOSX1 _8124_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf19),
    .D(_1593_[8]),
    .Q(\u_fir_pe1.mul [8])
);

DFFPOSX1 _8125_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf18),
    .D(_1593_[9]),
    .Q(\u_fir_pe1.mul [9])
);

DFFPOSX1 _8126_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf17),
    .D(_1593_[10]),
    .Q(\u_fir_pe1.mul [10])
);

DFFPOSX1 _8127_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf16),
    .D(_1593_[11]),
    .Q(\u_fir_pe1.mul [11])
);

DFFPOSX1 _8128_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf15),
    .D(_1593_[12]),
    .Q(\u_fir_pe1.mul [12])
);

DFFPOSX1 _8129_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf14),
    .D(_1593_[13]),
    .Q(\u_fir_pe1.mul [13])
);

DFFPOSX1 _8130_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf13),
    .D(_1593_[14]),
    .Q(\u_fir_pe1.mul [14])
);

DFFPOSX1 _8131_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf12),
    .D(_1593_[15]),
    .Q(\u_fir_pe1.mul [15])
);

NAND2X1 _8132_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [0]),
    .B(gnd),
    .Y(_2283_)
);

AND2X2 _8133_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [1]),
    .B(vdd),
    .Y(_2294_)
);

INVX1 _8134_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2294_),
    .Y(_2304_)
);

NOR2X1 _8135_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2283_),
    .B(_2304_),
    .Y(_2314_)
);

NAND2X1 _8136_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [1]),
    .Y(_2325_)
);

NOR2X1 _8137_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2283_),
    .B(_2325_),
    .Y(_2334_)
);

AOI22X1 _8138_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [0]),
    .B(gnd),
    .C(\X[2] [1]),
    .D(gnd),
    .Y(_2344_)
);

NOR2X1 _8139_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2344_),
    .B(_2334_),
    .Y(_2354_)
);

INVX1 _8140_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [2]),
    .Y(_2364_)
);

INVX2 _8141_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .Y(_2372_)
);

NOR2X1 _8142_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2364_),
    .B(_2372_),
    .Y(_2374_)
);

NAND2X1 _8143_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2374_),
    .B(_2354_),
    .Y(_2375_)
);

INVX1 _8144_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2375_),
    .Y(_2376_)
);

NOR2X1 _8145_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2374_),
    .B(_2354_),
    .Y(_2377_)
);

NOR2X1 _8146_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2377_),
    .B(_2376_),
    .Y(_2378_)
);

NAND2X1 _8147_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2314_),
    .B(_2378_),
    .Y(_2379_)
);

INVX1 _8148_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2379_),
    .Y(_2380_)
);

NAND2X1 _8149_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [3]),
    .Y(_2381_)
);

INVX1 _8150_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2381_),
    .Y(_2382_)
);

NAND2X1 _8151_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [2]),
    .Y(_1594_)
);

INVX1 _8152_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1594_),
    .Y(_1595_)
);

NAND2X1 _8153_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [0]),
    .Y(_1596_)
);

OR2X2 _8154_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2325_),
    .B(_1596_),
    .Y(_1597_)
);

AOI22X1 _8155_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [0]),
    .C(gnd),
    .D(\X[2] [1]),
    .Y(_1598_)
);

INVX1 _8156_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1598_),
    .Y(_1599_)
);

NAND3X1 _8157_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1595_),
    .B(_1599_),
    .C(_1597_),
    .Y(_1600_)
);

NOR2X1 _8158_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2325_),
    .B(_1596_),
    .Y(_1601_)
);

OAI21X1 _8159_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1598_),
    .B(_1601_),
    .C(_1594_),
    .Y(_1602_)
);

NAND3X1 _8160_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2334_),
    .B(_1602_),
    .C(_1600_),
    .Y(_1603_)
);

INVX1 _8161_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2334_),
    .Y(_1604_)
);

NAND3X1 _8162_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1594_),
    .B(_1599_),
    .C(_1597_),
    .Y(_1605_)
);

OAI21X1 _8163_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1598_),
    .B(_1601_),
    .C(_1595_),
    .Y(_1606_)
);

NAND3X1 _8164_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1604_),
    .B(_1606_),
    .C(_1605_),
    .Y(_1607_)
);

NAND3X1 _8165_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2382_),
    .B(_1607_),
    .C(_1603_),
    .Y(_1608_)
);

INVX2 _8166_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [3]),
    .Y(_1609_)
);

NAND2X1 _8167_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1607_),
    .B(_1603_),
    .Y(_1610_)
);

OAI21X1 _8168_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2372_),
    .B(_1609_),
    .C(_1610_),
    .Y(_1611_)
);

NAND2X1 _8169_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1608_),
    .B(_1611_),
    .Y(_1612_)
);

NAND2X1 _8170_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2375_),
    .B(_1612_),
    .Y(_1613_)
);

NAND3X1 _8171_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2376_),
    .B(_1608_),
    .C(_1611_),
    .Y(_1614_)
);

NAND3X1 _8172_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1614_),
    .B(_2380_),
    .C(_1613_),
    .Y(_1615_)
);

INVX1 _8173_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1615_),
    .Y(_1616_)
);

AOI21X1 _8174_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1613_),
    .B(_1614_),
    .C(_2380_),
    .Y(_1617_)
);

NOR2X1 _8175_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1617_),
    .B(_1616_),
    .Y(_2388_[3])
);

NAND2X1 _8176_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [0]),
    .B(vdd),
    .Y(_1618_)
);

NAND2X1 _8177_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [4]),
    .B(vdd),
    .Y(_1619_)
);

NOR2X1 _8178_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1618_),
    .B(_1619_),
    .Y(_1620_)
);

AOI22X1 _8179_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [0]),
    .B(vdd),
    .C(vdd),
    .D(\X[2] [4]),
    .Y(_1621_)
);

NOR2X1 _8180_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1621_),
    .B(_1620_),
    .Y(_1622_)
);

INVX1 _8181_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1622_),
    .Y(_1623_)
);

NAND2X1 _8182_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [0]),
    .B(gnd),
    .Y(_1624_)
);

NAND2X1 _8183_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [1]),
    .Y(_1625_)
);

OAI22X1 _8184_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1624_),
    .B(_1625_),
    .C(_1594_),
    .D(_1598_),
    .Y(_1626_)
);

NAND2X1 _8185_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [3]),
    .Y(_1627_)
);

INVX1 _8186_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1627_),
    .Y(_1628_)
);

AND2X2 _8187_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [1]),
    .Y(_1629_)
);

AND2X2 _8188_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [2]),
    .Y(_1630_)
);

NAND2X1 _8189_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1629_),
    .B(_1630_),
    .Y(_1631_)
);

AOI22X1 _8190_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [1]),
    .C(gnd),
    .D(\X[2] [2]),
    .Y(_1632_)
);

INVX1 _8191_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1632_),
    .Y(_1633_)
);

NAND3X1 _8192_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1628_),
    .B(_1633_),
    .C(_1631_),
    .Y(_1634_)
);

NAND3X1 _8193_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [2]),
    .C(_1625_),
    .Y(_1635_)
);

NAND2X1 _8194_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [2]),
    .Y(_1636_)
);

NAND3X1 _8195_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [1]),
    .C(_1636_),
    .Y(_1637_)
);

NAND3X1 _8196_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1627_),
    .B(_1635_),
    .C(_1637_),
    .Y(_1638_)
);

NAND3X1 _8197_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1626_),
    .B(_1638_),
    .C(_1634_),
    .Y(_1639_)
);

INVX1 _8198_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1626_),
    .Y(_1640_)
);

NAND2X1 _8199_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1638_),
    .B(_1634_),
    .Y(_1641_)
);

NAND2X1 _8200_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1640_),
    .B(_1641_),
    .Y(_1642_)
);

NAND3X1 _8201_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1623_),
    .B(_1639_),
    .C(_1642_),
    .Y(_1643_)
);

NAND2X1 _8202_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1626_),
    .B(_1641_),
    .Y(_1644_)
);

NAND3X1 _8203_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1634_),
    .B(_1638_),
    .C(_1640_),
    .Y(_1645_)
);

NAND3X1 _8204_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1622_),
    .B(_1645_),
    .C(_1644_),
    .Y(_1646_)
);

AOI22X1 _8205_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1603_),
    .B(_1608_),
    .C(_1643_),
    .D(_1646_),
    .Y(_1647_)
);

INVX1 _8206_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1647_),
    .Y(_1648_)
);

NAND2X1 _8207_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1603_),
    .B(_1608_),
    .Y(_1649_)
);

NAND2X1 _8208_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1643_),
    .B(_1646_),
    .Y(_1650_)
);

OR2X2 _8209_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1650_),
    .B(_1649_),
    .Y(_1651_)
);

NAND2X1 _8210_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1648_),
    .B(_1651_),
    .Y(_1652_)
);

OAI21X1 _8211_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2375_),
    .B(_1612_),
    .C(_1615_),
    .Y(_1653_)
);

OR2X2 _8212_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1653_),
    .B(_1652_),
    .Y(_1654_)
);

NAND3X1 _8213_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1622_),
    .B(_1639_),
    .C(_1642_),
    .Y(_1655_)
);

INVX1 _8214_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1639_),
    .Y(_1656_)
);

AOI21X1 _8215_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1634_),
    .B(_1638_),
    .C(_1626_),
    .Y(_1657_)
);

OAI21X1 _8216_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1657_),
    .B(_1656_),
    .C(_1623_),
    .Y(_1658_)
);

AOI21X1 _8217_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1655_),
    .B(_1658_),
    .C(_1649_),
    .Y(_1659_)
);

OAI21X1 _8218_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1647_),
    .B(_1659_),
    .C(_1653_),
    .Y(_1660_)
);

NAND2X1 _8219_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1660_),
    .B(_1654_),
    .Y(_2389_[4])
);

NOR2X1 _8220_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1615_),
    .B(_1652_),
    .Y(_1661_)
);

NOR3X1 _8221_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1647_),
    .B(_1614_),
    .C(_1659_),
    .Y(_1662_)
);

OAI21X1 _8222_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1623_),
    .B(_1657_),
    .C(_1639_),
    .Y(_1663_)
);

NAND2X1 _8223_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [0]),
    .B(gnd),
    .Y(_1664_)
);

INVX1 _8224_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1664_),
    .Y(_1665_)
);

AND2X2 _8225_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2]_5_bF$buf3 ),
    .Y(_1666_)
);

NAND2X1 _8226_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2294_),
    .B(_1666_),
    .Y(_1667_)
);

INVX2 _8227_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2]_5_bF$buf2 ),
    .Y(_1668_)
);

NAND2X1 _8228_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [1]),
    .B(vdd),
    .Y(_1669_)
);

OAI21X1 _8229_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2372_),
    .B(_1668_),
    .C(_1669_),
    .Y(_1670_)
);

NAND3X1 _8230_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1670_),
    .B(_1665_),
    .C(_1667_),
    .Y(_1671_)
);

NAND3X1 _8231_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2]_5_bF$buf1 ),
    .C(_1669_),
    .Y(_1672_)
);

NAND2X1 _8232_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2]_5_bF$buf0 ),
    .Y(_1673_)
);

NAND3X1 _8233_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [1]),
    .B(vdd),
    .C(_1673_),
    .Y(_1674_)
);

NAND3X1 _8234_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1664_),
    .B(_1672_),
    .C(_1674_),
    .Y(_1675_)
);

AND2X2 _8235_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1671_),
    .B(_1675_),
    .Y(_1676_)
);

NAND2X1 _8236_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [2]),
    .Y(_1677_)
);

OAI22X1 _8237_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2325_),
    .B(_1677_),
    .C(_1627_),
    .D(_1632_),
    .Y(_1678_)
);

NAND2X1 _8238_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [4]),
    .Y(_1679_)
);

INVX1 _8239_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1679_),
    .Y(_1680_)
);

AND2X2 _8240_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [3]),
    .Y(_1681_)
);

NAND2X1 _8241_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1630_),
    .B(_1681_),
    .Y(_1682_)
);

INVX1 _8242_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_1683_)
);

OAI21X1 _8243_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1683_),
    .B(_1609_),
    .C(_1677_),
    .Y(_1684_)
);

NAND3X1 _8244_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1680_),
    .B(_1684_),
    .C(_1682_),
    .Y(_1685_)
);

NAND3X1 _8245_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [3]),
    .C(_1677_),
    .Y(_1686_)
);

NAND2X1 _8246_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [3]),
    .Y(_1687_)
);

NAND3X1 _8247_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [2]),
    .C(_1687_),
    .Y(_1688_)
);

NAND3X1 _8248_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1679_),
    .B(_1686_),
    .C(_1688_),
    .Y(_1689_)
);

NAND3X1 _8249_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1678_),
    .B(_1689_),
    .C(_1685_),
    .Y(_1690_)
);

INVX1 _8250_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1678_),
    .Y(_1691_)
);

AOI21X1 _8251_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1686_),
    .B(_1688_),
    .C(_1679_),
    .Y(_1692_)
);

AOI22X1 _8252_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [4]),
    .C(_1682_),
    .D(_1684_),
    .Y(_1693_)
);

OAI21X1 _8253_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1692_),
    .B(_1693_),
    .C(_1691_),
    .Y(_1694_)
);

NAND3X1 _8254_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1690_),
    .B(_1676_),
    .C(_1694_),
    .Y(_1695_)
);

NAND2X1 _8255_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1675_),
    .B(_1671_),
    .Y(_1696_)
);

OAI21X1 _8256_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1692_),
    .B(_1693_),
    .C(_1678_),
    .Y(_1697_)
);

NAND3X1 _8257_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1689_),
    .B(_1685_),
    .C(_1691_),
    .Y(_1698_)
);

NAND3X1 _8258_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1696_),
    .B(_1698_),
    .C(_1697_),
    .Y(_1699_)
);

NAND3X1 _8259_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1695_),
    .B(_1699_),
    .C(_1663_),
    .Y(_1700_)
);

AOI21X1 _8260_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1622_),
    .B(_1642_),
    .C(_1656_),
    .Y(_1701_)
);

AOI21X1 _8261_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1697_),
    .B(_1698_),
    .C(_1696_),
    .Y(_1702_)
);

AOI21X1 _8262_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1694_),
    .B(_1690_),
    .C(_1676_),
    .Y(_1703_)
);

OAI21X1 _8263_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1702_),
    .B(_1703_),
    .C(_1701_),
    .Y(_1704_)
);

NAND3X1 _8264_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1620_),
    .B(_1700_),
    .C(_1704_),
    .Y(_1705_)
);

INVX1 _8265_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1620_),
    .Y(_1706_)
);

OAI21X1 _8266_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1702_),
    .B(_1703_),
    .C(_1663_),
    .Y(_1707_)
);

NAND3X1 _8267_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1695_),
    .B(_1699_),
    .C(_1701_),
    .Y(_1708_)
);

NAND3X1 _8268_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1706_),
    .B(_1707_),
    .C(_1708_),
    .Y(_1709_)
);

NAND3X1 _8269_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1647_),
    .B(_1705_),
    .C(_1709_),
    .Y(_1710_)
);

NAND3X1 _8270_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1706_),
    .B(_1700_),
    .C(_1704_),
    .Y(_1711_)
);

NAND3X1 _8271_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1620_),
    .B(_1707_),
    .C(_1708_),
    .Y(_1712_)
);

NAND3X1 _8272_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1648_),
    .B(_1711_),
    .C(_1712_),
    .Y(_1713_)
);

NAND3X1 _8273_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1710_),
    .B(_1713_),
    .C(_1662_),
    .Y(_1714_)
);

INVX1 _8274_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1614_),
    .Y(_1715_)
);

NAND3X1 _8275_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1715_),
    .B(_1648_),
    .C(_1651_),
    .Y(_1716_)
);

NAND3X1 _8276_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1648_),
    .B(_1705_),
    .C(_1709_),
    .Y(_1717_)
);

NAND3X1 _8277_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1647_),
    .B(_1711_),
    .C(_1712_),
    .Y(_1718_)
);

NAND3X1 _8278_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1717_),
    .B(_1718_),
    .C(_1716_),
    .Y(_1719_)
);

NAND3X1 _8279_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1714_),
    .B(_1719_),
    .C(_1661_),
    .Y(_1720_)
);

INVX1 _8280_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1661_),
    .Y(_1721_)
);

INVX1 _8281_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1714_),
    .Y(_1722_)
);

INVX1 _8282_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1719_),
    .Y(_1723_)
);

OAI21X1 _8283_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1722_),
    .B(_1723_),
    .C(_1721_),
    .Y(_1724_)
);

AND2X2 _8284_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1724_),
    .B(_1720_),
    .Y(_2390_[5])
);

AND2X2 _8285_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [0]),
    .B(gnd),
    .Y(_1725_)
);

NAND2X1 _8286_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2]_5_bF$buf3 ),
    .Y(_1726_)
);

OAI21X1 _8287_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2304_),
    .B(_1726_),
    .C(_1671_),
    .Y(_1727_)
);

OR2X2 _8288_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1727_),
    .B(_1725_),
    .Y(_1728_)
);

NAND2X1 _8289_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1725_),
    .B(_1727_),
    .Y(_1729_)
);

NAND2X1 _8290_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1729_),
    .B(_1728_),
    .Y(_1730_)
);

AOI21X1 _8291_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1685_),
    .B(_1689_),
    .C(_1678_),
    .Y(_1731_)
);

OAI21X1 _8292_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1696_),
    .B(_1731_),
    .C(_1690_),
    .Y(_1732_)
);

NAND2X1 _8293_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [1]),
    .B(gnd),
    .Y(_1733_)
);

INVX1 _8294_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1733_),
    .Y(_1734_)
);

AND2X2 _8295_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [2]),
    .B(vdd),
    .Y(_1735_)
);

AND2X2 _8296_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [6]),
    .Y(_1736_)
);

NAND2X1 _8297_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1735_),
    .B(_1736_),
    .Y(_1737_)
);

INVX2 _8298_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [6]),
    .Y(_1738_)
);

NAND2X1 _8299_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [2]),
    .B(vdd),
    .Y(_1739_)
);

OAI21X1 _8300_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2372_),
    .B(_1738_),
    .C(_1739_),
    .Y(_1740_)
);

NAND3X1 _8301_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1740_),
    .B(_1734_),
    .C(_1737_),
    .Y(_1741_)
);

NAND3X1 _8302_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [6]),
    .C(_1739_),
    .Y(_1742_)
);

NAND2X1 _8303_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [6]),
    .Y(_1743_)
);

NAND2X1 _8304_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1743_),
    .B(_1735_),
    .Y(_1744_)
);

NAND3X1 _8305_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1733_),
    .B(_1742_),
    .C(_1744_),
    .Y(_1745_)
);

AND2X2 _8306_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_),
    .B(_1745_),
    .Y(_1746_)
);

NAND2X1 _8307_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [3]),
    .Y(_1747_)
);

AOI22X1 _8308_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [2]),
    .C(gnd),
    .D(\X[2] [3]),
    .Y(_1748_)
);

OAI22X1 _8309_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1636_),
    .B(_1747_),
    .C(_1679_),
    .D(_1748_),
    .Y(_1749_)
);

NAND2X1 _8310_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2]_5_bF$buf2 ),
    .Y(_1750_)
);

INVX1 _8311_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1750_),
    .Y(_1751_)
);

AND2X2 _8312_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [4]),
    .Y(_1752_)
);

NAND2X1 _8313_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1681_),
    .B(_1752_),
    .Y(_1753_)
);

AOI22X1 _8314_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [3]),
    .C(gnd),
    .D(\X[2] [4]),
    .Y(_1754_)
);

INVX1 _8315_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1754_),
    .Y(_1755_)
);

NAND3X1 _8316_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1751_),
    .B(_1755_),
    .C(_1753_),
    .Y(_1756_)
);

NAND3X1 _8317_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [4]),
    .C(_1747_),
    .Y(_1757_)
);

NAND2X1 _8318_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [4]),
    .Y(_1758_)
);

NAND3X1 _8319_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [3]),
    .C(_1758_),
    .Y(_1759_)
);

NAND3X1 _8320_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1750_),
    .B(_1757_),
    .C(_1759_),
    .Y(_1760_)
);

NAND3X1 _8321_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1749_),
    .B(_1760_),
    .C(_1756_),
    .Y(_1761_)
);

INVX1 _8322_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1749_),
    .Y(_1762_)
);

AOI21X1 _8323_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1757_),
    .B(_1759_),
    .C(_1750_),
    .Y(_1763_)
);

AOI22X1 _8324_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2]_5_bF$buf1 ),
    .C(_1753_),
    .D(_1755_),
    .Y(_1764_)
);

OAI21X1 _8325_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1763_),
    .B(_1764_),
    .C(_1762_),
    .Y(_1765_)
);

NAND3X1 _8326_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1761_),
    .B(_1746_),
    .C(_1765_),
    .Y(_1766_)
);

NAND2X1 _8327_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1745_),
    .B(_1741_),
    .Y(_1767_)
);

OAI21X1 _8328_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1763_),
    .B(_1764_),
    .C(_1749_),
    .Y(_1768_)
);

NAND3X1 _8329_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1756_),
    .B(_1760_),
    .C(_1762_),
    .Y(_1769_)
);

NAND3X1 _8330_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1767_),
    .B(_1769_),
    .C(_1768_),
    .Y(_1770_)
);

NAND3X1 _8331_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1766_),
    .B(_1732_),
    .C(_1770_),
    .Y(_1771_)
);

INVX1 _8332_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1690_),
    .Y(_1772_)
);

AOI21X1 _8333_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1676_),
    .B(_1694_),
    .C(_1772_),
    .Y(_1773_)
);

AOI21X1 _8334_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1768_),
    .B(_1769_),
    .C(_1767_),
    .Y(_1774_)
);

AOI21X1 _8335_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1765_),
    .B(_1761_),
    .C(_1746_),
    .Y(_1775_)
);

OAI21X1 _8336_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1774_),
    .B(_1775_),
    .C(_1773_),
    .Y(_1776_)
);

NAND3X1 _8337_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1730_),
    .B(_1771_),
    .C(_1776_),
    .Y(_1777_)
);

AND2X2 _8338_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1728_),
    .B(_1729_),
    .Y(_1778_)
);

OAI21X1 _8339_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1774_),
    .B(_1775_),
    .C(_1732_),
    .Y(_1779_)
);

NAND3X1 _8340_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1766_),
    .B(_1770_),
    .C(_1773_),
    .Y(_1780_)
);

NAND3X1 _8341_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1778_),
    .B(_1779_),
    .C(_1780_),
    .Y(_1781_)
);

AOI22X1 _8342_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1705_),
    .B(_1700_),
    .C(_1777_),
    .D(_1781_),
    .Y(_1782_)
);

AOI21X1 _8343_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1695_),
    .B(_1699_),
    .C(_1663_),
    .Y(_1783_)
);

OAI21X1 _8344_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1706_),
    .B(_1783_),
    .C(_1700_),
    .Y(_1784_)
);

NAND3X1 _8345_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1778_),
    .B(_1771_),
    .C(_1776_),
    .Y(_1785_)
);

NAND3X1 _8346_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1730_),
    .B(_1779_),
    .C(_1780_),
    .Y(_1786_)
);

AOI21X1 _8347_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1786_),
    .B(_1785_),
    .C(_1784_),
    .Y(_1787_)
);

OAI21X1 _8348_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1787_),
    .B(_1782_),
    .C(_1710_),
    .Y(_1788_)
);

AOI21X1 _8349_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1712_),
    .B(_1711_),
    .C(_1648_),
    .Y(_1789_)
);

NAND3X1 _8350_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1784_),
    .B(_1785_),
    .C(_1786_),
    .Y(_1790_)
);

INVX1 _8351_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1700_),
    .Y(_1791_)
);

AOI21X1 _8352_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1620_),
    .B(_1704_),
    .C(_1791_),
    .Y(_1792_)
);

AOI21X1 _8353_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1780_),
    .B(_1779_),
    .C(_1730_),
    .Y(_1793_)
);

AOI21X1 _8354_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1776_),
    .B(_1771_),
    .C(_1778_),
    .Y(_1794_)
);

OAI21X1 _8355_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1793_),
    .B(_1794_),
    .C(_1792_),
    .Y(_1795_)
);

NAND3X1 _8356_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1789_),
    .B(_1790_),
    .C(_1795_),
    .Y(_1796_)
);

NAND2X1 _8357_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1796_),
    .B(_1788_),
    .Y(_1797_)
);

AOI21X1 _8358_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1714_),
    .B(_1720_),
    .C(_1797_),
    .Y(_1798_)
);

OAI21X1 _8359_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1723_),
    .B(_1721_),
    .C(_1714_),
    .Y(_1799_)
);

AOI21X1 _8360_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1788_),
    .B(_1796_),
    .C(_1799_),
    .Y(_1800_)
);

NOR2X1 _8361_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1798_),
    .B(_1800_),
    .Y(_2390_[6])
);

INVX1 _8362_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1796_),
    .Y(_1801_)
);

AOI21X1 _8363_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1766_),
    .B(_1770_),
    .C(_1732_),
    .Y(_1802_)
);

OAI21X1 _8364_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1730_),
    .B(_1802_),
    .C(_1771_),
    .Y(_1803_)
);

NAND2X1 _8365_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [0]),
    .B(gnd),
    .Y(_1804_)
);

INVX1 _8366_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1804_),
    .Y(_1805_)
);

NAND2X1 _8367_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [1]),
    .B(gnd),
    .Y(_1806_)
);

INVX1 _8368_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1806_),
    .Y(_1807_)
);

AND2X2 _8369_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1739_),
    .B(_1743_),
    .Y(_1808_)
);

OAI21X1 _8370_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1733_),
    .B(_1808_),
    .C(_1737_),
    .Y(_1809_)
);

NAND2X1 _8371_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1807_),
    .B(_1809_),
    .Y(_1810_)
);

NAND3X1 _8372_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1737_),
    .B(_1806_),
    .C(_1741_),
    .Y(_1811_)
);

NAND3X1 _8373_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1805_),
    .B(_1811_),
    .C(_1810_),
    .Y(_1812_)
);

AOI21X1 _8374_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_),
    .B(_1737_),
    .C(_1806_),
    .Y(_1813_)
);

NOR2X1 _8375_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1807_),
    .B(_1809_),
    .Y(_1814_)
);

OAI21X1 _8376_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1813_),
    .B(_1814_),
    .C(_1804_),
    .Y(_1815_)
);

NAND2X1 _8377_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1812_),
    .B(_1815_),
    .Y(_1816_)
);

AOI21X1 _8378_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1756_),
    .B(_1760_),
    .C(_1749_),
    .Y(_1817_)
);

OAI21X1 _8379_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1767_),
    .B(_1817_),
    .C(_1761_),
    .Y(_1818_)
);

NAND2X1 _8380_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [2]),
    .B(gnd),
    .Y(_1819_)
);

INVX1 _8381_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1819_),
    .Y(_1820_)
);

AND2X2 _8382_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [3]),
    .B(vdd),
    .Y(_1821_)
);

AND2X2 _8383_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [7]),
    .Y(_1822_)
);

NAND2X1 _8384_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1821_),
    .B(_1822_),
    .Y(_1823_)
);

AOI22X1 _8385_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [7]),
    .C(\X[2] [3]),
    .D(vdd),
    .Y(_1824_)
);

INVX1 _8386_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1824_),
    .Y(_1825_)
);

NAND3X1 _8387_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1820_),
    .B(_1825_),
    .C(_1823_),
    .Y(_1826_)
);

INVX1 _8388_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .Y(_1827_)
);

OAI21X1 _8389_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1609_),
    .B(_1827_),
    .C(_1822_),
    .Y(_1828_)
);

INVX1 _8390_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [7]),
    .Y(_1829_)
);

OAI21X1 _8391_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2372_),
    .B(_1829_),
    .C(_1821_),
    .Y(_1830_)
);

NAND3X1 _8392_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1819_),
    .B(_1828_),
    .C(_1830_),
    .Y(_1831_)
);

NAND2X1 _8393_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1826_),
    .B(_1831_),
    .Y(_1832_)
);

OAI21X1 _8394_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1750_),
    .B(_1754_),
    .C(_1753_),
    .Y(_1833_)
);

NAND2X1 _8395_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [6]),
    .Y(_1834_)
);

NAND2X1 _8396_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [4]),
    .Y(_1835_)
);

AND2X2 _8397_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2]_5_bF$buf0 ),
    .Y(_1836_)
);

NAND2X1 _8398_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1835_),
    .B(_1836_),
    .Y(_1837_)
);

OAI21X1 _8399_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1683_),
    .B(_1668_),
    .C(_1752_),
    .Y(_1838_)
);

AOI21X1 _8400_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1838_),
    .B(_1837_),
    .C(_1834_),
    .Y(_1839_)
);

INVX1 _8401_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1834_),
    .Y(_1840_)
);

NAND2X1 _8402_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1752_),
    .B(_1836_),
    .Y(_1841_)
);

AOI22X1 _8403_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [4]),
    .C(gnd),
    .D(\X[2]_5_bF$buf3 ),
    .Y(_1842_)
);

INVX1 _8404_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1842_),
    .Y(_1843_)
);

AOI21X1 _8405_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1841_),
    .B(_1843_),
    .C(_1840_),
    .Y(_1844_)
);

OAI21X1 _8406_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1844_),
    .B(_1839_),
    .C(_1833_),
    .Y(_1845_)
);

AOI22X1 _8407_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1681_),
    .B(_1752_),
    .C(_1755_),
    .D(_1751_),
    .Y(_1846_)
);

NAND3X1 _8408_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1840_),
    .B(_1843_),
    .C(_1841_),
    .Y(_1847_)
);

NAND2X1 _8409_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2]_5_bF$buf2 ),
    .Y(_1848_)
);

NOR2X1 _8410_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1835_),
    .B(_1848_),
    .Y(_1849_)
);

OAI21X1 _8411_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1842_),
    .B(_1849_),
    .C(_1834_),
    .Y(_1850_)
);

NAND3X1 _8412_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1847_),
    .B(_1846_),
    .C(_1850_),
    .Y(_1851_)
);

AOI21X1 _8413_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1845_),
    .B(_1851_),
    .C(_1832_),
    .Y(_1852_)
);

AND2X2 _8414_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1831_),
    .B(_1826_),
    .Y(_1853_)
);

NAND3X1 _8415_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1833_),
    .B(_1847_),
    .C(_1850_),
    .Y(_1854_)
);

OAI21X1 _8416_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1844_),
    .B(_1839_),
    .C(_1846_),
    .Y(_1855_)
);

AOI21X1 _8417_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1855_),
    .B(_1854_),
    .C(_1853_),
    .Y(_1856_)
);

OAI21X1 _8418_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1852_),
    .B(_1856_),
    .C(_1818_),
    .Y(_1857_)
);

INVX1 _8419_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1761_),
    .Y(_1858_)
);

AOI21X1 _8420_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1746_),
    .B(_1765_),
    .C(_1858_),
    .Y(_1859_)
);

NAND3X1 _8421_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1854_),
    .B(_1853_),
    .C(_1855_),
    .Y(_1860_)
);

NAND3X1 _8422_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1832_),
    .B(_1851_),
    .C(_1845_),
    .Y(_1861_)
);

NAND3X1 _8423_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1860_),
    .B(_1861_),
    .C(_1859_),
    .Y(_1862_)
);

AOI21X1 _8424_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1862_),
    .B(_1857_),
    .C(_1816_),
    .Y(_1863_)
);

AND2X2 _8425_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1815_),
    .B(_1812_),
    .Y(_1864_)
);

NAND3X1 _8426_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1818_),
    .B(_1860_),
    .C(_1861_),
    .Y(_1865_)
);

OAI21X1 _8427_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1852_),
    .B(_1856_),
    .C(_1859_),
    .Y(_1866_)
);

AOI21X1 _8428_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1866_),
    .B(_1865_),
    .C(_1864_),
    .Y(_1867_)
);

OAI21X1 _8429_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1867_),
    .B(_1863_),
    .C(_1803_),
    .Y(_1868_)
);

INVX1 _8430_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1771_),
    .Y(_1869_)
);

AOI21X1 _8431_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1778_),
    .B(_1776_),
    .C(_1869_),
    .Y(_1870_)
);

NAND3X1 _8432_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1865_),
    .B(_1864_),
    .C(_1866_),
    .Y(_1871_)
);

NAND3X1 _8433_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1816_),
    .B(_1857_),
    .C(_1862_),
    .Y(_1872_)
);

NAND3X1 _8434_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1871_),
    .B(_1872_),
    .C(_1870_),
    .Y(_1873_)
);

AOI21X1 _8435_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1873_),
    .B(_1868_),
    .C(_1729_),
    .Y(_1874_)
);

INVX1 _8436_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1729_),
    .Y(_1875_)
);

NAND3X1 _8437_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1803_),
    .B(_1871_),
    .C(_1872_),
    .Y(_1876_)
);

OAI21X1 _8438_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1863_),
    .B(_1867_),
    .C(_1870_),
    .Y(_1877_)
);

AOI21X1 _8439_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1877_),
    .B(_1876_),
    .C(_1875_),
    .Y(_1878_)
);

OAI21X1 _8440_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1878_),
    .B(_1874_),
    .C(_1790_),
    .Y(_1879_)
);

NAND3X1 _8441_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1875_),
    .B(_1876_),
    .C(_1877_),
    .Y(_1880_)
);

NAND3X1 _8442_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1729_),
    .B(_1868_),
    .C(_1873_),
    .Y(_1881_)
);

NAND3X1 _8443_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1782_),
    .B(_1880_),
    .C(_1881_),
    .Y(_1882_)
);

AND2X2 _8444_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1879_),
    .B(_1882_),
    .Y(_1883_)
);

OAI21X1 _8445_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1801_),
    .B(_1798_),
    .C(_1883_),
    .Y(_1884_)
);

NOR2X1 _8446_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1801_),
    .B(_1798_),
    .Y(_1885_)
);

AOI21X1 _8447_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1881_),
    .B(_1880_),
    .C(_1782_),
    .Y(_1886_)
);

INVX1 _8448_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1882_),
    .Y(_1887_)
);

OAI21X1 _8449_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1886_),
    .B(_1887_),
    .C(_1885_),
    .Y(_1888_)
);

AND2X2 _8450_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1888_),
    .B(_1884_),
    .Y(_2390_[7])
);

NAND3X1 _8451_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1879_),
    .B(_1882_),
    .C(_1798_),
    .Y(_1889_)
);

AOI21X1 _8452_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1801_),
    .B(_1879_),
    .C(_1887_),
    .Y(_1890_)
);

NAND2X1 _8453_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1890_),
    .B(_1889_),
    .Y(_1891_)
);

INVX1 _8454_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1876_),
    .Y(_1892_)
);

AOI21X1 _8455_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1875_),
    .B(_1877_),
    .C(_1892_),
    .Y(_1893_)
);

OAI21X1 _8456_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1804_),
    .B(_1814_),
    .C(_1810_),
    .Y(_1894_)
);

INVX1 _8457_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1894_),
    .Y(_1895_)
);

AOI21X1 _8458_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1860_),
    .B(_1861_),
    .C(_1818_),
    .Y(_1896_)
);

OAI21X1 _8459_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1816_),
    .B(_1896_),
    .C(_1865_),
    .Y(_1897_)
);

NAND2X1 _8460_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [1]),
    .B(gnd),
    .Y(_1898_)
);

INVX2 _8461_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_1899_)
);

NOR2X1 _8462_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2364_),
    .B(_1899_),
    .Y(_1900_)
);

OAI21X1 _8463_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1819_),
    .B(_1824_),
    .C(_1823_),
    .Y(_1901_)
);

NOR2X1 _8464_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1900_),
    .B(_1901_),
    .Y(_1902_)
);

AND2X2 _8465_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1901_),
    .B(_1900_),
    .Y(_1903_)
);

OAI21X1 _8466_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1902_),
    .B(_1903_),
    .C(_1898_),
    .Y(_1904_)
);

INVX1 _8467_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1898_),
    .Y(_1905_)
);

OR2X2 _8468_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1901_),
    .B(_1900_),
    .Y(_1906_)
);

NAND2X1 _8469_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1900_),
    .B(_1901_),
    .Y(_1907_)
);

NAND3X1 _8470_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1905_),
    .B(_1907_),
    .C(_1906_),
    .Y(_1908_)
);

NAND2X1 _8471_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1904_),
    .B(_1908_),
    .Y(_1909_)
);

AOI21X1 _8472_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1850_),
    .B(_1847_),
    .C(_1833_),
    .Y(_1910_)
);

OAI21X1 _8473_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1832_),
    .B(_1910_),
    .C(_1854_),
    .Y(_1911_)
);

NAND2X1 _8474_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [3]),
    .B(vdd),
    .Y(_1912_)
);

INVX1 _8475_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_1913_)
);

OAI21X1 _8476_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1609_),
    .B(_1913_),
    .C(_1619_),
    .Y(_1914_)
);

NAND2X1 _8477_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [4]),
    .B(gnd),
    .Y(_1915_)
);

OAI21X1 _8478_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1912_),
    .B(_1915_),
    .C(_1914_),
    .Y(_1916_)
);

OAI21X1 _8479_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1834_),
    .B(_1842_),
    .C(_1841_),
    .Y(_1917_)
);

NAND2X1 _8480_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [7]),
    .Y(_1918_)
);

NAND2X1 _8481_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2]_5_bF$buf1 ),
    .Y(_1919_)
);

NAND3X1 _8482_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [6]),
    .C(_1919_),
    .Y(_1920_)
);

AND2X2 _8483_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2]_5_bF$buf0 ),
    .Y(_1921_)
);

OAI21X1 _8484_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1683_),
    .B(_1738_),
    .C(_1921_),
    .Y(_1922_)
);

AOI21X1 _8485_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1922_),
    .B(_1920_),
    .C(_1918_),
    .Y(_1923_)
);

INVX1 _8486_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1918_),
    .Y(_1924_)
);

AND2X2 _8487_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [6]),
    .Y(_1925_)
);

NAND2X1 _8488_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1921_),
    .B(_1925_),
    .Y(_1926_)
);

NAND2X1 _8489_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [6]),
    .Y(_1927_)
);

NAND2X1 _8490_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1919_),
    .B(_1927_),
    .Y(_1928_)
);

AOI21X1 _8491_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1926_),
    .B(_1928_),
    .C(_1924_),
    .Y(_1929_)
);

OAI21X1 _8492_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1929_),
    .B(_1923_),
    .C(_1917_),
    .Y(_1930_)
);

AOI21X1 _8493_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1840_),
    .B(_1843_),
    .C(_1849_),
    .Y(_1931_)
);

NAND3X1 _8494_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1924_),
    .B(_1928_),
    .C(_1926_),
    .Y(_1932_)
);

NAND3X1 _8495_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1918_),
    .B(_1920_),
    .C(_1922_),
    .Y(_1933_)
);

NAND3X1 _8496_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1932_),
    .B(_1933_),
    .C(_1931_),
    .Y(_1934_)
);

AOI21X1 _8497_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1930_),
    .B(_1934_),
    .C(_1916_),
    .Y(_1935_)
);

INVX1 _8498_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1916_),
    .Y(_1936_)
);

NAND3X1 _8499_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1917_),
    .B(_1932_),
    .C(_1933_),
    .Y(_1937_)
);

OAI21X1 _8500_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1929_),
    .B(_1923_),
    .C(_1931_),
    .Y(_1938_)
);

AOI21X1 _8501_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1938_),
    .B(_1937_),
    .C(_1936_),
    .Y(_1939_)
);

OAI21X1 _8502_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1935_),
    .B(_1939_),
    .C(_1911_),
    .Y(_1940_)
);

INVX1 _8503_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1854_),
    .Y(_1941_)
);

AOI21X1 _8504_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1853_),
    .B(_1855_),
    .C(_1941_),
    .Y(_1942_)
);

NAND3X1 _8505_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1936_),
    .B(_1937_),
    .C(_1938_),
    .Y(_1943_)
);

NAND3X1 _8506_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1916_),
    .B(_1934_),
    .C(_1930_),
    .Y(_1944_)
);

NAND3X1 _8507_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1943_),
    .B(_1944_),
    .C(_1942_),
    .Y(_1945_)
);

AOI21X1 _8508_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1945_),
    .B(_1940_),
    .C(_1909_),
    .Y(_1946_)
);

AND2X2 _8509_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1908_),
    .B(_1904_),
    .Y(_1947_)
);

NAND3X1 _8510_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1943_),
    .B(_1944_),
    .C(_1911_),
    .Y(_1948_)
);

OAI21X1 _8511_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1935_),
    .B(_1939_),
    .C(_1942_),
    .Y(_1949_)
);

AOI21X1 _8512_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1949_),
    .B(_1948_),
    .C(_1947_),
    .Y(_1950_)
);

OAI21X1 _8513_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1950_),
    .B(_1946_),
    .C(_1897_),
    .Y(_1951_)
);

INVX1 _8514_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1865_),
    .Y(_1952_)
);

AOI21X1 _8515_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1864_),
    .B(_1866_),
    .C(_1952_),
    .Y(_1953_)
);

NAND3X1 _8516_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1947_),
    .B(_1948_),
    .C(_1949_),
    .Y(_1954_)
);

NAND3X1 _8517_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1909_),
    .B(_1940_),
    .C(_1945_),
    .Y(_1955_)
);

NAND3X1 _8518_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1954_),
    .B(_1955_),
    .C(_1953_),
    .Y(_1956_)
);

AOI21X1 _8519_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1951_),
    .B(_1956_),
    .C(_1895_),
    .Y(_1957_)
);

NAND3X1 _8520_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1897_),
    .B(_1954_),
    .C(_1955_),
    .Y(_1958_)
);

OAI21X1 _8521_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1950_),
    .B(_1946_),
    .C(_1953_),
    .Y(_1959_)
);

AOI21X1 _8522_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1959_),
    .B(_1958_),
    .C(_1894_),
    .Y(_1960_)
);

OAI21X1 _8523_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1960_),
    .B(_1957_),
    .C(_1893_),
    .Y(_1961_)
);

AOI21X1 _8524_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1872_),
    .B(_1871_),
    .C(_1803_),
    .Y(_1962_)
);

OAI21X1 _8525_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1729_),
    .B(_1962_),
    .C(_1876_),
    .Y(_1963_)
);

NAND3X1 _8526_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1894_),
    .B(_1958_),
    .C(_1959_),
    .Y(_1964_)
);

NAND3X1 _8527_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1895_),
    .B(_1956_),
    .C(_1951_),
    .Y(_1965_)
);

NAND3X1 _8528_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1963_),
    .B(_1964_),
    .C(_1965_),
    .Y(_1966_)
);

NAND2X1 _8529_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1966_),
    .B(_1961_),
    .Y(_1967_)
);

NAND2X1 _8530_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1967_),
    .B(_1891_),
    .Y(_1968_)
);

OAI21X1 _8531_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1796_),
    .B(_1886_),
    .C(_1882_),
    .Y(_1969_)
);

AOI21X1 _8532_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1883_),
    .B(_1798_),
    .C(_1969_),
    .Y(_1970_)
);

AND2X2 _8533_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1961_),
    .B(_1966_),
    .Y(_1971_)
);

NAND2X1 _8534_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1971_),
    .B(_1970_),
    .Y(_1972_)
);

NAND2X1 _8535_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1968_),
    .B(_1972_),
    .Y(_2390_[8])
);

INVX1 _8536_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1966_),
    .Y(_1973_)
);

AOI21X1 _8537_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1891_),
    .B(_1961_),
    .C(_1973_),
    .Y(_1974_)
);

AOI21X1 _8538_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1955_),
    .B(_1954_),
    .C(_1897_),
    .Y(_1975_)
);

OAI21X1 _8539_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1895_),
    .B(_1975_),
    .C(_1958_),
    .Y(_1976_)
);

OAI21X1 _8540_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1898_),
    .B(_1902_),
    .C(_1907_),
    .Y(_1977_)
);

AOI21X1 _8541_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1943_),
    .B(_1944_),
    .C(_1911_),
    .Y(_1978_)
);

OAI21X1 _8542_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1909_),
    .B(_1978_),
    .C(_1948_),
    .Y(_1979_)
);

NAND2X1 _8543_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [2]),
    .B(gnd),
    .Y(_1980_)
);

NOR2X1 _8544_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1912_),
    .B(_1915_),
    .Y(_1981_)
);

NAND2X1 _8545_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_1981_),
    .Y(_1982_)
);

INVX1 _8546_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1982_),
    .Y(_1983_)
);

AOI21X1 _8547_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [3]),
    .B(gnd),
    .C(_1981_),
    .Y(_1984_)
);

OAI21X1 _8548_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1984_),
    .B(_1983_),
    .C(_1980_),
    .Y(_1985_)
);

INVX1 _8549_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1980_),
    .Y(_1986_)
);

INVX1 _8550_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1984_),
    .Y(_1987_)
);

NAND3X1 _8551_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1986_),
    .B(_1982_),
    .C(_1987_),
    .Y(_1988_)
);

AND2X2 _8552_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1988_),
    .B(_1985_),
    .Y(_1989_)
);

AOI21X1 _8553_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1933_),
    .B(_1932_),
    .C(_1917_),
    .Y(_1990_)
);

OAI21X1 _8554_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1916_),
    .B(_1990_),
    .C(_1937_),
    .Y(_1991_)
);

NOR2X1 _8555_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1726_),
    .B(_1915_),
    .Y(_1992_)
);

AND2X2 _8556_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1726_),
    .B(_1915_),
    .Y(_1993_)
);

NOR2X1 _8557_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1992_),
    .B(_1993_),
    .Y(_1994_)
);

NAND2X1 _8558_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [6]),
    .Y(_1995_)
);

AOI22X1 _8559_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2]_5_bF$buf3 ),
    .C(gnd),
    .D(\X[2] [6]),
    .Y(_1996_)
);

OAI22X1 _8560_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1848_),
    .B(_1995_),
    .C(_1918_),
    .D(_1996_),
    .Y(_1997_)
);

AOI22X1 _8561_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [6]),
    .C(gnd),
    .D(\X[2] [7]),
    .Y(_1998_)
);

AND2X2 _8562_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [7]),
    .Y(_1999_)
);

AOI21X1 _8563_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1925_),
    .B(_1999_),
    .C(_1998_),
    .Y(_2000_)
);

NAND2X1 _8564_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2000_),
    .B(_1997_),
    .Y(_2001_)
);

AND2X2 _8565_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [6]),
    .Y(_2002_)
);

AOI22X1 _8566_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1836_),
    .B(_2002_),
    .C(_1928_),
    .D(_1924_),
    .Y(_2003_)
);

NAND2X1 _8567_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [7]),
    .Y(_2004_)
);

NAND2X1 _8568_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1995_),
    .B(_2004_),
    .Y(_2005_)
);

NAND2X1 _8569_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [7]),
    .Y(_2006_)
);

OAI21X1 _8570_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1927_),
    .B(_2006_),
    .C(_2005_),
    .Y(_2007_)
);

NAND2X1 _8571_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2007_),
    .B(_2003_),
    .Y(_2008_)
);

NAND3X1 _8572_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1994_),
    .B(_2001_),
    .C(_2008_),
    .Y(_2009_)
);

NAND2X1 _8573_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2]_5_bF$buf2 ),
    .B(gnd),
    .Y(_2010_)
);

INVX1 _8574_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [4]),
    .Y(_2011_)
);

OAI21X1 _8575_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2011_),
    .B(_1913_),
    .C(_1726_),
    .Y(_2012_)
);

OAI21X1 _8576_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1619_),
    .B(_2010_),
    .C(_2012_),
    .Y(_2013_)
);

NAND2X1 _8577_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1997_),
    .B(_2007_),
    .Y(_2014_)
);

NAND2X1 _8578_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2000_),
    .B(_2003_),
    .Y(_2015_)
);

NAND3X1 _8579_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2013_),
    .B(_2014_),
    .C(_2015_),
    .Y(_2016_)
);

NAND3X1 _8580_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2009_),
    .B(_2016_),
    .C(_1991_),
    .Y(_2017_)
);

NAND2X1 _8581_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2009_),
    .B(_2016_),
    .Y(_2018_)
);

NAND3X1 _8582_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1937_),
    .B(_1943_),
    .C(_2018_),
    .Y(_2019_)
);

NAND3X1 _8583_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1989_),
    .B(_2017_),
    .C(_2019_),
    .Y(_2020_)
);

NAND2X1 _8584_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1985_),
    .B(_1988_),
    .Y(_2021_)
);

AOI21X1 _8585_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1937_),
    .B(_1943_),
    .C(_2018_),
    .Y(_2022_)
);

AOI21X1 _8586_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2009_),
    .B(_2016_),
    .C(_1991_),
    .Y(_2023_)
);

OAI21X1 _8587_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2023_),
    .B(_2022_),
    .C(_2021_),
    .Y(_2024_)
);

NAND3X1 _8588_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2020_),
    .B(_2024_),
    .C(_1979_),
    .Y(_2025_)
);

INVX1 _8589_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1948_),
    .Y(_2026_)
);

AOI21X1 _8590_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1947_),
    .B(_1949_),
    .C(_2026_),
    .Y(_2027_)
);

INVX1 _8591_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2020_),
    .Y(_2028_)
);

AOI21X1 _8592_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2019_),
    .B(_2017_),
    .C(_1989_),
    .Y(_2029_)
);

OAI21X1 _8593_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2029_),
    .B(_2028_),
    .C(_2027_),
    .Y(_2030_)
);

NAND3X1 _8594_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1977_),
    .B(_2025_),
    .C(_2030_),
    .Y(_2031_)
);

INVX1 _8595_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1977_),
    .Y(_2032_)
);

INVX1 _8596_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2025_),
    .Y(_2033_)
);

AOI21X1 _8597_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2024_),
    .B(_2020_),
    .C(_1979_),
    .Y(_2034_)
);

OAI21X1 _8598_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2034_),
    .B(_2033_),
    .C(_2032_),
    .Y(_2035_)
);

NAND3X1 _8599_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1976_),
    .B(_2031_),
    .C(_2035_),
    .Y(_2036_)
);

INVX1 _8600_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1958_),
    .Y(_2037_)
);

AOI21X1 _8601_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1894_),
    .B(_1959_),
    .C(_2037_),
    .Y(_2038_)
);

OAI21X1 _8602_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2029_),
    .B(_2028_),
    .C(_1979_),
    .Y(_2039_)
);

NAND3X1 _8603_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2020_),
    .B(_2024_),
    .C(_2027_),
    .Y(_2040_)
);

AOI21X1 _8604_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2040_),
    .B(_2039_),
    .C(_2032_),
    .Y(_2041_)
);

AOI21X1 _8605_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2030_),
    .B(_2025_),
    .C(_1977_),
    .Y(_2042_)
);

OAI21X1 _8606_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2041_),
    .B(_2042_),
    .C(_2038_),
    .Y(_2043_)
);

AND2X2 _8607_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2043_),
    .B(_2036_),
    .Y(_2044_)
);

OR2X2 _8608_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1974_),
    .B(_2044_),
    .Y(_2045_)
);

NAND2X1 _8609_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2044_),
    .B(_1974_),
    .Y(_2046_)
);

NAND2X1 _8610_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2046_),
    .B(_2045_),
    .Y(_2390_[9])
);

NAND2X1 _8611_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2036_),
    .B(_2043_),
    .Y(_2047_)
);

NOR2X1 _8612_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1967_),
    .B(_2047_),
    .Y(_2048_)
);

NAND2X1 _8613_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2048_),
    .B(_1891_),
    .Y(_2049_)
);

AOI21X1 _8614_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2035_),
    .B(_2031_),
    .C(_1976_),
    .Y(_2050_)
);

AOI21X1 _8615_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1966_),
    .B(_2036_),
    .C(_2050_),
    .Y(_2051_)
);

INVX1 _8616_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2051_),
    .Y(_2052_)
);

OAI21X1 _8617_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2032_),
    .B(_2034_),
    .C(_2025_),
    .Y(_2053_)
);

OAI21X1 _8618_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1980_),
    .B(_1984_),
    .C(_1982_),
    .Y(_2054_)
);

OAI21X1 _8619_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2021_),
    .B(_2023_),
    .C(_2017_),
    .Y(_2055_)
);

INVX2 _8620_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_2056_)
);

NOR3X1 _8621_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1899_),
    .B(_1726_),
    .C(_1915_),
    .Y(_2057_)
);

OAI22X1 _8622_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2011_),
    .B(_1899_),
    .C(_1619_),
    .D(_2010_),
    .Y(_2058_)
);

INVX1 _8623_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2058_),
    .Y(_2059_)
);

OAI22X1 _8624_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1609_),
    .B(_2056_),
    .C(_2057_),
    .D(_2059_),
    .Y(_2060_)
);

NOR2X1 _8625_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1609_),
    .B(_2056_),
    .Y(_2061_)
);

NAND2X1 _8626_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_1992_),
    .Y(_2062_)
);

NAND3X1 _8627_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2061_),
    .B(_2058_),
    .C(_2062_),
    .Y(_2063_)
);

AND2X2 _8628_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2060_),
    .B(_2063_),
    .Y(_2064_)
);

NOR2X1 _8629_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2000_),
    .B(_1997_),
    .Y(_2065_)
);

OAI21X1 _8630_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2013_),
    .B(_2065_),
    .C(_2001_),
    .Y(_2066_)
);

NAND2X1 _8631_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [6]),
    .Y(_2067_)
);

NOR2X1 _8632_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2067_),
    .B(_2010_),
    .Y(_2068_)
);

AND2X2 _8633_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2067_),
    .B(_2010_),
    .Y(_2069_)
);

OAI22X1 _8634_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1925_),
    .B(_2006_),
    .C(_2068_),
    .D(_2069_),
    .Y(_2070_)
);

AND2X2 _8635_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[2] [6]),
    .Y(_2071_)
);

AND2X2 _8636_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2]_5_bF$buf1 ),
    .B(gnd),
    .Y(_2072_)
);

NAND2X1 _8637_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2071_),
    .B(_2072_),
    .Y(_2073_)
);

OAI21X1 _8638_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1668_),
    .B(_1913_),
    .C(_2067_),
    .Y(_2074_)
);

AOI21X1 _8639_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [6]),
    .C(_2006_),
    .Y(_2075_)
);

NAND3X1 _8640_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2074_),
    .B(_2075_),
    .C(_2073_),
    .Y(_2076_)
);

AND2X2 _8641_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2070_),
    .B(_2076_),
    .Y(_2077_)
);

NAND2X1 _8642_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2077_),
    .B(_2066_),
    .Y(_2078_)
);

NAND2X1 _8643_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2076_),
    .B(_2070_),
    .Y(_2079_)
);

NAND3X1 _8644_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2001_),
    .B(_2079_),
    .C(_2009_),
    .Y(_2080_)
);

NAND3X1 _8645_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2064_),
    .B(_2080_),
    .C(_2078_),
    .Y(_2081_)
);

NAND2X1 _8646_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2063_),
    .B(_2060_),
    .Y(_2082_)
);

NAND2X1 _8647_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2079_),
    .B(_2066_),
    .Y(_2083_)
);

NAND3X1 _8648_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2001_),
    .B(_2077_),
    .C(_2009_),
    .Y(_2084_)
);

NAND3X1 _8649_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2082_),
    .B(_2084_),
    .C(_2083_),
    .Y(_2085_)
);

NAND3X1 _8650_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2081_),
    .B(_2085_),
    .C(_2055_),
    .Y(_2086_)
);

NAND2X1 _8651_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2085_),
    .B(_2081_),
    .Y(_2087_)
);

NAND3X1 _8652_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2017_),
    .B(_2020_),
    .C(_2087_),
    .Y(_2088_)
);

NAND3X1 _8653_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2054_),
    .B(_2088_),
    .C(_2086_),
    .Y(_2089_)
);

INVX1 _8654_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2054_),
    .Y(_2090_)
);

NAND2X1 _8655_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2087_),
    .B(_2055_),
    .Y(_2091_)
);

AOI21X1 _8656_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1989_),
    .B(_2019_),
    .C(_2022_),
    .Y(_2092_)
);

AND2X2 _8657_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2081_),
    .B(_2085_),
    .Y(_2093_)
);

NAND2X1 _8658_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2092_),
    .B(_2093_),
    .Y(_2094_)
);

NAND3X1 _8659_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2090_),
    .B(_2091_),
    .C(_2094_),
    .Y(_2095_)
);

AOI21X1 _8660_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2089_),
    .B(_2095_),
    .C(_2053_),
    .Y(_2096_)
);

NAND2X1 _8661_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2089_),
    .B(_2095_),
    .Y(_2097_)
);

AOI21X1 _8662_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2025_),
    .B(_2031_),
    .C(_2097_),
    .Y(_2098_)
);

NOR2X1 _8663_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2096_),
    .B(_2098_),
    .Y(_2099_)
);

INVX1 _8664_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2099_),
    .Y(_2100_)
);

AOI21X1 _8665_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2049_),
    .B(_2052_),
    .C(_2100_),
    .Y(_2101_)
);

NAND2X1 _8666_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1971_),
    .B(_2044_),
    .Y(_2102_)
);

OAI21X1 _8667_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2102_),
    .B(_1970_),
    .C(_2052_),
    .Y(_2103_)
);

NOR2X1 _8668_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2099_),
    .B(_2103_),
    .Y(_2104_)
);

NOR2X1 _8669_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2101_),
    .B(_2104_),
    .Y(_2390_[10])
);

NAND3X1 _8670_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2089_),
    .B(_2095_),
    .C(_2053_),
    .Y(_2105_)
);

NAND2X1 _8671_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2099_),
    .B(_2103_),
    .Y(_2106_)
);

NOR2X1 _8672_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2087_),
    .B(_2092_),
    .Y(_2107_)
);

AOI21X1 _8673_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2054_),
    .B(_2088_),
    .C(_2107_),
    .Y(_2108_)
);

NAND2X1 _8674_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2062_),
    .B(_2063_),
    .Y(_2109_)
);

NAND2X1 _8675_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2078_),
    .B(_2081_),
    .Y(_2110_)
);

NOR3X1 _8676_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1899_),
    .B(_2067_),
    .C(_2010_),
    .Y(_2111_)
);

AOI22X1 _8677_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2]_5_bF$buf0 ),
    .B(gnd),
    .C(_2071_),
    .D(_2072_),
    .Y(_2112_)
);

OAI22X1 _8678_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2011_),
    .B(_2056_),
    .C(_2112_),
    .D(_2111_),
    .Y(_2113_)
);

NOR2X1 _8679_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2011_),
    .B(_2056_),
    .Y(_2114_)
);

NAND2X1 _8680_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_2068_),
    .Y(_2115_)
);

OAI21X1 _8681_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1668_),
    .B(_1899_),
    .C(_2073_),
    .Y(_2116_)
);

NAND3X1 _8682_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2114_),
    .B(_2115_),
    .C(_2116_),
    .Y(_2117_)
);

NAND2X1 _8683_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2113_),
    .B(_2117_),
    .Y(_2118_)
);

NAND2X1 _8684_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1925_),
    .B(_1999_),
    .Y(_2119_)
);

NAND2X1 _8685_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[2] [7]),
    .Y(_2120_)
);

OAI22X1 _8686_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1827_),
    .B(_1829_),
    .C(_1913_),
    .D(_1738_),
    .Y(_2121_)
);

OAI21X1 _8687_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2067_),
    .B(_2120_),
    .C(_2121_),
    .Y(_2122_)
);

NAND3X1 _8688_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2119_),
    .B(_2122_),
    .C(_2076_),
    .Y(_2123_)
);

INVX1 _8689_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2123_),
    .Y(_2124_)
);

AOI21X1 _8690_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2076_),
    .B(_2119_),
    .C(_2122_),
    .Y(_2125_)
);

OAI21X1 _8691_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2125_),
    .B(_2124_),
    .C(_2118_),
    .Y(_2126_)
);

AND2X2 _8692_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2117_),
    .B(_2113_),
    .Y(_2127_)
);

INVX1 _8693_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2125_),
    .Y(_2128_)
);

NAND3X1 _8694_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2123_),
    .B(_2128_),
    .C(_2127_),
    .Y(_2129_)
);

AND2X2 _8695_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2129_),
    .B(_2126_),
    .Y(_2130_)
);

NAND2X1 _8696_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2130_),
    .B(_2110_),
    .Y(_2131_)
);

AOI21X1 _8697_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2009_),
    .B(_2001_),
    .C(_2079_),
    .Y(_2132_)
);

AOI21X1 _8698_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2064_),
    .B(_2080_),
    .C(_2132_),
    .Y(_2133_)
);

NAND2X1 _8699_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2126_),
    .B(_2129_),
    .Y(_2134_)
);

NAND2X1 _8700_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2134_),
    .B(_2133_),
    .Y(_2135_)
);

NAND3X1 _8701_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2109_),
    .B(_2135_),
    .C(_2131_),
    .Y(_2136_)
);

INVX1 _8702_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2109_),
    .Y(_2137_)
);

NAND2X1 _8703_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2134_),
    .B(_2110_),
    .Y(_2138_)
);

NAND2X1 _8704_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2133_),
    .B(_2130_),
    .Y(_2139_)
);

NAND3X1 _8705_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2137_),
    .B(_2139_),
    .C(_2138_),
    .Y(_2140_)
);

NAND2X1 _8706_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2136_),
    .B(_2140_),
    .Y(_2141_)
);

NAND2X1 _8707_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2141_),
    .B(_2108_),
    .Y(_2142_)
);

AOI21X1 _8708_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2081_),
    .B(_2085_),
    .C(_2055_),
    .Y(_2143_)
);

OAI21X1 _8709_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2090_),
    .B(_2143_),
    .C(_2086_),
    .Y(_2144_)
);

NAND3X1 _8710_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2136_),
    .B(_2140_),
    .C(_2144_),
    .Y(_2145_)
);

NAND2X1 _8711_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2142_),
    .B(_2145_),
    .Y(_2146_)
);

INVX1 _8712_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2146_),
    .Y(_2147_)
);

NAND3X1 _8713_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2105_),
    .B(_2147_),
    .C(_2106_),
    .Y(_2148_)
);

OAI21X1 _8714_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2098_),
    .B(_2101_),
    .C(_2146_),
    .Y(_2149_)
);

NAND2X1 _8715_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2148_),
    .B(_2149_),
    .Y(_2390_[11])
);

NOR3X1 _8716_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2096_),
    .B(_2098_),
    .C(_2146_),
    .Y(_2150_)
);

NAND3X1 _8717_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2048_),
    .B(_2150_),
    .C(_1891_),
    .Y(_2151_)
);

OAI21X1 _8718_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2105_),
    .B(_2146_),
    .C(_2145_),
    .Y(_2152_)
);

AOI21X1 _8719_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2150_),
    .B(_2051_),
    .C(_2152_),
    .Y(_2153_)
);

AND2X2 _8720_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2136_),
    .B(_2131_),
    .Y(_2154_)
);

OAI21X1 _8721_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1899_),
    .B(_2073_),
    .C(_2117_),
    .Y(_2155_)
);

OAI21X1 _8722_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2124_),
    .B(_2118_),
    .C(_2128_),
    .Y(_2156_)
);

INVX1 _8723_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2156_),
    .Y(_2157_)
);

INVX1 _8724_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2120_),
    .Y(_2158_)
);

NOR2X1 _8725_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1668_),
    .B(_2056_),
    .Y(_2159_)
);

NOR2X1 _8726_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2067_),
    .B(_2120_),
    .Y(_2160_)
);

NOR2X1 _8727_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1738_),
    .B(_1899_),
    .Y(_2161_)
);

NOR2X1 _8728_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2161_),
    .B(_2160_),
    .Y(_2162_)
);

AOI21X1 _8729_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_2160_),
    .C(_2162_),
    .Y(_2163_)
);

OR2X2 _8730_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2163_),
    .B(_2159_),
    .Y(_2164_)
);

NAND2X1 _8731_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2159_),
    .B(_2163_),
    .Y(_2165_)
);

NAND3X1 _8732_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2158_),
    .B(_2165_),
    .C(_2164_),
    .Y(_2166_)
);

NOR2X1 _8733_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2159_),
    .B(_2163_),
    .Y(_2167_)
);

INVX1 _8734_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2165_),
    .Y(_2168_)
);

OAI21X1 _8735_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2167_),
    .B(_2168_),
    .C(_2120_),
    .Y(_2169_)
);

NAND2X1 _8736_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2166_),
    .B(_2169_),
    .Y(_2170_)
);

NAND2X1 _8737_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2157_),
    .B(_2170_),
    .Y(_2171_)
);

NAND3X1 _8738_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2156_),
    .B(_2166_),
    .C(_2169_),
    .Y(_2172_)
);

AOI21X1 _8739_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2171_),
    .B(_2172_),
    .C(_2155_),
    .Y(_2173_)
);

NAND3X1 _8740_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2155_),
    .B(_2172_),
    .C(_2171_),
    .Y(_2174_)
);

INVX1 _8741_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2174_),
    .Y(_2175_)
);

OAI21X1 _8742_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2173_),
    .B(_2175_),
    .C(_2154_),
    .Y(_2176_)
);

OR2X2 _8743_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2175_),
    .B(_2173_),
    .Y(_2177_)
);

OR2X2 _8744_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2177_),
    .B(_2154_),
    .Y(_2178_)
);

NAND2X1 _8745_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2176_),
    .B(_2178_),
    .Y(_2179_)
);

AOI21X1 _8746_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2151_),
    .B(_2153_),
    .C(_2179_),
    .Y(_2180_)
);

NAND3X1 _8747_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1971_),
    .B(_2044_),
    .C(_2150_),
    .Y(_2181_)
);

OAI21X1 _8748_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1970_),
    .B(_2181_),
    .C(_2153_),
    .Y(_2182_)
);

INVX1 _8749_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2179_),
    .Y(_2183_)
);

NOR2X1 _8750_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2183_),
    .B(_2182_),
    .Y(_2184_)
);

NOR2X1 _8751_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2180_),
    .B(_2184_),
    .Y(_2390_[12])
);

NOR2X1 _8752_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2154_),
    .B(_2177_),
    .Y(_2185_)
);

INVX1 _8753_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2160_),
    .Y(_2186_)
);

OAI21X1 _8754_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1899_),
    .B(_2186_),
    .C(_2165_),
    .Y(_2187_)
);

INVX1 _8755_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2187_),
    .Y(_2188_)
);

NOR2X1 _8756_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1829_),
    .B(_2056_),
    .Y(_2189_)
);

NAND2X1 _8757_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2161_),
    .B(_2189_),
    .Y(_2190_)
);

OAI22X1 _8758_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1738_),
    .B(_2056_),
    .C(_1899_),
    .D(_1829_),
    .Y(_2191_)
);

NAND2X1 _8759_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2191_),
    .B(_2190_),
    .Y(_2192_)
);

NAND2X1 _8760_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2192_),
    .B(_2166_),
    .Y(_2193_)
);

OR2X2 _8761_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2166_),
    .B(_2192_),
    .Y(_2194_)
);

NAND2X1 _8762_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2193_),
    .B(_2194_),
    .Y(_2195_)
);

NAND2X1 _8763_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2188_),
    .B(_2195_),
    .Y(_2196_)
);

OR2X2 _8764_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2195_),
    .B(_2188_),
    .Y(_2197_)
);

NAND2X1 _8765_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2196_),
    .B(_2197_),
    .Y(_2198_)
);

NAND3X1 _8766_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2172_),
    .B(_2174_),
    .C(_2198_),
    .Y(_2199_)
);

OAI21X1 _8767_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2157_),
    .B(_2170_),
    .C(_2174_),
    .Y(_2200_)
);

AND2X2 _8768_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2197_),
    .B(_2196_),
    .Y(_2201_)
);

NAND2X1 _8769_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2200_),
    .B(_2201_),
    .Y(_2202_)
);

NAND2X1 _8770_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2199_),
    .B(_2202_),
    .Y(_2203_)
);

OAI21X1 _8771_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2185_),
    .B(_2180_),
    .C(_2203_),
    .Y(_2204_)
);

NAND2X1 _8772_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2183_),
    .B(_2182_),
    .Y(_2205_)
);

AND2X2 _8773_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2202_),
    .B(_2199_),
    .Y(_2206_)
);

NAND3X1 _8774_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2178_),
    .B(_2206_),
    .C(_2205_),
    .Y(_2207_)
);

NAND2X1 _8775_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2207_),
    .B(_2204_),
    .Y(_2390_[13])
);

NAND3X1 _8776_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2176_),
    .B(_2178_),
    .C(_2206_),
    .Y(_2208_)
);

AOI21X1 _8777_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2151_),
    .B(_2153_),
    .C(_2208_),
    .Y(_2209_)
);

OAI21X1 _8778_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2178_),
    .B(_2203_),
    .C(_2202_),
    .Y(_2210_)
);

OAI21X1 _8779_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2188_),
    .B(_2195_),
    .C(_2194_),
    .Y(_2211_)
);

AND2X2 _8780_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2190_),
    .B(_2189_),
    .Y(_2212_)
);

OR2X2 _8781_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2211_),
    .B(_2212_),
    .Y(_2213_)
);

NAND2X1 _8782_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2212_),
    .B(_2211_),
    .Y(_2214_)
);

NAND2X1 _8783_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2214_),
    .B(_2213_),
    .Y(_2215_)
);

OAI21X1 _8784_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2210_),
    .B(_2209_),
    .C(_2215_),
    .Y(_2216_)
);

INVX1 _8785_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2176_),
    .Y(_2217_)
);

NOR3X1 _8786_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2217_),
    .B(_2185_),
    .C(_2203_),
    .Y(_2218_)
);

NAND2X1 _8787_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2218_),
    .B(_2182_),
    .Y(_2219_)
);

INVX1 _8788_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2210_),
    .Y(_2220_)
);

INVX1 _8789_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2215_),
    .Y(_2221_)
);

NAND3X1 _8790_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2220_),
    .B(_2221_),
    .C(_2219_),
    .Y(_2222_)
);

NAND2X1 _8791_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2222_),
    .B(_2216_),
    .Y(_2390_[14])
);

OAI21X1 _8792_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2210_),
    .B(_2209_),
    .C(_2221_),
    .Y(_2223_)
);

OAI21X1 _8793_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2161_),
    .B(_2211_),
    .C(_2189_),
    .Y(_2224_)
);

NAND2X1 _8794_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2224_),
    .B(_2223_),
    .Y(_2390_[15])
);

INVX1 _8795_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1618_),
    .Y(_2385_[0])
);

AND2X2 _8796_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [0]),
    .B(\u_fir_pe2.mul [0]),
    .Y(_2225_)
);

INVX1 _8797_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [1]),
    .Y(_2226_)
);

INVX1 _8798_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.mul [1]),
    .Y(_2227_)
);

NOR2X1 _8799_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2226_),
    .B(_2227_),
    .Y(_2228_)
);

NOR2X1 _8800_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [1]),
    .B(\u_fir_pe2.mul [1]),
    .Y(_2229_)
);

NOR2X1 _8801_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2229_),
    .B(_2228_),
    .Y(_2230_)
);

NAND2X1 _8802_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2225_),
    .B(_2230_),
    .Y(_2231_)
);

INVX1 _8803_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2231_),
    .Y(_2232_)
);

NOR2X1 _8804_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2225_),
    .B(_2230_),
    .Y(_2233_)
);

NOR2X1 _8805_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2233_),
    .B(_2232_),
    .Y(_2384_[1])
);

OAI21X1 _8806_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2226_),
    .B(_2227_),
    .C(_2231_),
    .Y(_2234_)
);

AND2X2 _8807_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [2]),
    .B(\u_fir_pe2.mul [2]),
    .Y(_2235_)
);

NOR2X1 _8808_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [2]),
    .B(\u_fir_pe2.mul [2]),
    .Y(_2236_)
);

OAI21X1 _8809_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2235_),
    .B(_2236_),
    .C(_2234_),
    .Y(_2237_)
);

INVX1 _8810_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2234_),
    .Y(_2238_)
);

NOR2X1 _8811_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2236_),
    .B(_2235_),
    .Y(_2239_)
);

NAND2X1 _8812_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2239_),
    .B(_2238_),
    .Y(_2240_)
);

NAND2X1 _8813_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2237_),
    .B(_2240_),
    .Y(_2384_[2])
);

AOI21X1 _8814_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2234_),
    .B(_2239_),
    .C(_2235_),
    .Y(_2241_)
);

INVX1 _8815_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [3]),
    .Y(_2242_)
);

INVX1 _8816_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.mul [3]),
    .Y(_2243_)
);

NOR2X1 _8817_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2242_),
    .B(_2243_),
    .Y(_2244_)
);

NOR2X1 _8818_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [3]),
    .B(\u_fir_pe2.mul [3]),
    .Y(_2245_)
);

NOR2X1 _8819_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2245_),
    .B(_2244_),
    .Y(_2246_)
);

NAND2X1 _8820_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2246_),
    .B(_2241_),
    .Y(_2247_)
);

OR2X2 _8821_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2241_),
    .B(_2246_),
    .Y(_2248_)
);

NAND2X1 _8822_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2247_),
    .B(_2248_),
    .Y(_2384_[3])
);

INVX1 _8823_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [4]),
    .Y(_2249_)
);

INVX1 _8824_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.mul [4]),
    .Y(_2250_)
);

NOR2X1 _8825_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2249_),
    .B(_2250_),
    .Y(_2251_)
);

NOR2X1 _8826_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [4]),
    .B(\u_fir_pe2.mul [4]),
    .Y(_2252_)
);

NOR2X1 _8827_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2252_),
    .B(_2251_),
    .Y(_2253_)
);

INVX1 _8828_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2244_),
    .Y(_2254_)
);

OAI21X1 _8829_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2245_),
    .B(_2241_),
    .C(_2254_),
    .Y(_2255_)
);

NAND2X1 _8830_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2253_),
    .B(_2255_),
    .Y(_2256_)
);

OR2X2 _8831_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2255_),
    .B(_2253_),
    .Y(_2257_)
);

AND2X2 _8832_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2257_),
    .B(_2256_),
    .Y(_2384_[4])
);

OAI21X1 _8833_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2249_),
    .B(_2250_),
    .C(_2256_),
    .Y(_2258_)
);

INVX1 _8834_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [5]),
    .Y(_2259_)
);

INVX1 _8835_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.mul [5]),
    .Y(_2260_)
);

NOR2X1 _8836_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2259_),
    .B(_2260_),
    .Y(_2261_)
);

NOR2X1 _8837_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [5]),
    .B(\u_fir_pe2.mul [5]),
    .Y(_2262_)
);

NOR2X1 _8838_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2262_),
    .B(_2261_),
    .Y(_2263_)
);

NAND2X1 _8839_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2263_),
    .B(_2258_),
    .Y(_2264_)
);

OR2X2 _8840_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2258_),
    .B(_2263_),
    .Y(_2265_)
);

AND2X2 _8841_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2265_),
    .B(_2264_),
    .Y(_2384_[5])
);

OAI21X1 _8842_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2259_),
    .B(_2260_),
    .C(_2264_),
    .Y(_2266_)
);

INVX1 _8843_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [6]),
    .Y(_2267_)
);

INVX1 _8844_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.mul [6]),
    .Y(_2268_)
);

NOR2X1 _8845_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2267_),
    .B(_2268_),
    .Y(_2269_)
);

NOR2X1 _8846_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [6]),
    .B(\u_fir_pe2.mul [6]),
    .Y(_2270_)
);

NOR2X1 _8847_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2270_),
    .B(_2269_),
    .Y(_2271_)
);

NAND2X1 _8848_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2271_),
    .B(_2266_),
    .Y(_2272_)
);

OR2X2 _8849_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2266_),
    .B(_2271_),
    .Y(_2273_)
);

AND2X2 _8850_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2273_),
    .B(_2272_),
    .Y(_2384_[6])
);

OAI21X1 _8851_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2267_),
    .B(_2268_),
    .C(_2272_),
    .Y(_2274_)
);

INVX1 _8852_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [7]),
    .Y(_2275_)
);

INVX1 _8853_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.mul [7]),
    .Y(_2276_)
);

NOR2X1 _8854_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2275_),
    .B(_2276_),
    .Y(_2277_)
);

NOR2X1 _8855_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [7]),
    .B(\u_fir_pe2.mul [7]),
    .Y(_2278_)
);

OAI21X1 _8856_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2277_),
    .B(_2278_),
    .C(_2274_),
    .Y(_2279_)
);

INVX1 _8857_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2274_),
    .Y(_2280_)
);

NOR2X1 _8858_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2278_),
    .B(_2277_),
    .Y(_2281_)
);

NAND2X1 _8859_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2281_),
    .B(_2280_),
    .Y(_2282_)
);

NAND2X1 _8860_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2279_),
    .B(_2282_),
    .Y(_2384_[7])
);

INVX1 _8861_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [8]),
    .Y(_2284_)
);

INVX1 _8862_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.mul [8]),
    .Y(_2285_)
);

NOR2X1 _8863_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2284_),
    .B(_2285_),
    .Y(_2286_)
);

NOR2X1 _8864_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [8]),
    .B(\u_fir_pe2.mul [8]),
    .Y(_2287_)
);

NAND2X1 _8865_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2251_),
    .B(_2263_),
    .Y(_2288_)
);

OAI21X1 _8866_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2259_),
    .B(_2260_),
    .C(_2288_),
    .Y(_2289_)
);

NAND2X1 _8867_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2269_),
    .B(_2281_),
    .Y(_2290_)
);

OAI21X1 _8868_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2275_),
    .B(_2276_),
    .C(_2290_),
    .Y(_2291_)
);

AND2X2 _8869_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2271_),
    .B(_2281_),
    .Y(_2292_)
);

AOI21X1 _8870_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2289_),
    .B(_2292_),
    .C(_2291_),
    .Y(_2293_)
);

AND2X2 _8871_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2253_),
    .B(_2263_),
    .Y(_2295_)
);

NAND3X1 _8872_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2295_),
    .B(_2292_),
    .C(_2255_),
    .Y(_2296_)
);

NAND2X1 _8873_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2293_),
    .B(_2296_),
    .Y(_2297_)
);

OAI21X1 _8874_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2286_),
    .B(_2287_),
    .C(_2297_),
    .Y(_2298_)
);

NOR2X1 _8875_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2287_),
    .B(_2286_),
    .Y(_2299_)
);

INVX1 _8876_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2297_),
    .Y(_2300_)
);

NAND2X1 _8877_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2299_),
    .B(_2300_),
    .Y(_2301_)
);

NAND2X1 _8878_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2298_),
    .B(_2301_),
    .Y(_2384_[8])
);

INVX1 _8879_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2286_),
    .Y(_2302_)
);

INVX1 _8880_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2299_),
    .Y(_2303_)
);

OAI21X1 _8881_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2303_),
    .B(_2300_),
    .C(_2302_),
    .Y(_2305_)
);

AND2X2 _8882_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [9]),
    .B(\u_fir_pe2.mul [9]),
    .Y(_2306_)
);

NOR2X1 _8883_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [9]),
    .B(\u_fir_pe2.mul [9]),
    .Y(_2307_)
);

NOR2X1 _8884_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2307_),
    .B(_2306_),
    .Y(_2308_)
);

INVX1 _8885_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2308_),
    .Y(_2309_)
);

OR2X2 _8886_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2305_),
    .B(_2309_),
    .Y(_2310_)
);

OAI21X1 _8887_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2306_),
    .B(_2307_),
    .C(_2305_),
    .Y(_2311_)
);

NAND2X1 _8888_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2311_),
    .B(_2310_),
    .Y(_2384_[9])
);

NOR2X1 _8889_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2309_),
    .B(_2303_),
    .Y(_2312_)
);

AOI21X1 _8890_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2308_),
    .B(_2286_),
    .C(_2306_),
    .Y(_2313_)
);

INVX1 _8891_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2313_),
    .Y(_2315_)
);

AOI21X1 _8892_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2297_),
    .B(_2312_),
    .C(_2315_),
    .Y(_2316_)
);

INVX1 _8893_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2316_),
    .Y(_2317_)
);

INVX1 _8894_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [10]),
    .Y(_2318_)
);

INVX1 _8895_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.mul [10]),
    .Y(_2319_)
);

NOR2X1 _8896_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2318_),
    .B(_2319_),
    .Y(_2320_)
);

NOR2X1 _8897_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [10]),
    .B(\u_fir_pe2.mul [10]),
    .Y(_2321_)
);

NOR2X1 _8898_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2321_),
    .B(_2320_),
    .Y(_2322_)
);

NAND2X1 _8899_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2322_),
    .B(_2317_),
    .Y(_2323_)
);

OAI21X1 _8900_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2320_),
    .B(_2321_),
    .C(_2316_),
    .Y(_2324_)
);

AND2X2 _8901_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2323_),
    .B(_2324_),
    .Y(_2384_[10])
);

OAI21X1 _8902_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2318_),
    .B(_2319_),
    .C(_2323_),
    .Y(_2326_)
);

AND2X2 _8903_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [11]),
    .B(\u_fir_pe2.mul [11]),
    .Y(_2327_)
);

NOR2X1 _8904_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [11]),
    .B(\u_fir_pe2.mul [11]),
    .Y(_2328_)
);

NOR2X1 _8905_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2328_),
    .B(_2327_),
    .Y(_2329_)
);

NOR2X1 _8906_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2329_),
    .B(_2326_),
    .Y(_2330_)
);

AND2X2 _8907_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2326_),
    .B(_2329_),
    .Y(_2331_)
);

NOR2X1 _8908_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2330_),
    .B(_2331_),
    .Y(_2384_[11])
);

AOI21X1 _8909_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2329_),
    .B(_2320_),
    .C(_2327_),
    .Y(_2332_)
);

NAND2X1 _8910_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2329_),
    .B(_2322_),
    .Y(_2333_)
);

OAI21X1 _8911_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2333_),
    .B(_2316_),
    .C(_2332_),
    .Y(_2335_)
);

INVX1 _8912_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [12]),
    .Y(_2336_)
);

INVX1 _8913_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.mul [12]),
    .Y(_2337_)
);

NOR2X1 _8914_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2336_),
    .B(_2337_),
    .Y(_2338_)
);

NOR2X1 _8915_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [12]),
    .B(\u_fir_pe2.mul [12]),
    .Y(_2339_)
);

NOR2X1 _8916_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2339_),
    .B(_2338_),
    .Y(_2340_)
);

NAND2X1 _8917_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2340_),
    .B(_2335_),
    .Y(_2341_)
);

OR2X2 _8918_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2335_),
    .B(_2340_),
    .Y(_2342_)
);

AND2X2 _8919_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2342_),
    .B(_2341_),
    .Y(_2384_[12])
);

OAI21X1 _8920_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2336_),
    .B(_2337_),
    .C(_2341_),
    .Y(_2343_)
);

INVX1 _8921_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [13]),
    .Y(_2345_)
);

INVX1 _8922_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.mul [13]),
    .Y(_2346_)
);

NOR2X1 _8923_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2345_),
    .B(_2346_),
    .Y(_2347_)
);

NOR2X1 _8924_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [13]),
    .B(\u_fir_pe2.mul [13]),
    .Y(_2348_)
);

NOR2X1 _8925_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2348_),
    .B(_2347_),
    .Y(_2349_)
);

NAND2X1 _8926_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2349_),
    .B(_2343_),
    .Y(_2350_)
);

OR2X2 _8927_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2343_),
    .B(_2349_),
    .Y(_2351_)
);

AND2X2 _8928_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2351_),
    .B(_2350_),
    .Y(_2384_[13])
);

OAI21X1 _8929_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2345_),
    .B(_2346_),
    .C(_2350_),
    .Y(_2352_)
);

INVX1 _8930_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [14]),
    .Y(_2353_)
);

INVX1 _8931_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.mul [14]),
    .Y(_2355_)
);

NOR2X1 _8932_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2353_),
    .B(_2355_),
    .Y(_2356_)
);

NOR2X1 _8933_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [14]),
    .B(\u_fir_pe2.mul [14]),
    .Y(_2357_)
);

NOR2X1 _8934_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2357_),
    .B(_2356_),
    .Y(_2358_)
);

AND2X2 _8935_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2352_),
    .B(_2358_),
    .Y(_2359_)
);

NOR2X1 _8936_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2358_),
    .B(_2352_),
    .Y(_2360_)
);

NOR2X1 _8937_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2360_),
    .B(_2359_),
    .Y(_2384_[14])
);

INVX1 _8938_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2356_),
    .Y(_2361_)
);

NAND2X1 _8939_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2358_),
    .B(_2352_),
    .Y(_2362_)
);

NAND2X1 _8940_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [15]),
    .B(\u_fir_pe2.mul [15]),
    .Y(_2363_)
);

OR2X2 _8941_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [15]),
    .B(\u_fir_pe2.mul [15]),
    .Y(_2365_)
);

NAND2X1 _8942_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2363_),
    .B(_2365_),
    .Y(_2366_)
);

INVX1 _8943_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2366_),
    .Y(_2367_)
);

NAND3X1 _8944_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2361_),
    .B(_2367_),
    .C(_2362_),
    .Y(_2368_)
);

OAI21X1 _8945_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2356_),
    .B(_2359_),
    .C(_2366_),
    .Y(_2369_)
);

NAND2X1 _8946_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2368_),
    .B(_2369_),
    .Y(_2384_[15])
);

NOR2X1 _8947_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe2.rYin [0]),
    .B(\u_fir_pe2.mul [0]),
    .Y(_2370_)
);

NOR2X1 _8948_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2370_),
    .B(_2225_),
    .Y(_2383_[0])
);

AOI21X1 _8949_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[2] [0]),
    .B(gnd),
    .C(_2294_),
    .Y(_2371_)
);

NOR2X1 _8950_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2371_),
    .B(_2314_),
    .Y(_2386_[1])
);

NOR2X1 _8951_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2314_),
    .B(_2378_),
    .Y(_2373_)
);

NOR2X1 _8952_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2373_),
    .B(_2380_),
    .Y(_2387_[2])
);

DFFPOSX1 _8953_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf11),
    .D(_2383_[0]),
    .Q(\Y[3] [0])
);

DFFPOSX1 _8954_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf10),
    .D(_2384_[1]),
    .Q(\Y[3] [1])
);

DFFPOSX1 _8955_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf9),
    .D(_2384_[2]),
    .Q(\Y[3] [2])
);

DFFPOSX1 _8956_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf8),
    .D(_2384_[3]),
    .Q(\Y[3] [3])
);

DFFPOSX1 _8957_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf7),
    .D(_2384_[4]),
    .Q(\Y[3] [4])
);

DFFPOSX1 _8958_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_2384_[5]),
    .Q(\Y[3] [5])
);

DFFPOSX1 _8959_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_2384_[6]),
    .Q(\Y[3] [6])
);

DFFPOSX1 _8960_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_2384_[7]),
    .Q(\Y[3] [7])
);

DFFPOSX1 _8961_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_2384_[8]),
    .Q(\Y[3] [8])
);

DFFPOSX1 _8962_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_2384_[9]),
    .Q(\Y[3] [9])
);

DFFPOSX1 _8963_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_2384_[10]),
    .Q(\Y[3] [10])
);

DFFPOSX1 _8964_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_2384_[11]),
    .Q(\Y[3] [11])
);

DFFPOSX1 _8965_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf57),
    .D(_2384_[12]),
    .Q(\Y[3] [12])
);

DFFPOSX1 _8966_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf56),
    .D(_2384_[13]),
    .Q(\Y[3] [13])
);

DFFPOSX1 _8967_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf55),
    .D(_2384_[14]),
    .Q(\Y[3] [14])
);

DFFPOSX1 _8968_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf54),
    .D(_2384_[15]),
    .Q(\Y[3] [15])
);

DFFPOSX1 _8969_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf53),
    .D(\X[2] [0]),
    .Q(\X[3] [0])
);

DFFPOSX1 _8970_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf52),
    .D(\X[2] [1]),
    .Q(\X[3] [1])
);

DFFPOSX1 _8971_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf51),
    .D(\X[2] [2]),
    .Q(\X[3] [2])
);

DFFPOSX1 _8972_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf50),
    .D(\X[2] [3]),
    .Q(\X[3] [3])
);

DFFPOSX1 _8973_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf49),
    .D(\X[2] [4]),
    .Q(\X[3] [4])
);

DFFPOSX1 _8974_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf48),
    .D(\X[2]_5_bF$buf3 ),
    .Q(\X[3] [5])
);

DFFPOSX1 _8975_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf47),
    .D(\X[2] [6]),
    .Q(\X[3] [6])
);

DFFPOSX1 _8976_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf46),
    .D(\X[2] [7]),
    .Q(\X[3] [7])
);

DFFPOSX1 _8977_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf45),
    .D(\Y[2] [0]),
    .Q(\u_fir_pe2.rYin [0])
);

DFFPOSX1 _8978_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf44),
    .D(\Y[2] [1]),
    .Q(\u_fir_pe2.rYin [1])
);

DFFPOSX1 _8979_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf43),
    .D(\Y[2] [2]),
    .Q(\u_fir_pe2.rYin [2])
);

DFFPOSX1 _8980_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf42),
    .D(\Y[2] [3]),
    .Q(\u_fir_pe2.rYin [3])
);

DFFPOSX1 _8981_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf41),
    .D(\Y[2] [4]),
    .Q(\u_fir_pe2.rYin [4])
);

DFFPOSX1 _8982_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf40),
    .D(\Y[2] [5]),
    .Q(\u_fir_pe2.rYin [5])
);

DFFPOSX1 _8983_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf39),
    .D(\Y[2] [6]),
    .Q(\u_fir_pe2.rYin [6])
);

DFFPOSX1 _8984_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf38),
    .D(\Y[2] [7]),
    .Q(\u_fir_pe2.rYin [7])
);

DFFPOSX1 _8985_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf37),
    .D(\Y[2] [8]),
    .Q(\u_fir_pe2.rYin [8])
);

DFFPOSX1 _8986_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf36),
    .D(\Y[2] [9]),
    .Q(\u_fir_pe2.rYin [9])
);

DFFPOSX1 _8987_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf35),
    .D(\Y[2] [10]),
    .Q(\u_fir_pe2.rYin [10])
);

DFFPOSX1 _8988_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf34),
    .D(\Y[2] [11]),
    .Q(\u_fir_pe2.rYin [11])
);

DFFPOSX1 _8989_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf33),
    .D(\Y[2] [12]),
    .Q(\u_fir_pe2.rYin [12])
);

DFFPOSX1 _8990_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf32),
    .D(\Y[2] [13]),
    .Q(\u_fir_pe2.rYin [13])
);

DFFPOSX1 _8991_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf31),
    .D(\Y[2] [14]),
    .Q(\u_fir_pe2.rYin [14])
);

DFFPOSX1 _8992_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf30),
    .D(\Y[2] [15]),
    .Q(\u_fir_pe2.rYin [15])
);

DFFPOSX1 _8993_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf29),
    .D(_2385_[0]),
    .Q(\u_fir_pe2.mul [0])
);

DFFPOSX1 _8994_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf28),
    .D(_2386_[1]),
    .Q(\u_fir_pe2.mul [1])
);

DFFPOSX1 _8995_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf27),
    .D(_2387_[2]),
    .Q(\u_fir_pe2.mul [2])
);

DFFPOSX1 _8996_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf26),
    .D(_2388_[3]),
    .Q(\u_fir_pe2.mul [3])
);

DFFPOSX1 _8997_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf25),
    .D(_2389_[4]),
    .Q(\u_fir_pe2.mul [4])
);

DFFPOSX1 _8998_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf24),
    .D(_2390_[5]),
    .Q(\u_fir_pe2.mul [5])
);

DFFPOSX1 _8999_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf23),
    .D(_2390_[6]),
    .Q(\u_fir_pe2.mul [6])
);

DFFPOSX1 _9000_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf22),
    .D(_2390_[7]),
    .Q(\u_fir_pe2.mul [7])
);

DFFPOSX1 _9001_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf21),
    .D(_2390_[8]),
    .Q(\u_fir_pe2.mul [8])
);

DFFPOSX1 _9002_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf20),
    .D(_2390_[9]),
    .Q(\u_fir_pe2.mul [9])
);

DFFPOSX1 _9003_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf19),
    .D(_2390_[10]),
    .Q(\u_fir_pe2.mul [10])
);

DFFPOSX1 _9004_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf18),
    .D(_2390_[11]),
    .Q(\u_fir_pe2.mul [11])
);

DFFPOSX1 _9005_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf17),
    .D(_2390_[12]),
    .Q(\u_fir_pe2.mul [12])
);

DFFPOSX1 _9006_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf16),
    .D(_2390_[13]),
    .Q(\u_fir_pe2.mul [13])
);

DFFPOSX1 _9007_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf15),
    .D(_2390_[14]),
    .Q(\u_fir_pe2.mul [14])
);

DFFPOSX1 _9008_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf14),
    .D(_2390_[15]),
    .Q(\u_fir_pe2.mul [15])
);

NAND2X1 _9009_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [0]),
    .B(vdd),
    .Y(_3080_)
);

AND2X2 _9010_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [1]),
    .B(gnd),
    .Y(_3091_)
);

INVX1 _9011_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3091_),
    .Y(_3101_)
);

NOR2X1 _9012_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3080_),
    .B(_3101_),
    .Y(_3111_)
);

NAND2X1 _9013_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [1]),
    .Y(_3122_)
);

NOR2X1 _9014_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3080_),
    .B(_3122_),
    .Y(_3131_)
);

AOI22X1 _9015_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [0]),
    .B(gnd),
    .C(\X[3] [1]),
    .D(vdd),
    .Y(_3141_)
);

NOR2X1 _9016_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3141_),
    .B(_3131_),
    .Y(_3151_)
);

INVX1 _9017_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [2]),
    .Y(_3161_)
);

INVX2 _9018_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_3169_)
);

NOR2X1 _9019_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3161_),
    .B(_3169_),
    .Y(_3171_)
);

NAND2X1 _9020_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3171_),
    .B(_3151_),
    .Y(_3172_)
);

INVX1 _9021_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3172_),
    .Y(_3173_)
);

NOR2X1 _9022_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3171_),
    .B(_3151_),
    .Y(_3174_)
);

NOR2X1 _9023_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3174_),
    .B(_3173_),
    .Y(_3175_)
);

NAND2X1 _9024_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3111_),
    .B(_3175_),
    .Y(_3176_)
);

INVX1 _9025_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3176_),
    .Y(_3177_)
);

NAND2X1 _9026_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [3]),
    .Y(_3178_)
);

INVX1 _9027_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3178_),
    .Y(_3179_)
);

NAND2X1 _9028_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[3] [2]),
    .Y(_2391_)
);

INVX1 _9029_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2391_),
    .Y(_2392_)
);

NAND2X1 _9030_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [0]),
    .Y(_2393_)
);

OR2X2 _9031_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3122_),
    .B(_2393_),
    .Y(_2394_)
);

AOI22X1 _9032_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [0]),
    .C(gnd),
    .D(\X[3] [1]),
    .Y(_2395_)
);

INVX1 _9033_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2395_),
    .Y(_2396_)
);

NAND3X1 _9034_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2392_),
    .B(_2396_),
    .C(_2394_),
    .Y(_2397_)
);

NOR2X1 _9035_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3122_),
    .B(_2393_),
    .Y(_2398_)
);

OAI21X1 _9036_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2395_),
    .B(_2398_),
    .C(_2391_),
    .Y(_2399_)
);

NAND3X1 _9037_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3131_),
    .B(_2399_),
    .C(_2397_),
    .Y(_2400_)
);

INVX1 _9038_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3131_),
    .Y(_2401_)
);

NAND3X1 _9039_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2391_),
    .B(_2396_),
    .C(_2394_),
    .Y(_2402_)
);

OAI21X1 _9040_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2395_),
    .B(_2398_),
    .C(_2392_),
    .Y(_2403_)
);

NAND3X1 _9041_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2401_),
    .B(_2403_),
    .C(_2402_),
    .Y(_2404_)
);

NAND3X1 _9042_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3179_),
    .B(_2404_),
    .C(_2400_),
    .Y(_2405_)
);

INVX2 _9043_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [3]),
    .Y(_2406_)
);

NAND2X1 _9044_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2404_),
    .B(_2400_),
    .Y(_2407_)
);

OAI21X1 _9045_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3169_),
    .B(_2406_),
    .C(_2407_),
    .Y(_2408_)
);

NAND2X1 _9046_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2405_),
    .B(_2408_),
    .Y(_2409_)
);

NAND2X1 _9047_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3172_),
    .B(_2409_),
    .Y(_2410_)
);

NAND3X1 _9048_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3173_),
    .B(_2405_),
    .C(_2408_),
    .Y(_2411_)
);

NAND3X1 _9049_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2411_),
    .B(_3177_),
    .C(_2410_),
    .Y(_2412_)
);

INVX1 _9050_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2412_),
    .Y(_2413_)
);

AOI21X1 _9051_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2410_),
    .B(_2411_),
    .C(_3177_),
    .Y(_2414_)
);

NOR2X1 _9052_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2414_),
    .B(_2413_),
    .Y(_3185_[3])
);

NAND2X1 _9053_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [0]),
    .B(gnd),
    .Y(_2415_)
);

NAND2X1 _9054_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [4]),
    .B(gnd),
    .Y(_2416_)
);

NOR2X1 _9055_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2415_),
    .B(_2416_),
    .Y(_2417_)
);

AOI22X1 _9056_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [0]),
    .B(gnd),
    .C(gnd),
    .D(\X[3] [4]),
    .Y(_2418_)
);

NOR2X1 _9057_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2418_),
    .B(_2417_),
    .Y(_2419_)
);

INVX1 _9058_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2419_),
    .Y(_2420_)
);

NAND2X1 _9059_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [0]),
    .B(gnd),
    .Y(_2421_)
);

NAND2X1 _9060_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [1]),
    .Y(_2422_)
);

OAI22X1 _9061_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2421_),
    .B(_2422_),
    .C(_2391_),
    .D(_2395_),
    .Y(_2423_)
);

NAND2X1 _9062_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[3] [3]),
    .Y(_2424_)
);

INVX1 _9063_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2424_),
    .Y(_2425_)
);

AND2X2 _9064_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [1]),
    .Y(_2426_)
);

AND2X2 _9065_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [2]),
    .Y(_2427_)
);

NAND2X1 _9066_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2426_),
    .B(_2427_),
    .Y(_2428_)
);

AOI22X1 _9067_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [1]),
    .C(gnd),
    .D(\X[3] [2]),
    .Y(_2429_)
);

INVX1 _9068_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2429_),
    .Y(_2430_)
);

NAND3X1 _9069_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2425_),
    .B(_2430_),
    .C(_2428_),
    .Y(_2431_)
);

NAND3X1 _9070_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [2]),
    .C(_2422_),
    .Y(_2432_)
);

NAND2X1 _9071_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [2]),
    .Y(_2433_)
);

NAND3X1 _9072_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [1]),
    .C(_2433_),
    .Y(_2434_)
);

NAND3X1 _9073_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2424_),
    .B(_2432_),
    .C(_2434_),
    .Y(_2435_)
);

NAND3X1 _9074_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2423_),
    .B(_2435_),
    .C(_2431_),
    .Y(_2436_)
);

INVX1 _9075_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2423_),
    .Y(_2437_)
);

NAND2X1 _9076_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2435_),
    .B(_2431_),
    .Y(_2438_)
);

NAND2X1 _9077_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2437_),
    .B(_2438_),
    .Y(_2439_)
);

NAND3X1 _9078_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2420_),
    .B(_2436_),
    .C(_2439_),
    .Y(_2440_)
);

NAND2X1 _9079_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2423_),
    .B(_2438_),
    .Y(_2441_)
);

NAND3X1 _9080_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2431_),
    .B(_2435_),
    .C(_2437_),
    .Y(_2442_)
);

NAND3X1 _9081_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2419_),
    .B(_2442_),
    .C(_2441_),
    .Y(_2443_)
);

AOI22X1 _9082_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2400_),
    .B(_2405_),
    .C(_2440_),
    .D(_2443_),
    .Y(_2444_)
);

INVX1 _9083_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2444_),
    .Y(_2445_)
);

NAND2X1 _9084_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2400_),
    .B(_2405_),
    .Y(_2446_)
);

NAND2X1 _9085_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2440_),
    .B(_2443_),
    .Y(_2447_)
);

OR2X2 _9086_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2447_),
    .B(_2446_),
    .Y(_2448_)
);

NAND2X1 _9087_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2445_),
    .B(_2448_),
    .Y(_2449_)
);

OAI21X1 _9088_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3172_),
    .B(_2409_),
    .C(_2412_),
    .Y(_2450_)
);

OR2X2 _9089_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2450_),
    .B(_2449_),
    .Y(_2451_)
);

NAND3X1 _9090_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2419_),
    .B(_2436_),
    .C(_2439_),
    .Y(_2452_)
);

INVX1 _9091_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2436_),
    .Y(_2453_)
);

AOI21X1 _9092_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2431_),
    .B(_2435_),
    .C(_2423_),
    .Y(_2454_)
);

OAI21X1 _9093_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2454_),
    .B(_2453_),
    .C(_2420_),
    .Y(_2455_)
);

AOI21X1 _9094_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2452_),
    .B(_2455_),
    .C(_2446_),
    .Y(_2456_)
);

OAI21X1 _9095_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2444_),
    .B(_2456_),
    .C(_2450_),
    .Y(_2457_)
);

NAND2X1 _9096_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2457_),
    .B(_2451_),
    .Y(_3186_[4])
);

NOR2X1 _9097_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2412_),
    .B(_2449_),
    .Y(_2458_)
);

NOR3X1 _9098_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2444_),
    .B(_2411_),
    .C(_2456_),
    .Y(_2459_)
);

OAI21X1 _9099_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2420_),
    .B(_2454_),
    .C(_2436_),
    .Y(_2460_)
);

NAND2X1 _9100_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [0]),
    .B(vdd),
    .Y(_2461_)
);

INVX1 _9101_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2461_),
    .Y(_2462_)
);

AND2X2 _9102_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3]_5_bF$buf3 ),
    .Y(_2463_)
);

NAND2X1 _9103_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3091_),
    .B(_2463_),
    .Y(_2464_)
);

INVX2 _9104_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3]_5_bF$buf2 ),
    .Y(_2465_)
);

NAND2X1 _9105_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [1]),
    .B(gnd),
    .Y(_2466_)
);

OAI21X1 _9106_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3169_),
    .B(_2465_),
    .C(_2466_),
    .Y(_2467_)
);

NAND3X1 _9107_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2467_),
    .B(_2462_),
    .C(_2464_),
    .Y(_2468_)
);

NAND3X1 _9108_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3]_5_bF$buf1 ),
    .C(_2466_),
    .Y(_2469_)
);

NAND2X1 _9109_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3]_5_bF$buf0 ),
    .Y(_2470_)
);

NAND3X1 _9110_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [1]),
    .B(gnd),
    .C(_2470_),
    .Y(_2471_)
);

NAND3X1 _9111_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2461_),
    .B(_2469_),
    .C(_2471_),
    .Y(_2472_)
);

AND2X2 _9112_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2468_),
    .B(_2472_),
    .Y(_2473_)
);

NAND2X1 _9113_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [2]),
    .Y(_2474_)
);

OAI22X1 _9114_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3122_),
    .B(_2474_),
    .C(_2424_),
    .D(_2429_),
    .Y(_2475_)
);

NAND2X1 _9115_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[3] [4]),
    .Y(_2476_)
);

INVX1 _9116_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2476_),
    .Y(_2477_)
);

AND2X2 _9117_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [3]),
    .Y(_2478_)
);

NAND2X1 _9118_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2427_),
    .B(_2478_),
    .Y(_2479_)
);

INVX1 _9119_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_2480_)
);

OAI21X1 _9120_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2480_),
    .B(_2406_),
    .C(_2474_),
    .Y(_2481_)
);

NAND3X1 _9121_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2477_),
    .B(_2481_),
    .C(_2479_),
    .Y(_2482_)
);

NAND3X1 _9122_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [3]),
    .C(_2474_),
    .Y(_2483_)
);

NAND2X1 _9123_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [3]),
    .Y(_2484_)
);

NAND3X1 _9124_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [2]),
    .C(_2484_),
    .Y(_2485_)
);

NAND3X1 _9125_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2476_),
    .B(_2483_),
    .C(_2485_),
    .Y(_2486_)
);

NAND3X1 _9126_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2475_),
    .B(_2486_),
    .C(_2482_),
    .Y(_2487_)
);

INVX1 _9127_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2475_),
    .Y(_2488_)
);

AOI21X1 _9128_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2483_),
    .B(_2485_),
    .C(_2476_),
    .Y(_2489_)
);

AOI22X1 _9129_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[3] [4]),
    .C(_2479_),
    .D(_2481_),
    .Y(_2490_)
);

OAI21X1 _9130_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2489_),
    .B(_2490_),
    .C(_2488_),
    .Y(_2491_)
);

NAND3X1 _9131_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2487_),
    .B(_2473_),
    .C(_2491_),
    .Y(_2492_)
);

NAND2X1 _9132_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2472_),
    .B(_2468_),
    .Y(_2493_)
);

OAI21X1 _9133_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2489_),
    .B(_2490_),
    .C(_2475_),
    .Y(_2494_)
);

NAND3X1 _9134_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2486_),
    .B(_2482_),
    .C(_2488_),
    .Y(_2495_)
);

NAND3X1 _9135_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2493_),
    .B(_2495_),
    .C(_2494_),
    .Y(_2496_)
);

NAND3X1 _9136_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2492_),
    .B(_2496_),
    .C(_2460_),
    .Y(_2497_)
);

AOI21X1 _9137_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2419_),
    .B(_2439_),
    .C(_2453_),
    .Y(_2498_)
);

AOI21X1 _9138_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2494_),
    .B(_2495_),
    .C(_2493_),
    .Y(_2499_)
);

AOI21X1 _9139_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2491_),
    .B(_2487_),
    .C(_2473_),
    .Y(_2500_)
);

OAI21X1 _9140_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2499_),
    .B(_2500_),
    .C(_2498_),
    .Y(_2501_)
);

NAND3X1 _9141_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2417_),
    .B(_2497_),
    .C(_2501_),
    .Y(_2502_)
);

INVX1 _9142_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2417_),
    .Y(_2503_)
);

OAI21X1 _9143_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2499_),
    .B(_2500_),
    .C(_2460_),
    .Y(_2504_)
);

NAND3X1 _9144_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2492_),
    .B(_2496_),
    .C(_2498_),
    .Y(_2505_)
);

NAND3X1 _9145_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2503_),
    .B(_2504_),
    .C(_2505_),
    .Y(_2506_)
);

NAND3X1 _9146_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2444_),
    .B(_2502_),
    .C(_2506_),
    .Y(_2507_)
);

NAND3X1 _9147_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2503_),
    .B(_2497_),
    .C(_2501_),
    .Y(_2508_)
);

NAND3X1 _9148_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2417_),
    .B(_2504_),
    .C(_2505_),
    .Y(_2509_)
);

NAND3X1 _9149_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2445_),
    .B(_2508_),
    .C(_2509_),
    .Y(_2510_)
);

NAND3X1 _9150_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2507_),
    .B(_2510_),
    .C(_2459_),
    .Y(_2511_)
);

INVX1 _9151_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2411_),
    .Y(_2512_)
);

NAND3X1 _9152_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2512_),
    .B(_2445_),
    .C(_2448_),
    .Y(_2513_)
);

NAND3X1 _9153_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2445_),
    .B(_2502_),
    .C(_2506_),
    .Y(_2514_)
);

NAND3X1 _9154_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2444_),
    .B(_2508_),
    .C(_2509_),
    .Y(_2515_)
);

NAND3X1 _9155_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2514_),
    .B(_2515_),
    .C(_2513_),
    .Y(_2516_)
);

NAND3X1 _9156_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2511_),
    .B(_2516_),
    .C(_2458_),
    .Y(_2517_)
);

INVX1 _9157_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2458_),
    .Y(_2518_)
);

INVX1 _9158_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2511_),
    .Y(_2519_)
);

INVX1 _9159_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2516_),
    .Y(_2520_)
);

OAI21X1 _9160_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2519_),
    .B(_2520_),
    .C(_2518_),
    .Y(_2521_)
);

AND2X2 _9161_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2521_),
    .B(_2517_),
    .Y(_3187_[5])
);

AND2X2 _9162_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [0]),
    .B(gnd),
    .Y(_2522_)
);

NAND2X1 _9163_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3]_5_bF$buf3 ),
    .Y(_2523_)
);

OAI21X1 _9164_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3101_),
    .B(_2523_),
    .C(_2468_),
    .Y(_2524_)
);

OR2X2 _9165_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2524_),
    .B(_2522_),
    .Y(_2525_)
);

NAND2X1 _9166_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2522_),
    .B(_2524_),
    .Y(_2526_)
);

NAND2X1 _9167_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2526_),
    .B(_2525_),
    .Y(_2527_)
);

AOI21X1 _9168_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2482_),
    .B(_2486_),
    .C(_2475_),
    .Y(_2528_)
);

OAI21X1 _9169_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2493_),
    .B(_2528_),
    .C(_2487_),
    .Y(_2529_)
);

NAND2X1 _9170_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [1]),
    .B(vdd),
    .Y(_2530_)
);

INVX1 _9171_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2530_),
    .Y(_2531_)
);

AND2X2 _9172_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [2]),
    .B(gnd),
    .Y(_2532_)
);

AND2X2 _9173_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [6]),
    .Y(_2533_)
);

NAND2X1 _9174_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2532_),
    .B(_2533_),
    .Y(_2534_)
);

INVX2 _9175_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [6]),
    .Y(_2535_)
);

NAND2X1 _9176_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [2]),
    .B(gnd),
    .Y(_2536_)
);

OAI21X1 _9177_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3169_),
    .B(_2535_),
    .C(_2536_),
    .Y(_2537_)
);

NAND3X1 _9178_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2537_),
    .B(_2531_),
    .C(_2534_),
    .Y(_2538_)
);

NAND3X1 _9179_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [6]),
    .C(_2536_),
    .Y(_2539_)
);

NAND2X1 _9180_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [6]),
    .Y(_2540_)
);

NAND2X1 _9181_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2540_),
    .B(_2532_),
    .Y(_2541_)
);

NAND3X1 _9182_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2530_),
    .B(_2539_),
    .C(_2541_),
    .Y(_2542_)
);

AND2X2 _9183_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2538_),
    .B(_2542_),
    .Y(_2543_)
);

NAND2X1 _9184_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [3]),
    .Y(_2544_)
);

AOI22X1 _9185_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [2]),
    .C(gnd),
    .D(\X[3] [3]),
    .Y(_2545_)
);

OAI22X1 _9186_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2433_),
    .B(_2544_),
    .C(_2476_),
    .D(_2545_),
    .Y(_2546_)
);

NAND2X1 _9187_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[3]_5_bF$buf2 ),
    .Y(_2547_)
);

INVX1 _9188_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2547_),
    .Y(_2548_)
);

AND2X2 _9189_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [4]),
    .Y(_2549_)
);

NAND2X1 _9190_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2478_),
    .B(_2549_),
    .Y(_2550_)
);

AOI22X1 _9191_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [3]),
    .C(gnd),
    .D(\X[3] [4]),
    .Y(_2551_)
);

INVX1 _9192_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2551_),
    .Y(_2552_)
);

NAND3X1 _9193_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2548_),
    .B(_2552_),
    .C(_2550_),
    .Y(_2553_)
);

NAND3X1 _9194_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [4]),
    .C(_2544_),
    .Y(_2554_)
);

NAND2X1 _9195_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [4]),
    .Y(_2555_)
);

NAND3X1 _9196_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [3]),
    .C(_2555_),
    .Y(_2556_)
);

NAND3X1 _9197_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2547_),
    .B(_2554_),
    .C(_2556_),
    .Y(_2557_)
);

NAND3X1 _9198_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2546_),
    .B(_2557_),
    .C(_2553_),
    .Y(_2558_)
);

INVX1 _9199_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2546_),
    .Y(_2559_)
);

AOI21X1 _9200_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2554_),
    .B(_2556_),
    .C(_2547_),
    .Y(_2560_)
);

AOI22X1 _9201_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[3]_5_bF$buf1 ),
    .C(_2550_),
    .D(_2552_),
    .Y(_2561_)
);

OAI21X1 _9202_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2560_),
    .B(_2561_),
    .C(_2559_),
    .Y(_2562_)
);

NAND3X1 _9203_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2558_),
    .B(_2543_),
    .C(_2562_),
    .Y(_2563_)
);

NAND2X1 _9204_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2542_),
    .B(_2538_),
    .Y(_2564_)
);

OAI21X1 _9205_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2560_),
    .B(_2561_),
    .C(_2546_),
    .Y(_2565_)
);

NAND3X1 _9206_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2553_),
    .B(_2557_),
    .C(_2559_),
    .Y(_2566_)
);

NAND3X1 _9207_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2564_),
    .B(_2566_),
    .C(_2565_),
    .Y(_2567_)
);

NAND3X1 _9208_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2563_),
    .B(_2529_),
    .C(_2567_),
    .Y(_2568_)
);

INVX1 _9209_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2487_),
    .Y(_2569_)
);

AOI21X1 _9210_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2473_),
    .B(_2491_),
    .C(_2569_),
    .Y(_2570_)
);

AOI21X1 _9211_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2565_),
    .B(_2566_),
    .C(_2564_),
    .Y(_2571_)
);

AOI21X1 _9212_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2562_),
    .B(_2558_),
    .C(_2543_),
    .Y(_2572_)
);

OAI21X1 _9213_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2571_),
    .B(_2572_),
    .C(_2570_),
    .Y(_2573_)
);

NAND3X1 _9214_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2527_),
    .B(_2568_),
    .C(_2573_),
    .Y(_2574_)
);

AND2X2 _9215_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2525_),
    .B(_2526_),
    .Y(_2575_)
);

OAI21X1 _9216_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2571_),
    .B(_2572_),
    .C(_2529_),
    .Y(_2576_)
);

NAND3X1 _9217_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2563_),
    .B(_2567_),
    .C(_2570_),
    .Y(_2577_)
);

NAND3X1 _9218_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2575_),
    .B(_2576_),
    .C(_2577_),
    .Y(_2578_)
);

AOI22X1 _9219_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2502_),
    .B(_2497_),
    .C(_2574_),
    .D(_2578_),
    .Y(_2579_)
);

AOI21X1 _9220_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2492_),
    .B(_2496_),
    .C(_2460_),
    .Y(_2580_)
);

OAI21X1 _9221_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2503_),
    .B(_2580_),
    .C(_2497_),
    .Y(_2581_)
);

NAND3X1 _9222_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2575_),
    .B(_2568_),
    .C(_2573_),
    .Y(_2582_)
);

NAND3X1 _9223_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2527_),
    .B(_2576_),
    .C(_2577_),
    .Y(_2583_)
);

AOI21X1 _9224_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2583_),
    .B(_2582_),
    .C(_2581_),
    .Y(_2584_)
);

OAI21X1 _9225_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2584_),
    .B(_2579_),
    .C(_2507_),
    .Y(_2585_)
);

AOI21X1 _9226_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2509_),
    .B(_2508_),
    .C(_2445_),
    .Y(_2586_)
);

NAND3X1 _9227_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2581_),
    .B(_2582_),
    .C(_2583_),
    .Y(_2587_)
);

INVX1 _9228_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2497_),
    .Y(_2588_)
);

AOI21X1 _9229_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2417_),
    .B(_2501_),
    .C(_2588_),
    .Y(_2589_)
);

AOI21X1 _9230_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2577_),
    .B(_2576_),
    .C(_2527_),
    .Y(_2590_)
);

AOI21X1 _9231_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2573_),
    .B(_2568_),
    .C(_2575_),
    .Y(_2591_)
);

OAI21X1 _9232_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2590_),
    .B(_2591_),
    .C(_2589_),
    .Y(_2592_)
);

NAND3X1 _9233_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2586_),
    .B(_2587_),
    .C(_2592_),
    .Y(_2593_)
);

NAND2X1 _9234_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2593_),
    .B(_2585_),
    .Y(_2594_)
);

AOI21X1 _9235_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2511_),
    .B(_2517_),
    .C(_2594_),
    .Y(_2595_)
);

OAI21X1 _9236_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2520_),
    .B(_2518_),
    .C(_2511_),
    .Y(_2596_)
);

AOI21X1 _9237_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2585_),
    .B(_2593_),
    .C(_2596_),
    .Y(_2597_)
);

NOR2X1 _9238_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2595_),
    .B(_2597_),
    .Y(_3187_[6])
);

INVX1 _9239_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2593_),
    .Y(_2598_)
);

AOI21X1 _9240_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2563_),
    .B(_2567_),
    .C(_2529_),
    .Y(_2599_)
);

OAI21X1 _9241_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2527_),
    .B(_2599_),
    .C(_2568_),
    .Y(_2600_)
);

NAND2X1 _9242_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [0]),
    .B(gnd),
    .Y(_2601_)
);

INVX1 _9243_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2601_),
    .Y(_2602_)
);

NAND2X1 _9244_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [1]),
    .B(gnd),
    .Y(_2603_)
);

INVX1 _9245_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2603_),
    .Y(_2604_)
);

AND2X2 _9246_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2536_),
    .B(_2540_),
    .Y(_2605_)
);

OAI21X1 _9247_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2530_),
    .B(_2605_),
    .C(_2534_),
    .Y(_2606_)
);

NAND2X1 _9248_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2604_),
    .B(_2606_),
    .Y(_2607_)
);

NAND3X1 _9249_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2534_),
    .B(_2603_),
    .C(_2538_),
    .Y(_2608_)
);

NAND3X1 _9250_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2602_),
    .B(_2608_),
    .C(_2607_),
    .Y(_2609_)
);

AOI21X1 _9251_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2538_),
    .B(_2534_),
    .C(_2603_),
    .Y(_2610_)
);

NOR2X1 _9252_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2604_),
    .B(_2606_),
    .Y(_2611_)
);

OAI21X1 _9253_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2610_),
    .B(_2611_),
    .C(_2601_),
    .Y(_2612_)
);

NAND2X1 _9254_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2609_),
    .B(_2612_),
    .Y(_2613_)
);

AOI21X1 _9255_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2553_),
    .B(_2557_),
    .C(_2546_),
    .Y(_2614_)
);

OAI21X1 _9256_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2564_),
    .B(_2614_),
    .C(_2558_),
    .Y(_2615_)
);

NAND2X1 _9257_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [2]),
    .B(vdd),
    .Y(_2616_)
);

INVX1 _9258_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2616_),
    .Y(_2617_)
);

AND2X2 _9259_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [3]),
    .B(gnd),
    .Y(_2618_)
);

AND2X2 _9260_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [7]),
    .Y(_2619_)
);

NAND2X1 _9261_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2618_),
    .B(_2619_),
    .Y(_2620_)
);

AOI22X1 _9262_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [7]),
    .C(\X[3] [3]),
    .D(gnd),
    .Y(_2621_)
);

INVX1 _9263_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2621_),
    .Y(_2622_)
);

NAND3X1 _9264_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2617_),
    .B(_2622_),
    .C(_2620_),
    .Y(_2623_)
);

INVX1 _9265_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_2624_)
);

OAI21X1 _9266_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2406_),
    .B(_2624_),
    .C(_2619_),
    .Y(_2625_)
);

INVX1 _9267_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [7]),
    .Y(_2626_)
);

OAI21X1 _9268_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3169_),
    .B(_2626_),
    .C(_2618_),
    .Y(_2627_)
);

NAND3X1 _9269_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2616_),
    .B(_2625_),
    .C(_2627_),
    .Y(_2628_)
);

NAND2X1 _9270_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2623_),
    .B(_2628_),
    .Y(_2629_)
);

OAI21X1 _9271_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2547_),
    .B(_2551_),
    .C(_2550_),
    .Y(_2630_)
);

NAND2X1 _9272_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[3] [6]),
    .Y(_2631_)
);

NAND2X1 _9273_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [4]),
    .Y(_2632_)
);

AND2X2 _9274_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3]_5_bF$buf0 ),
    .Y(_2633_)
);

NAND2X1 _9275_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2632_),
    .B(_2633_),
    .Y(_2634_)
);

OAI21X1 _9276_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2480_),
    .B(_2465_),
    .C(_2549_),
    .Y(_2635_)
);

AOI21X1 _9277_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2635_),
    .B(_2634_),
    .C(_2631_),
    .Y(_2636_)
);

INVX1 _9278_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2631_),
    .Y(_2637_)
);

NAND2X1 _9279_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2549_),
    .B(_2633_),
    .Y(_2638_)
);

AOI22X1 _9280_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [4]),
    .C(gnd),
    .D(\X[3]_5_bF$buf3 ),
    .Y(_2639_)
);

INVX1 _9281_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2639_),
    .Y(_2640_)
);

AOI21X1 _9282_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2638_),
    .B(_2640_),
    .C(_2637_),
    .Y(_2641_)
);

OAI21X1 _9283_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2641_),
    .B(_2636_),
    .C(_2630_),
    .Y(_2642_)
);

AOI22X1 _9284_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2478_),
    .B(_2549_),
    .C(_2552_),
    .D(_2548_),
    .Y(_2643_)
);

NAND3X1 _9285_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2637_),
    .B(_2640_),
    .C(_2638_),
    .Y(_2644_)
);

NAND2X1 _9286_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3]_5_bF$buf2 ),
    .Y(_2645_)
);

NOR2X1 _9287_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2632_),
    .B(_2645_),
    .Y(_2646_)
);

OAI21X1 _9288_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2639_),
    .B(_2646_),
    .C(_2631_),
    .Y(_2647_)
);

NAND3X1 _9289_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2644_),
    .B(_2643_),
    .C(_2647_),
    .Y(_2648_)
);

AOI21X1 _9290_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2642_),
    .B(_2648_),
    .C(_2629_),
    .Y(_2649_)
);

AND2X2 _9291_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2628_),
    .B(_2623_),
    .Y(_2650_)
);

NAND3X1 _9292_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2630_),
    .B(_2644_),
    .C(_2647_),
    .Y(_2651_)
);

OAI21X1 _9293_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2641_),
    .B(_2636_),
    .C(_2643_),
    .Y(_2652_)
);

AOI21X1 _9294_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2652_),
    .B(_2651_),
    .C(_2650_),
    .Y(_2653_)
);

OAI21X1 _9295_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2649_),
    .B(_2653_),
    .C(_2615_),
    .Y(_2654_)
);

INVX1 _9296_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2558_),
    .Y(_2655_)
);

AOI21X1 _9297_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2543_),
    .B(_2562_),
    .C(_2655_),
    .Y(_2656_)
);

NAND3X1 _9298_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2651_),
    .B(_2650_),
    .C(_2652_),
    .Y(_2657_)
);

NAND3X1 _9299_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2629_),
    .B(_2648_),
    .C(_2642_),
    .Y(_2658_)
);

NAND3X1 _9300_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2657_),
    .B(_2658_),
    .C(_2656_),
    .Y(_2659_)
);

AOI21X1 _9301_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2659_),
    .B(_2654_),
    .C(_2613_),
    .Y(_2660_)
);

AND2X2 _9302_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2612_),
    .B(_2609_),
    .Y(_2661_)
);

NAND3X1 _9303_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2615_),
    .B(_2657_),
    .C(_2658_),
    .Y(_2662_)
);

OAI21X1 _9304_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2649_),
    .B(_2653_),
    .C(_2656_),
    .Y(_2663_)
);

AOI21X1 _9305_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2663_),
    .B(_2662_),
    .C(_2661_),
    .Y(_2664_)
);

OAI21X1 _9306_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2664_),
    .B(_2660_),
    .C(_2600_),
    .Y(_2665_)
);

INVX1 _9307_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2568_),
    .Y(_2666_)
);

AOI21X1 _9308_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2575_),
    .B(_2573_),
    .C(_2666_),
    .Y(_2667_)
);

NAND3X1 _9309_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2662_),
    .B(_2661_),
    .C(_2663_),
    .Y(_2668_)
);

NAND3X1 _9310_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2613_),
    .B(_2654_),
    .C(_2659_),
    .Y(_2669_)
);

NAND3X1 _9311_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2668_),
    .B(_2669_),
    .C(_2667_),
    .Y(_2670_)
);

AOI21X1 _9312_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2670_),
    .B(_2665_),
    .C(_2526_),
    .Y(_2671_)
);

INVX1 _9313_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2526_),
    .Y(_2672_)
);

NAND3X1 _9314_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2600_),
    .B(_2668_),
    .C(_2669_),
    .Y(_2673_)
);

OAI21X1 _9315_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2660_),
    .B(_2664_),
    .C(_2667_),
    .Y(_2674_)
);

AOI21X1 _9316_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2674_),
    .B(_2673_),
    .C(_2672_),
    .Y(_2675_)
);

OAI21X1 _9317_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2675_),
    .B(_2671_),
    .C(_2587_),
    .Y(_2676_)
);

NAND3X1 _9318_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2672_),
    .B(_2673_),
    .C(_2674_),
    .Y(_2677_)
);

NAND3X1 _9319_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2526_),
    .B(_2665_),
    .C(_2670_),
    .Y(_2678_)
);

NAND3X1 _9320_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2579_),
    .B(_2677_),
    .C(_2678_),
    .Y(_2679_)
);

AND2X2 _9321_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2676_),
    .B(_2679_),
    .Y(_2680_)
);

OAI21X1 _9322_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2598_),
    .B(_2595_),
    .C(_2680_),
    .Y(_2681_)
);

NOR2X1 _9323_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2598_),
    .B(_2595_),
    .Y(_2682_)
);

AOI21X1 _9324_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2678_),
    .B(_2677_),
    .C(_2579_),
    .Y(_2683_)
);

INVX1 _9325_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2679_),
    .Y(_2684_)
);

OAI21X1 _9326_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2683_),
    .B(_2684_),
    .C(_2682_),
    .Y(_2685_)
);

AND2X2 _9327_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2685_),
    .B(_2681_),
    .Y(_3187_[7])
);

NAND3X1 _9328_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2676_),
    .B(_2679_),
    .C(_2595_),
    .Y(_2686_)
);

AOI21X1 _9329_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2598_),
    .B(_2676_),
    .C(_2684_),
    .Y(_2687_)
);

NAND2X1 _9330_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2687_),
    .B(_2686_),
    .Y(_2688_)
);

INVX1 _9331_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2673_),
    .Y(_2689_)
);

AOI21X1 _9332_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2672_),
    .B(_2674_),
    .C(_2689_),
    .Y(_2690_)
);

OAI21X1 _9333_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2601_),
    .B(_2611_),
    .C(_2607_),
    .Y(_2691_)
);

INVX1 _9334_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2691_),
    .Y(_2692_)
);

AOI21X1 _9335_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2657_),
    .B(_2658_),
    .C(_2615_),
    .Y(_2693_)
);

OAI21X1 _9336_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2613_),
    .B(_2693_),
    .C(_2662_),
    .Y(_2694_)
);

NAND2X1 _9337_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [1]),
    .B(gnd),
    .Y(_2695_)
);

INVX2 _9338_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_2696_)
);

NOR2X1 _9339_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3161_),
    .B(_2696_),
    .Y(_2697_)
);

OAI21X1 _9340_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2616_),
    .B(_2621_),
    .C(_2620_),
    .Y(_2698_)
);

NOR2X1 _9341_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2697_),
    .B(_2698_),
    .Y(_2699_)
);

AND2X2 _9342_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2698_),
    .B(_2697_),
    .Y(_2700_)
);

OAI21X1 _9343_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2699_),
    .B(_2700_),
    .C(_2695_),
    .Y(_2701_)
);

INVX1 _9344_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2695_),
    .Y(_2702_)
);

OR2X2 _9345_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2698_),
    .B(_2697_),
    .Y(_2703_)
);

NAND2X1 _9346_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2697_),
    .B(_2698_),
    .Y(_2704_)
);

NAND3X1 _9347_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2702_),
    .B(_2704_),
    .C(_2703_),
    .Y(_2705_)
);

NAND2X1 _9348_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2701_),
    .B(_2705_),
    .Y(_2706_)
);

AOI21X1 _9349_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2647_),
    .B(_2644_),
    .C(_2630_),
    .Y(_2707_)
);

OAI21X1 _9350_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2629_),
    .B(_2707_),
    .C(_2651_),
    .Y(_2708_)
);

NAND2X1 _9351_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [3]),
    .B(gnd),
    .Y(_2709_)
);

INVX1 _9352_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .Y(_2710_)
);

OAI21X1 _9353_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2406_),
    .B(_2710_),
    .C(_2416_),
    .Y(_2711_)
);

NAND2X1 _9354_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [4]),
    .B(vdd),
    .Y(_2712_)
);

OAI21X1 _9355_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2709_),
    .B(_2712_),
    .C(_2711_),
    .Y(_2713_)
);

OAI21X1 _9356_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2631_),
    .B(_2639_),
    .C(_2638_),
    .Y(_2714_)
);

NAND2X1 _9357_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[3] [7]),
    .Y(_2715_)
);

NAND2X1 _9358_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3]_5_bF$buf1 ),
    .Y(_2716_)
);

NAND3X1 _9359_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [6]),
    .C(_2716_),
    .Y(_2717_)
);

AND2X2 _9360_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3]_5_bF$buf0 ),
    .Y(_2718_)
);

OAI21X1 _9361_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2480_),
    .B(_2535_),
    .C(_2718_),
    .Y(_2719_)
);

AOI21X1 _9362_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2719_),
    .B(_2717_),
    .C(_2715_),
    .Y(_2720_)
);

INVX1 _9363_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2715_),
    .Y(_2721_)
);

AND2X2 _9364_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [6]),
    .Y(_2722_)
);

NAND2X1 _9365_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2718_),
    .B(_2722_),
    .Y(_2723_)
);

NAND2X1 _9366_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [6]),
    .Y(_2724_)
);

NAND2X1 _9367_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2716_),
    .B(_2724_),
    .Y(_2725_)
);

AOI21X1 _9368_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2723_),
    .B(_2725_),
    .C(_2721_),
    .Y(_2726_)
);

OAI21X1 _9369_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2726_),
    .B(_2720_),
    .C(_2714_),
    .Y(_2727_)
);

AOI21X1 _9370_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2637_),
    .B(_2640_),
    .C(_2646_),
    .Y(_2728_)
);

NAND3X1 _9371_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2721_),
    .B(_2725_),
    .C(_2723_),
    .Y(_2729_)
);

NAND3X1 _9372_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2715_),
    .B(_2717_),
    .C(_2719_),
    .Y(_2730_)
);

NAND3X1 _9373_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2729_),
    .B(_2730_),
    .C(_2728_),
    .Y(_2731_)
);

AOI21X1 _9374_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2727_),
    .B(_2731_),
    .C(_2713_),
    .Y(_2732_)
);

INVX1 _9375_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2713_),
    .Y(_2733_)
);

NAND3X1 _9376_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2714_),
    .B(_2729_),
    .C(_2730_),
    .Y(_2734_)
);

OAI21X1 _9377_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2726_),
    .B(_2720_),
    .C(_2728_),
    .Y(_2735_)
);

AOI21X1 _9378_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2735_),
    .B(_2734_),
    .C(_2733_),
    .Y(_2736_)
);

OAI21X1 _9379_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2732_),
    .B(_2736_),
    .C(_2708_),
    .Y(_2737_)
);

INVX1 _9380_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2651_),
    .Y(_2738_)
);

AOI21X1 _9381_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2650_),
    .B(_2652_),
    .C(_2738_),
    .Y(_2739_)
);

NAND3X1 _9382_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2733_),
    .B(_2734_),
    .C(_2735_),
    .Y(_2740_)
);

NAND3X1 _9383_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2713_),
    .B(_2731_),
    .C(_2727_),
    .Y(_2741_)
);

NAND3X1 _9384_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2740_),
    .B(_2741_),
    .C(_2739_),
    .Y(_2742_)
);

AOI21X1 _9385_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2742_),
    .B(_2737_),
    .C(_2706_),
    .Y(_2743_)
);

AND2X2 _9386_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2705_),
    .B(_2701_),
    .Y(_2744_)
);

NAND3X1 _9387_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2740_),
    .B(_2741_),
    .C(_2708_),
    .Y(_2745_)
);

OAI21X1 _9388_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2732_),
    .B(_2736_),
    .C(_2739_),
    .Y(_2746_)
);

AOI21X1 _9389_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2746_),
    .B(_2745_),
    .C(_2744_),
    .Y(_2747_)
);

OAI21X1 _9390_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2747_),
    .B(_2743_),
    .C(_2694_),
    .Y(_2748_)
);

INVX1 _9391_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2662_),
    .Y(_2749_)
);

AOI21X1 _9392_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2661_),
    .B(_2663_),
    .C(_2749_),
    .Y(_2750_)
);

NAND3X1 _9393_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2744_),
    .B(_2745_),
    .C(_2746_),
    .Y(_2751_)
);

NAND3X1 _9394_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2706_),
    .B(_2737_),
    .C(_2742_),
    .Y(_2752_)
);

NAND3X1 _9395_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2751_),
    .B(_2752_),
    .C(_2750_),
    .Y(_2753_)
);

AOI21X1 _9396_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2748_),
    .B(_2753_),
    .C(_2692_),
    .Y(_2754_)
);

NAND3X1 _9397_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2694_),
    .B(_2751_),
    .C(_2752_),
    .Y(_2755_)
);

OAI21X1 _9398_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2747_),
    .B(_2743_),
    .C(_2750_),
    .Y(_2756_)
);

AOI21X1 _9399_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2756_),
    .B(_2755_),
    .C(_2691_),
    .Y(_2757_)
);

OAI21X1 _9400_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2757_),
    .B(_2754_),
    .C(_2690_),
    .Y(_2758_)
);

AOI21X1 _9401_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2669_),
    .B(_2668_),
    .C(_2600_),
    .Y(_2759_)
);

OAI21X1 _9402_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2526_),
    .B(_2759_),
    .C(_2673_),
    .Y(_2760_)
);

NAND3X1 _9403_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2691_),
    .B(_2755_),
    .C(_2756_),
    .Y(_2761_)
);

NAND3X1 _9404_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2692_),
    .B(_2753_),
    .C(_2748_),
    .Y(_2762_)
);

NAND3X1 _9405_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2760_),
    .B(_2761_),
    .C(_2762_),
    .Y(_2763_)
);

NAND2X1 _9406_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2763_),
    .B(_2758_),
    .Y(_2764_)
);

NAND2X1 _9407_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2764_),
    .B(_2688_),
    .Y(_2765_)
);

OAI21X1 _9408_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2593_),
    .B(_2683_),
    .C(_2679_),
    .Y(_2766_)
);

AOI21X1 _9409_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2680_),
    .B(_2595_),
    .C(_2766_),
    .Y(_2767_)
);

AND2X2 _9410_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2758_),
    .B(_2763_),
    .Y(_2768_)
);

NAND2X1 _9411_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2768_),
    .B(_2767_),
    .Y(_2769_)
);

NAND2X1 _9412_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2765_),
    .B(_2769_),
    .Y(_3187_[8])
);

INVX1 _9413_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2763_),
    .Y(_2770_)
);

AOI21X1 _9414_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2688_),
    .B(_2758_),
    .C(_2770_),
    .Y(_2771_)
);

AOI21X1 _9415_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2752_),
    .B(_2751_),
    .C(_2694_),
    .Y(_2772_)
);

OAI21X1 _9416_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2692_),
    .B(_2772_),
    .C(_2755_),
    .Y(_2773_)
);

OAI21X1 _9417_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2695_),
    .B(_2699_),
    .C(_2704_),
    .Y(_2774_)
);

AOI21X1 _9418_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2740_),
    .B(_2741_),
    .C(_2708_),
    .Y(_2775_)
);

OAI21X1 _9419_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2706_),
    .B(_2775_),
    .C(_2745_),
    .Y(_2776_)
);

NAND2X1 _9420_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [2]),
    .B(gnd),
    .Y(_2777_)
);

NOR2X1 _9421_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2709_),
    .B(_2712_),
    .Y(_2778_)
);

NAND2X1 _9422_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_2778_),
    .Y(_2779_)
);

INVX1 _9423_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2779_),
    .Y(_2780_)
);

AOI21X1 _9424_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [3]),
    .B(gnd),
    .C(_2778_),
    .Y(_2781_)
);

OAI21X1 _9425_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2781_),
    .B(_2780_),
    .C(_2777_),
    .Y(_2782_)
);

INVX1 _9426_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2777_),
    .Y(_2783_)
);

INVX1 _9427_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2781_),
    .Y(_2784_)
);

NAND3X1 _9428_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2783_),
    .B(_2779_),
    .C(_2784_),
    .Y(_2785_)
);

AND2X2 _9429_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2785_),
    .B(_2782_),
    .Y(_2786_)
);

AOI21X1 _9430_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2730_),
    .B(_2729_),
    .C(_2714_),
    .Y(_2787_)
);

OAI21X1 _9431_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2713_),
    .B(_2787_),
    .C(_2734_),
    .Y(_2788_)
);

NOR2X1 _9432_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2523_),
    .B(_2712_),
    .Y(_2789_)
);

AND2X2 _9433_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2523_),
    .B(_2712_),
    .Y(_2790_)
);

NOR2X1 _9434_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2789_),
    .B(_2790_),
    .Y(_2791_)
);

NAND2X1 _9435_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [6]),
    .Y(_2792_)
);

AOI22X1 _9436_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3]_5_bF$buf3 ),
    .C(gnd),
    .D(\X[3] [6]),
    .Y(_2793_)
);

OAI22X1 _9437_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2645_),
    .B(_2792_),
    .C(_2715_),
    .D(_2793_),
    .Y(_2794_)
);

AOI22X1 _9438_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [6]),
    .C(gnd),
    .D(\X[3] [7]),
    .Y(_2795_)
);

AND2X2 _9439_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [7]),
    .Y(_2796_)
);

AOI21X1 _9440_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2722_),
    .B(_2796_),
    .C(_2795_),
    .Y(_2797_)
);

NAND2X1 _9441_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2797_),
    .B(_2794_),
    .Y(_2798_)
);

AND2X2 _9442_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [6]),
    .Y(_2799_)
);

AOI22X1 _9443_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2633_),
    .B(_2799_),
    .C(_2725_),
    .D(_2721_),
    .Y(_2800_)
);

NAND2X1 _9444_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [7]),
    .Y(_2801_)
);

NAND2X1 _9445_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2792_),
    .B(_2801_),
    .Y(_2802_)
);

NAND2X1 _9446_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [7]),
    .Y(_2803_)
);

OAI21X1 _9447_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2724_),
    .B(_2803_),
    .C(_2802_),
    .Y(_2804_)
);

NAND2X1 _9448_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2804_),
    .B(_2800_),
    .Y(_2805_)
);

NAND3X1 _9449_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2791_),
    .B(_2798_),
    .C(_2805_),
    .Y(_2806_)
);

NAND2X1 _9450_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3]_5_bF$buf2 ),
    .B(vdd),
    .Y(_2807_)
);

INVX1 _9451_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [4]),
    .Y(_2808_)
);

OAI21X1 _9452_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2808_),
    .B(_2710_),
    .C(_2523_),
    .Y(_2809_)
);

OAI21X1 _9453_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2416_),
    .B(_2807_),
    .C(_2809_),
    .Y(_2810_)
);

NAND2X1 _9454_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2794_),
    .B(_2804_),
    .Y(_2811_)
);

NAND2X1 _9455_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2797_),
    .B(_2800_),
    .Y(_2812_)
);

NAND3X1 _9456_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2810_),
    .B(_2811_),
    .C(_2812_),
    .Y(_2813_)
);

NAND3X1 _9457_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2806_),
    .B(_2813_),
    .C(_2788_),
    .Y(_2814_)
);

NAND2X1 _9458_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2806_),
    .B(_2813_),
    .Y(_2815_)
);

NAND3X1 _9459_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2734_),
    .B(_2740_),
    .C(_2815_),
    .Y(_2816_)
);

NAND3X1 _9460_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2786_),
    .B(_2814_),
    .C(_2816_),
    .Y(_2817_)
);

NAND2X1 _9461_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2782_),
    .B(_2785_),
    .Y(_2818_)
);

AOI21X1 _9462_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2734_),
    .B(_2740_),
    .C(_2815_),
    .Y(_2819_)
);

AOI21X1 _9463_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2806_),
    .B(_2813_),
    .C(_2788_),
    .Y(_2820_)
);

OAI21X1 _9464_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2820_),
    .B(_2819_),
    .C(_2818_),
    .Y(_2821_)
);

NAND3X1 _9465_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2817_),
    .B(_2821_),
    .C(_2776_),
    .Y(_2822_)
);

INVX1 _9466_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2745_),
    .Y(_2823_)
);

AOI21X1 _9467_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2744_),
    .B(_2746_),
    .C(_2823_),
    .Y(_2824_)
);

INVX1 _9468_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2817_),
    .Y(_2825_)
);

AOI21X1 _9469_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2816_),
    .B(_2814_),
    .C(_2786_),
    .Y(_2826_)
);

OAI21X1 _9470_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2826_),
    .B(_2825_),
    .C(_2824_),
    .Y(_2827_)
);

NAND3X1 _9471_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2774_),
    .B(_2822_),
    .C(_2827_),
    .Y(_2828_)
);

INVX1 _9472_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2774_),
    .Y(_2829_)
);

INVX1 _9473_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2822_),
    .Y(_2830_)
);

AOI21X1 _9474_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2821_),
    .B(_2817_),
    .C(_2776_),
    .Y(_2831_)
);

OAI21X1 _9475_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2831_),
    .B(_2830_),
    .C(_2829_),
    .Y(_2832_)
);

NAND3X1 _9476_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2773_),
    .B(_2828_),
    .C(_2832_),
    .Y(_2833_)
);

INVX1 _9477_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2755_),
    .Y(_2834_)
);

AOI21X1 _9478_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2691_),
    .B(_2756_),
    .C(_2834_),
    .Y(_2835_)
);

OAI21X1 _9479_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2826_),
    .B(_2825_),
    .C(_2776_),
    .Y(_2836_)
);

NAND3X1 _9480_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2817_),
    .B(_2821_),
    .C(_2824_),
    .Y(_2837_)
);

AOI21X1 _9481_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2837_),
    .B(_2836_),
    .C(_2829_),
    .Y(_2838_)
);

AOI21X1 _9482_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2827_),
    .B(_2822_),
    .C(_2774_),
    .Y(_2839_)
);

OAI21X1 _9483_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2838_),
    .B(_2839_),
    .C(_2835_),
    .Y(_2840_)
);

AND2X2 _9484_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2840_),
    .B(_2833_),
    .Y(_2841_)
);

OR2X2 _9485_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2771_),
    .B(_2841_),
    .Y(_2842_)
);

NAND2X1 _9486_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2841_),
    .B(_2771_),
    .Y(_2843_)
);

NAND2X1 _9487_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2843_),
    .B(_2842_),
    .Y(_3187_[9])
);

NAND2X1 _9488_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2833_),
    .B(_2840_),
    .Y(_2844_)
);

NOR2X1 _9489_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2764_),
    .B(_2844_),
    .Y(_2845_)
);

NAND2X1 _9490_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2845_),
    .B(_2688_),
    .Y(_2846_)
);

AOI21X1 _9491_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2832_),
    .B(_2828_),
    .C(_2773_),
    .Y(_2847_)
);

AOI21X1 _9492_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2763_),
    .B(_2833_),
    .C(_2847_),
    .Y(_2848_)
);

INVX1 _9493_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2848_),
    .Y(_2849_)
);

OAI21X1 _9494_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2829_),
    .B(_2831_),
    .C(_2822_),
    .Y(_2850_)
);

OAI21X1 _9495_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2777_),
    .B(_2781_),
    .C(_2779_),
    .Y(_2851_)
);

OAI21X1 _9496_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2818_),
    .B(_2820_),
    .C(_2814_),
    .Y(_2852_)
);

INVX2 _9497_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_2853_)
);

NOR3X1 _9498_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2696_),
    .B(_2523_),
    .C(_2712_),
    .Y(_2854_)
);

OAI22X1 _9499_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2808_),
    .B(_2696_),
    .C(_2416_),
    .D(_2807_),
    .Y(_2855_)
);

INVX1 _9500_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2855_),
    .Y(_2856_)
);

OAI22X1 _9501_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2406_),
    .B(_2853_),
    .C(_2854_),
    .D(_2856_),
    .Y(_2857_)
);

NOR2X1 _9502_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2406_),
    .B(_2853_),
    .Y(_2858_)
);

NAND2X1 _9503_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_2789_),
    .Y(_2859_)
);

NAND3X1 _9504_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2858_),
    .B(_2855_),
    .C(_2859_),
    .Y(_2860_)
);

AND2X2 _9505_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2857_),
    .B(_2860_),
    .Y(_2861_)
);

NOR2X1 _9506_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2797_),
    .B(_2794_),
    .Y(_2862_)
);

OAI21X1 _9507_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2810_),
    .B(_2862_),
    .C(_2798_),
    .Y(_2863_)
);

NAND2X1 _9508_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [6]),
    .Y(_2864_)
);

NOR2X1 _9509_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2864_),
    .B(_2807_),
    .Y(_2865_)
);

AND2X2 _9510_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2864_),
    .B(_2807_),
    .Y(_2866_)
);

OAI22X1 _9511_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2722_),
    .B(_2803_),
    .C(_2865_),
    .D(_2866_),
    .Y(_2867_)
);

AND2X2 _9512_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [6]),
    .Y(_2868_)
);

AND2X2 _9513_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3]_5_bF$buf1 ),
    .B(vdd),
    .Y(_2869_)
);

NAND2X1 _9514_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2868_),
    .B(_2869_),
    .Y(_2870_)
);

OAI21X1 _9515_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2465_),
    .B(_2710_),
    .C(_2864_),
    .Y(_2871_)
);

AOI21X1 _9516_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[3] [6]),
    .C(_2803_),
    .Y(_2872_)
);

NAND3X1 _9517_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2871_),
    .B(_2872_),
    .C(_2870_),
    .Y(_2873_)
);

AND2X2 _9518_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2867_),
    .B(_2873_),
    .Y(_2874_)
);

NAND2X1 _9519_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2874_),
    .B(_2863_),
    .Y(_2875_)
);

NAND2X1 _9520_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2873_),
    .B(_2867_),
    .Y(_2876_)
);

NAND3X1 _9521_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2798_),
    .B(_2876_),
    .C(_2806_),
    .Y(_2877_)
);

NAND3X1 _9522_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2861_),
    .B(_2877_),
    .C(_2875_),
    .Y(_2878_)
);

NAND2X1 _9523_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2860_),
    .B(_2857_),
    .Y(_2879_)
);

NAND2X1 _9524_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2876_),
    .B(_2863_),
    .Y(_2880_)
);

NAND3X1 _9525_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2798_),
    .B(_2874_),
    .C(_2806_),
    .Y(_2881_)
);

NAND3X1 _9526_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2879_),
    .B(_2881_),
    .C(_2880_),
    .Y(_2882_)
);

NAND3X1 _9527_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2878_),
    .B(_2882_),
    .C(_2852_),
    .Y(_2883_)
);

NAND2X1 _9528_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2882_),
    .B(_2878_),
    .Y(_2884_)
);

NAND3X1 _9529_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2814_),
    .B(_2817_),
    .C(_2884_),
    .Y(_2885_)
);

NAND3X1 _9530_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2851_),
    .B(_2885_),
    .C(_2883_),
    .Y(_2886_)
);

INVX1 _9531_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2851_),
    .Y(_2887_)
);

NAND2X1 _9532_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2884_),
    .B(_2852_),
    .Y(_2888_)
);

AOI21X1 _9533_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2786_),
    .B(_2816_),
    .C(_2819_),
    .Y(_2889_)
);

AND2X2 _9534_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2878_),
    .B(_2882_),
    .Y(_2890_)
);

NAND2X1 _9535_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2889_),
    .B(_2890_),
    .Y(_2891_)
);

NAND3X1 _9536_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2887_),
    .B(_2888_),
    .C(_2891_),
    .Y(_2892_)
);

AOI21X1 _9537_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2886_),
    .B(_2892_),
    .C(_2850_),
    .Y(_2893_)
);

NAND2X1 _9538_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2886_),
    .B(_2892_),
    .Y(_2894_)
);

AOI21X1 _9539_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2822_),
    .B(_2828_),
    .C(_2894_),
    .Y(_2895_)
);

NOR2X1 _9540_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2893_),
    .B(_2895_),
    .Y(_2896_)
);

INVX1 _9541_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2896_),
    .Y(_2897_)
);

AOI21X1 _9542_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2846_),
    .B(_2849_),
    .C(_2897_),
    .Y(_2898_)
);

NAND2X1 _9543_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2768_),
    .B(_2841_),
    .Y(_2899_)
);

OAI21X1 _9544_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2899_),
    .B(_2767_),
    .C(_2849_),
    .Y(_2900_)
);

NOR2X1 _9545_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2896_),
    .B(_2900_),
    .Y(_2901_)
);

NOR2X1 _9546_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2898_),
    .B(_2901_),
    .Y(_3187_[10])
);

NAND3X1 _9547_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2886_),
    .B(_2892_),
    .C(_2850_),
    .Y(_2902_)
);

NAND2X1 _9548_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2896_),
    .B(_2900_),
    .Y(_2903_)
);

NOR2X1 _9549_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2884_),
    .B(_2889_),
    .Y(_2904_)
);

AOI21X1 _9550_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2851_),
    .B(_2885_),
    .C(_2904_),
    .Y(_2905_)
);

NAND2X1 _9551_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2859_),
    .B(_2860_),
    .Y(_2906_)
);

NAND2X1 _9552_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2875_),
    .B(_2878_),
    .Y(_2907_)
);

NOR3X1 _9553_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2696_),
    .B(_2864_),
    .C(_2807_),
    .Y(_2908_)
);

AOI22X1 _9554_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3]_5_bF$buf0 ),
    .B(gnd),
    .C(_2868_),
    .D(_2869_),
    .Y(_2909_)
);

OAI22X1 _9555_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2808_),
    .B(_2853_),
    .C(_2909_),
    .D(_2908_),
    .Y(_2910_)
);

NOR2X1 _9556_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2808_),
    .B(_2853_),
    .Y(_2911_)
);

NAND2X1 _9557_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_2865_),
    .Y(_2912_)
);

OAI21X1 _9558_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2465_),
    .B(_2696_),
    .C(_2870_),
    .Y(_2913_)
);

NAND3X1 _9559_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2911_),
    .B(_2912_),
    .C(_2913_),
    .Y(_2914_)
);

NAND2X1 _9560_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2910_),
    .B(_2914_),
    .Y(_2915_)
);

NAND2X1 _9561_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2722_),
    .B(_2796_),
    .Y(_2916_)
);

NAND2X1 _9562_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[3] [7]),
    .Y(_2917_)
);

OAI22X1 _9563_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2624_),
    .B(_2626_),
    .C(_2710_),
    .D(_2535_),
    .Y(_2918_)
);

OAI21X1 _9564_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2864_),
    .B(_2917_),
    .C(_2918_),
    .Y(_2919_)
);

NAND3X1 _9565_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2916_),
    .B(_2919_),
    .C(_2873_),
    .Y(_2920_)
);

INVX1 _9566_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2920_),
    .Y(_2921_)
);

AOI21X1 _9567_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2873_),
    .B(_2916_),
    .C(_2919_),
    .Y(_2922_)
);

OAI21X1 _9568_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2922_),
    .B(_2921_),
    .C(_2915_),
    .Y(_2923_)
);

AND2X2 _9569_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2914_),
    .B(_2910_),
    .Y(_2924_)
);

INVX1 _9570_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2922_),
    .Y(_2925_)
);

NAND3X1 _9571_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2920_),
    .B(_2925_),
    .C(_2924_),
    .Y(_2926_)
);

AND2X2 _9572_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2926_),
    .B(_2923_),
    .Y(_2927_)
);

NAND2X1 _9573_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2927_),
    .B(_2907_),
    .Y(_2928_)
);

AOI21X1 _9574_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2806_),
    .B(_2798_),
    .C(_2876_),
    .Y(_2929_)
);

AOI21X1 _9575_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2861_),
    .B(_2877_),
    .C(_2929_),
    .Y(_2930_)
);

NAND2X1 _9576_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2923_),
    .B(_2926_),
    .Y(_2931_)
);

NAND2X1 _9577_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2931_),
    .B(_2930_),
    .Y(_2932_)
);

NAND3X1 _9578_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2906_),
    .B(_2932_),
    .C(_2928_),
    .Y(_2933_)
);

INVX1 _9579_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2906_),
    .Y(_2934_)
);

NAND2X1 _9580_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2931_),
    .B(_2907_),
    .Y(_2935_)
);

NAND2X1 _9581_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2930_),
    .B(_2927_),
    .Y(_2936_)
);

NAND3X1 _9582_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2934_),
    .B(_2936_),
    .C(_2935_),
    .Y(_2937_)
);

NAND2X1 _9583_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2933_),
    .B(_2937_),
    .Y(_2938_)
);

NAND2X1 _9584_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2938_),
    .B(_2905_),
    .Y(_2939_)
);

AOI21X1 _9585_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2878_),
    .B(_2882_),
    .C(_2852_),
    .Y(_2940_)
);

OAI21X1 _9586_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2887_),
    .B(_2940_),
    .C(_2883_),
    .Y(_2941_)
);

NAND3X1 _9587_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2933_),
    .B(_2937_),
    .C(_2941_),
    .Y(_2942_)
);

NAND2X1 _9588_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2939_),
    .B(_2942_),
    .Y(_2943_)
);

INVX1 _9589_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2943_),
    .Y(_2944_)
);

NAND3X1 _9590_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2902_),
    .B(_2944_),
    .C(_2903_),
    .Y(_2945_)
);

OAI21X1 _9591_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2895_),
    .B(_2898_),
    .C(_2943_),
    .Y(_2946_)
);

NAND2X1 _9592_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2945_),
    .B(_2946_),
    .Y(_3187_[11])
);

NOR3X1 _9593_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2893_),
    .B(_2895_),
    .C(_2943_),
    .Y(_2947_)
);

NAND3X1 _9594_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2845_),
    .B(_2947_),
    .C(_2688_),
    .Y(_2948_)
);

OAI21X1 _9595_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2902_),
    .B(_2943_),
    .C(_2942_),
    .Y(_2949_)
);

AOI21X1 _9596_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2947_),
    .B(_2848_),
    .C(_2949_),
    .Y(_2950_)
);

AND2X2 _9597_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2933_),
    .B(_2928_),
    .Y(_2951_)
);

OAI21X1 _9598_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2696_),
    .B(_2870_),
    .C(_2914_),
    .Y(_2952_)
);

OAI21X1 _9599_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2921_),
    .B(_2915_),
    .C(_2925_),
    .Y(_2953_)
);

INVX1 _9600_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2953_),
    .Y(_2954_)
);

INVX1 _9601_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2917_),
    .Y(_2955_)
);

NOR2X1 _9602_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2465_),
    .B(_2853_),
    .Y(_2956_)
);

NOR2X1 _9603_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2864_),
    .B(_2917_),
    .Y(_2957_)
);

NOR2X1 _9604_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2535_),
    .B(_2696_),
    .Y(_2958_)
);

NOR2X1 _9605_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2958_),
    .B(_2957_),
    .Y(_2959_)
);

AOI21X1 _9606_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(_2957_),
    .C(_2959_),
    .Y(_2960_)
);

OR2X2 _9607_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2960_),
    .B(_2956_),
    .Y(_2961_)
);

NAND2X1 _9608_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2956_),
    .B(_2960_),
    .Y(_2962_)
);

NAND3X1 _9609_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2955_),
    .B(_2962_),
    .C(_2961_),
    .Y(_2963_)
);

NOR2X1 _9610_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2956_),
    .B(_2960_),
    .Y(_2964_)
);

INVX1 _9611_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2962_),
    .Y(_2965_)
);

OAI21X1 _9612_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2964_),
    .B(_2965_),
    .C(_2917_),
    .Y(_2966_)
);

NAND2X1 _9613_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2963_),
    .B(_2966_),
    .Y(_2967_)
);

NAND2X1 _9614_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2954_),
    .B(_2967_),
    .Y(_2968_)
);

NAND3X1 _9615_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2953_),
    .B(_2963_),
    .C(_2966_),
    .Y(_2969_)
);

AOI21X1 _9616_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2968_),
    .B(_2969_),
    .C(_2952_),
    .Y(_2970_)
);

NAND3X1 _9617_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2952_),
    .B(_2969_),
    .C(_2968_),
    .Y(_2971_)
);

INVX1 _9618_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2971_),
    .Y(_2972_)
);

OAI21X1 _9619_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2970_),
    .B(_2972_),
    .C(_2951_),
    .Y(_2973_)
);

OR2X2 _9620_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2972_),
    .B(_2970_),
    .Y(_2974_)
);

OR2X2 _9621_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2974_),
    .B(_2951_),
    .Y(_2975_)
);

NAND2X1 _9622_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2973_),
    .B(_2975_),
    .Y(_2976_)
);

AOI21X1 _9623_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2948_),
    .B(_2950_),
    .C(_2976_),
    .Y(_2977_)
);

NAND3X1 _9624_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2768_),
    .B(_2841_),
    .C(_2947_),
    .Y(_2978_)
);

OAI21X1 _9625_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2767_),
    .B(_2978_),
    .C(_2950_),
    .Y(_2979_)
);

INVX1 _9626_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2976_),
    .Y(_2980_)
);

NOR2X1 _9627_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2980_),
    .B(_2979_),
    .Y(_2981_)
);

NOR2X1 _9628_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2977_),
    .B(_2981_),
    .Y(_3187_[12])
);

NOR2X1 _9629_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2951_),
    .B(_2974_),
    .Y(_2982_)
);

INVX1 _9630_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2957_),
    .Y(_2983_)
);

OAI21X1 _9631_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2696_),
    .B(_2983_),
    .C(_2962_),
    .Y(_2984_)
);

INVX1 _9632_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2984_),
    .Y(_2985_)
);

NOR2X1 _9633_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2626_),
    .B(_2853_),
    .Y(_2986_)
);

NAND2X1 _9634_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2958_),
    .B(_2986_),
    .Y(_2987_)
);

OAI22X1 _9635_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2535_),
    .B(_2853_),
    .C(_2696_),
    .D(_2626_),
    .Y(_2988_)
);

NAND2X1 _9636_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2988_),
    .B(_2987_),
    .Y(_2989_)
);

NAND2X1 _9637_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2989_),
    .B(_2963_),
    .Y(_2990_)
);

OR2X2 _9638_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2963_),
    .B(_2989_),
    .Y(_2991_)
);

NAND2X1 _9639_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2990_),
    .B(_2991_),
    .Y(_2992_)
);

NAND2X1 _9640_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2985_),
    .B(_2992_),
    .Y(_2993_)
);

OR2X2 _9641_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2992_),
    .B(_2985_),
    .Y(_2994_)
);

NAND2X1 _9642_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2993_),
    .B(_2994_),
    .Y(_2995_)
);

NAND3X1 _9643_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2969_),
    .B(_2971_),
    .C(_2995_),
    .Y(_2996_)
);

OAI21X1 _9644_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2954_),
    .B(_2967_),
    .C(_2971_),
    .Y(_2997_)
);

AND2X2 _9645_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2994_),
    .B(_2993_),
    .Y(_2998_)
);

NAND2X1 _9646_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2997_),
    .B(_2998_),
    .Y(_2999_)
);

NAND2X1 _9647_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2996_),
    .B(_2999_),
    .Y(_3000_)
);

OAI21X1 _9648_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2982_),
    .B(_2977_),
    .C(_3000_),
    .Y(_3001_)
);

NAND2X1 _9649_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2980_),
    .B(_2979_),
    .Y(_3002_)
);

AND2X2 _9650_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2999_),
    .B(_2996_),
    .Y(_3003_)
);

NAND3X1 _9651_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2975_),
    .B(_3003_),
    .C(_3002_),
    .Y(_3004_)
);

NAND2X1 _9652_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3004_),
    .B(_3001_),
    .Y(_3187_[13])
);

NAND3X1 _9653_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2973_),
    .B(_2975_),
    .C(_3003_),
    .Y(_3005_)
);

AOI21X1 _9654_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2948_),
    .B(_2950_),
    .C(_3005_),
    .Y(_3006_)
);

OAI21X1 _9655_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2975_),
    .B(_3000_),
    .C(_2999_),
    .Y(_3007_)
);

OAI21X1 _9656_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2985_),
    .B(_2992_),
    .C(_2991_),
    .Y(_3008_)
);

AND2X2 _9657_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2987_),
    .B(_2986_),
    .Y(_3009_)
);

OR2X2 _9658_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3008_),
    .B(_3009_),
    .Y(_3010_)
);

NAND2X1 _9659_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3009_),
    .B(_3008_),
    .Y(_3011_)
);

NAND2X1 _9660_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3011_),
    .B(_3010_),
    .Y(_3012_)
);

OAI21X1 _9661_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3007_),
    .B(_3006_),
    .C(_3012_),
    .Y(_3013_)
);

INVX1 _9662_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2973_),
    .Y(_3014_)
);

NOR3X1 _9663_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3014_),
    .B(_2982_),
    .C(_3000_),
    .Y(_3015_)
);

NAND2X1 _9664_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3015_),
    .B(_2979_),
    .Y(_3016_)
);

INVX1 _9665_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3007_),
    .Y(_3017_)
);

INVX1 _9666_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3012_),
    .Y(_3018_)
);

NAND3X1 _9667_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3017_),
    .B(_3018_),
    .C(_3016_),
    .Y(_3019_)
);

NAND2X1 _9668_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3019_),
    .B(_3013_),
    .Y(_3187_[14])
);

OAI21X1 _9669_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3007_),
    .B(_3006_),
    .C(_3018_),
    .Y(_3020_)
);

OAI21X1 _9670_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2958_),
    .B(_3008_),
    .C(_2986_),
    .Y(_3021_)
);

NAND2X1 _9671_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3021_),
    .B(_3020_),
    .Y(_3187_[15])
);

INVX1 _9672_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_2415_),
    .Y(_3182_[0])
);

AND2X2 _9673_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [0]),
    .B(\u_fir_pe3.mul [0]),
    .Y(_3022_)
);

INVX1 _9674_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [1]),
    .Y(_3023_)
);

INVX1 _9675_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.mul [1]),
    .Y(_3024_)
);

NOR2X1 _9676_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3023_),
    .B(_3024_),
    .Y(_3025_)
);

NOR2X1 _9677_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [1]),
    .B(\u_fir_pe3.mul [1]),
    .Y(_3026_)
);

NOR2X1 _9678_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3026_),
    .B(_3025_),
    .Y(_3027_)
);

NAND2X1 _9679_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3022_),
    .B(_3027_),
    .Y(_3028_)
);

INVX1 _9680_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3028_),
    .Y(_3029_)
);

NOR2X1 _9681_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3022_),
    .B(_3027_),
    .Y(_3030_)
);

NOR2X1 _9682_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3030_),
    .B(_3029_),
    .Y(_3181_[1])
);

OAI21X1 _9683_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3023_),
    .B(_3024_),
    .C(_3028_),
    .Y(_3031_)
);

AND2X2 _9684_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [2]),
    .B(\u_fir_pe3.mul [2]),
    .Y(_3032_)
);

NOR2X1 _9685_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [2]),
    .B(\u_fir_pe3.mul [2]),
    .Y(_3033_)
);

OAI21X1 _9686_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3032_),
    .B(_3033_),
    .C(_3031_),
    .Y(_3034_)
);

INVX1 _9687_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3031_),
    .Y(_3035_)
);

NOR2X1 _9688_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3033_),
    .B(_3032_),
    .Y(_3036_)
);

NAND2X1 _9689_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3036_),
    .B(_3035_),
    .Y(_3037_)
);

NAND2X1 _9690_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3034_),
    .B(_3037_),
    .Y(_3181_[2])
);

AOI21X1 _9691_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3031_),
    .B(_3036_),
    .C(_3032_),
    .Y(_3038_)
);

INVX1 _9692_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [3]),
    .Y(_3039_)
);

INVX1 _9693_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.mul [3]),
    .Y(_3040_)
);

NOR2X1 _9694_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3039_),
    .B(_3040_),
    .Y(_3041_)
);

NOR2X1 _9695_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [3]),
    .B(\u_fir_pe3.mul [3]),
    .Y(_3042_)
);

NOR2X1 _9696_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3042_),
    .B(_3041_),
    .Y(_3043_)
);

NAND2X1 _9697_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3043_),
    .B(_3038_),
    .Y(_3044_)
);

OR2X2 _9698_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3038_),
    .B(_3043_),
    .Y(_3045_)
);

NAND2X1 _9699_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3044_),
    .B(_3045_),
    .Y(_3181_[3])
);

INVX1 _9700_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [4]),
    .Y(_3046_)
);

INVX1 _9701_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.mul [4]),
    .Y(_3047_)
);

NOR2X1 _9702_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3046_),
    .B(_3047_),
    .Y(_3048_)
);

NOR2X1 _9703_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [4]),
    .B(\u_fir_pe3.mul [4]),
    .Y(_3049_)
);

NOR2X1 _9704_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3049_),
    .B(_3048_),
    .Y(_3050_)
);

INVX1 _9705_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3041_),
    .Y(_3051_)
);

OAI21X1 _9706_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3042_),
    .B(_3038_),
    .C(_3051_),
    .Y(_3052_)
);

NAND2X1 _9707_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3050_),
    .B(_3052_),
    .Y(_3053_)
);

OR2X2 _9708_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3052_),
    .B(_3050_),
    .Y(_3054_)
);

AND2X2 _9709_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3054_),
    .B(_3053_),
    .Y(_3181_[4])
);

OAI21X1 _9710_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3046_),
    .B(_3047_),
    .C(_3053_),
    .Y(_3055_)
);

INVX1 _9711_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [5]),
    .Y(_3056_)
);

INVX1 _9712_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.mul [5]),
    .Y(_3057_)
);

NOR2X1 _9713_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3056_),
    .B(_3057_),
    .Y(_3058_)
);

NOR2X1 _9714_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [5]),
    .B(\u_fir_pe3.mul [5]),
    .Y(_3059_)
);

NOR2X1 _9715_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3059_),
    .B(_3058_),
    .Y(_3060_)
);

NAND2X1 _9716_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3060_),
    .B(_3055_),
    .Y(_3061_)
);

OR2X2 _9717_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3055_),
    .B(_3060_),
    .Y(_3062_)
);

AND2X2 _9718_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3062_),
    .B(_3061_),
    .Y(_3181_[5])
);

OAI21X1 _9719_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3056_),
    .B(_3057_),
    .C(_3061_),
    .Y(_3063_)
);

INVX1 _9720_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [6]),
    .Y(_3064_)
);

INVX1 _9721_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.mul [6]),
    .Y(_3065_)
);

NOR2X1 _9722_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3064_),
    .B(_3065_),
    .Y(_3066_)
);

NOR2X1 _9723_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [6]),
    .B(\u_fir_pe3.mul [6]),
    .Y(_3067_)
);

NOR2X1 _9724_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3067_),
    .B(_3066_),
    .Y(_3068_)
);

NAND2X1 _9725_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3068_),
    .B(_3063_),
    .Y(_3069_)
);

OR2X2 _9726_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3063_),
    .B(_3068_),
    .Y(_3070_)
);

AND2X2 _9727_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3070_),
    .B(_3069_),
    .Y(_3181_[6])
);

OAI21X1 _9728_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3064_),
    .B(_3065_),
    .C(_3069_),
    .Y(_3071_)
);

INVX1 _9729_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [7]),
    .Y(_3072_)
);

INVX1 _9730_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.mul [7]),
    .Y(_3073_)
);

NOR2X1 _9731_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3072_),
    .B(_3073_),
    .Y(_3074_)
);

NOR2X1 _9732_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [7]),
    .B(\u_fir_pe3.mul [7]),
    .Y(_3075_)
);

OAI21X1 _9733_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3074_),
    .B(_3075_),
    .C(_3071_),
    .Y(_3076_)
);

INVX1 _9734_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3071_),
    .Y(_3077_)
);

NOR2X1 _9735_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3075_),
    .B(_3074_),
    .Y(_3078_)
);

NAND2X1 _9736_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3078_),
    .B(_3077_),
    .Y(_3079_)
);

NAND2X1 _9737_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3076_),
    .B(_3079_),
    .Y(_3181_[7])
);

INVX1 _9738_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [8]),
    .Y(_3081_)
);

INVX1 _9739_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.mul [8]),
    .Y(_3082_)
);

NOR2X1 _9740_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3081_),
    .B(_3082_),
    .Y(_3083_)
);

NOR2X1 _9741_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [8]),
    .B(\u_fir_pe3.mul [8]),
    .Y(_3084_)
);

NAND2X1 _9742_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3048_),
    .B(_3060_),
    .Y(_3085_)
);

OAI21X1 _9743_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3056_),
    .B(_3057_),
    .C(_3085_),
    .Y(_3086_)
);

NAND2X1 _9744_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3066_),
    .B(_3078_),
    .Y(_3087_)
);

OAI21X1 _9745_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3072_),
    .B(_3073_),
    .C(_3087_),
    .Y(_3088_)
);

AND2X2 _9746_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3068_),
    .B(_3078_),
    .Y(_3089_)
);

AOI21X1 _9747_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3086_),
    .B(_3089_),
    .C(_3088_),
    .Y(_3090_)
);

AND2X2 _9748_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3050_),
    .B(_3060_),
    .Y(_3092_)
);

NAND3X1 _9749_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3092_),
    .B(_3089_),
    .C(_3052_),
    .Y(_3093_)
);

NAND2X1 _9750_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3090_),
    .B(_3093_),
    .Y(_3094_)
);

OAI21X1 _9751_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3083_),
    .B(_3084_),
    .C(_3094_),
    .Y(_3095_)
);

NOR2X1 _9752_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3084_),
    .B(_3083_),
    .Y(_3096_)
);

INVX1 _9753_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3094_),
    .Y(_3097_)
);

NAND2X1 _9754_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3096_),
    .B(_3097_),
    .Y(_3098_)
);

NAND2X1 _9755_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3095_),
    .B(_3098_),
    .Y(_3181_[8])
);

INVX1 _9756_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3083_),
    .Y(_3099_)
);

INVX1 _9757_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3096_),
    .Y(_3100_)
);

OAI21X1 _9758_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3100_),
    .B(_3097_),
    .C(_3099_),
    .Y(_3102_)
);

AND2X2 _9759_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [9]),
    .B(\u_fir_pe3.mul [9]),
    .Y(_3103_)
);

NOR2X1 _9760_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [9]),
    .B(\u_fir_pe3.mul [9]),
    .Y(_3104_)
);

NOR2X1 _9761_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3104_),
    .B(_3103_),
    .Y(_3105_)
);

INVX1 _9762_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3105_),
    .Y(_3106_)
);

OR2X2 _9763_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3102_),
    .B(_3106_),
    .Y(_3107_)
);

OAI21X1 _9764_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3103_),
    .B(_3104_),
    .C(_3102_),
    .Y(_3108_)
);

NAND2X1 _9765_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3108_),
    .B(_3107_),
    .Y(_3181_[9])
);

NOR2X1 _9766_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3106_),
    .B(_3100_),
    .Y(_3109_)
);

AOI21X1 _9767_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3105_),
    .B(_3083_),
    .C(_3103_),
    .Y(_3110_)
);

INVX1 _9768_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3110_),
    .Y(_3112_)
);

AOI21X1 _9769_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3094_),
    .B(_3109_),
    .C(_3112_),
    .Y(_3113_)
);

INVX1 _9770_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3113_),
    .Y(_3114_)
);

INVX1 _9771_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [10]),
    .Y(_3115_)
);

INVX1 _9772_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.mul [10]),
    .Y(_3116_)
);

NOR2X1 _9773_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3115_),
    .B(_3116_),
    .Y(_3117_)
);

NOR2X1 _9774_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [10]),
    .B(\u_fir_pe3.mul [10]),
    .Y(_3118_)
);

NOR2X1 _9775_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3118_),
    .B(_3117_),
    .Y(_3119_)
);

NAND2X1 _9776_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3119_),
    .B(_3114_),
    .Y(_3120_)
);

OAI21X1 _9777_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3117_),
    .B(_3118_),
    .C(_3113_),
    .Y(_3121_)
);

AND2X2 _9778_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3120_),
    .B(_3121_),
    .Y(_3181_[10])
);

OAI21X1 _9779_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3115_),
    .B(_3116_),
    .C(_3120_),
    .Y(_3123_)
);

AND2X2 _9780_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [11]),
    .B(\u_fir_pe3.mul [11]),
    .Y(_3124_)
);

NOR2X1 _9781_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [11]),
    .B(\u_fir_pe3.mul [11]),
    .Y(_3125_)
);

NOR2X1 _9782_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3125_),
    .B(_3124_),
    .Y(_3126_)
);

NOR2X1 _9783_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3126_),
    .B(_3123_),
    .Y(_3127_)
);

AND2X2 _9784_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3123_),
    .B(_3126_),
    .Y(_3128_)
);

NOR2X1 _9785_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3127_),
    .B(_3128_),
    .Y(_3181_[11])
);

AOI21X1 _9786_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3126_),
    .B(_3117_),
    .C(_3124_),
    .Y(_3129_)
);

NAND2X1 _9787_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3126_),
    .B(_3119_),
    .Y(_3130_)
);

OAI21X1 _9788_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3130_),
    .B(_3113_),
    .C(_3129_),
    .Y(_3132_)
);

INVX1 _9789_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [12]),
    .Y(_3133_)
);

INVX1 _9790_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.mul [12]),
    .Y(_3134_)
);

NOR2X1 _9791_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3133_),
    .B(_3134_),
    .Y(_3135_)
);

NOR2X1 _9792_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [12]),
    .B(\u_fir_pe3.mul [12]),
    .Y(_3136_)
);

NOR2X1 _9793_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3136_),
    .B(_3135_),
    .Y(_3137_)
);

NAND2X1 _9794_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3137_),
    .B(_3132_),
    .Y(_3138_)
);

OR2X2 _9795_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3132_),
    .B(_3137_),
    .Y(_3139_)
);

AND2X2 _9796_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3139_),
    .B(_3138_),
    .Y(_3181_[12])
);

OAI21X1 _9797_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3133_),
    .B(_3134_),
    .C(_3138_),
    .Y(_3140_)
);

INVX1 _9798_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [13]),
    .Y(_3142_)
);

INVX1 _9799_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.mul [13]),
    .Y(_3143_)
);

NOR2X1 _9800_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3142_),
    .B(_3143_),
    .Y(_3144_)
);

NOR2X1 _9801_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [13]),
    .B(\u_fir_pe3.mul [13]),
    .Y(_3145_)
);

NOR2X1 _9802_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3145_),
    .B(_3144_),
    .Y(_3146_)
);

NAND2X1 _9803_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3146_),
    .B(_3140_),
    .Y(_3147_)
);

OR2X2 _9804_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3140_),
    .B(_3146_),
    .Y(_3148_)
);

AND2X2 _9805_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3148_),
    .B(_3147_),
    .Y(_3181_[13])
);

OAI21X1 _9806_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3142_),
    .B(_3143_),
    .C(_3147_),
    .Y(_3149_)
);

INVX1 _9807_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [14]),
    .Y(_3150_)
);

INVX1 _9808_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.mul [14]),
    .Y(_3152_)
);

NOR2X1 _9809_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3150_),
    .B(_3152_),
    .Y(_3153_)
);

NOR2X1 _9810_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [14]),
    .B(\u_fir_pe3.mul [14]),
    .Y(_3154_)
);

NOR2X1 _9811_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3154_),
    .B(_3153_),
    .Y(_3155_)
);

AND2X2 _9812_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3149_),
    .B(_3155_),
    .Y(_3156_)
);

NOR2X1 _9813_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3155_),
    .B(_3149_),
    .Y(_3157_)
);

NOR2X1 _9814_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3157_),
    .B(_3156_),
    .Y(_3181_[14])
);

INVX1 _9815_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3153_),
    .Y(_3158_)
);

NAND2X1 _9816_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3155_),
    .B(_3149_),
    .Y(_3159_)
);

NAND2X1 _9817_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [15]),
    .B(\u_fir_pe3.mul [15]),
    .Y(_3160_)
);

OR2X2 _9818_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [15]),
    .B(\u_fir_pe3.mul [15]),
    .Y(_3162_)
);

NAND2X1 _9819_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3160_),
    .B(_3162_),
    .Y(_3163_)
);

INVX1 _9820_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3163_),
    .Y(_3164_)
);

NAND3X1 _9821_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3158_),
    .B(_3164_),
    .C(_3159_),
    .Y(_3165_)
);

OAI21X1 _9822_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3153_),
    .B(_3156_),
    .C(_3163_),
    .Y(_3166_)
);

NAND2X1 _9823_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3165_),
    .B(_3166_),
    .Y(_3181_[15])
);

NOR2X1 _9824_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_fir_pe3.rYin [0]),
    .B(\u_fir_pe3.mul [0]),
    .Y(_3167_)
);

NOR2X1 _9825_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3167_),
    .B(_3022_),
    .Y(_3180_[0])
);

AOI21X1 _9826_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[3] [0]),
    .B(vdd),
    .C(_3091_),
    .Y(_3168_)
);

NOR2X1 _9827_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3168_),
    .B(_3111_),
    .Y(_3183_[1])
);

NOR2X1 _9828_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3111_),
    .B(_3175_),
    .Y(_3170_)
);

NOR2X1 _9829_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3170_),
    .B(_3177_),
    .Y(_3184_[2])
);

DFFPOSX1 _9830_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf13),
    .D(_3180_[0]),
    .Q(\Y[4] [0])
);

DFFPOSX1 _9831_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf12),
    .D(_3181_[1]),
    .Q(\Y[4] [1])
);

DFFPOSX1 _9832_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf11),
    .D(_3181_[2]),
    .Q(\Y[4] [2])
);

DFFPOSX1 _9833_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf10),
    .D(_3181_[3]),
    .Q(\Y[4] [3])
);

DFFPOSX1 _9834_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf9),
    .D(_3181_[4]),
    .Q(\Y[4] [4])
);

DFFPOSX1 _9835_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf8),
    .D(_3181_[5]),
    .Q(\Y[4] [5])
);

DFFPOSX1 _9836_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf7),
    .D(_3181_[6]),
    .Q(\Y[4] [6])
);

DFFPOSX1 _9837_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_3181_[7]),
    .Q(\Y[4] [7])
);

DFFPOSX1 _9838_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_3181_[8]),
    .Q(\Y[4] [8])
);

DFFPOSX1 _9839_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_3181_[9]),
    .Q(\Y[4] [9])
);

DFFPOSX1 _9840_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_3181_[10]),
    .Q(\Y[4] [10])
);

DFFPOSX1 _9841_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_3181_[11]),
    .Q(\Y[4] [11])
);

DFFPOSX1 _9842_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_3181_[12]),
    .Q(\Y[4] [12])
);

DFFPOSX1 _9843_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_3181_[13]),
    .Q(\Y[4] [13])
);

DFFPOSX1 _9844_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf57),
    .D(_3181_[14]),
    .Q(\Y[4] [14])
);

DFFPOSX1 _9845_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf56),
    .D(_3181_[15]),
    .Q(\Y[4] [15])
);

DFFPOSX1 _9846_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf55),
    .D(\X[3] [0]),
    .Q(\X[4] [0])
);

DFFPOSX1 _9847_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf54),
    .D(\X[3] [1]),
    .Q(\X[4] [1])
);

DFFPOSX1 _9848_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf53),
    .D(\X[3] [2]),
    .Q(\X[4] [2])
);

DFFPOSX1 _9849_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf52),
    .D(\X[3] [3]),
    .Q(\X[4] [3])
);

DFFPOSX1 _9850_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf51),
    .D(\X[3] [4]),
    .Q(\X[4] [4])
);

DFFPOSX1 _9851_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf50),
    .D(\X[3]_5_bF$buf3 ),
    .Q(\X[4] [5])
);

DFFPOSX1 _9852_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf49),
    .D(\X[3] [6]),
    .Q(\X[4] [6])
);

DFFPOSX1 _9853_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf48),
    .D(\X[3] [7]),
    .Q(\X[4] [7])
);

DFFPOSX1 _9854_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf47),
    .D(\Y[3] [0]),
    .Q(\u_fir_pe3.rYin [0])
);

DFFPOSX1 _9855_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf46),
    .D(\Y[3] [1]),
    .Q(\u_fir_pe3.rYin [1])
);

DFFPOSX1 _9856_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf45),
    .D(\Y[3] [2]),
    .Q(\u_fir_pe3.rYin [2])
);

DFFPOSX1 _9857_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf44),
    .D(\Y[3] [3]),
    .Q(\u_fir_pe3.rYin [3])
);

DFFPOSX1 _9858_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf43),
    .D(\Y[3] [4]),
    .Q(\u_fir_pe3.rYin [4])
);

DFFPOSX1 _9859_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf42),
    .D(\Y[3] [5]),
    .Q(\u_fir_pe3.rYin [5])
);

DFFPOSX1 _9860_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf41),
    .D(\Y[3] [6]),
    .Q(\u_fir_pe3.rYin [6])
);

DFFPOSX1 _9861_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf40),
    .D(\Y[3] [7]),
    .Q(\u_fir_pe3.rYin [7])
);

DFFPOSX1 _9862_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf39),
    .D(\Y[3] [8]),
    .Q(\u_fir_pe3.rYin [8])
);

DFFPOSX1 _9863_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf38),
    .D(\Y[3] [9]),
    .Q(\u_fir_pe3.rYin [9])
);

DFFPOSX1 _9864_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf37),
    .D(\Y[3] [10]),
    .Q(\u_fir_pe3.rYin [10])
);

DFFPOSX1 _9865_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf36),
    .D(\Y[3] [11]),
    .Q(\u_fir_pe3.rYin [11])
);

DFFPOSX1 _9866_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf35),
    .D(\Y[3] [12]),
    .Q(\u_fir_pe3.rYin [12])
);

DFFPOSX1 _9867_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf34),
    .D(\Y[3] [13]),
    .Q(\u_fir_pe3.rYin [13])
);

DFFPOSX1 _9868_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf33),
    .D(\Y[3] [14]),
    .Q(\u_fir_pe3.rYin [14])
);

DFFPOSX1 _9869_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf32),
    .D(\Y[3] [15]),
    .Q(\u_fir_pe3.rYin [15])
);

DFFPOSX1 _9870_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf31),
    .D(_3182_[0]),
    .Q(\u_fir_pe3.mul [0])
);

DFFPOSX1 _9871_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf30),
    .D(_3183_[1]),
    .Q(\u_fir_pe3.mul [1])
);

DFFPOSX1 _9872_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf29),
    .D(_3184_[2]),
    .Q(\u_fir_pe3.mul [2])
);

DFFPOSX1 _9873_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf28),
    .D(_3185_[3]),
    .Q(\u_fir_pe3.mul [3])
);

DFFPOSX1 _9874_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf27),
    .D(_3186_[4]),
    .Q(\u_fir_pe3.mul [4])
);

DFFPOSX1 _9875_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf26),
    .D(_3187_[5]),
    .Q(\u_fir_pe3.mul [5])
);

DFFPOSX1 _9876_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf25),
    .D(_3187_[6]),
    .Q(\u_fir_pe3.mul [6])
);

DFFPOSX1 _9877_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf24),
    .D(_3187_[7]),
    .Q(\u_fir_pe3.mul [7])
);

DFFPOSX1 _9878_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf23),
    .D(_3187_[8]),
    .Q(\u_fir_pe3.mul [8])
);

DFFPOSX1 _9879_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf22),
    .D(_3187_[9]),
    .Q(\u_fir_pe3.mul [9])
);

DFFPOSX1 _9880_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf21),
    .D(_3187_[10]),
    .Q(\u_fir_pe3.mul [10])
);

DFFPOSX1 _9881_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf20),
    .D(_3187_[11]),
    .Q(\u_fir_pe3.mul [11])
);

DFFPOSX1 _9882_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf19),
    .D(_3187_[12]),
    .Q(\u_fir_pe3.mul [12])
);

DFFPOSX1 _9883_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf18),
    .D(_3187_[13]),
    .Q(\u_fir_pe3.mul [13])
);

DFFPOSX1 _9884_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf17),
    .D(_3187_[14]),
    .Q(\u_fir_pe3.mul [14])
);

DFFPOSX1 _9885_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf16),
    .D(_3187_[15]),
    .Q(\u_fir_pe3.mul [15])
);

NAND2X1 _9886_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [0]),
    .B(vdd),
    .Y(_3877_)
);

AND2X2 _9887_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [1]),
    .B(gnd),
    .Y(_3888_)
);

INVX1 _9888_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3888_),
    .Y(_3898_)
);

NOR2X1 _9889_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3877_),
    .B(_3898_),
    .Y(_3908_)
);

NAND2X1 _9890_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [1]),
    .Y(_3919_)
);

NOR2X1 _9891_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3877_),
    .B(_3919_),
    .Y(_3928_)
);

AOI22X1 _9892_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [0]),
    .B(gnd),
    .C(\X[4] [1]),
    .D(vdd),
    .Y(_3938_)
);

NOR2X1 _9893_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3938_),
    .B(_3928_),
    .Y(_3948_)
);

INVX1 _9894_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [2]),
    .Y(_3958_)
);

INVX2 _9895_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_3966_)
);

NOR2X1 _9896_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3958_),
    .B(_3966_),
    .Y(_3968_)
);

NAND2X1 _9897_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3968_),
    .B(_3948_),
    .Y(_3969_)
);

INVX1 _9898_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3969_),
    .Y(_3970_)
);

NOR2X1 _9899_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3968_),
    .B(_3948_),
    .Y(_3971_)
);

NOR2X1 _9900_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3971_),
    .B(_3970_),
    .Y(_3972_)
);

NAND2X1 _9901_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3908_),
    .B(_3972_),
    .Y(_3973_)
);

INVX1 _9902_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3973_),
    .Y(_3974_)
);

NAND2X1 _9903_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [3]),
    .Y(_3975_)
);

INVX1 _9904_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3975_),
    .Y(_3976_)
);

NAND2X1 _9905_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[4] [2]),
    .Y(_3188_)
);

INVX1 _9906_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3188_),
    .Y(_3189_)
);

NAND2X1 _9907_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [0]),
    .Y(_3190_)
);

OR2X2 _9908_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3919_),
    .B(_3190_),
    .Y(_3191_)
);

AOI22X1 _9909_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [0]),
    .C(gnd),
    .D(\X[4] [1]),
    .Y(_3192_)
);

INVX1 _9910_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3192_),
    .Y(_3193_)
);

NAND3X1 _9911_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3189_),
    .B(_3193_),
    .C(_3191_),
    .Y(_3194_)
);

NOR2X1 _9912_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3919_),
    .B(_3190_),
    .Y(_3195_)
);

OAI21X1 _9913_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3192_),
    .B(_3195_),
    .C(_3188_),
    .Y(_3196_)
);

NAND3X1 _9914_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3928_),
    .B(_3196_),
    .C(_3194_),
    .Y(_3197_)
);

INVX1 _9915_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3928_),
    .Y(_3198_)
);

NAND3X1 _9916_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3188_),
    .B(_3193_),
    .C(_3191_),
    .Y(_3199_)
);

OAI21X1 _9917_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3192_),
    .B(_3195_),
    .C(_3189_),
    .Y(_3200_)
);

NAND3X1 _9918_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3198_),
    .B(_3200_),
    .C(_3199_),
    .Y(_3201_)
);

NAND3X1 _9919_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3976_),
    .B(_3201_),
    .C(_3197_),
    .Y(_3202_)
);

INVX2 _9920_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [3]),
    .Y(_3203_)
);

NAND2X1 _9921_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3201_),
    .B(_3197_),
    .Y(_3204_)
);

OAI21X1 _9922_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3966_),
    .B(_3203_),
    .C(_3204_),
    .Y(_3205_)
);

NAND2X1 _9923_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3202_),
    .B(_3205_),
    .Y(_3206_)
);

NAND2X1 _9924_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3969_),
    .B(_3206_),
    .Y(_3207_)
);

NAND3X1 _9925_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3970_),
    .B(_3202_),
    .C(_3205_),
    .Y(_3208_)
);

NAND3X1 _9926_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3208_),
    .B(_3974_),
    .C(_3207_),
    .Y(_3209_)
);

INVX1 _9927_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3209_),
    .Y(_3210_)
);

AOI21X1 _9928_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3207_),
    .B(_3208_),
    .C(_3974_),
    .Y(_3211_)
);

NOR2X1 _9929_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3211_),
    .B(_3210_),
    .Y(_3982_[3])
);

NAND2X1 _9930_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [0]),
    .B(gnd),
    .Y(_3212_)
);

NAND2X1 _9931_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [4]),
    .B(gnd),
    .Y(_3213_)
);

NOR2X1 _9932_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3212_),
    .B(_3213_),
    .Y(_3214_)
);

AOI22X1 _9933_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [0]),
    .B(gnd),
    .C(gnd),
    .D(\X[4] [4]),
    .Y(_3215_)
);

NOR2X1 _9934_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3215_),
    .B(_3214_),
    .Y(_3216_)
);

INVX1 _9935_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3216_),
    .Y(_3217_)
);

NAND2X1 _9936_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [0]),
    .B(gnd),
    .Y(_3218_)
);

NAND2X1 _9937_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [1]),
    .Y(_3219_)
);

OAI22X1 _9938_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3218_),
    .B(_3219_),
    .C(_3188_),
    .D(_3192_),
    .Y(_3220_)
);

NAND2X1 _9939_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[4] [3]),
    .Y(_3221_)
);

INVX1 _9940_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3221_),
    .Y(_3222_)
);

AND2X2 _9941_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [1]),
    .Y(_3223_)
);

AND2X2 _9942_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [2]),
    .Y(_3224_)
);

NAND2X1 _9943_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3223_),
    .B(_3224_),
    .Y(_3225_)
);

AOI22X1 _9944_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [1]),
    .C(gnd),
    .D(\X[4] [2]),
    .Y(_3226_)
);

INVX1 _9945_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3226_),
    .Y(_3227_)
);

NAND3X1 _9946_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3222_),
    .B(_3227_),
    .C(_3225_),
    .Y(_3228_)
);

NAND3X1 _9947_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [2]),
    .C(_3219_),
    .Y(_3229_)
);

NAND2X1 _9948_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [2]),
    .Y(_3230_)
);

NAND3X1 _9949_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [1]),
    .C(_3230_),
    .Y(_3231_)
);

NAND3X1 _9950_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3221_),
    .B(_3229_),
    .C(_3231_),
    .Y(_3232_)
);

NAND3X1 _9951_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3220_),
    .B(_3232_),
    .C(_3228_),
    .Y(_3233_)
);

INVX1 _9952_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3220_),
    .Y(_3234_)
);

NAND2X1 _9953_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3232_),
    .B(_3228_),
    .Y(_3235_)
);

NAND2X1 _9954_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3234_),
    .B(_3235_),
    .Y(_3236_)
);

NAND3X1 _9955_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3217_),
    .B(_3233_),
    .C(_3236_),
    .Y(_3237_)
);

NAND2X1 _9956_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3220_),
    .B(_3235_),
    .Y(_3238_)
);

NAND3X1 _9957_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3228_),
    .B(_3232_),
    .C(_3234_),
    .Y(_3239_)
);

NAND3X1 _9958_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3216_),
    .B(_3239_),
    .C(_3238_),
    .Y(_3240_)
);

AOI22X1 _9959_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3197_),
    .B(_3202_),
    .C(_3237_),
    .D(_3240_),
    .Y(_3241_)
);

INVX1 _9960_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3241_),
    .Y(_3242_)
);

NAND2X1 _9961_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3197_),
    .B(_3202_),
    .Y(_3243_)
);

NAND2X1 _9962_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3237_),
    .B(_3240_),
    .Y(_3244_)
);

OR2X2 _9963_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3244_),
    .B(_3243_),
    .Y(_3245_)
);

NAND2X1 _9964_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3242_),
    .B(_3245_),
    .Y(_3246_)
);

OAI21X1 _9965_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3969_),
    .B(_3206_),
    .C(_3209_),
    .Y(_3247_)
);

OR2X2 _9966_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3247_),
    .B(_3246_),
    .Y(_3248_)
);

NAND3X1 _9967_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3216_),
    .B(_3233_),
    .C(_3236_),
    .Y(_3249_)
);

INVX1 _9968_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3233_),
    .Y(_3250_)
);

AOI21X1 _9969_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3228_),
    .B(_3232_),
    .C(_3220_),
    .Y(_3251_)
);

OAI21X1 _9970_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3251_),
    .B(_3250_),
    .C(_3217_),
    .Y(_3252_)
);

AOI21X1 _9971_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3249_),
    .B(_3252_),
    .C(_3243_),
    .Y(_3253_)
);

OAI21X1 _9972_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3241_),
    .B(_3253_),
    .C(_3247_),
    .Y(_3254_)
);

NAND2X1 _9973_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3254_),
    .B(_3248_),
    .Y(_3983_[4])
);

NOR2X1 _9974_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3209_),
    .B(_3246_),
    .Y(_3255_)
);

NOR3X1 _9975_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3241_),
    .B(_3208_),
    .C(_3253_),
    .Y(_3256_)
);

OAI21X1 _9976_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3217_),
    .B(_3251_),
    .C(_3233_),
    .Y(_3257_)
);

NAND2X1 _9977_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [0]),
    .B(vdd),
    .Y(_3258_)
);

INVX1 _9978_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3258_),
    .Y(_3259_)
);

AND2X2 _9979_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4]_5_bF$buf2 ),
    .Y(_3260_)
);

NAND2X1 _9980_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3888_),
    .B(_3260_),
    .Y(_3261_)
);

INVX2 _9981_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4]_5_bF$buf1 ),
    .Y(_3262_)
);

NAND2X1 _9982_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [1]),
    .B(gnd),
    .Y(_3263_)
);

OAI21X1 _9983_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3966_),
    .B(_3262_),
    .C(_3263_),
    .Y(_3264_)
);

NAND3X1 _9984_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3264_),
    .B(_3259_),
    .C(_3261_),
    .Y(_3265_)
);

NAND3X1 _9985_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4]_5_bF$buf0 ),
    .C(_3263_),
    .Y(_3266_)
);

NAND2X1 _9986_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4]_5_bF$buf3 ),
    .Y(_3267_)
);

NAND3X1 _9987_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\X[4] [1]),
    .B(gnd),
    .C(_3267_),
    .Y(_3268_)
);

NAND3X1 _9988_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3258_),
    .B(_3266_),
    .C(_3268_),
    .Y(_3269_)
);

AND2X2 _9989_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3265_),
    .B(_3269_),
    .Y(_3270_)
);

NAND2X1 _9990_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [2]),
    .Y(_3271_)
);

OAI22X1 _9991_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3919_),
    .B(_3271_),
    .C(_3221_),
    .D(_3226_),
    .Y(_3272_)
);

NAND2X1 _9992_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(vdd),
    .B(\X[4] [4]),
    .Y(_3273_)
);

INVX1 _9993_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3273_),
    .Y(_3274_)
);

AND2X2 _9994_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [3]),
    .Y(_3275_)
);

NAND2X1 _9995_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3224_),
    .B(_3275_),
    .Y(_3276_)
);

INVX1 _9996_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .Y(_3277_)
);

OAI21X1 _9997_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3277_),
    .B(_3203_),
    .C(_3271_),
    .Y(_3278_)
);

NAND3X1 _9998_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_3274_),
    .B(_3278_),
    .C(_3276_),
    .Y(_3279_)
);

NAND3X1 _9999_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(gnd),
    .B(\X[4] [3]),
    .C(_3271_),
    .Y(_3280_)
);

endmodule
