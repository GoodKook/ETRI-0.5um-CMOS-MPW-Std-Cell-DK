magic
tech scmos
magscale 1 30
timestamp 1749790639
<< checkpaint >>
rect 9150 9150 180850 180850
<< metal1 >>
rect 50175 144100 57900 144145
rect 50175 142800 51100 144100
rect 139300 142900 139305 144290
rect 46300 136560 46800 136600
rect 46100 135115 46600 136560
rect 50175 135255 51465 142800
rect 137925 135180 139305 142900
rect 46100 99700 46615 135115
rect 46600 90300 46615 99700
rect 46100 53500 46615 90300
rect 142665 98400 143190 127275
rect 142665 91600 142700 98400
rect 142665 67988 143190 91600
rect 50040 46800 51465 55140
rect 137925 47000 139215 54810
rect 142666 53529 143188 67988
rect 50040 45400 51100 46800
rect 139200 45655 139215 47000
rect 50040 45368 57900 45400
<< m2contact >>
rect 51100 142800 57900 144100
rect 130800 142900 139300 144300
rect 46000 90300 46600 99700
rect 142700 91600 143300 98400
rect 51100 45400 57900 46800
rect 130800 45600 139200 47000
<< metal2 >>
rect 51100 144100 57900 145800
rect 44200 136600 48100 139300
rect 73300 138000 73700 145900
rect 86800 138700 87200 145900
rect 100300 139400 100700 145900
rect 92300 137100 92700 137700
rect 93000 137100 93400 138400
rect 93700 137100 94100 139100
rect 113800 138700 114200 145900
rect 97800 137100 98200 138400
rect 127300 138000 127700 145900
rect 130800 144300 139300 145800
rect 140500 140800 145900 141200
rect 98500 137100 98900 137700
rect 47600 136300 48100 136600
rect 140100 135200 144600 135500
rect 44600 126700 47900 127100
rect 44600 125800 45000 126700
rect 44100 123100 45000 125800
rect 140730 125800 140940 127395
rect 140730 125400 143600 125800
rect 48700 112300 49100 125400
rect 140730 125395 140940 125400
rect 145000 116500 145900 116900
rect 44100 109600 49100 112300
rect 144000 103000 145900 103400
rect 44100 90300 46000 99700
rect 143300 91600 145900 98400
rect 44100 82600 47800 85300
rect 44100 69100 45800 71800
rect 45400 62400 45800 69100
rect 47400 63400 47800 82600
rect 140200 75990 145900 76400
rect 140200 64700 140500 75990
rect 143600 62500 145900 62900
rect 45400 62100 48300 62400
rect 44100 55600 45800 58300
rect 143600 55600 144000 62500
rect 45400 53200 45800 55600
rect 141050 55300 144000 55600
rect 144500 59800 145900 60200
rect 47900 53200 48300 53700
rect 141300 53500 141700 53800
rect 144500 53500 144900 59800
rect 45400 52800 48300 53200
rect 104500 51700 105000 53200
rect 51100 44200 57900 45400
rect 76000 44100 76400 51300
rect 105300 50900 105700 53200
rect 89500 44100 89900 50500
rect 106000 50000 106500 53200
rect 108900 52500 109400 53200
rect 141300 53100 144900 53500
rect 103000 44200 103400 49600
rect 116400 44100 116900 52100
rect 130800 44200 139200 45600
<< m3contact >>
rect 93700 139100 94100 139400
rect 100300 139100 100700 139400
rect 86800 138400 87200 138700
rect 93000 138400 93400 138700
rect 73300 137700 73700 138000
rect 92300 137700 92700 138000
rect 97800 138400 98200 138700
rect 113800 138400 114200 138700
rect 140100 140800 140500 141200
rect 98500 137700 98900 138000
rect 127300 137700 127700 138000
rect 140100 136500 140500 136900
rect 144600 135000 145000 135500
rect 143600 125300 144000 125800
rect 144600 116500 145000 117000
rect 143600 103000 144000 103500
rect 76000 51300 76400 51700
rect 104500 51300 105000 51700
rect 89500 50500 89900 50900
rect 105200 50500 105700 50900
rect 108900 52100 109400 52500
rect 116400 52100 116900 52500
rect 103000 49600 103500 50000
rect 106000 49600 106500 50000
<< metal3 >>
rect 94100 139100 100300 139400
rect 87200 138400 93000 138700
rect 98200 138400 113800 138700
rect 73700 137700 92300 138000
rect 98900 137700 127300 138000
rect 140100 136900 140500 140800
rect 143600 103500 144000 125300
rect 144600 117000 145000 135000
rect 109400 52100 116400 52500
rect 76400 51300 104500 51700
rect 89900 50500 105200 50900
rect 103500 49600 106000 50000
use PIC  clk ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 62000 0 -1 171100
box -100 -9150 12100 25300
use PIC  down
timestamp 1569139307
transform 1 0 102500 0 -1 171100
box -100 -9150 12100 25300
use PIC  enable
timestamp 1569139307
transform 1 0 75500 0 -1 171100
box -100 -9150 12100 25300
use PVSS  GND ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 62000 0 1 18900
box 0 -9150 12000 25300
use POB8  hsync ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 102500 0 1 18900
box -100 -9150 12100 25300
use PIC  INV_IN
timestamp 1569139307
transform 0 -1 171100 1 0 129500
box -100 -9150 12100 25300
use PANA  INV_INA ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 0 1 18900 -1 0 87500
box -100 -9150 12095 25300
use POB8  INV_OUT1
timestamp 1569139307
transform 0 -1 171100 1 0 116000
box -100 -9150 12100 25300
use PANA  INV_OUT1A
timestamp 1569139307
transform 0 1 18900 -1 0 74000
box -100 -9150 12095 25300
use POB8  INV_OUT8
timestamp 1569139307
transform 0 -1 171100 1 0 102500
box -100 -9150 12100 25300
use PANA  INV_OUT8A
timestamp 1569139307
transform 0 1 18900 -1 0 60500
box -100 -9150 12095 25300
use IOFILLER18  IOFILLER18_0 ~/ETRI050_DesignKit/pads_ETRI
timestamp 1725930584
transform 0 -1 171100 -1 0 75646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_1
timestamp 1725930584
transform 0 -1 171098 -1 0 62146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_2
timestamp 1725930584
transform 0 -1 171100 -1 0 102646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_3
timestamp 1725930584
transform 0 -1 171100 -1 0 89146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_4
timestamp 1725930584
transform 0 -1 171102 -1 0 129646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_5
timestamp 1725930584
transform 0 -1 171100 -1 0 116146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_6
timestamp 1725930584
transform 1 0 73845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_7
timestamp 1725930584
transform 1 0 60345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_8
timestamp 1725930584
transform 1 0 100845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_9
timestamp 1725930584
transform 1 0 87345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_10
timestamp 1725930584
transform 1 0 127845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_11
timestamp 1725930584
transform 1 0 114345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_12
timestamp 1725930584
transform 0 1 18899 -1 0 75655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_13
timestamp 1725930584
transform 0 1 18899 -1 0 62155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_14
timestamp 1725930584
transform 0 1 18900 -1 0 102655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_15
timestamp 1725930584
transform 0 1 18900 -1 0 89155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_16
timestamp 1725930584
transform 1 0 73845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_17
timestamp 1725930584
transform 0 1 18897 -1 0 116155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_18
timestamp 1725930584
transform 0 1 18900 -1 0 129655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_19
timestamp 1725930584
transform 1 0 60345 0 -1 171101
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_20
timestamp 1725930584
transform 1 0 100845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_21
timestamp 1725930584
transform 1 0 87344 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_22
timestamp 1725930584
transform 1 0 127845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_23
timestamp 1725930584
transform 1 0 114345 0 -1 171100
box -60 0 1860 25060
use IOFILLER50  IOFILLER50_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 43621 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_1
timestamp 1569139307
transform 1 0 141360 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_2
timestamp 1569139307
transform 1 0 141345 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_3
timestamp 1569139307
transform 1 0 43638 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_4
timestamp 1569139307
transform 0 1 18900 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_5
timestamp 1569139307
transform 0 1 18900 -1 0 146379
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_6
timestamp 1569139307
transform 0 -1 171100 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_7
timestamp 1569139307
transform 0 -1 171100 -1 0 146346
box -35 0 5035 25060
use PIC  NAND_IN
timestamp 1569139307
transform 0 -1 171100 1 0 48500
box -100 -9150 12100 25300
use PANA  NAND_OUT1A
timestamp 1569139307
transform 0 1 18900 -1 0 128000
box -100 -9150 12095 25300
use POB8  NAND_OUT1
timestamp 1569139307
transform 0 -1 171100 1 0 62000
box -100 -9150 12100 25300
use PANA  NAND_OUT8A
timestamp 1569139307
transform 0 1 18900 -1 0 114500
box -100 -9150 12095 25300
use POB8  NAND_OUT8
timestamp 1569139307
transform 0 -1 171100 1 0 75500
box -100 -9150 12100 25300
use POB8  p_tick
timestamp 1569139307
transform 1 0 116000 0 1 18900
box -100 -9150 12100 25300
use PANA  PANA_0
timestamp 1569139307
transform 0 1 18900 -1 0 141500
box -100 -9150 12095 25300
use PCORNER  PCORNER_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 18900 0 1 18900
box 0 0 25300 25300
use PCORNER  PCORNER_1
timestamp 1569139307
transform 1 0 18900 0 -1 171100
box 0 0 25300 25300
use PCORNER  PCORNER_2
timestamp 1569139307
transform 0 -1 171100 1 0 18900
box 0 0 25300 25300
use PCORNER  PCORNER_3
timestamp 1569139307
transform -1 0 171100 0 -1 171100
box 0 0 25300 25300
use pong_pt1_Core  pong_pt1_Core_0
timestamp 1749783318
transform 1 0 51495 0 1 53490
box -5295 -360 91695 83745
use PVDD  PVDD_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 48500 0 1 18900
box 0 -9150 12000 25300
use PVDD  PVDD_1
timestamp 1569139307
transform 0 -1 171100 1 0 89000
box 0 -9150 12000 25300
use PVSS  PVSS_0
timestamp 1569139307
transform 1 0 129500 0 1 18900
box 0 -9150 12000 25300
use PVSS  PVSS_1
timestamp 1569139307
transform 1 0 129500 0 -1 171100
box 0 -9150 12000 25300
use PVSS  PVSS_2
timestamp 1569139307
transform 0 1 18900 -1 0 101000
box 0 -9150 12000 25300
use PIC  reset
timestamp 1569139307
transform 1 0 89000 0 -1 171100
box -100 -9150 12100 25300
use POB8  rgb
timestamp 1569139307
transform 1 0 75500 0 1 18900
box -100 -9150 12100 25300
use PIC  up
timestamp 1569139307
transform 1 0 116000 0 -1 171100
box -100 -9150 12100 25300
use PVDD  VCC
timestamp 1569139307
transform 1 0 48500 0 -1 171100
box 0 -9150 12000 25300
use POB8  vsync
timestamp 1569139307
transform 1 0 89000 0 1 18900
box -100 -9150 12100 25300
<< end >>
