magic
tech scmos
magscale 1 3
timestamp 1554524574
<< checkpaint >>
rect -56 -56 84 254
<< genericcontact >>
rect 11 180 17 186
rect 11 152 17 158
rect 11 124 17 130
rect 11 96 17 102
rect 11 68 17 74
rect 11 40 17 46
rect 11 12 17 18
<< metal1 >>
rect 4 4 24 194
<< end >>
