magic
tech scmos
magscale 1 2
timestamp 1727735028
<< nwell >>
rect -12 134 112 252
rect 18 130 54 134
<< ntransistor >>
rect 20 14 24 34
rect 40 14 44 34
rect 60 14 64 54
<< ptransistor >>
rect 20 146 24 226
rect 30 146 34 226
rect 50 146 54 226
<< ndiffusion >>
rect 48 34 60 54
rect 18 14 20 34
rect 24 14 26 34
rect 38 14 40 34
rect 44 14 46 34
rect 58 14 60 34
rect 64 14 66 54
<< pdiffusion >>
rect 18 146 20 226
rect 24 146 30 226
rect 34 146 36 226
rect 48 146 50 226
rect 54 146 56 226
<< ndcontact >>
rect 6 14 18 34
rect 26 14 38 34
rect 46 14 58 34
rect 66 14 78 54
<< pdcontact >>
rect 6 146 18 226
rect 36 146 48 226
rect 56 146 68 226
<< psubstratepcontact >>
rect -6 -6 106 6
<< nsubstratencontact >>
rect -6 234 106 246
<< polysilicon >>
rect 20 226 24 230
rect 30 226 34 230
rect 50 226 54 230
rect 20 142 24 146
rect 12 137 24 142
rect 12 89 16 137
rect 30 109 34 146
rect 50 138 54 146
rect 12 46 16 77
rect 30 47 34 97
rect 55 62 64 74
rect 60 54 64 62
rect 12 41 24 46
rect 30 41 44 47
rect 20 34 24 41
rect 40 34 44 41
rect 20 10 24 14
rect 40 10 44 14
rect 60 10 64 14
<< polycontact >>
rect 42 126 54 138
rect 24 97 36 109
rect 4 77 16 89
rect 43 62 55 74
<< metal1 >>
rect -6 246 106 248
rect -6 232 106 234
rect 36 226 48 232
rect 68 146 72 156
rect 6 138 14 146
rect 48 138 54 139
rect 6 130 42 138
rect 23 83 37 97
rect 3 63 17 77
rect 48 74 54 126
rect 63 117 72 146
rect 63 103 77 117
rect 32 62 43 68
rect 32 34 38 62
rect 70 54 77 103
rect 6 8 14 14
rect 46 8 58 14
rect -6 6 106 8
rect -6 -8 106 -6
<< m1p >>
rect 63 103 77 117
rect 23 83 37 97
rect 3 63 17 77
<< labels >>
rlabel metal1 63 103 77 117 0 Y
port 2 nsew signal output
rlabel metal1 -6 -8 106 8 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 23 83 37 97 0 B
port 1 nsew signal input
rlabel metal1 -6 232 106 248 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 3 63 17 77 0 A
port 0 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
