magic
tech scmos
magscale 1 2
timestamp 1706263538
<< metal1 >>
rect 506 507 520 508
rect 726 507 739 508
rect 834 507 844 508
rect 889 507 901 508
rect 501 506 527 507
rect 540 506 575 507
rect 498 505 530 506
rect 496 504 530 505
rect 494 503 530 504
rect 492 502 530 503
rect 490 501 530 502
rect 489 500 530 501
rect 488 499 530 500
rect 486 498 530 499
rect 485 496 530 498
rect 484 495 530 496
rect 483 494 530 495
rect 482 492 530 494
rect 481 491 530 492
rect 480 490 510 491
rect 521 490 530 491
rect 480 489 507 490
rect 524 489 530 490
rect 479 488 505 489
rect 527 488 530 489
rect 479 487 503 488
rect 529 487 530 488
rect 540 505 581 506
rect 540 504 584 505
rect 540 503 586 504
rect 540 502 587 503
rect 540 501 589 502
rect 540 500 590 501
rect 540 498 591 500
rect 540 497 592 498
rect 540 495 593 497
rect 540 493 594 495
rect 478 486 502 487
rect 478 484 501 486
rect 477 483 500 484
rect 477 481 499 483
rect 477 479 498 481
rect 476 477 498 479
rect 476 470 497 477
rect 540 476 560 493
rect 568 492 594 493
rect 570 491 594 492
rect 572 489 595 491
rect 573 487 595 489
rect 574 482 595 487
rect 573 480 595 482
rect 573 479 594 480
rect 572 478 594 479
rect 571 477 594 478
rect 569 476 593 477
rect 540 475 593 476
rect 540 473 592 475
rect 540 472 591 473
rect 540 470 590 472
rect 602 470 623 507
rect 476 466 498 470
rect 540 469 589 470
rect 540 468 587 469
rect 540 467 586 468
rect 540 466 585 467
rect 476 465 499 466
rect 477 464 499 465
rect 540 465 583 466
rect 540 464 581 465
rect 477 463 500 464
rect 540 463 578 464
rect 603 463 623 470
rect 641 467 662 507
rect 721 506 743 507
rect 718 505 744 506
rect 716 504 744 505
rect 714 503 744 504
rect 713 502 744 503
rect 711 501 744 502
rect 710 500 744 501
rect 709 499 744 500
rect 762 499 800 507
rect 830 506 848 507
rect 883 506 905 507
rect 827 505 851 506
rect 880 505 907 506
rect 825 504 852 505
rect 878 504 909 505
rect 824 503 854 504
rect 875 503 911 504
rect 822 502 855 503
rect 874 502 912 503
rect 821 501 856 502
rect 874 501 913 502
rect 820 500 857 501
rect 874 500 914 501
rect 820 499 858 500
rect 708 498 744 499
rect 707 496 744 498
rect 706 495 744 496
rect 705 493 744 495
rect 704 492 729 493
rect 741 492 744 493
rect 703 491 726 492
rect 761 491 800 499
rect 819 498 858 499
rect 874 498 915 500
rect 818 497 859 498
rect 817 496 859 497
rect 874 496 916 498
rect 817 495 860 496
rect 816 494 860 495
rect 816 493 861 494
rect 815 492 836 493
rect 840 492 861 493
rect 874 492 917 496
rect 1650 493 1706 494
rect 1642 492 1709 493
rect 815 491 835 492
rect 841 491 862 492
rect 703 490 724 491
rect 702 489 723 490
rect 702 488 722 489
rect 702 487 721 488
rect 701 486 721 487
rect 701 485 720 486
rect 701 484 719 485
rect 700 482 719 484
rect 727 483 736 484
rect 761 483 777 491
rect 815 490 834 491
rect 814 488 834 490
rect 842 489 862 491
rect 843 488 862 489
rect 874 491 885 492
rect 894 491 917 492
rect 1636 491 1712 492
rect 874 490 881 491
rect 896 490 918 491
rect 1632 490 1714 491
rect 874 489 879 490
rect 874 488 877 489
rect 897 488 918 490
rect 1567 489 1571 490
rect 1627 489 1716 490
rect 1563 488 1577 489
rect 1623 488 1718 489
rect 814 486 833 488
rect 724 482 739 483
rect 760 482 777 483
rect 813 483 833 486
rect 843 485 863 488
rect 874 487 875 488
rect 700 479 718 482
rect 722 481 741 482
rect 760 481 787 482
rect 721 480 742 481
rect 760 480 791 481
rect 720 479 743 480
rect 760 479 793 480
rect 813 479 832 483
rect 699 478 718 479
rect 719 478 744 479
rect 760 478 795 479
rect 699 477 745 478
rect 760 477 796 478
rect 699 475 746 477
rect 760 475 798 477
rect 699 473 747 475
rect 760 474 799 475
rect 760 473 800 474
rect 699 470 748 473
rect 699 469 722 470
rect 727 469 748 470
rect 760 470 801 473
rect 699 468 721 469
rect 728 468 749 469
rect 699 467 720 468
rect 641 463 661 467
rect 477 461 501 463
rect 540 462 573 463
rect 478 460 502 461
rect 478 459 503 460
rect 529 459 530 460
rect 478 458 505 459
rect 527 458 530 459
rect 479 457 507 458
rect 524 457 530 458
rect 479 456 510 457
rect 520 456 530 457
rect 480 454 530 456
rect 481 452 530 454
rect 482 451 530 452
rect 483 450 530 451
rect 484 449 530 450
rect 485 448 530 449
rect 486 447 530 448
rect 487 446 530 447
rect 488 445 530 446
rect 489 444 530 445
rect 491 443 530 444
rect 493 442 530 443
rect 495 441 528 442
rect 499 440 524 441
rect 540 440 560 462
rect 603 460 624 463
rect 640 460 661 463
rect 699 463 719 467
rect 729 466 749 468
rect 760 468 802 470
rect 760 467 762 468
rect 777 467 802 468
rect 812 467 832 479
rect 780 466 803 467
rect 699 461 718 463
rect 603 459 625 460
rect 639 459 661 460
rect 604 458 626 459
rect 638 458 660 459
rect 604 457 627 458
rect 637 457 660 458
rect 700 457 719 461
rect 730 458 749 466
rect 781 465 803 466
rect 782 464 803 465
rect 783 459 803 464
rect 813 463 832 467
rect 844 481 863 485
rect 898 485 918 488
rect 1561 487 1581 488
rect 1619 487 1719 488
rect 1560 486 1584 487
rect 1614 486 1721 487
rect 1558 485 1589 486
rect 1608 485 1722 486
rect 898 483 917 485
rect 1557 484 1724 485
rect 1556 483 1726 484
rect 897 481 917 483
rect 1555 482 1727 483
rect 1555 481 1728 482
rect 844 467 864 481
rect 896 480 917 481
rect 1554 480 1730 481
rect 896 479 916 480
rect 895 478 916 479
rect 1553 479 1731 480
rect 1553 478 1733 479
rect 894 477 915 478
rect 1553 477 1734 478
rect 893 476 915 477
rect 1552 476 1735 477
rect 891 475 914 476
rect 890 474 914 475
rect 1552 475 1736 476
rect 1552 474 1646 475
rect 1664 474 1738 475
rect 889 473 913 474
rect 1552 473 1581 474
rect 1585 473 1643 474
rect 1669 473 1739 474
rect 888 472 912 473
rect 1552 472 1574 473
rect 1592 472 1642 473
rect 1672 472 1740 473
rect 886 471 911 472
rect 1553 471 1571 472
rect 1596 471 1642 472
rect 1676 471 1741 472
rect 885 470 910 471
rect 1553 470 1569 471
rect 1598 470 1644 471
rect 1681 470 1742 471
rect 884 469 909 470
rect 1554 469 1568 470
rect 1600 469 1649 470
rect 1685 469 1743 470
rect 883 468 907 469
rect 1555 468 1566 469
rect 1601 468 1652 469
rect 1690 468 1744 469
rect 882 467 906 468
rect 1532 467 1537 468
rect 1557 467 1562 468
rect 1603 467 1656 468
rect 1697 467 1745 468
rect 844 463 863 467
rect 880 466 905 467
rect 1529 466 1540 467
rect 1604 466 1659 467
rect 1707 466 1746 467
rect 879 465 903 466
rect 1527 465 1543 466
rect 1604 465 1662 466
rect 1713 465 1747 466
rect 878 464 901 465
rect 1525 464 1544 465
rect 1605 464 1665 465
rect 1717 464 1748 465
rect 813 459 833 463
rect 843 460 863 463
rect 877 463 900 464
rect 1524 463 1546 464
rect 1573 463 1581 464
rect 1606 463 1668 464
rect 1721 463 1749 464
rect 877 462 899 463
rect 1523 462 1547 463
rect 1569 462 1584 463
rect 1606 462 1671 463
rect 1725 462 1750 463
rect 876 461 897 462
rect 1522 461 1548 462
rect 1567 461 1586 462
rect 1606 461 1675 462
rect 1728 461 1751 462
rect 875 460 896 461
rect 1521 460 1549 461
rect 1565 460 1588 461
rect 1607 460 1679 461
rect 1732 460 1751 461
rect 843 459 862 460
rect 875 459 895 460
rect 1520 459 1550 460
rect 1563 459 1589 460
rect 1607 459 1685 460
rect 1735 459 1752 460
rect 783 458 802 459
rect 604 456 629 457
rect 635 456 660 457
rect 701 456 720 457
rect 729 456 748 458
rect 782 457 802 458
rect 605 453 659 456
rect 701 455 721 456
rect 728 455 748 456
rect 701 454 722 455
rect 727 454 748 455
rect 758 456 759 457
rect 781 456 802 457
rect 758 455 762 456
rect 780 455 802 456
rect 814 458 833 459
rect 814 456 834 458
rect 842 456 862 459
rect 874 458 894 459
rect 1519 458 1551 459
rect 1561 458 1590 459
rect 1607 458 1702 459
rect 1738 458 1753 459
rect 873 457 893 458
rect 1519 457 1553 458
rect 1559 457 1591 458
rect 1607 457 1707 458
rect 1740 457 1753 458
rect 873 456 892 457
rect 1518 456 1591 457
rect 1606 456 1711 457
rect 1743 456 1754 457
rect 814 455 835 456
rect 841 455 861 456
rect 873 455 918 456
rect 758 454 766 455
rect 777 454 802 455
rect 815 454 836 455
rect 840 454 861 455
rect 606 451 658 453
rect 702 452 747 454
rect 758 452 801 454
rect 815 453 860 454
rect 816 452 860 453
rect 607 450 657 451
rect 703 450 746 452
rect 758 450 800 452
rect 816 451 859 452
rect 872 451 918 455
rect 1517 454 1592 456
rect 1516 453 1592 454
rect 1606 455 1714 456
rect 1746 455 1754 456
rect 1606 454 1717 455
rect 1748 454 1754 455
rect 1606 453 1720 454
rect 1750 453 1755 454
rect 1515 451 1592 453
rect 1605 452 1723 453
rect 1752 452 1755 453
rect 1605 451 1726 452
rect 1754 451 1755 452
rect 817 450 859 451
rect 608 448 656 450
rect 704 449 745 450
rect 758 449 799 450
rect 817 449 858 450
rect 704 448 744 449
rect 609 447 655 448
rect 705 447 744 448
rect 758 447 798 449
rect 818 448 858 449
rect 818 447 857 448
rect 610 446 654 447
rect 706 446 743 447
rect 758 446 797 447
rect 819 446 856 447
rect 611 445 653 446
rect 707 445 742 446
rect 758 445 796 446
rect 820 445 855 446
rect 612 444 652 445
rect 708 444 741 445
rect 758 444 794 445
rect 821 444 854 445
rect 614 443 650 444
rect 709 443 739 444
rect 758 443 793 444
rect 822 443 853 444
rect 616 442 648 443
rect 711 442 738 443
rect 758 442 791 443
rect 824 442 851 443
rect 618 441 646 442
rect 713 441 736 442
rect 758 441 789 442
rect 826 441 850 442
rect 620 440 643 441
rect 715 440 733 441
rect 762 440 786 441
rect 828 440 847 441
rect 871 440 918 451
rect 1514 450 1592 451
rect 1513 449 1592 450
rect 1604 450 1729 451
rect 1604 449 1732 450
rect 1512 448 1592 449
rect 1603 448 1735 449
rect 1511 447 1591 448
rect 1510 446 1591 447
rect 1603 447 1737 448
rect 1603 446 1740 447
rect 1509 445 1590 446
rect 1604 445 1743 446
rect 1508 444 1590 445
rect 1606 444 1745 445
rect 1507 443 1589 444
rect 1608 443 1748 444
rect 1506 442 1588 443
rect 1609 442 1750 443
rect 1505 441 1587 442
rect 1611 441 1664 442
rect 1667 441 1753 442
rect 1504 440 1586 441
rect 1612 440 1664 441
rect 1671 440 1755 441
rect 504 439 518 440
rect 625 439 638 440
rect 719 439 729 440
rect 769 439 782 440
rect 832 439 843 440
rect 1503 439 1585 440
rect 1614 439 1664 440
rect 1673 439 1757 440
rect 1501 438 1583 439
rect 1615 438 1665 439
rect 1676 438 1760 439
rect 1500 437 1540 438
rect 1545 437 1582 438
rect 1617 437 1665 438
rect 1678 437 1761 438
rect 1498 436 1535 437
rect 1544 436 1581 437
rect 1618 436 1665 437
rect 1681 436 1762 437
rect 1497 435 1531 436
rect 1542 435 1580 436
rect 1619 435 1665 436
rect 1683 435 1764 436
rect 1495 434 1528 435
rect 1541 434 1579 435
rect 1621 434 1665 435
rect 1685 434 1764 435
rect 1494 433 1524 434
rect 1539 433 1578 434
rect 1622 433 1666 434
rect 1688 433 1765 434
rect 1492 432 1521 433
rect 1538 432 1577 433
rect 1623 432 1666 433
rect 1690 432 1766 433
rect 1490 431 1519 432
rect 1536 431 1576 432
rect 1624 431 1667 432
rect 1693 431 1767 432
rect 1489 430 1517 431
rect 1534 430 1576 431
rect 1625 430 1667 431
rect 1695 430 1767 431
rect 1487 429 1516 430
rect 1532 429 1575 430
rect 1626 429 1668 430
rect 1699 429 1768 430
rect 1485 428 1514 429
rect 1531 428 1575 429
rect 1627 428 1669 429
rect 1703 428 1768 429
rect 1483 427 1512 428
rect 1529 427 1574 428
rect 1481 426 1510 427
rect 1528 426 1574 427
rect 1590 427 1593 428
rect 1600 427 1603 428
rect 1628 427 1670 428
rect 1709 427 1769 428
rect 1590 426 1608 427
rect 1629 426 1671 427
rect 1713 426 1769 427
rect 1479 425 1509 426
rect 1476 424 1508 425
rect 1527 424 1574 426
rect 1591 425 1611 426
rect 1630 425 1672 426
rect 1716 425 1770 426
rect 1591 424 1612 425
rect 1631 424 1674 425
rect 1718 424 1770 425
rect 1474 423 1507 424
rect 1514 423 1516 424
rect 1526 423 1575 424
rect 1473 422 1507 423
rect 1509 422 1516 423
rect 1525 422 1575 423
rect 1471 421 1516 422
rect 1469 420 1516 421
rect 1524 420 1575 422
rect 1592 423 1614 424
rect 1632 423 1675 424
rect 1721 423 1771 424
rect 1592 422 1615 423
rect 1633 422 1677 423
rect 1723 422 1771 423
rect 1592 421 1616 422
rect 1633 421 1679 422
rect 1725 421 1771 422
rect 1468 419 1517 420
rect 1466 418 1517 419
rect 1523 419 1575 420
rect 1593 419 1617 421
rect 1634 420 1681 421
rect 1727 420 1772 421
rect 1635 419 1683 420
rect 1729 419 1772 420
rect 1523 418 1576 419
rect 1465 417 1517 418
rect 1464 416 1518 417
rect 1522 416 1576 418
rect 1463 415 1519 416
rect 1521 415 1576 416
rect 1594 418 1618 419
rect 1636 418 1685 419
rect 1731 418 1772 419
rect 1594 416 1619 418
rect 1636 417 1688 418
rect 1732 417 1772 418
rect 1637 416 1692 417
rect 1734 416 1773 417
rect 1594 415 1620 416
rect 1638 415 1695 416
rect 1736 415 1773 416
rect 1462 414 1577 415
rect 1461 413 1577 414
rect 1460 411 1577 413
rect 1459 409 1577 411
rect 1595 413 1621 415
rect 1638 414 1699 415
rect 1737 414 1773 415
rect 1639 413 1703 414
rect 1739 413 1773 414
rect 1595 411 1622 413
rect 1640 412 1708 413
rect 1740 412 1774 413
rect 1640 411 1712 412
rect 1742 411 1774 412
rect 1595 409 1623 411
rect 1641 410 1715 411
rect 1743 410 1774 411
rect 1641 409 1717 410
rect 1744 409 1774 410
rect 1459 407 1578 409
rect 1459 406 1479 407
rect 1480 406 1578 407
rect 500 403 507 404
rect 522 403 529 404
rect 543 403 550 404
rect 497 402 509 403
rect 520 402 531 403
rect 540 402 552 403
rect 569 402 575 404
rect 496 401 510 402
rect 519 401 532 402
rect 496 400 511 401
rect 496 399 501 400
rect 503 399 511 400
rect 518 400 532 401
rect 539 401 553 402
rect 539 400 554 401
rect 568 400 575 402
rect 518 399 524 400
rect 526 399 533 400
rect 496 398 498 399
rect 505 398 511 399
rect 517 398 523 399
rect 527 398 533 399
rect 539 399 544 400
rect 546 399 554 400
rect 567 399 575 400
rect 539 398 541 399
rect 548 398 554 399
rect 506 395 512 398
rect 517 397 522 398
rect 506 394 511 395
rect 505 393 511 394
rect 504 392 511 393
rect 516 394 522 397
rect 528 395 534 398
rect 503 391 510 392
rect 502 390 509 391
rect 501 389 508 390
rect 499 388 507 389
rect 516 388 521 394
rect 498 387 506 388
rect 497 386 504 387
rect 496 385 503 386
rect 516 385 522 388
rect 529 387 534 395
rect 549 395 555 398
rect 566 397 575 399
rect 565 396 575 397
rect 564 395 569 396
rect 549 394 554 395
rect 564 394 568 395
rect 548 393 554 394
rect 563 393 568 394
rect 547 392 554 393
rect 562 392 567 393
rect 546 391 553 392
rect 562 391 566 392
rect 545 390 552 391
rect 561 390 566 391
rect 544 389 551 390
rect 560 389 565 390
rect 542 388 550 389
rect 559 388 564 389
rect 570 388 575 396
rect 541 387 549 388
rect 558 387 564 388
rect 569 387 575 388
rect 496 384 502 385
rect 517 384 522 385
rect 528 384 534 387
rect 540 386 547 387
rect 539 385 546 386
rect 539 384 545 385
rect 495 383 501 384
rect 517 383 523 384
rect 527 383 533 384
rect 495 378 512 383
rect 517 382 524 383
rect 526 382 533 383
rect 538 383 544 384
rect 558 383 578 387
rect 607 385 613 404
rect 687 403 692 404
rect 711 403 716 404
rect 736 403 745 404
rect 687 402 691 403
rect 712 402 717 403
rect 733 402 747 403
rect 686 401 691 402
rect 685 399 690 401
rect 713 400 718 402
rect 731 401 747 402
rect 730 400 747 401
rect 684 397 689 399
rect 714 398 719 400
rect 729 399 747 400
rect 728 398 737 399
rect 745 398 747 399
rect 622 396 629 397
rect 619 395 631 396
rect 619 394 632 395
rect 639 394 644 397
rect 648 396 653 397
rect 646 395 654 396
rect 645 394 655 395
rect 683 394 688 397
rect 701 396 708 397
rect 715 396 720 398
rect 728 397 735 398
rect 699 395 709 396
rect 697 394 709 395
rect 619 393 633 394
rect 619 392 622 393
rect 628 392 633 393
rect 639 393 656 394
rect 683 393 687 394
rect 696 393 709 394
rect 639 392 647 393
rect 648 392 656 393
rect 619 391 620 392
rect 628 390 634 392
rect 623 389 634 390
rect 620 388 634 389
rect 619 387 634 388
rect 618 386 624 387
rect 617 385 623 386
rect 629 385 634 387
rect 606 384 612 385
rect 600 383 601 384
rect 605 383 612 384
rect 518 381 532 382
rect 519 380 531 381
rect 520 379 530 380
rect 522 378 528 379
rect 538 378 555 383
rect 570 378 575 383
rect 600 382 612 383
rect 617 383 622 385
rect 628 383 634 385
rect 617 382 623 383
rect 627 382 634 383
rect 581 381 587 382
rect 600 381 611 382
rect 617 381 634 382
rect 581 378 586 381
rect 600 380 610 381
rect 618 380 634 381
rect 600 379 609 380
rect 619 379 627 380
rect 600 378 607 379
rect 620 378 625 379
rect 629 378 634 380
rect 639 391 645 392
rect 639 378 644 391
rect 650 390 656 392
rect 651 378 656 390
rect 662 383 665 384
rect 661 382 666 383
rect 682 382 687 393
rect 695 392 704 393
rect 706 392 709 393
rect 716 395 720 396
rect 727 396 734 397
rect 759 396 766 397
rect 781 396 789 397
rect 804 396 809 397
rect 727 395 733 396
rect 756 395 768 396
rect 779 395 791 396
rect 802 395 811 396
rect 812 395 817 406
rect 695 390 701 392
rect 716 391 721 395
rect 694 384 700 390
rect 717 385 721 391
rect 726 394 733 395
rect 755 394 770 395
rect 778 394 792 395
rect 801 394 817 395
rect 726 388 732 394
rect 754 393 770 394
rect 777 393 793 394
rect 800 393 817 394
rect 738 388 749 393
rect 754 392 761 393
rect 764 392 771 393
rect 776 392 784 393
rect 786 392 794 393
rect 753 390 759 392
rect 765 391 772 392
rect 776 391 782 392
rect 788 391 794 392
rect 799 392 807 393
rect 809 392 817 393
rect 799 391 805 392
rect 753 389 758 390
rect 766 389 772 391
rect 726 386 733 388
rect 695 383 701 384
rect 695 382 703 383
rect 706 382 709 383
rect 660 380 667 382
rect 661 379 666 380
rect 683 379 688 382
rect 696 381 709 382
rect 697 380 709 381
rect 716 380 721 385
rect 727 385 734 386
rect 727 384 735 385
rect 728 383 736 384
rect 743 383 749 388
rect 752 386 758 389
rect 767 386 772 389
rect 753 385 758 386
rect 753 383 759 385
rect 766 384 772 386
rect 775 384 781 391
rect 789 385 795 391
rect 789 384 794 385
rect 798 384 804 391
rect 811 390 817 392
rect 812 386 817 390
rect 811 384 817 386
rect 765 383 771 384
rect 728 382 749 383
rect 729 381 749 382
rect 754 382 761 383
rect 764 382 771 383
rect 776 383 782 384
rect 788 383 794 384
rect 776 382 784 383
rect 786 382 794 383
rect 799 383 805 384
rect 810 383 817 384
rect 799 382 807 383
rect 809 382 817 383
rect 754 381 770 382
rect 777 381 793 382
rect 799 381 817 382
rect 731 380 749 381
rect 755 380 769 381
rect 778 380 792 381
rect 800 380 817 381
rect 698 379 709 380
rect 662 378 665 379
rect 581 377 585 378
rect 684 377 689 379
rect 700 378 708 379
rect 715 378 720 380
rect 732 379 747 380
rect 756 379 768 380
rect 779 379 791 380
rect 801 379 810 380
rect 735 378 744 379
rect 759 378 766 379
rect 781 378 789 379
rect 803 378 808 379
rect 812 378 817 380
rect 823 393 828 404
rect 836 403 843 404
rect 836 402 842 403
rect 835 401 842 402
rect 834 400 841 401
rect 834 399 840 400
rect 833 398 839 399
rect 832 397 839 398
rect 832 396 838 397
rect 852 396 859 397
rect 874 396 882 397
rect 831 395 837 396
rect 849 395 861 396
rect 872 395 884 396
rect 830 394 837 395
rect 848 394 863 395
rect 871 394 885 395
rect 830 393 836 394
rect 847 393 863 394
rect 870 393 886 394
rect 823 390 835 393
rect 847 392 854 393
rect 857 392 864 393
rect 869 392 877 393
rect 879 392 887 393
rect 846 390 852 392
rect 858 391 865 392
rect 869 391 875 392
rect 881 391 887 392
rect 823 378 828 390
rect 829 389 836 390
rect 846 389 851 390
rect 859 389 865 391
rect 830 388 837 389
rect 831 387 837 388
rect 831 386 838 387
rect 845 386 851 389
rect 860 386 865 389
rect 832 385 839 386
rect 846 385 851 386
rect 833 383 840 385
rect 846 383 852 385
rect 859 384 865 386
rect 868 384 874 391
rect 882 385 888 391
rect 892 389 898 406
rect 1459 405 1477 406
rect 1479 405 1578 406
rect 1460 404 1475 405
rect 1478 404 1578 405
rect 1460 403 1473 404
rect 1477 403 1578 404
rect 1461 402 1470 403
rect 1476 402 1578 403
rect 1463 401 1466 402
rect 1475 401 1578 402
rect 1474 400 1578 401
rect 1473 399 1578 400
rect 1595 407 1624 409
rect 1642 408 1719 409
rect 1746 408 1774 409
rect 1642 407 1721 408
rect 1747 407 1774 408
rect 1595 404 1625 407
rect 1643 406 1722 407
rect 1748 406 1774 407
rect 1643 405 1724 406
rect 1749 405 1775 406
rect 1643 404 1726 405
rect 1751 404 1775 405
rect 1595 402 1626 404
rect 1644 403 1727 404
rect 1752 403 1775 404
rect 1644 402 1729 403
rect 1753 402 1775 403
rect 1595 400 1627 402
rect 1645 401 1730 402
rect 1754 401 1775 402
rect 1645 400 1731 401
rect 1755 400 1775 401
rect 1472 398 1577 399
rect 1595 398 1628 400
rect 1646 399 1733 400
rect 1756 399 1775 400
rect 1647 398 1734 399
rect 1757 398 1775 399
rect 1471 397 1577 398
rect 903 396 910 397
rect 1470 396 1577 397
rect 903 395 909 396
rect 1469 395 1577 396
rect 1594 396 1629 398
rect 1647 397 1735 398
rect 1758 397 1775 398
rect 1648 396 1737 397
rect 1759 396 1775 397
rect 902 394 908 395
rect 901 393 908 394
rect 1468 393 1576 395
rect 1594 394 1630 396
rect 1649 395 1738 396
rect 1760 395 1775 396
rect 1650 394 1739 395
rect 1594 393 1631 394
rect 1651 393 1740 394
rect 1761 393 1775 395
rect 901 392 907 393
rect 1467 392 1576 393
rect 900 391 906 392
rect 899 389 905 391
rect 1467 390 1575 392
rect 1593 391 1632 393
rect 1652 392 1742 393
rect 1762 392 1775 393
rect 1654 391 1743 392
rect 1763 391 1775 392
rect 1593 390 1633 391
rect 1656 390 1744 391
rect 1466 389 1574 390
rect 892 387 904 389
rect 1467 388 1574 389
rect 1592 388 1634 390
rect 1658 389 1745 390
rect 1764 389 1774 391
rect 1660 388 1746 389
rect 1765 388 1774 389
rect 1467 387 1573 388
rect 1592 387 1635 388
rect 1664 387 1747 388
rect 892 386 905 387
rect 1467 386 1572 387
rect 1592 386 1636 387
rect 1669 386 1748 387
rect 1766 386 1774 388
rect 882 384 887 385
rect 858 383 864 384
rect 834 382 841 383
rect 847 382 854 383
rect 857 382 864 383
rect 869 383 875 384
rect 881 383 887 384
rect 869 382 877 383
rect 879 382 887 383
rect 835 380 842 382
rect 847 381 863 382
rect 870 381 886 382
rect 848 380 862 381
rect 871 380 885 381
rect 836 379 843 380
rect 849 379 861 380
rect 872 379 884 380
rect 837 378 844 379
rect 852 378 859 379
rect 874 378 882 379
rect 892 378 898 386
rect 899 385 905 386
rect 1468 385 1572 386
rect 1591 385 1637 386
rect 1675 385 1749 386
rect 1767 385 1774 386
rect 900 384 906 385
rect 1468 384 1571 385
rect 1591 384 1639 385
rect 1681 384 1750 385
rect 900 383 907 384
rect 901 382 908 383
rect 1469 382 1570 384
rect 1590 383 1640 384
rect 1686 383 1751 384
rect 1768 383 1773 385
rect 1590 382 1642 383
rect 1689 382 1752 383
rect 1769 382 1773 383
rect 902 381 908 382
rect 1470 381 1569 382
rect 1590 381 1643 382
rect 1692 381 1753 382
rect 1769 381 1772 382
rect 902 380 909 381
rect 1470 380 1515 381
rect 1517 380 1568 381
rect 903 379 910 380
rect 1471 379 1513 380
rect 1519 379 1568 380
rect 1589 380 1645 381
rect 1695 380 1753 381
rect 1770 380 1772 381
rect 1589 379 1648 380
rect 1698 379 1754 380
rect 1770 379 1771 380
rect 904 378 910 379
rect 1472 378 1512 379
rect 1520 378 1567 379
rect 1588 378 1651 379
rect 1700 378 1755 379
rect 580 375 585 377
rect 685 376 689 377
rect 714 376 719 378
rect 1473 377 1511 378
rect 1521 377 1566 378
rect 1588 377 1655 378
rect 1703 377 1755 378
rect 1474 376 1510 377
rect 1521 376 1565 377
rect 1588 376 1660 377
rect 1705 376 1755 377
rect 685 375 690 376
rect 580 373 584 375
rect 686 373 691 375
rect 713 374 718 376
rect 1475 375 1509 376
rect 1522 375 1565 376
rect 1587 375 1665 376
rect 1708 375 1756 376
rect 1476 374 1506 375
rect 1522 374 1564 375
rect 1587 374 1671 375
rect 1711 374 1756 375
rect 712 373 717 374
rect 1477 373 1502 374
rect 1521 373 1564 374
rect 1586 373 1675 374
rect 1713 373 1756 374
rect 687 372 692 373
rect 711 372 716 373
rect 1479 372 1494 373
rect 1521 372 1563 373
rect 1586 372 1679 373
rect 1715 372 1757 373
rect 1484 371 1485 372
rect 1519 371 1562 372
rect 1516 370 1562 371
rect 1585 371 1681 372
rect 1716 371 1757 372
rect 1585 370 1684 371
rect 1718 370 1757 371
rect 1513 369 1561 370
rect 1584 369 1687 370
rect 1719 369 1757 370
rect 1509 368 1561 369
rect 1583 368 1689 369
rect 1720 368 1757 369
rect 1503 367 1560 368
rect 1583 367 1691 368
rect 1721 367 1758 368
rect 1494 366 1559 367
rect 1484 365 1559 366
rect 1582 366 1693 367
rect 1722 366 1758 367
rect 1582 365 1695 366
rect 1723 365 1758 366
rect 1482 364 1558 365
rect 1581 364 1697 365
rect 1724 364 1758 365
rect 1482 363 1557 364
rect 1481 362 1557 363
rect 1580 363 1699 364
rect 1725 363 1758 364
rect 1580 362 1700 363
rect 1726 362 1758 363
rect 1481 361 1556 362
rect 1579 361 1702 362
rect 1481 360 1555 361
rect 1578 360 1703 361
rect 1727 360 1758 362
rect 1481 359 1554 360
rect 1577 359 1704 360
rect 1728 359 1758 360
rect 1481 358 1553 359
rect 1577 358 1705 359
rect 1729 358 1758 359
rect 1481 357 1552 358
rect 1576 357 1706 358
rect 1482 356 1551 357
rect 1575 356 1707 357
rect 1730 356 1758 358
rect 1482 355 1550 356
rect 1574 355 1708 356
rect 1482 354 1549 355
rect 1573 354 1709 355
rect 1731 354 1758 356
rect 1483 353 1548 354
rect 1572 353 1710 354
rect 1732 353 1758 354
rect 471 352 692 353
rect 732 352 958 353
rect 994 352 1202 353
rect 1283 352 1350 353
rect 1483 352 1546 353
rect 1572 352 1711 353
rect 470 317 693 352
rect 732 351 959 352
rect 993 351 1208 352
rect 1283 351 1351 352
rect 731 317 960 351
rect 993 350 1211 351
rect 992 349 1213 350
rect 993 348 1215 349
rect 993 347 1217 348
rect 993 346 1218 347
rect 993 345 1220 346
rect 993 344 1221 345
rect 993 343 1222 344
rect 993 342 1223 343
rect 993 341 1224 342
rect 993 339 1225 341
rect 993 338 1226 339
rect 993 336 1227 338
rect 993 334 1228 336
rect 993 332 1229 334
rect 993 329 1230 332
rect 993 323 1231 329
rect 470 316 692 317
rect 732 316 959 317
rect 993 316 1232 323
rect 470 315 540 316
rect 811 315 881 316
rect 470 287 539 315
rect 470 286 540 287
rect 470 285 691 286
rect 470 284 692 285
rect 470 250 693 284
rect 470 249 692 250
rect 470 248 541 249
rect 543 248 545 249
rect 689 248 690 249
rect 470 247 540 248
rect 470 219 539 247
rect 470 218 540 219
rect 470 217 692 218
rect 470 209 693 217
rect 471 205 693 209
rect 472 202 693 205
rect 473 200 693 202
rect 474 198 693 200
rect 475 196 693 198
rect 476 195 693 196
rect 477 194 693 195
rect 478 192 693 194
rect 479 191 693 192
rect 480 190 693 191
rect 481 189 693 190
rect 482 188 693 189
rect 484 187 693 188
rect 485 186 693 187
rect 487 185 693 186
rect 489 184 693 185
rect 492 183 693 184
rect 494 182 693 183
rect 811 182 880 315
rect 993 185 1062 316
rect 1163 262 1232 316
rect 1085 261 1087 262
rect 1089 261 1159 262
rect 1160 261 1231 262
rect 1084 260 1166 261
rect 1085 259 1166 260
rect 1086 258 1166 259
rect 1087 257 1168 258
rect 1088 256 1169 257
rect 1089 255 1170 256
rect 1090 254 1170 255
rect 1091 253 1172 254
rect 1092 252 1173 253
rect 1093 251 1174 252
rect 1094 250 1175 251
rect 1095 249 1176 250
rect 1096 248 1177 249
rect 1097 247 1178 248
rect 1098 246 1179 247
rect 1099 245 1180 246
rect 1100 244 1181 245
rect 1101 243 1182 244
rect 1102 242 1183 243
rect 1103 241 1184 242
rect 1104 240 1185 241
rect 1105 239 1186 240
rect 1106 238 1187 239
rect 1107 237 1188 238
rect 1108 236 1189 237
rect 1109 235 1190 236
rect 1110 234 1191 235
rect 1111 233 1192 234
rect 1112 232 1193 233
rect 1113 231 1194 232
rect 1114 230 1195 231
rect 1115 229 1196 230
rect 1116 228 1197 229
rect 1117 227 1198 228
rect 1118 226 1199 227
rect 1119 225 1200 226
rect 1120 224 1201 225
rect 1121 223 1202 224
rect 1122 222 1203 223
rect 1123 221 1204 222
rect 1124 220 1205 221
rect 1125 219 1206 220
rect 1126 218 1207 219
rect 1127 217 1208 218
rect 1128 216 1209 217
rect 1129 215 1210 216
rect 1130 214 1211 215
rect 1131 213 1212 214
rect 1132 212 1213 213
rect 1133 211 1214 212
rect 1134 210 1215 211
rect 1135 209 1216 210
rect 1136 208 1217 209
rect 1137 207 1218 208
rect 1138 206 1219 207
rect 1139 205 1220 206
rect 1140 204 1221 205
rect 1141 203 1223 204
rect 1142 202 1223 203
rect 1143 201 1225 202
rect 1144 200 1225 201
rect 1145 199 1227 200
rect 1146 198 1227 199
rect 1147 197 1229 198
rect 1148 196 1229 197
rect 1149 195 1231 196
rect 1150 194 1231 195
rect 1151 193 1233 194
rect 1152 192 1233 193
rect 1153 191 1235 192
rect 1154 190 1235 191
rect 1155 189 1237 190
rect 1156 188 1237 189
rect 1157 187 1239 188
rect 1158 186 1239 187
rect 1159 185 1241 186
rect 992 183 1062 185
rect 1160 184 1241 185
rect 1161 183 1243 184
rect 1282 183 1351 351
rect 1484 351 1545 352
rect 1571 351 1631 352
rect 1640 351 1711 352
rect 1733 351 1758 353
rect 1484 350 1543 351
rect 1570 350 1629 351
rect 1644 350 1712 351
rect 1485 349 1541 350
rect 1568 349 1628 350
rect 1646 349 1713 350
rect 1734 349 1758 351
rect 1486 348 1539 349
rect 1567 348 1627 349
rect 1648 348 1713 349
rect 1486 347 1537 348
rect 1566 347 1626 348
rect 1650 347 1714 348
rect 1735 347 1758 349
rect 1487 346 1535 347
rect 1565 346 1625 347
rect 1651 346 1714 347
rect 1736 346 1758 347
rect 1488 345 1533 346
rect 1564 345 1625 346
rect 1653 345 1715 346
rect 1736 345 1757 346
rect 1488 344 1530 345
rect 1562 344 1624 345
rect 1654 344 1715 345
rect 1489 343 1527 344
rect 1561 343 1624 344
rect 1655 343 1716 344
rect 1737 343 1757 345
rect 1489 342 1524 343
rect 1560 342 1623 343
rect 1656 342 1716 343
rect 1490 341 1522 342
rect 1558 341 1623 342
rect 1657 341 1716 342
rect 1490 340 1518 341
rect 1556 340 1623 341
rect 1658 340 1717 341
rect 1738 340 1757 343
rect 1490 339 1515 340
rect 1555 339 1622 340
rect 1659 339 1717 340
rect 1491 338 1512 339
rect 1553 338 1622 339
rect 1660 338 1717 339
rect 1739 338 1756 340
rect 1491 337 1509 338
rect 1551 337 1622 338
rect 1661 337 1717 338
rect 1492 336 1506 337
rect 1549 336 1621 337
rect 1662 336 1717 337
rect 1492 335 1503 336
rect 1547 335 1621 336
rect 1663 335 1717 336
rect 1740 336 1756 338
rect 1740 335 1755 336
rect 1493 334 1500 335
rect 1545 334 1621 335
rect 1638 334 1640 335
rect 1663 334 1718 335
rect 1543 333 1620 334
rect 1638 333 1641 334
rect 1540 332 1620 333
rect 1538 331 1620 332
rect 1637 332 1642 333
rect 1664 332 1718 334
rect 1741 333 1755 335
rect 1741 332 1754 333
rect 1536 330 1619 331
rect 1637 330 1643 332
rect 1665 330 1717 332
rect 1533 329 1619 330
rect 1636 329 1644 330
rect 1531 328 1618 329
rect 1636 328 1645 329
rect 1666 328 1717 330
rect 1742 330 1754 332
rect 1742 329 1753 330
rect 1529 327 1618 328
rect 1635 327 1645 328
rect 1526 326 1617 327
rect 1635 326 1646 327
rect 1667 326 1717 328
rect 1743 328 1753 329
rect 1743 326 1752 328
rect 1524 325 1617 326
rect 1522 324 1616 325
rect 1634 324 1647 326
rect 1520 323 1616 324
rect 1518 322 1615 323
rect 1633 322 1648 324
rect 1668 323 1716 326
rect 1744 324 1751 326
rect 1516 321 1615 322
rect 1632 321 1649 322
rect 1669 321 1715 323
rect 1744 322 1750 324
rect 1745 321 1749 322
rect 1515 320 1614 321
rect 1632 320 1650 321
rect 1513 319 1614 320
rect 1512 318 1613 319
rect 1631 318 1650 320
rect 1669 319 1714 321
rect 1745 320 1748 321
rect 1745 319 1747 320
rect 1670 318 1713 319
rect 1745 318 1746 319
rect 1510 317 1613 318
rect 1509 316 1612 317
rect 1630 316 1651 318
rect 1670 316 1712 318
rect 1508 315 1611 316
rect 1507 314 1611 315
rect 1629 314 1652 316
rect 1670 315 1711 316
rect 1506 313 1610 314
rect 1628 313 1652 314
rect 1671 314 1710 315
rect 1505 312 1609 313
rect 1504 311 1608 312
rect 1628 311 1653 313
rect 1671 312 1709 314
rect 1671 311 1708 312
rect 1503 310 1607 311
rect 1502 309 1607 310
rect 1627 310 1653 311
rect 1672 310 1707 311
rect 1627 309 1654 310
rect 1502 308 1606 309
rect 1501 307 1605 308
rect 1626 307 1654 309
rect 1500 306 1604 307
rect 1625 306 1654 307
rect 1672 309 1706 310
rect 1672 308 1705 309
rect 1672 307 1704 308
rect 1672 306 1703 307
rect 1730 306 1731 307
rect 1500 305 1603 306
rect 1625 305 1655 306
rect 1499 304 1602 305
rect 1624 304 1655 305
rect 1672 305 1702 306
rect 1729 305 1731 306
rect 1672 304 1700 305
rect 1728 304 1731 305
rect 1499 303 1601 304
rect 1498 302 1600 303
rect 1623 302 1655 304
rect 1498 301 1599 302
rect 1622 301 1655 302
rect 1673 303 1699 304
rect 1727 303 1732 304
rect 1673 302 1698 303
rect 1726 302 1732 303
rect 1673 301 1696 302
rect 1725 301 1732 302
rect 1497 300 1598 301
rect 1497 299 1597 300
rect 1621 299 1656 301
rect 1496 298 1596 299
rect 1620 298 1656 299
rect 1496 297 1595 298
rect 1619 297 1656 298
rect 1495 296 1594 297
rect 1495 295 1593 296
rect 1618 295 1656 297
rect 1673 300 1695 301
rect 1724 300 1732 301
rect 1673 299 1693 300
rect 1723 299 1732 300
rect 1673 298 1692 299
rect 1722 298 1732 299
rect 1673 297 1690 298
rect 1721 297 1732 298
rect 1673 296 1688 297
rect 1720 296 1733 297
rect 1673 295 1687 296
rect 1719 295 1733 296
rect 1495 294 1591 295
rect 1617 294 1656 295
rect 1495 293 1590 294
rect 1616 293 1656 294
rect 1494 292 1589 293
rect 1615 292 1656 293
rect 1494 291 1587 292
rect 1614 291 1656 292
rect 1494 290 1586 291
rect 1613 290 1656 291
rect 1494 289 1584 290
rect 1612 289 1656 290
rect 1672 294 1685 295
rect 1718 294 1733 295
rect 1672 293 1683 294
rect 1716 293 1733 294
rect 1672 292 1681 293
rect 1715 292 1733 293
rect 1672 291 1678 292
rect 1714 291 1733 292
rect 1672 290 1676 291
rect 1713 290 1733 291
rect 1672 289 1673 290
rect 1711 289 1733 290
rect 1494 288 1583 289
rect 1611 288 1656 289
rect 1710 288 1733 289
rect 1493 287 1581 288
rect 1610 287 1656 288
rect 1708 287 1733 288
rect 1493 286 1579 287
rect 1608 286 1656 287
rect 1707 286 1733 287
rect 1493 285 1577 286
rect 1607 285 1656 286
rect 1705 285 1733 286
rect 1493 284 1575 285
rect 1606 284 1656 285
rect 1704 284 1733 285
rect 1493 283 1574 284
rect 1605 283 1656 284
rect 1702 283 1733 284
rect 1493 282 1571 283
rect 1603 282 1656 283
rect 1701 282 1733 283
rect 1493 281 1569 282
rect 1602 281 1655 282
rect 1699 281 1733 282
rect 1493 280 1567 281
rect 1600 280 1655 281
rect 1697 280 1733 281
rect 1493 279 1565 280
rect 1599 279 1655 280
rect 1695 279 1733 280
rect 1493 278 1563 279
rect 1597 278 1655 279
rect 1694 278 1733 279
rect 1493 277 1560 278
rect 1595 277 1655 278
rect 1692 277 1733 278
rect 1493 276 1558 277
rect 1594 276 1655 277
rect 1690 276 1732 277
rect 1493 275 1556 276
rect 1592 275 1654 276
rect 1688 275 1732 276
rect 1493 274 1553 275
rect 1590 274 1654 275
rect 1685 274 1732 275
rect 1493 273 1551 274
rect 1588 273 1654 274
rect 1683 273 1732 274
rect 1493 272 1549 273
rect 1586 272 1654 273
rect 1681 272 1732 273
rect 1493 271 1547 272
rect 1584 271 1653 272
rect 1678 271 1732 272
rect 1494 270 1545 271
rect 1582 270 1653 271
rect 1676 270 1732 271
rect 1494 269 1544 270
rect 1581 269 1653 270
rect 1673 269 1731 270
rect 1494 268 1542 269
rect 1579 268 1653 269
rect 1670 268 1731 269
rect 1494 267 1541 268
rect 1577 267 1652 268
rect 1667 267 1731 268
rect 1494 266 1540 267
rect 1575 266 1652 267
rect 1663 266 1731 267
rect 1494 265 1538 266
rect 1573 265 1652 266
rect 1659 265 1730 266
rect 1495 264 1537 265
rect 1571 264 1730 265
rect 1495 263 1536 264
rect 1569 263 1730 264
rect 1495 262 1535 263
rect 1568 262 1730 263
rect 1495 261 1534 262
rect 1566 261 1729 262
rect 1496 259 1533 261
rect 1564 260 1729 261
rect 1563 259 1729 260
rect 1496 258 1532 259
rect 1561 258 1728 259
rect 1497 256 1531 258
rect 1560 257 1728 258
rect 1558 256 1728 257
rect 1497 255 1530 256
rect 1557 255 1727 256
rect 1498 254 1530 255
rect 1556 254 1727 255
rect 1498 253 1529 254
rect 1554 253 1726 254
rect 1499 252 1529 253
rect 1553 252 1726 253
rect 1499 250 1528 252
rect 1552 251 1726 252
rect 1551 250 1725 251
rect 1500 248 1527 250
rect 1550 249 1616 250
rect 1617 249 1725 250
rect 1549 248 1614 249
rect 1501 247 1527 248
rect 1548 247 1613 248
rect 1617 247 1724 249
rect 1501 246 1526 247
rect 1547 246 1611 247
rect 1617 246 1723 247
rect 1502 244 1526 246
rect 1546 245 1609 246
rect 1616 245 1723 246
rect 1546 244 1608 245
rect 1616 244 1722 245
rect 1503 243 1526 244
rect 1545 243 1606 244
rect 1615 243 1722 244
rect 1503 242 1525 243
rect 1544 242 1605 243
rect 1615 242 1721 243
rect 1504 241 1525 242
rect 1505 239 1525 241
rect 1543 241 1603 242
rect 1543 240 1601 241
rect 1614 240 1720 242
rect 1542 239 1600 240
rect 1613 239 1719 240
rect 1506 237 1524 239
rect 1541 238 1598 239
rect 1612 238 1719 239
rect 1541 237 1597 238
rect 1612 237 1718 238
rect 1507 236 1524 237
rect 1508 234 1524 236
rect 1540 236 1595 237
rect 1611 236 1717 237
rect 1540 235 1594 236
rect 1610 235 1717 236
rect 1509 233 1524 234
rect 1539 234 1592 235
rect 1610 234 1716 235
rect 1539 233 1591 234
rect 1609 233 1715 234
rect 1510 232 1524 233
rect 1511 231 1524 232
rect 1538 232 1590 233
rect 1608 232 1657 233
rect 1658 232 1715 233
rect 1538 231 1589 232
rect 1607 231 1656 232
rect 1657 231 1714 232
rect 1512 229 1523 231
rect 1513 228 1523 229
rect 1537 230 1587 231
rect 1607 230 1654 231
rect 1657 230 1713 231
rect 1537 229 1586 230
rect 1606 229 1653 230
rect 1537 228 1585 229
rect 1605 228 1651 229
rect 1656 228 1712 230
rect 1514 227 1523 228
rect 1515 226 1523 227
rect 1516 225 1523 226
rect 1536 227 1584 228
rect 1604 227 1650 228
rect 1655 227 1711 228
rect 1536 226 1583 227
rect 1604 226 1649 227
rect 1655 226 1710 227
rect 1536 225 1582 226
rect 1603 225 1648 226
rect 1654 225 1709 226
rect 1517 224 1523 225
rect 1518 223 1523 224
rect 1519 222 1523 223
rect 1520 221 1523 222
rect 1535 224 1581 225
rect 1602 224 1646 225
rect 1654 224 1708 225
rect 1535 222 1580 224
rect 1601 223 1645 224
rect 1653 223 1707 224
rect 1601 222 1644 223
rect 1535 221 1579 222
rect 1600 221 1643 222
rect 1653 221 1706 223
rect 1521 220 1523 221
rect 1522 219 1523 220
rect 1534 220 1578 221
rect 1599 220 1642 221
rect 1652 220 1705 221
rect 1534 219 1577 220
rect 1599 219 1641 220
rect 1652 219 1704 220
rect 1534 217 1576 219
rect 1598 218 1640 219
rect 1652 218 1703 219
rect 1598 217 1639 218
rect 1652 217 1702 218
rect 1534 216 1575 217
rect 1597 216 1639 217
rect 1651 216 1701 217
rect 1533 214 1574 216
rect 1597 215 1638 216
rect 1651 215 1700 216
rect 1596 214 1637 215
rect 1651 214 1699 215
rect 1533 212 1573 214
rect 1596 213 1636 214
rect 1595 212 1636 213
rect 1651 213 1698 214
rect 1651 212 1697 213
rect 1533 210 1572 212
rect 1595 211 1635 212
rect 1650 211 1695 212
rect 1595 210 1634 211
rect 1533 207 1571 210
rect 1594 209 1634 210
rect 1650 210 1694 211
rect 1650 209 1693 210
rect 1594 208 1633 209
rect 1593 207 1633 208
rect 1650 208 1692 209
rect 1650 207 1691 208
rect 1533 206 1570 207
rect 1534 204 1570 206
rect 1593 206 1632 207
rect 1650 206 1690 207
rect 1593 205 1631 206
rect 1650 205 1688 206
rect 1534 203 1569 204
rect 1535 201 1569 203
rect 1592 203 1631 205
rect 1649 204 1687 205
rect 1649 203 1686 204
rect 1592 201 1630 203
rect 1649 202 1685 203
rect 1649 201 1683 202
rect 1536 200 1569 201
rect 1536 199 1568 200
rect 1537 197 1568 199
rect 1538 196 1568 197
rect 1591 198 1629 201
rect 1649 200 1682 201
rect 1649 199 1681 200
rect 1649 198 1679 199
rect 1591 196 1628 198
rect 1539 194 1568 196
rect 1540 193 1568 194
rect 1541 192 1568 193
rect 1542 190 1568 192
rect 1543 189 1568 190
rect 1544 188 1568 189
rect 1545 187 1568 188
rect 1546 186 1568 187
rect 1548 185 1568 186
rect 1549 184 1568 185
rect 1550 183 1568 184
rect 993 182 1061 183
rect 1162 182 1243 183
rect 1283 182 1351 183
rect 1552 182 1568 183
rect 1590 195 1628 196
rect 1649 197 1678 198
rect 1649 196 1676 197
rect 1649 195 1675 196
rect 1590 191 1627 195
rect 1649 194 1674 195
rect 1649 193 1672 194
rect 1649 192 1671 193
rect 1649 191 1670 192
rect 1590 185 1626 191
rect 1649 190 1669 191
rect 1649 189 1668 190
rect 1649 188 1667 189
rect 1650 187 1666 188
rect 1650 185 1665 187
rect 501 181 691 182
rect 813 181 878 182
rect 1163 181 1245 182
rect 1284 181 1350 182
rect 1553 181 1569 182
rect 1164 180 1245 181
rect 1554 180 1569 181
rect 1165 179 1247 180
rect 1556 179 1569 180
rect 1590 179 1625 185
rect 1650 184 1664 185
rect 1650 183 1663 184
rect 1650 181 1662 183
rect 1650 180 1661 181
rect 1166 178 1247 179
rect 1557 178 1569 179
rect 1167 177 1249 178
rect 1558 177 1569 178
rect 1168 176 1249 177
rect 1560 176 1569 177
rect 1169 175 1251 176
rect 1561 175 1570 176
rect 1170 174 1251 175
rect 1562 174 1570 175
rect 1591 174 1625 179
rect 1651 178 1660 180
rect 1651 177 1659 178
rect 1651 176 1658 177
rect 1171 173 1253 174
rect 1563 173 1570 174
rect 1172 172 1254 173
rect 1565 172 1570 173
rect 1173 171 1255 172
rect 1566 171 1571 172
rect 1592 171 1625 174
rect 1652 175 1658 176
rect 1652 173 1657 175
rect 1652 172 1656 173
rect 1174 170 1255 171
rect 1567 170 1571 171
rect 1569 169 1571 170
rect 1593 169 1625 171
rect 1653 171 1656 172
rect 1653 169 1655 171
rect 1570 168 1571 169
rect 1594 167 1625 169
rect 1595 166 1625 167
rect 1595 165 1626 166
rect 1596 163 1626 165
rect 1597 161 1626 163
rect 1598 160 1626 161
rect 1599 158 1627 160
rect 1600 157 1627 158
rect 1601 156 1627 157
rect 1602 155 1627 156
rect 1603 154 1628 155
rect 1604 153 1628 154
rect 1605 152 1628 153
rect 1606 151 1628 152
rect 1607 150 1629 151
rect 1608 149 1629 150
rect 1609 148 1629 149
rect 1610 147 1630 148
rect 1611 146 1630 147
rect 1613 145 1630 146
rect 1614 144 1631 145
rect 1615 143 1631 144
rect 1617 142 1631 143
rect 1618 141 1632 142
rect 1301 140 1314 141
rect 1620 140 1632 141
rect 487 139 511 140
rect 528 139 537 140
rect 734 139 743 140
rect 831 139 839 140
rect 486 137 512 139
rect 486 136 511 137
rect 486 133 512 136
rect 487 131 511 133
rect 477 127 522 128
rect 476 119 522 127
rect 477 118 521 119
rect 528 118 538 139
rect 584 136 638 137
rect 583 130 639 136
rect 683 134 720 135
rect 583 127 638 130
rect 627 121 638 127
rect 682 126 721 134
rect 683 125 720 126
rect 695 124 708 125
rect 695 123 707 124
rect 696 121 707 123
rect 733 122 743 139
rect 781 131 821 132
rect 781 125 822 131
rect 780 123 822 125
rect 781 122 822 123
rect 720 121 743 122
rect 795 121 807 122
rect 627 120 637 121
rect 528 117 539 118
rect 541 117 542 118
rect 543 117 545 118
rect 626 117 637 120
rect 695 119 707 121
rect 695 117 708 119
rect 493 115 506 116
rect 489 114 509 115
rect 487 113 512 114
rect 485 112 513 113
rect 483 111 515 112
rect 482 110 516 111
rect 481 109 517 110
rect 480 108 517 109
rect 480 107 518 108
rect 528 107 547 117
rect 626 114 636 117
rect 695 116 709 117
rect 694 114 709 116
rect 625 110 636 114
rect 693 113 710 114
rect 693 112 711 113
rect 719 112 743 121
rect 796 116 807 121
rect 692 111 712 112
rect 691 110 712 111
rect 624 109 636 110
rect 690 109 714 110
rect 576 108 646 109
rect 689 108 715 109
rect 479 106 496 107
rect 503 106 519 107
rect 479 105 492 106
rect 506 105 519 106
rect 478 104 491 105
rect 507 104 519 105
rect 478 99 490 104
rect 508 103 519 104
rect 528 106 539 107
rect 508 102 520 103
rect 508 101 519 102
rect 508 99 520 101
rect 479 98 491 99
rect 507 98 519 99
rect 479 97 493 98
rect 505 97 519 98
rect 480 96 496 97
rect 502 96 518 97
rect 480 95 518 96
rect 481 94 517 95
rect 482 93 516 94
rect 483 92 515 93
rect 484 91 514 92
rect 486 90 513 91
rect 488 89 510 90
rect 490 88 508 89
rect 487 83 497 84
rect 486 72 498 83
rect 528 82 538 106
rect 575 100 647 108
rect 688 107 716 108
rect 687 106 717 107
rect 686 105 701 106
rect 703 105 719 106
rect 685 104 700 105
rect 703 104 720 105
rect 683 103 700 104
rect 704 103 723 104
rect 682 102 699 103
rect 705 102 723 103
rect 680 101 698 102
rect 706 101 723 102
rect 678 100 697 101
rect 707 100 723 101
rect 576 99 646 100
rect 677 99 696 100
rect 709 99 722 100
rect 603 98 615 99
rect 678 98 695 99
rect 710 98 721 99
rect 604 88 614 98
rect 679 97 694 98
rect 711 97 721 98
rect 680 96 693 97
rect 712 96 720 97
rect 680 95 691 96
rect 715 95 719 96
rect 681 94 690 95
rect 716 94 719 95
rect 682 93 688 94
rect 683 92 687 93
rect 604 87 615 88
rect 584 86 637 87
rect 528 81 537 82
rect 583 77 638 86
rect 584 76 638 77
rect 486 71 538 72
rect 486 63 540 71
rect 487 62 540 63
rect 628 61 638 76
rect 691 73 701 88
rect 733 82 743 112
rect 795 111 807 116
rect 795 108 808 111
rect 794 107 808 108
rect 830 110 840 139
rect 886 130 940 138
rect 998 137 1007 138
rect 998 130 1008 137
rect 886 129 898 130
rect 900 129 901 130
rect 935 129 937 130
rect 886 128 897 129
rect 886 127 896 128
rect 886 126 897 127
rect 886 125 939 126
rect 886 119 940 125
rect 997 124 1008 130
rect 997 123 1009 124
rect 996 120 1009 123
rect 886 118 939 119
rect 886 117 898 118
rect 996 117 1010 120
rect 886 116 897 117
rect 995 116 1011 117
rect 886 115 896 116
rect 994 115 1011 116
rect 886 114 897 115
rect 994 114 1012 115
rect 886 113 898 114
rect 900 113 901 114
rect 938 113 939 114
rect 993 113 1012 114
rect 830 109 842 110
rect 844 109 845 110
rect 846 109 848 110
rect 794 105 809 107
rect 793 102 809 105
rect 793 101 810 102
rect 792 100 811 101
rect 791 98 811 100
rect 830 99 850 109
rect 886 105 941 113
rect 992 112 1013 113
rect 992 111 1014 112
rect 991 110 1015 111
rect 990 109 1016 110
rect 990 108 1017 109
rect 988 106 1002 108
rect 1004 107 1018 108
rect 1004 106 1019 107
rect 986 105 1001 106
rect 1005 105 1021 106
rect 887 104 940 105
rect 985 104 1000 105
rect 1006 104 1022 105
rect 907 101 919 104
rect 984 103 999 104
rect 1007 103 1024 104
rect 983 102 998 103
rect 1008 102 1026 103
rect 981 101 998 102
rect 1009 101 1026 102
rect 906 100 919 101
rect 980 100 997 101
rect 1010 100 1026 101
rect 879 99 904 100
rect 905 99 920 100
rect 921 99 944 100
rect 945 99 947 100
rect 978 99 996 100
rect 1011 99 1026 100
rect 830 98 849 99
rect 877 98 948 99
rect 978 98 995 99
rect 1012 98 1025 99
rect 791 97 812 98
rect 790 96 813 97
rect 789 95 813 96
rect 789 94 814 95
rect 788 93 801 94
rect 803 93 815 94
rect 787 91 800 93
rect 803 92 816 93
rect 803 91 817 92
rect 786 90 799 91
rect 804 90 818 91
rect 785 89 799 90
rect 805 89 819 90
rect 784 88 798 89
rect 805 88 820 89
rect 783 87 797 88
rect 806 87 821 88
rect 782 86 797 87
rect 807 86 822 87
rect 781 85 796 86
rect 807 85 823 86
rect 780 84 795 85
rect 808 84 824 85
rect 778 83 794 84
rect 809 83 825 84
rect 777 82 793 83
rect 810 82 824 83
rect 776 81 793 82
rect 811 81 823 82
rect 776 80 792 81
rect 812 80 822 81
rect 777 79 791 80
rect 813 79 822 80
rect 777 78 790 79
rect 814 78 821 79
rect 779 77 789 78
rect 816 77 820 78
rect 779 76 788 77
rect 817 76 819 77
rect 781 75 786 76
rect 782 74 785 75
rect 691 72 702 73
rect 691 62 745 72
rect 830 61 840 98
rect 877 91 949 98
rect 978 97 994 98
rect 1014 97 1024 98
rect 979 96 993 97
rect 1015 96 1024 97
rect 980 95 991 96
rect 1017 95 1023 96
rect 981 94 990 95
rect 1018 94 1022 95
rect 982 93 989 94
rect 983 92 988 93
rect 984 91 986 92
rect 877 90 948 91
rect 912 87 913 88
rect 993 87 998 88
rect 999 87 1001 88
rect 902 86 923 87
rect 896 85 929 86
rect 894 84 932 85
rect 891 83 934 84
rect 890 82 936 83
rect 888 81 937 82
rect 887 80 938 81
rect 886 79 940 80
rect 885 78 940 79
rect 885 77 903 78
rect 922 77 941 78
rect 884 76 900 77
rect 926 76 941 77
rect 884 71 897 76
rect 928 75 942 76
rect 929 74 942 75
rect 930 73 942 74
rect 929 71 942 73
rect 884 70 898 71
rect 928 70 942 71
rect 992 73 1002 87
rect 1034 82 1044 140
rect 1135 139 1144 140
rect 1297 139 1318 140
rect 1103 137 1104 138
rect 1096 136 1107 137
rect 1093 135 1111 136
rect 1091 134 1112 135
rect 1090 133 1114 134
rect 1089 132 1115 133
rect 1088 131 1116 132
rect 1087 130 1117 131
rect 1134 130 1145 139
rect 1296 138 1319 139
rect 1294 137 1321 138
rect 1293 136 1322 137
rect 1086 129 1145 130
rect 1085 128 1145 129
rect 1084 127 1100 128
rect 1103 127 1145 128
rect 1084 126 1098 127
rect 1106 126 1145 127
rect 1187 126 1243 136
rect 1292 135 1323 136
rect 1291 134 1324 135
rect 1290 133 1325 134
rect 1289 132 1325 133
rect 1289 131 1302 132
rect 1313 131 1326 132
rect 1289 130 1301 131
rect 1314 130 1326 131
rect 1289 129 1300 130
rect 1315 129 1327 130
rect 1084 125 1096 126
rect 1108 125 1145 126
rect 1231 125 1243 126
rect 1083 124 1095 125
rect 1109 124 1145 125
rect 1232 124 1242 125
rect 1083 123 1094 124
rect 1082 122 1094 123
rect 1110 122 1145 124
rect 1082 120 1093 122
rect 1111 120 1145 122
rect 1082 113 1092 120
rect 1111 119 1122 120
rect 1134 119 1145 120
rect 1112 114 1122 119
rect 1135 118 1145 119
rect 1134 114 1145 118
rect 1231 119 1242 124
rect 1288 123 1299 129
rect 1316 127 1327 129
rect 1317 125 1327 127
rect 1316 123 1327 125
rect 1289 122 1300 123
rect 1315 122 1327 123
rect 1289 121 1302 122
rect 1313 121 1326 122
rect 1289 120 1303 121
rect 1312 120 1326 121
rect 1289 119 1325 120
rect 1231 115 1241 119
rect 1290 118 1325 119
rect 1291 117 1324 118
rect 1291 116 1323 117
rect 1293 115 1322 116
rect 1082 112 1093 113
rect 1111 112 1145 114
rect 1082 110 1094 112
rect 1110 110 1145 112
rect 1230 111 1241 115
rect 1294 114 1321 115
rect 1296 113 1319 114
rect 1297 112 1318 113
rect 1302 111 1314 112
rect 1230 110 1240 111
rect 1083 109 1094 110
rect 1109 109 1145 110
rect 1083 108 1096 109
rect 1108 108 1145 109
rect 1084 107 1097 108
rect 1107 107 1145 108
rect 1084 106 1099 107
rect 1105 106 1145 107
rect 1084 105 1145 106
rect 1085 104 1145 105
rect 1229 108 1240 110
rect 1330 109 1334 110
rect 1323 108 1335 109
rect 1229 104 1239 108
rect 1283 106 1335 108
rect 1086 103 1118 104
rect 1134 103 1145 104
rect 1228 103 1239 104
rect 1087 102 1117 103
rect 1135 102 1145 103
rect 1180 102 1250 103
rect 1088 101 1116 102
rect 1089 100 1115 101
rect 1090 99 1113 100
rect 1092 98 1112 99
rect 1094 97 1109 98
rect 1096 96 1107 97
rect 1092 73 1102 88
rect 1134 83 1145 102
rect 1179 94 1251 102
rect 1282 100 1335 106
rect 1282 99 1331 100
rect 1283 98 1324 99
rect 1298 97 1310 98
rect 1337 97 1347 140
rect 1622 139 1632 140
rect 1623 138 1633 139
rect 1625 137 1633 138
rect 1627 136 1634 137
rect 1629 135 1634 136
rect 1632 134 1635 135
rect 1638 102 1651 103
rect 1412 99 1433 102
rect 1439 99 1457 102
rect 1462 100 1482 102
rect 1463 99 1482 100
rect 1490 99 1506 102
rect 1512 100 1533 102
rect 1542 100 1560 102
rect 1564 101 1578 102
rect 1596 101 1613 102
rect 1634 101 1656 102
rect 1564 100 1579 101
rect 1596 100 1614 101
rect 1631 100 1658 101
rect 1512 99 1532 100
rect 1543 99 1560 100
rect 1565 99 1579 100
rect 1597 99 1613 100
rect 1629 99 1640 100
rect 1647 99 1658 100
rect 1684 99 1705 102
rect 1712 100 1733 102
rect 1713 99 1733 100
rect 1742 100 1774 102
rect 1742 99 1775 100
rect 1785 99 1818 102
rect 1416 98 1429 99
rect 1443 98 1453 99
rect 1466 98 1479 99
rect 1494 98 1503 99
rect 1516 98 1529 99
rect 1546 98 1557 99
rect 1568 98 1580 99
rect 1601 98 1610 99
rect 1628 98 1637 99
rect 1650 98 1658 99
rect 1688 98 1701 99
rect 1717 98 1729 99
rect 1746 98 1757 99
rect 1766 98 1775 99
rect 1789 98 1801 99
rect 1809 98 1818 99
rect 1417 97 1428 98
rect 1443 97 1450 98
rect 1467 97 1478 98
rect 1494 97 1501 98
rect 1517 97 1528 98
rect 1547 97 1556 98
rect 1570 97 1581 98
rect 1602 97 1609 98
rect 1626 97 1636 98
rect 1651 97 1659 98
rect 1689 97 1700 98
rect 1717 97 1728 98
rect 1299 96 1310 97
rect 1180 93 1250 94
rect 1207 92 1219 93
rect 1135 82 1144 83
rect 992 72 1003 73
rect 1092 72 1103 73
rect 992 71 1045 72
rect 885 69 901 70
rect 925 69 941 70
rect 885 68 905 69
rect 922 68 941 69
rect 886 67 940 68
rect 887 66 940 67
rect 888 65 939 66
rect 889 64 938 65
rect 891 63 936 64
rect 892 62 934 63
rect 992 62 1046 71
rect 1092 62 1146 72
rect 895 61 931 62
rect 1208 61 1219 92
rect 1299 85 1309 96
rect 1322 95 1324 96
rect 1327 95 1334 96
rect 1336 95 1347 97
rect 1321 94 1347 95
rect 1320 87 1347 94
rect 1321 86 1347 87
rect 1336 85 1347 86
rect 1300 84 1302 85
rect 1303 84 1308 85
rect 1294 81 1304 82
rect 1294 72 1305 81
rect 1337 80 1347 85
rect 1418 81 1427 97
rect 1442 96 1449 97
rect 1468 96 1479 97
rect 1442 95 1447 96
rect 1469 95 1479 96
rect 1494 96 1500 97
rect 1494 95 1499 96
rect 1441 94 1446 95
rect 1469 94 1480 95
rect 1494 94 1498 95
rect 1440 93 1445 94
rect 1470 93 1480 94
rect 1493 93 1498 94
rect 1439 92 1444 93
rect 1470 92 1481 93
rect 1493 92 1497 93
rect 1439 91 1443 92
rect 1471 91 1481 92
rect 1492 91 1497 92
rect 1438 90 1442 91
rect 1437 89 1441 90
rect 1472 89 1482 91
rect 1492 90 1496 91
rect 1436 88 1440 89
rect 1435 87 1439 88
rect 1473 87 1483 89
rect 1491 88 1495 90
rect 1434 86 1438 87
rect 1433 85 1437 86
rect 1474 85 1484 87
rect 1490 86 1494 88
rect 1489 85 1493 86
rect 1432 84 1436 85
rect 1475 84 1485 85
rect 1489 84 1492 85
rect 1431 83 1437 84
rect 1430 82 1437 83
rect 1476 83 1485 84
rect 1488 83 1492 84
rect 1476 82 1486 83
rect 1488 82 1491 83
rect 1428 81 1438 82
rect 1477 81 1486 82
rect 1487 81 1491 82
rect 1418 80 1439 81
rect 1477 80 1490 81
rect 1418 78 1440 80
rect 1478 79 1490 80
rect 1478 78 1489 79
rect 1294 71 1348 72
rect 1294 63 1349 71
rect 1294 62 1348 63
rect 1418 62 1427 78
rect 1429 77 1441 78
rect 1430 76 1442 77
rect 1431 75 1442 76
rect 1432 74 1443 75
rect 1432 73 1444 74
rect 1433 72 1445 73
rect 1434 71 1445 72
rect 1434 70 1446 71
rect 1435 69 1447 70
rect 1436 67 1448 69
rect 1437 66 1449 67
rect 1438 65 1450 66
rect 1439 64 1451 65
rect 1439 63 1452 64
rect 1440 62 1452 63
rect 1417 61 1428 62
rect 1441 61 1454 62
rect 1479 61 1489 78
rect 1517 73 1527 97
rect 1548 92 1555 97
rect 1570 96 1582 97
rect 1571 95 1583 96
rect 1571 94 1584 95
rect 1571 92 1585 94
rect 1548 91 1554 92
rect 1549 73 1554 91
rect 1518 71 1527 73
rect 1518 67 1528 71
rect 1548 69 1554 73
rect 1571 91 1586 92
rect 1603 91 1608 97
rect 1625 96 1634 97
rect 1652 96 1659 97
rect 1624 95 1633 96
rect 1653 95 1659 96
rect 1623 94 1632 95
rect 1654 94 1659 95
rect 1622 93 1632 94
rect 1621 92 1631 93
rect 1655 92 1659 94
rect 1571 90 1587 91
rect 1548 68 1553 69
rect 1519 65 1529 67
rect 1547 65 1553 68
rect 1519 64 1530 65
rect 1546 64 1552 65
rect 1520 63 1531 64
rect 1545 63 1552 64
rect 1571 64 1575 90
rect 1576 89 1588 90
rect 1577 88 1589 89
rect 1577 87 1590 88
rect 1578 86 1591 87
rect 1579 85 1592 86
rect 1580 84 1592 85
rect 1581 83 1593 84
rect 1582 82 1594 83
rect 1583 81 1595 82
rect 1583 80 1596 81
rect 1584 79 1597 80
rect 1585 78 1598 79
rect 1586 77 1599 78
rect 1587 76 1599 77
rect 1588 75 1600 76
rect 1588 74 1601 75
rect 1589 73 1602 74
rect 1590 72 1603 73
rect 1604 72 1607 91
rect 1620 90 1630 92
rect 1619 87 1629 90
rect 1656 89 1659 92
rect 1690 95 1700 97
rect 1618 86 1629 87
rect 1618 84 1628 86
rect 1617 74 1628 84
rect 1690 83 1699 95
rect 1718 83 1728 97
rect 1690 79 1728 83
rect 1642 78 1662 79
rect 1690 78 1700 79
rect 1642 76 1663 78
rect 1645 75 1661 76
rect 1648 74 1660 75
rect 1591 71 1607 72
rect 1592 70 1607 71
rect 1618 70 1629 74
rect 1649 72 1659 74
rect 1593 68 1607 70
rect 1619 68 1630 70
rect 1594 67 1607 68
rect 1595 66 1607 67
rect 1620 66 1631 68
rect 1596 65 1607 66
rect 1621 65 1632 66
rect 1597 64 1607 65
rect 1622 64 1633 65
rect 1571 63 1576 64
rect 1520 62 1532 63
rect 1544 62 1551 63
rect 1521 61 1534 62
rect 1542 61 1551 62
rect 1570 61 1576 63
rect 1598 62 1607 64
rect 1623 63 1633 64
rect 1650 63 1659 72
rect 1624 62 1634 63
rect 1599 61 1607 62
rect 1625 61 1636 62
rect 628 60 637 61
rect 831 60 839 61
rect 897 60 929 61
rect 1209 60 1218 61
rect 1417 60 1429 61
rect 1441 60 1455 61
rect 1478 60 1490 61
rect 1522 60 1550 61
rect 1569 60 1577 61
rect 1600 60 1607 61
rect 1626 60 1637 61
rect 1649 60 1659 63
rect 1690 63 1699 78
rect 1690 62 1700 63
rect 1689 61 1700 62
rect 1718 61 1728 79
rect 1747 82 1757 98
rect 1769 97 1775 98
rect 1770 96 1775 97
rect 1771 94 1775 96
rect 1772 91 1775 94
rect 1769 86 1771 87
rect 1768 83 1771 86
rect 1767 82 1771 83
rect 1747 78 1771 82
rect 1747 61 1757 78
rect 1767 77 1771 78
rect 1768 74 1771 77
rect 1769 73 1771 74
rect 1790 82 1800 98
rect 1812 97 1818 98
rect 1813 96 1818 97
rect 1814 94 1818 96
rect 1815 91 1818 94
rect 1812 85 1815 87
rect 1811 83 1815 85
rect 1810 82 1815 83
rect 1790 78 1815 82
rect 1776 68 1778 69
rect 1775 66 1778 68
rect 1774 64 1778 66
rect 1773 63 1778 64
rect 1772 62 1777 63
rect 1771 61 1777 62
rect 1790 62 1800 78
rect 1810 77 1815 78
rect 1811 75 1815 77
rect 1812 73 1815 75
rect 1819 68 1822 69
rect 1818 67 1822 68
rect 1818 66 1821 67
rect 1817 64 1821 66
rect 1816 63 1821 64
rect 1815 62 1821 63
rect 1790 61 1801 62
rect 1814 61 1820 62
rect 1689 60 1701 61
rect 1717 60 1729 61
rect 1746 60 1759 61
rect 1769 60 1777 61
rect 1789 60 1802 61
rect 1812 60 1820 61
rect 904 59 923 60
rect 1413 59 1433 60
rect 1442 59 1458 60
rect 1474 59 1494 60
rect 1523 59 1549 60
rect 1566 59 1581 60
rect 1601 59 1607 60
rect 1628 59 1640 60
rect 1648 59 1659 60
rect 1685 59 1704 60
rect 1713 59 1733 60
rect 1412 57 1433 59
rect 1443 57 1458 59
rect 1473 57 1496 59
rect 1524 58 1548 59
rect 1526 57 1546 58
rect 1565 57 1582 59
rect 1602 58 1607 59
rect 1630 58 1659 59
rect 1529 56 1543 57
rect 1603 56 1607 58
rect 1632 57 1656 58
rect 1684 57 1705 59
rect 1712 57 1733 59
rect 1741 58 1777 60
rect 1785 59 1820 60
rect 1784 58 1820 59
rect 1741 57 1776 58
rect 1784 57 1819 58
rect 1636 56 1651 57
rect 499 45 502 46
rect 712 45 715 46
rect 766 45 768 46
rect 1188 45 1191 46
rect 479 42 493 43
rect 478 39 494 42
rect 478 38 493 39
rect 478 37 485 38
rect 478 32 484 37
rect 478 31 485 32
rect 478 29 492 31
rect 478 27 493 29
rect 478 25 492 27
rect 478 24 485 25
rect 478 18 484 24
rect 478 17 492 18
rect 478 16 493 17
rect 478 13 494 16
rect 497 13 502 45
rect 611 44 613 45
rect 545 40 548 41
rect 543 39 548 40
rect 609 39 614 44
rect 512 35 517 36
rect 531 35 536 36
rect 542 35 548 39
rect 610 38 614 39
rect 563 35 565 36
rect 573 35 578 36
rect 596 35 601 36
rect 624 35 629 36
rect 638 35 643 36
rect 663 35 669 36
rect 687 35 690 36
rect 704 35 707 36
rect 710 35 716 45
rect 728 42 746 43
rect 727 41 746 42
rect 727 39 747 41
rect 727 38 746 39
rect 733 37 741 38
rect 510 34 519 35
rect 529 34 538 35
rect 540 34 551 35
rect 555 34 558 35
rect 561 34 566 35
rect 571 34 580 35
rect 589 34 592 35
rect 594 34 602 35
rect 610 34 614 35
rect 622 34 631 35
rect 636 34 645 35
rect 660 34 671 35
rect 678 34 692 35
rect 701 34 716 35
rect 508 33 520 34
rect 528 33 552 34
rect 508 32 521 33
rect 527 32 552 33
rect 507 31 521 32
rect 526 31 552 32
rect 506 30 522 31
rect 526 30 538 31
rect 540 30 551 31
rect 554 30 566 34
rect 570 33 582 34
rect 569 32 582 33
rect 568 31 583 32
rect 588 31 604 34
rect 568 30 584 31
rect 506 29 512 30
rect 516 29 522 30
rect 506 27 511 29
rect 506 26 512 27
rect 517 26 522 29
rect 525 28 532 30
rect 525 27 531 28
rect 506 23 523 26
rect 506 21 522 23
rect 524 21 530 27
rect 506 19 511 21
rect 524 20 531 21
rect 525 19 531 20
rect 506 18 512 19
rect 525 18 532 19
rect 542 18 548 30
rect 554 29 574 30
rect 578 29 584 30
rect 588 30 605 31
rect 554 28 562 29
rect 566 28 573 29
rect 578 28 585 29
rect 554 27 561 28
rect 506 17 513 18
rect 518 17 521 18
rect 526 17 533 18
rect 536 17 538 18
rect 507 15 522 17
rect 526 16 538 17
rect 542 17 549 18
rect 542 16 552 17
rect 526 15 539 16
rect 543 15 552 16
rect 508 14 521 15
rect 527 14 539 15
rect 509 13 521 14
rect 528 13 539 14
rect 544 13 552 15
rect 554 13 560 27
rect 566 19 572 28
rect 579 26 585 28
rect 580 22 585 26
rect 579 19 585 22
rect 566 18 573 19
rect 578 18 585 19
rect 588 28 595 30
rect 599 28 605 30
rect 567 17 574 18
rect 577 17 584 18
rect 568 16 584 17
rect 568 15 583 16
rect 569 14 582 15
rect 570 13 581 14
rect 588 13 594 28
rect 600 13 605 28
rect 609 13 614 34
rect 621 33 631 34
rect 620 32 631 33
rect 634 32 646 34
rect 660 33 672 34
rect 678 33 693 34
rect 700 33 716 34
rect 619 31 631 32
rect 633 31 646 32
rect 659 32 673 33
rect 619 30 630 31
rect 633 30 645 31
rect 659 30 674 32
rect 618 28 625 30
rect 633 29 639 30
rect 659 29 662 30
rect 668 29 674 30
rect 632 28 639 29
rect 660 28 661 29
rect 618 25 624 28
rect 633 27 639 28
rect 669 27 674 29
rect 633 26 641 27
rect 663 26 674 27
rect 633 25 643 26
rect 661 25 674 26
rect 618 22 623 25
rect 634 24 644 25
rect 660 24 674 25
rect 634 23 645 24
rect 659 23 674 24
rect 635 22 646 23
rect 618 19 624 22
rect 638 21 646 22
rect 639 20 646 21
rect 658 22 674 23
rect 658 21 664 22
rect 658 20 663 21
rect 669 20 674 22
rect 618 18 625 19
rect 618 17 626 18
rect 629 17 631 18
rect 634 17 636 18
rect 640 17 646 20
rect 657 18 663 20
rect 668 18 674 20
rect 619 15 632 17
rect 620 14 632 15
rect 621 13 632 14
rect 633 15 646 17
rect 658 17 664 18
rect 667 17 674 18
rect 658 15 674 17
rect 633 14 645 15
rect 659 14 674 15
rect 633 13 644 14
rect 660 13 674 14
rect 678 31 694 33
rect 678 30 695 31
rect 699 30 716 33
rect 678 29 685 30
rect 688 29 695 30
rect 678 26 684 29
rect 479 12 493 13
rect 498 12 502 13
rect 511 12 520 13
rect 529 12 538 13
rect 545 12 552 13
rect 555 12 559 13
rect 571 12 580 13
rect 589 12 593 13
rect 600 12 604 13
rect 610 12 614 13
rect 622 12 631 13
rect 634 12 643 13
rect 660 12 667 13
rect 670 12 673 13
rect 678 12 683 26
rect 689 13 695 29
rect 698 29 705 30
rect 708 29 716 30
rect 698 25 704 29
rect 709 27 716 29
rect 698 22 703 25
rect 698 19 704 22
rect 710 20 716 27
rect 698 18 705 19
rect 709 18 716 20
rect 698 17 706 18
rect 708 17 716 18
rect 699 15 716 17
rect 700 14 716 15
rect 701 13 716 14
rect 734 13 740 37
rect 750 35 755 36
rect 748 34 757 35
rect 747 33 758 34
rect 746 32 759 33
rect 745 31 759 32
rect 745 30 760 31
rect 744 29 750 30
rect 744 27 749 29
rect 755 28 760 30
rect 743 26 750 27
rect 755 26 761 28
rect 743 22 761 26
rect 743 21 760 22
rect 743 20 750 21
rect 744 19 749 20
rect 744 18 750 19
rect 744 17 751 18
rect 756 17 760 18
rect 745 15 760 17
rect 746 14 760 15
rect 747 13 759 14
rect 764 13 769 45
rect 933 44 936 45
rect 991 44 993 45
rect 1187 44 1192 45
rect 1278 44 1280 45
rect 932 39 937 44
rect 979 40 982 41
rect 978 39 982 40
rect 989 39 994 44
rect 1066 42 1078 43
rect 933 38 936 39
rect 977 36 982 39
rect 990 38 994 39
rect 1065 41 1080 42
rect 1065 40 1081 41
rect 1065 38 1082 40
rect 1065 37 1072 38
rect 1074 37 1082 38
rect 779 35 783 36
rect 798 35 803 36
rect 814 35 818 36
rect 837 35 840 36
rect 847 35 851 36
rect 867 35 871 36
rect 878 35 882 36
rect 919 35 924 36
rect 947 35 952 36
rect 961 35 967 36
rect 976 35 983 36
rect 1005 35 1010 36
rect 1029 35 1032 36
rect 1045 35 1050 36
rect 776 34 785 35
rect 796 34 805 35
rect 811 34 821 35
rect 829 34 833 35
rect 835 34 842 35
rect 846 34 853 35
rect 860 34 873 35
rect 876 34 884 35
rect 891 34 895 35
rect 902 34 906 35
rect 911 34 915 35
rect 917 34 925 35
rect 932 34 936 35
rect 945 34 954 35
rect 959 34 969 35
rect 974 34 986 35
rect 990 34 994 35
rect 1003 34 1012 35
rect 1020 34 1024 35
rect 1026 34 1034 35
rect 1043 34 1052 35
rect 775 32 787 34
rect 795 33 805 34
rect 810 33 822 34
rect 829 33 843 34
rect 844 33 854 34
rect 794 32 805 33
rect 774 31 788 32
rect 773 30 788 31
rect 793 31 805 32
rect 809 32 823 33
rect 809 31 824 32
rect 793 30 804 31
rect 808 30 825 31
rect 773 29 779 30
rect 783 29 789 30
rect 773 27 778 29
rect 772 26 778 27
rect 784 26 789 29
rect 792 29 799 30
rect 807 29 814 30
rect 818 29 825 30
rect 792 28 798 29
rect 772 21 789 26
rect 772 19 778 21
rect 791 20 797 28
rect 807 26 813 29
rect 819 27 825 29
rect 829 30 855 33
rect 829 27 835 30
rect 839 29 846 30
rect 849 29 855 30
rect 807 24 812 26
rect 806 23 812 24
rect 807 22 812 23
rect 791 19 798 20
rect 807 19 813 22
rect 820 21 826 27
rect 773 18 779 19
rect 792 18 799 19
rect 807 18 814 19
rect 819 18 825 21
rect 773 17 780 18
rect 784 17 788 18
rect 792 17 800 18
rect 803 17 805 18
rect 807 17 815 18
rect 818 17 825 18
rect 773 16 789 17
rect 774 15 788 16
rect 793 15 805 17
rect 808 16 824 17
rect 775 14 788 15
rect 794 14 805 15
rect 809 15 824 16
rect 809 14 823 15
rect 776 13 788 14
rect 795 13 805 14
rect 811 13 822 14
rect 829 13 834 27
rect 839 13 845 29
rect 850 15 855 29
rect 859 31 885 34
rect 859 30 886 31
rect 859 29 866 30
rect 869 29 877 30
rect 850 14 856 15
rect 850 13 855 14
rect 859 13 865 29
rect 869 27 876 29
rect 880 28 886 30
rect 870 13 875 27
rect 881 15 886 28
rect 890 19 895 34
rect 901 19 907 34
rect 890 18 896 19
rect 900 18 907 19
rect 890 17 897 18
rect 899 17 907 18
rect 890 15 907 17
rect 880 14 886 15
rect 891 14 907 15
rect 881 13 886 14
rect 892 13 907 14
rect 911 33 926 34
rect 911 30 927 33
rect 911 29 918 30
rect 921 29 928 30
rect 911 26 917 29
rect 911 15 916 26
rect 911 14 917 15
rect 690 12 694 13
rect 702 12 709 13
rect 711 12 715 13
rect 735 12 739 13
rect 748 12 758 13
rect 765 12 769 13
rect 777 12 787 13
rect 796 12 805 13
rect 812 12 821 13
rect 829 12 833 13
rect 840 12 844 13
rect 851 12 855 13
rect 860 12 864 13
rect 871 12 874 13
rect 881 12 885 13
rect 893 12 900 13
rect 903 12 906 13
rect 911 12 916 14
rect 922 13 928 29
rect 932 13 937 34
rect 944 33 954 34
rect 943 32 954 33
rect 942 31 954 32
rect 957 33 970 34
rect 957 31 971 33
rect 974 31 987 34
rect 941 30 953 31
rect 957 30 972 31
rect 975 30 986 31
rect 941 29 948 30
rect 958 29 960 30
rect 966 29 972 30
rect 941 28 947 29
rect 940 27 947 28
rect 967 27 972 29
rect 940 20 946 27
rect 961 26 972 27
rect 959 25 972 26
rect 957 24 972 25
rect 956 22 972 24
rect 956 21 962 22
rect 940 19 947 20
rect 941 18 947 19
rect 955 18 961 21
rect 967 20 972 22
rect 966 18 972 20
rect 941 17 949 18
rect 952 17 954 18
rect 942 15 954 17
rect 956 17 962 18
rect 965 17 972 18
rect 956 15 972 17
rect 977 20 982 30
rect 977 18 983 20
rect 977 17 984 18
rect 977 16 986 17
rect 943 14 954 15
rect 944 13 954 14
rect 957 13 972 15
rect 978 14 987 16
rect 979 13 987 14
rect 989 13 994 34
rect 1001 33 1013 34
rect 1020 33 1035 34
rect 1041 33 1052 34
rect 1000 32 1014 33
rect 1019 32 1036 33
rect 1000 31 1015 32
rect 999 30 1015 31
rect 1020 30 1036 32
rect 1040 30 1052 33
rect 1065 31 1071 37
rect 1075 36 1082 37
rect 1076 35 1082 36
rect 1092 35 1096 36
rect 1109 35 1115 36
rect 1126 35 1131 36
rect 1145 35 1150 36
rect 1167 35 1169 36
rect 1177 35 1183 36
rect 1187 35 1193 44
rect 1218 42 1223 43
rect 1196 35 1199 36
rect 1077 33 1082 35
rect 1090 34 1099 35
rect 1107 34 1117 35
rect 1124 34 1133 35
rect 1142 34 1152 35
rect 1160 34 1163 35
rect 1166 34 1170 35
rect 1175 34 1184 35
rect 1187 34 1201 35
rect 1076 31 1082 33
rect 1088 32 1100 34
rect 1106 33 1117 34
rect 1123 33 1134 34
rect 1087 31 1101 32
rect 1105 31 1117 33
rect 1122 32 1135 33
rect 1121 31 1136 32
rect 1065 30 1072 31
rect 1074 30 1082 31
rect 1086 30 1102 31
rect 998 29 1005 30
rect 1009 29 1016 30
rect 998 26 1004 29
rect 1010 27 1016 29
rect 1019 29 1027 30
rect 1030 29 1036 30
rect 1019 27 1026 29
rect 1011 26 1016 27
rect 1020 26 1026 27
rect 998 21 1003 26
rect 1011 21 1017 26
rect 998 19 1004 21
rect 1011 20 1016 21
rect 1020 20 1025 26
rect 1031 25 1037 29
rect 1039 27 1046 30
rect 1065 29 1081 30
rect 1086 29 1092 30
rect 1096 29 1102 30
rect 1105 30 1112 31
rect 1113 30 1116 31
rect 1121 30 1128 31
rect 1129 30 1136 31
rect 1105 29 1110 30
rect 1032 24 1037 25
rect 1040 26 1048 27
rect 1040 25 1050 26
rect 1040 24 1051 25
rect 1065 24 1080 29
rect 1086 26 1091 29
rect 1097 26 1102 29
rect 1104 28 1110 29
rect 1120 28 1126 30
rect 1131 29 1136 30
rect 1141 31 1154 34
rect 1141 30 1155 31
rect 1141 29 1143 30
rect 1149 29 1155 30
rect 1131 28 1137 29
rect 1104 27 1111 28
rect 1120 27 1125 28
rect 1132 27 1137 28
rect 1150 27 1155 29
rect 1104 26 1113 27
rect 1120 26 1126 27
rect 1131 26 1137 27
rect 1144 26 1155 27
rect 1085 25 1102 26
rect 1105 25 1115 26
rect 998 18 1005 19
rect 1010 18 1016 20
rect 998 17 1006 18
rect 1008 17 1016 18
rect 1019 17 1025 20
rect 1031 17 1037 24
rect 1041 23 1052 24
rect 1042 22 1053 23
rect 1045 21 1053 22
rect 1046 20 1053 21
rect 1047 18 1053 20
rect 999 16 1015 17
rect 1000 15 1014 16
rect 1020 15 1025 17
rect 1032 16 1037 17
rect 1001 14 1014 15
rect 1019 14 1026 15
rect 1002 13 1013 14
rect 1020 13 1025 14
rect 1031 13 1037 16
rect 1040 17 1042 18
rect 1046 17 1053 18
rect 1040 16 1053 17
rect 1040 14 1052 16
rect 1040 13 1051 14
rect 1065 13 1071 24
rect 1074 23 1081 24
rect 1075 22 1081 23
rect 1085 22 1103 25
rect 1105 24 1116 25
rect 1106 23 1117 24
rect 1107 22 1117 23
rect 1075 20 1082 22
rect 1085 21 1102 22
rect 1110 21 1118 22
rect 1085 20 1091 21
rect 1111 20 1118 21
rect 1076 18 1082 20
rect 1086 19 1091 20
rect 1086 18 1092 19
rect 1112 18 1118 20
rect 1120 21 1137 26
rect 1142 25 1155 26
rect 1141 24 1155 25
rect 1140 22 1155 24
rect 1139 21 1145 22
rect 1120 18 1126 21
rect 1134 18 1135 19
rect 1139 18 1144 21
rect 1150 19 1155 22
rect 1149 18 1155 19
rect 1076 17 1083 18
rect 1086 17 1093 18
rect 1098 17 1102 18
rect 1077 15 1083 17
rect 1087 15 1102 17
rect 1105 17 1107 18
rect 1111 17 1118 18
rect 1105 16 1118 17
rect 1121 17 1127 18
rect 1132 17 1136 18
rect 1105 15 1117 16
rect 1121 15 1136 17
rect 1139 17 1145 18
rect 1148 17 1155 18
rect 1139 15 1155 17
rect 1159 30 1170 34
rect 1174 33 1185 34
rect 1187 33 1202 34
rect 1173 32 1184 33
rect 1172 30 1184 32
rect 1187 31 1203 33
rect 1187 30 1204 31
rect 1159 29 1169 30
rect 1171 29 1179 30
rect 1159 27 1166 29
rect 1171 28 1178 29
rect 1187 28 1194 30
rect 1198 28 1204 30
rect 1077 14 1084 15
rect 1088 14 1101 15
rect 1104 14 1116 15
rect 1122 14 1136 15
rect 1140 14 1156 15
rect 1078 13 1084 14
rect 1089 13 1101 14
rect 1105 13 1116 14
rect 1123 13 1136 14
rect 1141 13 1156 14
rect 1159 13 1165 27
rect 1171 26 1177 28
rect 1171 22 1176 26
rect 1171 19 1177 22
rect 1171 18 1178 19
rect 1171 17 1179 18
rect 1183 17 1184 18
rect 1172 16 1185 17
rect 1173 14 1185 16
rect 1174 13 1185 14
rect 1187 13 1193 28
rect 1199 13 1204 28
rect 1217 15 1223 42
rect 1267 40 1270 41
rect 1265 36 1270 40
rect 1277 39 1282 44
rect 1290 40 1293 41
rect 1324 40 1327 41
rect 1277 38 1281 39
rect 1288 36 1293 40
rect 1323 39 1327 40
rect 1236 35 1240 36
rect 1252 35 1258 36
rect 1265 35 1271 36
rect 1287 35 1293 36
rect 1322 36 1327 39
rect 1659 37 1665 38
rect 1695 37 1697 38
rect 1712 37 1714 38
rect 1491 36 1501 37
rect 1506 36 1514 37
rect 1521 36 1528 37
rect 1536 36 1545 37
rect 1552 36 1562 37
rect 1570 36 1580 37
rect 1585 36 1593 37
rect 1601 36 1616 37
rect 1626 36 1641 37
rect 1657 36 1667 37
rect 1676 36 1686 37
rect 1695 36 1714 37
rect 1722 36 1732 37
rect 1735 36 1743 37
rect 1322 35 1328 36
rect 1339 35 1344 36
rect 1493 35 1499 36
rect 1508 35 1513 36
rect 1523 35 1529 36
rect 1539 35 1543 36
rect 1554 35 1560 36
rect 1572 35 1579 36
rect 1587 35 1591 36
rect 1228 34 1241 35
rect 1250 34 1259 35
rect 1262 34 1273 35
rect 1227 32 1243 34
rect 1249 33 1259 34
rect 1248 32 1260 33
rect 1227 30 1244 32
rect 1227 28 1234 30
rect 1238 28 1244 30
rect 1217 14 1224 15
rect 1217 13 1223 14
rect 1227 13 1233 28
rect 1239 15 1244 28
rect 1247 30 1259 32
rect 1261 31 1274 34
rect 1262 30 1273 31
rect 1247 28 1253 30
rect 1247 27 1254 28
rect 1247 26 1256 27
rect 1247 25 1258 26
rect 1248 24 1259 25
rect 1249 23 1260 24
rect 1250 22 1260 23
rect 1252 21 1261 22
rect 1254 20 1261 21
rect 1255 18 1261 20
rect 1248 17 1250 18
rect 1254 17 1261 18
rect 1265 20 1270 30
rect 1265 17 1271 20
rect 1247 15 1260 17
rect 1265 16 1274 17
rect 1265 15 1275 16
rect 1239 14 1245 15
rect 1247 14 1259 15
rect 1266 14 1275 15
rect 923 12 927 13
rect 933 12 936 13
rect 945 12 954 13
rect 959 12 965 13
rect 968 12 972 13
rect 980 12 986 13
rect 990 12 994 13
rect 1003 12 1011 13
rect 1020 12 1024 13
rect 1032 12 1036 13
rect 1040 12 1050 13
rect 1066 12 1070 13
rect 1078 12 1083 13
rect 1090 12 1100 13
rect 1106 12 1115 13
rect 1125 12 1135 13
rect 1142 12 1149 13
rect 1152 12 1155 13
rect 1160 12 1164 13
rect 1176 12 1184 13
rect 1188 12 1192 13
rect 1200 12 1203 13
rect 1218 12 1223 13
rect 1228 12 1231 13
rect 1239 12 1244 14
rect 1247 13 1258 14
rect 1267 13 1275 14
rect 1277 13 1282 35
rect 1285 33 1297 35
rect 1284 31 1297 33
rect 1285 30 1297 31
rect 1288 18 1293 30
rect 1300 19 1305 35
rect 1312 34 1316 35
rect 1311 19 1317 34
rect 1319 33 1331 35
rect 1337 34 1346 35
rect 1494 34 1499 35
rect 1336 33 1347 34
rect 1319 32 1332 33
rect 1335 32 1348 33
rect 1319 30 1331 32
rect 1335 31 1349 32
rect 1334 30 1349 31
rect 1300 18 1306 19
rect 1310 18 1317 19
rect 1288 17 1294 18
rect 1300 17 1307 18
rect 1309 17 1317 18
rect 1288 16 1297 17
rect 1300 16 1317 17
rect 1322 20 1327 30
rect 1334 29 1339 30
rect 1344 29 1349 30
rect 1333 26 1339 29
rect 1345 27 1350 29
rect 1344 26 1350 27
rect 1333 23 1351 26
rect 1494 24 1498 34
rect 1509 33 1512 35
rect 1524 34 1530 35
rect 1539 34 1542 35
rect 1524 33 1531 34
rect 1333 21 1350 23
rect 1322 18 1328 20
rect 1333 18 1339 21
rect 1494 20 1499 24
rect 1509 20 1511 33
rect 1524 31 1532 33
rect 1495 19 1500 20
rect 1508 19 1510 20
rect 1347 18 1348 19
rect 1495 18 1501 19
rect 1507 18 1510 19
rect 1524 19 1526 31
rect 1527 30 1533 31
rect 1528 29 1534 30
rect 1529 28 1535 29
rect 1530 27 1536 28
rect 1531 26 1537 27
rect 1531 25 1538 26
rect 1532 24 1539 25
rect 1540 24 1542 34
rect 1533 23 1542 24
rect 1534 22 1542 23
rect 1535 21 1542 22
rect 1536 19 1542 21
rect 1524 18 1527 19
rect 1537 18 1542 19
rect 1555 18 1560 35
rect 1573 34 1578 35
rect 1573 33 1579 34
rect 1574 31 1579 33
rect 1587 33 1590 35
rect 1587 31 1589 33
rect 1575 28 1580 31
rect 1586 29 1588 31
rect 1586 28 1587 29
rect 1576 26 1581 28
rect 1585 26 1587 28
rect 1603 28 1608 36
rect 1613 35 1616 36
rect 1628 35 1634 36
rect 1636 35 1642 36
rect 1656 35 1659 36
rect 1664 35 1667 36
rect 1678 35 1684 36
rect 1614 34 1617 35
rect 1628 34 1633 35
rect 1615 32 1617 34
rect 1613 28 1615 30
rect 1603 26 1615 28
rect 1577 23 1582 26
rect 1584 23 1586 26
rect 1578 21 1585 23
rect 1579 18 1584 21
rect 1603 18 1608 26
rect 1613 24 1615 26
rect 1614 23 1615 24
rect 1629 27 1633 34
rect 1638 32 1643 35
rect 1655 34 1659 35
rect 1655 33 1658 34
rect 1665 33 1667 35
rect 1639 30 1643 32
rect 1654 32 1658 33
rect 1666 32 1667 33
rect 1654 31 1659 32
rect 1654 30 1660 31
rect 1638 28 1643 30
rect 1655 29 1661 30
rect 1655 28 1663 29
rect 1637 27 1642 28
rect 1656 27 1665 28
rect 1629 26 1634 27
rect 1635 26 1640 27
rect 1657 26 1666 27
rect 1629 25 1640 26
rect 1658 25 1667 26
rect 1617 21 1618 22
rect 1616 19 1618 21
rect 1629 19 1633 25
rect 1635 24 1640 25
rect 1660 24 1668 25
rect 1636 23 1641 24
rect 1662 23 1668 24
rect 1636 22 1642 23
rect 1663 22 1668 23
rect 1637 21 1642 22
rect 1654 21 1655 22
rect 1637 20 1643 21
rect 1615 18 1618 19
rect 1322 17 1329 18
rect 1334 17 1341 18
rect 1346 17 1349 18
rect 1496 17 1503 18
rect 1505 17 1509 18
rect 1523 17 1527 18
rect 1538 17 1542 18
rect 1554 17 1560 18
rect 1322 16 1332 17
rect 1334 16 1349 17
rect 1497 16 1508 17
rect 1521 16 1530 17
rect 1539 16 1542 17
rect 1552 16 1562 17
rect 1580 16 1583 18
rect 1602 17 1609 18
rect 1614 17 1618 18
rect 1628 18 1633 19
rect 1638 19 1643 20
rect 1654 20 1656 21
rect 1638 18 1644 19
rect 1654 18 1657 20
rect 1664 19 1668 22
rect 1664 18 1667 19
rect 1679 18 1684 35
rect 1695 35 1698 36
rect 1695 34 1697 35
rect 1695 33 1696 34
rect 1694 32 1696 33
rect 1695 31 1696 32
rect 1702 18 1707 36
rect 1710 35 1714 36
rect 1724 35 1730 36
rect 1711 34 1714 35
rect 1712 32 1714 34
rect 1725 33 1730 35
rect 1737 35 1741 36
rect 1737 34 1740 35
rect 1737 33 1739 34
rect 1726 31 1731 33
rect 1736 31 1738 33
rect 1727 30 1732 31
rect 1728 29 1732 30
rect 1735 29 1737 31
rect 1728 28 1733 29
rect 1734 28 1736 29
rect 1729 27 1736 28
rect 1729 26 1735 27
rect 1730 18 1735 26
rect 1628 17 1634 18
rect 1639 17 1645 18
rect 1654 17 1658 18
rect 1663 17 1666 18
rect 1678 17 1684 18
rect 1701 17 1707 18
rect 1729 17 1735 18
rect 1600 16 1617 17
rect 1626 16 1636 17
rect 1640 16 1646 17
rect 1655 16 1665 17
rect 1676 16 1686 17
rect 1699 16 1710 17
rect 1727 16 1738 17
rect 1289 13 1298 16
rect 1301 14 1317 16
rect 1323 14 1332 16
rect 1335 15 1349 16
rect 1498 15 1506 16
rect 1540 15 1542 16
rect 1580 15 1582 16
rect 1643 15 1646 16
rect 1657 15 1663 16
rect 1336 14 1349 15
rect 1302 13 1317 14
rect 1324 13 1332 14
rect 1337 13 1349 14
rect 1248 12 1257 13
rect 1267 12 1274 13
rect 1278 12 1281 13
rect 1290 12 1297 13
rect 1303 12 1310 13
rect 1313 12 1316 13
rect 1325 12 1331 13
rect 1338 12 1348 13
<< metal2 >>
rect 508 505 522 506
rect 728 505 741 506
rect 836 505 846 506
rect 891 505 903 506
rect 503 504 529 505
rect 542 504 577 505
rect 500 503 532 504
rect 498 502 532 503
rect 496 501 532 502
rect 494 500 532 501
rect 492 499 532 500
rect 491 498 532 499
rect 490 497 532 498
rect 488 496 532 497
rect 487 494 532 496
rect 486 493 532 494
rect 485 492 532 493
rect 484 490 532 492
rect 483 489 532 490
rect 482 488 512 489
rect 523 488 532 489
rect 482 487 509 488
rect 526 487 532 488
rect 481 486 507 487
rect 529 486 532 487
rect 481 485 505 486
rect 531 485 532 486
rect 542 503 583 504
rect 542 502 586 503
rect 542 501 588 502
rect 542 500 589 501
rect 542 499 591 500
rect 542 498 592 499
rect 542 496 593 498
rect 542 495 594 496
rect 542 493 595 495
rect 542 491 596 493
rect 480 484 504 485
rect 480 482 503 484
rect 479 481 502 482
rect 479 479 501 481
rect 479 477 500 479
rect 478 475 500 477
rect 478 468 499 475
rect 542 474 562 491
rect 570 490 596 491
rect 572 489 596 490
rect 574 487 597 489
rect 575 485 597 487
rect 576 480 597 485
rect 575 478 597 480
rect 575 477 596 478
rect 574 476 596 477
rect 573 475 596 476
rect 571 474 595 475
rect 542 473 595 474
rect 542 471 594 473
rect 542 470 593 471
rect 542 468 592 470
rect 604 468 625 505
rect 478 464 500 468
rect 542 467 591 468
rect 542 466 589 467
rect 542 465 588 466
rect 542 464 587 465
rect 478 463 501 464
rect 479 462 501 463
rect 542 463 585 464
rect 542 462 583 463
rect 479 461 502 462
rect 542 461 580 462
rect 605 461 625 468
rect 643 465 664 505
rect 723 504 745 505
rect 720 503 746 504
rect 718 502 746 503
rect 716 501 746 502
rect 715 500 746 501
rect 713 499 746 500
rect 712 498 746 499
rect 711 497 746 498
rect 764 497 802 505
rect 832 504 850 505
rect 885 504 907 505
rect 829 503 853 504
rect 882 503 909 504
rect 827 502 854 503
rect 880 502 911 503
rect 826 501 856 502
rect 877 501 913 502
rect 824 500 857 501
rect 876 500 914 501
rect 823 499 858 500
rect 876 499 915 500
rect 822 498 859 499
rect 876 498 916 499
rect 822 497 860 498
rect 710 496 746 497
rect 709 494 746 496
rect 708 493 746 494
rect 707 491 746 493
rect 706 490 731 491
rect 743 490 746 491
rect 705 489 728 490
rect 763 489 802 497
rect 821 496 860 497
rect 876 496 917 498
rect 820 495 861 496
rect 819 494 861 495
rect 876 494 918 496
rect 819 493 862 494
rect 818 492 862 493
rect 818 491 863 492
rect 817 490 838 491
rect 842 490 863 491
rect 876 490 919 494
rect 1652 491 1708 492
rect 1644 490 1711 491
rect 817 489 837 490
rect 843 489 864 490
rect 705 488 726 489
rect 704 487 725 488
rect 704 486 724 487
rect 704 485 723 486
rect 703 484 723 485
rect 703 483 722 484
rect 703 482 721 483
rect 702 480 721 482
rect 729 481 738 482
rect 763 481 779 489
rect 817 488 836 489
rect 816 486 836 488
rect 844 487 864 489
rect 845 486 864 487
rect 876 489 887 490
rect 896 489 919 490
rect 1638 489 1714 490
rect 876 488 883 489
rect 898 488 920 489
rect 1634 488 1716 489
rect 876 487 881 488
rect 876 486 879 487
rect 899 486 920 488
rect 1569 487 1573 488
rect 1629 487 1718 488
rect 1565 486 1579 487
rect 1625 486 1720 487
rect 816 484 835 486
rect 726 480 741 481
rect 762 480 779 481
rect 815 481 835 484
rect 845 483 865 486
rect 876 485 877 486
rect 702 477 720 480
rect 724 479 743 480
rect 762 479 789 480
rect 723 478 744 479
rect 762 478 793 479
rect 722 477 745 478
rect 762 477 795 478
rect 815 477 834 481
rect 701 476 720 477
rect 721 476 746 477
rect 762 476 797 477
rect 701 475 747 476
rect 762 475 798 476
rect 701 473 748 475
rect 762 473 800 475
rect 701 471 749 473
rect 762 472 801 473
rect 762 471 802 472
rect 701 468 750 471
rect 701 467 724 468
rect 729 467 750 468
rect 762 468 803 471
rect 701 466 723 467
rect 730 466 751 467
rect 701 465 722 466
rect 643 461 663 465
rect 479 459 503 461
rect 542 460 575 461
rect 480 458 504 459
rect 480 457 505 458
rect 531 457 532 458
rect 480 456 507 457
rect 529 456 532 457
rect 481 455 509 456
rect 526 455 532 456
rect 481 454 512 455
rect 522 454 532 455
rect 482 452 532 454
rect 483 450 532 452
rect 484 449 532 450
rect 485 448 532 449
rect 486 447 532 448
rect 487 446 532 447
rect 488 445 532 446
rect 489 444 532 445
rect 490 443 532 444
rect 491 442 532 443
rect 493 441 532 442
rect 495 440 532 441
rect 497 439 530 440
rect 501 438 526 439
rect 542 438 562 460
rect 605 458 626 461
rect 642 458 663 461
rect 701 461 721 465
rect 731 464 751 466
rect 762 466 804 468
rect 762 465 764 466
rect 779 465 804 466
rect 814 465 834 477
rect 782 464 805 465
rect 701 459 720 461
rect 605 457 627 458
rect 641 457 663 458
rect 606 456 628 457
rect 640 456 662 457
rect 606 455 629 456
rect 639 455 662 456
rect 702 455 721 459
rect 732 456 751 464
rect 783 463 805 464
rect 784 462 805 463
rect 785 457 805 462
rect 815 461 834 465
rect 846 479 865 483
rect 900 483 920 486
rect 1563 485 1583 486
rect 1621 485 1721 486
rect 1562 484 1586 485
rect 1616 484 1723 485
rect 1560 483 1591 484
rect 1610 483 1724 484
rect 900 481 919 483
rect 1559 482 1726 483
rect 1558 481 1728 482
rect 899 479 919 481
rect 1557 480 1729 481
rect 1557 479 1730 480
rect 846 465 866 479
rect 898 478 919 479
rect 1556 478 1732 479
rect 898 477 918 478
rect 897 476 918 477
rect 1555 477 1733 478
rect 1555 476 1735 477
rect 896 475 917 476
rect 1555 475 1736 476
rect 895 474 917 475
rect 1554 474 1737 475
rect 893 473 916 474
rect 892 472 916 473
rect 1554 473 1738 474
rect 1554 472 1648 473
rect 1666 472 1740 473
rect 891 471 915 472
rect 1554 471 1583 472
rect 1587 471 1645 472
rect 1671 471 1741 472
rect 890 470 914 471
rect 1554 470 1576 471
rect 1594 470 1644 471
rect 1674 470 1742 471
rect 888 469 913 470
rect 1555 469 1573 470
rect 1598 469 1644 470
rect 1678 469 1743 470
rect 887 468 912 469
rect 1555 468 1571 469
rect 1600 468 1646 469
rect 1683 468 1744 469
rect 886 467 911 468
rect 1556 467 1570 468
rect 1602 467 1651 468
rect 1687 467 1745 468
rect 885 466 909 467
rect 1557 466 1568 467
rect 1603 466 1654 467
rect 1692 466 1746 467
rect 884 465 908 466
rect 1534 465 1539 466
rect 1559 465 1564 466
rect 1605 465 1658 466
rect 1699 465 1747 466
rect 846 461 865 465
rect 882 464 907 465
rect 1531 464 1542 465
rect 1606 464 1661 465
rect 1709 464 1748 465
rect 881 463 905 464
rect 1529 463 1545 464
rect 1606 463 1664 464
rect 1715 463 1749 464
rect 880 462 903 463
rect 1527 462 1546 463
rect 1607 462 1667 463
rect 1719 462 1750 463
rect 815 457 835 461
rect 845 458 865 461
rect 879 461 902 462
rect 1526 461 1548 462
rect 1575 461 1583 462
rect 1608 461 1670 462
rect 1723 461 1751 462
rect 879 460 901 461
rect 1525 460 1549 461
rect 1571 460 1586 461
rect 1608 460 1673 461
rect 1727 460 1752 461
rect 878 459 899 460
rect 1524 459 1550 460
rect 1569 459 1588 460
rect 1608 459 1677 460
rect 1730 459 1753 460
rect 877 458 898 459
rect 1523 458 1551 459
rect 1567 458 1590 459
rect 1609 458 1681 459
rect 1734 458 1753 459
rect 845 457 864 458
rect 877 457 897 458
rect 1522 457 1552 458
rect 1565 457 1591 458
rect 1609 457 1687 458
rect 1737 457 1754 458
rect 785 456 804 457
rect 606 454 631 455
rect 637 454 662 455
rect 703 454 722 455
rect 731 454 750 456
rect 784 455 804 456
rect 607 451 661 454
rect 703 453 723 454
rect 730 453 750 454
rect 703 452 724 453
rect 729 452 750 453
rect 760 454 761 455
rect 783 454 804 455
rect 760 453 764 454
rect 782 453 804 454
rect 816 456 835 457
rect 816 454 836 456
rect 844 454 864 457
rect 876 456 896 457
rect 1521 456 1553 457
rect 1563 456 1592 457
rect 1609 456 1704 457
rect 1740 456 1755 457
rect 875 455 895 456
rect 1521 455 1555 456
rect 1561 455 1593 456
rect 1609 455 1709 456
rect 1742 455 1755 456
rect 875 454 894 455
rect 1520 454 1593 455
rect 1608 454 1713 455
rect 1745 454 1756 455
rect 816 453 837 454
rect 843 453 863 454
rect 875 453 920 454
rect 760 452 768 453
rect 779 452 804 453
rect 817 452 838 453
rect 842 452 863 453
rect 608 449 660 451
rect 704 450 749 452
rect 760 450 803 452
rect 817 451 862 452
rect 818 450 862 451
rect 609 448 659 449
rect 705 448 748 450
rect 760 448 802 450
rect 818 449 861 450
rect 874 449 920 453
rect 1519 452 1594 454
rect 1518 451 1594 452
rect 1608 453 1716 454
rect 1748 453 1756 454
rect 1608 452 1719 453
rect 1750 452 1756 453
rect 1608 451 1722 452
rect 1752 451 1757 452
rect 1517 449 1594 451
rect 1607 450 1725 451
rect 1754 450 1757 451
rect 1607 449 1728 450
rect 1756 449 1757 450
rect 819 448 861 449
rect 610 446 658 448
rect 706 447 747 448
rect 760 447 801 448
rect 819 447 860 448
rect 706 446 746 447
rect 611 445 657 446
rect 707 445 746 446
rect 760 445 800 447
rect 820 446 860 447
rect 820 445 859 446
rect 612 444 656 445
rect 708 444 745 445
rect 760 444 799 445
rect 821 444 858 445
rect 613 443 655 444
rect 709 443 744 444
rect 760 443 798 444
rect 822 443 857 444
rect 614 442 654 443
rect 710 442 743 443
rect 760 442 796 443
rect 823 442 856 443
rect 616 441 652 442
rect 711 441 741 442
rect 760 441 795 442
rect 824 441 855 442
rect 618 440 650 441
rect 713 440 740 441
rect 760 440 793 441
rect 826 440 853 441
rect 620 439 648 440
rect 715 439 738 440
rect 760 439 791 440
rect 828 439 852 440
rect 622 438 645 439
rect 717 438 735 439
rect 764 438 788 439
rect 830 438 849 439
rect 873 438 920 449
rect 1516 448 1594 449
rect 1515 447 1594 448
rect 1606 448 1731 449
rect 1606 447 1734 448
rect 1514 446 1594 447
rect 1605 446 1737 447
rect 1513 445 1593 446
rect 1512 444 1593 445
rect 1605 445 1739 446
rect 1605 444 1742 445
rect 1511 443 1592 444
rect 1606 443 1745 444
rect 1510 442 1592 443
rect 1608 442 1747 443
rect 1509 441 1591 442
rect 1610 441 1750 442
rect 1508 440 1590 441
rect 1611 440 1752 441
rect 1507 439 1589 440
rect 1613 439 1666 440
rect 1669 439 1755 440
rect 1506 438 1588 439
rect 1614 438 1666 439
rect 1673 438 1757 439
rect 506 437 520 438
rect 627 437 640 438
rect 721 437 731 438
rect 771 437 784 438
rect 834 437 845 438
rect 1505 437 1587 438
rect 1616 437 1666 438
rect 1675 437 1759 438
rect 1503 436 1585 437
rect 1617 436 1667 437
rect 1678 436 1762 437
rect 1502 435 1542 436
rect 1547 435 1584 436
rect 1619 435 1667 436
rect 1680 435 1763 436
rect 1500 434 1537 435
rect 1546 434 1583 435
rect 1620 434 1667 435
rect 1683 434 1764 435
rect 1499 433 1533 434
rect 1544 433 1582 434
rect 1621 433 1667 434
rect 1685 433 1766 434
rect 1497 432 1530 433
rect 1543 432 1581 433
rect 1623 432 1667 433
rect 1687 432 1766 433
rect 1496 431 1526 432
rect 1541 431 1580 432
rect 1624 431 1668 432
rect 1690 431 1767 432
rect 1494 430 1523 431
rect 1540 430 1579 431
rect 1625 430 1668 431
rect 1692 430 1768 431
rect 1492 429 1521 430
rect 1538 429 1578 430
rect 1626 429 1669 430
rect 1695 429 1769 430
rect 1491 428 1519 429
rect 1536 428 1578 429
rect 1627 428 1669 429
rect 1697 428 1769 429
rect 1489 427 1518 428
rect 1534 427 1577 428
rect 1628 427 1670 428
rect 1701 427 1770 428
rect 1487 426 1516 427
rect 1533 426 1577 427
rect 1629 426 1671 427
rect 1705 426 1770 427
rect 1485 425 1514 426
rect 1531 425 1576 426
rect 1483 424 1512 425
rect 1530 424 1576 425
rect 1592 425 1595 426
rect 1602 425 1605 426
rect 1630 425 1672 426
rect 1711 425 1771 426
rect 1592 424 1610 425
rect 1631 424 1673 425
rect 1715 424 1771 425
rect 1481 423 1511 424
rect 1478 422 1510 423
rect 1529 422 1576 424
rect 1593 423 1613 424
rect 1632 423 1674 424
rect 1718 423 1772 424
rect 1593 422 1614 423
rect 1633 422 1676 423
rect 1720 422 1772 423
rect 1476 421 1509 422
rect 1516 421 1518 422
rect 1528 421 1577 422
rect 1475 420 1509 421
rect 1511 420 1518 421
rect 1527 420 1577 421
rect 1473 419 1518 420
rect 1471 418 1518 419
rect 1526 418 1577 420
rect 1594 421 1616 422
rect 1634 421 1677 422
rect 1723 421 1773 422
rect 1594 420 1617 421
rect 1635 420 1679 421
rect 1725 420 1773 421
rect 1594 419 1618 420
rect 1635 419 1681 420
rect 1727 419 1773 420
rect 1470 417 1519 418
rect 1468 416 1519 417
rect 1525 417 1577 418
rect 1595 417 1619 419
rect 1636 418 1683 419
rect 1729 418 1774 419
rect 1637 417 1685 418
rect 1731 417 1774 418
rect 1525 416 1578 417
rect 1467 415 1519 416
rect 1466 414 1520 415
rect 1524 414 1578 416
rect 1465 413 1521 414
rect 1523 413 1578 414
rect 1596 416 1620 417
rect 1638 416 1687 417
rect 1733 416 1774 417
rect 1596 414 1621 416
rect 1638 415 1690 416
rect 1734 415 1774 416
rect 1639 414 1694 415
rect 1736 414 1775 415
rect 1596 413 1622 414
rect 1640 413 1697 414
rect 1738 413 1775 414
rect 1464 412 1579 413
rect 1463 411 1579 412
rect 1462 409 1579 411
rect 1461 407 1579 409
rect 1597 411 1623 413
rect 1640 412 1701 413
rect 1739 412 1775 413
rect 1641 411 1705 412
rect 1741 411 1775 412
rect 1597 409 1624 411
rect 1642 410 1710 411
rect 1742 410 1776 411
rect 1642 409 1714 410
rect 1744 409 1776 410
rect 1597 407 1625 409
rect 1643 408 1717 409
rect 1745 408 1776 409
rect 1643 407 1719 408
rect 1746 407 1776 408
rect 1461 405 1580 407
rect 1461 404 1481 405
rect 1482 404 1580 405
rect 502 401 509 402
rect 524 401 531 402
rect 545 401 552 402
rect 499 400 511 401
rect 522 400 533 401
rect 542 400 554 401
rect 571 400 577 402
rect 498 399 512 400
rect 521 399 534 400
rect 498 398 513 399
rect 498 397 503 398
rect 505 397 513 398
rect 520 398 534 399
rect 541 399 555 400
rect 541 398 556 399
rect 570 398 577 400
rect 520 397 526 398
rect 528 397 535 398
rect 498 396 500 397
rect 507 396 513 397
rect 519 396 525 397
rect 529 396 535 397
rect 541 397 546 398
rect 548 397 556 398
rect 569 397 577 398
rect 541 396 543 397
rect 550 396 556 397
rect 508 393 514 396
rect 519 395 524 396
rect 508 392 513 393
rect 507 391 513 392
rect 506 390 513 391
rect 518 392 524 395
rect 530 393 536 396
rect 505 389 512 390
rect 504 388 511 389
rect 503 387 510 388
rect 501 386 509 387
rect 518 386 523 392
rect 500 385 508 386
rect 499 384 506 385
rect 498 383 505 384
rect 518 383 524 386
rect 531 385 536 393
rect 551 393 557 396
rect 568 395 577 397
rect 567 394 577 395
rect 566 393 571 394
rect 551 392 556 393
rect 566 392 570 393
rect 550 391 556 392
rect 565 391 570 392
rect 549 390 556 391
rect 564 390 569 391
rect 548 389 555 390
rect 564 389 568 390
rect 547 388 554 389
rect 563 388 568 389
rect 546 387 553 388
rect 562 387 567 388
rect 544 386 552 387
rect 561 386 566 387
rect 572 386 577 394
rect 543 385 551 386
rect 560 385 566 386
rect 571 385 577 386
rect 498 382 504 383
rect 519 382 524 383
rect 530 382 536 385
rect 542 384 549 385
rect 541 383 548 384
rect 541 382 547 383
rect 497 381 503 382
rect 519 381 525 382
rect 529 381 535 382
rect 497 376 514 381
rect 519 380 526 381
rect 528 380 535 381
rect 540 381 546 382
rect 560 381 580 385
rect 609 383 615 402
rect 689 401 694 402
rect 713 401 718 402
rect 738 401 747 402
rect 689 400 693 401
rect 714 400 719 401
rect 735 400 749 401
rect 688 399 693 400
rect 687 397 692 399
rect 715 398 720 400
rect 733 399 749 400
rect 732 398 749 399
rect 686 395 691 397
rect 716 396 721 398
rect 731 397 749 398
rect 730 396 739 397
rect 747 396 749 397
rect 624 394 631 395
rect 621 393 633 394
rect 621 392 634 393
rect 641 392 646 395
rect 650 394 655 395
rect 648 393 656 394
rect 647 392 657 393
rect 685 392 690 395
rect 703 394 710 395
rect 717 394 722 396
rect 730 395 737 396
rect 701 393 711 394
rect 699 392 711 393
rect 621 391 635 392
rect 621 390 624 391
rect 630 390 635 391
rect 641 391 658 392
rect 685 391 689 392
rect 698 391 711 392
rect 641 390 649 391
rect 650 390 658 391
rect 621 389 622 390
rect 630 388 636 390
rect 625 387 636 388
rect 622 386 636 387
rect 621 385 636 386
rect 620 384 626 385
rect 619 383 625 384
rect 631 383 636 385
rect 608 382 614 383
rect 602 381 603 382
rect 607 381 614 382
rect 520 379 534 380
rect 521 378 533 379
rect 522 377 532 378
rect 524 376 530 377
rect 540 376 557 381
rect 572 376 577 381
rect 602 380 614 381
rect 619 381 624 383
rect 630 381 636 383
rect 619 380 625 381
rect 629 380 636 381
rect 583 379 589 380
rect 602 379 613 380
rect 619 379 636 380
rect 583 376 588 379
rect 602 378 612 379
rect 620 378 636 379
rect 602 377 611 378
rect 621 377 629 378
rect 602 376 609 377
rect 622 376 627 377
rect 631 376 636 378
rect 641 389 647 390
rect 641 376 646 389
rect 652 388 658 390
rect 653 376 658 388
rect 664 381 667 382
rect 663 380 668 381
rect 684 380 689 391
rect 697 390 706 391
rect 708 390 711 391
rect 718 393 722 394
rect 729 394 736 395
rect 761 394 768 395
rect 783 394 791 395
rect 806 394 811 395
rect 729 393 735 394
rect 758 393 770 394
rect 781 393 793 394
rect 804 393 813 394
rect 814 393 819 404
rect 697 388 703 390
rect 718 389 723 393
rect 696 382 702 388
rect 719 383 723 389
rect 728 392 735 393
rect 757 392 772 393
rect 780 392 794 393
rect 803 392 819 393
rect 728 386 734 392
rect 756 391 772 392
rect 779 391 795 392
rect 802 391 819 392
rect 740 386 751 391
rect 756 390 763 391
rect 766 390 773 391
rect 778 390 786 391
rect 788 390 796 391
rect 755 388 761 390
rect 767 389 774 390
rect 778 389 784 390
rect 790 389 796 390
rect 801 390 809 391
rect 811 390 819 391
rect 801 389 807 390
rect 755 387 760 388
rect 768 387 774 389
rect 728 384 735 386
rect 697 381 703 382
rect 697 380 705 381
rect 708 380 711 381
rect 662 378 669 380
rect 663 377 668 378
rect 685 377 690 380
rect 698 379 711 380
rect 699 378 711 379
rect 718 378 723 383
rect 729 383 736 384
rect 729 382 737 383
rect 730 381 738 382
rect 745 381 751 386
rect 754 384 760 387
rect 769 384 774 387
rect 755 383 760 384
rect 755 381 761 383
rect 768 382 774 384
rect 777 382 783 389
rect 791 383 797 389
rect 791 382 796 383
rect 800 382 806 389
rect 813 388 819 390
rect 814 384 819 388
rect 813 382 819 384
rect 767 381 773 382
rect 730 380 751 381
rect 731 379 751 380
rect 756 380 763 381
rect 766 380 773 381
rect 778 381 784 382
rect 790 381 796 382
rect 778 380 786 381
rect 788 380 796 381
rect 801 381 807 382
rect 812 381 819 382
rect 801 380 809 381
rect 811 380 819 381
rect 756 379 772 380
rect 779 379 795 380
rect 801 379 819 380
rect 733 378 751 379
rect 757 378 771 379
rect 780 378 794 379
rect 802 378 819 379
rect 700 377 711 378
rect 664 376 667 377
rect 583 375 587 376
rect 686 375 691 377
rect 702 376 710 377
rect 717 376 722 378
rect 734 377 749 378
rect 758 377 770 378
rect 781 377 793 378
rect 803 377 812 378
rect 737 376 746 377
rect 761 376 768 377
rect 783 376 791 377
rect 805 376 810 377
rect 814 376 819 378
rect 825 391 830 402
rect 838 401 845 402
rect 838 400 844 401
rect 837 399 844 400
rect 836 398 843 399
rect 836 397 842 398
rect 835 396 841 397
rect 834 395 841 396
rect 834 394 840 395
rect 854 394 861 395
rect 876 394 884 395
rect 833 393 839 394
rect 851 393 863 394
rect 874 393 886 394
rect 832 392 839 393
rect 850 392 865 393
rect 873 392 887 393
rect 832 391 838 392
rect 849 391 865 392
rect 872 391 888 392
rect 825 388 837 391
rect 849 390 856 391
rect 859 390 866 391
rect 871 390 879 391
rect 881 390 889 391
rect 848 388 854 390
rect 860 389 867 390
rect 871 389 877 390
rect 883 389 889 390
rect 825 376 830 388
rect 831 387 838 388
rect 848 387 853 388
rect 861 387 867 389
rect 832 386 839 387
rect 833 385 839 386
rect 833 384 840 385
rect 847 384 853 387
rect 862 384 867 387
rect 834 383 841 384
rect 848 383 853 384
rect 835 381 842 383
rect 848 381 854 383
rect 861 382 867 384
rect 870 382 876 389
rect 884 383 890 389
rect 894 387 900 404
rect 1461 403 1479 404
rect 1481 403 1580 404
rect 1462 402 1477 403
rect 1480 402 1580 403
rect 1462 401 1475 402
rect 1479 401 1580 402
rect 1463 400 1472 401
rect 1478 400 1580 401
rect 1465 399 1468 400
rect 1477 399 1580 400
rect 1476 398 1580 399
rect 1475 397 1580 398
rect 1597 405 1626 407
rect 1644 406 1721 407
rect 1748 406 1776 407
rect 1644 405 1723 406
rect 1749 405 1776 406
rect 1597 402 1627 405
rect 1645 404 1724 405
rect 1750 404 1776 405
rect 1645 403 1726 404
rect 1751 403 1777 404
rect 1645 402 1728 403
rect 1753 402 1777 403
rect 1597 400 1628 402
rect 1646 401 1729 402
rect 1754 401 1777 402
rect 1646 400 1731 401
rect 1755 400 1777 401
rect 1597 398 1629 400
rect 1647 399 1732 400
rect 1756 399 1777 400
rect 1647 398 1733 399
rect 1757 398 1777 399
rect 1474 396 1579 397
rect 1597 396 1630 398
rect 1648 397 1735 398
rect 1758 397 1777 398
rect 1649 396 1736 397
rect 1759 396 1777 397
rect 1473 395 1579 396
rect 905 394 912 395
rect 1472 394 1579 395
rect 905 393 911 394
rect 1471 393 1579 394
rect 1596 394 1631 396
rect 1649 395 1737 396
rect 1760 395 1777 396
rect 1650 394 1739 395
rect 1761 394 1777 395
rect 904 392 910 393
rect 903 391 910 392
rect 1470 391 1578 393
rect 1596 392 1632 394
rect 1651 393 1740 394
rect 1762 393 1777 394
rect 1652 392 1741 393
rect 1596 391 1633 392
rect 1653 391 1742 392
rect 1763 391 1777 393
rect 903 390 909 391
rect 1469 390 1578 391
rect 902 389 908 390
rect 901 387 907 389
rect 1469 388 1577 390
rect 1595 389 1634 391
rect 1654 390 1744 391
rect 1764 390 1777 391
rect 1656 389 1745 390
rect 1765 389 1777 390
rect 1595 388 1635 389
rect 1658 388 1746 389
rect 1468 387 1576 388
rect 894 385 906 387
rect 1469 386 1576 387
rect 1594 386 1636 388
rect 1660 387 1747 388
rect 1766 387 1776 389
rect 1662 386 1748 387
rect 1767 386 1776 387
rect 1469 385 1575 386
rect 1594 385 1637 386
rect 1666 385 1749 386
rect 894 384 907 385
rect 1469 384 1574 385
rect 1594 384 1638 385
rect 1671 384 1750 385
rect 1768 384 1776 386
rect 884 382 889 383
rect 860 381 866 382
rect 836 380 843 381
rect 849 380 856 381
rect 859 380 866 381
rect 871 381 877 382
rect 883 381 889 382
rect 871 380 879 381
rect 881 380 889 381
rect 837 378 844 380
rect 849 379 865 380
rect 872 379 888 380
rect 850 378 864 379
rect 873 378 887 379
rect 838 377 845 378
rect 851 377 863 378
rect 874 377 886 378
rect 839 376 846 377
rect 854 376 861 377
rect 876 376 884 377
rect 894 376 900 384
rect 901 383 907 384
rect 1470 383 1574 384
rect 1593 383 1639 384
rect 1677 383 1751 384
rect 1769 383 1776 384
rect 902 382 908 383
rect 1470 382 1573 383
rect 1593 382 1641 383
rect 1683 382 1752 383
rect 902 381 909 382
rect 903 380 910 381
rect 1471 380 1572 382
rect 1592 381 1642 382
rect 1688 381 1753 382
rect 1770 381 1775 383
rect 1592 380 1644 381
rect 1691 380 1754 381
rect 1771 380 1775 381
rect 904 379 910 380
rect 1472 379 1571 380
rect 1592 379 1645 380
rect 1694 379 1755 380
rect 1771 379 1774 380
rect 904 378 911 379
rect 1472 378 1517 379
rect 1519 378 1570 379
rect 905 377 912 378
rect 1473 377 1515 378
rect 1521 377 1570 378
rect 1591 378 1647 379
rect 1697 378 1755 379
rect 1772 378 1774 379
rect 1591 377 1650 378
rect 1700 377 1756 378
rect 1772 377 1773 378
rect 906 376 912 377
rect 1474 376 1514 377
rect 1522 376 1569 377
rect 1590 376 1653 377
rect 1702 376 1757 377
rect 582 373 587 375
rect 687 374 691 375
rect 716 374 721 376
rect 1475 375 1513 376
rect 1523 375 1568 376
rect 1590 375 1657 376
rect 1705 375 1757 376
rect 1476 374 1512 375
rect 1523 374 1567 375
rect 1590 374 1662 375
rect 1707 374 1757 375
rect 687 373 692 374
rect 582 371 586 373
rect 688 371 693 373
rect 715 372 720 374
rect 1477 373 1511 374
rect 1524 373 1567 374
rect 1589 373 1667 374
rect 1710 373 1758 374
rect 1478 372 1508 373
rect 1524 372 1566 373
rect 1589 372 1673 373
rect 1713 372 1758 373
rect 714 371 719 372
rect 1479 371 1504 372
rect 1523 371 1566 372
rect 1588 371 1677 372
rect 1715 371 1758 372
rect 689 370 694 371
rect 713 370 718 371
rect 1481 370 1496 371
rect 1523 370 1565 371
rect 1588 370 1681 371
rect 1717 370 1759 371
rect 1486 369 1487 370
rect 1521 369 1564 370
rect 1518 368 1564 369
rect 1587 369 1683 370
rect 1718 369 1759 370
rect 1587 368 1686 369
rect 1720 368 1759 369
rect 1515 367 1563 368
rect 1586 367 1689 368
rect 1721 367 1759 368
rect 1511 366 1563 367
rect 1585 366 1691 367
rect 1722 366 1759 367
rect 1505 365 1562 366
rect 1585 365 1693 366
rect 1723 365 1760 366
rect 1496 364 1561 365
rect 1486 363 1561 364
rect 1584 364 1695 365
rect 1724 364 1760 365
rect 1584 363 1697 364
rect 1725 363 1760 364
rect 1484 362 1560 363
rect 1583 362 1699 363
rect 1726 362 1760 363
rect 1484 361 1559 362
rect 1483 360 1559 361
rect 1582 361 1701 362
rect 1727 361 1760 362
rect 1582 360 1702 361
rect 1728 360 1760 361
rect 1483 359 1558 360
rect 1581 359 1704 360
rect 1483 358 1557 359
rect 1580 358 1705 359
rect 1729 358 1760 360
rect 1483 357 1556 358
rect 1579 357 1706 358
rect 1730 357 1760 358
rect 1483 356 1555 357
rect 1579 356 1707 357
rect 1731 356 1760 357
rect 1483 355 1554 356
rect 1578 355 1708 356
rect 1484 354 1553 355
rect 1577 354 1709 355
rect 1732 354 1760 356
rect 1484 353 1552 354
rect 1576 353 1710 354
rect 1484 352 1551 353
rect 1575 352 1711 353
rect 1733 352 1760 354
rect 1485 351 1550 352
rect 1574 351 1712 352
rect 1734 351 1760 352
rect 473 350 694 351
rect 734 350 960 351
rect 996 350 1204 351
rect 1285 350 1352 351
rect 1485 350 1548 351
rect 1574 350 1713 351
rect 472 315 695 350
rect 734 349 961 350
rect 995 349 1210 350
rect 1285 349 1353 350
rect 733 315 962 349
rect 995 348 1213 349
rect 994 347 1215 348
rect 995 346 1217 347
rect 995 345 1219 346
rect 995 344 1220 345
rect 995 343 1222 344
rect 995 342 1223 343
rect 995 341 1224 342
rect 995 340 1225 341
rect 995 339 1226 340
rect 995 337 1227 339
rect 995 336 1228 337
rect 995 334 1229 336
rect 995 332 1230 334
rect 995 330 1231 332
rect 995 327 1232 330
rect 995 321 1233 327
rect 472 314 694 315
rect 734 314 961 315
rect 995 314 1234 321
rect 472 313 542 314
rect 813 313 883 314
rect 472 285 541 313
rect 472 284 542 285
rect 472 283 693 284
rect 472 282 694 283
rect 472 248 695 282
rect 472 247 694 248
rect 472 246 543 247
rect 545 246 547 247
rect 691 246 692 247
rect 472 245 542 246
rect 472 217 541 245
rect 472 216 542 217
rect 472 215 694 216
rect 472 207 695 215
rect 473 203 695 207
rect 474 200 695 203
rect 475 198 695 200
rect 476 196 695 198
rect 477 194 695 196
rect 478 193 695 194
rect 479 192 695 193
rect 480 190 695 192
rect 481 189 695 190
rect 482 188 695 189
rect 483 187 695 188
rect 484 186 695 187
rect 486 185 695 186
rect 487 184 695 185
rect 489 183 695 184
rect 491 182 695 183
rect 494 181 695 182
rect 496 180 695 181
rect 813 180 882 313
rect 995 183 1064 314
rect 1165 260 1234 314
rect 1087 259 1089 260
rect 1091 259 1161 260
rect 1162 259 1233 260
rect 1086 258 1168 259
rect 1087 257 1168 258
rect 1088 256 1168 257
rect 1089 255 1170 256
rect 1090 254 1171 255
rect 1091 253 1172 254
rect 1092 252 1172 253
rect 1093 251 1174 252
rect 1094 250 1175 251
rect 1095 249 1176 250
rect 1096 248 1177 249
rect 1097 247 1178 248
rect 1098 246 1179 247
rect 1099 245 1180 246
rect 1100 244 1181 245
rect 1101 243 1182 244
rect 1102 242 1183 243
rect 1103 241 1184 242
rect 1104 240 1185 241
rect 1105 239 1186 240
rect 1106 238 1187 239
rect 1107 237 1188 238
rect 1108 236 1189 237
rect 1109 235 1190 236
rect 1110 234 1191 235
rect 1111 233 1192 234
rect 1112 232 1193 233
rect 1113 231 1194 232
rect 1114 230 1195 231
rect 1115 229 1196 230
rect 1116 228 1197 229
rect 1117 227 1198 228
rect 1118 226 1199 227
rect 1119 225 1200 226
rect 1120 224 1201 225
rect 1121 223 1202 224
rect 1122 222 1203 223
rect 1123 221 1204 222
rect 1124 220 1205 221
rect 1125 219 1206 220
rect 1126 218 1207 219
rect 1127 217 1208 218
rect 1128 216 1209 217
rect 1129 215 1210 216
rect 1130 214 1211 215
rect 1131 213 1212 214
rect 1132 212 1213 213
rect 1133 211 1214 212
rect 1134 210 1215 211
rect 1135 209 1216 210
rect 1136 208 1217 209
rect 1137 207 1218 208
rect 1138 206 1219 207
rect 1139 205 1220 206
rect 1140 204 1221 205
rect 1141 203 1222 204
rect 1142 202 1223 203
rect 1143 201 1225 202
rect 1144 200 1225 201
rect 1145 199 1227 200
rect 1146 198 1227 199
rect 1147 197 1229 198
rect 1148 196 1229 197
rect 1149 195 1231 196
rect 1150 194 1231 195
rect 1151 193 1233 194
rect 1152 192 1233 193
rect 1153 191 1235 192
rect 1154 190 1235 191
rect 1155 189 1237 190
rect 1156 188 1237 189
rect 1157 187 1239 188
rect 1158 186 1239 187
rect 1159 185 1241 186
rect 1160 184 1241 185
rect 1161 183 1243 184
rect 994 181 1064 183
rect 1162 182 1243 183
rect 1163 181 1245 182
rect 1284 181 1353 349
rect 1486 349 1547 350
rect 1573 349 1633 350
rect 1642 349 1713 350
rect 1735 349 1760 351
rect 1486 348 1545 349
rect 1572 348 1631 349
rect 1646 348 1714 349
rect 1487 347 1543 348
rect 1570 347 1630 348
rect 1648 347 1715 348
rect 1736 347 1760 349
rect 1488 346 1541 347
rect 1569 346 1629 347
rect 1650 346 1715 347
rect 1488 345 1539 346
rect 1568 345 1628 346
rect 1652 345 1716 346
rect 1737 345 1760 347
rect 1489 344 1537 345
rect 1567 344 1627 345
rect 1653 344 1716 345
rect 1738 344 1760 345
rect 1490 343 1535 344
rect 1566 343 1627 344
rect 1655 343 1717 344
rect 1738 343 1759 344
rect 1490 342 1532 343
rect 1564 342 1626 343
rect 1656 342 1717 343
rect 1491 341 1529 342
rect 1563 341 1626 342
rect 1657 341 1718 342
rect 1739 341 1759 343
rect 1491 340 1526 341
rect 1562 340 1625 341
rect 1658 340 1718 341
rect 1492 339 1524 340
rect 1560 339 1625 340
rect 1659 339 1718 340
rect 1492 338 1520 339
rect 1558 338 1625 339
rect 1660 338 1719 339
rect 1740 338 1759 341
rect 1492 337 1517 338
rect 1557 337 1624 338
rect 1661 337 1719 338
rect 1493 336 1514 337
rect 1555 336 1624 337
rect 1662 336 1719 337
rect 1741 336 1758 338
rect 1493 335 1511 336
rect 1553 335 1624 336
rect 1663 335 1719 336
rect 1494 334 1508 335
rect 1551 334 1623 335
rect 1664 334 1719 335
rect 1494 333 1505 334
rect 1549 333 1623 334
rect 1665 333 1719 334
rect 1742 334 1758 336
rect 1742 333 1757 334
rect 1495 332 1502 333
rect 1547 332 1623 333
rect 1640 332 1642 333
rect 1665 332 1720 333
rect 1545 331 1622 332
rect 1640 331 1643 332
rect 1542 330 1622 331
rect 1540 329 1622 330
rect 1639 330 1644 331
rect 1666 330 1720 332
rect 1743 331 1757 333
rect 1743 330 1756 331
rect 1538 328 1621 329
rect 1639 328 1645 330
rect 1667 328 1719 330
rect 1535 327 1621 328
rect 1638 327 1646 328
rect 1533 326 1620 327
rect 1638 326 1647 327
rect 1668 326 1719 328
rect 1744 328 1756 330
rect 1744 327 1755 328
rect 1531 325 1620 326
rect 1637 325 1647 326
rect 1528 324 1619 325
rect 1637 324 1648 325
rect 1669 324 1719 326
rect 1745 326 1755 327
rect 1745 324 1754 326
rect 1526 323 1619 324
rect 1524 322 1618 323
rect 1636 322 1649 324
rect 1522 321 1618 322
rect 1520 320 1617 321
rect 1635 320 1650 322
rect 1670 321 1718 324
rect 1746 322 1753 324
rect 1518 319 1617 320
rect 1634 319 1651 320
rect 1671 319 1717 321
rect 1746 320 1752 322
rect 1747 319 1751 320
rect 1517 318 1616 319
rect 1634 318 1652 319
rect 1515 317 1616 318
rect 1514 316 1615 317
rect 1633 316 1652 318
rect 1671 317 1716 319
rect 1747 318 1750 319
rect 1747 317 1749 318
rect 1672 316 1715 317
rect 1747 316 1748 317
rect 1512 315 1615 316
rect 1511 314 1614 315
rect 1632 314 1653 316
rect 1672 314 1714 316
rect 1510 313 1613 314
rect 1509 312 1613 313
rect 1631 312 1654 314
rect 1672 313 1713 314
rect 1508 311 1612 312
rect 1630 311 1654 312
rect 1673 312 1712 313
rect 1507 310 1611 311
rect 1506 309 1610 310
rect 1630 309 1655 311
rect 1673 310 1711 312
rect 1673 309 1710 310
rect 1505 308 1609 309
rect 1504 307 1609 308
rect 1629 308 1655 309
rect 1674 308 1709 309
rect 1629 307 1656 308
rect 1504 306 1608 307
rect 1503 305 1607 306
rect 1628 305 1656 307
rect 1502 304 1606 305
rect 1627 304 1656 305
rect 1674 307 1708 308
rect 1674 306 1707 307
rect 1674 305 1706 306
rect 1674 304 1705 305
rect 1732 304 1733 305
rect 1502 303 1605 304
rect 1627 303 1657 304
rect 1501 302 1604 303
rect 1626 302 1657 303
rect 1674 303 1704 304
rect 1731 303 1733 304
rect 1674 302 1702 303
rect 1730 302 1733 303
rect 1501 301 1603 302
rect 1500 300 1602 301
rect 1625 300 1657 302
rect 1500 299 1601 300
rect 1624 299 1657 300
rect 1675 301 1701 302
rect 1729 301 1734 302
rect 1675 300 1700 301
rect 1728 300 1734 301
rect 1675 299 1698 300
rect 1727 299 1734 300
rect 1499 298 1600 299
rect 1499 297 1599 298
rect 1623 297 1658 299
rect 1498 296 1598 297
rect 1622 296 1658 297
rect 1498 295 1597 296
rect 1621 295 1658 296
rect 1497 294 1596 295
rect 1497 293 1595 294
rect 1620 293 1658 295
rect 1675 298 1697 299
rect 1726 298 1734 299
rect 1675 297 1695 298
rect 1725 297 1734 298
rect 1675 296 1694 297
rect 1724 296 1734 297
rect 1675 295 1692 296
rect 1723 295 1734 296
rect 1675 294 1690 295
rect 1722 294 1735 295
rect 1675 293 1689 294
rect 1721 293 1735 294
rect 1497 292 1593 293
rect 1619 292 1658 293
rect 1497 291 1592 292
rect 1618 291 1658 292
rect 1496 290 1591 291
rect 1617 290 1658 291
rect 1496 289 1589 290
rect 1616 289 1658 290
rect 1496 288 1588 289
rect 1615 288 1658 289
rect 1496 287 1586 288
rect 1614 287 1658 288
rect 1674 292 1687 293
rect 1720 292 1735 293
rect 1674 291 1685 292
rect 1718 291 1735 292
rect 1674 290 1683 291
rect 1717 290 1735 291
rect 1674 289 1680 290
rect 1716 289 1735 290
rect 1674 288 1678 289
rect 1715 288 1735 289
rect 1674 287 1675 288
rect 1713 287 1735 288
rect 1496 286 1585 287
rect 1613 286 1658 287
rect 1712 286 1735 287
rect 1495 285 1583 286
rect 1612 285 1658 286
rect 1710 285 1735 286
rect 1495 284 1581 285
rect 1610 284 1658 285
rect 1709 284 1735 285
rect 1495 283 1579 284
rect 1609 283 1658 284
rect 1707 283 1735 284
rect 1495 282 1577 283
rect 1608 282 1658 283
rect 1706 282 1735 283
rect 1495 281 1576 282
rect 1607 281 1658 282
rect 1704 281 1735 282
rect 1495 280 1573 281
rect 1605 280 1658 281
rect 1703 280 1735 281
rect 1495 279 1571 280
rect 1604 279 1657 280
rect 1701 279 1735 280
rect 1495 278 1569 279
rect 1602 278 1657 279
rect 1699 278 1735 279
rect 1495 277 1567 278
rect 1601 277 1657 278
rect 1697 277 1735 278
rect 1495 276 1565 277
rect 1599 276 1657 277
rect 1696 276 1735 277
rect 1495 275 1562 276
rect 1597 275 1657 276
rect 1694 275 1735 276
rect 1495 274 1560 275
rect 1596 274 1657 275
rect 1692 274 1734 275
rect 1495 273 1558 274
rect 1594 273 1656 274
rect 1690 273 1734 274
rect 1495 272 1555 273
rect 1592 272 1656 273
rect 1687 272 1734 273
rect 1495 271 1553 272
rect 1590 271 1656 272
rect 1685 271 1734 272
rect 1495 270 1551 271
rect 1588 270 1656 271
rect 1683 270 1734 271
rect 1495 269 1549 270
rect 1586 269 1655 270
rect 1680 269 1734 270
rect 1496 268 1547 269
rect 1584 268 1655 269
rect 1678 268 1734 269
rect 1496 267 1546 268
rect 1583 267 1655 268
rect 1675 267 1733 268
rect 1496 266 1544 267
rect 1581 266 1655 267
rect 1672 266 1733 267
rect 1496 265 1543 266
rect 1579 265 1654 266
rect 1669 265 1733 266
rect 1496 264 1542 265
rect 1577 264 1654 265
rect 1665 264 1733 265
rect 1496 263 1540 264
rect 1575 263 1654 264
rect 1661 263 1732 264
rect 1497 262 1539 263
rect 1573 262 1732 263
rect 1497 261 1538 262
rect 1571 261 1732 262
rect 1497 260 1537 261
rect 1570 260 1732 261
rect 1497 259 1536 260
rect 1568 259 1731 260
rect 1498 257 1535 259
rect 1566 258 1731 259
rect 1565 257 1731 258
rect 1498 256 1534 257
rect 1563 256 1730 257
rect 1499 254 1533 256
rect 1562 255 1730 256
rect 1560 254 1730 255
rect 1499 253 1532 254
rect 1559 253 1729 254
rect 1500 252 1532 253
rect 1558 252 1729 253
rect 1500 251 1531 252
rect 1556 251 1728 252
rect 1501 250 1531 251
rect 1555 250 1728 251
rect 1501 248 1530 250
rect 1554 249 1728 250
rect 1553 248 1727 249
rect 1502 246 1529 248
rect 1552 247 1618 248
rect 1619 247 1727 248
rect 1551 246 1616 247
rect 1503 245 1529 246
rect 1550 245 1615 246
rect 1619 245 1726 247
rect 1503 244 1528 245
rect 1549 244 1613 245
rect 1619 244 1725 245
rect 1504 242 1528 244
rect 1548 243 1611 244
rect 1618 243 1725 244
rect 1548 242 1610 243
rect 1618 242 1724 243
rect 1505 241 1528 242
rect 1547 241 1608 242
rect 1617 241 1724 242
rect 1505 240 1527 241
rect 1546 240 1607 241
rect 1617 240 1723 241
rect 1506 239 1527 240
rect 1507 237 1527 239
rect 1545 239 1605 240
rect 1545 238 1603 239
rect 1616 238 1722 240
rect 1544 237 1602 238
rect 1615 237 1721 238
rect 1508 235 1526 237
rect 1543 236 1600 237
rect 1614 236 1721 237
rect 1543 235 1599 236
rect 1614 235 1720 236
rect 1509 234 1526 235
rect 1510 232 1526 234
rect 1542 234 1597 235
rect 1613 234 1719 235
rect 1542 233 1596 234
rect 1612 233 1719 234
rect 1511 231 1526 232
rect 1541 232 1594 233
rect 1612 232 1718 233
rect 1541 231 1593 232
rect 1611 231 1717 232
rect 1512 230 1526 231
rect 1513 229 1526 230
rect 1540 230 1592 231
rect 1610 230 1659 231
rect 1660 230 1717 231
rect 1540 229 1591 230
rect 1609 229 1658 230
rect 1659 229 1716 230
rect 1514 227 1525 229
rect 1515 226 1525 227
rect 1539 228 1589 229
rect 1609 228 1656 229
rect 1659 228 1715 229
rect 1539 227 1588 228
rect 1608 227 1655 228
rect 1539 226 1587 227
rect 1607 226 1653 227
rect 1658 226 1714 228
rect 1516 225 1525 226
rect 1517 224 1525 225
rect 1518 223 1525 224
rect 1538 225 1586 226
rect 1606 225 1652 226
rect 1657 225 1713 226
rect 1538 224 1585 225
rect 1606 224 1651 225
rect 1657 224 1712 225
rect 1538 223 1584 224
rect 1605 223 1650 224
rect 1656 223 1711 224
rect 1519 222 1525 223
rect 1520 221 1525 222
rect 1521 220 1525 221
rect 1522 219 1525 220
rect 1537 222 1583 223
rect 1604 222 1648 223
rect 1656 222 1710 223
rect 1537 220 1582 222
rect 1603 221 1647 222
rect 1655 221 1709 222
rect 1603 220 1646 221
rect 1537 219 1581 220
rect 1602 219 1645 220
rect 1655 219 1708 221
rect 1523 218 1525 219
rect 1524 217 1525 218
rect 1536 218 1580 219
rect 1601 218 1644 219
rect 1654 218 1707 219
rect 1536 217 1579 218
rect 1601 217 1643 218
rect 1654 217 1706 218
rect 1536 215 1578 217
rect 1600 216 1642 217
rect 1654 216 1705 217
rect 1600 215 1641 216
rect 1654 215 1704 216
rect 1536 214 1577 215
rect 1599 214 1641 215
rect 1653 214 1703 215
rect 1535 212 1576 214
rect 1599 213 1640 214
rect 1653 213 1702 214
rect 1598 212 1639 213
rect 1653 212 1701 213
rect 1535 210 1575 212
rect 1598 211 1638 212
rect 1597 210 1638 211
rect 1653 211 1700 212
rect 1653 210 1699 211
rect 1535 208 1574 210
rect 1597 209 1637 210
rect 1652 209 1697 210
rect 1597 208 1636 209
rect 1535 205 1573 208
rect 1596 207 1636 208
rect 1652 208 1696 209
rect 1652 207 1695 208
rect 1596 206 1635 207
rect 1595 205 1635 206
rect 1652 206 1694 207
rect 1652 205 1693 206
rect 1535 204 1572 205
rect 1536 202 1572 204
rect 1595 204 1634 205
rect 1652 204 1692 205
rect 1595 203 1633 204
rect 1652 203 1690 204
rect 1536 201 1571 202
rect 1537 199 1571 201
rect 1594 201 1633 203
rect 1651 202 1689 203
rect 1651 201 1688 202
rect 1594 199 1632 201
rect 1651 200 1687 201
rect 1651 199 1685 200
rect 1538 198 1571 199
rect 1538 197 1570 198
rect 1539 195 1570 197
rect 1540 194 1570 195
rect 1593 196 1631 199
rect 1651 198 1684 199
rect 1651 197 1683 198
rect 1651 196 1681 197
rect 1593 194 1630 196
rect 1541 192 1570 194
rect 1542 191 1570 192
rect 1543 190 1570 191
rect 1544 188 1570 190
rect 1545 187 1570 188
rect 1546 186 1570 187
rect 1547 185 1570 186
rect 1548 184 1570 185
rect 1550 183 1570 184
rect 1551 182 1570 183
rect 1552 181 1570 182
rect 995 180 1063 181
rect 1164 180 1245 181
rect 1285 180 1353 181
rect 1554 180 1570 181
rect 1592 193 1630 194
rect 1651 195 1680 196
rect 1651 194 1678 195
rect 1651 193 1677 194
rect 1592 189 1629 193
rect 1651 192 1676 193
rect 1651 191 1674 192
rect 1651 190 1673 191
rect 1651 189 1672 190
rect 1592 183 1628 189
rect 1651 188 1671 189
rect 1651 187 1670 188
rect 1651 186 1669 187
rect 1652 185 1668 186
rect 1652 183 1667 185
rect 503 179 693 180
rect 815 179 880 180
rect 1165 179 1247 180
rect 1286 179 1352 180
rect 1555 179 1571 180
rect 1166 178 1247 179
rect 1556 178 1571 179
rect 1167 177 1249 178
rect 1558 177 1571 178
rect 1592 177 1627 183
rect 1652 182 1666 183
rect 1652 181 1665 182
rect 1652 179 1664 181
rect 1652 178 1663 179
rect 1168 176 1249 177
rect 1559 176 1571 177
rect 1169 175 1251 176
rect 1560 175 1571 176
rect 1170 174 1251 175
rect 1562 174 1571 175
rect 1171 173 1253 174
rect 1563 173 1572 174
rect 1172 172 1253 173
rect 1564 172 1572 173
rect 1593 172 1627 177
rect 1653 176 1662 178
rect 1653 175 1661 176
rect 1653 174 1660 175
rect 1173 171 1255 172
rect 1565 171 1572 172
rect 1174 170 1256 171
rect 1567 170 1572 171
rect 1175 169 1257 170
rect 1568 169 1573 170
rect 1594 169 1627 172
rect 1654 173 1660 174
rect 1654 171 1659 173
rect 1654 170 1658 171
rect 1176 168 1257 169
rect 1569 168 1573 169
rect 1571 167 1573 168
rect 1595 167 1627 169
rect 1655 169 1658 170
rect 1655 167 1657 169
rect 1572 166 1573 167
rect 1596 165 1627 167
rect 1597 164 1627 165
rect 1597 163 1628 164
rect 1598 161 1628 163
rect 1599 159 1628 161
rect 1600 158 1628 159
rect 1601 156 1629 158
rect 1602 155 1629 156
rect 1603 154 1629 155
rect 1604 153 1629 154
rect 1605 152 1630 153
rect 1606 151 1630 152
rect 1607 150 1630 151
rect 1608 149 1630 150
rect 1609 148 1631 149
rect 1610 147 1631 148
rect 1611 146 1631 147
rect 1612 145 1632 146
rect 1613 144 1632 145
rect 1615 143 1632 144
rect 1616 142 1633 143
rect 1617 141 1633 142
rect 1619 140 1633 141
rect 1620 139 1634 140
rect 1303 138 1316 139
rect 1622 138 1634 139
rect 489 137 513 138
rect 530 137 539 138
rect 736 137 745 138
rect 833 137 841 138
rect 488 135 514 137
rect 488 134 513 135
rect 488 131 514 134
rect 489 129 513 131
rect 479 125 524 126
rect 478 117 524 125
rect 479 116 523 117
rect 530 116 540 137
rect 586 134 640 135
rect 585 128 641 134
rect 685 132 722 133
rect 585 125 640 128
rect 629 119 640 125
rect 684 124 723 132
rect 685 123 722 124
rect 697 122 710 123
rect 697 121 709 122
rect 698 119 709 121
rect 735 120 745 137
rect 783 129 823 130
rect 783 123 824 129
rect 782 121 824 123
rect 783 120 824 121
rect 722 119 745 120
rect 797 119 809 120
rect 629 118 639 119
rect 530 115 541 116
rect 543 115 544 116
rect 545 115 547 116
rect 628 115 639 118
rect 697 117 709 119
rect 697 115 710 117
rect 495 113 508 114
rect 491 112 511 113
rect 489 111 514 112
rect 487 110 515 111
rect 485 109 517 110
rect 484 108 518 109
rect 483 107 519 108
rect 482 106 519 107
rect 482 105 520 106
rect 530 105 549 115
rect 628 112 638 115
rect 697 114 711 115
rect 696 112 711 114
rect 627 108 638 112
rect 695 111 712 112
rect 695 110 713 111
rect 721 110 745 119
rect 798 114 809 119
rect 694 109 714 110
rect 693 108 714 109
rect 626 107 638 108
rect 692 107 716 108
rect 578 106 648 107
rect 691 106 717 107
rect 481 104 498 105
rect 505 104 521 105
rect 481 103 494 104
rect 508 103 521 104
rect 480 102 493 103
rect 509 102 521 103
rect 480 97 492 102
rect 510 101 521 102
rect 530 104 541 105
rect 510 100 522 101
rect 510 99 521 100
rect 510 97 522 99
rect 481 96 493 97
rect 509 96 521 97
rect 481 95 495 96
rect 507 95 521 96
rect 482 94 498 95
rect 504 94 520 95
rect 482 93 520 94
rect 483 92 519 93
rect 484 91 518 92
rect 485 90 517 91
rect 486 89 516 90
rect 488 88 515 89
rect 490 87 512 88
rect 492 86 510 87
rect 489 81 499 82
rect 488 70 500 81
rect 530 80 540 104
rect 577 98 649 106
rect 690 105 718 106
rect 689 104 719 105
rect 688 103 703 104
rect 705 103 721 104
rect 687 102 702 103
rect 705 102 722 103
rect 685 101 702 102
rect 706 101 725 102
rect 684 100 701 101
rect 707 100 725 101
rect 682 99 700 100
rect 708 99 725 100
rect 680 98 699 99
rect 709 98 725 99
rect 578 97 648 98
rect 679 97 698 98
rect 711 97 724 98
rect 605 96 617 97
rect 680 96 697 97
rect 712 96 723 97
rect 606 86 616 96
rect 681 95 696 96
rect 713 95 723 96
rect 682 94 695 95
rect 714 94 722 95
rect 682 93 693 94
rect 717 93 721 94
rect 683 92 692 93
rect 718 92 721 93
rect 684 91 690 92
rect 685 90 689 91
rect 606 85 617 86
rect 586 84 639 85
rect 530 79 539 80
rect 585 75 640 84
rect 586 74 640 75
rect 488 69 540 70
rect 488 61 542 69
rect 489 60 542 61
rect 630 59 640 74
rect 693 71 703 86
rect 735 80 745 110
rect 797 109 809 114
rect 797 106 810 109
rect 796 105 810 106
rect 832 108 842 137
rect 888 128 942 136
rect 1000 135 1009 136
rect 1000 128 1010 135
rect 888 127 900 128
rect 902 127 903 128
rect 937 127 939 128
rect 888 126 899 127
rect 888 125 898 126
rect 888 124 899 125
rect 888 123 941 124
rect 888 117 942 123
rect 999 122 1010 128
rect 999 121 1011 122
rect 998 118 1011 121
rect 888 116 941 117
rect 888 115 900 116
rect 998 115 1012 118
rect 888 114 899 115
rect 997 114 1013 115
rect 888 113 898 114
rect 996 113 1013 114
rect 888 112 899 113
rect 996 112 1014 113
rect 888 111 900 112
rect 902 111 903 112
rect 940 111 941 112
rect 995 111 1014 112
rect 832 107 844 108
rect 846 107 847 108
rect 848 107 850 108
rect 796 103 811 105
rect 795 100 811 103
rect 795 99 812 100
rect 794 98 813 99
rect 793 96 813 98
rect 832 97 852 107
rect 888 103 943 111
rect 994 110 1015 111
rect 994 109 1016 110
rect 993 108 1017 109
rect 992 107 1018 108
rect 992 106 1019 107
rect 990 104 1004 106
rect 1006 105 1020 106
rect 1006 104 1021 105
rect 988 103 1003 104
rect 1007 103 1023 104
rect 889 102 942 103
rect 987 102 1002 103
rect 1008 102 1024 103
rect 909 99 921 102
rect 986 101 1001 102
rect 1009 101 1026 102
rect 985 100 1000 101
rect 1010 100 1028 101
rect 983 99 1000 100
rect 1011 99 1028 100
rect 908 98 921 99
rect 982 98 999 99
rect 1012 98 1028 99
rect 881 97 906 98
rect 907 97 922 98
rect 923 97 946 98
rect 947 97 949 98
rect 980 97 998 98
rect 1013 97 1028 98
rect 832 96 851 97
rect 879 96 950 97
rect 980 96 997 97
rect 1014 96 1027 97
rect 793 95 814 96
rect 792 94 815 95
rect 791 93 815 94
rect 791 92 816 93
rect 790 91 803 92
rect 805 91 817 92
rect 789 89 802 91
rect 805 90 818 91
rect 805 89 819 90
rect 788 88 801 89
rect 806 88 820 89
rect 787 87 801 88
rect 807 87 821 88
rect 786 86 800 87
rect 807 86 822 87
rect 785 85 799 86
rect 808 85 823 86
rect 784 84 799 85
rect 809 84 824 85
rect 783 83 798 84
rect 809 83 825 84
rect 782 82 797 83
rect 810 82 826 83
rect 780 81 796 82
rect 811 81 827 82
rect 779 80 795 81
rect 812 80 826 81
rect 778 79 795 80
rect 813 79 825 80
rect 778 78 794 79
rect 814 78 824 79
rect 779 77 793 78
rect 815 77 824 78
rect 779 76 792 77
rect 816 76 823 77
rect 781 75 791 76
rect 818 75 822 76
rect 781 74 790 75
rect 819 74 821 75
rect 783 73 788 74
rect 784 72 787 73
rect 693 70 704 71
rect 693 60 747 70
rect 832 59 842 96
rect 879 89 951 96
rect 980 95 996 96
rect 1016 95 1026 96
rect 981 94 995 95
rect 1017 94 1026 95
rect 982 93 993 94
rect 1019 93 1025 94
rect 983 92 992 93
rect 1020 92 1024 93
rect 984 91 991 92
rect 985 90 990 91
rect 986 89 988 90
rect 879 88 950 89
rect 914 85 915 86
rect 995 85 1000 86
rect 1001 85 1003 86
rect 904 84 925 85
rect 898 83 931 84
rect 896 82 934 83
rect 893 81 936 82
rect 892 80 938 81
rect 890 79 939 80
rect 889 78 940 79
rect 888 77 942 78
rect 887 76 942 77
rect 887 75 905 76
rect 924 75 943 76
rect 886 74 902 75
rect 928 74 943 75
rect 886 69 899 74
rect 930 73 944 74
rect 931 72 944 73
rect 932 71 944 72
rect 931 69 944 71
rect 886 68 900 69
rect 930 68 944 69
rect 994 71 1004 85
rect 1036 80 1046 138
rect 1137 137 1146 138
rect 1299 137 1320 138
rect 1105 135 1106 136
rect 1098 134 1109 135
rect 1095 133 1113 134
rect 1093 132 1114 133
rect 1092 131 1116 132
rect 1091 130 1117 131
rect 1090 129 1118 130
rect 1089 128 1119 129
rect 1136 128 1147 137
rect 1298 136 1321 137
rect 1296 135 1323 136
rect 1295 134 1324 135
rect 1088 127 1147 128
rect 1087 126 1147 127
rect 1086 125 1102 126
rect 1105 125 1147 126
rect 1086 124 1100 125
rect 1108 124 1147 125
rect 1189 124 1245 134
rect 1294 133 1325 134
rect 1293 132 1326 133
rect 1292 131 1327 132
rect 1291 130 1327 131
rect 1291 129 1304 130
rect 1315 129 1328 130
rect 1291 128 1303 129
rect 1316 128 1328 129
rect 1291 127 1302 128
rect 1317 127 1329 128
rect 1086 123 1098 124
rect 1110 123 1147 124
rect 1233 123 1245 124
rect 1085 122 1097 123
rect 1111 122 1147 123
rect 1234 122 1244 123
rect 1085 121 1096 122
rect 1084 120 1096 121
rect 1112 120 1147 122
rect 1084 118 1095 120
rect 1113 118 1147 120
rect 1084 111 1094 118
rect 1113 117 1124 118
rect 1136 117 1147 118
rect 1114 112 1124 117
rect 1137 116 1147 117
rect 1136 112 1147 116
rect 1233 117 1244 122
rect 1290 121 1301 127
rect 1318 125 1329 127
rect 1319 123 1329 125
rect 1318 121 1329 123
rect 1291 120 1302 121
rect 1317 120 1329 121
rect 1291 119 1304 120
rect 1315 119 1328 120
rect 1291 118 1305 119
rect 1314 118 1328 119
rect 1291 117 1327 118
rect 1233 113 1243 117
rect 1292 116 1327 117
rect 1293 115 1326 116
rect 1293 114 1325 115
rect 1295 113 1324 114
rect 1084 110 1095 111
rect 1113 110 1147 112
rect 1084 108 1096 110
rect 1112 108 1147 110
rect 1232 109 1243 113
rect 1296 112 1323 113
rect 1298 111 1321 112
rect 1299 110 1320 111
rect 1304 109 1316 110
rect 1232 108 1242 109
rect 1085 107 1096 108
rect 1111 107 1147 108
rect 1085 106 1098 107
rect 1110 106 1147 107
rect 1086 105 1099 106
rect 1109 105 1147 106
rect 1086 104 1101 105
rect 1107 104 1147 105
rect 1086 103 1147 104
rect 1087 102 1147 103
rect 1231 106 1242 108
rect 1332 107 1336 108
rect 1325 106 1337 107
rect 1231 102 1241 106
rect 1285 104 1337 106
rect 1088 101 1120 102
rect 1136 101 1147 102
rect 1230 101 1241 102
rect 1089 100 1119 101
rect 1137 100 1147 101
rect 1182 100 1252 101
rect 1090 99 1118 100
rect 1091 98 1117 99
rect 1092 97 1115 98
rect 1094 96 1114 97
rect 1096 95 1111 96
rect 1098 94 1109 95
rect 1094 71 1104 86
rect 1136 81 1147 100
rect 1181 92 1253 100
rect 1284 98 1337 104
rect 1284 97 1333 98
rect 1285 96 1326 97
rect 1300 95 1312 96
rect 1339 95 1349 138
rect 1624 137 1634 138
rect 1625 136 1635 137
rect 1627 135 1635 136
rect 1629 134 1636 135
rect 1631 133 1636 134
rect 1634 132 1637 133
rect 1640 100 1653 101
rect 1414 97 1435 100
rect 1441 97 1459 100
rect 1464 98 1484 100
rect 1465 97 1484 98
rect 1492 97 1508 100
rect 1514 98 1535 100
rect 1544 98 1562 100
rect 1566 99 1580 100
rect 1598 99 1615 100
rect 1636 99 1658 100
rect 1566 98 1581 99
rect 1598 98 1616 99
rect 1633 98 1660 99
rect 1514 97 1534 98
rect 1545 97 1562 98
rect 1567 97 1581 98
rect 1599 97 1615 98
rect 1631 97 1642 98
rect 1649 97 1660 98
rect 1686 97 1707 100
rect 1714 98 1735 100
rect 1715 97 1735 98
rect 1744 98 1776 100
rect 1744 97 1777 98
rect 1787 97 1820 100
rect 1418 96 1431 97
rect 1445 96 1455 97
rect 1468 96 1481 97
rect 1496 96 1505 97
rect 1518 96 1531 97
rect 1548 96 1559 97
rect 1570 96 1582 97
rect 1603 96 1612 97
rect 1630 96 1639 97
rect 1652 96 1660 97
rect 1690 96 1703 97
rect 1719 96 1731 97
rect 1748 96 1759 97
rect 1768 96 1777 97
rect 1791 96 1803 97
rect 1811 96 1820 97
rect 1419 95 1430 96
rect 1445 95 1452 96
rect 1469 95 1480 96
rect 1496 95 1503 96
rect 1519 95 1530 96
rect 1549 95 1558 96
rect 1572 95 1583 96
rect 1604 95 1611 96
rect 1628 95 1638 96
rect 1653 95 1661 96
rect 1691 95 1702 96
rect 1719 95 1730 96
rect 1301 94 1312 95
rect 1182 91 1252 92
rect 1209 90 1221 91
rect 1137 80 1146 81
rect 994 70 1005 71
rect 1094 70 1105 71
rect 994 69 1047 70
rect 887 67 903 68
rect 927 67 943 68
rect 887 66 907 67
rect 924 66 943 67
rect 888 65 942 66
rect 889 64 942 65
rect 890 63 941 64
rect 891 62 940 63
rect 893 61 938 62
rect 894 60 936 61
rect 994 60 1048 69
rect 1094 60 1148 70
rect 897 59 933 60
rect 1210 59 1221 90
rect 1301 83 1311 94
rect 1324 93 1326 94
rect 1329 93 1336 94
rect 1338 93 1349 95
rect 1323 92 1349 93
rect 1322 85 1349 92
rect 1323 84 1349 85
rect 1338 83 1349 84
rect 1302 82 1304 83
rect 1305 82 1310 83
rect 1296 79 1306 80
rect 1296 70 1307 79
rect 1339 78 1349 83
rect 1420 79 1429 95
rect 1444 94 1451 95
rect 1470 94 1481 95
rect 1444 93 1449 94
rect 1471 93 1481 94
rect 1496 94 1502 95
rect 1496 93 1501 94
rect 1443 92 1448 93
rect 1471 92 1482 93
rect 1496 92 1500 93
rect 1442 91 1447 92
rect 1472 91 1482 92
rect 1495 91 1500 92
rect 1441 90 1446 91
rect 1472 90 1483 91
rect 1495 90 1499 91
rect 1441 89 1445 90
rect 1473 89 1483 90
rect 1494 89 1499 90
rect 1440 88 1444 89
rect 1439 87 1443 88
rect 1474 87 1484 89
rect 1494 88 1498 89
rect 1438 86 1442 87
rect 1437 85 1441 86
rect 1475 85 1485 87
rect 1493 86 1497 88
rect 1436 84 1440 85
rect 1435 83 1439 84
rect 1476 83 1486 85
rect 1492 84 1496 86
rect 1491 83 1495 84
rect 1434 82 1438 83
rect 1477 82 1487 83
rect 1491 82 1494 83
rect 1433 81 1439 82
rect 1432 80 1439 81
rect 1478 81 1487 82
rect 1490 81 1494 82
rect 1478 80 1488 81
rect 1490 80 1493 81
rect 1430 79 1440 80
rect 1479 79 1488 80
rect 1489 79 1493 80
rect 1420 78 1441 79
rect 1479 78 1492 79
rect 1420 76 1442 78
rect 1480 77 1492 78
rect 1480 76 1491 77
rect 1296 69 1350 70
rect 1296 61 1351 69
rect 1296 60 1350 61
rect 1420 60 1429 76
rect 1431 75 1443 76
rect 1432 74 1444 75
rect 1433 73 1444 74
rect 1434 72 1445 73
rect 1434 71 1446 72
rect 1435 70 1447 71
rect 1436 69 1447 70
rect 1436 68 1448 69
rect 1437 67 1449 68
rect 1438 65 1450 67
rect 1439 64 1451 65
rect 1440 63 1452 64
rect 1441 62 1453 63
rect 1441 61 1454 62
rect 1442 60 1454 61
rect 1419 59 1430 60
rect 1443 59 1456 60
rect 1481 59 1491 76
rect 1519 71 1529 95
rect 1550 90 1557 95
rect 1572 94 1584 95
rect 1573 93 1585 94
rect 1573 92 1586 93
rect 1573 90 1587 92
rect 1550 89 1556 90
rect 1551 71 1556 89
rect 1520 69 1529 71
rect 1520 65 1530 69
rect 1550 67 1556 71
rect 1573 89 1588 90
rect 1605 89 1610 95
rect 1627 94 1636 95
rect 1654 94 1661 95
rect 1626 93 1635 94
rect 1655 93 1661 94
rect 1625 92 1634 93
rect 1656 92 1661 93
rect 1624 91 1634 92
rect 1623 90 1633 91
rect 1657 90 1661 92
rect 1573 88 1589 89
rect 1550 66 1555 67
rect 1521 63 1531 65
rect 1549 63 1555 66
rect 1521 62 1532 63
rect 1548 62 1554 63
rect 1522 61 1533 62
rect 1547 61 1554 62
rect 1573 62 1577 88
rect 1578 87 1590 88
rect 1579 86 1591 87
rect 1579 85 1592 86
rect 1580 84 1593 85
rect 1581 83 1594 84
rect 1582 82 1594 83
rect 1583 81 1595 82
rect 1584 80 1596 81
rect 1585 79 1597 80
rect 1585 78 1598 79
rect 1586 77 1599 78
rect 1587 76 1600 77
rect 1588 75 1601 76
rect 1589 74 1601 75
rect 1590 73 1602 74
rect 1590 72 1603 73
rect 1591 71 1604 72
rect 1592 70 1605 71
rect 1606 70 1609 89
rect 1622 88 1632 90
rect 1621 85 1631 88
rect 1658 87 1661 90
rect 1692 93 1702 95
rect 1620 84 1631 85
rect 1620 82 1630 84
rect 1619 72 1630 82
rect 1692 81 1701 93
rect 1720 81 1730 95
rect 1692 77 1730 81
rect 1644 76 1664 77
rect 1692 76 1702 77
rect 1644 74 1665 76
rect 1647 73 1663 74
rect 1650 72 1662 73
rect 1593 69 1609 70
rect 1594 68 1609 69
rect 1620 68 1631 72
rect 1651 70 1661 72
rect 1595 66 1609 68
rect 1621 66 1632 68
rect 1596 65 1609 66
rect 1597 64 1609 65
rect 1622 64 1633 66
rect 1598 63 1609 64
rect 1623 63 1634 64
rect 1599 62 1609 63
rect 1624 62 1635 63
rect 1573 61 1578 62
rect 1522 60 1534 61
rect 1546 60 1553 61
rect 1523 59 1536 60
rect 1544 59 1553 60
rect 1572 59 1578 61
rect 1600 60 1609 62
rect 1625 61 1635 62
rect 1652 61 1661 70
rect 1626 60 1636 61
rect 1601 59 1609 60
rect 1627 59 1638 60
rect 630 58 639 59
rect 833 58 841 59
rect 899 58 931 59
rect 1211 58 1220 59
rect 1419 58 1431 59
rect 1443 58 1457 59
rect 1480 58 1492 59
rect 1524 58 1552 59
rect 1571 58 1579 59
rect 1602 58 1609 59
rect 1628 58 1639 59
rect 1651 58 1661 61
rect 1692 61 1701 76
rect 1692 60 1702 61
rect 1691 59 1702 60
rect 1720 59 1730 77
rect 1749 80 1759 96
rect 1771 95 1777 96
rect 1772 94 1777 95
rect 1773 92 1777 94
rect 1774 89 1777 92
rect 1771 84 1773 85
rect 1770 81 1773 84
rect 1769 80 1773 81
rect 1749 76 1773 80
rect 1749 59 1759 76
rect 1769 75 1773 76
rect 1770 72 1773 75
rect 1771 71 1773 72
rect 1792 80 1802 96
rect 1814 95 1820 96
rect 1815 94 1820 95
rect 1816 92 1820 94
rect 1817 89 1820 92
rect 1814 83 1817 85
rect 1813 81 1817 83
rect 1812 80 1817 81
rect 1792 76 1817 80
rect 1778 66 1780 67
rect 1777 64 1780 66
rect 1776 62 1780 64
rect 1775 61 1780 62
rect 1774 60 1779 61
rect 1773 59 1779 60
rect 1792 60 1802 76
rect 1812 75 1817 76
rect 1813 73 1817 75
rect 1814 71 1817 73
rect 1821 66 1824 67
rect 1820 65 1824 66
rect 1820 64 1823 65
rect 1819 62 1823 64
rect 1818 61 1823 62
rect 1817 60 1823 61
rect 1792 59 1803 60
rect 1816 59 1822 60
rect 1691 58 1703 59
rect 1719 58 1731 59
rect 1748 58 1761 59
rect 1771 58 1779 59
rect 1791 58 1804 59
rect 1814 58 1822 59
rect 906 57 925 58
rect 1415 57 1435 58
rect 1444 57 1460 58
rect 1476 57 1496 58
rect 1525 57 1551 58
rect 1568 57 1583 58
rect 1603 57 1609 58
rect 1630 57 1642 58
rect 1650 57 1661 58
rect 1687 57 1706 58
rect 1715 57 1735 58
rect 1414 55 1435 57
rect 1445 55 1460 57
rect 1475 55 1498 57
rect 1526 56 1550 57
rect 1528 55 1548 56
rect 1567 55 1584 57
rect 1604 56 1609 57
rect 1632 56 1661 57
rect 1531 54 1545 55
rect 1605 54 1609 56
rect 1634 55 1658 56
rect 1686 55 1707 57
rect 1714 55 1735 57
rect 1743 56 1779 58
rect 1787 57 1822 58
rect 1786 56 1822 57
rect 1743 55 1778 56
rect 1786 55 1821 56
rect 1638 54 1653 55
rect 501 43 504 44
rect 714 43 717 44
rect 768 43 770 44
rect 1190 43 1193 44
rect 481 40 495 41
rect 480 37 496 40
rect 480 36 495 37
rect 480 35 487 36
rect 480 30 486 35
rect 480 29 487 30
rect 480 27 494 29
rect 480 25 495 27
rect 480 23 494 25
rect 480 22 487 23
rect 480 16 486 22
rect 480 15 494 16
rect 480 14 495 15
rect 480 11 496 14
rect 499 11 504 43
rect 613 42 615 43
rect 547 38 550 39
rect 545 37 550 38
rect 611 37 616 42
rect 514 33 519 34
rect 533 33 538 34
rect 544 33 550 37
rect 612 36 616 37
rect 565 33 567 34
rect 575 33 580 34
rect 598 33 603 34
rect 626 33 631 34
rect 640 33 645 34
rect 665 33 671 34
rect 689 33 692 34
rect 706 33 709 34
rect 712 33 718 43
rect 730 40 748 41
rect 729 39 748 40
rect 729 37 749 39
rect 729 36 748 37
rect 735 35 743 36
rect 512 32 521 33
rect 531 32 540 33
rect 542 32 553 33
rect 557 32 560 33
rect 563 32 568 33
rect 573 32 582 33
rect 591 32 594 33
rect 596 32 604 33
rect 612 32 616 33
rect 624 32 633 33
rect 638 32 647 33
rect 662 32 673 33
rect 680 32 694 33
rect 703 32 718 33
rect 510 31 522 32
rect 530 31 554 32
rect 510 30 523 31
rect 529 30 554 31
rect 509 29 523 30
rect 528 29 554 30
rect 508 28 524 29
rect 528 28 540 29
rect 542 28 553 29
rect 556 28 568 32
rect 572 31 584 32
rect 571 30 584 31
rect 570 29 585 30
rect 590 29 606 32
rect 570 28 586 29
rect 508 27 514 28
rect 518 27 524 28
rect 508 25 513 27
rect 508 24 514 25
rect 519 24 524 27
rect 527 26 534 28
rect 527 25 533 26
rect 508 21 525 24
rect 508 19 524 21
rect 526 19 532 25
rect 508 17 513 19
rect 526 18 533 19
rect 527 17 533 18
rect 508 16 514 17
rect 527 16 534 17
rect 544 16 550 28
rect 556 27 576 28
rect 580 27 586 28
rect 590 28 607 29
rect 556 26 564 27
rect 568 26 575 27
rect 580 26 587 27
rect 556 25 563 26
rect 508 15 515 16
rect 520 15 523 16
rect 528 15 535 16
rect 538 15 540 16
rect 509 13 524 15
rect 528 14 540 15
rect 544 15 551 16
rect 544 14 554 15
rect 528 13 541 14
rect 545 13 554 14
rect 510 12 523 13
rect 529 12 541 13
rect 511 11 523 12
rect 530 11 541 12
rect 546 11 554 13
rect 556 11 562 25
rect 568 17 574 26
rect 581 24 587 26
rect 582 20 587 24
rect 581 17 587 20
rect 568 16 575 17
rect 580 16 587 17
rect 590 26 597 28
rect 601 26 607 28
rect 569 15 576 16
rect 579 15 586 16
rect 570 14 586 15
rect 570 13 585 14
rect 571 12 584 13
rect 572 11 583 12
rect 590 11 596 26
rect 602 11 607 26
rect 611 11 616 32
rect 623 31 633 32
rect 622 30 633 31
rect 636 30 648 32
rect 662 31 674 32
rect 680 31 695 32
rect 702 31 718 32
rect 621 29 633 30
rect 635 29 648 30
rect 661 30 675 31
rect 621 28 632 29
rect 635 28 647 29
rect 661 28 676 30
rect 620 26 627 28
rect 635 27 641 28
rect 661 27 664 28
rect 670 27 676 28
rect 634 26 641 27
rect 662 26 663 27
rect 620 23 626 26
rect 635 25 641 26
rect 671 25 676 27
rect 635 24 643 25
rect 665 24 676 25
rect 635 23 645 24
rect 663 23 676 24
rect 620 20 625 23
rect 636 22 646 23
rect 662 22 676 23
rect 636 21 647 22
rect 661 21 676 22
rect 637 20 648 21
rect 620 17 626 20
rect 640 19 648 20
rect 641 18 648 19
rect 660 20 676 21
rect 660 19 666 20
rect 660 18 665 19
rect 671 18 676 20
rect 620 16 627 17
rect 620 15 628 16
rect 631 15 633 16
rect 636 15 638 16
rect 642 15 648 18
rect 659 16 665 18
rect 670 16 676 18
rect 621 13 634 15
rect 622 12 634 13
rect 623 11 634 12
rect 635 13 648 15
rect 660 15 666 16
rect 669 15 676 16
rect 660 13 676 15
rect 635 12 647 13
rect 661 12 676 13
rect 635 11 646 12
rect 662 11 676 12
rect 680 29 696 31
rect 680 28 697 29
rect 701 28 718 31
rect 680 27 687 28
rect 690 27 697 28
rect 680 24 686 27
rect 481 10 495 11
rect 500 10 504 11
rect 513 10 522 11
rect 531 10 540 11
rect 547 10 554 11
rect 557 10 561 11
rect 573 10 582 11
rect 591 10 595 11
rect 602 10 606 11
rect 612 10 616 11
rect 624 10 633 11
rect 636 10 645 11
rect 662 10 669 11
rect 672 10 675 11
rect 680 10 685 24
rect 691 11 697 27
rect 700 27 707 28
rect 710 27 718 28
rect 700 23 706 27
rect 711 25 718 27
rect 700 20 705 23
rect 700 17 706 20
rect 712 18 718 25
rect 700 16 707 17
rect 711 16 718 18
rect 700 15 708 16
rect 710 15 718 16
rect 701 13 718 15
rect 702 12 718 13
rect 703 11 718 12
rect 736 11 742 35
rect 752 33 757 34
rect 750 32 759 33
rect 749 31 760 32
rect 748 30 761 31
rect 747 29 761 30
rect 747 28 762 29
rect 746 27 752 28
rect 746 25 751 27
rect 757 26 762 28
rect 745 24 752 25
rect 757 24 763 26
rect 745 20 763 24
rect 745 19 762 20
rect 745 18 752 19
rect 746 17 751 18
rect 746 16 752 17
rect 746 15 753 16
rect 758 15 762 16
rect 747 13 762 15
rect 748 12 762 13
rect 749 11 761 12
rect 766 11 771 43
rect 935 42 938 43
rect 993 42 995 43
rect 1189 42 1194 43
rect 1280 42 1282 43
rect 934 37 939 42
rect 981 38 984 39
rect 980 37 984 38
rect 991 37 996 42
rect 1068 40 1080 41
rect 935 36 938 37
rect 979 34 984 37
rect 992 36 996 37
rect 1067 39 1082 40
rect 1067 38 1083 39
rect 1067 36 1084 38
rect 1067 35 1074 36
rect 1076 35 1084 36
rect 781 33 785 34
rect 800 33 805 34
rect 816 33 820 34
rect 839 33 842 34
rect 849 33 853 34
rect 869 33 873 34
rect 880 33 884 34
rect 921 33 926 34
rect 949 33 954 34
rect 963 33 969 34
rect 978 33 985 34
rect 1007 33 1012 34
rect 1031 33 1034 34
rect 1047 33 1052 34
rect 778 32 787 33
rect 798 32 807 33
rect 813 32 823 33
rect 831 32 835 33
rect 837 32 844 33
rect 848 32 855 33
rect 862 32 875 33
rect 878 32 886 33
rect 893 32 897 33
rect 904 32 908 33
rect 913 32 917 33
rect 919 32 927 33
rect 934 32 938 33
rect 947 32 956 33
rect 961 32 971 33
rect 976 32 988 33
rect 992 32 996 33
rect 1005 32 1014 33
rect 1022 32 1026 33
rect 1028 32 1036 33
rect 1045 32 1054 33
rect 777 30 789 32
rect 797 31 807 32
rect 812 31 824 32
rect 831 31 845 32
rect 846 31 856 32
rect 796 30 807 31
rect 776 29 790 30
rect 775 28 790 29
rect 795 29 807 30
rect 811 30 825 31
rect 811 29 826 30
rect 795 28 806 29
rect 810 28 827 29
rect 775 27 781 28
rect 785 27 791 28
rect 775 25 780 27
rect 774 24 780 25
rect 786 24 791 27
rect 794 27 801 28
rect 809 27 816 28
rect 820 27 827 28
rect 794 26 800 27
rect 774 19 791 24
rect 774 17 780 19
rect 793 18 799 26
rect 809 24 815 27
rect 821 25 827 27
rect 831 28 857 31
rect 831 25 837 28
rect 841 27 848 28
rect 851 27 857 28
rect 809 22 814 24
rect 808 21 814 22
rect 809 20 814 21
rect 793 17 800 18
rect 809 17 815 20
rect 822 19 828 25
rect 775 16 781 17
rect 794 16 801 17
rect 809 16 816 17
rect 821 16 827 19
rect 775 15 782 16
rect 786 15 790 16
rect 794 15 802 16
rect 805 15 807 16
rect 809 15 817 16
rect 820 15 827 16
rect 775 14 791 15
rect 776 13 790 14
rect 795 13 807 15
rect 810 14 826 15
rect 777 12 790 13
rect 796 12 807 13
rect 811 13 826 14
rect 811 12 825 13
rect 778 11 790 12
rect 797 11 807 12
rect 813 11 824 12
rect 831 11 836 25
rect 841 11 847 27
rect 852 13 857 27
rect 861 29 887 32
rect 861 28 888 29
rect 861 27 868 28
rect 871 27 879 28
rect 852 12 858 13
rect 852 11 857 12
rect 861 11 867 27
rect 871 25 878 27
rect 882 26 888 28
rect 872 11 877 25
rect 883 13 888 26
rect 892 17 897 32
rect 903 17 909 32
rect 892 16 898 17
rect 902 16 909 17
rect 892 15 899 16
rect 901 15 909 16
rect 892 13 909 15
rect 882 12 888 13
rect 893 12 909 13
rect 883 11 888 12
rect 894 11 909 12
rect 913 31 928 32
rect 913 28 929 31
rect 913 27 920 28
rect 923 27 930 28
rect 913 24 919 27
rect 913 13 918 24
rect 913 12 919 13
rect 692 10 696 11
rect 704 10 711 11
rect 713 10 717 11
rect 737 10 741 11
rect 750 10 760 11
rect 767 10 771 11
rect 779 10 789 11
rect 798 10 807 11
rect 814 10 823 11
rect 831 10 835 11
rect 842 10 846 11
rect 853 10 857 11
rect 862 10 866 11
rect 873 10 876 11
rect 883 10 887 11
rect 895 10 902 11
rect 905 10 908 11
rect 913 10 918 12
rect 924 11 930 27
rect 934 11 939 32
rect 946 31 956 32
rect 945 30 956 31
rect 944 29 956 30
rect 959 31 972 32
rect 959 29 973 31
rect 976 29 989 32
rect 943 28 955 29
rect 959 28 974 29
rect 977 28 988 29
rect 943 27 950 28
rect 960 27 962 28
rect 968 27 974 28
rect 943 26 949 27
rect 942 25 949 26
rect 969 25 974 27
rect 942 18 948 25
rect 963 24 974 25
rect 961 23 974 24
rect 959 22 974 23
rect 958 20 974 22
rect 958 19 964 20
rect 942 17 949 18
rect 943 16 949 17
rect 957 16 963 19
rect 969 18 974 20
rect 968 16 974 18
rect 943 15 951 16
rect 954 15 956 16
rect 944 13 956 15
rect 958 15 964 16
rect 967 15 974 16
rect 958 13 974 15
rect 979 18 984 28
rect 979 16 985 18
rect 979 15 986 16
rect 979 14 988 15
rect 945 12 956 13
rect 946 11 956 12
rect 959 11 974 13
rect 980 12 989 14
rect 981 11 989 12
rect 991 11 996 32
rect 1003 31 1015 32
rect 1022 31 1037 32
rect 1043 31 1054 32
rect 1002 30 1016 31
rect 1021 30 1038 31
rect 1002 29 1017 30
rect 1001 28 1017 29
rect 1022 28 1038 30
rect 1042 28 1054 31
rect 1067 29 1073 35
rect 1077 34 1084 35
rect 1078 33 1084 34
rect 1094 33 1098 34
rect 1111 33 1117 34
rect 1128 33 1133 34
rect 1147 33 1152 34
rect 1169 33 1171 34
rect 1179 33 1185 34
rect 1189 33 1195 42
rect 1220 40 1225 41
rect 1198 33 1201 34
rect 1079 31 1084 33
rect 1092 32 1101 33
rect 1109 32 1119 33
rect 1126 32 1135 33
rect 1144 32 1154 33
rect 1162 32 1165 33
rect 1168 32 1172 33
rect 1177 32 1186 33
rect 1189 32 1203 33
rect 1078 29 1084 31
rect 1090 30 1102 32
rect 1108 31 1119 32
rect 1125 31 1136 32
rect 1089 29 1103 30
rect 1107 29 1119 31
rect 1124 30 1137 31
rect 1123 29 1138 30
rect 1067 28 1074 29
rect 1076 28 1084 29
rect 1088 28 1104 29
rect 1000 27 1007 28
rect 1011 27 1018 28
rect 1000 24 1006 27
rect 1012 25 1018 27
rect 1021 27 1029 28
rect 1032 27 1038 28
rect 1021 25 1028 27
rect 1013 24 1018 25
rect 1022 24 1028 25
rect 1000 19 1005 24
rect 1013 19 1019 24
rect 1000 17 1006 19
rect 1013 18 1018 19
rect 1022 18 1027 24
rect 1033 23 1039 27
rect 1041 25 1048 28
rect 1067 27 1083 28
rect 1088 27 1094 28
rect 1098 27 1104 28
rect 1107 28 1114 29
rect 1115 28 1118 29
rect 1123 28 1130 29
rect 1131 28 1138 29
rect 1107 27 1112 28
rect 1034 22 1039 23
rect 1042 24 1050 25
rect 1042 23 1052 24
rect 1042 22 1053 23
rect 1067 22 1082 27
rect 1088 24 1093 27
rect 1099 24 1104 27
rect 1106 26 1112 27
rect 1122 26 1128 28
rect 1133 27 1138 28
rect 1143 29 1156 32
rect 1143 28 1157 29
rect 1143 27 1145 28
rect 1151 27 1157 28
rect 1133 26 1139 27
rect 1106 25 1113 26
rect 1122 25 1127 26
rect 1134 25 1139 26
rect 1152 25 1157 27
rect 1106 24 1115 25
rect 1122 24 1128 25
rect 1133 24 1139 25
rect 1146 24 1157 25
rect 1087 23 1104 24
rect 1107 23 1117 24
rect 1000 16 1007 17
rect 1012 16 1018 18
rect 1000 15 1008 16
rect 1010 15 1018 16
rect 1021 15 1027 18
rect 1033 15 1039 22
rect 1043 21 1054 22
rect 1044 20 1055 21
rect 1047 19 1055 20
rect 1048 18 1055 19
rect 1049 16 1055 18
rect 1001 14 1017 15
rect 1002 13 1016 14
rect 1022 13 1027 15
rect 1034 14 1039 15
rect 1003 12 1016 13
rect 1021 12 1028 13
rect 1004 11 1015 12
rect 1022 11 1027 12
rect 1033 11 1039 14
rect 1042 15 1044 16
rect 1048 15 1055 16
rect 1042 14 1055 15
rect 1042 12 1054 14
rect 1042 11 1053 12
rect 1067 11 1073 22
rect 1076 21 1083 22
rect 1077 20 1083 21
rect 1087 20 1105 23
rect 1107 22 1118 23
rect 1108 21 1119 22
rect 1109 20 1119 21
rect 1077 18 1084 20
rect 1087 19 1104 20
rect 1112 19 1120 20
rect 1087 18 1093 19
rect 1113 18 1120 19
rect 1078 16 1084 18
rect 1088 17 1093 18
rect 1088 16 1094 17
rect 1114 16 1120 18
rect 1122 19 1139 24
rect 1144 23 1157 24
rect 1143 22 1157 23
rect 1142 20 1157 22
rect 1141 19 1147 20
rect 1122 16 1128 19
rect 1136 16 1137 17
rect 1141 16 1146 19
rect 1152 17 1157 20
rect 1151 16 1157 17
rect 1078 15 1085 16
rect 1088 15 1095 16
rect 1100 15 1104 16
rect 1079 13 1085 15
rect 1089 13 1104 15
rect 1107 15 1109 16
rect 1113 15 1120 16
rect 1107 14 1120 15
rect 1123 15 1129 16
rect 1134 15 1138 16
rect 1107 13 1119 14
rect 1123 13 1138 15
rect 1141 15 1147 16
rect 1150 15 1157 16
rect 1141 13 1157 15
rect 1161 28 1172 32
rect 1176 31 1187 32
rect 1189 31 1204 32
rect 1175 30 1186 31
rect 1174 28 1186 30
rect 1189 29 1205 31
rect 1189 28 1206 29
rect 1161 27 1171 28
rect 1173 27 1181 28
rect 1161 25 1168 27
rect 1173 26 1180 27
rect 1189 26 1196 28
rect 1200 26 1206 28
rect 1079 12 1086 13
rect 1090 12 1103 13
rect 1106 12 1118 13
rect 1124 12 1138 13
rect 1142 12 1158 13
rect 1080 11 1086 12
rect 1091 11 1103 12
rect 1107 11 1118 12
rect 1125 11 1138 12
rect 1143 11 1158 12
rect 1161 11 1167 25
rect 1173 24 1179 26
rect 1173 20 1178 24
rect 1173 17 1179 20
rect 1173 16 1180 17
rect 1173 15 1181 16
rect 1185 15 1186 16
rect 1174 14 1187 15
rect 1175 12 1187 14
rect 1176 11 1187 12
rect 1189 11 1195 26
rect 1201 11 1206 26
rect 1219 13 1225 40
rect 1269 38 1272 39
rect 1267 34 1272 38
rect 1279 37 1284 42
rect 1292 38 1295 39
rect 1326 38 1329 39
rect 1279 36 1283 37
rect 1290 34 1295 38
rect 1325 37 1329 38
rect 1238 33 1242 34
rect 1254 33 1260 34
rect 1267 33 1273 34
rect 1289 33 1295 34
rect 1324 34 1329 37
rect 1661 35 1667 36
rect 1697 35 1699 36
rect 1714 35 1716 36
rect 1493 34 1503 35
rect 1508 34 1516 35
rect 1523 34 1530 35
rect 1538 34 1547 35
rect 1554 34 1564 35
rect 1572 34 1582 35
rect 1587 34 1595 35
rect 1603 34 1618 35
rect 1628 34 1643 35
rect 1659 34 1669 35
rect 1678 34 1688 35
rect 1697 34 1716 35
rect 1724 34 1734 35
rect 1737 34 1745 35
rect 1324 33 1330 34
rect 1341 33 1346 34
rect 1495 33 1501 34
rect 1510 33 1515 34
rect 1525 33 1531 34
rect 1541 33 1545 34
rect 1556 33 1562 34
rect 1574 33 1581 34
rect 1589 33 1593 34
rect 1230 32 1243 33
rect 1252 32 1261 33
rect 1264 32 1275 33
rect 1229 30 1245 32
rect 1251 31 1261 32
rect 1250 30 1262 31
rect 1229 28 1246 30
rect 1229 26 1236 28
rect 1240 26 1246 28
rect 1219 12 1226 13
rect 1219 11 1225 12
rect 1229 11 1235 26
rect 1241 13 1246 26
rect 1249 28 1261 30
rect 1263 29 1276 32
rect 1264 28 1275 29
rect 1249 26 1255 28
rect 1249 25 1256 26
rect 1249 24 1258 25
rect 1249 23 1260 24
rect 1250 22 1261 23
rect 1251 21 1262 22
rect 1252 20 1262 21
rect 1254 19 1263 20
rect 1256 18 1263 19
rect 1257 16 1263 18
rect 1250 15 1252 16
rect 1256 15 1263 16
rect 1267 18 1272 28
rect 1267 15 1273 18
rect 1249 13 1262 15
rect 1267 14 1276 15
rect 1267 13 1277 14
rect 1241 12 1247 13
rect 1249 12 1261 13
rect 1268 12 1277 13
rect 925 10 929 11
rect 935 10 938 11
rect 947 10 956 11
rect 961 10 967 11
rect 970 10 974 11
rect 982 10 988 11
rect 992 10 996 11
rect 1005 10 1013 11
rect 1022 10 1026 11
rect 1034 10 1038 11
rect 1042 10 1052 11
rect 1068 10 1072 11
rect 1080 10 1085 11
rect 1092 10 1102 11
rect 1108 10 1117 11
rect 1127 10 1137 11
rect 1144 10 1151 11
rect 1154 10 1157 11
rect 1162 10 1166 11
rect 1178 10 1186 11
rect 1190 10 1194 11
rect 1202 10 1205 11
rect 1220 10 1225 11
rect 1230 10 1233 11
rect 1241 10 1246 12
rect 1249 11 1260 12
rect 1269 11 1277 12
rect 1279 11 1284 33
rect 1287 31 1299 33
rect 1286 29 1299 31
rect 1287 28 1299 29
rect 1290 16 1295 28
rect 1302 17 1307 33
rect 1314 32 1318 33
rect 1313 17 1319 32
rect 1321 31 1333 33
rect 1339 32 1348 33
rect 1496 32 1501 33
rect 1338 31 1349 32
rect 1321 30 1334 31
rect 1337 30 1350 31
rect 1321 28 1333 30
rect 1337 29 1351 30
rect 1336 28 1351 29
rect 1302 16 1308 17
rect 1312 16 1319 17
rect 1290 15 1296 16
rect 1302 15 1309 16
rect 1311 15 1319 16
rect 1290 14 1299 15
rect 1302 14 1319 15
rect 1324 18 1329 28
rect 1336 27 1341 28
rect 1346 27 1351 28
rect 1335 24 1341 27
rect 1347 25 1352 27
rect 1346 24 1352 25
rect 1335 21 1353 24
rect 1496 22 1500 32
rect 1511 31 1514 33
rect 1526 32 1532 33
rect 1541 32 1544 33
rect 1526 31 1533 32
rect 1335 19 1352 21
rect 1324 16 1330 18
rect 1335 16 1341 19
rect 1496 18 1501 22
rect 1511 18 1513 31
rect 1526 29 1534 31
rect 1497 17 1502 18
rect 1510 17 1512 18
rect 1349 16 1350 17
rect 1497 16 1503 17
rect 1509 16 1512 17
rect 1526 17 1528 29
rect 1529 28 1535 29
rect 1530 27 1536 28
rect 1531 26 1537 27
rect 1532 25 1538 26
rect 1533 24 1539 25
rect 1533 23 1540 24
rect 1534 22 1541 23
rect 1542 22 1544 32
rect 1535 21 1544 22
rect 1536 20 1544 21
rect 1537 19 1544 20
rect 1538 17 1544 19
rect 1526 16 1529 17
rect 1539 16 1544 17
rect 1557 16 1562 33
rect 1575 32 1580 33
rect 1575 31 1581 32
rect 1576 29 1581 31
rect 1589 31 1592 33
rect 1589 29 1591 31
rect 1577 26 1582 29
rect 1588 27 1590 29
rect 1588 26 1589 27
rect 1578 24 1583 26
rect 1587 24 1589 26
rect 1605 26 1610 34
rect 1615 33 1618 34
rect 1630 33 1636 34
rect 1638 33 1644 34
rect 1658 33 1661 34
rect 1666 33 1669 34
rect 1680 33 1686 34
rect 1616 32 1619 33
rect 1630 32 1635 33
rect 1617 30 1619 32
rect 1615 26 1617 28
rect 1605 24 1617 26
rect 1579 21 1584 24
rect 1586 21 1588 24
rect 1580 19 1587 21
rect 1581 16 1586 19
rect 1605 16 1610 24
rect 1615 22 1617 24
rect 1616 21 1617 22
rect 1631 25 1635 32
rect 1640 30 1645 33
rect 1657 32 1661 33
rect 1657 31 1660 32
rect 1667 31 1669 33
rect 1641 28 1645 30
rect 1656 30 1660 31
rect 1668 30 1669 31
rect 1656 29 1661 30
rect 1656 28 1662 29
rect 1640 26 1645 28
rect 1657 27 1663 28
rect 1657 26 1665 27
rect 1639 25 1644 26
rect 1658 25 1667 26
rect 1631 24 1636 25
rect 1637 24 1642 25
rect 1659 24 1668 25
rect 1631 23 1642 24
rect 1660 23 1669 24
rect 1619 19 1620 20
rect 1618 17 1620 19
rect 1631 17 1635 23
rect 1637 22 1642 23
rect 1662 22 1670 23
rect 1638 21 1643 22
rect 1664 21 1670 22
rect 1638 20 1644 21
rect 1665 20 1670 21
rect 1639 19 1644 20
rect 1656 19 1657 20
rect 1639 18 1645 19
rect 1617 16 1620 17
rect 1324 15 1331 16
rect 1336 15 1343 16
rect 1348 15 1351 16
rect 1498 15 1505 16
rect 1507 15 1511 16
rect 1525 15 1529 16
rect 1540 15 1544 16
rect 1556 15 1562 16
rect 1324 14 1334 15
rect 1336 14 1351 15
rect 1499 14 1510 15
rect 1523 14 1532 15
rect 1541 14 1544 15
rect 1554 14 1564 15
rect 1582 14 1585 16
rect 1604 15 1611 16
rect 1616 15 1620 16
rect 1630 16 1635 17
rect 1640 17 1645 18
rect 1656 18 1658 19
rect 1640 16 1646 17
rect 1656 16 1659 18
rect 1666 17 1670 20
rect 1666 16 1669 17
rect 1681 16 1686 33
rect 1697 33 1700 34
rect 1697 32 1699 33
rect 1697 31 1698 32
rect 1696 30 1698 31
rect 1697 29 1698 30
rect 1704 16 1709 34
rect 1712 33 1716 34
rect 1726 33 1732 34
rect 1713 32 1716 33
rect 1714 30 1716 32
rect 1727 31 1732 33
rect 1739 33 1743 34
rect 1739 32 1742 33
rect 1739 31 1741 32
rect 1728 29 1733 31
rect 1738 29 1740 31
rect 1729 28 1734 29
rect 1730 27 1734 28
rect 1737 27 1739 29
rect 1730 26 1735 27
rect 1736 26 1738 27
rect 1731 25 1738 26
rect 1731 24 1737 25
rect 1732 16 1737 24
rect 1630 15 1636 16
rect 1641 15 1647 16
rect 1656 15 1660 16
rect 1665 15 1668 16
rect 1680 15 1686 16
rect 1703 15 1709 16
rect 1731 15 1737 16
rect 1602 14 1619 15
rect 1628 14 1638 15
rect 1642 14 1648 15
rect 1657 14 1667 15
rect 1678 14 1688 15
rect 1701 14 1712 15
rect 1729 14 1740 15
rect 1291 11 1300 14
rect 1303 12 1319 14
rect 1325 12 1334 14
rect 1337 13 1351 14
rect 1500 13 1508 14
rect 1542 13 1544 14
rect 1582 13 1584 14
rect 1645 13 1648 14
rect 1659 13 1665 14
rect 1338 12 1351 13
rect 1304 11 1319 12
rect 1326 11 1334 12
rect 1339 11 1351 12
rect 1250 10 1259 11
rect 1269 10 1276 11
rect 1280 10 1283 11
rect 1292 10 1299 11
rect 1305 10 1312 11
rect 1315 10 1318 11
rect 1327 10 1333 11
rect 1340 10 1350 11
<< metal3 >>
rect 510 503 524 504
rect 730 503 743 504
rect 838 503 848 504
rect 893 503 905 504
rect 505 502 531 503
rect 544 502 579 503
rect 502 501 534 502
rect 500 500 534 501
rect 498 499 534 500
rect 496 498 534 499
rect 494 497 534 498
rect 493 496 534 497
rect 492 495 534 496
rect 490 494 534 495
rect 489 492 534 494
rect 488 491 534 492
rect 487 490 534 491
rect 486 488 534 490
rect 485 487 534 488
rect 484 486 514 487
rect 525 486 534 487
rect 484 485 511 486
rect 528 485 534 486
rect 483 484 509 485
rect 531 484 534 485
rect 483 483 507 484
rect 533 483 534 484
rect 544 501 585 502
rect 544 500 588 501
rect 544 499 590 500
rect 544 498 591 499
rect 544 497 593 498
rect 544 496 594 497
rect 544 494 595 496
rect 544 493 596 494
rect 544 491 597 493
rect 544 489 598 491
rect 482 482 506 483
rect 482 480 505 482
rect 481 479 504 480
rect 481 477 503 479
rect 481 475 502 477
rect 480 473 502 475
rect 480 466 501 473
rect 544 472 564 489
rect 572 488 598 489
rect 574 487 598 488
rect 576 485 599 487
rect 577 483 599 485
rect 578 478 599 483
rect 577 476 599 478
rect 577 475 598 476
rect 576 474 598 475
rect 575 473 598 474
rect 573 472 597 473
rect 544 471 597 472
rect 544 469 596 471
rect 544 468 595 469
rect 544 466 594 468
rect 606 466 627 503
rect 480 462 502 466
rect 544 465 593 466
rect 544 464 591 465
rect 544 463 590 464
rect 544 462 589 463
rect 480 461 503 462
rect 481 460 503 461
rect 544 461 587 462
rect 544 460 585 461
rect 481 459 504 460
rect 544 459 582 460
rect 607 459 627 466
rect 645 463 666 503
rect 725 502 747 503
rect 722 501 748 502
rect 720 500 748 501
rect 718 499 748 500
rect 717 498 748 499
rect 715 497 748 498
rect 714 496 748 497
rect 713 495 748 496
rect 766 495 804 503
rect 834 502 852 503
rect 887 502 909 503
rect 831 501 855 502
rect 884 501 911 502
rect 829 500 856 501
rect 882 500 913 501
rect 828 499 858 500
rect 879 499 915 500
rect 826 498 859 499
rect 878 498 916 499
rect 825 497 860 498
rect 878 497 917 498
rect 824 496 861 497
rect 878 496 918 497
rect 824 495 862 496
rect 712 494 748 495
rect 711 492 748 494
rect 710 491 748 492
rect 709 489 748 491
rect 708 488 733 489
rect 745 488 748 489
rect 707 487 730 488
rect 765 487 804 495
rect 823 494 862 495
rect 878 494 919 496
rect 822 493 863 494
rect 821 492 863 493
rect 878 492 920 494
rect 821 491 864 492
rect 820 490 864 491
rect 820 489 865 490
rect 819 488 840 489
rect 844 488 865 489
rect 878 488 921 492
rect 1654 489 1710 490
rect 1646 488 1713 489
rect 819 487 839 488
rect 845 487 866 488
rect 707 486 728 487
rect 706 485 727 486
rect 706 484 726 485
rect 706 483 725 484
rect 705 482 725 483
rect 705 481 724 482
rect 705 480 723 481
rect 704 478 723 480
rect 731 479 740 480
rect 765 479 781 487
rect 819 486 838 487
rect 818 484 838 486
rect 846 485 866 487
rect 847 484 866 485
rect 878 487 889 488
rect 898 487 921 488
rect 1640 487 1716 488
rect 878 486 885 487
rect 900 486 922 487
rect 1636 486 1718 487
rect 878 485 883 486
rect 878 484 881 485
rect 901 484 922 486
rect 1571 485 1575 486
rect 1631 485 1720 486
rect 1567 484 1581 485
rect 1627 484 1722 485
rect 818 482 837 484
rect 728 478 743 479
rect 764 478 781 479
rect 817 479 837 482
rect 847 481 867 484
rect 878 483 879 484
rect 704 475 722 478
rect 726 477 745 478
rect 764 477 791 478
rect 725 476 746 477
rect 764 476 795 477
rect 724 475 747 476
rect 764 475 797 476
rect 817 475 836 479
rect 703 474 722 475
rect 723 474 748 475
rect 764 474 799 475
rect 703 473 749 474
rect 764 473 800 474
rect 703 471 750 473
rect 764 471 802 473
rect 703 469 751 471
rect 764 470 803 471
rect 764 469 804 470
rect 703 466 752 469
rect 703 465 726 466
rect 731 465 752 466
rect 764 466 805 469
rect 703 464 725 465
rect 732 464 753 465
rect 703 463 724 464
rect 645 459 665 463
rect 481 457 505 459
rect 544 458 577 459
rect 482 456 506 457
rect 482 455 507 456
rect 533 455 534 456
rect 482 454 509 455
rect 531 454 534 455
rect 483 453 511 454
rect 528 453 534 454
rect 483 452 514 453
rect 524 452 534 453
rect 484 450 534 452
rect 485 448 534 450
rect 486 447 534 448
rect 487 446 534 447
rect 488 445 534 446
rect 489 444 534 445
rect 490 443 534 444
rect 491 442 534 443
rect 492 441 534 442
rect 493 440 534 441
rect 495 439 534 440
rect 497 438 534 439
rect 499 437 532 438
rect 503 436 528 437
rect 544 436 564 458
rect 607 456 628 459
rect 644 456 665 459
rect 703 459 723 463
rect 733 462 753 464
rect 764 464 806 466
rect 764 463 766 464
rect 781 463 806 464
rect 816 463 836 475
rect 784 462 807 463
rect 703 457 722 459
rect 607 455 629 456
rect 643 455 665 456
rect 608 454 630 455
rect 642 454 664 455
rect 608 453 631 454
rect 641 453 664 454
rect 704 453 723 457
rect 734 454 753 462
rect 785 461 807 462
rect 786 460 807 461
rect 787 455 807 460
rect 817 459 836 463
rect 848 477 867 481
rect 902 481 922 484
rect 1565 483 1585 484
rect 1623 483 1723 484
rect 1564 482 1588 483
rect 1618 482 1725 483
rect 1562 481 1593 482
rect 1612 481 1726 482
rect 902 479 921 481
rect 1561 480 1728 481
rect 1560 479 1730 480
rect 901 477 921 479
rect 1559 478 1731 479
rect 1559 477 1732 478
rect 848 463 868 477
rect 900 476 921 477
rect 1558 476 1734 477
rect 900 475 920 476
rect 899 474 920 475
rect 1557 475 1735 476
rect 1557 474 1737 475
rect 898 473 919 474
rect 1557 473 1738 474
rect 897 472 919 473
rect 1556 472 1739 473
rect 895 471 918 472
rect 894 470 918 471
rect 1556 471 1740 472
rect 1556 470 1650 471
rect 1668 470 1742 471
rect 893 469 917 470
rect 1556 469 1585 470
rect 1589 469 1647 470
rect 1673 469 1743 470
rect 892 468 916 469
rect 1556 468 1578 469
rect 1596 468 1646 469
rect 1676 468 1744 469
rect 890 467 915 468
rect 1557 467 1575 468
rect 1600 467 1646 468
rect 1680 467 1745 468
rect 889 466 914 467
rect 1557 466 1573 467
rect 1602 466 1648 467
rect 1685 466 1746 467
rect 888 465 913 466
rect 1558 465 1572 466
rect 1604 465 1653 466
rect 1689 465 1747 466
rect 887 464 911 465
rect 1559 464 1570 465
rect 1605 464 1656 465
rect 1694 464 1748 465
rect 886 463 910 464
rect 1536 463 1541 464
rect 1561 463 1566 464
rect 1607 463 1660 464
rect 1701 463 1749 464
rect 848 459 867 463
rect 884 462 909 463
rect 1533 462 1544 463
rect 1608 462 1663 463
rect 1711 462 1750 463
rect 883 461 907 462
rect 1531 461 1547 462
rect 1608 461 1666 462
rect 1717 461 1751 462
rect 882 460 905 461
rect 1529 460 1548 461
rect 1609 460 1669 461
rect 1721 460 1752 461
rect 817 455 837 459
rect 847 456 867 459
rect 881 459 904 460
rect 1528 459 1550 460
rect 1577 459 1585 460
rect 1610 459 1672 460
rect 1725 459 1753 460
rect 881 458 903 459
rect 1527 458 1551 459
rect 1573 458 1588 459
rect 1610 458 1675 459
rect 1729 458 1754 459
rect 880 457 901 458
rect 1526 457 1552 458
rect 1571 457 1590 458
rect 1610 457 1679 458
rect 1732 457 1755 458
rect 879 456 900 457
rect 1525 456 1553 457
rect 1569 456 1592 457
rect 1611 456 1683 457
rect 1736 456 1755 457
rect 847 455 866 456
rect 879 455 899 456
rect 1524 455 1554 456
rect 1567 455 1593 456
rect 1611 455 1689 456
rect 1739 455 1756 456
rect 787 454 806 455
rect 608 452 633 453
rect 639 452 664 453
rect 705 452 724 453
rect 733 452 752 454
rect 786 453 806 454
rect 609 449 663 452
rect 705 451 725 452
rect 732 451 752 452
rect 705 450 726 451
rect 731 450 752 451
rect 762 452 763 453
rect 785 452 806 453
rect 762 451 766 452
rect 784 451 806 452
rect 818 454 837 455
rect 818 452 838 454
rect 846 452 866 455
rect 878 454 898 455
rect 1523 454 1555 455
rect 1565 454 1594 455
rect 1611 454 1706 455
rect 1742 454 1757 455
rect 877 453 897 454
rect 1523 453 1557 454
rect 1563 453 1595 454
rect 1611 453 1711 454
rect 1744 453 1757 454
rect 877 452 896 453
rect 1522 452 1595 453
rect 1610 452 1715 453
rect 1747 452 1758 453
rect 818 451 839 452
rect 845 451 865 452
rect 877 451 922 452
rect 762 450 770 451
rect 781 450 806 451
rect 819 450 840 451
rect 844 450 865 451
rect 610 447 662 449
rect 706 448 751 450
rect 762 448 805 450
rect 819 449 864 450
rect 820 448 864 449
rect 611 446 661 447
rect 707 446 750 448
rect 762 446 804 448
rect 820 447 863 448
rect 876 447 922 451
rect 1521 450 1596 452
rect 1520 449 1596 450
rect 1610 451 1718 452
rect 1750 451 1758 452
rect 1610 450 1721 451
rect 1752 450 1758 451
rect 1610 449 1724 450
rect 1754 449 1759 450
rect 1519 447 1596 449
rect 1609 448 1727 449
rect 1756 448 1759 449
rect 1609 447 1730 448
rect 1758 447 1759 448
rect 821 446 863 447
rect 612 444 660 446
rect 708 445 749 446
rect 762 445 803 446
rect 821 445 862 446
rect 708 444 748 445
rect 613 443 659 444
rect 709 443 748 444
rect 762 443 802 445
rect 822 444 862 445
rect 822 443 861 444
rect 614 442 658 443
rect 710 442 747 443
rect 762 442 801 443
rect 823 442 860 443
rect 615 441 657 442
rect 711 441 746 442
rect 762 441 800 442
rect 824 441 859 442
rect 616 440 656 441
rect 712 440 745 441
rect 762 440 798 441
rect 825 440 858 441
rect 618 439 654 440
rect 713 439 743 440
rect 762 439 797 440
rect 826 439 857 440
rect 620 438 652 439
rect 715 438 742 439
rect 762 438 795 439
rect 828 438 855 439
rect 622 437 650 438
rect 717 437 740 438
rect 762 437 793 438
rect 830 437 854 438
rect 624 436 647 437
rect 719 436 737 437
rect 766 436 790 437
rect 832 436 851 437
rect 875 436 922 447
rect 1518 446 1596 447
rect 1517 445 1596 446
rect 1608 446 1733 447
rect 1608 445 1736 446
rect 1516 444 1596 445
rect 1607 444 1739 445
rect 1515 443 1595 444
rect 1514 442 1595 443
rect 1607 443 1741 444
rect 1607 442 1744 443
rect 1513 441 1594 442
rect 1608 441 1747 442
rect 1512 440 1594 441
rect 1610 440 1749 441
rect 1511 439 1593 440
rect 1612 439 1752 440
rect 1510 438 1592 439
rect 1613 438 1754 439
rect 1509 437 1591 438
rect 1615 437 1668 438
rect 1671 437 1757 438
rect 1508 436 1590 437
rect 1616 436 1668 437
rect 1675 436 1759 437
rect 508 435 522 436
rect 629 435 642 436
rect 723 435 733 436
rect 773 435 786 436
rect 836 435 847 436
rect 1507 435 1589 436
rect 1618 435 1668 436
rect 1677 435 1761 436
rect 1505 434 1587 435
rect 1619 434 1669 435
rect 1680 434 1764 435
rect 1504 433 1544 434
rect 1549 433 1586 434
rect 1621 433 1669 434
rect 1682 433 1765 434
rect 1502 432 1539 433
rect 1548 432 1585 433
rect 1622 432 1669 433
rect 1685 432 1766 433
rect 1501 431 1535 432
rect 1546 431 1584 432
rect 1623 431 1669 432
rect 1687 431 1768 432
rect 1499 430 1532 431
rect 1545 430 1583 431
rect 1625 430 1669 431
rect 1689 430 1768 431
rect 1498 429 1528 430
rect 1543 429 1582 430
rect 1626 429 1670 430
rect 1692 429 1769 430
rect 1496 428 1525 429
rect 1542 428 1581 429
rect 1627 428 1670 429
rect 1694 428 1770 429
rect 1494 427 1523 428
rect 1540 427 1580 428
rect 1628 427 1671 428
rect 1697 427 1771 428
rect 1493 426 1521 427
rect 1538 426 1580 427
rect 1629 426 1671 427
rect 1699 426 1771 427
rect 1491 425 1520 426
rect 1536 425 1579 426
rect 1630 425 1672 426
rect 1703 425 1772 426
rect 1489 424 1518 425
rect 1535 424 1579 425
rect 1631 424 1673 425
rect 1707 424 1772 425
rect 1487 423 1516 424
rect 1533 423 1578 424
rect 1485 422 1514 423
rect 1532 422 1578 423
rect 1594 423 1597 424
rect 1604 423 1607 424
rect 1632 423 1674 424
rect 1713 423 1773 424
rect 1594 422 1612 423
rect 1633 422 1675 423
rect 1717 422 1773 423
rect 1483 421 1513 422
rect 1480 420 1512 421
rect 1531 420 1578 422
rect 1595 421 1615 422
rect 1634 421 1676 422
rect 1720 421 1774 422
rect 1595 420 1616 421
rect 1635 420 1678 421
rect 1722 420 1774 421
rect 1478 419 1511 420
rect 1518 419 1520 420
rect 1530 419 1579 420
rect 1477 418 1511 419
rect 1513 418 1520 419
rect 1529 418 1579 419
rect 1475 417 1520 418
rect 1473 416 1520 417
rect 1528 416 1579 418
rect 1596 419 1618 420
rect 1636 419 1679 420
rect 1725 419 1775 420
rect 1596 418 1619 419
rect 1637 418 1681 419
rect 1727 418 1775 419
rect 1596 417 1620 418
rect 1637 417 1683 418
rect 1729 417 1775 418
rect 1472 415 1521 416
rect 1470 414 1521 415
rect 1527 415 1579 416
rect 1597 415 1621 417
rect 1638 416 1685 417
rect 1731 416 1776 417
rect 1639 415 1687 416
rect 1733 415 1776 416
rect 1527 414 1580 415
rect 1469 413 1521 414
rect 1468 412 1522 413
rect 1526 412 1580 414
rect 1467 411 1523 412
rect 1525 411 1580 412
rect 1598 414 1622 415
rect 1640 414 1689 415
rect 1735 414 1776 415
rect 1598 412 1623 414
rect 1640 413 1692 414
rect 1736 413 1776 414
rect 1641 412 1696 413
rect 1738 412 1777 413
rect 1598 411 1624 412
rect 1642 411 1699 412
rect 1740 411 1777 412
rect 1466 410 1581 411
rect 1465 409 1581 410
rect 1464 407 1581 409
rect 1463 405 1581 407
rect 1599 409 1625 411
rect 1642 410 1703 411
rect 1741 410 1777 411
rect 1643 409 1707 410
rect 1743 409 1777 410
rect 1599 407 1626 409
rect 1644 408 1712 409
rect 1744 408 1778 409
rect 1644 407 1716 408
rect 1746 407 1778 408
rect 1599 405 1627 407
rect 1645 406 1719 407
rect 1747 406 1778 407
rect 1645 405 1721 406
rect 1748 405 1778 406
rect 1463 403 1582 405
rect 1463 402 1483 403
rect 1484 402 1582 403
rect 504 399 511 400
rect 526 399 533 400
rect 547 399 554 400
rect 501 398 513 399
rect 524 398 535 399
rect 544 398 556 399
rect 573 398 579 400
rect 500 397 514 398
rect 523 397 536 398
rect 500 396 515 397
rect 500 395 505 396
rect 507 395 515 396
rect 522 396 536 397
rect 543 397 557 398
rect 543 396 558 397
rect 572 396 579 398
rect 522 395 528 396
rect 530 395 537 396
rect 500 394 502 395
rect 509 394 515 395
rect 521 394 527 395
rect 531 394 537 395
rect 543 395 548 396
rect 550 395 558 396
rect 571 395 579 396
rect 543 394 545 395
rect 552 394 558 395
rect 510 391 516 394
rect 521 393 526 394
rect 510 390 515 391
rect 509 389 515 390
rect 508 388 515 389
rect 520 390 526 393
rect 532 391 538 394
rect 507 387 514 388
rect 506 386 513 387
rect 505 385 512 386
rect 503 384 511 385
rect 520 384 525 390
rect 502 383 510 384
rect 501 382 508 383
rect 500 381 507 382
rect 520 381 526 384
rect 533 383 538 391
rect 553 391 559 394
rect 570 393 579 395
rect 569 392 579 393
rect 568 391 573 392
rect 553 390 558 391
rect 568 390 572 391
rect 552 389 558 390
rect 567 389 572 390
rect 551 388 558 389
rect 566 388 571 389
rect 550 387 557 388
rect 566 387 570 388
rect 549 386 556 387
rect 565 386 570 387
rect 548 385 555 386
rect 564 385 569 386
rect 546 384 554 385
rect 563 384 568 385
rect 574 384 579 392
rect 545 383 553 384
rect 562 383 568 384
rect 573 383 579 384
rect 500 380 506 381
rect 521 380 526 381
rect 532 380 538 383
rect 544 382 551 383
rect 543 381 550 382
rect 543 380 549 381
rect 499 379 505 380
rect 521 379 527 380
rect 531 379 537 380
rect 499 374 516 379
rect 521 378 528 379
rect 530 378 537 379
rect 542 379 548 380
rect 562 379 582 383
rect 611 381 617 400
rect 691 399 696 400
rect 715 399 720 400
rect 740 399 749 400
rect 691 398 695 399
rect 716 398 721 399
rect 737 398 751 399
rect 690 397 695 398
rect 689 395 694 397
rect 717 396 722 398
rect 735 397 751 398
rect 734 396 751 397
rect 688 393 693 395
rect 718 394 723 396
rect 733 395 751 396
rect 732 394 741 395
rect 749 394 751 395
rect 626 392 633 393
rect 623 391 635 392
rect 623 390 636 391
rect 643 390 648 393
rect 652 392 657 393
rect 650 391 658 392
rect 649 390 659 391
rect 687 390 692 393
rect 705 392 712 393
rect 719 392 724 394
rect 732 393 739 394
rect 703 391 713 392
rect 701 390 713 391
rect 623 389 637 390
rect 623 388 626 389
rect 632 388 637 389
rect 643 389 660 390
rect 687 389 691 390
rect 700 389 713 390
rect 643 388 651 389
rect 652 388 660 389
rect 623 387 624 388
rect 632 386 638 388
rect 627 385 638 386
rect 624 384 638 385
rect 623 383 638 384
rect 622 382 628 383
rect 621 381 627 382
rect 633 381 638 383
rect 610 380 616 381
rect 604 379 605 380
rect 609 379 616 380
rect 522 377 536 378
rect 523 376 535 377
rect 524 375 534 376
rect 526 374 532 375
rect 542 374 559 379
rect 574 374 579 379
rect 604 378 616 379
rect 621 379 626 381
rect 632 379 638 381
rect 621 378 627 379
rect 631 378 638 379
rect 585 377 591 378
rect 604 377 615 378
rect 621 377 638 378
rect 585 374 590 377
rect 604 376 614 377
rect 622 376 638 377
rect 604 375 613 376
rect 623 375 631 376
rect 604 374 611 375
rect 624 374 629 375
rect 633 374 638 376
rect 643 387 649 388
rect 643 374 648 387
rect 654 386 660 388
rect 655 374 660 386
rect 666 379 669 380
rect 665 378 670 379
rect 686 378 691 389
rect 699 388 708 389
rect 710 388 713 389
rect 720 391 724 392
rect 731 392 738 393
rect 763 392 770 393
rect 785 392 793 393
rect 808 392 813 393
rect 731 391 737 392
rect 760 391 772 392
rect 783 391 795 392
rect 806 391 815 392
rect 816 391 821 402
rect 699 386 705 388
rect 720 387 725 391
rect 698 380 704 386
rect 721 381 725 387
rect 730 390 737 391
rect 759 390 774 391
rect 782 390 796 391
rect 805 390 821 391
rect 730 384 736 390
rect 758 389 774 390
rect 781 389 797 390
rect 804 389 821 390
rect 742 384 753 389
rect 758 388 765 389
rect 768 388 775 389
rect 780 388 788 389
rect 790 388 798 389
rect 757 386 763 388
rect 769 387 776 388
rect 780 387 786 388
rect 792 387 798 388
rect 803 388 811 389
rect 813 388 821 389
rect 803 387 809 388
rect 757 385 762 386
rect 770 385 776 387
rect 730 382 737 384
rect 699 379 705 380
rect 699 378 707 379
rect 710 378 713 379
rect 664 376 671 378
rect 665 375 670 376
rect 687 375 692 378
rect 700 377 713 378
rect 701 376 713 377
rect 720 376 725 381
rect 731 381 738 382
rect 731 380 739 381
rect 732 379 740 380
rect 747 379 753 384
rect 756 382 762 385
rect 771 382 776 385
rect 757 381 762 382
rect 757 379 763 381
rect 770 380 776 382
rect 779 380 785 387
rect 793 381 799 387
rect 793 380 798 381
rect 802 380 808 387
rect 815 386 821 388
rect 816 382 821 386
rect 815 380 821 382
rect 769 379 775 380
rect 732 378 753 379
rect 733 377 753 378
rect 758 378 765 379
rect 768 378 775 379
rect 780 379 786 380
rect 792 379 798 380
rect 780 378 788 379
rect 790 378 798 379
rect 803 379 809 380
rect 814 379 821 380
rect 803 378 811 379
rect 813 378 821 379
rect 758 377 774 378
rect 781 377 797 378
rect 803 377 821 378
rect 735 376 753 377
rect 759 376 773 377
rect 782 376 796 377
rect 804 376 821 377
rect 702 375 713 376
rect 666 374 669 375
rect 585 373 589 374
rect 688 373 693 375
rect 704 374 712 375
rect 719 374 724 376
rect 736 375 751 376
rect 760 375 772 376
rect 783 375 795 376
rect 805 375 814 376
rect 739 374 748 375
rect 763 374 770 375
rect 785 374 793 375
rect 807 374 812 375
rect 816 374 821 376
rect 827 389 832 400
rect 840 399 847 400
rect 840 398 846 399
rect 839 397 846 398
rect 838 396 845 397
rect 838 395 844 396
rect 837 394 843 395
rect 836 393 843 394
rect 836 392 842 393
rect 856 392 863 393
rect 878 392 886 393
rect 835 391 841 392
rect 853 391 865 392
rect 876 391 888 392
rect 834 390 841 391
rect 852 390 867 391
rect 875 390 889 391
rect 834 389 840 390
rect 851 389 867 390
rect 874 389 890 390
rect 827 386 839 389
rect 851 388 858 389
rect 861 388 868 389
rect 873 388 881 389
rect 883 388 891 389
rect 850 386 856 388
rect 862 387 869 388
rect 873 387 879 388
rect 885 387 891 388
rect 827 374 832 386
rect 833 385 840 386
rect 850 385 855 386
rect 863 385 869 387
rect 834 384 841 385
rect 835 383 841 384
rect 835 382 842 383
rect 849 382 855 385
rect 864 382 869 385
rect 836 381 843 382
rect 850 381 855 382
rect 837 379 844 381
rect 850 379 856 381
rect 863 380 869 382
rect 872 380 878 387
rect 886 381 892 387
rect 896 385 902 402
rect 1463 401 1481 402
rect 1483 401 1582 402
rect 1464 400 1479 401
rect 1482 400 1582 401
rect 1464 399 1477 400
rect 1481 399 1582 400
rect 1465 398 1474 399
rect 1480 398 1582 399
rect 1467 397 1470 398
rect 1479 397 1582 398
rect 1478 396 1582 397
rect 1477 395 1582 396
rect 1599 403 1628 405
rect 1646 404 1723 405
rect 1750 404 1778 405
rect 1646 403 1725 404
rect 1751 403 1778 404
rect 1599 400 1629 403
rect 1647 402 1726 403
rect 1752 402 1778 403
rect 1647 401 1728 402
rect 1753 401 1779 402
rect 1647 400 1730 401
rect 1755 400 1779 401
rect 1599 398 1630 400
rect 1648 399 1731 400
rect 1756 399 1779 400
rect 1648 398 1733 399
rect 1757 398 1779 399
rect 1599 396 1631 398
rect 1649 397 1734 398
rect 1758 397 1779 398
rect 1649 396 1735 397
rect 1759 396 1779 397
rect 1476 394 1581 395
rect 1599 394 1632 396
rect 1650 395 1737 396
rect 1760 395 1779 396
rect 1651 394 1738 395
rect 1761 394 1779 395
rect 1475 393 1581 394
rect 907 392 914 393
rect 1474 392 1581 393
rect 907 391 913 392
rect 1473 391 1581 392
rect 1598 392 1633 394
rect 1651 393 1739 394
rect 1762 393 1779 394
rect 1652 392 1741 393
rect 1763 392 1779 393
rect 906 390 912 391
rect 905 389 912 390
rect 1472 389 1580 391
rect 1598 390 1634 392
rect 1653 391 1742 392
rect 1764 391 1779 392
rect 1654 390 1743 391
rect 1598 389 1635 390
rect 1655 389 1744 390
rect 1765 389 1779 391
rect 905 388 911 389
rect 1471 388 1580 389
rect 904 387 910 388
rect 903 385 909 387
rect 1471 386 1579 388
rect 1597 387 1636 389
rect 1656 388 1746 389
rect 1766 388 1779 389
rect 1658 387 1747 388
rect 1767 387 1779 388
rect 1597 386 1637 387
rect 1660 386 1748 387
rect 1470 385 1578 386
rect 896 383 908 385
rect 1471 384 1578 385
rect 1596 384 1638 386
rect 1662 385 1749 386
rect 1768 385 1778 387
rect 1664 384 1750 385
rect 1769 384 1778 385
rect 1471 383 1577 384
rect 1596 383 1639 384
rect 1668 383 1751 384
rect 896 382 909 383
rect 1471 382 1576 383
rect 1596 382 1640 383
rect 1673 382 1752 383
rect 1770 382 1778 384
rect 886 380 891 381
rect 862 379 868 380
rect 838 378 845 379
rect 851 378 858 379
rect 861 378 868 379
rect 873 379 879 380
rect 885 379 891 380
rect 873 378 881 379
rect 883 378 891 379
rect 839 376 846 378
rect 851 377 867 378
rect 874 377 890 378
rect 852 376 866 377
rect 875 376 889 377
rect 840 375 847 376
rect 853 375 865 376
rect 876 375 888 376
rect 841 374 848 375
rect 856 374 863 375
rect 878 374 886 375
rect 896 374 902 382
rect 903 381 909 382
rect 1472 381 1576 382
rect 1595 381 1641 382
rect 1679 381 1753 382
rect 1771 381 1778 382
rect 904 380 910 381
rect 1472 380 1575 381
rect 1595 380 1643 381
rect 1685 380 1754 381
rect 904 379 911 380
rect 905 378 912 379
rect 1473 378 1574 380
rect 1594 379 1644 380
rect 1690 379 1755 380
rect 1772 379 1777 381
rect 1594 378 1646 379
rect 1693 378 1756 379
rect 1773 378 1777 379
rect 906 377 912 378
rect 1474 377 1573 378
rect 1594 377 1647 378
rect 1696 377 1757 378
rect 1773 377 1776 378
rect 906 376 913 377
rect 1474 376 1519 377
rect 1521 376 1572 377
rect 907 375 914 376
rect 1475 375 1517 376
rect 1523 375 1572 376
rect 1593 376 1649 377
rect 1699 376 1757 377
rect 1774 376 1776 377
rect 1593 375 1652 376
rect 1702 375 1758 376
rect 1774 375 1775 376
rect 908 374 914 375
rect 1476 374 1516 375
rect 1524 374 1571 375
rect 1592 374 1655 375
rect 1704 374 1759 375
rect 584 371 589 373
rect 689 372 693 373
rect 718 372 723 374
rect 1477 373 1515 374
rect 1525 373 1570 374
rect 1592 373 1659 374
rect 1707 373 1759 374
rect 1478 372 1514 373
rect 1525 372 1569 373
rect 1592 372 1664 373
rect 1709 372 1759 373
rect 689 371 694 372
rect 584 369 588 371
rect 690 369 695 371
rect 717 370 722 372
rect 1479 371 1513 372
rect 1526 371 1569 372
rect 1591 371 1669 372
rect 1712 371 1760 372
rect 1480 370 1510 371
rect 1526 370 1568 371
rect 1591 370 1675 371
rect 1715 370 1760 371
rect 716 369 721 370
rect 1481 369 1506 370
rect 1525 369 1568 370
rect 1590 369 1679 370
rect 1717 369 1760 370
rect 691 368 696 369
rect 715 368 720 369
rect 1483 368 1498 369
rect 1525 368 1567 369
rect 1590 368 1683 369
rect 1719 368 1761 369
rect 1488 367 1489 368
rect 1523 367 1566 368
rect 1520 366 1566 367
rect 1589 367 1685 368
rect 1720 367 1761 368
rect 1589 366 1688 367
rect 1722 366 1761 367
rect 1517 365 1565 366
rect 1588 365 1691 366
rect 1723 365 1761 366
rect 1513 364 1565 365
rect 1587 364 1693 365
rect 1724 364 1761 365
rect 1507 363 1564 364
rect 1587 363 1695 364
rect 1725 363 1762 364
rect 1498 362 1563 363
rect 1488 361 1563 362
rect 1586 362 1697 363
rect 1726 362 1762 363
rect 1586 361 1699 362
rect 1727 361 1762 362
rect 1486 360 1562 361
rect 1585 360 1701 361
rect 1728 360 1762 361
rect 1486 359 1561 360
rect 1485 358 1561 359
rect 1584 359 1703 360
rect 1729 359 1762 360
rect 1584 358 1704 359
rect 1730 358 1762 359
rect 1485 357 1560 358
rect 1583 357 1706 358
rect 1485 356 1559 357
rect 1582 356 1707 357
rect 1731 356 1762 358
rect 1485 355 1558 356
rect 1581 355 1708 356
rect 1732 355 1762 356
rect 1485 354 1557 355
rect 1581 354 1709 355
rect 1733 354 1762 355
rect 1485 353 1556 354
rect 1580 353 1710 354
rect 1486 352 1555 353
rect 1579 352 1711 353
rect 1734 352 1762 354
rect 1486 351 1554 352
rect 1578 351 1712 352
rect 1486 350 1553 351
rect 1577 350 1713 351
rect 1735 350 1762 352
rect 1487 349 1552 350
rect 1576 349 1714 350
rect 1736 349 1762 350
rect 475 348 696 349
rect 736 348 962 349
rect 998 348 1206 349
rect 1287 348 1354 349
rect 1487 348 1550 349
rect 1576 348 1715 349
rect 474 313 697 348
rect 736 347 963 348
rect 997 347 1212 348
rect 1287 347 1355 348
rect 735 313 964 347
rect 997 346 1215 347
rect 996 345 1217 346
rect 997 344 1219 345
rect 997 343 1221 344
rect 997 342 1222 343
rect 997 341 1224 342
rect 997 340 1225 341
rect 997 339 1226 340
rect 997 338 1227 339
rect 997 337 1228 338
rect 997 335 1229 337
rect 997 334 1230 335
rect 997 332 1231 334
rect 997 330 1232 332
rect 997 328 1233 330
rect 997 325 1234 328
rect 997 319 1235 325
rect 474 312 696 313
rect 736 312 963 313
rect 997 312 1236 319
rect 474 311 544 312
rect 815 311 885 312
rect 474 283 543 311
rect 474 282 544 283
rect 474 281 695 282
rect 474 280 696 281
rect 474 246 697 280
rect 474 245 696 246
rect 474 244 545 245
rect 547 244 549 245
rect 693 244 694 245
rect 474 243 544 244
rect 474 215 543 243
rect 474 214 544 215
rect 474 213 696 214
rect 474 205 697 213
rect 475 201 697 205
rect 476 198 697 201
rect 477 196 697 198
rect 478 194 697 196
rect 479 192 697 194
rect 480 191 697 192
rect 481 190 697 191
rect 482 188 697 190
rect 483 187 697 188
rect 484 186 697 187
rect 485 185 697 186
rect 486 184 697 185
rect 488 183 697 184
rect 489 182 697 183
rect 491 181 697 182
rect 493 180 697 181
rect 496 179 697 180
rect 498 178 697 179
rect 815 178 884 311
rect 997 181 1066 312
rect 1167 258 1236 312
rect 1089 257 1091 258
rect 1093 257 1163 258
rect 1164 257 1235 258
rect 1088 256 1170 257
rect 1089 255 1170 256
rect 1090 254 1170 255
rect 1091 253 1172 254
rect 1092 252 1173 253
rect 1093 251 1174 252
rect 1094 250 1174 251
rect 1095 249 1176 250
rect 1096 248 1177 249
rect 1097 247 1178 248
rect 1098 246 1179 247
rect 1099 245 1180 246
rect 1100 244 1181 245
rect 1101 243 1182 244
rect 1102 242 1183 243
rect 1103 241 1184 242
rect 1104 240 1185 241
rect 1105 239 1186 240
rect 1106 238 1187 239
rect 1107 237 1188 238
rect 1108 236 1189 237
rect 1109 235 1190 236
rect 1110 234 1191 235
rect 1111 233 1192 234
rect 1112 232 1193 233
rect 1113 231 1194 232
rect 1114 230 1195 231
rect 1115 229 1196 230
rect 1116 228 1197 229
rect 1117 227 1198 228
rect 1118 226 1199 227
rect 1119 225 1200 226
rect 1120 224 1201 225
rect 1121 223 1202 224
rect 1122 222 1203 223
rect 1123 221 1204 222
rect 1124 220 1205 221
rect 1125 219 1206 220
rect 1126 218 1207 219
rect 1127 217 1208 218
rect 1128 216 1209 217
rect 1129 215 1210 216
rect 1130 214 1211 215
rect 1131 213 1212 214
rect 1132 212 1213 213
rect 1133 211 1214 212
rect 1134 210 1215 211
rect 1135 209 1216 210
rect 1136 208 1217 209
rect 1137 207 1218 208
rect 1138 206 1219 207
rect 1139 205 1220 206
rect 1140 204 1221 205
rect 1141 203 1222 204
rect 1142 202 1223 203
rect 1143 201 1224 202
rect 1144 200 1225 201
rect 1145 199 1227 200
rect 1146 198 1227 199
rect 1147 197 1229 198
rect 1148 196 1229 197
rect 1149 195 1231 196
rect 1150 194 1231 195
rect 1151 193 1233 194
rect 1152 192 1233 193
rect 1153 191 1235 192
rect 1154 190 1235 191
rect 1155 189 1237 190
rect 1156 188 1237 189
rect 1157 187 1239 188
rect 1158 186 1239 187
rect 1159 185 1241 186
rect 1160 184 1241 185
rect 1161 183 1243 184
rect 1162 182 1243 183
rect 1163 181 1245 182
rect 996 179 1066 181
rect 1164 180 1245 181
rect 1165 179 1247 180
rect 1286 179 1355 347
rect 1488 347 1549 348
rect 1575 347 1635 348
rect 1644 347 1715 348
rect 1737 347 1762 349
rect 1488 346 1547 347
rect 1574 346 1633 347
rect 1648 346 1716 347
rect 1489 345 1545 346
rect 1572 345 1632 346
rect 1650 345 1717 346
rect 1738 345 1762 347
rect 1490 344 1543 345
rect 1571 344 1631 345
rect 1652 344 1717 345
rect 1490 343 1541 344
rect 1570 343 1630 344
rect 1654 343 1718 344
rect 1739 343 1762 345
rect 1491 342 1539 343
rect 1569 342 1629 343
rect 1655 342 1718 343
rect 1740 342 1762 343
rect 1492 341 1537 342
rect 1568 341 1629 342
rect 1657 341 1719 342
rect 1740 341 1761 342
rect 1492 340 1534 341
rect 1566 340 1628 341
rect 1658 340 1719 341
rect 1493 339 1531 340
rect 1565 339 1628 340
rect 1659 339 1720 340
rect 1741 339 1761 341
rect 1493 338 1528 339
rect 1564 338 1627 339
rect 1660 338 1720 339
rect 1494 337 1526 338
rect 1562 337 1627 338
rect 1661 337 1720 338
rect 1494 336 1522 337
rect 1560 336 1627 337
rect 1662 336 1721 337
rect 1742 336 1761 339
rect 1494 335 1519 336
rect 1559 335 1626 336
rect 1663 335 1721 336
rect 1495 334 1516 335
rect 1557 334 1626 335
rect 1664 334 1721 335
rect 1743 334 1760 336
rect 1495 333 1513 334
rect 1555 333 1626 334
rect 1665 333 1721 334
rect 1496 332 1510 333
rect 1553 332 1625 333
rect 1666 332 1721 333
rect 1496 331 1507 332
rect 1551 331 1625 332
rect 1667 331 1721 332
rect 1744 332 1760 334
rect 1744 331 1759 332
rect 1497 330 1504 331
rect 1549 330 1625 331
rect 1642 330 1644 331
rect 1667 330 1722 331
rect 1547 329 1624 330
rect 1642 329 1645 330
rect 1544 328 1624 329
rect 1542 327 1624 328
rect 1641 328 1646 329
rect 1668 328 1722 330
rect 1745 329 1759 331
rect 1745 328 1758 329
rect 1540 326 1623 327
rect 1641 326 1647 328
rect 1669 326 1721 328
rect 1537 325 1623 326
rect 1640 325 1648 326
rect 1535 324 1622 325
rect 1640 324 1649 325
rect 1670 324 1721 326
rect 1746 326 1758 328
rect 1746 325 1757 326
rect 1533 323 1622 324
rect 1639 323 1649 324
rect 1530 322 1621 323
rect 1639 322 1650 323
rect 1671 322 1721 324
rect 1747 324 1757 325
rect 1747 322 1756 324
rect 1528 321 1621 322
rect 1526 320 1620 321
rect 1638 320 1651 322
rect 1524 319 1620 320
rect 1522 318 1619 319
rect 1637 318 1652 320
rect 1672 319 1720 322
rect 1748 320 1755 322
rect 1520 317 1619 318
rect 1636 317 1653 318
rect 1673 317 1719 319
rect 1748 318 1754 320
rect 1749 317 1753 318
rect 1519 316 1618 317
rect 1636 316 1654 317
rect 1517 315 1618 316
rect 1516 314 1617 315
rect 1635 314 1654 316
rect 1673 315 1718 317
rect 1749 316 1752 317
rect 1749 315 1751 316
rect 1674 314 1717 315
rect 1749 314 1750 315
rect 1514 313 1617 314
rect 1513 312 1616 313
rect 1634 312 1655 314
rect 1674 312 1716 314
rect 1512 311 1615 312
rect 1511 310 1615 311
rect 1633 310 1656 312
rect 1674 311 1715 312
rect 1510 309 1614 310
rect 1632 309 1656 310
rect 1675 310 1714 311
rect 1509 308 1613 309
rect 1508 307 1612 308
rect 1632 307 1657 309
rect 1675 308 1713 310
rect 1675 307 1712 308
rect 1507 306 1611 307
rect 1506 305 1611 306
rect 1631 306 1657 307
rect 1676 306 1711 307
rect 1631 305 1658 306
rect 1506 304 1610 305
rect 1505 303 1609 304
rect 1630 303 1658 305
rect 1504 302 1608 303
rect 1629 302 1658 303
rect 1676 305 1710 306
rect 1676 304 1709 305
rect 1676 303 1708 304
rect 1676 302 1707 303
rect 1734 302 1735 303
rect 1504 301 1607 302
rect 1629 301 1659 302
rect 1503 300 1606 301
rect 1628 300 1659 301
rect 1676 301 1706 302
rect 1733 301 1735 302
rect 1676 300 1704 301
rect 1732 300 1735 301
rect 1503 299 1605 300
rect 1502 298 1604 299
rect 1627 298 1659 300
rect 1502 297 1603 298
rect 1626 297 1659 298
rect 1677 299 1703 300
rect 1731 299 1736 300
rect 1677 298 1702 299
rect 1730 298 1736 299
rect 1677 297 1700 298
rect 1729 297 1736 298
rect 1501 296 1602 297
rect 1501 295 1601 296
rect 1625 295 1660 297
rect 1500 294 1600 295
rect 1624 294 1660 295
rect 1500 293 1599 294
rect 1623 293 1660 294
rect 1499 292 1598 293
rect 1499 291 1597 292
rect 1622 291 1660 293
rect 1677 296 1699 297
rect 1728 296 1736 297
rect 1677 295 1697 296
rect 1727 295 1736 296
rect 1677 294 1696 295
rect 1726 294 1736 295
rect 1677 293 1694 294
rect 1725 293 1736 294
rect 1677 292 1692 293
rect 1724 292 1737 293
rect 1677 291 1691 292
rect 1723 291 1737 292
rect 1499 290 1595 291
rect 1621 290 1660 291
rect 1499 289 1594 290
rect 1620 289 1660 290
rect 1498 288 1593 289
rect 1619 288 1660 289
rect 1498 287 1591 288
rect 1618 287 1660 288
rect 1498 286 1590 287
rect 1617 286 1660 287
rect 1498 285 1588 286
rect 1616 285 1660 286
rect 1676 290 1689 291
rect 1722 290 1737 291
rect 1676 289 1687 290
rect 1720 289 1737 290
rect 1676 288 1685 289
rect 1719 288 1737 289
rect 1676 287 1682 288
rect 1718 287 1737 288
rect 1676 286 1680 287
rect 1717 286 1737 287
rect 1676 285 1677 286
rect 1715 285 1737 286
rect 1498 284 1587 285
rect 1615 284 1660 285
rect 1714 284 1737 285
rect 1497 283 1585 284
rect 1614 283 1660 284
rect 1712 283 1737 284
rect 1497 282 1583 283
rect 1612 282 1660 283
rect 1711 282 1737 283
rect 1497 281 1581 282
rect 1611 281 1660 282
rect 1709 281 1737 282
rect 1497 280 1579 281
rect 1610 280 1660 281
rect 1708 280 1737 281
rect 1497 279 1578 280
rect 1609 279 1660 280
rect 1706 279 1737 280
rect 1497 278 1575 279
rect 1607 278 1660 279
rect 1705 278 1737 279
rect 1497 277 1573 278
rect 1606 277 1659 278
rect 1703 277 1737 278
rect 1497 276 1571 277
rect 1604 276 1659 277
rect 1701 276 1737 277
rect 1497 275 1569 276
rect 1603 275 1659 276
rect 1699 275 1737 276
rect 1497 274 1567 275
rect 1601 274 1659 275
rect 1698 274 1737 275
rect 1497 273 1564 274
rect 1599 273 1659 274
rect 1696 273 1737 274
rect 1497 272 1562 273
rect 1598 272 1659 273
rect 1694 272 1736 273
rect 1497 271 1560 272
rect 1596 271 1658 272
rect 1692 271 1736 272
rect 1497 270 1557 271
rect 1594 270 1658 271
rect 1689 270 1736 271
rect 1497 269 1555 270
rect 1592 269 1658 270
rect 1687 269 1736 270
rect 1497 268 1553 269
rect 1590 268 1658 269
rect 1685 268 1736 269
rect 1497 267 1551 268
rect 1588 267 1657 268
rect 1682 267 1736 268
rect 1498 266 1549 267
rect 1586 266 1657 267
rect 1680 266 1736 267
rect 1498 265 1548 266
rect 1585 265 1657 266
rect 1677 265 1735 266
rect 1498 264 1546 265
rect 1583 264 1657 265
rect 1674 264 1735 265
rect 1498 263 1545 264
rect 1581 263 1656 264
rect 1671 263 1735 264
rect 1498 262 1544 263
rect 1579 262 1656 263
rect 1667 262 1735 263
rect 1498 261 1542 262
rect 1577 261 1656 262
rect 1663 261 1734 262
rect 1499 260 1541 261
rect 1575 260 1734 261
rect 1499 259 1540 260
rect 1573 259 1734 260
rect 1499 258 1539 259
rect 1572 258 1734 259
rect 1499 257 1538 258
rect 1570 257 1733 258
rect 1500 255 1537 257
rect 1568 256 1733 257
rect 1567 255 1733 256
rect 1500 254 1536 255
rect 1565 254 1732 255
rect 1501 252 1535 254
rect 1564 253 1732 254
rect 1562 252 1732 253
rect 1501 251 1534 252
rect 1561 251 1731 252
rect 1502 250 1534 251
rect 1560 250 1731 251
rect 1502 249 1533 250
rect 1558 249 1730 250
rect 1503 248 1533 249
rect 1557 248 1730 249
rect 1503 246 1532 248
rect 1556 247 1730 248
rect 1555 246 1729 247
rect 1504 244 1531 246
rect 1554 245 1620 246
rect 1621 245 1729 246
rect 1553 244 1618 245
rect 1505 243 1531 244
rect 1552 243 1617 244
rect 1621 243 1728 245
rect 1505 242 1530 243
rect 1551 242 1615 243
rect 1621 242 1727 243
rect 1506 240 1530 242
rect 1550 241 1613 242
rect 1620 241 1727 242
rect 1550 240 1612 241
rect 1620 240 1726 241
rect 1507 239 1530 240
rect 1549 239 1610 240
rect 1619 239 1726 240
rect 1507 238 1529 239
rect 1548 238 1609 239
rect 1619 238 1725 239
rect 1508 237 1529 238
rect 1509 235 1529 237
rect 1547 237 1607 238
rect 1547 236 1605 237
rect 1618 236 1724 238
rect 1546 235 1604 236
rect 1617 235 1723 236
rect 1510 233 1528 235
rect 1545 234 1602 235
rect 1616 234 1723 235
rect 1545 233 1601 234
rect 1616 233 1722 234
rect 1511 232 1528 233
rect 1512 230 1528 232
rect 1544 232 1599 233
rect 1615 232 1721 233
rect 1544 231 1598 232
rect 1614 231 1721 232
rect 1513 229 1528 230
rect 1543 230 1596 231
rect 1614 230 1720 231
rect 1543 229 1595 230
rect 1613 229 1719 230
rect 1514 228 1528 229
rect 1515 227 1528 228
rect 1542 228 1594 229
rect 1612 228 1661 229
rect 1662 228 1719 229
rect 1542 227 1593 228
rect 1611 227 1660 228
rect 1661 227 1718 228
rect 1516 225 1527 227
rect 1517 224 1527 225
rect 1541 226 1591 227
rect 1611 226 1658 227
rect 1661 226 1717 227
rect 1541 225 1590 226
rect 1610 225 1657 226
rect 1541 224 1589 225
rect 1609 224 1655 225
rect 1660 224 1716 226
rect 1518 223 1527 224
rect 1519 222 1527 223
rect 1520 221 1527 222
rect 1540 223 1588 224
rect 1608 223 1654 224
rect 1659 223 1715 224
rect 1540 222 1587 223
rect 1608 222 1653 223
rect 1659 222 1714 223
rect 1540 221 1586 222
rect 1607 221 1652 222
rect 1658 221 1713 222
rect 1521 220 1527 221
rect 1522 219 1527 220
rect 1523 218 1527 219
rect 1524 217 1527 218
rect 1539 220 1585 221
rect 1606 220 1650 221
rect 1658 220 1712 221
rect 1539 218 1584 220
rect 1605 219 1649 220
rect 1657 219 1711 220
rect 1605 218 1648 219
rect 1539 217 1583 218
rect 1604 217 1647 218
rect 1657 217 1710 219
rect 1525 216 1527 217
rect 1526 215 1527 216
rect 1538 216 1582 217
rect 1603 216 1646 217
rect 1656 216 1709 217
rect 1538 215 1581 216
rect 1603 215 1645 216
rect 1656 215 1708 216
rect 1538 213 1580 215
rect 1602 214 1644 215
rect 1656 214 1707 215
rect 1602 213 1643 214
rect 1656 213 1706 214
rect 1538 212 1579 213
rect 1601 212 1643 213
rect 1655 212 1705 213
rect 1537 210 1578 212
rect 1601 211 1642 212
rect 1655 211 1704 212
rect 1600 210 1641 211
rect 1655 210 1703 211
rect 1537 208 1577 210
rect 1600 209 1640 210
rect 1599 208 1640 209
rect 1655 209 1702 210
rect 1655 208 1701 209
rect 1537 206 1576 208
rect 1599 207 1639 208
rect 1654 207 1699 208
rect 1599 206 1638 207
rect 1537 203 1575 206
rect 1598 205 1638 206
rect 1654 206 1698 207
rect 1654 205 1697 206
rect 1598 204 1637 205
rect 1597 203 1637 204
rect 1654 204 1696 205
rect 1654 203 1695 204
rect 1537 202 1574 203
rect 1538 200 1574 202
rect 1597 202 1636 203
rect 1654 202 1694 203
rect 1597 201 1635 202
rect 1654 201 1692 202
rect 1538 199 1573 200
rect 1539 197 1573 199
rect 1596 199 1635 201
rect 1653 200 1691 201
rect 1653 199 1690 200
rect 1596 197 1634 199
rect 1653 198 1689 199
rect 1653 197 1687 198
rect 1540 196 1573 197
rect 1540 195 1572 196
rect 1541 193 1572 195
rect 1542 192 1572 193
rect 1595 194 1633 197
rect 1653 196 1686 197
rect 1653 195 1685 196
rect 1653 194 1683 195
rect 1595 192 1632 194
rect 1543 190 1572 192
rect 1544 189 1572 190
rect 1545 188 1572 189
rect 1546 186 1572 188
rect 1547 185 1572 186
rect 1548 184 1572 185
rect 1549 183 1572 184
rect 1550 182 1572 183
rect 1552 181 1572 182
rect 1553 180 1572 181
rect 1554 179 1572 180
rect 997 178 1065 179
rect 1166 178 1247 179
rect 1287 178 1355 179
rect 1556 178 1572 179
rect 1594 191 1632 192
rect 1653 193 1682 194
rect 1653 192 1680 193
rect 1653 191 1679 192
rect 1594 187 1631 191
rect 1653 190 1678 191
rect 1653 189 1676 190
rect 1653 188 1675 189
rect 1653 187 1674 188
rect 1594 181 1630 187
rect 1653 186 1673 187
rect 1653 185 1672 186
rect 1653 184 1671 185
rect 1654 183 1670 184
rect 1654 181 1669 183
rect 505 177 695 178
rect 817 177 882 178
rect 1167 177 1249 178
rect 1288 177 1354 178
rect 1557 177 1573 178
rect 1168 176 1249 177
rect 1558 176 1573 177
rect 1169 175 1251 176
rect 1560 175 1573 176
rect 1594 175 1629 181
rect 1654 180 1668 181
rect 1654 179 1667 180
rect 1654 177 1666 179
rect 1654 176 1665 177
rect 1170 174 1251 175
rect 1561 174 1573 175
rect 1171 173 1253 174
rect 1562 173 1573 174
rect 1172 172 1253 173
rect 1564 172 1573 173
rect 1173 171 1255 172
rect 1565 171 1574 172
rect 1174 170 1255 171
rect 1566 170 1574 171
rect 1595 170 1629 175
rect 1655 174 1664 176
rect 1655 173 1663 174
rect 1655 172 1662 173
rect 1175 169 1257 170
rect 1567 169 1574 170
rect 1176 168 1258 169
rect 1569 168 1574 169
rect 1177 167 1259 168
rect 1570 167 1575 168
rect 1596 167 1629 170
rect 1656 171 1662 172
rect 1656 169 1661 171
rect 1656 168 1660 169
rect 1178 166 1259 167
rect 1571 166 1575 167
rect 1573 165 1575 166
rect 1597 165 1629 167
rect 1657 167 1660 168
rect 1657 165 1659 167
rect 1574 164 1575 165
rect 1598 163 1629 165
rect 1599 162 1629 163
rect 1599 161 1630 162
rect 1600 159 1630 161
rect 1601 157 1630 159
rect 1602 156 1630 157
rect 1603 154 1631 156
rect 1604 153 1631 154
rect 1605 152 1631 153
rect 1606 151 1631 152
rect 1607 150 1632 151
rect 1608 149 1632 150
rect 1609 148 1632 149
rect 1610 147 1632 148
rect 1611 146 1633 147
rect 1612 145 1633 146
rect 1613 144 1633 145
rect 1614 143 1634 144
rect 1615 142 1634 143
rect 1617 141 1634 142
rect 1618 140 1635 141
rect 1619 139 1635 140
rect 1621 138 1635 139
rect 1622 137 1636 138
rect 1305 136 1318 137
rect 1624 136 1636 137
rect 491 135 515 136
rect 532 135 541 136
rect 738 135 747 136
rect 835 135 843 136
rect 490 133 516 135
rect 490 132 515 133
rect 490 129 516 132
rect 491 127 515 129
rect 481 123 526 124
rect 480 115 526 123
rect 481 114 525 115
rect 532 114 542 135
rect 588 132 642 133
rect 587 126 643 132
rect 687 130 724 131
rect 587 123 642 126
rect 631 117 642 123
rect 686 122 725 130
rect 687 121 724 122
rect 699 120 712 121
rect 699 119 711 120
rect 700 117 711 119
rect 737 118 747 135
rect 785 127 825 128
rect 785 121 826 127
rect 784 119 826 121
rect 785 118 826 119
rect 724 117 747 118
rect 799 117 811 118
rect 631 116 641 117
rect 532 113 543 114
rect 545 113 546 114
rect 547 113 549 114
rect 630 113 641 116
rect 699 115 711 117
rect 699 113 712 115
rect 497 111 510 112
rect 493 110 513 111
rect 491 109 516 110
rect 489 108 517 109
rect 487 107 519 108
rect 486 106 520 107
rect 485 105 521 106
rect 484 104 521 105
rect 484 103 522 104
rect 532 103 551 113
rect 630 110 640 113
rect 699 112 713 113
rect 698 110 713 112
rect 629 106 640 110
rect 697 109 714 110
rect 697 108 715 109
rect 723 108 747 117
rect 800 112 811 117
rect 696 107 716 108
rect 695 106 716 107
rect 628 105 640 106
rect 694 105 718 106
rect 580 104 650 105
rect 693 104 719 105
rect 483 102 500 103
rect 507 102 523 103
rect 483 101 496 102
rect 510 101 523 102
rect 482 100 495 101
rect 511 100 523 101
rect 482 95 494 100
rect 512 99 523 100
rect 532 102 543 103
rect 512 98 524 99
rect 512 97 523 98
rect 512 95 524 97
rect 483 94 495 95
rect 511 94 523 95
rect 483 93 497 94
rect 509 93 523 94
rect 484 92 500 93
rect 506 92 522 93
rect 484 91 522 92
rect 485 90 521 91
rect 486 89 520 90
rect 487 88 519 89
rect 488 87 518 88
rect 490 86 517 87
rect 492 85 514 86
rect 494 84 512 85
rect 491 79 501 80
rect 490 68 502 79
rect 532 78 542 102
rect 579 96 651 104
rect 692 103 720 104
rect 691 102 721 103
rect 690 101 705 102
rect 707 101 723 102
rect 689 100 704 101
rect 707 100 724 101
rect 687 99 704 100
rect 708 99 727 100
rect 686 98 703 99
rect 709 98 727 99
rect 684 97 702 98
rect 710 97 727 98
rect 682 96 701 97
rect 711 96 727 97
rect 580 95 650 96
rect 681 95 700 96
rect 713 95 726 96
rect 607 94 619 95
rect 682 94 699 95
rect 714 94 725 95
rect 608 84 618 94
rect 683 93 698 94
rect 715 93 725 94
rect 684 92 697 93
rect 716 92 724 93
rect 684 91 695 92
rect 719 91 723 92
rect 685 90 694 91
rect 720 90 723 91
rect 686 89 692 90
rect 687 88 691 89
rect 608 83 619 84
rect 588 82 641 83
rect 532 77 541 78
rect 587 73 642 82
rect 588 72 642 73
rect 490 67 542 68
rect 490 59 544 67
rect 491 58 544 59
rect 632 57 642 72
rect 695 69 705 84
rect 737 78 747 108
rect 799 107 811 112
rect 799 104 812 107
rect 798 103 812 104
rect 834 106 844 135
rect 890 126 944 134
rect 1002 133 1011 134
rect 1002 126 1012 133
rect 890 125 902 126
rect 904 125 905 126
rect 939 125 941 126
rect 890 124 901 125
rect 890 123 900 124
rect 890 122 901 123
rect 890 121 943 122
rect 890 115 944 121
rect 1001 120 1012 126
rect 1001 119 1013 120
rect 1000 116 1013 119
rect 890 114 943 115
rect 890 113 902 114
rect 1000 113 1014 116
rect 890 112 901 113
rect 999 112 1015 113
rect 890 111 900 112
rect 998 111 1015 112
rect 890 110 901 111
rect 998 110 1016 111
rect 890 109 902 110
rect 904 109 905 110
rect 942 109 943 110
rect 997 109 1016 110
rect 834 105 846 106
rect 848 105 849 106
rect 850 105 852 106
rect 798 101 813 103
rect 797 98 813 101
rect 797 97 814 98
rect 796 96 815 97
rect 795 94 815 96
rect 834 95 854 105
rect 890 101 945 109
rect 996 108 1017 109
rect 996 107 1018 108
rect 995 106 1019 107
rect 994 105 1020 106
rect 994 104 1021 105
rect 992 102 1006 104
rect 1008 103 1022 104
rect 1008 102 1023 103
rect 990 101 1005 102
rect 1009 101 1025 102
rect 891 100 944 101
rect 989 100 1004 101
rect 1010 100 1026 101
rect 911 97 923 100
rect 988 99 1003 100
rect 1011 99 1028 100
rect 987 98 1002 99
rect 1012 98 1030 99
rect 985 97 1002 98
rect 1013 97 1030 98
rect 910 96 923 97
rect 984 96 1001 97
rect 1014 96 1030 97
rect 883 95 908 96
rect 909 95 924 96
rect 925 95 948 96
rect 949 95 951 96
rect 982 95 1000 96
rect 1015 95 1030 96
rect 834 94 853 95
rect 881 94 952 95
rect 982 94 999 95
rect 1016 94 1029 95
rect 795 93 816 94
rect 794 92 817 93
rect 793 91 817 92
rect 793 90 818 91
rect 792 89 805 90
rect 807 89 819 90
rect 791 87 804 89
rect 807 88 820 89
rect 807 87 821 88
rect 790 86 803 87
rect 808 86 822 87
rect 789 85 803 86
rect 809 85 823 86
rect 788 84 802 85
rect 809 84 824 85
rect 787 83 801 84
rect 810 83 825 84
rect 786 82 801 83
rect 811 82 826 83
rect 785 81 800 82
rect 811 81 827 82
rect 784 80 799 81
rect 812 80 828 81
rect 782 79 798 80
rect 813 79 829 80
rect 781 78 797 79
rect 814 78 828 79
rect 780 77 797 78
rect 815 77 827 78
rect 780 76 796 77
rect 816 76 826 77
rect 781 75 795 76
rect 817 75 826 76
rect 781 74 794 75
rect 818 74 825 75
rect 783 73 793 74
rect 820 73 824 74
rect 783 72 792 73
rect 821 72 823 73
rect 785 71 790 72
rect 786 70 789 71
rect 695 68 706 69
rect 695 58 749 68
rect 834 57 844 94
rect 881 87 953 94
rect 982 93 998 94
rect 1018 93 1028 94
rect 983 92 997 93
rect 1019 92 1028 93
rect 984 91 995 92
rect 1021 91 1027 92
rect 985 90 994 91
rect 1022 90 1026 91
rect 986 89 993 90
rect 987 88 992 89
rect 988 87 990 88
rect 881 86 952 87
rect 916 83 917 84
rect 997 83 1002 84
rect 1003 83 1005 84
rect 906 82 927 83
rect 900 81 933 82
rect 898 80 936 81
rect 895 79 938 80
rect 894 78 940 79
rect 892 77 941 78
rect 891 76 942 77
rect 890 75 944 76
rect 889 74 944 75
rect 889 73 907 74
rect 926 73 945 74
rect 888 72 904 73
rect 930 72 945 73
rect 888 67 901 72
rect 932 71 946 72
rect 933 70 946 71
rect 934 69 946 70
rect 933 67 946 69
rect 888 66 902 67
rect 932 66 946 67
rect 996 69 1006 83
rect 1038 78 1048 136
rect 1139 135 1148 136
rect 1301 135 1322 136
rect 1107 133 1108 134
rect 1100 132 1111 133
rect 1097 131 1115 132
rect 1095 130 1116 131
rect 1094 129 1118 130
rect 1093 128 1119 129
rect 1092 127 1120 128
rect 1091 126 1121 127
rect 1138 126 1149 135
rect 1300 134 1323 135
rect 1298 133 1325 134
rect 1297 132 1326 133
rect 1090 125 1149 126
rect 1089 124 1149 125
rect 1088 123 1104 124
rect 1107 123 1149 124
rect 1088 122 1102 123
rect 1110 122 1149 123
rect 1191 122 1247 132
rect 1296 131 1327 132
rect 1295 130 1328 131
rect 1294 129 1329 130
rect 1293 128 1329 129
rect 1293 127 1306 128
rect 1317 127 1330 128
rect 1293 126 1305 127
rect 1318 126 1330 127
rect 1293 125 1304 126
rect 1319 125 1331 126
rect 1088 121 1100 122
rect 1112 121 1149 122
rect 1235 121 1247 122
rect 1087 120 1099 121
rect 1113 120 1149 121
rect 1236 120 1246 121
rect 1087 119 1098 120
rect 1086 118 1098 119
rect 1114 118 1149 120
rect 1086 116 1097 118
rect 1115 116 1149 118
rect 1086 109 1096 116
rect 1115 115 1126 116
rect 1138 115 1149 116
rect 1116 110 1126 115
rect 1139 114 1149 115
rect 1138 110 1149 114
rect 1235 115 1246 120
rect 1292 119 1303 125
rect 1320 123 1331 125
rect 1321 121 1331 123
rect 1320 119 1331 121
rect 1293 118 1304 119
rect 1319 118 1331 119
rect 1293 117 1306 118
rect 1317 117 1330 118
rect 1293 116 1307 117
rect 1316 116 1330 117
rect 1293 115 1329 116
rect 1235 111 1245 115
rect 1294 114 1329 115
rect 1295 113 1328 114
rect 1295 112 1327 113
rect 1297 111 1326 112
rect 1086 108 1097 109
rect 1115 108 1149 110
rect 1086 106 1098 108
rect 1114 106 1149 108
rect 1234 107 1245 111
rect 1298 110 1325 111
rect 1300 109 1323 110
rect 1301 108 1322 109
rect 1306 107 1318 108
rect 1234 106 1244 107
rect 1087 105 1098 106
rect 1113 105 1149 106
rect 1087 104 1100 105
rect 1112 104 1149 105
rect 1088 103 1101 104
rect 1111 103 1149 104
rect 1088 102 1103 103
rect 1109 102 1149 103
rect 1088 101 1149 102
rect 1089 100 1149 101
rect 1233 104 1244 106
rect 1334 105 1338 106
rect 1327 104 1339 105
rect 1233 100 1243 104
rect 1287 102 1339 104
rect 1090 99 1122 100
rect 1138 99 1149 100
rect 1232 99 1243 100
rect 1091 98 1121 99
rect 1139 98 1149 99
rect 1184 98 1254 99
rect 1092 97 1120 98
rect 1093 96 1119 97
rect 1094 95 1117 96
rect 1096 94 1116 95
rect 1098 93 1113 94
rect 1100 92 1111 93
rect 1096 69 1106 84
rect 1138 79 1149 98
rect 1183 90 1255 98
rect 1286 96 1339 102
rect 1286 95 1335 96
rect 1287 94 1328 95
rect 1302 93 1314 94
rect 1341 93 1351 136
rect 1626 135 1636 136
rect 1627 134 1637 135
rect 1629 133 1637 134
rect 1631 132 1638 133
rect 1633 131 1638 132
rect 1636 130 1639 131
rect 1642 98 1655 99
rect 1416 95 1437 98
rect 1443 95 1461 98
rect 1466 96 1486 98
rect 1467 95 1486 96
rect 1494 95 1510 98
rect 1516 96 1537 98
rect 1546 96 1564 98
rect 1568 97 1582 98
rect 1600 97 1617 98
rect 1638 97 1660 98
rect 1568 96 1583 97
rect 1600 96 1618 97
rect 1635 96 1662 97
rect 1516 95 1536 96
rect 1547 95 1564 96
rect 1569 95 1583 96
rect 1601 95 1617 96
rect 1633 95 1644 96
rect 1651 95 1662 96
rect 1688 95 1709 98
rect 1716 96 1737 98
rect 1717 95 1737 96
rect 1746 96 1778 98
rect 1746 95 1779 96
rect 1789 95 1822 98
rect 1420 94 1433 95
rect 1447 94 1457 95
rect 1470 94 1483 95
rect 1498 94 1507 95
rect 1520 94 1533 95
rect 1550 94 1561 95
rect 1572 94 1584 95
rect 1605 94 1614 95
rect 1632 94 1641 95
rect 1654 94 1662 95
rect 1692 94 1705 95
rect 1721 94 1733 95
rect 1750 94 1761 95
rect 1770 94 1779 95
rect 1793 94 1805 95
rect 1813 94 1822 95
rect 1421 93 1432 94
rect 1447 93 1454 94
rect 1471 93 1482 94
rect 1498 93 1505 94
rect 1521 93 1532 94
rect 1551 93 1560 94
rect 1574 93 1585 94
rect 1606 93 1613 94
rect 1630 93 1640 94
rect 1655 93 1663 94
rect 1693 93 1704 94
rect 1721 93 1732 94
rect 1303 92 1314 93
rect 1184 89 1254 90
rect 1211 88 1223 89
rect 1139 78 1148 79
rect 996 68 1007 69
rect 1096 68 1107 69
rect 996 67 1049 68
rect 889 65 905 66
rect 929 65 945 66
rect 889 64 909 65
rect 926 64 945 65
rect 890 63 944 64
rect 891 62 944 63
rect 892 61 943 62
rect 893 60 942 61
rect 895 59 940 60
rect 896 58 938 59
rect 996 58 1050 67
rect 1096 58 1150 68
rect 899 57 935 58
rect 1212 57 1223 88
rect 1303 81 1313 92
rect 1326 91 1328 92
rect 1331 91 1338 92
rect 1340 91 1351 93
rect 1325 90 1351 91
rect 1324 83 1351 90
rect 1325 82 1351 83
rect 1340 81 1351 82
rect 1304 80 1306 81
rect 1307 80 1312 81
rect 1298 77 1308 78
rect 1298 68 1309 77
rect 1341 76 1351 81
rect 1422 77 1431 93
rect 1446 92 1453 93
rect 1472 92 1483 93
rect 1446 91 1451 92
rect 1473 91 1483 92
rect 1498 92 1504 93
rect 1498 91 1503 92
rect 1445 90 1450 91
rect 1473 90 1484 91
rect 1498 90 1502 91
rect 1444 89 1449 90
rect 1474 89 1484 90
rect 1497 89 1502 90
rect 1443 88 1448 89
rect 1474 88 1485 89
rect 1497 88 1501 89
rect 1443 87 1447 88
rect 1475 87 1485 88
rect 1496 87 1501 88
rect 1442 86 1446 87
rect 1441 85 1445 86
rect 1476 85 1486 87
rect 1496 86 1500 87
rect 1440 84 1444 85
rect 1439 83 1443 84
rect 1477 83 1487 85
rect 1495 84 1499 86
rect 1438 82 1442 83
rect 1437 81 1441 82
rect 1478 81 1488 83
rect 1494 82 1498 84
rect 1493 81 1497 82
rect 1436 80 1440 81
rect 1479 80 1489 81
rect 1493 80 1496 81
rect 1435 79 1441 80
rect 1434 78 1441 79
rect 1480 79 1489 80
rect 1492 79 1496 80
rect 1480 78 1490 79
rect 1492 78 1495 79
rect 1432 77 1442 78
rect 1481 77 1490 78
rect 1491 77 1495 78
rect 1422 76 1443 77
rect 1481 76 1494 77
rect 1422 74 1444 76
rect 1482 75 1494 76
rect 1482 74 1493 75
rect 1298 67 1352 68
rect 1298 59 1353 67
rect 1298 58 1352 59
rect 1422 58 1431 74
rect 1433 73 1445 74
rect 1434 72 1446 73
rect 1435 71 1446 72
rect 1436 70 1447 71
rect 1436 69 1448 70
rect 1437 68 1449 69
rect 1438 67 1449 68
rect 1438 66 1450 67
rect 1439 65 1451 66
rect 1440 63 1452 65
rect 1441 62 1453 63
rect 1442 61 1454 62
rect 1443 60 1455 61
rect 1443 59 1456 60
rect 1444 58 1456 59
rect 1421 57 1432 58
rect 1445 57 1458 58
rect 1483 57 1493 74
rect 1521 69 1531 93
rect 1552 88 1559 93
rect 1574 92 1586 93
rect 1575 91 1587 92
rect 1575 90 1588 91
rect 1575 88 1589 90
rect 1552 87 1558 88
rect 1553 69 1558 87
rect 1522 67 1531 69
rect 1522 63 1532 67
rect 1552 65 1558 69
rect 1575 87 1590 88
rect 1607 87 1612 93
rect 1629 92 1638 93
rect 1656 92 1663 93
rect 1628 91 1637 92
rect 1657 91 1663 92
rect 1627 90 1636 91
rect 1658 90 1663 91
rect 1626 89 1636 90
rect 1625 88 1635 89
rect 1659 88 1663 90
rect 1575 86 1591 87
rect 1552 64 1557 65
rect 1523 61 1533 63
rect 1551 61 1557 64
rect 1523 60 1534 61
rect 1550 60 1556 61
rect 1524 59 1535 60
rect 1549 59 1556 60
rect 1575 60 1579 86
rect 1580 85 1592 86
rect 1581 84 1593 85
rect 1581 83 1594 84
rect 1582 82 1595 83
rect 1583 81 1596 82
rect 1584 80 1596 81
rect 1585 79 1597 80
rect 1586 78 1598 79
rect 1587 77 1599 78
rect 1587 76 1600 77
rect 1588 75 1601 76
rect 1589 74 1602 75
rect 1590 73 1603 74
rect 1591 72 1603 73
rect 1592 71 1604 72
rect 1592 70 1605 71
rect 1593 69 1606 70
rect 1594 68 1607 69
rect 1608 68 1611 87
rect 1624 86 1634 88
rect 1623 83 1633 86
rect 1660 85 1663 88
rect 1694 91 1704 93
rect 1622 82 1633 83
rect 1622 80 1632 82
rect 1621 70 1632 80
rect 1694 79 1703 91
rect 1722 79 1732 93
rect 1694 75 1732 79
rect 1646 74 1666 75
rect 1694 74 1704 75
rect 1646 72 1667 74
rect 1649 71 1665 72
rect 1652 70 1664 71
rect 1595 67 1611 68
rect 1596 66 1611 67
rect 1622 66 1633 70
rect 1653 68 1663 70
rect 1597 64 1611 66
rect 1623 64 1634 66
rect 1598 63 1611 64
rect 1599 62 1611 63
rect 1624 62 1635 64
rect 1600 61 1611 62
rect 1625 61 1636 62
rect 1601 60 1611 61
rect 1626 60 1637 61
rect 1575 59 1580 60
rect 1524 58 1536 59
rect 1548 58 1555 59
rect 1525 57 1538 58
rect 1546 57 1555 58
rect 1574 57 1580 59
rect 1602 58 1611 60
rect 1627 59 1637 60
rect 1654 59 1663 68
rect 1628 58 1638 59
rect 1603 57 1611 58
rect 1629 57 1640 58
rect 632 56 641 57
rect 835 56 843 57
rect 901 56 933 57
rect 1213 56 1222 57
rect 1421 56 1433 57
rect 1445 56 1459 57
rect 1482 56 1494 57
rect 1526 56 1554 57
rect 1573 56 1581 57
rect 1604 56 1611 57
rect 1630 56 1641 57
rect 1653 56 1663 59
rect 1694 59 1703 74
rect 1694 58 1704 59
rect 1693 57 1704 58
rect 1722 57 1732 75
rect 1751 78 1761 94
rect 1773 93 1779 94
rect 1774 92 1779 93
rect 1775 90 1779 92
rect 1776 87 1779 90
rect 1773 82 1775 83
rect 1772 79 1775 82
rect 1771 78 1775 79
rect 1751 74 1775 78
rect 1751 57 1761 74
rect 1771 73 1775 74
rect 1772 70 1775 73
rect 1773 69 1775 70
rect 1794 78 1804 94
rect 1816 93 1822 94
rect 1817 92 1822 93
rect 1818 90 1822 92
rect 1819 87 1822 90
rect 1816 81 1819 83
rect 1815 79 1819 81
rect 1814 78 1819 79
rect 1794 74 1819 78
rect 1780 64 1782 65
rect 1779 62 1782 64
rect 1778 60 1782 62
rect 1777 59 1782 60
rect 1776 58 1781 59
rect 1775 57 1781 58
rect 1794 58 1804 74
rect 1814 73 1819 74
rect 1815 71 1819 73
rect 1816 69 1819 71
rect 1823 64 1826 65
rect 1822 63 1826 64
rect 1822 62 1825 63
rect 1821 60 1825 62
rect 1820 59 1825 60
rect 1819 58 1825 59
rect 1794 57 1805 58
rect 1818 57 1824 58
rect 1693 56 1705 57
rect 1721 56 1733 57
rect 1750 56 1763 57
rect 1773 56 1781 57
rect 1793 56 1806 57
rect 1816 56 1824 57
rect 908 55 927 56
rect 1417 55 1437 56
rect 1446 55 1462 56
rect 1478 55 1498 56
rect 1527 55 1553 56
rect 1570 55 1585 56
rect 1605 55 1611 56
rect 1632 55 1644 56
rect 1652 55 1663 56
rect 1689 55 1708 56
rect 1717 55 1737 56
rect 1416 53 1437 55
rect 1447 53 1462 55
rect 1477 53 1500 55
rect 1528 54 1552 55
rect 1530 53 1550 54
rect 1569 53 1586 55
rect 1606 54 1611 55
rect 1634 54 1663 55
rect 1533 52 1547 53
rect 1607 52 1611 54
rect 1636 53 1660 54
rect 1688 53 1709 55
rect 1716 53 1737 55
rect 1745 54 1781 56
rect 1789 55 1824 56
rect 1788 54 1824 55
rect 1745 53 1780 54
rect 1788 53 1823 54
rect 1640 52 1655 53
rect 503 41 506 42
rect 716 41 719 42
rect 770 41 772 42
rect 1192 41 1195 42
rect 483 38 497 39
rect 482 35 498 38
rect 482 34 497 35
rect 482 33 489 34
rect 482 28 488 33
rect 482 27 489 28
rect 482 25 496 27
rect 482 23 497 25
rect 482 21 496 23
rect 482 20 489 21
rect 482 14 488 20
rect 482 13 496 14
rect 482 12 497 13
rect 482 9 498 12
rect 501 9 506 41
rect 615 40 617 41
rect 549 36 552 37
rect 547 35 552 36
rect 613 35 618 40
rect 516 31 521 32
rect 535 31 540 32
rect 546 31 552 35
rect 614 34 618 35
rect 567 31 569 32
rect 577 31 582 32
rect 600 31 605 32
rect 628 31 633 32
rect 642 31 647 32
rect 667 31 673 32
rect 691 31 694 32
rect 708 31 711 32
rect 714 31 720 41
rect 732 38 750 39
rect 731 37 750 38
rect 731 35 751 37
rect 731 34 750 35
rect 737 33 745 34
rect 514 30 523 31
rect 533 30 542 31
rect 544 30 555 31
rect 559 30 562 31
rect 565 30 570 31
rect 575 30 584 31
rect 593 30 596 31
rect 598 30 606 31
rect 614 30 618 31
rect 626 30 635 31
rect 640 30 649 31
rect 664 30 675 31
rect 682 30 696 31
rect 705 30 720 31
rect 512 29 524 30
rect 532 29 556 30
rect 512 28 525 29
rect 531 28 556 29
rect 511 27 525 28
rect 530 27 556 28
rect 510 26 526 27
rect 530 26 542 27
rect 544 26 555 27
rect 558 26 570 30
rect 574 29 586 30
rect 573 28 586 29
rect 572 27 587 28
rect 592 27 608 30
rect 572 26 588 27
rect 510 25 516 26
rect 520 25 526 26
rect 510 23 515 25
rect 510 22 516 23
rect 521 22 526 25
rect 529 24 536 26
rect 529 23 535 24
rect 510 19 527 22
rect 510 17 526 19
rect 528 17 534 23
rect 510 15 515 17
rect 528 16 535 17
rect 529 15 535 16
rect 510 14 516 15
rect 529 14 536 15
rect 546 14 552 26
rect 558 25 578 26
rect 582 25 588 26
rect 592 26 609 27
rect 558 24 566 25
rect 570 24 577 25
rect 582 24 589 25
rect 558 23 565 24
rect 510 13 517 14
rect 522 13 525 14
rect 530 13 537 14
rect 540 13 542 14
rect 511 11 526 13
rect 530 12 542 13
rect 546 13 553 14
rect 546 12 556 13
rect 530 11 543 12
rect 547 11 556 12
rect 512 10 525 11
rect 531 10 543 11
rect 513 9 525 10
rect 532 9 543 10
rect 548 9 556 11
rect 558 9 564 23
rect 570 15 576 24
rect 583 22 589 24
rect 584 18 589 22
rect 583 15 589 18
rect 570 14 577 15
rect 582 14 589 15
rect 592 24 599 26
rect 603 24 609 26
rect 571 13 578 14
rect 581 13 588 14
rect 572 12 588 13
rect 572 11 587 12
rect 573 10 586 11
rect 574 9 585 10
rect 592 9 598 24
rect 604 9 609 24
rect 613 9 618 30
rect 625 29 635 30
rect 624 28 635 29
rect 638 28 650 30
rect 664 29 676 30
rect 682 29 697 30
rect 704 29 720 30
rect 623 27 635 28
rect 637 27 650 28
rect 663 28 677 29
rect 623 26 634 27
rect 637 26 649 27
rect 663 26 678 28
rect 622 24 629 26
rect 637 25 643 26
rect 663 25 666 26
rect 672 25 678 26
rect 636 24 643 25
rect 664 24 665 25
rect 622 21 628 24
rect 637 23 643 24
rect 673 23 678 25
rect 637 22 645 23
rect 667 22 678 23
rect 637 21 647 22
rect 665 21 678 22
rect 622 18 627 21
rect 638 20 648 21
rect 664 20 678 21
rect 638 19 649 20
rect 663 19 678 20
rect 639 18 650 19
rect 622 15 628 18
rect 642 17 650 18
rect 643 16 650 17
rect 662 18 678 19
rect 662 17 668 18
rect 662 16 667 17
rect 673 16 678 18
rect 622 14 629 15
rect 622 13 630 14
rect 633 13 635 14
rect 638 13 640 14
rect 644 13 650 16
rect 661 14 667 16
rect 672 14 678 16
rect 623 11 636 13
rect 624 10 636 11
rect 625 9 636 10
rect 637 11 650 13
rect 662 13 668 14
rect 671 13 678 14
rect 662 11 678 13
rect 637 10 649 11
rect 663 10 678 11
rect 637 9 648 10
rect 664 9 678 10
rect 682 27 698 29
rect 682 26 699 27
rect 703 26 720 29
rect 682 25 689 26
rect 692 25 699 26
rect 682 22 688 25
rect 483 8 497 9
rect 502 8 506 9
rect 515 8 524 9
rect 533 8 542 9
rect 549 8 556 9
rect 559 8 563 9
rect 575 8 584 9
rect 593 8 597 9
rect 604 8 608 9
rect 614 8 618 9
rect 626 8 635 9
rect 638 8 647 9
rect 664 8 671 9
rect 674 8 677 9
rect 682 8 687 22
rect 693 9 699 25
rect 702 25 709 26
rect 712 25 720 26
rect 702 21 708 25
rect 713 23 720 25
rect 702 18 707 21
rect 702 15 708 18
rect 714 16 720 23
rect 702 14 709 15
rect 713 14 720 16
rect 702 13 710 14
rect 712 13 720 14
rect 703 11 720 13
rect 704 10 720 11
rect 705 9 720 10
rect 738 9 744 33
rect 754 31 759 32
rect 752 30 761 31
rect 751 29 762 30
rect 750 28 763 29
rect 749 27 763 28
rect 749 26 764 27
rect 748 25 754 26
rect 748 23 753 25
rect 759 24 764 26
rect 747 22 754 23
rect 759 22 765 24
rect 747 18 765 22
rect 747 17 764 18
rect 747 16 754 17
rect 748 15 753 16
rect 748 14 754 15
rect 748 13 755 14
rect 760 13 764 14
rect 749 11 764 13
rect 750 10 764 11
rect 751 9 763 10
rect 768 9 773 41
rect 937 40 940 41
rect 995 40 997 41
rect 1191 40 1196 41
rect 1282 40 1284 41
rect 936 35 941 40
rect 983 36 986 37
rect 982 35 986 36
rect 993 35 998 40
rect 1070 38 1082 39
rect 937 34 940 35
rect 981 32 986 35
rect 994 34 998 35
rect 1069 37 1084 38
rect 1069 36 1085 37
rect 1069 34 1086 36
rect 1069 33 1076 34
rect 1078 33 1086 34
rect 783 31 787 32
rect 802 31 807 32
rect 818 31 822 32
rect 841 31 844 32
rect 851 31 855 32
rect 871 31 875 32
rect 882 31 886 32
rect 923 31 928 32
rect 951 31 956 32
rect 965 31 971 32
rect 980 31 987 32
rect 1009 31 1014 32
rect 1033 31 1036 32
rect 1049 31 1054 32
rect 780 30 789 31
rect 800 30 809 31
rect 815 30 825 31
rect 833 30 837 31
rect 839 30 846 31
rect 850 30 857 31
rect 864 30 877 31
rect 880 30 888 31
rect 895 30 899 31
rect 906 30 910 31
rect 915 30 919 31
rect 921 30 929 31
rect 936 30 940 31
rect 949 30 958 31
rect 963 30 973 31
rect 978 30 990 31
rect 994 30 998 31
rect 1007 30 1016 31
rect 1024 30 1028 31
rect 1030 30 1038 31
rect 1047 30 1056 31
rect 779 28 791 30
rect 799 29 809 30
rect 814 29 826 30
rect 833 29 847 30
rect 848 29 858 30
rect 798 28 809 29
rect 778 27 792 28
rect 777 26 792 27
rect 797 27 809 28
rect 813 28 827 29
rect 813 27 828 28
rect 797 26 808 27
rect 812 26 829 27
rect 777 25 783 26
rect 787 25 793 26
rect 777 23 782 25
rect 776 22 782 23
rect 788 22 793 25
rect 796 25 803 26
rect 811 25 818 26
rect 822 25 829 26
rect 796 24 802 25
rect 776 17 793 22
rect 776 15 782 17
rect 795 16 801 24
rect 811 22 817 25
rect 823 23 829 25
rect 833 26 859 29
rect 833 23 839 26
rect 843 25 850 26
rect 853 25 859 26
rect 811 20 816 22
rect 810 19 816 20
rect 811 18 816 19
rect 795 15 802 16
rect 811 15 817 18
rect 824 17 830 23
rect 777 14 783 15
rect 796 14 803 15
rect 811 14 818 15
rect 823 14 829 17
rect 777 13 784 14
rect 788 13 792 14
rect 796 13 804 14
rect 807 13 809 14
rect 811 13 819 14
rect 822 13 829 14
rect 777 12 793 13
rect 778 11 792 12
rect 797 11 809 13
rect 812 12 828 13
rect 779 10 792 11
rect 798 10 809 11
rect 813 11 828 12
rect 813 10 827 11
rect 780 9 792 10
rect 799 9 809 10
rect 815 9 826 10
rect 833 9 838 23
rect 843 9 849 25
rect 854 11 859 25
rect 863 27 889 30
rect 863 26 890 27
rect 863 25 870 26
rect 873 25 881 26
rect 854 10 860 11
rect 854 9 859 10
rect 863 9 869 25
rect 873 23 880 25
rect 884 24 890 26
rect 874 9 879 23
rect 885 11 890 24
rect 894 15 899 30
rect 905 15 911 30
rect 894 14 900 15
rect 904 14 911 15
rect 894 13 901 14
rect 903 13 911 14
rect 894 11 911 13
rect 884 10 890 11
rect 895 10 911 11
rect 885 9 890 10
rect 896 9 911 10
rect 915 29 930 30
rect 915 26 931 29
rect 915 25 922 26
rect 925 25 932 26
rect 915 22 921 25
rect 915 11 920 22
rect 915 10 921 11
rect 694 8 698 9
rect 706 8 713 9
rect 715 8 719 9
rect 739 8 743 9
rect 752 8 762 9
rect 769 8 773 9
rect 781 8 791 9
rect 800 8 809 9
rect 816 8 825 9
rect 833 8 837 9
rect 844 8 848 9
rect 855 8 859 9
rect 864 8 868 9
rect 875 8 878 9
rect 885 8 889 9
rect 897 8 904 9
rect 907 8 910 9
rect 915 8 920 10
rect 926 9 932 25
rect 936 9 941 30
rect 948 29 958 30
rect 947 28 958 29
rect 946 27 958 28
rect 961 29 974 30
rect 961 27 975 29
rect 978 27 991 30
rect 945 26 957 27
rect 961 26 976 27
rect 979 26 990 27
rect 945 25 952 26
rect 962 25 964 26
rect 970 25 976 26
rect 945 24 951 25
rect 944 23 951 24
rect 971 23 976 25
rect 944 16 950 23
rect 965 22 976 23
rect 963 21 976 22
rect 961 20 976 21
rect 960 18 976 20
rect 960 17 966 18
rect 944 15 951 16
rect 945 14 951 15
rect 959 14 965 17
rect 971 16 976 18
rect 970 14 976 16
rect 945 13 953 14
rect 956 13 958 14
rect 946 11 958 13
rect 960 13 966 14
rect 969 13 976 14
rect 960 11 976 13
rect 981 16 986 26
rect 981 14 987 16
rect 981 13 988 14
rect 981 12 990 13
rect 947 10 958 11
rect 948 9 958 10
rect 961 9 976 11
rect 982 10 991 12
rect 983 9 991 10
rect 993 9 998 30
rect 1005 29 1017 30
rect 1024 29 1039 30
rect 1045 29 1056 30
rect 1004 28 1018 29
rect 1023 28 1040 29
rect 1004 27 1019 28
rect 1003 26 1019 27
rect 1024 26 1040 28
rect 1044 26 1056 29
rect 1069 27 1075 33
rect 1079 32 1086 33
rect 1080 31 1086 32
rect 1096 31 1100 32
rect 1113 31 1119 32
rect 1130 31 1135 32
rect 1149 31 1154 32
rect 1171 31 1173 32
rect 1181 31 1187 32
rect 1191 31 1197 40
rect 1222 38 1227 39
rect 1200 31 1203 32
rect 1081 29 1086 31
rect 1094 30 1103 31
rect 1111 30 1121 31
rect 1128 30 1137 31
rect 1146 30 1156 31
rect 1164 30 1167 31
rect 1170 30 1174 31
rect 1179 30 1188 31
rect 1191 30 1205 31
rect 1080 27 1086 29
rect 1092 28 1104 30
rect 1110 29 1121 30
rect 1127 29 1138 30
rect 1091 27 1105 28
rect 1109 27 1121 29
rect 1126 28 1139 29
rect 1125 27 1140 28
rect 1069 26 1076 27
rect 1078 26 1086 27
rect 1090 26 1106 27
rect 1002 25 1009 26
rect 1013 25 1020 26
rect 1002 22 1008 25
rect 1014 23 1020 25
rect 1023 25 1031 26
rect 1034 25 1040 26
rect 1023 23 1030 25
rect 1015 22 1020 23
rect 1024 22 1030 23
rect 1002 17 1007 22
rect 1015 17 1021 22
rect 1002 15 1008 17
rect 1015 16 1020 17
rect 1024 16 1029 22
rect 1035 21 1041 25
rect 1043 23 1050 26
rect 1069 25 1085 26
rect 1090 25 1096 26
rect 1100 25 1106 26
rect 1109 26 1116 27
rect 1117 26 1120 27
rect 1125 26 1132 27
rect 1133 26 1140 27
rect 1109 25 1114 26
rect 1036 20 1041 21
rect 1044 22 1052 23
rect 1044 21 1054 22
rect 1044 20 1055 21
rect 1069 20 1084 25
rect 1090 22 1095 25
rect 1101 22 1106 25
rect 1108 24 1114 25
rect 1124 24 1130 26
rect 1135 25 1140 26
rect 1145 27 1158 30
rect 1145 26 1159 27
rect 1145 25 1147 26
rect 1153 25 1159 26
rect 1135 24 1141 25
rect 1108 23 1115 24
rect 1124 23 1129 24
rect 1136 23 1141 24
rect 1154 23 1159 25
rect 1108 22 1117 23
rect 1124 22 1130 23
rect 1135 22 1141 23
rect 1148 22 1159 23
rect 1089 21 1106 22
rect 1109 21 1119 22
rect 1002 14 1009 15
rect 1014 14 1020 16
rect 1002 13 1010 14
rect 1012 13 1020 14
rect 1023 13 1029 16
rect 1035 13 1041 20
rect 1045 19 1056 20
rect 1046 18 1057 19
rect 1049 17 1057 18
rect 1050 16 1057 17
rect 1051 14 1057 16
rect 1003 12 1019 13
rect 1004 11 1018 12
rect 1024 11 1029 13
rect 1036 12 1041 13
rect 1005 10 1018 11
rect 1023 10 1030 11
rect 1006 9 1017 10
rect 1024 9 1029 10
rect 1035 9 1041 12
rect 1044 13 1046 14
rect 1050 13 1057 14
rect 1044 12 1057 13
rect 1044 10 1056 12
rect 1044 9 1055 10
rect 1069 9 1075 20
rect 1078 19 1085 20
rect 1079 18 1085 19
rect 1089 18 1107 21
rect 1109 20 1120 21
rect 1110 19 1121 20
rect 1111 18 1121 19
rect 1079 16 1086 18
rect 1089 17 1106 18
rect 1114 17 1122 18
rect 1089 16 1095 17
rect 1115 16 1122 17
rect 1080 14 1086 16
rect 1090 15 1095 16
rect 1090 14 1096 15
rect 1116 14 1122 16
rect 1124 17 1141 22
rect 1146 21 1159 22
rect 1145 20 1159 21
rect 1144 18 1159 20
rect 1143 17 1149 18
rect 1124 14 1130 17
rect 1138 14 1139 15
rect 1143 14 1148 17
rect 1154 15 1159 18
rect 1153 14 1159 15
rect 1080 13 1087 14
rect 1090 13 1097 14
rect 1102 13 1106 14
rect 1081 11 1087 13
rect 1091 11 1106 13
rect 1109 13 1111 14
rect 1115 13 1122 14
rect 1109 12 1122 13
rect 1125 13 1131 14
rect 1136 13 1140 14
rect 1109 11 1121 12
rect 1125 11 1140 13
rect 1143 13 1149 14
rect 1152 13 1159 14
rect 1143 11 1159 13
rect 1163 26 1174 30
rect 1178 29 1189 30
rect 1191 29 1206 30
rect 1177 28 1188 29
rect 1176 26 1188 28
rect 1191 27 1207 29
rect 1191 26 1208 27
rect 1163 25 1173 26
rect 1175 25 1183 26
rect 1163 23 1170 25
rect 1175 24 1182 25
rect 1191 24 1198 26
rect 1202 24 1208 26
rect 1081 10 1088 11
rect 1092 10 1105 11
rect 1108 10 1120 11
rect 1126 10 1140 11
rect 1144 10 1160 11
rect 1082 9 1088 10
rect 1093 9 1105 10
rect 1109 9 1120 10
rect 1127 9 1140 10
rect 1145 9 1160 10
rect 1163 9 1169 23
rect 1175 22 1181 24
rect 1175 18 1180 22
rect 1175 15 1181 18
rect 1175 14 1182 15
rect 1175 13 1183 14
rect 1187 13 1188 14
rect 1176 12 1189 13
rect 1177 10 1189 12
rect 1178 9 1189 10
rect 1191 9 1197 24
rect 1203 9 1208 24
rect 1221 11 1227 38
rect 1271 36 1274 37
rect 1269 32 1274 36
rect 1281 35 1286 40
rect 1294 36 1297 37
rect 1328 36 1331 37
rect 1281 34 1285 35
rect 1292 32 1297 36
rect 1327 35 1331 36
rect 1240 31 1244 32
rect 1256 31 1262 32
rect 1269 31 1275 32
rect 1291 31 1297 32
rect 1326 32 1331 35
rect 1663 33 1669 34
rect 1699 33 1701 34
rect 1716 33 1718 34
rect 1495 32 1505 33
rect 1510 32 1518 33
rect 1525 32 1532 33
rect 1540 32 1549 33
rect 1556 32 1566 33
rect 1574 32 1584 33
rect 1589 32 1597 33
rect 1605 32 1620 33
rect 1630 32 1645 33
rect 1661 32 1671 33
rect 1680 32 1690 33
rect 1699 32 1718 33
rect 1726 32 1736 33
rect 1739 32 1747 33
rect 1326 31 1332 32
rect 1343 31 1348 32
rect 1497 31 1503 32
rect 1512 31 1517 32
rect 1527 31 1533 32
rect 1543 31 1547 32
rect 1558 31 1564 32
rect 1576 31 1583 32
rect 1591 31 1595 32
rect 1232 30 1245 31
rect 1254 30 1263 31
rect 1266 30 1277 31
rect 1231 28 1247 30
rect 1253 29 1263 30
rect 1252 28 1264 29
rect 1231 26 1248 28
rect 1231 24 1238 26
rect 1242 24 1248 26
rect 1221 10 1228 11
rect 1221 9 1227 10
rect 1231 9 1237 24
rect 1243 11 1248 24
rect 1251 26 1263 28
rect 1265 27 1278 30
rect 1266 26 1277 27
rect 1251 24 1257 26
rect 1251 23 1258 24
rect 1251 22 1260 23
rect 1251 21 1262 22
rect 1252 20 1263 21
rect 1253 19 1264 20
rect 1254 18 1264 19
rect 1256 17 1265 18
rect 1258 16 1265 17
rect 1259 14 1265 16
rect 1252 13 1254 14
rect 1258 13 1265 14
rect 1269 16 1274 26
rect 1269 13 1275 16
rect 1251 11 1264 13
rect 1269 12 1278 13
rect 1269 11 1279 12
rect 1243 10 1249 11
rect 1251 10 1263 11
rect 1270 10 1279 11
rect 927 8 931 9
rect 937 8 940 9
rect 949 8 958 9
rect 963 8 969 9
rect 972 8 976 9
rect 984 8 990 9
rect 994 8 998 9
rect 1007 8 1015 9
rect 1024 8 1028 9
rect 1036 8 1040 9
rect 1044 8 1054 9
rect 1070 8 1074 9
rect 1082 8 1087 9
rect 1094 8 1104 9
rect 1110 8 1119 9
rect 1129 8 1139 9
rect 1146 8 1153 9
rect 1156 8 1159 9
rect 1164 8 1168 9
rect 1180 8 1188 9
rect 1192 8 1196 9
rect 1204 8 1207 9
rect 1222 8 1227 9
rect 1232 8 1235 9
rect 1243 8 1248 10
rect 1251 9 1262 10
rect 1271 9 1279 10
rect 1281 9 1286 31
rect 1289 29 1301 31
rect 1288 27 1301 29
rect 1289 26 1301 27
rect 1292 14 1297 26
rect 1304 15 1309 31
rect 1316 30 1320 31
rect 1315 15 1321 30
rect 1323 29 1335 31
rect 1341 30 1350 31
rect 1498 30 1503 31
rect 1340 29 1351 30
rect 1323 28 1336 29
rect 1339 28 1352 29
rect 1323 26 1335 28
rect 1339 27 1353 28
rect 1338 26 1353 27
rect 1304 14 1310 15
rect 1314 14 1321 15
rect 1292 13 1298 14
rect 1304 13 1311 14
rect 1313 13 1321 14
rect 1292 12 1301 13
rect 1304 12 1321 13
rect 1326 16 1331 26
rect 1338 25 1343 26
rect 1348 25 1353 26
rect 1337 22 1343 25
rect 1349 23 1354 25
rect 1348 22 1354 23
rect 1337 19 1355 22
rect 1498 20 1502 30
rect 1513 29 1516 31
rect 1528 30 1534 31
rect 1543 30 1546 31
rect 1528 29 1535 30
rect 1337 17 1354 19
rect 1326 14 1332 16
rect 1337 14 1343 17
rect 1498 16 1503 20
rect 1513 16 1515 29
rect 1528 27 1536 29
rect 1499 15 1504 16
rect 1512 15 1514 16
rect 1351 14 1352 15
rect 1499 14 1505 15
rect 1511 14 1514 15
rect 1528 15 1530 27
rect 1531 26 1537 27
rect 1532 25 1538 26
rect 1533 24 1539 25
rect 1534 23 1540 24
rect 1535 22 1541 23
rect 1535 21 1542 22
rect 1536 20 1543 21
rect 1544 20 1546 30
rect 1537 19 1546 20
rect 1538 18 1546 19
rect 1539 17 1546 18
rect 1540 15 1546 17
rect 1528 14 1531 15
rect 1541 14 1546 15
rect 1559 14 1564 31
rect 1577 30 1582 31
rect 1577 29 1583 30
rect 1578 27 1583 29
rect 1591 29 1594 31
rect 1591 27 1593 29
rect 1579 24 1584 27
rect 1590 25 1592 27
rect 1590 24 1591 25
rect 1580 22 1585 24
rect 1589 22 1591 24
rect 1607 24 1612 32
rect 1617 31 1620 32
rect 1632 31 1638 32
rect 1640 31 1646 32
rect 1660 31 1663 32
rect 1668 31 1671 32
rect 1682 31 1688 32
rect 1618 30 1621 31
rect 1632 30 1637 31
rect 1619 28 1621 30
rect 1617 24 1619 26
rect 1607 22 1619 24
rect 1581 19 1586 22
rect 1588 19 1590 22
rect 1582 17 1589 19
rect 1583 14 1588 17
rect 1607 14 1612 22
rect 1617 20 1619 22
rect 1618 19 1619 20
rect 1633 23 1637 30
rect 1642 28 1647 31
rect 1659 30 1663 31
rect 1659 29 1662 30
rect 1669 29 1671 31
rect 1643 26 1647 28
rect 1658 28 1662 29
rect 1670 28 1671 29
rect 1658 27 1663 28
rect 1658 26 1664 27
rect 1642 24 1647 26
rect 1659 25 1665 26
rect 1659 24 1667 25
rect 1641 23 1646 24
rect 1660 23 1669 24
rect 1633 22 1638 23
rect 1639 22 1644 23
rect 1661 22 1670 23
rect 1633 21 1644 22
rect 1662 21 1671 22
rect 1621 17 1622 18
rect 1620 15 1622 17
rect 1633 15 1637 21
rect 1639 20 1644 21
rect 1664 20 1672 21
rect 1640 19 1645 20
rect 1666 19 1672 20
rect 1640 18 1646 19
rect 1667 18 1672 19
rect 1641 17 1646 18
rect 1658 17 1659 18
rect 1641 16 1647 17
rect 1619 14 1622 15
rect 1326 13 1333 14
rect 1338 13 1345 14
rect 1350 13 1353 14
rect 1500 13 1507 14
rect 1509 13 1513 14
rect 1527 13 1531 14
rect 1542 13 1546 14
rect 1558 13 1564 14
rect 1326 12 1336 13
rect 1338 12 1353 13
rect 1501 12 1512 13
rect 1525 12 1534 13
rect 1543 12 1546 13
rect 1556 12 1566 13
rect 1584 12 1587 14
rect 1606 13 1613 14
rect 1618 13 1622 14
rect 1632 14 1637 15
rect 1642 15 1647 16
rect 1658 16 1660 17
rect 1642 14 1648 15
rect 1658 14 1661 16
rect 1668 15 1672 18
rect 1668 14 1671 15
rect 1683 14 1688 31
rect 1699 31 1702 32
rect 1699 30 1701 31
rect 1699 29 1700 30
rect 1698 28 1700 29
rect 1699 27 1700 28
rect 1706 14 1711 32
rect 1714 31 1718 32
rect 1728 31 1734 32
rect 1715 30 1718 31
rect 1716 28 1718 30
rect 1729 29 1734 31
rect 1741 31 1745 32
rect 1741 30 1744 31
rect 1741 29 1743 30
rect 1730 27 1735 29
rect 1740 27 1742 29
rect 1731 26 1736 27
rect 1732 25 1736 26
rect 1739 25 1741 27
rect 1732 24 1737 25
rect 1738 24 1740 25
rect 1733 23 1740 24
rect 1733 22 1739 23
rect 1734 14 1739 22
rect 1632 13 1638 14
rect 1643 13 1649 14
rect 1658 13 1662 14
rect 1667 13 1670 14
rect 1682 13 1688 14
rect 1705 13 1711 14
rect 1733 13 1739 14
rect 1604 12 1621 13
rect 1630 12 1640 13
rect 1644 12 1650 13
rect 1659 12 1669 13
rect 1680 12 1690 13
rect 1703 12 1714 13
rect 1731 12 1742 13
rect 1293 9 1302 12
rect 1305 10 1321 12
rect 1327 10 1336 12
rect 1339 11 1353 12
rect 1502 11 1510 12
rect 1544 11 1546 12
rect 1584 11 1586 12
rect 1647 11 1650 12
rect 1661 11 1667 12
rect 1340 10 1353 11
rect 1306 9 1321 10
rect 1328 9 1336 10
rect 1341 9 1353 10
rect 1252 8 1261 9
rect 1271 8 1278 9
rect 1282 8 1285 9
rect 1294 8 1301 9
rect 1307 8 1314 9
rect 1317 8 1320 9
rect 1329 8 1335 9
rect 1342 8 1352 9
<< end >>
