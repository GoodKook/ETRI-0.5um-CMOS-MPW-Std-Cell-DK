magic
tech scmos
timestamp 1740666625
<< end >>
