magic
tech scmos
magscale 1 2
timestamp 1724155847
<< metal1 >>
rect -63 5218 -3 5478
rect 5810 5462 5903 5478
rect 3167 5413 3173 5427
rect 1467 5397 1493 5403
rect 2727 5397 2813 5403
rect 3300 5383 3313 5387
rect 3297 5373 3313 5383
rect 3297 5343 3303 5373
rect 3277 5337 3303 5343
rect 3277 5327 3283 5337
rect 3267 5317 3283 5327
rect 3267 5313 3280 5317
rect 5347 5317 5413 5323
rect 1707 5277 1773 5283
rect -63 5202 30 5218
rect -63 4698 -3 5202
rect 4767 5097 4833 5103
rect 60 5083 73 5087
rect 57 5073 73 5083
rect 1653 5083 1667 5093
rect 1653 5080 1683 5083
rect 1657 5077 1683 5080
rect 57 5047 63 5073
rect 57 5037 73 5047
rect 60 5033 73 5037
rect 1677 5043 1683 5077
rect 1917 5047 1923 5073
rect 1677 5040 1703 5043
rect 1677 5037 1707 5040
rect 1693 5027 1707 5037
rect 1907 5033 1933 5047
rect 5843 4958 5903 5462
rect 5810 4942 5903 4958
rect 3107 4897 3133 4903
rect 1113 4883 1127 4893
rect 5727 4897 5773 4903
rect 1113 4880 1173 4883
rect 1117 4877 1173 4880
rect 2927 4877 2963 4883
rect 1127 4857 1153 4863
rect 1260 4863 1273 4867
rect 1257 4853 1273 4863
rect 1400 4863 1413 4867
rect 1397 4853 1413 4863
rect 1257 4827 1263 4853
rect 1257 4817 1273 4827
rect 1260 4813 1273 4817
rect 127 4797 193 4803
rect 1397 4803 1403 4853
rect 2957 4827 2963 4877
rect 3100 4863 3113 4867
rect 2947 4817 2963 4827
rect 3097 4853 3113 4863
rect 3220 4863 3233 4867
rect 3217 4853 3233 4863
rect 3600 4863 3613 4867
rect 3597 4853 3613 4863
rect 5727 4863 5740 4867
rect 5727 4853 5743 4863
rect 3097 4827 3103 4853
rect 3097 4817 3113 4827
rect 2947 4813 2960 4817
rect 3100 4813 3113 4817
rect 1347 4797 1403 4803
rect 3217 4803 3223 4853
rect 3597 4827 3603 4853
rect 5737 4827 5743 4853
rect 3587 4817 3603 4827
rect 3587 4813 3600 4817
rect 5727 4817 5743 4827
rect 5727 4813 5740 4817
rect 3217 4797 3253 4803
rect -63 4682 30 4698
rect -63 4178 -3 4682
rect 4447 4597 4513 4603
rect 1747 4577 1793 4583
rect 2367 4577 2413 4583
rect 2587 4577 2673 4583
rect 4517 4577 4553 4583
rect 1507 4563 1520 4567
rect 1613 4563 1627 4573
rect 1507 4553 1523 4563
rect 1613 4560 1643 4563
rect 1617 4557 1643 4560
rect 1517 4527 1523 4553
rect 1637 4527 1643 4557
rect 1727 4563 1740 4567
rect 3200 4566 3220 4567
rect 1727 4553 1743 4563
rect 1517 4517 1533 4527
rect 1520 4513 1533 4517
rect 1637 4517 1653 4527
rect 1640 4513 1653 4517
rect 1737 4526 1743 4553
rect 3207 4563 3220 4566
rect 3460 4563 3473 4567
rect 3207 4553 3223 4563
rect 3217 4527 3223 4553
rect 3457 4553 3473 4563
rect 3947 4563 3960 4567
rect 3947 4553 3963 4563
rect 4247 4557 4273 4563
rect 4467 4563 4480 4567
rect 4517 4563 4523 4577
rect 4880 4563 4893 4567
rect 4467 4553 4483 4563
rect 3207 4517 3223 4527
rect 3207 4513 3220 4517
rect 3457 4523 3463 4553
rect 3427 4517 3463 4523
rect 3957 4527 3963 4553
rect 3957 4517 3973 4527
rect 3960 4513 3973 4517
rect 4477 4503 4483 4553
rect 4497 4557 4523 4563
rect 4497 4527 4503 4557
rect 4877 4553 4893 4563
rect 5620 4563 5633 4567
rect 5617 4553 5633 4563
rect 4877 4527 4883 4553
rect 5617 4527 5623 4553
rect 4497 4517 4513 4527
rect 4500 4513 4513 4517
rect 4877 4517 4893 4527
rect 4880 4513 4893 4517
rect 5607 4517 5623 4527
rect 5607 4513 5620 4517
rect 4447 4497 4483 4503
rect 2380 4486 2393 4487
rect 2387 4473 2393 4486
rect 3927 4477 3993 4483
rect 5027 4477 5073 4483
rect 5843 4438 5903 4942
rect 5810 4422 5903 4438
rect 5707 4383 5720 4387
rect 5707 4373 5723 4383
rect 967 4357 1013 4363
rect 247 4343 260 4347
rect 247 4333 263 4343
rect 627 4343 640 4347
rect 4020 4343 4033 4347
rect 627 4333 643 4343
rect 257 4307 263 4333
rect 637 4307 643 4333
rect 4017 4333 4033 4343
rect 4980 4343 4993 4347
rect 4977 4333 4993 4343
rect 5187 4343 5200 4347
rect 5187 4333 5203 4343
rect 4017 4307 4023 4333
rect 257 4297 273 4307
rect 260 4293 273 4297
rect 637 4297 653 4307
rect 640 4293 653 4297
rect 4007 4297 4023 4307
rect 4007 4293 4020 4297
rect 1327 4277 1373 4283
rect 1827 4277 1913 4283
rect 3127 4277 3153 4283
rect 4977 4283 4983 4333
rect 5197 4307 5203 4333
rect 5197 4297 5213 4307
rect 5200 4293 5213 4297
rect 5717 4303 5723 4373
rect 5717 4297 5743 4303
rect 4927 4277 4983 4283
rect 5167 4277 5193 4283
rect 3987 4257 4053 4263
rect 5737 4246 5743 4297
rect -63 4162 30 4178
rect -63 3658 -3 4162
rect 507 4057 553 4063
rect 2507 4057 2613 4063
rect 3307 4057 3353 4063
rect 3427 4057 3473 4063
rect 3927 4057 3993 4063
rect 5087 4057 5113 4063
rect 5207 4057 5233 4063
rect 5740 4063 5753 4067
rect 5737 4053 5753 4063
rect 320 4043 333 4047
rect 317 4033 333 4043
rect 407 4043 420 4047
rect 3060 4043 3073 4047
rect 407 4033 423 4043
rect 317 4007 323 4033
rect 307 3997 323 4007
rect 417 4003 423 4033
rect 3057 4033 3073 4043
rect 3947 4043 3960 4047
rect 3947 4033 3963 4043
rect 5367 4043 5380 4047
rect 5737 4043 5743 4053
rect 5367 4033 5383 4043
rect 3057 4007 3063 4033
rect 3957 4007 3963 4033
rect 5377 4007 5383 4033
rect 417 3997 443 4003
rect 3057 3997 3073 4007
rect 307 3993 320 3997
rect 437 3987 443 3997
rect 3060 3993 3073 3997
rect 3947 3997 3963 4007
rect 3947 3993 3960 3997
rect 5367 3997 5383 4007
rect 5717 4037 5743 4043
rect 5717 4007 5723 4037
rect 5717 3997 5733 4007
rect 5367 3993 5380 3997
rect 5720 3993 5733 3997
rect 437 3977 453 3987
rect 440 3973 453 3977
rect 3927 3957 3973 3963
rect 5843 3918 5903 4422
rect 5810 3902 5903 3918
rect 1567 3837 1633 3843
rect 2287 3837 2333 3843
rect 547 3823 560 3827
rect 700 3823 713 3827
rect 547 3813 563 3823
rect 557 3787 563 3813
rect 547 3777 563 3787
rect 697 3813 713 3823
rect 827 3823 840 3827
rect 827 3813 843 3823
rect 1327 3817 1353 3823
rect 1467 3823 1480 3827
rect 1467 3813 1483 3823
rect 1867 3823 1880 3827
rect 2040 3823 2053 3827
rect 1867 3813 1883 3823
rect 697 3787 703 3813
rect 837 3787 843 3813
rect 1477 3787 1483 3813
rect 697 3777 713 3787
rect 547 3773 560 3777
rect 700 3773 713 3777
rect 837 3777 853 3787
rect 840 3773 853 3777
rect 1467 3777 1483 3787
rect 1877 3787 1883 3813
rect 2037 3813 2053 3823
rect 3880 3823 3893 3827
rect 3877 3813 3893 3823
rect 5413 3823 5427 3833
rect 5397 3820 5427 3823
rect 5397 3817 5423 3820
rect 1877 3777 1893 3787
rect 1467 3773 1480 3777
rect 1880 3773 1893 3777
rect 2037 3783 2043 3813
rect 2017 3780 2043 3783
rect 2013 3777 2043 3780
rect 3877 3787 3883 3813
rect 4613 3787 4627 3793
rect 5397 3787 5403 3817
rect 5787 3823 5800 3827
rect 5787 3813 5803 3823
rect 5797 3787 5803 3813
rect 3877 3777 3893 3787
rect 2013 3767 2027 3777
rect 3880 3773 3893 3777
rect 4613 3780 4633 3787
rect 4617 3777 4633 3780
rect 4620 3773 4633 3777
rect 5387 3777 5403 3787
rect 5387 3773 5400 3777
rect 5787 3777 5803 3787
rect 5787 3773 5800 3777
rect 647 3757 753 3763
rect -63 3642 30 3658
rect -63 3138 -3 3642
rect 5647 3557 5713 3563
rect 1587 3537 1623 3543
rect 1617 3487 1623 3537
rect 5107 3537 5143 3543
rect 5137 3523 5143 3537
rect 5137 3517 5163 3523
rect 5157 3487 5163 3517
rect 5417 3517 5453 3523
rect 5417 3487 5423 3517
rect 1607 3477 1623 3487
rect 1607 3473 1620 3477
rect 2067 3477 2093 3483
rect 5147 3477 5163 3487
rect 5147 3473 5160 3477
rect 5407 3477 5423 3487
rect 5677 3487 5683 3533
rect 5787 3517 5813 3523
rect 5677 3477 5693 3487
rect 5407 3473 5420 3477
rect 5680 3473 5693 3477
rect 3987 3457 4033 3463
rect 5843 3398 5903 3902
rect 5810 3382 5903 3398
rect 1247 3357 1273 3363
rect 1067 3337 1133 3343
rect 647 3317 673 3323
rect 4737 3317 4773 3323
rect 167 3297 193 3303
rect 957 3297 993 3303
rect 957 3247 963 3297
rect 4737 3303 4743 3317
rect 4860 3303 4873 3307
rect 4717 3297 4743 3303
rect 4717 3267 4723 3297
rect 4707 3257 4723 3267
rect 4857 3293 4873 3303
rect 4857 3263 4863 3293
rect 4837 3260 4863 3263
rect 4833 3257 4863 3260
rect 4707 3253 4720 3257
rect 4833 3247 4847 3257
rect 287 3237 313 3243
rect 3247 3237 3313 3243
rect 5347 3237 5453 3243
rect -63 3122 30 3138
rect -63 2618 -3 3122
rect 3407 3017 3513 3023
rect 1287 3003 1300 3007
rect 1287 2993 1303 3003
rect 1297 2967 1303 2993
rect 1287 2957 1303 2967
rect 1287 2953 1300 2957
rect 5347 2937 5393 2943
rect 5407 2937 5453 2943
rect 5843 2878 5903 3382
rect 5810 2862 5903 2878
rect 4913 2823 4927 2833
rect 4913 2820 4973 2823
rect 4917 2817 4973 2820
rect 2607 2797 2633 2803
rect 1420 2783 1433 2787
rect 1417 2773 1433 2783
rect 1647 2783 1660 2787
rect 2173 2783 2187 2793
rect 1647 2773 1663 2783
rect 1417 2743 1423 2773
rect 1387 2737 1423 2743
rect 1657 2747 1663 2773
rect 2157 2780 2187 2783
rect 2157 2777 2183 2780
rect 2157 2747 2163 2777
rect 1657 2737 1673 2747
rect 1660 2733 1673 2737
rect 2147 2737 2163 2747
rect 2147 2733 2160 2737
rect 5787 2737 5813 2743
rect 4087 2717 4113 2723
rect -63 2602 30 2618
rect -63 2098 -3 2602
rect 2867 2517 2913 2523
rect 5107 2497 5143 2503
rect 3560 2483 3573 2487
rect 3557 2473 3573 2483
rect 4587 2483 4600 2487
rect 4720 2483 4733 2487
rect 4587 2473 4603 2483
rect 3557 2443 3563 2473
rect 4597 2447 4603 2473
rect 4717 2473 4733 2483
rect 4827 2483 4840 2487
rect 4827 2473 4843 2483
rect 4967 2483 4980 2487
rect 5137 2483 5143 2497
rect 5767 2497 5803 2503
rect 4967 2473 4983 2483
rect 5137 2477 5163 2483
rect 4717 2447 4723 2473
rect 3527 2437 3563 2443
rect 4587 2437 4603 2447
rect 4587 2433 4600 2437
rect 4707 2437 4723 2447
rect 4837 2447 4843 2473
rect 4837 2437 4853 2447
rect 4707 2433 4720 2437
rect 4840 2433 4853 2437
rect 4977 2443 4983 2473
rect 5157 2447 5163 2477
rect 5553 2447 5567 2453
rect 5797 2447 5803 2497
rect 4977 2437 5013 2443
rect 5147 2437 5163 2447
rect 5147 2433 5160 2437
rect 5247 2437 5293 2443
rect 5547 2440 5567 2447
rect 5547 2437 5563 2440
rect 5547 2433 5560 2437
rect 5787 2437 5803 2447
rect 5787 2433 5800 2437
rect 5843 2358 5903 2862
rect 5810 2342 5903 2358
rect 1227 2277 1313 2283
rect 3907 2277 3953 2283
rect 4447 2277 4473 2283
rect 4487 2277 4533 2283
rect 2060 2263 2073 2267
rect 2057 2253 2073 2263
rect 3560 2263 3573 2267
rect 3557 2253 3573 2263
rect 3820 2263 3833 2267
rect 3817 2253 3833 2263
rect 4220 2263 4233 2267
rect 4217 2253 4233 2263
rect 4347 2263 4360 2267
rect 4347 2253 4363 2263
rect 4597 2263 4603 2293
rect 5467 2277 5513 2283
rect 4467 2257 4503 2263
rect 4597 2257 4623 2263
rect 2057 2223 2063 2253
rect 2037 2217 2063 2223
rect 2333 2227 2347 2233
rect 3557 2227 3563 2253
rect 3817 2227 3823 2253
rect 2333 2220 2353 2227
rect 2337 2217 2353 2220
rect 2037 2207 2043 2217
rect 2340 2213 2353 2217
rect 3557 2217 3573 2227
rect 3560 2213 3573 2217
rect 3807 2217 3823 2227
rect 4217 2227 4223 2253
rect 4357 2227 4363 2253
rect 4497 2227 4503 2257
rect 4617 2227 4623 2257
rect 4887 2263 4900 2267
rect 4887 2253 4903 2263
rect 5027 2263 5040 2267
rect 5200 2263 5213 2267
rect 5027 2253 5043 2263
rect 4217 2217 4233 2227
rect 3807 2213 3820 2217
rect 4220 2213 4233 2217
rect 4357 2217 4373 2227
rect 4360 2213 4373 2217
rect 4497 2217 4513 2227
rect 4500 2213 4513 2217
rect 4607 2217 4623 2227
rect 4897 2227 4903 2253
rect 5037 2227 5043 2253
rect 4897 2217 4913 2227
rect 4607 2213 4620 2217
rect 4900 2213 4913 2217
rect 5027 2217 5043 2227
rect 5197 2253 5213 2263
rect 5447 2263 5460 2267
rect 5447 2253 5463 2263
rect 5197 2227 5203 2253
rect 5197 2217 5213 2227
rect 5027 2213 5040 2217
rect 5200 2213 5213 2217
rect 5457 2223 5463 2253
rect 5457 2217 5483 2223
rect 2027 2197 2043 2207
rect 2027 2193 2040 2197
rect 3407 2197 3473 2203
rect 3647 2197 3683 2203
rect 3677 2183 3683 2197
rect 3787 2197 3853 2203
rect 4447 2197 4473 2203
rect 5477 2203 5483 2217
rect 5613 2223 5627 2233
rect 5587 2220 5627 2223
rect 5587 2217 5623 2220
rect 5477 2197 5533 2203
rect 3677 2177 3733 2183
rect 5697 2167 5703 2193
rect 4587 2157 4633 2163
rect -63 2082 30 2098
rect -63 1578 -3 2082
rect 4607 2017 4633 2023
rect 187 1977 253 1983
rect 1447 1977 1483 1983
rect 680 1963 693 1967
rect 677 1953 693 1963
rect 1087 1963 1100 1967
rect 1087 1953 1103 1963
rect 1347 1963 1360 1967
rect 1477 1963 1483 1977
rect 1587 1977 1613 1983
rect 1887 1977 1933 1983
rect 3047 1977 3093 1983
rect 3577 1977 3633 1983
rect 1620 1963 1633 1967
rect 1347 1953 1363 1963
rect 1477 1957 1503 1963
rect 677 1927 683 1953
rect 667 1917 683 1927
rect 1097 1927 1103 1953
rect 1357 1927 1363 1953
rect 1497 1927 1503 1957
rect 1097 1917 1113 1927
rect 667 1913 680 1917
rect 1100 1913 1113 1917
rect 1357 1917 1373 1927
rect 1360 1913 1373 1917
rect 1487 1917 1503 1927
rect 1617 1953 1633 1963
rect 1767 1963 1780 1967
rect 1880 1963 1893 1967
rect 1767 1953 1783 1963
rect 1617 1927 1623 1953
rect 1617 1917 1633 1927
rect 1487 1913 1500 1917
rect 1620 1913 1633 1917
rect 1777 1903 1783 1953
rect 1877 1953 1893 1963
rect 2420 1963 2433 1967
rect 2417 1953 2433 1963
rect 2937 1957 2973 1963
rect 1877 1927 1883 1953
rect 2417 1927 2423 1953
rect 2937 1927 2943 1957
rect 1877 1917 1893 1927
rect 1880 1913 1893 1917
rect 2407 1917 2423 1927
rect 2407 1913 2420 1917
rect 2927 1917 2943 1927
rect 2927 1913 2940 1917
rect 1777 1897 1813 1903
rect 3577 1867 3583 1977
rect 4607 1977 4693 1983
rect 5327 1977 5393 1983
rect 5767 1977 5813 1983
rect 3600 1963 3613 1967
rect 3597 1953 3613 1963
rect 3727 1963 3740 1967
rect 3880 1963 3893 1967
rect 3727 1953 3743 1963
rect 3597 1887 3603 1953
rect 3737 1927 3743 1953
rect 3727 1917 3743 1927
rect 3877 1953 3893 1963
rect 4140 1963 4153 1967
rect 4137 1953 4153 1963
rect 4260 1963 4273 1967
rect 4257 1953 4273 1963
rect 4767 1963 4780 1967
rect 4767 1953 4783 1963
rect 5027 1963 5040 1967
rect 5027 1953 5043 1963
rect 5307 1963 5320 1967
rect 5307 1953 5323 1963
rect 3727 1913 3740 1917
rect 3877 1887 3883 1953
rect 4137 1903 4143 1953
rect 4257 1927 4263 1953
rect 4247 1917 4263 1927
rect 4517 1927 4523 1953
rect 4777 1927 4783 1953
rect 5037 1927 5043 1953
rect 5317 1927 5323 1953
rect 4517 1917 4533 1927
rect 4247 1913 4260 1917
rect 4520 1913 4533 1917
rect 4777 1917 4793 1927
rect 4780 1913 4793 1917
rect 5037 1917 5053 1927
rect 5040 1913 5053 1917
rect 5307 1917 5323 1927
rect 5307 1913 5320 1917
rect 4137 1897 4173 1903
rect 3877 1877 3893 1887
rect 3880 1873 3893 1877
rect 4947 1877 4973 1883
rect 5843 1838 5903 2342
rect 5810 1822 5903 1838
rect 2027 1743 2040 1747
rect 2027 1733 2043 1743
rect 2327 1743 2340 1747
rect 2327 1733 2343 1743
rect 2447 1743 2460 1747
rect 2560 1743 2573 1747
rect 2447 1733 2463 1743
rect 2037 1707 2043 1733
rect 2027 1697 2043 1707
rect 2027 1693 2040 1697
rect 287 1677 413 1683
rect 2167 1677 2253 1683
rect 2337 1683 2343 1733
rect 2457 1707 2463 1733
rect 2447 1697 2463 1707
rect 2557 1733 2573 1743
rect 2827 1743 2840 1747
rect 2827 1733 2843 1743
rect 2557 1707 2563 1733
rect 2557 1697 2573 1707
rect 2447 1693 2460 1697
rect 2560 1693 2573 1697
rect 2837 1703 2843 1733
rect 2817 1697 2843 1703
rect 2817 1687 2823 1697
rect 2307 1677 2343 1683
rect 2807 1677 2823 1687
rect 2857 1687 2863 1753
rect 3220 1743 3233 1747
rect 3217 1733 3233 1743
rect 3347 1743 3360 1747
rect 3780 1743 3793 1747
rect 3347 1733 3363 1743
rect 3217 1707 3223 1733
rect 3357 1707 3363 1733
rect 3777 1733 3793 1743
rect 3920 1746 3940 1747
rect 3920 1743 3933 1746
rect 3917 1733 3933 1743
rect 3777 1707 3783 1733
rect 3917 1707 3923 1733
rect 4047 1743 4060 1747
rect 4047 1733 4063 1743
rect 4147 1743 4160 1747
rect 4273 1743 4287 1752
rect 4147 1733 4163 1743
rect 4273 1740 4313 1743
rect 4277 1737 4313 1740
rect 4427 1743 4440 1747
rect 4560 1743 4573 1747
rect 4427 1733 4443 1743
rect 3217 1697 3233 1707
rect 3220 1693 3233 1697
rect 3347 1697 3363 1707
rect 3347 1693 3360 1697
rect 3767 1697 3783 1707
rect 3767 1693 3780 1697
rect 3907 1697 3923 1707
rect 4057 1707 4063 1733
rect 4157 1707 4163 1733
rect 4057 1697 4073 1707
rect 3907 1693 3920 1697
rect 4060 1693 4073 1697
rect 4147 1697 4163 1707
rect 4437 1703 4443 1733
rect 4557 1733 4573 1743
rect 4800 1743 4813 1747
rect 4797 1733 4813 1743
rect 5100 1743 5113 1747
rect 4927 1737 4963 1743
rect 4557 1707 4563 1733
rect 4437 1697 4463 1703
rect 4557 1697 4573 1707
rect 4147 1693 4160 1697
rect 4457 1687 4463 1697
rect 4560 1693 4573 1697
rect 2857 1677 2873 1687
rect 2807 1673 2820 1677
rect 2860 1673 2873 1677
rect 3147 1677 3173 1683
rect 3867 1677 3933 1683
rect 4457 1677 4473 1687
rect 4460 1673 4473 1677
rect 4797 1683 4803 1733
rect 4957 1707 4963 1737
rect 5097 1733 5113 1743
rect 5220 1743 5233 1747
rect 5217 1733 5233 1743
rect 5640 1743 5653 1747
rect 5637 1733 5653 1743
rect 5097 1707 5103 1733
rect 4957 1697 4973 1707
rect 4960 1693 4973 1697
rect 5087 1697 5103 1707
rect 5217 1707 5223 1733
rect 5637 1707 5643 1733
rect 5217 1697 5233 1707
rect 5087 1693 5100 1697
rect 5220 1693 5233 1697
rect 5637 1697 5653 1707
rect 5640 1693 5653 1697
rect 4767 1677 4803 1683
rect 4127 1657 4213 1663
rect 5327 1637 5373 1643
rect -63 1562 30 1578
rect -63 1058 -3 1562
rect 3867 1537 3893 1543
rect 4347 1477 4413 1483
rect 5707 1477 5773 1483
rect 127 1457 193 1463
rect 2267 1457 2313 1463
rect 2667 1457 2733 1463
rect 4087 1463 4100 1467
rect 4087 1453 4103 1463
rect 1340 1443 1353 1447
rect 1337 1433 1353 1443
rect 1587 1443 1600 1447
rect 1587 1433 1603 1443
rect 2127 1443 2140 1447
rect 2560 1443 2573 1447
rect 2127 1433 2143 1443
rect 1337 1407 1343 1433
rect 1597 1407 1603 1433
rect 2137 1407 2143 1433
rect 2557 1433 2573 1443
rect 2820 1443 2833 1447
rect 2817 1433 2833 1443
rect 4097 1443 4103 1453
rect 4477 1457 4533 1463
rect 4477 1447 4483 1457
rect 5697 1457 5753 1463
rect 4097 1437 4123 1443
rect 2557 1407 2563 1433
rect 2817 1407 2823 1433
rect 1337 1397 1353 1407
rect 1340 1393 1353 1397
rect 1597 1397 1613 1407
rect 1600 1393 1613 1397
rect 2137 1397 2153 1407
rect 2140 1393 2153 1397
rect 2557 1397 2573 1407
rect 2560 1393 2573 1397
rect 2807 1397 2823 1407
rect 4117 1407 4123 1437
rect 4487 1443 4500 1447
rect 5080 1443 5093 1447
rect 4487 1433 4503 1443
rect 4497 1407 4503 1433
rect 4117 1397 4133 1407
rect 2807 1393 2820 1397
rect 4120 1393 4133 1397
rect 4487 1397 4503 1407
rect 5077 1433 5093 1443
rect 5540 1443 5553 1447
rect 5537 1433 5553 1443
rect 5077 1407 5083 1433
rect 5537 1407 5543 1433
rect 5077 1397 5093 1407
rect 4487 1393 4500 1397
rect 5080 1393 5093 1397
rect 5527 1397 5543 1407
rect 5697 1407 5703 1457
rect 5697 1397 5713 1407
rect 5527 1393 5540 1397
rect 5700 1393 5713 1397
rect 5207 1377 5233 1383
rect 5407 1377 5453 1383
rect 4253 1343 4267 1353
rect 4207 1340 4267 1343
rect 4207 1337 4263 1340
rect 5843 1318 5903 1822
rect 5810 1302 5903 1318
rect 167 1237 233 1243
rect 847 1237 873 1243
rect 1327 1237 1393 1243
rect 1487 1237 1533 1243
rect 2140 1223 2153 1227
rect 2137 1213 2153 1223
rect 2273 1223 2287 1233
rect 2257 1220 2287 1223
rect 3997 1237 4053 1243
rect 2257 1217 2283 1220
rect 2137 1183 2143 1213
rect 2257 1187 2263 1217
rect 2137 1177 2163 1183
rect 2157 1167 2163 1177
rect 2247 1177 2263 1187
rect 3733 1187 3747 1193
rect 3997 1187 4003 1237
rect 4767 1237 4793 1243
rect 4257 1217 4293 1223
rect 3733 1180 3753 1187
rect 3737 1177 3753 1180
rect 2247 1173 2260 1177
rect 3740 1173 3753 1177
rect 3997 1177 4013 1187
rect 4000 1173 4013 1177
rect 4257 1167 4263 1217
rect 4687 1223 4700 1227
rect 4687 1213 4703 1223
rect 4907 1223 4920 1227
rect 4907 1213 4923 1223
rect 4697 1187 4703 1213
rect 4687 1177 4703 1187
rect 4917 1183 4923 1213
rect 5057 1187 5063 1233
rect 5447 1220 5503 1223
rect 5447 1217 5507 1220
rect 5493 1207 5507 1217
rect 4917 1177 4953 1183
rect 4687 1173 4700 1177
rect 5057 1177 5073 1187
rect 5060 1173 5073 1177
rect 807 1157 873 1163
rect 1507 1157 1573 1163
rect 1627 1157 1673 1163
rect 2157 1163 2173 1167
rect 2107 1157 2173 1163
rect 2160 1153 2173 1157
rect 2367 1157 2413 1163
rect 3527 1157 3573 1163
rect 3847 1157 3913 1163
rect 4247 1157 4263 1167
rect 4247 1153 4260 1157
rect 407 1137 433 1143
rect 3247 1137 3313 1143
rect -63 1042 30 1058
rect -63 538 -3 1042
rect 987 977 1033 983
rect 1187 977 1213 983
rect 567 957 593 963
rect 1527 957 1613 963
rect 2393 963 2407 973
rect 2393 960 2473 963
rect 2397 957 2473 960
rect 107 937 213 943
rect 1107 937 1173 943
rect 1547 937 1613 943
rect 3587 937 3653 943
rect 320 923 333 927
rect 317 913 333 923
rect 2307 923 2320 927
rect 2307 913 2323 923
rect 2427 923 2440 927
rect 2427 913 2443 923
rect 173 887 187 893
rect 317 887 323 913
rect 173 880 193 887
rect 177 877 193 880
rect 180 873 193 877
rect 307 877 323 887
rect 307 873 320 877
rect 127 857 173 863
rect 2317 863 2323 913
rect 2437 886 2443 913
rect 2677 917 2713 923
rect 2677 866 2683 917
rect 3080 923 3093 927
rect 3077 913 3093 923
rect 3367 923 3380 927
rect 3533 923 3547 933
rect 4267 937 4373 943
rect 5447 937 5493 943
rect 5547 937 5673 943
rect 3367 913 3383 923
rect 3077 887 3083 913
rect 3067 877 3083 887
rect 3377 887 3383 913
rect 3517 920 3547 923
rect 3517 917 3543 920
rect 3377 877 3393 887
rect 3067 873 3080 877
rect 3380 873 3393 877
rect 2287 857 2323 863
rect 3517 863 3523 917
rect 4677 906 4683 933
rect 5087 923 5100 927
rect 5240 923 5253 927
rect 5087 913 5103 923
rect 5097 887 5103 913
rect 5237 913 5253 923
rect 5360 923 5373 927
rect 5357 913 5373 923
rect 5237 887 5243 913
rect 5357 887 5363 913
rect 5097 877 5113 887
rect 5100 873 5113 877
rect 5237 877 5253 887
rect 5240 873 5253 877
rect 5347 877 5363 887
rect 5347 873 5360 877
rect 3467 857 3523 863
rect 5843 798 5903 1302
rect 5810 782 5903 798
rect 117 703 123 733
rect 147 717 193 723
rect 117 697 143 703
rect 137 667 143 697
rect 407 703 420 707
rect 673 703 687 713
rect 713 703 727 713
rect 2277 717 2313 723
rect 407 693 423 703
rect 673 700 727 703
rect 677 697 723 700
rect 137 657 153 667
rect 140 653 153 657
rect 417 663 423 693
rect 697 667 703 697
rect 827 703 840 707
rect 1400 703 1413 707
rect 827 693 843 703
rect 837 667 843 693
rect 397 657 423 663
rect 397 643 403 657
rect 687 657 703 667
rect 687 653 700 657
rect 827 657 843 667
rect 1397 693 1413 703
rect 1527 703 1540 707
rect 1680 703 1693 707
rect 1527 693 1543 703
rect 827 653 840 657
rect 367 637 403 643
rect 487 637 553 643
rect 1397 643 1403 693
rect 1537 667 1543 693
rect 1677 693 1693 703
rect 1840 703 1853 707
rect 1837 693 1853 703
rect 1980 703 1993 707
rect 1977 693 1993 703
rect 2120 703 2133 707
rect 2117 693 2133 703
rect 1677 667 1683 693
rect 1837 683 1843 693
rect 1817 677 1843 683
rect 1817 667 1823 677
rect 1977 667 1983 693
rect 1527 657 1543 667
rect 1527 653 1540 657
rect 1667 657 1683 667
rect 1667 653 1680 657
rect 1807 657 1823 667
rect 1807 653 1820 657
rect 1967 657 1983 667
rect 2117 667 2123 693
rect 2277 667 2283 717
rect 2507 703 2520 707
rect 2507 693 2523 703
rect 2787 703 2800 707
rect 2787 693 2803 703
rect 2927 703 2940 707
rect 2927 693 2943 703
rect 3067 703 3080 707
rect 3100 703 3113 707
rect 3067 693 3083 703
rect 2517 667 2523 693
rect 2797 667 2803 693
rect 2117 657 2133 667
rect 1967 653 1980 657
rect 2120 653 2133 657
rect 2277 657 2293 667
rect 2280 653 2293 657
rect 2517 657 2533 667
rect 2520 653 2533 657
rect 2797 657 2813 667
rect 2800 653 2813 657
rect 2937 663 2943 693
rect 3077 667 3083 693
rect 2937 657 2963 663
rect 1347 637 1403 643
rect 1767 637 1833 643
rect 2087 637 2153 643
rect 2227 637 2273 643
rect 2487 637 2593 643
rect 2957 643 2963 657
rect 3067 657 3083 667
rect 3097 693 3113 703
rect 3227 703 3240 707
rect 3380 703 3393 707
rect 3227 693 3243 703
rect 3097 667 3103 693
rect 3237 667 3243 693
rect 3377 693 3393 703
rect 3467 703 3480 707
rect 4440 703 4453 707
rect 3467 693 3483 703
rect 3377 667 3383 693
rect 3477 667 3483 693
rect 4437 693 4453 703
rect 5140 703 5153 707
rect 5137 693 5153 703
rect 5420 703 5433 707
rect 5417 693 5433 703
rect 5547 703 5560 707
rect 5547 693 5563 703
rect 4437 667 4443 693
rect 3097 657 3113 667
rect 3067 653 3080 657
rect 3100 653 3113 657
rect 3227 657 3243 667
rect 3227 653 3240 657
rect 3367 657 3383 667
rect 3367 653 3380 657
rect 3467 657 3483 667
rect 3467 653 3480 657
rect 4427 657 4443 667
rect 5137 667 5143 693
rect 5137 657 5153 667
rect 4427 653 4440 657
rect 5140 653 5153 657
rect 5417 663 5423 693
rect 5557 667 5563 693
rect 5397 657 5423 663
rect 2957 637 3013 643
rect 3967 637 3993 643
rect 4107 637 4153 643
rect 4167 637 4213 643
rect 4367 637 4473 643
rect 5397 643 5403 657
rect 5547 657 5563 667
rect 5547 653 5560 657
rect 5347 637 5403 643
rect -63 522 30 538
rect -63 18 -3 522
rect 267 417 353 423
rect 847 417 893 423
rect 1187 417 1213 423
rect 1497 417 1533 423
rect 200 403 213 407
rect 197 393 213 403
rect 1497 403 1503 417
rect 1637 417 1673 423
rect 1637 403 1643 417
rect 2127 417 2233 423
rect 2807 417 2863 423
rect 1477 397 1503 403
rect 1617 397 1643 403
rect 197 367 203 393
rect 1477 367 1483 397
rect 1617 367 1623 397
rect 1847 403 1860 407
rect 2300 403 2313 407
rect 1847 393 1863 403
rect 1857 367 1863 393
rect 197 357 213 367
rect 200 353 213 357
rect 1467 357 1483 367
rect 1467 353 1480 357
rect 1607 357 1623 367
rect 1607 353 1620 357
rect 1847 357 1863 367
rect 2297 393 2313 403
rect 2707 403 2720 407
rect 2707 393 2723 403
rect 2297 367 2303 393
rect 2717 367 2723 393
rect 2857 367 2863 417
rect 3087 417 3123 423
rect 2987 403 3000 407
rect 3117 403 3123 417
rect 4567 417 4673 423
rect 5133 403 5147 413
rect 2987 393 3003 403
rect 3117 397 3143 403
rect 5133 400 5163 403
rect 5137 397 5163 400
rect 2997 367 3003 393
rect 2297 357 2313 367
rect 1847 353 1860 357
rect 2300 353 2313 357
rect 2707 357 2723 367
rect 2707 353 2720 357
rect 2847 357 2863 367
rect 2847 353 2860 357
rect 2987 357 3003 367
rect 2987 353 3000 357
rect 3137 343 3143 397
rect 5157 367 5163 397
rect 5147 357 5163 367
rect 5437 363 5443 413
rect 5417 357 5443 363
rect 5147 353 5160 357
rect 3107 337 3143 343
rect 3407 337 3453 343
rect 5417 343 5423 357
rect 5387 337 5423 343
rect 3147 326 3160 327
rect 3147 313 3153 326
rect 5843 278 5903 782
rect 5810 262 5903 278
rect 2327 237 2353 243
rect 1327 217 1373 223
rect 5327 217 5353 223
rect 2617 197 2693 203
rect 1100 183 1113 187
rect 1097 173 1113 183
rect 2200 183 2213 187
rect 2197 173 2213 183
rect 1097 143 1103 173
rect 2197 143 2203 173
rect 1077 137 1103 143
rect 2177 137 2203 143
rect 2617 143 2623 197
rect 5067 197 5133 203
rect 2747 183 2760 187
rect 3820 183 3833 187
rect 2747 180 2763 183
rect 2747 173 2767 180
rect 2753 166 2767 173
rect 3817 173 3833 183
rect 4100 183 4113 187
rect 4097 173 4113 183
rect 4660 183 4673 187
rect 4657 173 4673 183
rect 3817 143 3823 173
rect 4097 147 4103 173
rect 2617 137 2643 143
rect 3817 140 3843 143
rect 3817 137 3847 140
rect 467 117 613 123
rect 1077 123 1083 137
rect 1027 117 1083 123
rect 2177 123 2183 137
rect 2637 127 2643 137
rect 3833 127 3847 137
rect 4087 137 4103 147
rect 4657 143 4663 173
rect 4637 137 4663 143
rect 4087 133 4100 137
rect 2127 117 2183 123
rect 2547 117 2613 123
rect 2637 125 2660 127
rect 2637 117 2653 125
rect 2640 113 2653 117
rect 3487 117 3513 123
rect 4167 117 4233 123
rect 4637 123 4643 137
rect 4607 117 4643 123
rect 5007 117 5113 123
rect 5507 117 5573 123
rect 687 97 713 103
rect 2547 97 2613 103
rect -63 2 30 18
rect 5843 2 5903 262
<< m2contact >>
rect 3153 5413 3167 5427
rect 3173 5413 3187 5427
rect 1453 5393 1467 5407
rect 1493 5393 1507 5407
rect 2713 5393 2727 5407
rect 2813 5393 2827 5407
rect 3313 5373 3327 5387
rect 3253 5313 3267 5327
rect 5333 5313 5347 5327
rect 5413 5313 5427 5327
rect 1693 5273 1707 5287
rect 1773 5272 1787 5286
rect 1653 5093 1667 5107
rect 4753 5093 4767 5107
rect 4833 5093 4847 5107
rect 73 5073 87 5087
rect 73 5033 87 5047
rect 1913 5073 1927 5087
rect 1893 5033 1907 5047
rect 1933 5033 1947 5047
rect 1693 5013 1707 5027
rect 1113 4893 1127 4907
rect 3093 4893 3107 4907
rect 3133 4893 3147 4907
rect 5713 4892 5727 4906
rect 5773 4893 5787 4907
rect 1173 4873 1187 4887
rect 2913 4874 2927 4888
rect 1113 4852 1127 4866
rect 1153 4853 1167 4867
rect 1273 4853 1287 4867
rect 1413 4853 1427 4867
rect 1273 4813 1287 4827
rect 113 4793 127 4807
rect 193 4793 207 4807
rect 1333 4793 1347 4807
rect 2933 4813 2947 4827
rect 3113 4853 3127 4867
rect 3233 4853 3247 4867
rect 3613 4853 3627 4867
rect 5713 4853 5727 4867
rect 3113 4813 3127 4827
rect 3573 4813 3587 4827
rect 5713 4813 5727 4827
rect 3253 4793 3267 4807
rect 4433 4593 4447 4607
rect 4513 4593 4527 4607
rect 1613 4573 1627 4587
rect 1733 4573 1747 4587
rect 1793 4573 1807 4587
rect 2353 4573 2367 4587
rect 2413 4573 2427 4587
rect 2573 4573 2587 4587
rect 2673 4574 2687 4588
rect 1493 4553 1507 4567
rect 1713 4553 1727 4567
rect 1533 4513 1547 4527
rect 1653 4513 1667 4527
rect 3193 4552 3207 4566
rect 3473 4553 3487 4567
rect 3933 4553 3947 4567
rect 4233 4553 4247 4567
rect 4273 4553 4287 4567
rect 4453 4553 4467 4567
rect 4553 4573 4567 4587
rect 1733 4512 1747 4526
rect 3193 4513 3207 4527
rect 3413 4513 3427 4527
rect 3973 4513 3987 4527
rect 4433 4493 4447 4507
rect 4893 4553 4907 4567
rect 5633 4553 5647 4567
rect 4513 4513 4527 4527
rect 4893 4513 4907 4527
rect 5593 4513 5607 4527
rect 2373 4472 2387 4486
rect 2393 4473 2407 4487
rect 3913 4473 3927 4487
rect 3993 4473 4007 4487
rect 5013 4473 5027 4487
rect 5073 4473 5087 4487
rect 5693 4373 5707 4387
rect 953 4353 967 4367
rect 1013 4353 1027 4367
rect 233 4333 247 4347
rect 613 4333 627 4347
rect 4033 4333 4047 4347
rect 4993 4333 5007 4347
rect 5173 4333 5187 4347
rect 273 4293 287 4307
rect 653 4293 667 4307
rect 3993 4293 4007 4307
rect 1313 4273 1327 4287
rect 1373 4273 1387 4287
rect 1813 4273 1827 4287
rect 1913 4273 1927 4287
rect 3113 4273 3127 4287
rect 3153 4273 3167 4287
rect 4913 4273 4927 4287
rect 5213 4293 5227 4307
rect 5153 4271 5167 4285
rect 5193 4273 5207 4287
rect 3973 4253 3987 4267
rect 4053 4252 4067 4266
rect 5733 4232 5747 4246
rect 493 4053 507 4067
rect 553 4053 567 4067
rect 2493 4053 2507 4067
rect 2613 4053 2627 4067
rect 3293 4053 3307 4067
rect 3353 4053 3367 4067
rect 3413 4053 3427 4067
rect 3473 4052 3487 4066
rect 3913 4053 3927 4067
rect 3993 4053 4007 4067
rect 5073 4053 5087 4067
rect 5113 4053 5127 4067
rect 5193 4053 5207 4067
rect 5233 4053 5247 4067
rect 5753 4053 5767 4067
rect 333 4033 347 4047
rect 393 4033 407 4047
rect 293 3993 307 4007
rect 3073 4033 3087 4047
rect 3933 4033 3947 4047
rect 5353 4033 5367 4047
rect 3073 3993 3087 4007
rect 3933 3993 3947 4007
rect 5353 3993 5367 4007
rect 5733 3993 5747 4007
rect 453 3973 467 3987
rect 3913 3953 3927 3967
rect 3973 3953 3987 3967
rect 1553 3833 1567 3847
rect 1633 3833 1647 3847
rect 2273 3833 2287 3847
rect 2333 3833 2347 3847
rect 5413 3833 5427 3847
rect 533 3813 547 3827
rect 533 3773 547 3787
rect 713 3813 727 3827
rect 813 3813 827 3827
rect 1313 3813 1327 3827
rect 1353 3813 1367 3827
rect 1453 3813 1467 3827
rect 1853 3813 1867 3827
rect 713 3773 727 3787
rect 853 3773 867 3787
rect 1453 3773 1467 3787
rect 2053 3813 2067 3827
rect 3893 3813 3907 3827
rect 1893 3773 1907 3787
rect 4613 3793 4627 3807
rect 5773 3813 5787 3827
rect 3893 3773 3907 3787
rect 4633 3773 4647 3787
rect 5373 3773 5387 3787
rect 5773 3773 5787 3787
rect 633 3753 647 3767
rect 753 3753 767 3767
rect 2013 3753 2027 3767
rect 5633 3553 5647 3567
rect 5713 3553 5727 3567
rect 1573 3533 1587 3547
rect 5093 3533 5107 3547
rect 5673 3533 5687 3547
rect 5453 3513 5467 3527
rect 1593 3473 1607 3487
rect 2053 3473 2067 3487
rect 2093 3473 2107 3487
rect 5133 3473 5147 3487
rect 5393 3473 5407 3487
rect 5773 3513 5787 3527
rect 5813 3513 5827 3527
rect 5693 3473 5707 3487
rect 3973 3453 3987 3467
rect 4033 3453 4047 3467
rect 1233 3353 1247 3367
rect 1273 3353 1287 3367
rect 1053 3333 1067 3347
rect 1133 3333 1147 3347
rect 633 3313 647 3327
rect 673 3313 687 3327
rect 153 3293 167 3307
rect 193 3293 207 3307
rect 993 3293 1007 3307
rect 4773 3313 4787 3327
rect 4693 3253 4707 3267
rect 4873 3293 4887 3307
rect 273 3233 287 3247
rect 313 3233 327 3247
rect 953 3233 967 3247
rect 3233 3233 3247 3247
rect 3313 3233 3327 3247
rect 4833 3233 4847 3247
rect 5333 3233 5347 3247
rect 5453 3233 5467 3247
rect 3393 3012 3407 3026
rect 3513 3013 3527 3027
rect 1273 2993 1287 3007
rect 1273 2953 1287 2967
rect 5333 2933 5347 2947
rect 5393 2933 5407 2947
rect 5453 2933 5467 2947
rect 4913 2833 4927 2847
rect 4973 2813 4987 2827
rect 2173 2793 2187 2807
rect 2593 2793 2607 2807
rect 2633 2793 2647 2807
rect 1433 2773 1447 2787
rect 1633 2773 1647 2787
rect 1373 2733 1387 2747
rect 1673 2733 1687 2747
rect 2133 2733 2147 2747
rect 5773 2733 5787 2747
rect 5813 2733 5827 2747
rect 4073 2713 4087 2727
rect 4113 2713 4127 2727
rect 2853 2513 2867 2527
rect 2913 2513 2927 2527
rect 5093 2493 5107 2507
rect 3573 2473 3587 2487
rect 4573 2473 4587 2487
rect 3513 2433 3527 2447
rect 4733 2473 4747 2487
rect 4813 2473 4827 2487
rect 4953 2473 4967 2487
rect 5753 2493 5767 2507
rect 4573 2433 4587 2447
rect 4693 2433 4707 2447
rect 4853 2433 4867 2447
rect 5553 2453 5567 2467
rect 5013 2433 5027 2447
rect 5133 2433 5147 2447
rect 5233 2433 5247 2447
rect 5293 2433 5307 2447
rect 5533 2433 5547 2447
rect 5773 2433 5787 2447
rect 4593 2293 4607 2307
rect 1213 2274 1227 2288
rect 1313 2273 1327 2287
rect 3893 2273 3907 2287
rect 3953 2273 3967 2287
rect 4433 2273 4447 2287
rect 4473 2273 4487 2287
rect 4533 2273 4547 2287
rect 2073 2253 2087 2267
rect 3573 2253 3587 2267
rect 3833 2253 3847 2267
rect 4233 2253 4247 2267
rect 4333 2253 4347 2267
rect 4453 2253 4467 2267
rect 5453 2273 5467 2287
rect 5513 2272 5527 2286
rect 2333 2233 2347 2247
rect 2353 2213 2367 2227
rect 3573 2213 3587 2227
rect 3793 2213 3807 2227
rect 4873 2253 4887 2267
rect 5013 2253 5027 2267
rect 4233 2213 4247 2227
rect 4373 2213 4387 2227
rect 4513 2213 4527 2227
rect 4593 2213 4607 2227
rect 4913 2213 4927 2227
rect 5013 2213 5027 2227
rect 5213 2253 5227 2267
rect 5433 2253 5447 2267
rect 5213 2213 5227 2227
rect 5613 2233 5627 2247
rect 2013 2193 2027 2207
rect 3393 2193 3407 2207
rect 3473 2193 3487 2207
rect 3633 2193 3647 2207
rect 3773 2191 3787 2205
rect 3853 2193 3867 2207
rect 4433 2193 4447 2207
rect 4473 2193 4487 2207
rect 5573 2213 5587 2227
rect 5533 2191 5547 2205
rect 5693 2193 5707 2207
rect 3733 2173 3747 2187
rect 4573 2152 4587 2166
rect 4633 2153 4647 2167
rect 5693 2153 5707 2167
rect 4593 2013 4607 2027
rect 4633 2013 4647 2027
rect 173 1973 187 1987
rect 253 1973 267 1987
rect 1433 1973 1447 1987
rect 693 1953 707 1967
rect 1073 1953 1087 1967
rect 1333 1953 1347 1967
rect 1573 1973 1587 1987
rect 1613 1973 1627 1987
rect 1873 1973 1887 1987
rect 1933 1973 1947 1987
rect 3033 1973 3047 1987
rect 3093 1973 3107 1987
rect 653 1913 667 1927
rect 1113 1913 1127 1927
rect 1373 1913 1387 1927
rect 1473 1913 1487 1927
rect 1633 1953 1647 1967
rect 1753 1953 1767 1967
rect 1633 1913 1647 1927
rect 1893 1953 1907 1967
rect 2433 1953 2447 1967
rect 2973 1953 2987 1967
rect 1893 1913 1907 1927
rect 2393 1913 2407 1927
rect 2913 1913 2927 1927
rect 1813 1891 1827 1905
rect 3633 1973 3647 1987
rect 4593 1973 4607 1987
rect 4693 1973 4707 1987
rect 5313 1973 5327 1987
rect 5393 1973 5407 1987
rect 5753 1973 5767 1987
rect 5813 1973 5827 1987
rect 3613 1953 3627 1967
rect 3713 1953 3727 1967
rect 3713 1913 3727 1927
rect 3893 1953 3907 1967
rect 4153 1953 4167 1967
rect 4273 1953 4287 1967
rect 4513 1953 4527 1967
rect 4753 1953 4767 1967
rect 5013 1953 5027 1967
rect 5293 1953 5307 1967
rect 4233 1913 4247 1927
rect 4533 1913 4547 1927
rect 4793 1913 4807 1927
rect 5053 1913 5067 1927
rect 5293 1913 5307 1927
rect 4173 1893 4187 1907
rect 3593 1873 3607 1887
rect 3893 1873 3907 1887
rect 4933 1873 4947 1887
rect 4973 1873 4987 1887
rect 3573 1853 3587 1867
rect 2853 1753 2867 1767
rect 2013 1733 2027 1747
rect 2313 1733 2327 1747
rect 2433 1733 2447 1747
rect 2013 1693 2027 1707
rect 273 1673 287 1687
rect 413 1673 427 1687
rect 2153 1673 2167 1687
rect 2253 1671 2267 1685
rect 2293 1671 2307 1685
rect 2433 1693 2447 1707
rect 2573 1733 2587 1747
rect 2813 1733 2827 1747
rect 2573 1693 2587 1707
rect 2793 1673 2807 1687
rect 4273 1752 4287 1766
rect 3233 1733 3247 1747
rect 3333 1733 3347 1747
rect 3793 1733 3807 1747
rect 3933 1732 3947 1746
rect 4033 1733 4047 1747
rect 4133 1733 4147 1747
rect 4313 1733 4327 1747
rect 4413 1733 4427 1747
rect 3233 1693 3247 1707
rect 3333 1693 3347 1707
rect 3753 1693 3767 1707
rect 3893 1693 3907 1707
rect 4073 1693 4087 1707
rect 4133 1693 4147 1707
rect 4573 1733 4587 1747
rect 4813 1733 4827 1747
rect 4913 1733 4927 1747
rect 4573 1693 4587 1707
rect 2873 1673 2887 1687
rect 3133 1671 3147 1685
rect 3173 1673 3187 1687
rect 3853 1673 3867 1687
rect 3933 1673 3947 1687
rect 4473 1673 4487 1687
rect 4753 1673 4767 1687
rect 5113 1733 5127 1747
rect 5233 1733 5247 1747
rect 5653 1733 5667 1747
rect 4973 1693 4987 1707
rect 5073 1693 5087 1707
rect 5233 1693 5247 1707
rect 5653 1693 5667 1707
rect 4113 1653 4127 1667
rect 4213 1653 4227 1667
rect 5313 1633 5327 1647
rect 5373 1633 5387 1647
rect 3853 1533 3867 1547
rect 3893 1533 3907 1547
rect 4333 1473 4347 1487
rect 4413 1473 4427 1487
rect 5693 1473 5707 1487
rect 5773 1473 5787 1487
rect 113 1453 127 1467
rect 193 1453 207 1467
rect 2253 1453 2267 1467
rect 2313 1453 2327 1467
rect 2653 1453 2667 1467
rect 2733 1453 2747 1467
rect 4073 1453 4087 1467
rect 1353 1433 1367 1447
rect 1573 1433 1587 1447
rect 2113 1433 2127 1447
rect 2573 1433 2587 1447
rect 2833 1433 2847 1447
rect 4533 1453 4547 1467
rect 1353 1393 1367 1407
rect 1613 1393 1627 1407
rect 2153 1393 2167 1407
rect 2573 1393 2587 1407
rect 2793 1393 2807 1407
rect 4473 1433 4487 1447
rect 4133 1393 4147 1407
rect 4473 1393 4487 1407
rect 5093 1433 5107 1447
rect 5553 1433 5567 1447
rect 5093 1393 5107 1407
rect 5513 1393 5527 1407
rect 5753 1453 5767 1467
rect 5713 1393 5727 1407
rect 5193 1373 5207 1387
rect 5233 1373 5247 1387
rect 5393 1373 5407 1387
rect 5453 1371 5467 1385
rect 4253 1353 4267 1367
rect 4193 1333 4207 1347
rect 153 1233 167 1247
rect 233 1233 247 1247
rect 833 1233 847 1247
rect 873 1233 887 1247
rect 1313 1233 1327 1247
rect 1393 1233 1407 1247
rect 1473 1232 1487 1246
rect 1533 1233 1547 1247
rect 2273 1233 2287 1247
rect 2153 1213 2167 1227
rect 2233 1173 2247 1187
rect 3733 1193 3747 1207
rect 4053 1234 4067 1248
rect 4753 1234 4767 1248
rect 4793 1233 4807 1247
rect 5053 1233 5067 1247
rect 3753 1173 3767 1187
rect 4013 1173 4027 1187
rect 4293 1213 4307 1227
rect 4673 1213 4687 1227
rect 4893 1213 4907 1227
rect 4673 1173 4687 1187
rect 5433 1213 5447 1227
rect 5493 1193 5507 1207
rect 4953 1173 4967 1187
rect 5073 1173 5087 1187
rect 793 1153 807 1167
rect 873 1153 887 1167
rect 1493 1153 1507 1167
rect 1573 1153 1587 1167
rect 1613 1153 1627 1167
rect 1673 1153 1687 1167
rect 2093 1153 2107 1167
rect 2173 1153 2187 1167
rect 2353 1153 2367 1167
rect 2413 1153 2427 1167
rect 3513 1153 3527 1167
rect 3573 1153 3587 1167
rect 3833 1153 3847 1167
rect 3913 1153 3927 1167
rect 4233 1153 4247 1167
rect 393 1133 407 1147
rect 433 1132 447 1146
rect 3233 1133 3247 1147
rect 3313 1133 3327 1147
rect 973 973 987 987
rect 1033 973 1047 987
rect 1173 973 1187 987
rect 1213 973 1227 987
rect 2393 973 2407 987
rect 553 953 567 967
rect 593 953 607 967
rect 1513 953 1527 967
rect 1613 953 1627 967
rect 2473 953 2487 967
rect 93 933 107 947
rect 213 933 227 947
rect 1093 934 1107 948
rect 1173 933 1187 947
rect 1533 933 1547 947
rect 1613 932 1627 946
rect 3533 933 3547 947
rect 3573 933 3587 947
rect 333 913 347 927
rect 2293 913 2307 927
rect 2413 913 2427 927
rect 173 893 187 907
rect 193 873 207 887
rect 293 873 307 887
rect 113 853 127 867
rect 173 853 187 867
rect 2273 853 2287 867
rect 2433 872 2447 886
rect 2713 913 2727 927
rect 3093 913 3107 927
rect 3353 913 3367 927
rect 3653 932 3667 946
rect 4253 933 4267 947
rect 4373 933 4387 947
rect 4673 933 4687 947
rect 5433 933 5447 947
rect 5493 933 5507 947
rect 5533 933 5547 947
rect 3053 873 3067 887
rect 3393 873 3407 887
rect 2673 852 2687 866
rect 3453 853 3467 867
rect 5673 932 5687 946
rect 5073 913 5087 927
rect 4673 892 4687 906
rect 5253 913 5267 927
rect 5373 913 5387 927
rect 5113 873 5127 887
rect 5253 873 5267 887
rect 5333 873 5347 887
rect 113 733 127 747
rect 133 713 147 727
rect 193 713 207 727
rect 673 713 687 727
rect 393 693 407 707
rect 713 713 727 727
rect 153 653 167 667
rect 813 693 827 707
rect 353 633 367 647
rect 673 653 687 667
rect 813 653 827 667
rect 1413 693 1427 707
rect 1513 693 1527 707
rect 473 633 487 647
rect 553 633 567 647
rect 1333 633 1347 647
rect 1693 693 1707 707
rect 1853 693 1867 707
rect 1993 693 2007 707
rect 2133 693 2147 707
rect 1513 653 1527 667
rect 1653 653 1667 667
rect 1793 653 1807 667
rect 1953 653 1967 667
rect 2313 714 2327 728
rect 2493 693 2507 707
rect 2773 693 2787 707
rect 2913 693 2927 707
rect 3053 693 3067 707
rect 2133 653 2147 667
rect 2293 653 2307 667
rect 2533 653 2547 667
rect 2813 653 2827 667
rect 1753 633 1767 647
rect 1833 633 1847 647
rect 2073 633 2087 647
rect 2153 633 2167 647
rect 2213 633 2227 647
rect 2273 633 2287 647
rect 2473 633 2487 647
rect 2593 633 2607 647
rect 3053 653 3067 667
rect 3113 693 3127 707
rect 3213 693 3227 707
rect 3393 693 3407 707
rect 3453 693 3467 707
rect 4453 693 4467 707
rect 5153 693 5167 707
rect 5433 693 5447 707
rect 5533 693 5547 707
rect 3113 653 3127 667
rect 3213 653 3227 667
rect 3353 653 3367 667
rect 3453 653 3467 667
rect 4413 653 4427 667
rect 5153 653 5167 667
rect 3013 631 3027 645
rect 3953 633 3967 647
rect 3993 633 4007 647
rect 4093 633 4107 647
rect 4153 633 4167 647
rect 4213 633 4227 647
rect 4353 633 4367 647
rect 4473 633 4487 647
rect 5333 633 5347 647
rect 5533 653 5547 667
rect 253 413 267 427
rect 353 413 367 427
rect 833 413 847 427
rect 893 413 907 427
rect 1173 413 1187 427
rect 1213 413 1227 427
rect 213 393 227 407
rect 1533 413 1547 427
rect 1673 413 1687 427
rect 2113 413 2127 427
rect 2233 413 2247 427
rect 2793 413 2807 427
rect 1833 393 1847 407
rect 213 353 227 367
rect 1453 353 1467 367
rect 1593 353 1607 367
rect 1833 353 1847 367
rect 2313 393 2327 407
rect 2693 393 2707 407
rect 3073 413 3087 427
rect 2973 393 2987 407
rect 4553 413 4567 427
rect 4673 413 4687 427
rect 5133 413 5147 427
rect 5433 413 5447 427
rect 2313 353 2327 367
rect 2693 353 2707 367
rect 2833 353 2847 367
rect 2973 353 2987 367
rect 3093 333 3107 347
rect 5133 353 5147 367
rect 3393 333 3407 347
rect 3453 331 3467 345
rect 5373 333 5387 347
rect 3133 313 3147 327
rect 3153 312 3167 326
rect 2313 233 2327 247
rect 2353 233 2367 247
rect 1313 213 1327 227
rect 1373 213 1387 227
rect 5313 213 5327 227
rect 5353 213 5367 227
rect 1113 173 1127 187
rect 2213 173 2227 187
rect 2693 193 2707 207
rect 5053 193 5067 207
rect 5133 193 5147 207
rect 2733 173 2747 187
rect 2753 152 2767 166
rect 3833 173 3847 187
rect 4113 173 4127 187
rect 4673 173 4687 187
rect 453 113 467 127
rect 613 113 627 127
rect 1013 113 1027 127
rect 2113 113 2127 127
rect 4073 133 4087 147
rect 2533 113 2547 127
rect 2613 113 2627 127
rect 2653 111 2667 125
rect 3473 113 3487 127
rect 3513 113 3527 127
rect 3833 113 3847 127
rect 4153 113 4167 127
rect 4233 113 4247 127
rect 4593 113 4607 127
rect 4993 111 5007 125
rect 5113 113 5127 127
rect 5493 113 5507 127
rect 5573 113 5587 127
rect 673 93 687 107
rect 713 93 727 107
rect 2533 92 2547 106
rect 2613 92 2627 106
<< metal2 >>
rect 653 5380 667 5393
rect 656 5376 663 5380
rect 36 5247 43 5343
rect 96 5336 123 5343
rect 116 5187 123 5336
rect 76 5087 83 5173
rect 276 5147 283 5353
rect 616 5347 623 5374
rect 316 5340 323 5343
rect 313 5327 327 5340
rect 353 5323 367 5333
rect 336 5320 367 5323
rect 336 5316 363 5320
rect 56 4867 63 5074
rect 276 5076 283 5133
rect 73 5027 87 5033
rect 96 4947 103 5043
rect 196 5007 203 5074
rect 216 4947 223 5033
rect 256 5007 263 5043
rect 316 4907 323 5073
rect 336 5047 343 5316
rect 556 5247 563 5343
rect 676 5327 683 5343
rect 676 5287 683 5313
rect 756 5287 763 5393
rect 1036 5347 1043 5523
rect 2096 5487 2103 5523
rect 2216 5487 2223 5523
rect 2836 5487 2843 5523
rect 1376 5347 1383 5413
rect 1453 5407 1467 5413
rect 1507 5396 1563 5403
rect 1556 5376 1563 5396
rect 796 5287 803 5343
rect 553 5080 567 5093
rect 556 5076 563 5080
rect 596 5076 603 5233
rect 456 5043 463 5074
rect 416 4987 423 5043
rect 456 5036 483 5043
rect 236 4856 243 4893
rect 56 4387 63 4813
rect 76 4567 83 4823
rect 116 4820 123 4823
rect 113 4807 127 4820
rect 156 4787 163 4853
rect 276 4826 283 4893
rect 476 4856 483 5036
rect 496 4947 503 5043
rect 696 5007 703 5233
rect 573 4860 587 4873
rect 576 4856 583 4860
rect 416 4826 423 4853
rect 216 4807 223 4823
rect 207 4796 223 4807
rect 207 4793 220 4796
rect 376 4607 383 4823
rect 496 4787 503 4823
rect 656 4727 663 4973
rect 716 4967 723 5273
rect 816 5027 823 5093
rect 716 4856 723 4913
rect 756 4887 763 4953
rect 753 4860 767 4873
rect 756 4856 763 4860
rect 696 4787 703 4823
rect 796 4767 803 4993
rect 836 4887 843 5343
rect 956 5340 963 5343
rect 953 5327 967 5340
rect 1136 5340 1143 5343
rect 956 5247 963 5313
rect 976 5087 983 5133
rect 916 5076 963 5083
rect 896 5040 903 5043
rect 893 5027 907 5040
rect 936 4987 943 5033
rect 856 4856 863 4973
rect 956 4947 963 5076
rect 996 5076 1003 5113
rect 1036 5076 1043 5213
rect 1076 5187 1083 5332
rect 1133 5327 1147 5340
rect 1136 5267 1143 5313
rect 1476 5287 1483 5374
rect 1616 5346 1623 5373
rect 1476 5247 1483 5273
rect 1656 5247 1663 5343
rect 1696 5287 1703 5343
rect 1736 5307 1743 5353
rect 1856 5346 1863 5413
rect 1776 5307 1783 5343
rect 1836 5287 1843 5313
rect 1780 5286 1800 5287
rect 1787 5273 1793 5286
rect 1296 5207 1303 5233
rect 1056 5040 1063 5043
rect 1053 5027 1067 5040
rect 976 4923 983 4953
rect 956 4916 983 4923
rect 893 4860 907 4873
rect 896 4856 903 4860
rect 116 4556 123 4593
rect 436 4556 443 4593
rect 696 4556 703 4653
rect 796 4643 803 4753
rect 776 4636 803 4643
rect 736 4568 743 4633
rect 776 4556 783 4636
rect 156 4526 163 4553
rect 276 4527 283 4554
rect 196 4487 203 4523
rect 276 4447 283 4513
rect 396 4487 403 4554
rect 516 4527 523 4554
rect 220 4343 233 4347
rect 216 4336 233 4343
rect 220 4333 233 4336
rect 316 4336 323 4373
rect 256 4306 263 4333
rect 116 4127 123 4303
rect 276 4048 283 4293
rect 336 4283 343 4303
rect 316 4276 343 4283
rect 76 4036 103 4043
rect 76 3983 83 4036
rect 196 4006 203 4033
rect 76 3976 103 3983
rect 96 3816 103 3976
rect 136 3967 143 4003
rect 256 3987 263 4003
rect 236 3816 243 3893
rect 256 3867 263 3973
rect 296 3907 303 3993
rect 316 3987 323 4276
rect 356 4183 363 4293
rect 336 4176 363 4183
rect 336 4047 343 4176
rect 376 4167 383 4433
rect 396 4407 403 4473
rect 556 4427 563 4523
rect 596 4520 603 4523
rect 593 4507 607 4520
rect 656 4467 663 4554
rect 473 4343 487 4353
rect 456 4340 487 4343
rect 456 4336 483 4340
rect 376 4047 383 4113
rect 376 4036 393 4047
rect 380 4033 393 4036
rect 156 3787 163 3814
rect 76 3707 83 3783
rect 296 3786 303 3853
rect 316 3847 323 3952
rect 56 3696 73 3703
rect 16 2787 23 3613
rect 56 3527 63 3696
rect 116 3527 123 3772
rect 96 3516 113 3523
rect 56 3307 63 3473
rect 76 3467 83 3483
rect 136 3480 143 3483
rect 133 3467 147 3480
rect 76 3327 83 3453
rect 96 3296 103 3353
rect 156 3266 163 3293
rect 76 3260 83 3263
rect 36 2807 43 3013
rect 56 2867 63 3253
rect 73 3247 87 3260
rect 116 3027 123 3263
rect 136 3007 143 3193
rect 176 3083 183 3393
rect 196 3367 203 3733
rect 216 3707 223 3783
rect 316 3747 323 3833
rect 356 3816 363 3893
rect 396 3827 403 3873
rect 376 3747 383 3783
rect 396 3667 403 3773
rect 416 3543 423 4153
rect 476 4036 483 4073
rect 496 4067 503 4393
rect 556 4336 563 4373
rect 616 4347 623 4373
rect 576 4207 583 4303
rect 456 4000 463 4003
rect 436 3827 443 3993
rect 453 3987 467 4000
rect 496 3927 503 4003
rect 453 3820 467 3833
rect 456 3816 463 3820
rect 496 3816 503 3873
rect 536 3827 543 3873
rect 436 3567 443 3773
rect 520 3783 533 3787
rect 516 3776 533 3783
rect 520 3773 533 3776
rect 536 3627 543 3693
rect 416 3536 443 3543
rect 313 3520 327 3533
rect 316 3516 323 3520
rect 216 3323 223 3513
rect 196 3320 223 3323
rect 193 3316 223 3320
rect 193 3307 207 3316
rect 256 3296 263 3453
rect 356 3407 363 3533
rect 436 3528 443 3536
rect 460 3486 480 3487
rect 467 3483 480 3486
rect 467 3476 483 3483
rect 467 3473 480 3476
rect 536 3403 543 3553
rect 516 3396 543 3403
rect 476 3308 483 3373
rect 516 3296 523 3396
rect 556 3303 563 4053
rect 636 4036 643 4353
rect 693 4340 707 4353
rect 716 4347 723 4523
rect 756 4423 763 4513
rect 896 4443 903 4713
rect 956 4647 963 4916
rect 996 4903 1003 5013
rect 1116 5007 1123 5173
rect 1136 5088 1143 5133
rect 1176 5076 1183 5113
rect 1216 5076 1223 5173
rect 1256 5076 1263 5133
rect 1296 5076 1303 5193
rect 1136 5027 1143 5074
rect 1196 4967 1203 5043
rect 976 4896 1003 4903
rect 976 4823 983 4896
rect 1113 4887 1127 4893
rect 976 4816 1003 4823
rect 1016 4820 1023 4823
rect 996 4607 1003 4816
rect 1013 4807 1027 4820
rect 1076 4767 1083 4823
rect 1116 4787 1123 4852
rect 996 4526 1003 4593
rect 1016 4568 1023 4653
rect 1096 4556 1103 4593
rect 896 4436 923 4443
rect 736 4416 763 4423
rect 696 4336 703 4340
rect 736 4336 743 4416
rect 916 4367 923 4436
rect 956 4367 963 4413
rect 1016 4367 1023 4554
rect 1076 4467 1083 4523
rect 1136 4507 1143 4913
rect 1156 4867 1163 4893
rect 1173 4860 1187 4873
rect 1216 4868 1223 5013
rect 1236 4987 1243 5043
rect 1176 4856 1183 4860
rect 1276 4867 1283 4993
rect 1256 4727 1263 4854
rect 1296 4856 1303 4893
rect 1336 4856 1343 4893
rect 1276 4623 1283 4813
rect 1276 4616 1303 4623
rect 1233 4560 1247 4573
rect 1236 4556 1243 4560
rect 1196 4467 1203 4523
rect 656 4267 663 4293
rect 576 3827 583 3913
rect 616 3887 623 4003
rect 656 3983 663 4193
rect 676 4103 683 4303
rect 836 4296 863 4303
rect 836 4267 843 4296
rect 916 4127 923 4303
rect 956 4267 963 4353
rect 976 4306 983 4353
rect 1093 4340 1107 4353
rect 1096 4336 1103 4340
rect 1056 4267 1063 4303
rect 676 4096 703 4103
rect 636 3976 663 3983
rect 636 3863 643 3976
rect 616 3856 643 3863
rect 616 3816 623 3856
rect 656 3816 663 3913
rect 676 3827 683 4073
rect 696 3927 703 4096
rect 756 4000 763 4003
rect 753 3987 767 4000
rect 816 3987 823 4034
rect 636 3767 643 3783
rect 696 3767 703 3873
rect 716 3827 723 3853
rect 736 3816 743 3913
rect 776 3816 783 3853
rect 816 3827 823 3973
rect 876 3887 883 4003
rect 936 4000 943 4003
rect 933 3987 947 4000
rect 996 3867 1003 4253
rect 1116 4036 1123 4113
rect 1016 3967 1023 4013
rect 836 3786 843 3853
rect 1036 3843 1043 3993
rect 1016 3836 1043 3843
rect 1016 3816 1023 3836
rect 1056 3816 1063 3853
rect 1156 3847 1163 4453
rect 1276 4447 1283 4573
rect 1176 4307 1183 4373
rect 1296 4367 1303 4616
rect 1336 4556 1343 4793
rect 1356 4727 1363 4823
rect 1396 4767 1403 5113
rect 1416 5046 1423 5133
rect 1516 5047 1523 5074
rect 1536 5043 1543 5113
rect 1616 5076 1623 5113
rect 1653 5088 1667 5093
rect 1666 5080 1667 5088
rect 1756 5076 1763 5133
rect 1536 5036 1563 5043
rect 1416 4947 1423 4993
rect 1416 4867 1423 4933
rect 1436 4868 1443 4953
rect 1456 4820 1463 4823
rect 1453 4807 1467 4820
rect 1276 4127 1283 4303
rect 1296 4267 1303 4293
rect 1316 4287 1323 4333
rect 1236 4036 1243 4073
rect 1336 4063 1343 4493
rect 1376 4447 1383 4523
rect 1396 4407 1403 4713
rect 1476 4687 1483 4813
rect 1416 4526 1423 4573
rect 1496 4567 1503 4893
rect 1556 4856 1563 5036
rect 1656 4967 1663 5013
rect 1676 5007 1683 5074
rect 1693 5027 1707 5033
rect 1676 4947 1683 4993
rect 1596 4856 1603 4893
rect 1676 4856 1683 4893
rect 1516 4816 1543 4823
rect 1576 4820 1583 4823
rect 1696 4820 1703 4823
rect 1516 4727 1523 4816
rect 1573 4807 1587 4820
rect 1693 4807 1707 4820
rect 1747 4816 1763 4823
rect 1516 4467 1523 4713
rect 1613 4567 1627 4573
rect 1536 4487 1543 4513
rect 1600 4523 1613 4527
rect 1596 4516 1613 4523
rect 1600 4513 1613 4516
rect 1396 4336 1403 4372
rect 1376 4300 1383 4303
rect 1373 4287 1387 4300
rect 1416 4227 1423 4303
rect 1476 4267 1483 4453
rect 1376 4067 1383 4213
rect 1496 4167 1503 4353
rect 1556 4343 1563 4433
rect 1556 4336 1583 4343
rect 1336 4056 1363 4063
rect 1216 3967 1223 4003
rect 1276 3967 1283 4003
rect 1336 3927 1343 4033
rect 756 3780 763 3783
rect 796 3780 803 3783
rect 633 3747 647 3753
rect 576 3543 583 3593
rect 576 3536 603 3543
rect 596 3516 603 3536
rect 653 3520 667 3533
rect 656 3516 663 3520
rect 696 3486 703 3593
rect 716 3587 723 3773
rect 753 3767 767 3780
rect 793 3767 807 3780
rect 956 3786 963 3813
rect 1196 3786 1203 3813
rect 856 3747 863 3773
rect 896 3516 903 3753
rect 916 3747 923 3783
rect 1036 3707 1043 3783
rect 936 3516 943 3553
rect 756 3447 763 3483
rect 596 3307 603 3353
rect 556 3296 583 3303
rect 276 3260 283 3263
rect 273 3247 287 3260
rect 316 3247 323 3293
rect 356 3207 363 3252
rect 396 3167 403 3263
rect 436 3127 443 3294
rect 156 3076 183 3083
rect 156 3027 163 3076
rect 156 2996 163 3013
rect 16 1907 23 2733
rect 36 2687 43 2743
rect 96 2740 103 2743
rect 93 2727 107 2740
rect 136 2507 143 2853
rect 156 2587 163 2793
rect 216 2776 223 2873
rect 276 2687 283 3013
rect 336 2803 343 2952
rect 376 2903 383 3113
rect 576 3067 583 3296
rect 633 3300 647 3313
rect 673 3308 687 3313
rect 636 3296 643 3300
rect 716 3296 723 3373
rect 396 2927 403 2993
rect 376 2896 403 2903
rect 316 2796 343 2803
rect 316 2776 323 2796
rect 396 2747 403 2896
rect 496 2807 503 3053
rect 676 3047 683 3294
rect 736 3260 743 3263
rect 733 3247 747 3260
rect 796 3207 803 3433
rect 856 3387 863 3514
rect 916 3447 923 3483
rect 876 3336 883 3393
rect 816 3296 843 3303
rect 816 3247 823 3296
rect 956 3263 963 3353
rect 976 3267 983 3333
rect 996 3307 1003 3573
rect 1016 3527 1023 3593
rect 1036 3516 1043 3653
rect 1076 3516 1083 3573
rect 1096 3547 1103 3783
rect 1216 3687 1223 3913
rect 1276 3816 1283 3853
rect 1296 3827 1303 3873
rect 1356 3827 1363 4056
rect 1456 4036 1463 4113
rect 1056 3447 1063 3483
rect 1136 3483 1143 3573
rect 1216 3516 1223 3593
rect 1116 3476 1143 3483
rect 1196 3480 1203 3483
rect 1056 3347 1063 3433
rect 1007 3296 1023 3303
rect 936 3256 963 3263
rect 576 2996 583 3032
rect 636 2967 643 2994
rect 556 2823 563 2963
rect 716 2927 723 2963
rect 776 2927 783 2994
rect 796 2963 803 3093
rect 856 3008 863 3193
rect 867 2996 883 3003
rect 876 2967 883 2996
rect 796 2956 823 2963
rect 556 2816 583 2823
rect 487 2783 500 2787
rect 487 2776 503 2783
rect 487 2773 500 2776
rect 73 2488 87 2493
rect 196 2446 203 2573
rect 276 2567 283 2673
rect 316 2476 323 2553
rect 376 2476 383 2553
rect 456 2507 463 2732
rect 556 2507 563 2793
rect 576 2746 583 2816
rect 816 2776 823 2956
rect 916 2947 923 3013
rect 956 2996 963 3233
rect 1096 3207 1103 3294
rect 996 3027 1003 3193
rect 993 3000 1007 3013
rect 996 2996 1003 3000
rect 1036 2963 1043 3173
rect 1076 3008 1083 3073
rect 1116 3067 1123 3476
rect 1193 3467 1207 3480
rect 1216 3387 1223 3433
rect 1136 3263 1143 3333
rect 1236 3287 1243 3353
rect 1136 3256 1163 3263
rect 1016 2956 1043 2963
rect 1096 2960 1103 2963
rect 896 2807 903 2893
rect 956 2816 963 2933
rect 616 2723 623 2743
rect 596 2716 623 2723
rect 76 2256 83 2413
rect 216 2307 223 2473
rect 116 2256 123 2293
rect 96 2107 103 2223
rect 167 1973 173 1987
rect 113 1960 127 1973
rect 196 1963 203 2254
rect 496 2256 503 2493
rect 596 2287 603 2716
rect 676 2687 683 2743
rect 776 2547 783 2743
rect 673 2480 687 2493
rect 676 2476 683 2480
rect 616 2387 623 2473
rect 716 2446 723 2493
rect 776 2476 783 2533
rect 856 2476 863 2673
rect 1016 2667 1023 2956
rect 1093 2947 1107 2960
rect 1156 2947 1163 3233
rect 1216 3227 1223 3263
rect 1216 3187 1223 3213
rect 1256 3207 1263 3673
rect 1316 3587 1323 3813
rect 1336 3787 1343 3814
rect 1416 3816 1423 3873
rect 1453 3827 1467 3833
rect 1496 3823 1503 4153
rect 1516 4007 1523 4253
rect 1576 4247 1583 4336
rect 1596 4287 1603 4393
rect 1636 4207 1643 4753
rect 1696 4556 1703 4753
rect 1716 4567 1723 4673
rect 1736 4547 1743 4573
rect 1756 4567 1763 4816
rect 1776 4807 1783 4853
rect 1796 4727 1803 5233
rect 1916 5087 1923 5343
rect 2016 5163 2023 5373
rect 2036 5287 2043 5473
rect 2096 5376 2103 5413
rect 2116 5307 2123 5343
rect 2016 5156 2043 5163
rect 1996 5107 2003 5133
rect 1880 5043 1893 5047
rect 1836 5040 1843 5043
rect 1833 5027 1847 5040
rect 1876 5036 1893 5043
rect 1880 5033 1893 5036
rect 1916 4887 1923 5052
rect 1947 5043 1960 5047
rect 1947 5036 1963 5043
rect 1947 5033 1960 5036
rect 1833 4860 1847 4873
rect 1836 4856 1843 4860
rect 1876 4856 1923 4863
rect 1793 4568 1807 4573
rect 1833 4560 1847 4573
rect 1856 4563 1863 4823
rect 1916 4767 1923 4856
rect 1936 4847 1943 4913
rect 2016 4896 2023 5113
rect 2036 4927 2043 5156
rect 2056 4927 2063 5193
rect 2076 5076 2083 5273
rect 2056 4856 2083 4863
rect 1936 4820 1963 4823
rect 1933 4816 1963 4820
rect 1933 4807 1947 4816
rect 2076 4767 2083 4856
rect 1836 4556 1843 4560
rect 1856 4556 1883 4563
rect 1667 4523 1680 4527
rect 1667 4516 1683 4523
rect 1667 4513 1680 4516
rect 1656 4127 1663 4303
rect 1696 4167 1703 4473
rect 1736 4227 1743 4512
rect 1756 4296 1783 4303
rect 1756 4187 1763 4296
rect 1816 4287 1823 4523
rect 1876 4363 1883 4556
rect 1996 4527 2003 4573
rect 1916 4367 1923 4523
rect 1876 4356 1903 4363
rect 1896 4336 1903 4356
rect 1936 4336 1943 4473
rect 2016 4367 2023 4593
rect 2056 4568 2063 4693
rect 2096 4647 2103 4913
rect 2156 4856 2163 5373
rect 2176 5347 2183 5473
rect 2587 5416 2613 5423
rect 2636 5407 2643 5433
rect 2593 5380 2607 5393
rect 2596 5376 2603 5380
rect 2196 5076 2203 5213
rect 2276 5207 2283 5343
rect 2636 5307 2643 5393
rect 2367 5116 2393 5123
rect 2373 5080 2387 5093
rect 2376 5076 2383 5080
rect 2256 5007 2263 5043
rect 2196 4856 2203 4913
rect 2236 4826 2243 4913
rect 2296 4868 2303 5074
rect 2396 5023 2403 5032
rect 2376 5016 2403 5023
rect 2136 4767 2143 4823
rect 2176 4787 2183 4823
rect 2336 4787 2343 4893
rect 2376 4868 2383 5016
rect 2436 5007 2443 5133
rect 2496 5088 2503 5293
rect 2656 5267 2663 5473
rect 2876 5447 2883 5523
rect 3256 5487 3263 5523
rect 2713 5407 2727 5413
rect 2736 5376 2743 5433
rect 2813 5407 2827 5413
rect 2596 5076 2603 5173
rect 2676 5088 2683 5293
rect 2476 5007 2483 5043
rect 2476 4927 2483 4993
rect 2516 4967 2523 5032
rect 2416 4856 2423 4893
rect 2556 4887 2563 5073
rect 2696 5046 2703 5193
rect 2756 5076 2763 5133
rect 2796 5087 2803 5393
rect 2816 5376 2843 5383
rect 2816 5207 2823 5376
rect 3016 5347 3023 5433
rect 2816 5046 2823 5153
rect 2856 5076 2863 5253
rect 2916 5207 2923 5343
rect 2976 5336 3003 5343
rect 2996 5267 3003 5336
rect 3036 5307 3043 5453
rect 3147 5413 3153 5427
rect 3187 5416 3213 5423
rect 3193 5388 3207 5393
rect 3236 5376 3243 5453
rect 3136 5323 3143 5374
rect 3127 5316 3143 5323
rect 2656 5007 2663 5043
rect 2736 5007 2743 5043
rect 2396 4803 2403 4823
rect 2396 4796 2423 4803
rect 2096 4556 2103 4593
rect 2136 4556 2143 4633
rect 2236 4487 2243 4554
rect 2256 4387 2263 4753
rect 2356 4526 2363 4573
rect 2376 4507 2383 4593
rect 2416 4587 2423 4796
rect 2416 4556 2423 4573
rect 2456 4556 2463 4733
rect 2476 4727 2483 4854
rect 2516 4727 2523 4823
rect 2556 4787 2563 4823
rect 2596 4667 2603 4873
rect 2636 4856 2643 4953
rect 2367 4486 2380 4487
rect 2367 4473 2373 4486
rect 2407 4473 2413 4487
rect 2013 4340 2027 4353
rect 2073 4340 2087 4353
rect 2016 4336 2023 4340
rect 2076 4336 2083 4340
rect 1876 4227 1883 4303
rect 1916 4300 1923 4303
rect 1913 4287 1927 4300
rect 1576 4036 1583 4073
rect 1656 4036 1663 4113
rect 1756 4087 1763 4173
rect 1556 3847 1563 3992
rect 1756 3927 1763 4034
rect 1596 3867 1603 3893
rect 1776 3887 1783 4213
rect 1896 4048 1903 4273
rect 1976 4036 1983 4253
rect 2036 4227 2043 4303
rect 2016 4048 2023 4193
rect 1476 3816 1503 3823
rect 1440 3783 1453 3787
rect 1276 3367 1283 3533
rect 1313 3520 1327 3533
rect 1316 3516 1323 3520
rect 1396 3407 1403 3783
rect 1436 3776 1453 3783
rect 1440 3773 1453 3776
rect 1476 3528 1483 3816
rect 1596 3787 1603 3853
rect 1516 3707 1523 3772
rect 1296 3296 1303 3333
rect 1356 3207 1363 3263
rect 1276 3007 1283 3053
rect 1093 2780 1107 2793
rect 1136 2787 1143 2893
rect 1176 2787 1183 2953
rect 1216 2867 1223 2963
rect 1276 2847 1283 2953
rect 1096 2776 1103 2780
rect 1193 2780 1207 2793
rect 1196 2776 1203 2780
rect 1236 2776 1243 2833
rect 1036 2746 1043 2773
rect 796 2387 803 2443
rect 956 2407 963 2474
rect 1076 2446 1083 2732
rect 976 2387 983 2433
rect 533 2260 547 2273
rect 536 2256 543 2260
rect 216 2226 223 2253
rect 256 2107 263 2223
rect 296 2216 323 2223
rect 253 1968 267 1973
rect 116 1956 123 1960
rect 176 1956 203 1963
rect 16 1407 23 1692
rect 36 1647 43 1954
rect 176 1923 183 1956
rect 96 1867 103 1923
rect 136 1916 183 1923
rect 236 1903 243 1923
rect 276 1920 283 1923
rect 216 1896 243 1903
rect 273 1907 287 1920
rect 316 1907 323 2216
rect 376 2107 383 2223
rect 416 2167 423 2223
rect 456 2187 463 2253
rect 416 1967 423 2153
rect 516 2147 523 2223
rect 556 2187 563 2223
rect 616 2147 623 2293
rect 953 2260 967 2273
rect 956 2256 963 2260
rect 676 2220 683 2223
rect 673 2207 687 2220
rect 516 2107 523 2133
rect 136 1776 143 1893
rect 56 1623 63 1734
rect 36 1616 63 1623
rect 36 1367 43 1616
rect 76 1507 83 1633
rect 76 1436 83 1493
rect 113 1448 127 1453
rect 16 887 23 1293
rect 36 1186 43 1233
rect 96 1216 103 1353
rect 156 1347 163 1633
rect 196 1467 203 1893
rect 216 1867 223 1896
rect 216 1647 223 1853
rect 296 1736 303 1853
rect 356 1703 363 1753
rect 276 1700 283 1703
rect 273 1687 287 1700
rect 316 1696 363 1703
rect 256 1436 263 1673
rect 296 1403 303 1493
rect 376 1443 383 1833
rect 416 1736 423 1813
rect 436 1807 443 1953
rect 536 1926 543 2033
rect 696 1967 703 2173
rect 716 2027 723 2223
rect 756 2167 763 2253
rect 816 2187 823 2212
rect 853 2207 867 2212
rect 896 2147 903 2254
rect 1016 2226 1023 2293
rect 1076 2256 1083 2333
rect 1096 2307 1103 2533
rect 1176 2483 1183 2733
rect 1256 2740 1263 2743
rect 1253 2727 1267 2740
rect 1296 2707 1303 3193
rect 1336 3008 1343 3113
rect 1496 3107 1503 3633
rect 1536 3516 1543 3693
rect 1576 3547 1583 3713
rect 1576 3516 1583 3533
rect 1596 3528 1603 3573
rect 1556 3407 1563 3483
rect 1516 3207 1523 3393
rect 1596 3303 1603 3473
rect 1616 3467 1623 3873
rect 1636 3783 1643 3833
rect 1696 3816 1723 3823
rect 1636 3776 1663 3783
rect 1716 3647 1723 3816
rect 1736 3816 1783 3823
rect 1816 3816 1823 3913
rect 1836 3867 1843 4003
rect 1856 3827 1863 3993
rect 1896 3927 1903 4034
rect 1956 3907 1963 4003
rect 1996 3967 2003 4003
rect 1976 3828 1983 3853
rect 1736 3707 1743 3816
rect 1636 3347 1643 3593
rect 1716 3587 1723 3633
rect 1736 3627 1743 3693
rect 1716 3387 1723 3443
rect 1776 3407 1783 3613
rect 1796 3387 1803 3783
rect 1836 3707 1843 3783
rect 1876 3727 1883 3814
rect 1916 3780 1923 3783
rect 1896 3687 1903 3773
rect 1913 3767 1927 3780
rect 1996 3747 2003 3783
rect 2013 3767 2027 3773
rect 2036 3763 2043 3993
rect 2056 3967 2063 4003
rect 2136 3907 2143 4373
rect 2256 4223 2263 4303
rect 2236 4216 2263 4223
rect 2236 4187 2243 4216
rect 2236 4127 2243 4173
rect 2236 4036 2243 4113
rect 2276 4006 2283 4093
rect 2296 4087 2303 4373
rect 2316 4307 2323 4334
rect 2336 4306 2343 4393
rect 2436 4348 2443 4433
rect 2496 4343 2503 4653
rect 2573 4560 2587 4573
rect 2576 4556 2583 4560
rect 2556 4487 2563 4523
rect 2596 4487 2603 4523
rect 2636 4467 2643 4793
rect 2656 4767 2663 4823
rect 2656 4607 2663 4673
rect 2696 4647 2703 4893
rect 2756 4856 2763 4953
rect 2736 4787 2743 4812
rect 2796 4767 2803 4993
rect 2876 4856 2883 5013
rect 2896 4907 2903 5043
rect 2916 4888 2923 5193
rect 2936 5027 2943 5133
rect 2956 5087 2963 5253
rect 2987 5136 3013 5143
rect 2996 5076 3003 5113
rect 2976 4947 2983 5043
rect 3076 4967 3083 5113
rect 3116 5076 3123 5313
rect 3156 5247 3163 5353
rect 3296 5343 3303 5473
rect 3313 5387 3327 5393
rect 3476 5376 3483 5523
rect 4516 5516 4543 5523
rect 4616 5516 4643 5523
rect 3776 5388 3783 5413
rect 3836 5376 3843 5413
rect 3416 5346 3423 5373
rect 3216 5340 3223 5343
rect 3256 5340 3263 5343
rect 3213 5327 3227 5340
rect 3253 5327 3267 5340
rect 3276 5336 3303 5343
rect 3176 5087 3183 5113
rect 3133 4907 3147 4913
rect 3087 4893 3093 4907
rect 2856 4820 2863 4823
rect 2853 4807 2867 4820
rect 2956 4826 2963 4893
rect 3116 4867 3123 4893
rect 3176 4867 3183 5033
rect 3256 4987 3263 5173
rect 2696 4616 2743 4623
rect 2696 4587 2703 4616
rect 2687 4578 2703 4587
rect 2687 4574 2700 4578
rect 2680 4573 2700 4574
rect 2716 4556 2723 4593
rect 2736 4587 2743 4616
rect 2476 4336 2503 4343
rect 2536 4336 2543 4393
rect 2416 4283 2423 4303
rect 2396 4276 2423 4283
rect 2396 4227 2403 4276
rect 2056 3827 2063 3893
rect 2236 3816 2243 3973
rect 2273 3827 2287 3833
rect 2036 3756 2053 3763
rect 1853 3467 1867 3472
rect 1576 3296 1603 3303
rect 1776 3296 1803 3303
rect 1576 2996 1583 3173
rect 1356 2907 1363 2963
rect 1396 2907 1403 2963
rect 1476 2927 1483 2993
rect 1496 2907 1503 2933
rect 1616 2867 1623 3252
rect 1796 3227 1803 3296
rect 1636 2966 1643 3073
rect 1696 2996 1703 3113
rect 1816 3067 1823 3393
rect 1736 2996 1783 3003
rect 1816 2996 1823 3053
rect 1836 3047 1843 3293
rect 1856 3008 1863 3373
rect 1896 3367 1903 3483
rect 1916 3336 1923 3472
rect 1936 3427 1943 3733
rect 1996 3647 2003 3733
rect 2056 3487 2063 3753
rect 2116 3747 2123 3783
rect 2136 3707 2143 3773
rect 2156 3747 2163 3814
rect 1976 3387 1983 3483
rect 2056 3383 2063 3413
rect 2076 3407 2083 3673
rect 2216 3607 2223 3783
rect 2296 3727 2303 4073
rect 2316 3827 2323 3953
rect 2336 3927 2343 4003
rect 2376 3887 2383 4003
rect 2347 3843 2360 3847
rect 2347 3833 2363 3843
rect 2356 3816 2363 3833
rect 2416 3828 2423 4233
rect 2476 4107 2483 4336
rect 2556 4283 2563 4303
rect 2536 4276 2563 4283
rect 2480 4063 2493 4067
rect 2476 4053 2493 4063
rect 2476 4036 2483 4053
rect 2453 3987 2467 3992
rect 2376 3747 2383 3783
rect 2336 3607 2343 3713
rect 2396 3627 2403 3753
rect 2176 3487 2183 3514
rect 2056 3376 2083 3383
rect 2016 3308 2023 3353
rect 2076 3147 2083 3376
rect 1696 2907 1703 2933
rect 1716 2927 1723 2963
rect 1776 2907 1783 2996
rect 1896 2966 1903 3033
rect 1360 2743 1373 2747
rect 1356 2736 1373 2743
rect 1360 2733 1373 2736
rect 1396 2727 1403 2774
rect 1416 2746 1423 2793
rect 1447 2783 1460 2787
rect 1447 2776 1463 2783
rect 1493 2780 1507 2793
rect 1496 2776 1503 2780
rect 1447 2773 1460 2776
rect 1633 2787 1647 2793
rect 1176 2476 1193 2483
rect 1256 2476 1263 2533
rect 1196 2447 1203 2474
rect 1276 2407 1283 2443
rect 1356 2407 1363 2693
rect 1476 2667 1483 2743
rect 1536 2727 1543 2773
rect 1656 2746 1663 2773
rect 1576 2687 1583 2743
rect 1656 2707 1663 2732
rect 1673 2727 1687 2733
rect 1396 2476 1403 2533
rect 1736 2507 1743 2553
rect 1676 2476 1703 2483
rect 1476 2427 1483 2453
rect 1267 2376 1293 2383
rect 1207 2274 1213 2287
rect 1200 2273 1220 2274
rect 1327 2283 1340 2287
rect 1327 2273 1343 2283
rect 1336 2256 1343 2273
rect 936 2187 943 2212
rect 1096 2187 1103 2223
rect 1216 2220 1223 2223
rect 1213 2207 1227 2220
rect 816 2027 823 2133
rect 856 2047 863 2093
rect 640 1923 653 1927
rect 496 1847 503 1912
rect 596 1827 603 1923
rect 636 1916 653 1923
rect 640 1913 653 1916
rect 676 1867 683 1954
rect 816 1927 823 2013
rect 856 1956 863 2033
rect 896 1956 903 2053
rect 696 1827 703 1913
rect 436 1767 443 1793
rect 436 1687 443 1703
rect 427 1676 443 1687
rect 427 1673 440 1676
rect 476 1487 483 1813
rect 596 1787 603 1813
rect 616 1748 623 1813
rect 656 1736 663 1773
rect 696 1736 703 1813
rect 736 1747 743 1923
rect 776 1920 783 1923
rect 773 1907 787 1920
rect 876 1920 883 1923
rect 873 1907 887 1920
rect 956 1907 963 2013
rect 1013 1960 1027 1973
rect 1016 1956 1023 1960
rect 1076 1967 1083 2053
rect 1153 1968 1167 1973
rect 1036 1920 1043 1923
rect 376 1436 403 1443
rect 436 1436 443 1473
rect 496 1463 503 1693
rect 536 1667 543 1703
rect 616 1627 623 1734
rect 856 1747 863 1793
rect 716 1700 723 1703
rect 476 1456 503 1463
rect 476 1436 483 1456
rect 396 1406 403 1436
rect 536 1407 543 1613
rect 596 1436 603 1513
rect 147 1233 153 1247
rect 176 1227 183 1393
rect 196 1307 203 1403
rect 236 1347 243 1403
rect 276 1396 303 1403
rect 233 1220 247 1233
rect 276 1228 283 1396
rect 356 1383 363 1403
rect 336 1376 363 1383
rect 236 1216 243 1220
rect 36 367 43 1172
rect 93 928 107 933
rect 153 923 167 933
rect 136 920 167 923
rect 136 916 163 920
rect 176 907 183 1172
rect 256 1127 263 1183
rect 336 1167 343 1376
rect 456 1228 463 1403
rect 616 1287 623 1403
rect 656 1327 663 1393
rect 676 1307 683 1692
rect 713 1687 727 1700
rect 756 1587 763 1733
rect 896 1706 903 1773
rect 956 1736 963 1853
rect 996 1787 1003 1912
rect 1033 1907 1047 1920
rect 1096 1847 1103 1954
rect 1216 1923 1223 2053
rect 1256 2007 1263 2212
rect 1296 2187 1303 2254
rect 1393 2207 1407 2212
rect 1336 1967 1343 2173
rect 1436 1987 1443 2413
rect 1496 2367 1503 2474
rect 1616 2436 1643 2443
rect 1476 2256 1483 2293
rect 1556 2267 1563 2413
rect 1636 2307 1643 2436
rect 1676 2347 1683 2476
rect 1796 2476 1803 2593
rect 1836 2567 1843 2963
rect 1896 2807 1903 2952
rect 1976 2907 1983 2953
rect 2016 2907 2023 3053
rect 2036 2996 2043 3133
rect 1856 2687 1863 2774
rect 1956 2667 1963 2743
rect 1956 2607 1963 2653
rect 1896 2367 1903 2573
rect 2016 2446 2023 2793
rect 2036 2787 2043 2833
rect 2056 2807 2063 2893
rect 2076 2867 2083 2963
rect 2096 2907 2103 3473
rect 2116 3367 2123 3483
rect 2216 3463 2223 3483
rect 2216 3456 2243 3463
rect 2196 3260 2203 3263
rect 2193 3247 2207 3260
rect 2196 3187 2203 3233
rect 2236 3087 2243 3456
rect 2256 3287 2263 3483
rect 2316 3427 2323 3514
rect 2336 3263 2343 3593
rect 2416 3587 2423 3673
rect 2436 3647 2443 3913
rect 2496 3847 2503 4003
rect 2536 3847 2543 4276
rect 2576 4036 2583 4153
rect 2596 4067 2603 4452
rect 2656 4447 2663 4513
rect 2696 4487 2703 4523
rect 2776 4523 2783 4713
rect 2756 4516 2783 4523
rect 2656 4336 2663 4393
rect 2636 4267 2643 4303
rect 2676 4283 2683 4303
rect 2676 4276 2703 4283
rect 2696 4207 2703 4276
rect 2716 4227 2723 4293
rect 2736 4287 2743 4334
rect 2613 4040 2627 4053
rect 2676 4048 2683 4173
rect 2756 4147 2763 4516
rect 2796 4348 2803 4753
rect 2816 4407 2823 4633
rect 2836 4627 2843 4693
rect 2896 4607 2903 4673
rect 2833 4560 2847 4573
rect 2836 4556 2843 4560
rect 2896 4556 2903 4593
rect 2836 4336 2843 4453
rect 2936 4367 2943 4813
rect 2996 4807 3003 4823
rect 2956 4407 2963 4653
rect 2976 4556 2983 4733
rect 2996 4587 3003 4793
rect 3036 4787 3043 4812
rect 3096 4707 3103 4853
rect 3156 4820 3163 4823
rect 3113 4807 3127 4813
rect 3153 4807 3167 4820
rect 3176 4747 3183 4813
rect 3016 4503 3023 4523
rect 2996 4496 3023 4503
rect 2616 4036 2623 4040
rect 2756 4043 2763 4073
rect 2736 4036 2763 4043
rect 2596 4000 2603 4003
rect 2593 3987 2607 4000
rect 2533 3820 2547 3833
rect 2636 3823 2643 4003
rect 2776 3847 2783 4033
rect 2796 4007 2803 4273
rect 2816 4227 2823 4303
rect 2876 4300 2883 4303
rect 2873 4287 2887 4300
rect 2936 4296 2963 4303
rect 2536 3816 2543 3820
rect 2616 3816 2643 3823
rect 2856 3823 2863 3992
rect 2896 3887 2903 4073
rect 2916 4007 2923 4193
rect 2956 4107 2963 4296
rect 2976 4287 2983 4353
rect 2996 4247 3003 4496
rect 3036 4447 3043 4573
rect 3096 4568 3103 4693
rect 3196 4587 3203 4973
rect 3276 4947 3283 5336
rect 3496 5227 3503 5343
rect 3716 5340 3723 5343
rect 3296 5083 3303 5133
rect 3436 5088 3443 5193
rect 3516 5103 3523 5173
rect 3496 5096 3523 5103
rect 3296 5076 3323 5083
rect 3496 5076 3503 5096
rect 3216 4827 3223 4913
rect 3236 4867 3243 4933
rect 3256 4868 3263 4893
rect 3296 4887 3303 4993
rect 3296 4856 3303 4873
rect 3336 4823 3343 4873
rect 3396 4856 3403 5033
rect 3536 4856 3543 4893
rect 3556 4887 3563 5213
rect 3616 5007 3623 5043
rect 3656 5007 3663 5332
rect 3713 5327 3727 5340
rect 3716 5207 3723 5313
rect 3736 5307 3743 5373
rect 3776 5347 3783 5374
rect 3676 5043 3683 5074
rect 3676 5036 3703 5043
rect 3616 4967 3623 4993
rect 3336 4816 3383 4823
rect 3256 4727 3263 4793
rect 3180 4566 3200 4567
rect 3180 4563 3193 4566
rect 3176 4556 3193 4563
rect 3180 4553 3193 4556
rect 3216 4527 3223 4713
rect 3276 4556 3283 4633
rect 3056 4427 3063 4512
rect 3116 4447 3123 4523
rect 3193 4503 3207 4513
rect 3176 4500 3207 4503
rect 3176 4496 3203 4500
rect 3056 4336 3103 4343
rect 2996 4207 3003 4233
rect 3096 4187 3103 4336
rect 3116 4287 3123 4433
rect 3176 4336 3183 4496
rect 3316 4487 3323 4673
rect 3396 4568 3403 4733
rect 3476 4707 3483 4833
rect 3560 4823 3573 4827
rect 3516 4820 3523 4823
rect 3513 4807 3527 4820
rect 3556 4816 3573 4823
rect 3560 4813 3573 4816
rect 3596 4667 3603 4873
rect 3613 4867 3627 4873
rect 3696 4868 3703 5036
rect 3736 4967 3743 5043
rect 3756 4947 3763 4993
rect 3676 4787 3683 4823
rect 3336 4467 3343 4513
rect 3413 4507 3427 4513
rect 3436 4427 3443 4593
rect 3156 4300 3163 4303
rect 3153 4287 3167 4300
rect 3196 4187 3203 4303
rect 2953 4048 2967 4053
rect 3056 3907 3063 4034
rect 3087 4043 3100 4047
rect 3087 4036 3103 4043
rect 3133 4040 3147 4053
rect 3176 4047 3183 4133
rect 3136 4036 3143 4040
rect 3087 4033 3100 4036
rect 3196 4007 3203 4093
rect 3236 4067 3243 4393
rect 3296 4336 3303 4393
rect 3456 4343 3463 4633
rect 3487 4563 3500 4567
rect 3487 4556 3503 4563
rect 3536 4556 3543 4633
rect 3596 4587 3603 4613
rect 3487 4553 3500 4556
rect 3656 4527 3663 4593
rect 3516 4487 3523 4523
rect 3596 4467 3603 4523
rect 3456 4336 3483 4343
rect 3276 4247 3283 4303
rect 3316 4283 3323 4303
rect 3376 4300 3383 4303
rect 3296 4276 3323 4283
rect 3373 4287 3387 4300
rect 3296 4147 3303 4276
rect 3256 4036 3263 4093
rect 3293 4040 3307 4053
rect 3316 4047 3323 4193
rect 3296 4036 3303 4040
rect 2856 3816 2883 3823
rect 2616 3786 2623 3816
rect 2876 3786 2883 3816
rect 2496 3780 2503 3783
rect 2493 3767 2507 3780
rect 2896 3587 2903 3873
rect 3016 3816 3023 3873
rect 3076 3828 3083 3993
rect 3156 3967 3163 4003
rect 3236 3947 3243 4003
rect 3076 3786 3083 3814
rect 3096 3687 3103 3873
rect 3296 3816 3303 3973
rect 3336 3947 3343 4233
rect 3353 4047 3367 4053
rect 3376 4036 3383 4173
rect 3416 4067 3423 4093
rect 3476 4087 3483 4336
rect 3596 4247 3603 4353
rect 3656 4336 3663 4413
rect 3676 4367 3683 4653
rect 3696 4563 3703 4673
rect 3736 4647 3743 4893
rect 3776 4887 3783 5193
rect 3816 5087 3823 5273
rect 3856 5207 3863 5343
rect 3956 5307 3963 5353
rect 3976 5127 3983 5413
rect 4316 5346 4323 5393
rect 3996 5336 4023 5343
rect 4076 5340 4083 5343
rect 3996 5287 4003 5336
rect 4073 5327 4087 5340
rect 4416 5340 4423 5343
rect 4413 5327 4427 5340
rect 4456 5307 4463 5353
rect 4476 5347 4483 5393
rect 4536 5376 4543 5516
rect 4636 5376 4643 5516
rect 5336 5376 5383 5383
rect 5456 5376 5463 5413
rect 3836 5076 3843 5113
rect 4016 5088 4023 5153
rect 3796 4868 3803 5033
rect 3896 5036 3913 5043
rect 3896 4847 3903 4873
rect 3767 4823 3780 4827
rect 3767 4813 3783 4823
rect 3776 4707 3783 4813
rect 3696 4556 3723 4563
rect 3776 4556 3783 4593
rect 3796 4567 3803 4653
rect 3736 4348 3743 4433
rect 3816 4336 3823 4793
rect 3836 4367 3843 4693
rect 3896 4643 3903 4833
rect 3916 4747 3923 5033
rect 3936 5007 3943 5074
rect 3996 5040 4003 5043
rect 3993 5027 4007 5040
rect 4047 5016 4073 5023
rect 3956 4820 3963 4823
rect 3953 4807 3967 4820
rect 3876 4636 3903 4643
rect 3876 4587 3883 4636
rect 3933 4567 3947 4573
rect 3956 4526 3963 4613
rect 3976 4567 3983 4733
rect 4013 4560 4027 4573
rect 4056 4567 4063 4993
rect 4076 4747 4083 4933
rect 4116 4863 4123 5133
rect 4233 5080 4247 5093
rect 4236 5076 4243 5080
rect 4136 5007 4143 5074
rect 4096 4856 4123 4863
rect 4016 4556 4023 4560
rect 3876 4487 3883 4523
rect 3987 4523 4000 4527
rect 3987 4516 4003 4523
rect 3987 4513 4000 4516
rect 3887 4476 3903 4483
rect 3413 4040 3427 4053
rect 3416 4036 3423 4040
rect 3456 4006 3463 4053
rect 3476 3967 3483 4052
rect 3533 4040 3547 4053
rect 3536 4036 3543 4040
rect 3347 3936 3363 3943
rect 2416 3486 2423 3573
rect 2473 3528 2487 3533
rect 2593 3520 2607 3533
rect 2596 3516 2603 3520
rect 2713 3520 2727 3533
rect 3036 3528 3043 3573
rect 2716 3516 2723 3520
rect 2436 3383 2443 3513
rect 2496 3407 2503 3483
rect 2436 3376 2463 3383
rect 2316 3256 2343 3263
rect 2436 3260 2443 3263
rect 2433 3247 2447 3260
rect 2153 3000 2167 3013
rect 2156 2996 2163 3000
rect 2196 2996 2203 3033
rect 2236 2966 2243 3033
rect 2273 3000 2287 3013
rect 2276 2996 2283 3000
rect 2316 2996 2323 3113
rect 2296 2927 2303 2963
rect 2416 2867 2423 3013
rect 2056 2776 2063 2793
rect 2096 2776 2103 2833
rect 2376 2827 2383 2853
rect 2120 2743 2133 2747
rect 2116 2736 2133 2743
rect 2120 2733 2133 2736
rect 2156 2746 2163 2793
rect 2173 2787 2187 2793
rect 2036 2443 2043 2732
rect 2196 2687 2203 2743
rect 2276 2707 2283 2774
rect 2336 2707 2343 2743
rect 2436 2727 2443 3233
rect 2456 3027 2463 3376
rect 2556 3327 2563 3514
rect 2493 3300 2507 3313
rect 2496 3296 2503 3300
rect 2576 3247 2583 3453
rect 2616 3427 2623 3483
rect 2676 3387 2683 3514
rect 2736 3447 2743 3483
rect 2776 3427 2783 3473
rect 2896 3467 2903 3514
rect 3036 3487 3043 3514
rect 2716 3287 2723 3333
rect 2736 3267 2743 3313
rect 2896 3303 2903 3453
rect 3056 3407 3063 3653
rect 3196 3647 3203 3783
rect 3116 3463 3123 3483
rect 3096 3456 3123 3463
rect 2887 3296 2903 3303
rect 2936 3296 2943 3333
rect 2976 3296 2983 3393
rect 2676 3260 2683 3263
rect 2673 3247 2687 3260
rect 2556 3236 2573 3243
rect 2556 3003 2563 3236
rect 2816 3087 2823 3263
rect 2536 2996 2563 3003
rect 2636 2996 2643 3033
rect 2676 2996 2683 3073
rect 2736 2967 2743 2994
rect 2696 2927 2703 2963
rect 2876 2927 2883 3294
rect 2956 3243 2963 3263
rect 2936 3236 2963 3243
rect 2896 2966 2903 3033
rect 2936 3008 2943 3236
rect 3076 3227 3083 3294
rect 3076 3167 3083 3213
rect 3096 3083 3103 3456
rect 3156 3407 3163 3633
rect 3356 3607 3363 3936
rect 3496 3927 3503 4003
rect 3376 3887 3383 3913
rect 3476 3823 3483 3893
rect 3476 3816 3493 3823
rect 3376 3707 3383 3813
rect 3416 3747 3423 3772
rect 3456 3647 3463 3713
rect 3216 3516 3223 3553
rect 3196 3480 3203 3483
rect 3193 3467 3207 3480
rect 3236 3427 3243 3472
rect 3336 3467 3343 3573
rect 3236 3263 3243 3392
rect 3296 3296 3303 3353
rect 3356 3327 3363 3593
rect 3456 3516 3463 3633
rect 3496 3347 3503 3533
rect 3516 3467 3523 3613
rect 3556 3547 3563 4073
rect 3576 3667 3583 4153
rect 3596 4003 3603 4193
rect 3616 4187 3623 4313
rect 3656 4036 3663 4193
rect 3676 4147 3683 4303
rect 3716 4043 3723 4073
rect 3736 4067 3743 4334
rect 3876 4306 3883 4393
rect 3896 4347 3903 4476
rect 3916 4407 3923 4473
rect 3936 4363 3943 4433
rect 3916 4356 3943 4363
rect 3916 4336 3923 4356
rect 3956 4336 3963 4393
rect 3976 4387 3983 4492
rect 4007 4473 4013 4487
rect 3716 4036 3743 4043
rect 3773 4040 3787 4053
rect 3776 4036 3783 4040
rect 3596 3996 3623 4003
rect 3753 3987 3767 3992
rect 3716 3786 3723 3813
rect 3676 3727 3683 3783
rect 3736 3587 3743 3913
rect 3836 3887 3843 4303
rect 3936 4283 3943 4303
rect 3936 4276 3953 4283
rect 3856 4047 3863 4133
rect 3916 4067 3923 4193
rect 3893 4040 3907 4053
rect 3936 4047 3943 4253
rect 3896 4036 3903 4040
rect 3876 4000 3883 4003
rect 3873 3987 3887 4000
rect 3896 3827 3903 3933
rect 3916 3887 3923 3953
rect 3936 3947 3943 3993
rect 3956 3967 3963 4273
rect 3996 4267 4003 4293
rect 3976 4147 3983 4253
rect 3996 4107 4003 4173
rect 4016 4167 4023 4433
rect 4036 4427 4043 4523
rect 4056 4403 4063 4513
rect 4036 4396 4063 4403
rect 4036 4347 4043 4396
rect 4076 4336 4083 4473
rect 4096 4447 4103 4856
rect 4136 4747 4143 4823
rect 4156 4787 4163 4853
rect 4276 4567 4283 5233
rect 4516 5147 4523 5343
rect 4616 5247 4623 5343
rect 4676 5207 4683 5374
rect 4716 5307 4723 5343
rect 4796 5287 4803 5343
rect 4296 4827 4303 5093
rect 4436 5043 4443 5073
rect 4556 5043 4563 5113
rect 4616 5076 4623 5133
rect 4356 5007 4363 5043
rect 4396 5036 4443 5043
rect 4476 4927 4483 5043
rect 4516 5036 4563 5043
rect 4376 4820 4383 4823
rect 4296 4747 4303 4813
rect 4373 4807 4387 4820
rect 4416 4767 4423 4823
rect 4296 4556 4303 4613
rect 4416 4607 4423 4753
rect 4456 4727 4463 4873
rect 4516 4856 4523 4953
rect 4496 4820 4503 4823
rect 4493 4807 4507 4820
rect 4556 4767 4563 4913
rect 4576 4887 4583 5033
rect 4596 4927 4603 5043
rect 4656 4947 4663 5074
rect 4676 5047 4683 5193
rect 4756 5107 4763 5133
rect 4816 5127 4823 5153
rect 4836 5107 4843 5133
rect 4756 5076 4763 5093
rect 4856 5088 4863 5233
rect 4896 5207 4903 5343
rect 4976 5343 4983 5374
rect 4956 5336 4983 5343
rect 4816 5046 4823 5073
rect 4916 5046 4923 5153
rect 4956 5088 4963 5336
rect 5096 5287 5103 5343
rect 5136 5247 5143 5374
rect 5376 5347 5383 5376
rect 5696 5376 5703 5413
rect 4736 5007 4743 5043
rect 5016 5046 5023 5093
rect 5113 5088 5127 5093
rect 5156 5046 5163 5173
rect 5196 5147 5203 5343
rect 5416 5340 5423 5343
rect 5316 5327 5323 5332
rect 5316 5316 5333 5327
rect 5320 5313 5333 5316
rect 5376 5187 5383 5333
rect 5413 5327 5427 5340
rect 5476 5167 5483 5343
rect 5516 5127 5523 5374
rect 5636 5346 5643 5374
rect 5456 5076 5463 5113
rect 4616 4856 4623 4893
rect 4656 4856 4663 4933
rect 4696 4827 4703 4893
rect 4733 4860 4747 4873
rect 4736 4856 4743 4860
rect 4776 4856 4783 4893
rect 4816 4887 4823 5032
rect 4916 4947 4923 4993
rect 4576 4816 4603 4823
rect 4636 4820 4643 4823
rect 4436 4568 4443 4593
rect 4456 4567 4463 4613
rect 4176 4423 4183 4483
rect 4176 4416 4203 4423
rect 4116 4367 4123 4393
rect 4056 4300 4063 4303
rect 4053 4287 4067 4300
rect 4096 4267 4103 4292
rect 3976 4047 3983 4073
rect 3993 4040 4007 4053
rect 4036 4048 4043 4233
rect 4056 4127 4063 4252
rect 3996 4036 4003 4040
rect 4156 4043 4163 4113
rect 4196 4043 4203 4416
rect 4236 4343 4243 4553
rect 4316 4487 4323 4523
rect 4356 4487 4363 4554
rect 4216 4336 4243 4343
rect 4216 4147 4223 4336
rect 4316 4300 4323 4303
rect 4313 4287 4327 4300
rect 4376 4247 4383 4453
rect 4436 4336 4443 4493
rect 4476 4467 4483 4653
rect 4496 4467 4503 4713
rect 4516 4607 4523 4633
rect 4576 4627 4583 4816
rect 4633 4807 4647 4820
rect 4676 4787 4683 4813
rect 4756 4787 4763 4823
rect 4816 4747 4823 4823
rect 4553 4560 4567 4573
rect 4556 4556 4563 4560
rect 4596 4556 4603 4593
rect 4516 4443 4523 4513
rect 4616 4483 4623 4513
rect 4587 4476 4623 4483
rect 4496 4436 4523 4443
rect 4496 4407 4503 4436
rect 4416 4267 4423 4303
rect 4456 4227 4463 4303
rect 4556 4296 4583 4303
rect 4493 4287 4507 4292
rect 4136 4036 4163 4043
rect 4176 4036 4203 4043
rect 3956 3927 3963 3953
rect 3973 3947 3987 3953
rect 4016 3923 4023 4003
rect 3996 3916 4023 3923
rect 3776 3707 3783 3783
rect 3816 3763 3823 3783
rect 3816 3756 3843 3763
rect 3816 3687 3823 3713
rect 3836 3707 3843 3756
rect 3876 3747 3883 3814
rect 3953 3820 3967 3833
rect 3996 3827 4003 3916
rect 4056 3907 4063 3993
rect 4176 3947 4183 4036
rect 3956 3816 3963 3820
rect 4016 3816 4023 3893
rect 3576 3516 3583 3553
rect 3516 3327 3523 3453
rect 3196 3256 3243 3263
rect 3316 3260 3323 3263
rect 3313 3247 3327 3260
rect 3087 3076 3103 3083
rect 3076 2996 3083 3073
rect 3236 3027 3243 3233
rect 3233 3000 3247 3013
rect 3236 2996 3243 3000
rect 2476 2788 2483 2853
rect 2647 2796 2703 2803
rect 2596 2767 2603 2793
rect 2696 2776 2703 2796
rect 2556 2740 2563 2743
rect 2553 2727 2567 2740
rect 2616 2727 2623 2773
rect 2456 2667 2463 2713
rect 2096 2476 2103 2513
rect 2176 2447 2183 2474
rect 2036 2436 2063 2443
rect 1456 1968 1463 2013
rect 1536 1956 1543 2173
rect 1576 2067 1583 2293
rect 1756 2256 1763 2293
rect 1816 2226 1823 2293
rect 1616 2187 1623 2223
rect 1656 2216 1683 2223
rect 1573 1960 1587 1973
rect 1576 1956 1583 1960
rect 1116 1736 1123 1913
rect 1136 1887 1143 1923
rect 1176 1916 1223 1923
rect 796 1567 803 1703
rect 756 1436 763 1473
rect 696 1367 703 1393
rect 536 1228 543 1253
rect 213 920 227 933
rect 253 928 267 933
rect 216 916 223 920
rect 336 927 343 1153
rect 396 1147 403 1183
rect 436 1180 443 1183
rect 433 1167 447 1180
rect 416 928 423 1013
rect 116 880 123 883
rect 113 867 127 880
rect 280 883 293 887
rect 116 747 123 773
rect 76 696 83 733
rect 136 727 143 853
rect 136 667 143 713
rect 156 707 163 813
rect 176 807 183 853
rect 196 787 203 873
rect 216 747 223 853
rect 236 807 243 883
rect 276 876 293 883
rect 280 873 293 876
rect 316 803 323 914
rect 436 927 443 1132
rect 496 1127 503 1214
rect 336 827 343 873
rect 316 796 343 803
rect 193 700 207 713
rect 196 696 203 700
rect 156 523 163 653
rect 276 663 283 793
rect 316 727 323 796
rect 336 743 343 796
rect 356 767 363 883
rect 456 867 463 1113
rect 596 967 603 1233
rect 616 1227 623 1273
rect 653 1220 667 1233
rect 656 1216 663 1220
rect 696 1216 703 1353
rect 736 1307 743 1403
rect 776 1267 783 1403
rect 816 1323 823 1473
rect 836 1447 843 1633
rect 976 1627 983 1703
rect 1036 1647 1043 1734
rect 1096 1627 1103 1703
rect 1176 1703 1183 1873
rect 1216 1847 1223 1873
rect 1256 1807 1263 1923
rect 1276 1736 1283 1833
rect 1296 1747 1303 1793
rect 1316 1767 1323 1893
rect 1356 1847 1363 1933
rect 1387 1923 1400 1927
rect 1387 1916 1403 1923
rect 1387 1913 1400 1916
rect 1436 1887 1443 1923
rect 1176 1696 1203 1703
rect 1133 1687 1147 1692
rect 916 1436 923 1493
rect 847 1403 860 1407
rect 847 1396 863 1403
rect 847 1393 860 1396
rect 856 1327 863 1373
rect 816 1316 843 1323
rect 816 1216 823 1273
rect 836 1247 843 1316
rect 856 1227 863 1313
rect 896 1287 903 1403
rect 936 1327 943 1353
rect 636 1107 643 1183
rect 676 1127 683 1183
rect 736 1007 743 1213
rect 796 1180 803 1183
rect 793 1167 807 1180
rect 876 1167 883 1233
rect 936 1216 943 1313
rect 956 1223 963 1573
rect 1016 1436 1023 1473
rect 996 1400 1003 1403
rect 993 1387 1007 1400
rect 1036 1307 1043 1403
rect 1076 1367 1083 1493
rect 1116 1436 1123 1573
rect 1156 1436 1163 1473
rect 1136 1400 1143 1403
rect 1133 1387 1147 1400
rect 1196 1387 1203 1696
rect 1216 1667 1223 1703
rect 1316 1667 1323 1753
rect 1356 1736 1363 1833
rect 1380 1703 1393 1707
rect 1376 1696 1393 1703
rect 1380 1693 1393 1696
rect 1416 1647 1423 1853
rect 1436 1747 1443 1873
rect 1476 1867 1483 1913
rect 1496 1827 1503 1954
rect 1473 1740 1487 1753
rect 1476 1736 1483 1740
rect 1276 1436 1283 1513
rect 956 1216 983 1223
rect 1033 1220 1047 1233
rect 1036 1216 1043 1220
rect 516 916 523 953
rect 556 928 563 953
rect 636 947 643 993
rect 976 987 983 1216
rect 336 740 363 743
rect 336 736 367 740
rect 353 727 367 736
rect 376 696 383 853
rect 396 707 403 753
rect 276 656 323 663
rect 356 660 363 663
rect 156 516 183 523
rect 156 396 163 473
rect 176 407 183 516
rect 256 507 263 653
rect 353 647 367 660
rect 416 567 423 853
rect 496 807 503 883
rect 596 867 603 932
rect 696 928 703 953
rect 453 700 467 713
rect 493 700 507 713
rect 456 696 463 700
rect 496 696 503 700
rect 476 660 483 663
rect 473 647 487 660
rect 516 627 523 663
rect 116 307 123 333
rect 136 267 143 363
rect 96 176 103 253
rect 196 176 203 473
rect 216 407 223 433
rect 253 400 267 413
rect 256 396 263 400
rect 336 367 343 433
rect 216 327 223 353
rect 256 147 263 333
rect 276 327 283 363
rect 316 307 323 333
rect 356 327 363 413
rect 416 396 423 493
rect 516 403 523 493
rect 536 427 543 653
rect 556 647 563 853
rect 596 696 603 813
rect 636 767 643 883
rect 676 847 683 872
rect 696 727 703 813
rect 736 807 743 914
rect 756 747 763 873
rect 776 863 783 883
rect 776 856 803 863
rect 673 708 687 713
rect 616 660 623 663
rect 613 647 627 660
rect 696 666 703 713
rect 713 707 727 713
rect 796 708 803 856
rect 816 807 823 883
rect 816 707 823 733
rect 676 627 683 653
rect 736 660 743 663
rect 733 647 747 660
rect 776 607 783 663
rect 816 607 823 653
rect 836 647 843 753
rect 856 747 863 813
rect 876 767 883 953
rect 976 916 983 952
rect 1016 886 1023 1183
rect 1076 1147 1083 1233
rect 896 807 903 873
rect 916 847 923 883
rect 896 696 903 793
rect 976 696 983 773
rect 1013 700 1027 713
rect 1036 707 1043 973
rect 1096 948 1103 1373
rect 1196 1307 1203 1373
rect 1216 1287 1223 1393
rect 1256 1367 1263 1403
rect 1176 987 1183 1183
rect 1196 1107 1203 1233
rect 1216 987 1223 1273
rect 1256 1247 1263 1353
rect 1316 1347 1323 1473
rect 1336 1387 1343 1633
rect 1376 1447 1383 1533
rect 1456 1507 1463 1703
rect 1536 1703 1543 1873
rect 1556 1847 1563 1923
rect 1596 1847 1603 1913
rect 1616 1887 1623 1973
rect 1636 1967 1643 2013
rect 1656 1968 1663 2113
rect 1676 1987 1683 2216
rect 1736 2167 1743 2223
rect 1696 1956 1703 2013
rect 1736 1987 1743 2153
rect 1776 2127 1783 2212
rect 1836 2207 1843 2353
rect 1916 2303 1923 2413
rect 1916 2296 1943 2303
rect 1876 2256 1883 2293
rect 1756 1967 1763 2053
rect 1836 2047 1843 2093
rect 1896 2027 1903 2223
rect 1873 1968 1887 1973
rect 1740 1963 1753 1967
rect 1736 1956 1753 1963
rect 1740 1953 1753 1956
rect 1896 1967 1903 2013
rect 1916 1987 1923 2193
rect 1936 2167 1943 2296
rect 1976 2167 1983 2223
rect 2016 2216 2043 2223
rect 1976 2007 1983 2153
rect 1636 1807 1643 1913
rect 1676 1887 1683 1912
rect 1756 1887 1763 1912
rect 1876 1907 1883 1954
rect 1933 1960 1947 1973
rect 1996 1963 2003 2193
rect 1936 1956 1943 1960
rect 1976 1956 2003 1963
rect 1907 1923 1920 1927
rect 1907 1916 1923 1923
rect 1907 1913 1920 1916
rect 1516 1696 1543 1703
rect 1367 1436 1383 1447
rect 1416 1436 1423 1473
rect 1516 1448 1523 1696
rect 1656 1703 1663 1833
rect 1636 1696 1663 1703
rect 1536 1547 1543 1673
rect 1367 1433 1380 1436
rect 1556 1436 1563 1473
rect 1576 1447 1583 1613
rect 1276 1228 1283 1333
rect 1313 1220 1327 1233
rect 1356 1227 1363 1393
rect 1316 1216 1323 1220
rect 1256 987 1263 1172
rect 1296 1127 1303 1183
rect 1347 1176 1363 1183
rect 1076 767 1083 883
rect 1116 880 1123 883
rect 1113 867 1127 880
rect 1176 823 1183 933
rect 1216 916 1223 973
rect 1276 923 1283 993
rect 1256 916 1283 923
rect 1236 880 1243 883
rect 1233 867 1247 880
rect 1156 816 1183 823
rect 1156 767 1163 816
rect 1296 787 1303 893
rect 1016 696 1023 700
rect 876 660 883 663
rect 873 647 887 660
rect 936 627 943 673
rect 776 447 783 473
rect 516 396 543 403
rect 316 176 323 293
rect 416 283 423 313
rect 436 307 443 363
rect 416 276 453 283
rect 436 227 443 253
rect 436 176 443 213
rect 476 176 483 293
rect 496 207 503 394
rect 556 360 563 363
rect 596 360 603 363
rect 553 347 567 360
rect 593 347 607 360
rect 576 316 613 323
rect 576 287 583 316
rect 596 176 603 293
rect 636 207 643 413
rect 673 400 687 413
rect 676 396 683 400
rect 696 327 703 363
rect 736 327 743 363
rect 756 247 763 353
rect 696 187 703 213
rect 636 176 683 183
rect 116 107 123 143
rect 336 107 343 143
rect 456 140 463 143
rect 453 127 467 140
rect 496 107 503 143
rect 536 47 543 173
rect 576 107 583 132
rect 613 127 627 132
rect 676 107 683 176
rect 736 176 743 213
rect 776 176 783 433
rect 856 427 863 473
rect 956 447 963 653
rect 996 607 1003 663
rect 1056 647 1063 733
rect 1096 696 1103 753
rect 1136 696 1143 733
rect 1176 696 1183 773
rect 1316 747 1323 1133
rect 1356 916 1363 1176
rect 1376 1167 1383 1373
rect 1393 1227 1407 1233
rect 1436 1216 1443 1333
rect 1476 1267 1483 1434
rect 1536 1327 1543 1392
rect 1596 1307 1603 1573
rect 1636 1487 1643 1696
rect 1676 1627 1683 1734
rect 1656 1567 1663 1593
rect 1696 1587 1703 1753
rect 1756 1748 1763 1873
rect 1716 1700 1723 1703
rect 1713 1687 1727 1700
rect 1776 1507 1783 1703
rect 1796 1487 1803 1734
rect 1816 1687 1823 1891
rect 1836 1563 1843 1893
rect 1896 1867 1903 1913
rect 1856 1736 1863 1793
rect 1836 1556 1853 1563
rect 1856 1448 1863 1553
rect 1627 1403 1640 1407
rect 1627 1396 1643 1403
rect 1627 1393 1640 1396
rect 1676 1327 1683 1403
rect 1473 1228 1487 1232
rect 1416 1107 1423 1183
rect 1396 928 1403 1053
rect 833 400 847 413
rect 836 396 843 400
rect 893 407 907 413
rect 976 396 983 453
rect 1016 408 1023 493
rect 816 307 823 363
rect 956 327 963 363
rect 996 307 1003 352
rect 1056 287 1063 553
rect 1096 427 1103 633
rect 1116 547 1123 652
rect 1156 627 1163 652
rect 1196 467 1203 593
rect 1093 400 1107 413
rect 1096 396 1103 400
rect 1136 396 1143 433
rect 1216 427 1223 693
rect 1236 666 1243 733
rect 1336 727 1343 813
rect 1356 708 1363 853
rect 1376 787 1383 883
rect 1416 827 1423 873
rect 1436 847 1443 1153
rect 1456 1147 1463 1183
rect 1496 1180 1503 1183
rect 1493 1167 1507 1180
rect 1476 1156 1493 1163
rect 1476 987 1483 1156
rect 1496 1107 1503 1132
rect 1536 1067 1543 1233
rect 1556 1227 1563 1293
rect 1736 1287 1743 1434
rect 1573 1167 1587 1172
rect 1616 1167 1623 1183
rect 1547 1056 1563 1063
rect 1496 916 1503 1033
rect 1516 967 1523 1053
rect 1533 920 1547 933
rect 1556 927 1563 1056
rect 1536 916 1543 920
rect 1476 880 1483 883
rect 1473 867 1487 880
rect 1576 847 1583 1113
rect 1616 967 1623 1153
rect 1636 943 1643 1133
rect 1656 1127 1663 1214
rect 1676 1167 1683 1253
rect 1756 1216 1763 1293
rect 1627 936 1643 943
rect 1616 916 1623 932
rect 1676 916 1683 973
rect 1596 886 1603 913
rect 1376 663 1383 694
rect 1336 647 1343 663
rect 1356 656 1383 663
rect 1396 663 1403 733
rect 1416 707 1423 753
rect 1476 696 1483 753
rect 1516 707 1523 813
rect 1396 656 1423 663
rect 1276 447 1283 573
rect 1336 527 1343 633
rect 1173 407 1187 413
rect 1196 396 1243 403
rect 1276 396 1283 433
rect 756 123 763 143
rect 736 116 763 123
rect 736 107 743 116
rect 816 107 823 193
rect 856 176 863 233
rect 896 176 903 253
rect 1036 227 1043 253
rect 993 180 1007 193
rect 996 176 1003 180
rect 1036 176 1043 213
rect 1116 187 1123 363
rect 1156 203 1163 253
rect 1136 196 1163 203
rect 1136 176 1143 196
rect 1176 187 1183 313
rect 1096 146 1103 173
rect 1196 147 1203 396
rect 1256 360 1263 363
rect 1253 347 1267 360
rect 1316 227 1323 273
rect 1336 267 1343 413
rect 1356 407 1363 656
rect 1373 400 1387 413
rect 1416 408 1423 656
rect 1496 567 1503 613
rect 1516 567 1523 653
rect 1536 427 1543 833
rect 1576 807 1583 833
rect 1696 807 1703 1172
rect 1716 1067 1723 1183
rect 1716 767 1723 953
rect 1747 923 1760 927
rect 1747 916 1763 923
rect 1747 913 1760 916
rect 1776 847 1783 883
rect 1776 767 1783 833
rect 1576 696 1583 733
rect 1616 696 1623 733
rect 1656 587 1663 653
rect 1676 607 1683 753
rect 1707 703 1720 707
rect 1707 696 1723 703
rect 1756 696 1763 733
rect 1776 727 1783 753
rect 1796 707 1803 773
rect 1707 693 1720 696
rect 1736 643 1743 652
rect 1716 636 1743 643
rect 1676 507 1683 593
rect 1716 587 1723 636
rect 1736 547 1743 613
rect 1596 447 1603 493
rect 1376 396 1383 400
rect 1553 400 1567 413
rect 1556 396 1563 400
rect 1396 267 1403 352
rect 1416 287 1423 313
rect 1436 307 1443 352
rect 1456 283 1463 353
rect 1436 276 1463 283
rect 1236 176 1243 213
rect 1273 180 1287 193
rect 1276 176 1283 180
rect 1336 147 1343 213
rect 1356 187 1363 253
rect 1436 227 1443 276
rect 1376 176 1383 213
rect 1456 183 1463 233
rect 1476 207 1483 393
rect 1580 363 1593 367
rect 1496 287 1503 313
rect 1536 267 1543 363
rect 1576 356 1593 363
rect 1580 353 1593 356
rect 1616 327 1623 473
rect 1673 400 1687 413
rect 1676 396 1683 400
rect 1756 363 1763 633
rect 1796 587 1803 653
rect 1816 623 1823 1353
rect 1836 1167 1843 1392
rect 1876 1367 1883 1653
rect 1896 1627 1903 1703
rect 1916 1667 1923 1893
rect 1956 1827 1963 1923
rect 2016 1747 2023 2193
rect 2036 2067 2043 2216
rect 2036 1927 2043 2032
rect 1896 1347 1903 1613
rect 1916 1436 1923 1473
rect 1936 1467 1943 1734
rect 1976 1687 1983 1703
rect 1976 1587 1983 1673
rect 1916 1256 1923 1373
rect 1956 1367 1963 1403
rect 1956 1307 1963 1353
rect 1976 1223 1983 1473
rect 1996 1387 2003 1653
rect 2016 1627 2023 1693
rect 2036 1527 2043 1793
rect 2056 1667 2063 2436
rect 2076 2387 2083 2443
rect 2116 2440 2123 2443
rect 2113 2427 2127 2440
rect 2187 2436 2203 2443
rect 2076 2267 2083 2313
rect 2096 2287 2103 2353
rect 2136 2220 2143 2223
rect 2096 2187 2103 2212
rect 2133 2207 2147 2220
rect 2176 2207 2183 2373
rect 2196 2226 2203 2436
rect 2236 2256 2243 2413
rect 2336 2387 2343 2613
rect 2456 2476 2463 2653
rect 2356 2447 2363 2474
rect 2496 2387 2503 2573
rect 2616 2527 2623 2713
rect 2676 2707 2683 2743
rect 2756 2527 2763 2913
rect 2956 2887 2963 2963
rect 2956 2807 2963 2873
rect 2776 2746 2783 2773
rect 2896 2746 2903 2773
rect 2816 2740 2823 2743
rect 2813 2727 2827 2740
rect 2916 2547 2923 2793
rect 2976 2776 2983 2813
rect 2996 2787 3003 2993
rect 3156 2967 3163 2994
rect 3096 2927 3103 2963
rect 3007 2776 3023 2783
rect 2936 2627 2943 2743
rect 3096 2707 3103 2913
rect 3216 2787 3223 2963
rect 3256 2927 3263 2963
rect 3296 2803 3303 3193
rect 3316 2947 3323 3113
rect 3396 3047 3403 3313
rect 3436 3227 3443 3263
rect 3380 3026 3400 3027
rect 3380 3023 3393 3026
rect 3376 3013 3393 3023
rect 3376 2996 3383 3013
rect 3356 2947 3363 2963
rect 3276 2796 3303 2803
rect 3276 2746 3283 2796
rect 3336 2776 3343 2813
rect 3356 2783 3363 2933
rect 3356 2776 3383 2783
rect 3196 2647 3203 2732
rect 2913 2527 2927 2533
rect 2516 2407 2523 2474
rect 2656 2446 2663 2513
rect 2696 2476 2703 2513
rect 2856 2476 2863 2513
rect 2976 2507 2983 2533
rect 2976 2476 2983 2493
rect 3036 2476 3043 2633
rect 3136 2527 3143 2573
rect 2716 2407 2723 2443
rect 2276 2256 2283 2313
rect 2336 2247 2343 2333
rect 2376 2256 2383 2373
rect 2416 2256 2423 2293
rect 2576 2267 2583 2373
rect 2596 2268 2603 2353
rect 2776 2307 2783 2473
rect 2956 2440 2963 2443
rect 2176 2147 2183 2193
rect 2076 1956 2083 1993
rect 2116 1983 2123 2113
rect 2136 2047 2143 2073
rect 2196 2047 2203 2212
rect 2256 2167 2263 2223
rect 2267 2156 2283 2163
rect 2116 1976 2143 1983
rect 2116 1807 2123 1923
rect 2136 1787 2143 1976
rect 2156 1748 2163 2013
rect 2196 1956 2203 2012
rect 2236 1956 2243 2033
rect 2076 1587 2083 1703
rect 2156 1687 2163 1734
rect 2176 1707 2183 1773
rect 2216 1743 2223 1912
rect 2196 1736 2223 1743
rect 2236 1736 2243 1853
rect 2276 1803 2283 2156
rect 2296 1967 2303 2223
rect 2476 2226 2483 2253
rect 2316 1956 2323 2213
rect 2356 1956 2363 2213
rect 2396 2087 2403 2223
rect 2256 1796 2283 1803
rect 2256 1767 2263 1796
rect 2276 1736 2283 1773
rect 2316 1747 2323 1893
rect 2336 1867 2343 1923
rect 2416 1926 2423 2133
rect 2436 1967 2443 2173
rect 2516 2147 2523 2223
rect 2556 2187 2563 2212
rect 2556 2087 2563 2113
rect 2456 1956 2463 2033
rect 2596 1956 2603 2173
rect 2656 1987 2663 2253
rect 2676 2226 2683 2293
rect 2036 1436 2043 1492
rect 2116 1447 2123 1553
rect 1956 1216 1983 1223
rect 1856 916 1863 973
rect 1896 916 1903 1113
rect 2016 1087 2023 1393
rect 2056 1327 2063 1403
rect 2096 1396 2123 1403
rect 2096 1247 2103 1313
rect 2116 1307 2123 1396
rect 2136 1347 2143 1453
rect 2176 1436 2183 1613
rect 2196 1467 2203 1736
rect 2256 1467 2263 1671
rect 2053 1220 2067 1233
rect 2056 1216 2063 1220
rect 1936 886 1943 973
rect 2036 967 2043 1183
rect 2096 1180 2103 1183
rect 2093 1167 2107 1180
rect 2087 1083 2100 1087
rect 2087 1073 2103 1083
rect 1836 647 1843 793
rect 1856 707 1863 853
rect 1876 787 1883 883
rect 2076 883 2083 1033
rect 2096 967 2103 1073
rect 2116 1027 2123 1253
rect 2156 1227 2163 1393
rect 2196 1267 2203 1403
rect 2236 1347 2243 1403
rect 2136 1183 2143 1214
rect 2236 1227 2243 1312
rect 2276 1263 2283 1453
rect 2296 1447 2303 1671
rect 2336 1467 2343 1753
rect 2356 1747 2363 1793
rect 2396 1783 2403 1913
rect 2376 1780 2403 1783
rect 2373 1776 2403 1780
rect 2373 1767 2387 1776
rect 2436 1747 2443 1853
rect 2476 1827 2483 1923
rect 2536 1847 2543 1954
rect 2616 1887 2623 1923
rect 2516 1748 2523 1813
rect 2576 1747 2583 1873
rect 2616 1736 2623 1773
rect 2676 1767 2683 2153
rect 2696 1947 2703 2033
rect 2736 2007 2743 2133
rect 2776 2107 2783 2223
rect 2816 2187 2823 2273
rect 2736 1956 2743 1993
rect 2776 1968 2783 2013
rect 2796 1747 2803 1853
rect 2816 1807 2823 2173
rect 2796 1736 2813 1747
rect 2800 1733 2813 1736
rect 2356 1696 2383 1703
rect 2356 1647 2363 1696
rect 2356 1607 2363 1633
rect 2313 1440 2327 1453
rect 2376 1443 2383 1673
rect 2316 1436 2323 1440
rect 2356 1436 2383 1443
rect 2336 1267 2343 1392
rect 2396 1307 2403 1473
rect 2416 1327 2423 1513
rect 2436 1447 2443 1693
rect 2456 1463 2463 1733
rect 2496 1467 2503 1703
rect 2556 1567 2563 1733
rect 2456 1456 2483 1463
rect 2476 1436 2483 1456
rect 2576 1447 2583 1693
rect 2636 1667 2643 1703
rect 2656 1467 2663 1673
rect 2696 1667 2703 1733
rect 2736 1667 2743 1703
rect 2256 1256 2283 1263
rect 2136 1176 2163 1183
rect 2176 1180 2183 1183
rect 2136 1027 2143 1113
rect 2156 947 2163 1176
rect 2173 1167 2187 1180
rect 2216 1147 2223 1172
rect 2176 1007 2183 1132
rect 2236 1127 2243 1173
rect 1876 696 1883 752
rect 1936 747 1943 872
rect 2036 807 2043 883
rect 2076 876 2123 883
rect 1956 707 1963 773
rect 1816 616 1843 623
rect 1816 467 1823 593
rect 1836 407 1843 616
rect 1856 587 1863 653
rect 1896 627 1903 663
rect 1976 666 1983 753
rect 2007 703 2020 707
rect 2007 696 2023 703
rect 2053 700 2067 713
rect 2096 707 2103 876
rect 2056 696 2063 700
rect 2007 693 2020 696
rect 1876 567 1883 593
rect 1956 527 1963 653
rect 2076 660 2083 663
rect 2073 647 2087 660
rect 1656 327 1663 363
rect 1696 327 1703 363
rect 1736 356 1763 363
rect 1456 176 1503 183
rect 916 140 923 143
rect 1016 140 1023 143
rect 913 127 927 140
rect 1013 127 1027 140
rect 727 96 743 107
rect 727 93 740 96
rect 1436 47 1443 113
rect 1476 47 1483 176
rect 1616 146 1623 193
rect 1596 136 1613 143
rect 1636 87 1643 233
rect 1736 176 1743 356
rect 1856 366 1863 433
rect 1896 396 1903 493
rect 2116 487 2123 853
rect 2136 707 2143 793
rect 2156 767 2163 883
rect 2176 727 2183 873
rect 2196 827 2203 1113
rect 2236 928 2243 1033
rect 2256 947 2263 1256
rect 2273 1228 2287 1233
rect 2296 1216 2303 1253
rect 2356 1247 2363 1293
rect 2356 1180 2363 1183
rect 2353 1167 2367 1180
rect 2416 1167 2423 1273
rect 2436 1216 2443 1393
rect 2456 1287 2463 1403
rect 2476 1267 2483 1353
rect 2536 1347 2543 1393
rect 2556 1367 2563 1434
rect 2633 1440 2647 1453
rect 2676 1447 2683 1493
rect 2636 1436 2643 1440
rect 2573 1383 2587 1393
rect 2573 1380 2603 1383
rect 2576 1376 2603 1380
rect 2353 1147 2367 1153
rect 2300 1103 2313 1107
rect 2296 1093 2313 1103
rect 2296 927 2303 1093
rect 2280 923 2293 927
rect 2276 916 2293 923
rect 2280 913 2293 916
rect 2256 863 2263 883
rect 2236 856 2263 863
rect 2176 696 2183 713
rect 2216 696 2223 793
rect 2236 727 2243 856
rect 2256 707 2263 833
rect 2156 660 2163 663
rect 2136 567 2143 653
rect 2153 647 2167 660
rect 2196 627 2203 663
rect 2276 647 2283 853
rect 2296 703 2303 813
rect 2316 728 2323 1053
rect 2336 1027 2343 1073
rect 2356 1047 2363 1112
rect 2476 1067 2483 1183
rect 2496 1047 2503 1293
rect 2516 1287 2523 1313
rect 2596 1216 2603 1376
rect 2616 1347 2623 1403
rect 2696 1403 2703 1593
rect 2716 1527 2723 1573
rect 2756 1463 2763 1633
rect 2776 1467 2783 1703
rect 2796 1507 2803 1673
rect 2816 1627 2823 1693
rect 2747 1456 2763 1463
rect 2736 1436 2743 1453
rect 2780 1443 2793 1447
rect 2776 1436 2793 1443
rect 2780 1433 2793 1436
rect 2676 1396 2703 1403
rect 2436 1040 2483 1043
rect 2436 1036 2487 1040
rect 2336 927 2343 992
rect 2356 916 2363 1012
rect 2393 967 2407 973
rect 2416 927 2423 973
rect 2436 907 2443 1036
rect 2473 1027 2487 1036
rect 2456 987 2463 1013
rect 2516 967 2523 1053
rect 2487 953 2493 967
rect 2516 916 2523 953
rect 2556 927 2563 1183
rect 2576 886 2583 933
rect 2596 923 2603 1113
rect 2616 947 2623 1253
rect 2656 1243 2663 1392
rect 2676 1287 2683 1396
rect 2756 1367 2763 1403
rect 2796 1347 2803 1393
rect 2636 1236 2663 1243
rect 2636 1167 2643 1236
rect 2676 1223 2683 1273
rect 2696 1247 2703 1273
rect 2656 1216 2683 1223
rect 2656 943 2663 1216
rect 2696 1027 2703 1153
rect 2716 987 2723 1183
rect 2736 1027 2743 1053
rect 2656 936 2683 943
rect 2596 916 2623 923
rect 2336 847 2343 873
rect 2496 880 2503 883
rect 2296 696 2313 703
rect 2356 703 2363 853
rect 2376 767 2383 872
rect 2433 867 2447 872
rect 2493 867 2507 880
rect 2596 867 2603 916
rect 2676 887 2683 936
rect 2713 927 2727 933
rect 2736 916 2743 1013
rect 2756 947 2763 1332
rect 2796 1223 2803 1293
rect 2816 1267 2823 1553
rect 2836 1447 2843 2293
rect 2876 2256 2883 2333
rect 2896 2287 2903 2433
rect 2953 2427 2967 2440
rect 2996 2347 3003 2443
rect 3136 2427 3143 2473
rect 2996 2227 3003 2333
rect 3136 2267 3143 2333
rect 3156 2307 3163 2593
rect 3276 2447 3283 2732
rect 3296 2707 3303 2743
rect 3436 2707 3443 3173
rect 3476 3127 3483 3263
rect 3556 3187 3563 3413
rect 3596 3367 3603 3483
rect 3656 3427 3663 3553
rect 3716 3516 3723 3553
rect 3476 3087 3483 3113
rect 3513 3000 3527 3013
rect 3516 2996 3523 3000
rect 3496 2960 3503 2963
rect 3493 2947 3507 2960
rect 3536 2867 3543 2963
rect 3576 2947 3583 3333
rect 3596 3207 3603 3263
rect 3456 2746 3463 2853
rect 3596 2723 3603 3153
rect 3576 2716 3603 2723
rect 3476 2607 3483 2693
rect 3316 2476 3323 2513
rect 3476 2507 3483 2593
rect 3353 2480 3367 2493
rect 3356 2476 3363 2480
rect 3473 2480 3487 2493
rect 3516 2487 3523 2513
rect 3476 2476 3483 2480
rect 3216 2347 3223 2443
rect 3336 2440 3343 2443
rect 2896 2167 2903 2223
rect 2916 2087 2923 2213
rect 3016 2167 3023 2253
rect 3036 2216 3063 2223
rect 3116 2220 3123 2223
rect 3036 2167 3043 2216
rect 3113 2207 3127 2220
rect 3116 2107 3123 2193
rect 3136 2087 3143 2213
rect 3236 2207 3243 2433
rect 3333 2427 3347 2440
rect 3396 2427 3403 2474
rect 3456 2407 3463 2443
rect 3513 2423 3527 2433
rect 3496 2420 3527 2423
rect 3496 2416 3523 2420
rect 2916 2043 2923 2073
rect 2907 2036 2923 2043
rect 2896 1956 2903 2033
rect 2956 2016 2973 2023
rect 2856 1767 2863 1833
rect 2916 1827 2923 1913
rect 2936 1767 2943 1933
rect 2956 1847 2963 2016
rect 2973 2003 2987 2013
rect 2973 2000 3003 2003
rect 2976 1996 3003 2000
rect 2973 1967 2987 1973
rect 2996 1956 3003 1996
rect 3033 1968 3047 1973
rect 3046 1960 3047 1968
rect 3056 1967 3063 2053
rect 3156 2047 3163 2093
rect 3236 2043 3243 2193
rect 3256 2047 3263 2333
rect 3376 2267 3383 2393
rect 3276 2143 3283 2213
rect 3356 2187 3363 2223
rect 3396 2207 3403 2293
rect 3416 2223 3423 2373
rect 3496 2256 3503 2416
rect 3516 2327 3523 2393
rect 3536 2267 3543 2653
rect 3556 2387 3563 2693
rect 3576 2487 3583 2716
rect 3616 2707 3623 3033
rect 3636 3008 3643 3294
rect 3676 3266 3683 3313
rect 3696 3127 3703 3483
rect 3716 3347 3723 3413
rect 3736 3307 3743 3472
rect 3756 3303 3763 3393
rect 3776 3367 3783 3553
rect 3833 3520 3847 3533
rect 3836 3516 3843 3520
rect 3816 3407 3823 3483
rect 3756 3296 3783 3303
rect 3856 3266 3863 3433
rect 3896 3407 3903 3773
rect 3936 3647 3943 3783
rect 4016 3627 4023 3653
rect 3953 3520 3967 3533
rect 3956 3516 3963 3520
rect 3936 3447 3943 3483
rect 3976 3480 3983 3483
rect 3973 3467 3987 3480
rect 4016 3307 4023 3473
rect 4036 3467 4043 3593
rect 4056 3527 4063 3633
rect 4076 3567 4083 3853
rect 4136 3847 4143 3933
rect 4196 3847 4203 4013
rect 4296 4006 4303 4073
rect 4096 3786 4103 3833
rect 4096 3516 4103 3713
rect 4116 3667 4123 3733
rect 4196 3687 4203 3772
rect 4216 3687 4223 3733
rect 4236 3727 4243 3913
rect 4156 3523 4163 3593
rect 4176 3587 4183 3633
rect 4196 3607 4203 3673
rect 4236 3607 4243 3713
rect 4256 3707 4263 3933
rect 4316 3847 4323 4133
rect 4356 4036 4363 4073
rect 4436 4007 4443 4053
rect 4476 4036 4483 4093
rect 4496 4067 4503 4113
rect 4576 4107 4583 4296
rect 4596 4187 4603 4453
rect 4636 4423 4643 4733
rect 4916 4707 4923 4933
rect 4936 4907 4943 5033
rect 5056 4967 5063 5043
rect 5276 5046 5283 5073
rect 5187 5036 5203 5043
rect 4996 4856 5003 4913
rect 4936 4807 4943 4853
rect 5056 4787 5063 4893
rect 5136 4856 5143 4893
rect 5176 4827 5183 5033
rect 5236 4856 5243 4973
rect 5216 4787 5223 4823
rect 4856 4567 4863 4633
rect 4756 4526 4763 4553
rect 4676 4520 4683 4523
rect 4673 4507 4687 4520
rect 4676 4427 4683 4493
rect 4616 4416 4643 4423
rect 4616 4306 4623 4416
rect 4676 4336 4683 4373
rect 4796 4348 4803 4523
rect 4836 4427 4843 4523
rect 4876 4467 4883 4693
rect 4896 4567 4903 4593
rect 4936 4556 4943 4593
rect 4907 4523 4920 4527
rect 4907 4516 4923 4523
rect 4907 4513 4920 4516
rect 4956 4507 4963 4523
rect 4836 4387 4843 4413
rect 4956 4367 4963 4493
rect 4916 4336 4963 4343
rect 4516 4048 4523 4073
rect 4636 4036 4643 4153
rect 4696 4147 4703 4273
rect 4776 4167 4783 4292
rect 4836 4143 4843 4333
rect 4956 4307 4963 4336
rect 4936 4296 4953 4303
rect 4816 4136 4843 4143
rect 4696 4036 4703 4133
rect 4496 3967 4503 4003
rect 4556 3967 4563 4034
rect 4656 4000 4663 4003
rect 4653 3987 4667 4000
rect 4276 3787 4283 3833
rect 4516 3816 4543 3823
rect 4156 3516 4183 3523
rect 4233 3520 4247 3533
rect 4236 3516 4243 3520
rect 4276 3487 4283 3533
rect 4076 3427 4083 3483
rect 4096 3336 4103 3453
rect 4296 3447 4303 3753
rect 4316 3687 4323 3783
rect 4336 3767 4343 3813
rect 4416 3776 4433 3783
rect 4396 3487 4403 3514
rect 4296 3336 4303 3393
rect 4416 3347 4423 3776
rect 4496 3727 4503 3773
rect 4516 3647 4523 3816
rect 4576 3747 4583 3783
rect 4596 3567 4603 3973
rect 4796 3967 4803 4093
rect 4816 4006 4823 4136
rect 4916 3927 4923 4273
rect 4936 4006 4943 4296
rect 4976 4227 4983 4453
rect 4996 4347 5003 4513
rect 5016 4487 5023 4773
rect 5036 4526 5043 4593
rect 5136 4567 5143 4673
rect 5156 4556 5163 4733
rect 5076 4503 5083 4523
rect 5076 4496 5103 4503
rect 5036 4336 5043 4413
rect 4996 4036 5003 4073
rect 5076 4067 5083 4473
rect 5096 4427 5103 4496
rect 5173 4347 5187 4353
rect 5116 4187 5123 4303
rect 5196 4287 5203 4433
rect 5216 4347 5223 4473
rect 5256 4447 5263 4554
rect 5276 4526 5283 4973
rect 5316 4927 5323 5043
rect 5356 4987 5363 5043
rect 5396 4967 5403 5074
rect 5636 5043 5643 5332
rect 5716 5127 5723 5343
rect 5436 5007 5443 5043
rect 5476 5007 5483 5043
rect 5616 5036 5643 5043
rect 5316 4856 5323 4913
rect 5436 4816 5463 4823
rect 5376 4747 5383 4812
rect 5456 4727 5463 4816
rect 5376 4427 5383 4533
rect 5396 4336 5403 4713
rect 5476 4707 5483 4953
rect 5496 4827 5503 5013
rect 5556 4856 5563 4893
rect 5616 4827 5623 5036
rect 5656 5007 5663 5073
rect 5716 4927 5723 5043
rect 5707 4906 5720 4907
rect 5707 4893 5713 4906
rect 5756 4903 5763 5113
rect 5736 4896 5763 4903
rect 5713 4867 5727 4872
rect 5636 4816 5663 4823
rect 5436 4487 5443 4512
rect 5436 4427 5443 4473
rect 5476 4467 5483 4523
rect 5516 4447 5523 4693
rect 5576 4556 5583 4593
rect 5556 4487 5563 4523
rect 5436 4336 5443 4373
rect 5556 4347 5563 4433
rect 5227 4303 5240 4307
rect 5227 4296 5243 4303
rect 5227 4293 5240 4296
rect 5113 4040 5127 4053
rect 5116 4036 5123 4040
rect 5156 4036 5163 4271
rect 5176 4067 5183 4173
rect 5193 4040 5207 4053
rect 5196 4036 5203 4040
rect 5016 3967 5023 4003
rect 4653 3820 4667 3833
rect 4656 3816 4663 3820
rect 4856 3827 4863 3913
rect 5076 3907 5083 4032
rect 4613 3807 4627 3813
rect 4756 3786 4763 3813
rect 4616 3607 4623 3772
rect 4636 3707 4643 3773
rect 4796 3780 4803 3783
rect 4836 3780 4843 3783
rect 4673 3767 4687 3772
rect 4793 3767 4807 3780
rect 4833 3767 4847 3780
rect 4856 3667 4863 3773
rect 4876 3727 4883 3783
rect 4936 3776 4963 3783
rect 4956 3707 4963 3776
rect 4976 3767 4983 3814
rect 4996 3683 5003 3893
rect 5076 3707 5083 3753
rect 4996 3676 5023 3683
rect 4496 3516 4503 3553
rect 4616 3516 4623 3593
rect 4476 3447 4483 3483
rect 4676 3483 4683 3633
rect 4736 3567 4743 3593
rect 4736 3516 4743 3553
rect 4676 3476 4703 3483
rect 4036 3296 4063 3303
rect 3776 2996 3783 3033
rect 3876 2967 3883 3213
rect 4036 3087 4043 3296
rect 4196 3266 4203 3333
rect 4616 3308 4623 3393
rect 4676 3308 4683 3333
rect 4156 3256 4183 3263
rect 4176 3127 4183 3256
rect 4216 3256 4243 3263
rect 4216 3167 4223 3256
rect 3936 2996 3943 3073
rect 4016 3008 4023 3033
rect 3676 2827 3683 2963
rect 3696 2776 3703 2813
rect 3656 2547 3663 2743
rect 3596 2476 3603 2533
rect 3656 2483 3663 2533
rect 3676 2527 3683 2693
rect 3796 2667 3803 2963
rect 3916 2927 3923 2963
rect 3956 2887 3963 2963
rect 4016 2927 4023 2994
rect 4116 2967 4123 3113
rect 4216 2996 4223 3153
rect 4336 2996 4343 3033
rect 4056 2927 4063 2963
rect 3816 2747 3823 2813
rect 3716 2488 3723 2553
rect 3756 2507 3763 2593
rect 3656 2476 3683 2483
rect 3416 2216 3443 2223
rect 3476 2220 3483 2223
rect 3276 2136 3303 2143
rect 3216 2036 3243 2043
rect 3076 1926 3083 1993
rect 3096 1987 3103 2013
rect 3176 1956 3183 2033
rect 3216 1956 3223 2036
rect 3296 1967 3303 2136
rect 3416 2127 3423 2193
rect 2856 1687 2863 1732
rect 2876 1700 2883 1703
rect 2873 1687 2887 1700
rect 2876 1647 2883 1673
rect 2856 1436 2863 1513
rect 2876 1467 2883 1493
rect 2896 1448 2903 1673
rect 2936 1667 2943 1703
rect 2936 1587 2943 1632
rect 2956 1567 2963 1793
rect 2976 1607 2983 1913
rect 3016 1763 3023 1923
rect 3156 1920 3163 1923
rect 3153 1907 3167 1920
rect 3056 1827 3063 1853
rect 3016 1756 3043 1763
rect 3036 1748 3043 1756
rect 3156 1736 3163 1872
rect 3196 1827 3203 1913
rect 3196 1748 3203 1813
rect 2996 1507 3003 1673
rect 2836 1247 2843 1393
rect 2776 1216 2803 1223
rect 2776 923 2783 1216
rect 2856 1183 2863 1214
rect 2876 1207 2883 1392
rect 2936 1243 2943 1473
rect 2996 1463 3003 1493
rect 3016 1487 3023 1703
rect 3036 1487 3043 1533
rect 3056 1527 3063 1553
rect 2996 1456 3023 1463
rect 3016 1436 3023 1456
rect 2996 1323 3003 1403
rect 2976 1316 3003 1323
rect 2976 1287 2983 1316
rect 2936 1240 2983 1243
rect 2936 1236 2987 1240
rect 2973 1227 2987 1236
rect 2996 1186 3003 1293
rect 2836 1103 2843 1183
rect 2856 1176 2883 1183
rect 2836 1096 2863 1103
rect 2836 1007 2843 1073
rect 2856 1067 2863 1096
rect 2876 1087 2883 1176
rect 2776 916 2803 923
rect 2656 847 2663 883
rect 2356 696 2383 703
rect 2416 696 2423 753
rect 2187 616 2203 627
rect 2213 627 2227 633
rect 2187 613 2200 616
rect 1836 307 1843 353
rect 1656 127 1663 174
rect 1796 167 1803 293
rect 1956 267 1963 363
rect 1853 180 1867 193
rect 1976 188 1983 333
rect 2016 307 2023 453
rect 2113 400 2127 413
rect 2116 396 2123 400
rect 2156 366 2163 493
rect 2196 408 2203 473
rect 2236 427 2243 453
rect 2233 400 2247 413
rect 2276 407 2283 612
rect 2296 547 2303 653
rect 2236 396 2243 400
rect 2316 407 2323 473
rect 2336 467 2343 663
rect 2376 627 2383 696
rect 2496 707 2503 753
rect 2413 603 2427 613
rect 2436 607 2443 663
rect 2476 660 2483 663
rect 2473 647 2487 660
rect 2387 600 2427 603
rect 2387 596 2423 600
rect 2456 587 2463 613
rect 2376 503 2383 553
rect 2396 527 2403 573
rect 2376 496 2403 503
rect 2356 427 2363 493
rect 2056 360 2063 363
rect 2053 347 2067 360
rect 2216 360 2223 363
rect 1856 176 1863 180
rect 2016 176 2023 213
rect 1916 146 1923 173
rect 2056 146 2063 233
rect 2136 176 2143 293
rect 2176 187 2183 353
rect 2213 347 2227 360
rect 2256 223 2263 363
rect 2296 327 2303 394
rect 2376 396 2383 473
rect 2396 447 2403 496
rect 2416 407 2423 533
rect 2316 307 2323 353
rect 2396 327 2403 363
rect 2436 363 2443 553
rect 2496 547 2503 653
rect 2516 607 2523 793
rect 2576 708 2583 753
rect 2676 707 2683 852
rect 2696 783 2703 913
rect 2756 880 2763 883
rect 2753 867 2767 880
rect 2696 776 2723 783
rect 2616 696 2663 703
rect 2456 447 2463 493
rect 2536 487 2543 653
rect 2556 607 2563 663
rect 2593 647 2607 652
rect 2496 396 2503 473
rect 2536 396 2543 433
rect 2556 407 2563 533
rect 2436 356 2483 363
rect 2416 287 2423 353
rect 2436 327 2443 356
rect 2476 307 2483 333
rect 2516 287 2523 363
rect 2576 307 2583 433
rect 2636 396 2643 433
rect 2656 423 2663 696
rect 2696 696 2703 753
rect 2716 727 2723 776
rect 2736 696 2743 753
rect 2776 707 2783 873
rect 2796 847 2803 916
rect 2796 783 2803 833
rect 2816 827 2823 973
rect 2836 916 2843 993
rect 2896 967 2903 1113
rect 2916 1107 2923 1183
rect 3016 1163 3023 1333
rect 3036 1267 3043 1392
rect 3076 1347 3083 1734
rect 3093 1682 3107 1693
rect 3176 1700 3183 1703
rect 3173 1687 3187 1700
rect 3093 1680 3133 1682
rect 3096 1675 3133 1680
rect 3196 1667 3203 1692
rect 3096 1447 3103 1593
rect 3116 1587 3123 1633
rect 3116 1487 3123 1513
rect 3156 1436 3163 1473
rect 3076 1216 3083 1293
rect 3096 1287 3103 1393
rect 3136 1383 3143 1403
rect 3136 1376 3163 1383
rect 3116 1187 3123 1253
rect 3036 1163 3043 1183
rect 3016 1156 3043 1163
rect 2896 953 2913 967
rect 2896 916 2903 953
rect 2856 880 2863 883
rect 2853 867 2867 880
rect 2796 776 2823 783
rect 2796 687 2803 753
rect 2816 707 2823 776
rect 2836 747 2843 813
rect 2916 767 2923 914
rect 2936 807 2943 1073
rect 2956 1027 2963 1113
rect 3016 1107 3023 1156
rect 3066 1153 3067 1160
rect 3053 1143 3067 1153
rect 3036 1140 3067 1143
rect 3036 1136 3063 1140
rect 3036 1067 3043 1136
rect 2996 947 3003 993
rect 3016 916 3023 1013
rect 3036 1007 3043 1032
rect 3056 987 3063 1073
rect 2996 827 3003 883
rect 2976 776 3023 783
rect 2976 747 2983 776
rect 2996 708 3003 753
rect 3016 747 3023 776
rect 2900 703 2913 707
rect 2896 696 2913 703
rect 2900 693 2913 696
rect 3056 707 3063 873
rect 2676 447 2683 653
rect 2656 416 2683 423
rect 2676 408 2683 416
rect 2696 407 2703 633
rect 2716 507 2723 663
rect 2756 627 2763 663
rect 2776 487 2783 653
rect 2816 487 2823 653
rect 2916 527 2923 652
rect 2936 627 2943 694
rect 2956 507 2963 633
rect 2976 627 2983 663
rect 3053 647 3067 653
rect 3016 607 3023 631
rect 3016 507 3023 572
rect 2616 360 2623 363
rect 2296 247 2303 273
rect 2296 236 2313 247
rect 2300 233 2313 236
rect 2256 220 2283 223
rect 2256 216 2287 220
rect 2196 146 2203 213
rect 2273 207 2287 216
rect 2266 193 2267 200
rect 2213 187 2227 193
rect 2253 180 2267 193
rect 2256 176 2263 180
rect 1656 67 1663 113
rect 1836 107 1843 143
rect 1956 107 1963 132
rect 1996 47 2003 143
rect 2116 140 2123 143
rect 2113 127 2127 140
rect 2136 67 2143 93
rect 2196 67 2203 132
rect 2236 107 2243 143
rect 2336 27 2343 273
rect 2536 263 2543 293
rect 2507 256 2543 263
rect 2367 233 2373 247
rect 2376 47 2383 113
rect 2396 107 2403 143
rect 2476 127 2483 233
rect 2516 176 2523 213
rect 2556 188 2563 233
rect 2596 187 2603 353
rect 2613 347 2627 360
rect 2656 343 2663 363
rect 2636 336 2663 343
rect 2533 127 2547 132
rect 2513 107 2527 113
rect 2576 107 2583 132
rect 2616 127 2623 273
rect 2636 267 2643 336
rect 2676 303 2683 333
rect 2656 296 2683 303
rect 2656 207 2663 296
rect 2676 176 2683 273
rect 2696 207 2703 353
rect 2716 347 2723 472
rect 2793 427 2807 433
rect 2773 400 2787 413
rect 2953 408 2967 413
rect 2776 396 2783 400
rect 2976 407 2983 453
rect 2736 307 2743 353
rect 2756 247 2763 363
rect 2796 327 2803 363
rect 2756 187 2763 233
rect 2813 188 2827 193
rect 2720 183 2733 187
rect 2716 176 2733 183
rect 2720 173 2733 176
rect 2836 183 2843 353
rect 2856 327 2863 394
rect 2896 243 2903 363
rect 2936 307 2943 363
rect 2876 236 2903 243
rect 2876 187 2883 236
rect 2836 176 2863 183
rect 2696 140 2703 143
rect 2693 127 2707 140
rect 2513 106 2540 107
rect 2513 100 2533 106
rect 2516 96 2533 100
rect 2520 93 2533 96
rect 2620 106 2633 107
rect 2627 93 2633 106
rect 2456 -24 2463 13
rect 2536 -24 2543 33
rect 2656 27 2663 111
rect 2676 63 2683 93
rect 2676 56 2703 63
rect 2696 43 2703 56
rect 2736 47 2743 133
rect 2756 107 2763 152
rect 2796 140 2803 143
rect 2793 127 2807 140
rect 2696 36 2723 43
rect 2576 -24 2583 13
rect 2676 -17 2683 33
rect 2716 23 2723 36
rect 2753 23 2767 33
rect 2716 20 2767 23
rect 2716 16 2763 20
rect 2656 -24 2683 -17
rect 2696 -24 2703 13
rect 2856 -17 2863 176
rect 2896 176 2903 213
rect 2936 176 2943 233
rect 2976 227 2983 353
rect 2996 27 3003 473
rect 3036 427 3043 553
rect 3056 396 3063 433
rect 3076 427 3083 1153
rect 3096 987 3103 1183
rect 3136 1167 3143 1353
rect 3156 1227 3163 1376
rect 3176 1307 3183 1403
rect 3216 1367 3223 1833
rect 3236 1747 3243 1813
rect 3276 1763 3283 1873
rect 3296 1787 3303 1913
rect 3316 1763 3323 2093
rect 3336 1827 3343 2113
rect 3396 1887 3403 1923
rect 3436 1847 3443 2216
rect 3473 2207 3487 2220
rect 3516 2187 3523 2212
rect 3556 2167 3563 2273
rect 3576 2267 3583 2413
rect 3616 2307 3623 2443
rect 3676 2307 3683 2476
rect 3756 2476 3763 2493
rect 3776 2487 3783 2573
rect 3607 2283 3620 2287
rect 3607 2273 3623 2283
rect 3616 2256 3623 2273
rect 3676 2263 3683 2293
rect 3656 2256 3703 2263
rect 3756 2256 3763 2333
rect 3796 2267 3803 2593
rect 3896 2507 3903 2613
rect 3916 2547 3923 2732
rect 3893 2480 3907 2493
rect 3936 2487 3943 2713
rect 3956 2667 3963 2774
rect 3976 2727 3983 2913
rect 4196 2887 4203 2963
rect 4256 2887 4263 2994
rect 4376 2967 4383 3294
rect 4416 3167 4423 3263
rect 4436 2996 4443 3233
rect 4516 3207 4523 3293
rect 4616 3143 4623 3294
rect 4716 3267 4723 3413
rect 4756 3387 4763 3573
rect 4776 3447 4783 3514
rect 4916 3487 4923 3553
rect 4996 3527 5003 3653
rect 4816 3427 4823 3483
rect 4976 3447 4983 3483
rect 4773 3300 4787 3313
rect 4776 3296 4783 3300
rect 4816 3296 4823 3373
rect 4656 3260 4663 3263
rect 4653 3247 4667 3260
rect 4693 3247 4707 3253
rect 4756 3227 4763 3263
rect 4833 3247 4847 3252
rect 4856 3227 4863 3433
rect 4873 3307 4887 3313
rect 4896 3296 4903 3393
rect 4996 3383 5003 3473
rect 5016 3467 5023 3676
rect 5076 3567 5083 3633
rect 5076 3516 5083 3553
rect 5096 3547 5103 3772
rect 5116 3747 5123 3973
rect 5176 3867 5183 4003
rect 5236 3927 5243 4053
rect 5256 4043 5263 4113
rect 5276 4107 5283 4303
rect 5316 4267 5323 4333
rect 5356 4227 5363 4273
rect 5256 4036 5283 4043
rect 5356 4047 5363 4213
rect 5340 4003 5353 4007
rect 5336 4000 5353 4003
rect 5333 3993 5353 4000
rect 5376 4003 5383 4303
rect 5416 4300 5423 4303
rect 5413 4287 5427 4300
rect 5576 4303 5583 4453
rect 5407 4256 5433 4263
rect 5456 4047 5463 4293
rect 5476 4147 5483 4303
rect 5536 4300 5543 4303
rect 5533 4287 5547 4300
rect 5556 4296 5583 4303
rect 5407 4043 5420 4047
rect 5407 4036 5423 4043
rect 5407 4034 5420 4036
rect 5400 4033 5420 4034
rect 5476 4036 5483 4133
rect 5533 4040 5547 4053
rect 5556 4047 5563 4296
rect 5536 4036 5543 4040
rect 5376 3996 5403 4003
rect 5333 3987 5347 3993
rect 5116 3667 5123 3733
rect 5136 3603 5143 3814
rect 5236 3783 5243 3853
rect 5216 3776 5243 3783
rect 5256 3783 5263 3873
rect 5356 3816 5363 3913
rect 5376 3827 5383 3973
rect 5256 3776 5303 3783
rect 5127 3596 5143 3603
rect 5116 3516 5123 3593
rect 5056 3480 5063 3483
rect 5053 3467 5067 3480
rect 5133 3463 5147 3473
rect 5116 3460 5147 3463
rect 5116 3456 5143 3460
rect 4996 3376 5023 3383
rect 4933 3300 4947 3313
rect 4936 3296 4943 3300
rect 4956 3260 4963 3263
rect 4953 3247 4967 3260
rect 4616 3136 4643 3143
rect 4536 2996 4543 3073
rect 4616 3003 4623 3033
rect 4596 2996 4623 3003
rect 4007 2816 4043 2823
rect 4036 2803 4043 2816
rect 4376 2807 4383 2833
rect 4036 2796 4063 2803
rect 4013 2780 4027 2793
rect 4016 2776 4023 2780
rect 4056 2776 4063 2796
rect 4076 2740 4083 2743
rect 4036 2627 4043 2732
rect 4073 2727 4087 2740
rect 4116 2727 4123 2773
rect 4056 2667 4063 2713
rect 3896 2476 3903 2480
rect 3816 2447 3823 2474
rect 3956 2476 3963 2533
rect 3876 2440 3883 2443
rect 3833 2423 3847 2433
rect 3816 2420 3847 2423
rect 3873 2427 3887 2440
rect 3916 2436 3933 2443
rect 3816 2416 3843 2420
rect 3696 2226 3703 2256
rect 3456 1927 3463 2073
rect 3276 1756 3303 1763
rect 3316 1760 3343 1763
rect 3316 1756 3347 1760
rect 3296 1736 3303 1756
rect 3333 1747 3347 1756
rect 3236 1447 3243 1693
rect 3276 1607 3283 1703
rect 3336 1647 3343 1693
rect 3356 1667 3363 1793
rect 3376 1507 3383 1773
rect 3416 1736 3423 1773
rect 3476 1723 3483 1973
rect 3496 1956 3503 2093
rect 3536 1907 3543 1923
rect 3576 1907 3583 2213
rect 3636 2220 3643 2223
rect 3633 2207 3647 2220
rect 3596 2027 3603 2113
rect 3616 1967 3623 2053
rect 3696 2003 3703 2133
rect 3736 2067 3743 2173
rect 3727 2053 3743 2067
rect 3736 2047 3743 2053
rect 3636 2000 3703 2003
rect 3633 1996 3703 2000
rect 3633 1987 3647 1996
rect 3653 1960 3667 1973
rect 3700 1963 3713 1967
rect 3656 1956 3663 1960
rect 3696 1956 3713 1963
rect 3700 1953 3713 1956
rect 3596 1903 3603 1953
rect 3596 1896 3623 1903
rect 3536 1767 3543 1893
rect 3573 1867 3587 1872
rect 3576 1807 3583 1853
rect 3556 1736 3563 1793
rect 3596 1736 3603 1873
rect 3616 1867 3623 1896
rect 3476 1716 3503 1723
rect 3296 1436 3303 1473
rect 3116 1047 3123 1133
rect 3176 1087 3183 1183
rect 3216 1163 3223 1183
rect 3196 1156 3223 1163
rect 3107 923 3120 927
rect 3107 916 3123 923
rect 3156 916 3163 1013
rect 3196 967 3203 1156
rect 3236 1047 3243 1133
rect 3256 1047 3263 1373
rect 3276 1327 3283 1403
rect 3356 1406 3363 1473
rect 3396 1436 3403 1692
rect 3456 1647 3463 1703
rect 3476 1406 3483 1693
rect 3496 1687 3503 1716
rect 3516 1696 3543 1703
rect 3576 1700 3583 1703
rect 3516 1448 3523 1696
rect 3573 1687 3587 1700
rect 3556 1507 3563 1553
rect 3576 1467 3583 1533
rect 3573 1440 3587 1453
rect 3576 1436 3583 1440
rect 3596 1406 3603 1573
rect 3316 1307 3323 1393
rect 3336 1267 3343 1333
rect 3376 1216 3383 1253
rect 3276 1186 3283 1213
rect 3276 1147 3283 1172
rect 3333 1147 3347 1153
rect 3327 1140 3347 1147
rect 3327 1136 3343 1140
rect 3327 1133 3340 1136
rect 3356 1087 3363 1183
rect 3396 1083 3403 1173
rect 3376 1076 3403 1083
rect 3216 947 3223 973
rect 3236 923 3243 1033
rect 3256 1007 3263 1033
rect 3216 916 3263 923
rect 3296 916 3303 1013
rect 3336 987 3343 1073
rect 3107 913 3120 916
rect 3136 847 3143 883
rect 3176 847 3183 872
rect 3096 408 3103 833
rect 3116 707 3123 753
rect 3136 696 3143 793
rect 3196 787 3203 873
rect 3216 707 3223 916
rect 3356 927 3363 1033
rect 3116 507 3123 653
rect 3156 607 3163 663
rect 3196 427 3203 652
rect 3216 507 3223 653
rect 3236 527 3243 873
rect 3276 807 3283 883
rect 3276 767 3283 793
rect 3316 767 3323 883
rect 3276 696 3283 732
rect 3356 727 3363 873
rect 3376 767 3383 1076
rect 3396 967 3403 1053
rect 3416 947 3423 1353
rect 3436 1007 3443 1313
rect 3456 1227 3463 1293
rect 3476 1248 3483 1392
rect 3616 1367 3623 1533
rect 3516 1228 3523 1333
rect 3636 1327 3643 1873
rect 3716 1867 3723 1913
rect 3716 1827 3723 1853
rect 3656 1467 3663 1793
rect 3676 1747 3683 1773
rect 3716 1736 3723 1792
rect 3736 1767 3743 1954
rect 3756 1887 3763 2173
rect 3776 2107 3783 2191
rect 3796 2083 3803 2213
rect 3816 2187 3823 2416
rect 3836 2267 3843 2393
rect 3880 2283 3893 2287
rect 3876 2273 3893 2283
rect 3876 2256 3883 2273
rect 3916 2263 3923 2293
rect 3936 2287 3943 2433
rect 4056 2427 4063 2473
rect 4076 2363 4083 2653
rect 4096 2647 4103 2693
rect 4196 2607 4203 2743
rect 4236 2683 4243 2793
rect 4276 2727 4283 2743
rect 4236 2676 4253 2683
rect 4136 2436 4163 2443
rect 4156 2387 4163 2436
rect 4176 2363 4183 2513
rect 4256 2488 4263 2673
rect 4276 2587 4283 2713
rect 4336 2687 4343 2793
rect 4373 2780 4387 2793
rect 4376 2776 4383 2780
rect 4396 2687 4403 2743
rect 4296 2476 4303 2513
rect 4076 2356 4103 2363
rect 3916 2256 3943 2263
rect 3936 2223 3943 2256
rect 3956 2226 3963 2273
rect 4056 2256 4063 2293
rect 3856 2220 3863 2223
rect 3853 2207 3867 2220
rect 3896 2216 3943 2223
rect 4036 2203 4043 2212
rect 4016 2196 4043 2203
rect 3816 2087 3823 2133
rect 3776 2076 3803 2083
rect 3776 1968 3783 2076
rect 3776 1706 3783 1793
rect 3796 1747 3803 1833
rect 3816 1787 3823 1923
rect 3856 1787 3863 2093
rect 3876 1907 3883 2173
rect 3996 2067 4003 2173
rect 3907 1963 3920 1967
rect 3907 1956 3923 1963
rect 3907 1953 3920 1956
rect 3876 1736 3883 1853
rect 3896 1827 3903 1873
rect 3676 1487 3683 1673
rect 3696 1627 3703 1692
rect 3476 928 3483 1153
rect 3496 1147 3503 1183
rect 3576 1167 3583 1313
rect 3616 1247 3623 1293
rect 3676 1216 3683 1313
rect 3716 1243 3723 1653
rect 3736 1427 3743 1692
rect 3756 1543 3763 1693
rect 3856 1700 3863 1703
rect 3853 1687 3867 1700
rect 3836 1587 3843 1613
rect 3856 1607 3863 1673
rect 3896 1547 3903 1693
rect 3916 1667 3923 1893
rect 3936 1767 3943 1923
rect 3996 1787 4003 1953
rect 4016 1843 4023 2196
rect 4036 2007 4043 2133
rect 4056 2087 4063 2193
rect 4096 2147 4103 2356
rect 4156 2356 4183 2363
rect 4156 2256 4163 2356
rect 4196 2267 4203 2293
rect 4136 2220 4143 2223
rect 4056 1956 4063 2073
rect 4096 1987 4103 2112
rect 4116 2007 4123 2213
rect 4133 2207 4147 2220
rect 4093 1960 4107 1973
rect 4096 1956 4103 1960
rect 4036 1863 4043 1913
rect 4036 1856 4063 1863
rect 4016 1836 4043 1843
rect 3940 1746 3960 1747
rect 3947 1743 3960 1746
rect 3947 1736 3963 1743
rect 3947 1733 3960 1736
rect 4036 1747 4043 1836
rect 4016 1700 4023 1703
rect 3936 1647 3943 1673
rect 3756 1536 3773 1543
rect 3776 1436 3783 1533
rect 3836 1436 3843 1533
rect 3736 1267 3743 1413
rect 3796 1327 3803 1392
rect 3716 1236 3743 1243
rect 3736 1207 3743 1236
rect 3796 1216 3803 1253
rect 3396 823 3403 873
rect 3416 847 3423 883
rect 3456 880 3463 883
rect 3453 867 3467 880
rect 3436 827 3443 853
rect 3516 847 3523 1153
rect 3616 1087 3623 1133
rect 3656 967 3663 1183
rect 3696 1067 3703 1183
rect 3736 1067 3743 1172
rect 3756 1087 3763 1173
rect 3696 1027 3703 1053
rect 3533 928 3547 933
rect 3573 928 3587 933
rect 3396 816 3423 823
rect 3213 423 3227 433
rect 3236 423 3243 513
rect 3256 487 3263 653
rect 3336 660 3343 663
rect 3333 647 3347 660
rect 3356 627 3363 653
rect 3376 647 3383 753
rect 3396 707 3403 753
rect 3416 727 3423 816
rect 3436 696 3443 813
rect 3453 707 3467 713
rect 3456 627 3463 653
rect 3213 420 3243 423
rect 3216 416 3243 420
rect 3016 267 3023 353
rect 3096 176 3103 333
rect 3136 327 3143 393
rect 3156 366 3163 413
rect 3216 396 3223 416
rect 3253 400 3267 413
rect 3256 396 3263 400
rect 3160 326 3173 327
rect 3167 313 3173 326
rect 3196 303 3203 363
rect 3236 327 3243 352
rect 3176 296 3203 303
rect 3176 267 3183 296
rect 3296 287 3303 413
rect 3336 360 3343 363
rect 3333 347 3347 360
rect 3396 347 3403 613
rect 3476 607 3483 773
rect 3556 767 3563 883
rect 3576 708 3583 773
rect 3596 767 3603 833
rect 3636 827 3643 873
rect 3656 847 3663 932
rect 3736 916 3743 953
rect 3776 927 3783 993
rect 3616 707 3623 793
rect 3516 660 3523 663
rect 3513 647 3527 660
rect 3436 396 3443 513
rect 3536 367 3543 573
rect 3556 567 3563 663
rect 3596 607 3603 652
rect 3636 587 3643 753
rect 3676 743 3683 873
rect 3696 787 3703 853
rect 3716 767 3723 883
rect 3756 827 3763 883
rect 3676 736 3693 743
rect 3696 696 3703 733
rect 3776 703 3783 873
rect 3796 747 3803 1093
rect 3816 1067 3823 1183
rect 3833 1147 3847 1153
rect 3856 1107 3863 1533
rect 3876 1406 3883 1473
rect 3916 1436 3923 1573
rect 3876 1227 3883 1293
rect 3896 1216 3903 1313
rect 3956 1287 3963 1373
rect 3976 1287 3983 1692
rect 4013 1687 4027 1700
rect 4056 1667 4063 1856
rect 4076 1748 4083 1923
rect 4116 1847 4123 1873
rect 4136 1867 4143 2033
rect 4156 1967 4163 2113
rect 4216 1956 4223 2353
rect 4236 2307 4243 2443
rect 4256 2267 4263 2413
rect 4276 2307 4283 2443
rect 4336 2427 4343 2573
rect 4356 2487 4363 2653
rect 4416 2567 4423 2613
rect 4436 2587 4443 2774
rect 4556 2747 4563 2952
rect 4616 2947 4623 2973
rect 4636 2927 4643 3136
rect 4676 3008 4683 3073
rect 4716 3008 4723 3033
rect 4836 2996 4883 3003
rect 4916 2996 4923 3053
rect 4956 2996 4963 3073
rect 4696 2960 4703 2963
rect 4693 2947 4707 2960
rect 4756 2907 4763 2994
rect 4876 2967 4883 2996
rect 4816 2927 4823 2963
rect 4996 2927 5003 3294
rect 5016 3027 5023 3376
rect 5116 3266 5123 3456
rect 5156 3363 5163 3733
rect 5196 3528 5203 3553
rect 5136 3356 5163 3363
rect 5096 3167 5103 3263
rect 5076 2996 5083 3033
rect 5116 3007 5123 3252
rect 5136 3047 5143 3356
rect 5176 3327 5183 3473
rect 5256 3447 5263 3473
rect 5276 3427 5283 3776
rect 5336 3747 5343 3783
rect 5396 3783 5403 3996
rect 5576 3987 5583 4273
rect 5413 3828 5427 3833
rect 5436 3816 5443 3873
rect 5396 3776 5423 3783
rect 5373 3763 5387 3773
rect 5373 3760 5393 3763
rect 5376 3756 5393 3760
rect 5316 3516 5323 3593
rect 5356 3516 5363 3573
rect 5396 3527 5403 3753
rect 5416 3487 5423 3776
rect 5516 3747 5523 3893
rect 5380 3483 5393 3487
rect 5376 3476 5393 3483
rect 5380 3473 5393 3476
rect 5436 3463 5443 3733
rect 5536 3547 5543 3973
rect 5596 3963 5603 4513
rect 5616 4467 5623 4593
rect 5636 4567 5643 4816
rect 5696 4687 5703 4823
rect 5696 4556 5703 4593
rect 5716 4567 5723 4813
rect 5676 4487 5683 4523
rect 5656 4336 5663 4413
rect 5676 4387 5683 4433
rect 5693 4387 5707 4393
rect 5716 4363 5723 4513
rect 5696 4356 5723 4363
rect 5676 4047 5683 4293
rect 5647 4003 5660 4007
rect 5647 3996 5663 4003
rect 5647 3993 5660 3996
rect 5576 3956 5603 3963
rect 5576 3907 5583 3956
rect 5596 3816 5603 3913
rect 5576 3707 5583 3783
rect 5616 3667 5623 3783
rect 5467 3523 5480 3527
rect 5467 3516 5483 3523
rect 5467 3513 5480 3516
rect 5416 3456 5443 3463
rect 5196 3296 5203 3413
rect 5236 3308 5243 3333
rect 5156 3256 5183 3263
rect 5156 3247 5163 3256
rect 4767 2836 4793 2843
rect 4596 2788 4603 2833
rect 4636 2776 4643 2833
rect 4776 2776 4783 2813
rect 4816 2787 4823 2892
rect 4476 2740 4483 2743
rect 4456 2483 4463 2733
rect 4473 2727 4487 2740
rect 4516 2687 4523 2743
rect 4436 2476 4463 2483
rect 4336 2367 4343 2413
rect 4376 2407 4383 2443
rect 4247 2256 4263 2267
rect 4247 2253 4260 2256
rect 4333 2267 4347 2273
rect 4236 1967 4243 2213
rect 4276 2147 4283 2223
rect 4316 2167 4323 2223
rect 4336 2187 4343 2213
rect 4316 2087 4323 2153
rect 4276 1967 4283 2073
rect 4336 1967 4343 2173
rect 4136 1827 4143 1853
rect 4113 1748 4127 1753
rect 4136 1747 4143 1773
rect 4036 1436 4043 1513
rect 4076 1467 4083 1693
rect 4096 1443 4103 1473
rect 4076 1436 4103 1443
rect 4016 1400 4023 1403
rect 4013 1387 4027 1400
rect 3916 1180 3923 1183
rect 3816 927 3823 1053
rect 3856 916 3863 1053
rect 3876 967 3883 1172
rect 3913 1167 3927 1180
rect 3956 1127 3963 1172
rect 3976 1027 3983 1073
rect 3996 1067 4003 1253
rect 4056 1248 4063 1403
rect 4116 1387 4123 1653
rect 4136 1627 4143 1693
rect 4156 1567 4163 1913
rect 4233 1907 4247 1913
rect 4176 1747 4183 1893
rect 4256 1867 4263 1953
rect 4256 1736 4263 1832
rect 4276 1787 4283 1913
rect 4356 1883 4363 2373
rect 4416 2367 4423 2443
rect 4433 2260 4447 2273
rect 4456 2267 4463 2413
rect 4476 2303 4483 2573
rect 4516 2507 4523 2673
rect 4536 2476 4543 2693
rect 4573 2487 4587 2493
rect 4516 2440 4523 2443
rect 4513 2427 4527 2440
rect 4596 2443 4603 2633
rect 4616 2587 4623 2743
rect 4656 2707 4663 2743
rect 4676 2587 4683 2733
rect 4696 2647 4703 2753
rect 4756 2567 4763 2743
rect 4616 2487 4623 2533
rect 4736 2487 4743 2533
rect 4776 2503 4783 2713
rect 4796 2567 4803 2743
rect 4776 2496 4803 2503
rect 4753 2480 4767 2493
rect 4756 2476 4763 2480
rect 4796 2476 4803 2496
rect 4816 2487 4823 2733
rect 4596 2436 4623 2443
rect 4556 2423 4563 2432
rect 4536 2416 4563 2423
rect 4476 2296 4503 2303
rect 4436 2256 4443 2260
rect 4376 2187 4383 2213
rect 4416 2147 4423 2223
rect 4476 2207 4483 2273
rect 4376 2007 4383 2053
rect 4396 2047 4403 2113
rect 4436 1968 4443 2193
rect 4476 2107 4483 2172
rect 4476 1956 4483 2013
rect 4496 1967 4503 2296
rect 4536 2287 4543 2416
rect 4576 2407 4583 2433
rect 4576 2307 4583 2333
rect 4596 2307 4603 2413
rect 4616 2367 4623 2436
rect 4676 2367 4683 2443
rect 4696 2387 4703 2433
rect 4716 2387 4723 2473
rect 4836 2427 4843 2873
rect 4907 2833 4913 2847
rect 5016 2827 5023 2953
rect 5056 2927 5063 2963
rect 4913 2807 4927 2812
rect 4913 2800 4933 2807
rect 4916 2796 4933 2800
rect 4920 2793 4933 2796
rect 4900 2746 4920 2747
rect 4900 2743 4913 2746
rect 4896 2736 4913 2743
rect 4900 2733 4913 2736
rect 4856 2707 4863 2733
rect 4956 2743 4963 2813
rect 4973 2803 4987 2813
rect 4973 2800 5003 2803
rect 4976 2796 5003 2800
rect 4996 2776 5003 2796
rect 4956 2736 4983 2743
rect 5036 2740 5043 2743
rect 5033 2727 5047 2740
rect 4876 2476 4883 2533
rect 4916 2488 4923 2553
rect 4956 2487 4963 2573
rect 4853 2423 4867 2433
rect 4853 2420 4883 2423
rect 4856 2416 4883 2420
rect 4567 2296 4583 2307
rect 4567 2293 4580 2296
rect 4516 1967 4523 2213
rect 4536 2127 4543 2223
rect 4576 2203 4583 2223
rect 4556 2200 4583 2203
rect 4556 2196 4587 2200
rect 4536 2047 4543 2113
rect 4556 2087 4563 2196
rect 4573 2187 4587 2196
rect 4576 2027 4583 2152
rect 4596 2127 4603 2213
rect 4596 2027 4603 2053
rect 4593 1960 4607 1973
rect 4616 1963 4623 2353
rect 4636 2167 4643 2293
rect 4676 2268 4683 2332
rect 4656 2167 4663 2223
rect 4736 2103 4743 2413
rect 4876 2267 4883 2416
rect 4896 2407 4903 2443
rect 4936 2347 4943 2443
rect 4976 2427 4983 2633
rect 5056 2527 5063 2833
rect 5076 2727 5083 2933
rect 5096 2747 5103 2963
rect 5136 2887 5143 3012
rect 5156 2947 5163 3233
rect 5216 3207 5223 3252
rect 5216 2996 5223 3033
rect 5256 2963 5263 3213
rect 5276 3167 5283 3353
rect 5356 3296 5363 3393
rect 5336 3260 5343 3263
rect 5333 3247 5347 3260
rect 5376 3027 5383 3263
rect 5313 3000 5327 3013
rect 5316 2996 5323 3000
rect 5127 2796 5153 2803
rect 5196 2747 5203 2963
rect 5236 2956 5263 2963
rect 4756 2127 4763 2254
rect 4796 2147 4803 2223
rect 4736 2096 4763 2103
rect 4647 2013 4653 2027
rect 4676 1968 4683 1993
rect 4696 1987 4703 2033
rect 4596 1956 4603 1960
rect 4616 1956 4643 1963
rect 4376 1907 4383 1953
rect 4416 1920 4423 1923
rect 4456 1920 4463 1923
rect 4413 1907 4427 1920
rect 4453 1907 4467 1920
rect 4356 1876 4383 1883
rect 4273 1748 4287 1752
rect 4176 1547 4183 1693
rect 4213 1667 4227 1673
rect 4236 1667 4243 1703
rect 4296 1667 4303 1813
rect 4376 1767 4383 1876
rect 4313 1747 4327 1753
rect 4416 1747 4423 1833
rect 4336 1627 4343 1703
rect 4376 1647 4383 1703
rect 4147 1406 4160 1407
rect 4147 1393 4153 1406
rect 4116 1247 4123 1333
rect 4136 1327 4143 1393
rect 4216 1387 4223 1473
rect 4256 1447 4263 1573
rect 4027 1183 4040 1187
rect 4027 1176 4043 1183
rect 4027 1173 4040 1176
rect 3896 916 3903 1013
rect 3936 886 3943 973
rect 3956 927 3963 953
rect 3976 916 3983 1013
rect 4016 928 4023 1033
rect 3836 880 3843 883
rect 3833 867 3847 880
rect 3956 847 3963 873
rect 3756 696 3783 703
rect 3816 696 3823 813
rect 3856 707 3863 833
rect 3573 400 3587 413
rect 3756 408 3763 696
rect 3876 666 3883 793
rect 3796 507 3803 663
rect 3956 660 3963 663
rect 3836 467 3843 652
rect 3953 647 3967 660
rect 3976 587 3983 653
rect 3996 647 4003 733
rect 4016 666 4023 753
rect 4056 747 4063 1153
rect 4076 1027 4083 1183
rect 4076 927 4083 1013
rect 4136 923 4143 1253
rect 4156 1183 4163 1371
rect 4196 1287 4203 1333
rect 4236 1327 4243 1434
rect 4296 1436 4303 1513
rect 4336 1487 4343 1572
rect 4376 1547 4383 1633
rect 4416 1587 4423 1693
rect 4436 1647 4443 1853
rect 4476 1787 4483 1873
rect 4496 1763 4503 1913
rect 4516 1887 4523 1932
rect 4536 1807 4543 1913
rect 4476 1756 4503 1763
rect 4476 1736 4483 1756
rect 4456 1667 4463 1693
rect 4333 1440 4347 1452
rect 4356 1447 4363 1533
rect 4396 1503 4403 1553
rect 4387 1496 4403 1503
rect 4336 1436 4343 1440
rect 4253 1347 4267 1353
rect 4196 1216 4203 1273
rect 4156 1176 4173 1183
rect 4236 1180 4243 1183
rect 4233 1167 4247 1180
rect 4256 1167 4263 1293
rect 4196 1047 4203 1153
rect 4276 1087 4283 1353
rect 4296 1227 4303 1313
rect 4316 1287 4323 1403
rect 4376 1367 4383 1493
rect 4416 1487 4423 1513
rect 4476 1487 4483 1673
rect 4496 1627 4503 1703
rect 4460 1443 4473 1447
rect 4456 1436 4473 1443
rect 4460 1433 4473 1436
rect 4356 1127 4363 1183
rect 4376 1147 4383 1173
rect 4216 967 4223 993
rect 4136 916 4163 923
rect 4156 807 4163 916
rect 4253 920 4267 933
rect 4256 916 4263 920
rect 4096 660 4103 663
rect 4093 647 4107 660
rect 3996 607 4003 633
rect 4136 487 4143 653
rect 4156 647 4163 733
rect 4196 708 4203 883
rect 4296 827 4303 1093
rect 4376 947 4383 1133
rect 4396 1127 4403 1393
rect 4456 1216 4463 1333
rect 4476 1307 4483 1393
rect 4496 1327 4503 1573
rect 4536 1467 4543 1692
rect 4556 1547 4563 1873
rect 4576 1747 4583 1923
rect 4636 1767 4643 1956
rect 4756 1967 4763 2096
rect 4696 1887 4703 1923
rect 4736 1867 4743 1923
rect 4776 1887 4783 2033
rect 4796 1968 4803 1993
rect 4816 1956 4823 2033
rect 4856 2007 4863 2173
rect 4876 2087 4883 2213
rect 4896 2147 4903 2313
rect 4996 2307 5003 2513
rect 5076 2507 5083 2653
rect 5136 2647 5143 2713
rect 5216 2707 5223 2933
rect 5093 2507 5107 2513
rect 5093 2480 5107 2493
rect 5096 2476 5103 2480
rect 4956 2256 4963 2293
rect 5016 2267 5023 2433
rect 5036 2347 5043 2443
rect 4916 2103 4923 2213
rect 4936 2127 4943 2223
rect 4916 2096 4943 2103
rect 4876 2047 4883 2073
rect 4716 1768 4723 1793
rect 4576 1647 4583 1693
rect 4596 1587 4603 1703
rect 4616 1540 4653 1543
rect 4613 1536 4653 1540
rect 4613 1527 4627 1536
rect 4676 1487 4683 1753
rect 4756 1736 4763 1773
rect 4796 1703 4803 1913
rect 4836 1903 4843 1912
rect 4816 1896 4843 1903
rect 4816 1747 4823 1896
rect 4836 1736 4843 1793
rect 4876 1736 4883 1833
rect 4916 1747 4923 1993
rect 4936 1887 4943 2096
rect 4956 1967 4963 2033
rect 4996 2007 5003 2173
rect 5016 1967 5023 2213
rect 4973 1863 4987 1873
rect 4973 1860 5003 1863
rect 4976 1856 5003 1860
rect 4736 1687 4743 1703
rect 4776 1696 4803 1703
rect 4736 1676 4753 1687
rect 4740 1673 4753 1676
rect 4527 1443 4540 1447
rect 4527 1436 4543 1443
rect 4527 1433 4540 1436
rect 4556 1347 4563 1403
rect 4596 1367 4603 1393
rect 4493 1220 4507 1233
rect 4536 1223 4543 1313
rect 4596 1267 4603 1353
rect 4616 1287 4623 1453
rect 4636 1447 4643 1473
rect 4696 1463 4703 1673
rect 4736 1507 4743 1573
rect 4676 1456 4703 1463
rect 4676 1436 4683 1456
rect 4713 1440 4727 1453
rect 4736 1447 4743 1493
rect 4716 1436 4723 1440
rect 4636 1267 4643 1393
rect 4656 1347 4663 1403
rect 4496 1216 4503 1220
rect 4536 1216 4563 1223
rect 4556 1186 4563 1216
rect 4676 1227 4683 1253
rect 4396 1007 4403 1113
rect 4476 1107 4483 1183
rect 4516 1127 4523 1183
rect 4556 1127 4563 1172
rect 4576 1067 4583 1173
rect 4616 1107 4623 1183
rect 4656 1147 4663 1183
rect 4476 1027 4483 1053
rect 4616 1027 4623 1093
rect 4333 928 4347 933
rect 4376 916 4383 933
rect 4476 916 4483 1013
rect 4516 916 4523 993
rect 4576 886 4583 1013
rect 4676 947 4683 1173
rect 4696 967 4703 1403
rect 4736 1247 4743 1393
rect 4756 1248 4763 1473
rect 4776 1227 4783 1696
rect 4856 1700 4863 1703
rect 4816 1507 4823 1693
rect 4853 1687 4867 1700
rect 4896 1647 4903 1703
rect 4916 1383 4923 1693
rect 4896 1376 4923 1383
rect 4836 1360 4843 1363
rect 4833 1347 4847 1360
rect 4716 1147 4723 1173
rect 4736 1107 4743 1183
rect 4796 1107 4803 1233
rect 4816 1227 4823 1333
rect 4856 1216 4863 1253
rect 4896 1227 4903 1376
rect 4936 1243 4943 1753
rect 4956 1547 4963 1813
rect 4996 1736 5003 1856
rect 5036 1768 5043 2293
rect 5056 2226 5063 2413
rect 5136 2407 5143 2433
rect 5156 2347 5163 2693
rect 5236 2523 5243 2956
rect 5296 2847 5303 2963
rect 5336 2960 5343 2963
rect 5333 2947 5347 2960
rect 5396 2947 5403 3252
rect 5416 3227 5423 3456
rect 5476 3296 5483 3433
rect 5496 3367 5503 3472
rect 5456 3247 5463 3263
rect 5453 3227 5467 3233
rect 5496 3027 5503 3263
rect 5536 3027 5543 3533
rect 5556 3527 5563 3553
rect 5596 3516 5603 3573
rect 5627 3553 5633 3567
rect 5633 3520 5647 3532
rect 5656 3523 5663 3973
rect 5676 3927 5683 3993
rect 5696 3847 5703 4356
rect 5736 4343 5743 4896
rect 5776 4856 5783 4893
rect 5796 4447 5803 4812
rect 5716 4336 5743 4343
rect 5756 4336 5763 4373
rect 5716 3887 5723 4336
rect 5836 4347 5843 4913
rect 5736 4267 5743 4293
rect 5776 4283 5783 4303
rect 5816 4300 5823 4303
rect 5813 4287 5827 4300
rect 5776 4276 5803 4283
rect 5736 4047 5743 4232
rect 5756 4067 5763 4093
rect 5776 4036 5783 4253
rect 5796 4183 5803 4276
rect 5796 4176 5823 4183
rect 5756 4000 5763 4003
rect 5736 3963 5743 3993
rect 5753 3987 5767 4000
rect 5736 3956 5763 3963
rect 5756 3816 5763 3956
rect 5776 3827 5783 3873
rect 5676 3547 5683 3773
rect 5696 3667 5703 3783
rect 5796 3786 5803 3993
rect 5636 3516 5643 3520
rect 5656 3516 5673 3523
rect 5716 3516 5723 3553
rect 5776 3527 5783 3773
rect 5576 3447 5583 3483
rect 5676 3483 5683 3512
rect 5796 3487 5803 3733
rect 5816 3647 5823 4176
rect 5656 3476 5683 3483
rect 5656 3407 5663 3476
rect 5656 3336 5663 3393
rect 5696 3367 5703 3473
rect 5416 2887 5423 2993
rect 5456 2947 5463 2963
rect 5293 2780 5307 2793
rect 5296 2776 5303 2780
rect 5316 2707 5323 2743
rect 5336 2647 5343 2873
rect 5456 2847 5463 2933
rect 5496 2907 5503 2952
rect 5536 2947 5543 3013
rect 5556 2907 5563 3294
rect 5576 2996 5583 3213
rect 5636 2996 5643 3033
rect 5656 2966 5663 2993
rect 5416 2776 5423 2813
rect 5396 2667 5403 2732
rect 5436 2707 5443 2743
rect 5236 2516 5263 2523
rect 5196 2387 5203 2432
rect 5116 2256 5123 2293
rect 5076 2027 5083 2153
rect 5096 2087 5103 2223
rect 5196 2223 5203 2333
rect 5236 2323 5243 2433
rect 5256 2427 5263 2516
rect 5276 2488 5283 2513
rect 5296 2447 5303 2513
rect 5216 2316 5243 2323
rect 5216 2267 5223 2316
rect 5256 2307 5263 2373
rect 5296 2267 5303 2412
rect 5436 2407 5443 2473
rect 5456 2443 5463 2633
rect 5476 2487 5483 2873
rect 5553 2820 5567 2833
rect 5676 2823 5683 2893
rect 5696 2847 5703 3073
rect 5736 3008 5743 3353
rect 5816 3087 5823 3513
rect 5776 3008 5783 3033
rect 5756 2960 5763 2963
rect 5753 2947 5767 2960
rect 5556 2816 5563 2820
rect 5676 2816 5703 2823
rect 5496 2776 5523 2783
rect 5496 2747 5503 2776
rect 5696 2776 5703 2816
rect 5616 2736 5643 2743
rect 5516 2507 5523 2713
rect 5636 2707 5643 2736
rect 5656 2687 5663 2774
rect 5716 2723 5723 2743
rect 5756 2740 5763 2743
rect 5696 2716 5723 2723
rect 5753 2727 5767 2740
rect 5556 2547 5563 2673
rect 5520 2483 5533 2487
rect 5516 2476 5533 2483
rect 5520 2474 5533 2476
rect 5520 2473 5540 2474
rect 5556 2467 5563 2533
rect 5696 2447 5703 2716
rect 5756 2607 5763 2653
rect 5756 2507 5763 2533
rect 5776 2487 5783 2733
rect 5456 2436 5483 2443
rect 5336 2347 5343 2373
rect 5376 2307 5383 2403
rect 5336 2267 5343 2293
rect 5373 2260 5387 2272
rect 5376 2256 5383 2260
rect 5416 2256 5423 2313
rect 5436 2267 5443 2333
rect 5476 2307 5483 2436
rect 5496 2347 5503 2432
rect 5516 2307 5523 2353
rect 5536 2327 5543 2433
rect 5536 2287 5543 2313
rect 5176 2216 5203 2223
rect 5153 2127 5167 2133
rect 5147 2120 5167 2127
rect 5147 2116 5163 2120
rect 5147 2113 5160 2116
rect 5056 1967 5063 1993
rect 5096 1987 5103 2033
rect 5096 1976 5113 1987
rect 5100 1973 5113 1976
rect 5136 1956 5143 2033
rect 5156 1967 5163 2013
rect 5056 1807 5063 1913
rect 5076 1887 5083 1923
rect 4976 1527 4983 1693
rect 4996 1467 5003 1493
rect 5016 1487 5023 1513
rect 4967 1436 4983 1443
rect 5036 1436 5043 1673
rect 4956 1267 4963 1434
rect 4916 1236 4943 1243
rect 4627 936 4663 943
rect 4656 927 4663 936
rect 4656 926 4680 927
rect 4656 916 4673 926
rect 4660 913 4673 916
rect 4756 916 4763 993
rect 4276 707 4283 753
rect 4396 723 4403 883
rect 4496 880 4503 883
rect 4493 867 4507 880
rect 4376 716 4403 723
rect 4376 708 4383 716
rect 4296 696 4343 703
rect 4216 660 4223 663
rect 4213 647 4227 660
rect 4256 567 4263 663
rect 4296 527 4303 696
rect 3576 396 3583 400
rect 3196 176 3203 273
rect 3256 203 3263 233
rect 3256 196 3283 203
rect 3256 147 3263 174
rect 3016 136 3043 143
rect 3016 47 3023 136
rect 3036 43 3043 93
rect 3056 67 3063 113
rect 3076 87 3083 143
rect 3176 140 3183 143
rect 3173 127 3187 140
rect 3276 107 3283 196
rect 3316 176 3323 253
rect 3396 146 3403 253
rect 3456 176 3463 331
rect 3496 247 3503 363
rect 3556 176 3563 253
rect 3596 176 3603 213
rect 3636 187 3643 353
rect 3356 87 3363 143
rect 3476 140 3483 143
rect 3473 127 3487 140
rect 3516 127 3523 173
rect 3476 87 3483 113
rect 3576 87 3583 143
rect 3616 107 3623 143
rect 3656 107 3663 394
rect 3796 366 3803 393
rect 3696 227 3703 363
rect 3736 267 3743 363
rect 3716 47 3723 143
rect 3036 36 3073 43
rect 2836 -24 2863 -17
rect 3816 -17 3823 293
rect 3836 187 3843 352
rect 3896 307 3903 453
rect 3976 396 3983 433
rect 3916 366 3923 393
rect 4056 363 4063 433
rect 4096 423 4103 473
rect 4113 423 4127 433
rect 4096 420 4127 423
rect 4096 416 4123 420
rect 4116 396 4123 416
rect 4296 396 4303 433
rect 4316 403 4323 653
rect 4436 666 4443 853
rect 4453 707 4467 713
rect 4536 696 4543 753
rect 4353 647 4367 652
rect 4316 396 4343 403
rect 3896 176 3903 253
rect 3956 207 3963 352
rect 3996 203 4003 363
rect 4056 356 4103 363
rect 4136 327 4143 363
rect 4236 267 4243 352
rect 4276 327 4283 363
rect 4316 287 4323 353
rect 4296 207 4303 233
rect 3976 196 4003 203
rect 3976 183 3983 196
rect 3956 176 3983 183
rect 3833 127 3847 132
rect 3916 107 3923 132
rect 3956 47 3963 176
rect 3976 27 3983 132
rect 4076 87 4083 133
rect 4096 107 4103 174
rect 4127 183 4140 187
rect 4127 176 4143 183
rect 4127 173 4140 176
rect 4316 176 4323 273
rect 4336 227 4343 396
rect 4356 343 4363 433
rect 4376 407 4383 553
rect 4416 423 4423 653
rect 4476 660 4483 663
rect 4396 416 4423 423
rect 4396 396 4403 416
rect 4436 396 4443 652
rect 4473 647 4487 660
rect 4576 567 4583 793
rect 4636 696 4643 793
rect 4676 728 4683 892
rect 4816 807 4823 1173
rect 4836 1127 4843 1183
rect 4896 943 4903 1073
rect 4916 1047 4923 1236
rect 5016 1216 5023 1253
rect 5036 1223 5043 1353
rect 5056 1247 5063 1703
rect 5076 1367 5083 1693
rect 5096 1687 5103 1853
rect 5116 1827 5123 1923
rect 5156 1867 5163 1913
rect 5176 1787 5183 2216
rect 5216 2183 5223 2213
rect 5236 2187 5243 2223
rect 5276 2216 5303 2223
rect 5216 2176 5233 2183
rect 5196 2107 5203 2153
rect 5196 1967 5203 2053
rect 5236 1956 5243 1993
rect 5296 1967 5303 2216
rect 5336 2216 5363 2223
rect 5316 2127 5323 2213
rect 5336 2187 5343 2216
rect 5393 2207 5407 2212
rect 5316 1987 5323 2033
rect 5336 2027 5343 2173
rect 5216 1920 5223 1923
rect 5213 1907 5227 1920
rect 5116 1747 5123 1773
rect 5236 1747 5243 1873
rect 5296 1863 5303 1913
rect 5316 1887 5323 1973
rect 5333 1963 5347 1973
rect 5356 1968 5363 2133
rect 5436 2107 5443 2213
rect 5456 2147 5463 2273
rect 5513 2260 5527 2272
rect 5516 2256 5523 2260
rect 5556 2256 5563 2432
rect 5576 2327 5583 2353
rect 5576 2267 5583 2292
rect 5496 2187 5503 2223
rect 5333 1960 5353 1963
rect 5336 1956 5353 1960
rect 5393 1960 5407 1973
rect 5396 1956 5403 1960
rect 5296 1856 5323 1863
rect 5256 1736 5263 1793
rect 5296 1748 5303 1793
rect 5316 1767 5323 1856
rect 5336 1827 5343 1853
rect 5216 1706 5223 1733
rect 5136 1647 5143 1703
rect 5096 1447 5103 1613
rect 5196 1587 5203 1673
rect 5236 1603 5243 1693
rect 5236 1596 5263 1603
rect 5116 1436 5123 1553
rect 5156 1436 5163 1473
rect 5196 1448 5203 1573
rect 5136 1400 5143 1403
rect 5096 1327 5103 1393
rect 5133 1387 5147 1400
rect 5236 1387 5243 1573
rect 5116 1247 5123 1333
rect 5036 1216 5063 1223
rect 4936 1027 4943 1213
rect 4896 936 4923 943
rect 4916 916 4923 936
rect 4836 887 4843 914
rect 4896 880 4903 883
rect 4836 847 4843 873
rect 4893 867 4907 880
rect 4356 336 4383 343
rect 4356 187 4363 313
rect 4376 283 4383 336
rect 4456 307 4463 363
rect 4496 347 4503 553
rect 4616 547 4623 663
rect 4656 627 4663 663
rect 4556 427 4563 473
rect 4716 447 4723 713
rect 4556 396 4563 413
rect 4516 307 4523 352
rect 4536 327 4543 363
rect 4376 276 4403 283
rect 4153 127 4167 132
rect 4236 127 4243 173
rect 4376 107 4383 253
rect 4396 187 4403 276
rect 4436 176 4443 253
rect 4473 180 4487 193
rect 4476 176 4483 180
rect 4456 107 4463 143
rect 4516 146 4523 233
rect 4613 188 4627 193
rect 4636 183 4643 433
rect 4673 400 4687 413
rect 4756 408 4763 593
rect 4776 587 4783 663
rect 4856 607 4863 753
rect 4916 708 4923 753
rect 4956 708 4963 1173
rect 4996 1007 5003 1172
rect 5056 1007 5063 1216
rect 5136 1216 5143 1253
rect 4976 996 4993 1003
rect 4976 927 4983 996
rect 5056 916 5063 953
rect 5076 927 5083 1173
rect 5116 923 5123 1183
rect 5156 1087 5163 1172
rect 5107 916 5123 923
rect 5176 916 5183 1053
rect 5196 1047 5203 1373
rect 5256 1367 5263 1596
rect 5276 1347 5283 1703
rect 5316 1696 5343 1703
rect 5336 1667 5343 1696
rect 5326 1653 5327 1660
rect 5313 1647 5327 1653
rect 5356 1587 5363 1893
rect 5376 1867 5383 1923
rect 5376 1827 5383 1853
rect 5416 1847 5423 1923
rect 5416 1736 5423 1812
rect 5436 1767 5443 1913
rect 5456 1847 5463 2112
rect 5476 1967 5483 2113
rect 5516 1956 5523 2053
rect 5536 1987 5543 2191
rect 5576 2127 5583 2213
rect 5596 1947 5603 2393
rect 5616 2367 5623 2443
rect 5760 2443 5773 2447
rect 5756 2436 5773 2443
rect 5760 2433 5773 2436
rect 5616 2247 5623 2313
rect 5636 2256 5643 2293
rect 5676 2283 5683 2353
rect 5696 2307 5703 2433
rect 5676 2276 5703 2283
rect 5436 1683 5443 1703
rect 5416 1676 5443 1683
rect 5387 1633 5393 1647
rect 5416 1587 5423 1676
rect 5496 1667 5503 1912
rect 5536 1847 5543 1923
rect 5576 1827 5583 1913
rect 5536 1736 5543 1793
rect 5616 1787 5623 2212
rect 5636 1956 5643 2193
rect 5676 2147 5683 2223
rect 5696 2207 5703 2276
rect 5716 2207 5723 2433
rect 5696 1956 5703 2153
rect 5656 1867 5663 1923
rect 5656 1747 5663 1813
rect 5696 1767 5703 1893
rect 5636 1703 5643 1734
rect 5716 1747 5723 1973
rect 5516 1647 5523 1693
rect 5556 1683 5563 1703
rect 5596 1696 5643 1703
rect 5536 1676 5563 1683
rect 5356 1436 5383 1443
rect 5376 1406 5383 1436
rect 5336 1387 5343 1403
rect 5396 1387 5403 1453
rect 5436 1448 5443 1593
rect 5536 1547 5543 1676
rect 5496 1487 5503 1513
rect 5476 1436 5483 1473
rect 5327 1376 5343 1387
rect 5327 1373 5340 1376
rect 5213 1223 5227 1233
rect 5213 1220 5243 1223
rect 5216 1216 5243 1220
rect 5216 1147 5223 1173
rect 5256 1147 5263 1183
rect 5316 1107 5323 1333
rect 5336 1227 5343 1253
rect 5376 1216 5383 1353
rect 5436 1227 5443 1353
rect 5356 1087 5363 1172
rect 5096 883 5103 914
rect 5076 876 5103 883
rect 4987 856 5013 863
rect 5076 747 5083 876
rect 5156 880 5163 883
rect 5116 767 5123 873
rect 5153 867 5167 880
rect 5093 700 5107 713
rect 5096 696 5103 700
rect 4896 587 4903 663
rect 4916 567 4923 613
rect 4676 396 4683 400
rect 4767 396 4783 403
rect 4816 396 4823 433
rect 4676 187 4683 253
rect 4696 227 4703 293
rect 4736 267 4743 363
rect 4776 267 4783 396
rect 4956 396 4963 533
rect 4896 367 4903 394
rect 4996 366 5003 693
rect 5136 666 5143 753
rect 5156 707 5163 813
rect 5196 767 5203 883
rect 5236 827 5243 993
rect 5256 927 5263 1073
rect 5396 1067 5403 1183
rect 5436 1147 5443 1173
rect 5436 1047 5443 1133
rect 5456 1127 5463 1371
rect 5496 1343 5503 1403
rect 5516 1367 5523 1393
rect 5496 1336 5523 1343
rect 5316 928 5323 953
rect 5173 700 5187 713
rect 5176 696 5183 700
rect 5256 703 5263 873
rect 5296 807 5303 883
rect 5276 756 5323 763
rect 5276 727 5283 756
rect 5296 707 5303 733
rect 5256 696 5283 703
rect 5016 656 5043 663
rect 4796 247 4803 293
rect 4636 176 4663 183
rect 4496 27 4503 133
rect 4596 140 4603 143
rect 4593 127 4607 140
rect 4593 107 4607 113
rect 4656 87 4663 176
rect 4736 176 4743 213
rect 4796 146 4803 233
rect 4876 176 4883 253
rect 4936 243 4943 352
rect 5016 327 5023 656
rect 5133 408 5147 413
rect 5116 360 5123 363
rect 5113 347 5127 360
rect 4916 236 4943 243
rect 4716 140 4723 143
rect 4713 127 4727 140
rect 4836 87 4843 143
rect 4896 140 4903 143
rect 4893 127 4907 140
rect 4916 47 4923 236
rect 4976 176 4983 273
rect 5136 247 5143 353
rect 5056 207 5063 233
rect 5053 187 5067 193
rect 4936 127 4943 153
rect 4980 125 5000 127
rect 4987 113 4993 125
rect 5036 107 5043 143
rect 5076 107 5083 213
rect 5156 207 5163 653
rect 5216 396 5223 513
rect 5236 467 5243 663
rect 5276 647 5283 696
rect 5316 696 5323 756
rect 5336 727 5343 873
rect 5356 767 5363 1033
rect 5376 927 5383 973
rect 5476 947 5483 1233
rect 5496 1223 5503 1313
rect 5516 1287 5523 1336
rect 5536 1307 5543 1493
rect 5556 1447 5563 1553
rect 5616 1436 5623 1696
rect 5696 1700 5703 1703
rect 5653 1687 5667 1693
rect 5693 1687 5707 1700
rect 5696 1406 5703 1473
rect 5716 1443 5723 1693
rect 5736 1507 5743 2293
rect 5796 2287 5803 2833
rect 5816 2747 5823 2994
rect 5816 2667 5823 2693
rect 5836 2643 5843 4293
rect 5816 2636 5843 2643
rect 5756 2167 5763 2193
rect 5776 2147 5783 2173
rect 5816 1987 5823 2636
rect 5836 2487 5843 2613
rect 5836 2327 5843 2433
rect 5756 1467 5763 1973
rect 5776 1487 5783 1773
rect 5796 1567 5803 1933
rect 5816 1907 5823 1952
rect 5716 1436 5743 1443
rect 5816 1447 5823 1853
rect 5636 1327 5643 1403
rect 5616 1247 5623 1293
rect 5656 1283 5663 1373
rect 5647 1276 5663 1283
rect 5496 1216 5523 1223
rect 5496 987 5503 1193
rect 5636 1183 5643 1273
rect 5616 1176 5643 1183
rect 5420 943 5433 947
rect 5416 933 5433 943
rect 5416 916 5423 933
rect 5396 847 5403 872
rect 5376 723 5383 793
rect 5356 716 5383 723
rect 5356 696 5363 716
rect 5396 707 5403 773
rect 5336 660 5343 663
rect 5376 660 5383 663
rect 5333 647 5347 660
rect 5373 647 5387 660
rect 5376 607 5383 633
rect 5236 427 5243 453
rect 5256 408 5263 593
rect 5133 180 5147 193
rect 5136 176 5143 180
rect 5176 176 5183 313
rect 5276 188 5283 353
rect 5296 347 5303 553
rect 5316 407 5323 433
rect 5416 403 5423 713
rect 5433 707 5447 713
rect 5476 708 5483 933
rect 5493 928 5507 933
rect 5533 928 5547 933
rect 5573 920 5587 933
rect 5596 927 5603 1093
rect 5576 916 5583 920
rect 5496 727 5503 773
rect 5516 767 5523 883
rect 5556 807 5563 883
rect 5596 847 5603 873
rect 5536 796 5553 803
rect 5536 707 5543 796
rect 5616 787 5623 1013
rect 5636 927 5643 1033
rect 5656 987 5663 1233
rect 5676 1223 5683 1313
rect 5716 1307 5723 1393
rect 5756 1247 5763 1293
rect 5676 1216 5703 1223
rect 5676 1067 5683 1193
rect 5816 1183 5823 1273
rect 5796 1176 5823 1183
rect 5836 1163 5843 2273
rect 5816 1156 5843 1163
rect 5676 967 5683 1053
rect 5673 920 5687 932
rect 5676 916 5683 920
rect 5716 916 5723 953
rect 5576 703 5583 773
rect 5556 696 5583 703
rect 5593 700 5607 713
rect 5636 708 5643 793
rect 5676 783 5683 833
rect 5696 807 5703 883
rect 5676 776 5703 783
rect 5596 696 5603 700
rect 5436 427 5443 653
rect 5456 627 5463 663
rect 5416 396 5443 403
rect 5476 396 5483 633
rect 5496 607 5503 663
rect 5536 627 5543 653
rect 5556 447 5563 696
rect 5336 360 5343 363
rect 5376 360 5383 363
rect 5316 227 5323 353
rect 5333 347 5347 360
rect 5373 347 5387 360
rect 5376 267 5383 333
rect 5416 247 5423 353
rect 5116 140 5123 143
rect 5113 127 5127 140
rect 5216 107 5223 173
rect 5316 147 5323 192
rect 5356 176 5363 213
rect 5436 188 5443 396
rect 5456 287 5463 353
rect 5496 327 5503 363
rect 5476 176 5483 213
rect 5516 176 5523 253
rect 5536 247 5543 363
rect 5576 327 5583 613
rect 5616 467 5623 663
rect 5656 660 5663 663
rect 5653 647 5667 660
rect 5636 396 5643 453
rect 5656 427 5663 633
rect 5676 408 5683 653
rect 5696 627 5703 776
rect 5756 696 5763 973
rect 5796 667 5803 1113
rect 5547 236 5563 243
rect 5556 187 5563 236
rect 5576 183 5583 273
rect 5596 207 5603 293
rect 5576 176 5623 183
rect 5656 176 5663 352
rect 5676 207 5683 333
rect 5696 183 5703 233
rect 5716 207 5723 573
rect 5816 427 5823 1156
rect 5753 400 5767 413
rect 5756 396 5763 400
rect 5776 327 5783 363
rect 5836 327 5843 1133
rect 5696 176 5723 183
rect 5773 180 5787 193
rect 5776 176 5783 180
rect 5496 140 5503 143
rect 5493 127 5507 140
rect 5576 127 5583 176
rect 5716 147 5723 176
rect 3816 -24 3843 -17
<< m3contact >>
rect 653 5393 667 5407
rect 753 5393 767 5407
rect 213 5374 227 5388
rect 333 5374 347 5388
rect 373 5374 387 5388
rect 613 5374 627 5388
rect 693 5374 707 5388
rect 273 5353 287 5367
rect 33 5233 47 5247
rect 73 5173 87 5187
rect 113 5173 127 5187
rect 53 5074 67 5088
rect 313 5313 327 5327
rect 353 5333 367 5347
rect 493 5332 507 5346
rect 273 5133 287 5147
rect 113 5074 127 5088
rect 153 5074 167 5088
rect 193 5074 207 5088
rect 233 5074 247 5088
rect 73 5013 87 5027
rect 133 5032 147 5046
rect 313 5073 327 5087
rect 213 5033 227 5047
rect 193 4993 207 5007
rect 253 4993 267 5007
rect 93 4933 107 4947
rect 213 4933 227 4947
rect 613 5333 627 5347
rect 713 5332 727 5346
rect 673 5313 687 5327
rect 813 5374 827 5388
rect 2033 5473 2047 5487
rect 2093 5473 2107 5487
rect 2173 5473 2187 5487
rect 2213 5473 2227 5487
rect 2653 5473 2667 5487
rect 2833 5473 2847 5487
rect 1373 5413 1387 5427
rect 1453 5413 1467 5427
rect 1853 5413 1867 5427
rect 1313 5374 1327 5388
rect 1413 5374 1427 5388
rect 1473 5374 1487 5388
rect 1513 5374 1527 5388
rect 673 5273 687 5287
rect 713 5273 727 5287
rect 753 5273 767 5287
rect 793 5273 807 5287
rect 553 5233 567 5247
rect 593 5233 607 5247
rect 693 5233 707 5247
rect 553 5093 567 5107
rect 393 5074 407 5088
rect 453 5074 467 5088
rect 513 5074 527 5088
rect 653 5074 667 5088
rect 333 5033 347 5047
rect 373 5032 387 5046
rect 413 4973 427 4987
rect 233 4893 247 4907
rect 273 4893 287 4907
rect 313 4893 327 4907
rect 53 4853 67 4867
rect 93 4854 107 4868
rect 153 4853 167 4867
rect 193 4854 207 4868
rect 53 4813 67 4827
rect 313 4854 327 4868
rect 353 4854 367 4868
rect 413 4853 427 4867
rect 533 5032 547 5046
rect 693 4993 707 5007
rect 653 4973 667 4987
rect 493 4933 507 4947
rect 573 4873 587 4887
rect 613 4854 627 4868
rect 273 4812 287 4826
rect 333 4812 347 4826
rect 153 4773 167 4787
rect 413 4812 427 4826
rect 453 4812 467 4826
rect 593 4812 607 4826
rect 493 4773 507 4787
rect 813 5093 827 5107
rect 773 5032 787 5046
rect 813 5013 827 5027
rect 793 4993 807 5007
rect 713 4953 727 4967
rect 753 4953 767 4967
rect 713 4913 727 4927
rect 753 4873 767 4887
rect 733 4812 747 4826
rect 693 4773 707 4787
rect 1033 5333 1047 5347
rect 1073 5332 1087 5346
rect 953 5313 967 5327
rect 953 5233 967 5247
rect 1033 5213 1047 5227
rect 973 5133 987 5147
rect 873 5074 887 5088
rect 993 5113 1007 5127
rect 933 5033 947 5047
rect 893 5013 907 5027
rect 853 4973 867 4987
rect 933 4973 947 4987
rect 833 4873 847 4887
rect 973 5073 987 5087
rect 1193 5332 1207 5346
rect 1373 5333 1387 5347
rect 1433 5332 1447 5346
rect 1133 5313 1147 5327
rect 1613 5373 1627 5387
rect 1673 5374 1687 5388
rect 1793 5374 1807 5388
rect 1733 5353 1747 5367
rect 1533 5332 1547 5346
rect 1573 5332 1587 5346
rect 1613 5332 1627 5346
rect 1473 5273 1487 5287
rect 1133 5253 1147 5267
rect 1933 5374 1947 5388
rect 2013 5373 2027 5387
rect 1813 5332 1827 5346
rect 1853 5332 1867 5346
rect 1833 5313 1847 5327
rect 1733 5293 1747 5307
rect 1773 5293 1787 5307
rect 1793 5272 1807 5286
rect 1833 5273 1847 5287
rect 1293 5233 1307 5247
rect 1473 5233 1487 5247
rect 1653 5233 1667 5247
rect 1793 5233 1807 5247
rect 1293 5193 1307 5207
rect 1073 5173 1087 5187
rect 1113 5173 1127 5187
rect 1213 5173 1227 5187
rect 1073 5074 1087 5088
rect 1013 5032 1027 5046
rect 993 5013 1007 5027
rect 1053 5013 1067 5027
rect 973 4953 987 4967
rect 953 4933 967 4947
rect 893 4873 907 4887
rect 833 4812 847 4826
rect 793 4753 807 4767
rect 653 4713 667 4727
rect 693 4653 707 4667
rect 113 4593 127 4607
rect 373 4593 387 4607
rect 433 4593 447 4607
rect 73 4553 87 4567
rect 153 4553 167 4567
rect 213 4554 227 4568
rect 273 4554 287 4568
rect 313 4554 327 4568
rect 353 4554 367 4568
rect 393 4554 407 4568
rect 473 4554 487 4568
rect 513 4554 527 4568
rect 573 4554 587 4568
rect 613 4554 627 4568
rect 653 4554 667 4568
rect 733 4633 747 4647
rect 893 4713 907 4727
rect 733 4554 747 4568
rect 833 4554 847 4568
rect 93 4512 107 4526
rect 153 4512 167 4526
rect 233 4512 247 4526
rect 273 4513 287 4527
rect 193 4473 207 4487
rect 333 4512 347 4526
rect 453 4512 467 4526
rect 513 4513 527 4527
rect 393 4473 407 4487
rect 273 4433 287 4447
rect 373 4433 387 4447
rect 53 4373 67 4387
rect 313 4373 327 4387
rect 93 4334 107 4348
rect 253 4333 267 4347
rect 73 4292 87 4306
rect 193 4292 207 4306
rect 253 4292 267 4306
rect 113 4113 127 4127
rect 293 4292 307 4306
rect 353 4293 367 4307
rect 153 4034 167 4048
rect 193 4033 207 4047
rect 233 4034 247 4048
rect 273 4034 287 4048
rect 193 3992 207 4006
rect 253 3973 267 3987
rect 133 3953 147 3967
rect 233 3893 247 3907
rect 153 3814 167 3828
rect 193 3814 207 3828
rect 593 4493 607 4507
rect 653 4453 667 4467
rect 553 4413 567 4427
rect 393 4393 407 4407
rect 493 4393 507 4407
rect 473 4353 487 4367
rect 413 4334 427 4348
rect 433 4292 447 4306
rect 373 4153 387 4167
rect 413 4153 427 4167
rect 373 4113 387 4127
rect 353 3992 367 4006
rect 313 3973 327 3987
rect 313 3952 327 3966
rect 293 3893 307 3907
rect 253 3853 267 3867
rect 293 3853 307 3867
rect 113 3772 127 3786
rect 153 3773 167 3787
rect 353 3893 367 3907
rect 313 3833 327 3847
rect 13 3613 27 3627
rect 73 3693 87 3707
rect 193 3733 207 3747
rect 53 3513 67 3527
rect 113 3513 127 3527
rect 53 3473 67 3487
rect 73 3453 87 3467
rect 133 3453 147 3467
rect 173 3393 187 3407
rect 93 3353 107 3367
rect 73 3313 87 3327
rect 53 3293 67 3307
rect 53 3253 67 3267
rect 33 3013 47 3027
rect 73 3233 87 3247
rect 153 3252 167 3266
rect 133 3193 147 3207
rect 113 3013 127 3027
rect 73 2994 87 3008
rect 253 3772 267 3786
rect 293 3772 307 3786
rect 393 3873 407 3887
rect 393 3813 407 3827
rect 393 3773 407 3787
rect 313 3733 327 3747
rect 373 3733 387 3747
rect 213 3693 227 3707
rect 393 3653 407 3667
rect 313 3533 327 3547
rect 353 3533 367 3547
rect 473 4073 487 4087
rect 553 4373 567 4387
rect 613 4373 627 4387
rect 593 4334 607 4348
rect 633 4353 647 4367
rect 693 4353 707 4367
rect 533 4292 547 4306
rect 573 4193 587 4207
rect 433 3993 447 4007
rect 493 3913 507 3927
rect 493 3873 507 3887
rect 533 3873 547 3887
rect 453 3833 467 3847
rect 433 3813 447 3827
rect 433 3773 447 3787
rect 473 3772 487 3786
rect 533 3693 547 3707
rect 533 3613 547 3627
rect 433 3553 447 3567
rect 533 3553 547 3567
rect 213 3513 227 3527
rect 253 3514 267 3528
rect 193 3353 207 3367
rect 253 3453 267 3467
rect 213 3294 227 3308
rect 433 3514 447 3528
rect 413 3472 427 3486
rect 453 3472 467 3486
rect 353 3393 367 3407
rect 473 3373 487 3387
rect 313 3293 327 3307
rect 373 3294 387 3308
rect 433 3294 447 3308
rect 473 3294 487 3308
rect 573 4034 587 4048
rect 753 4513 767 4527
rect 1133 5133 1147 5147
rect 1173 5113 1187 5127
rect 1133 5074 1147 5088
rect 1253 5133 1267 5147
rect 1413 5133 1427 5147
rect 1753 5133 1767 5147
rect 1393 5113 1407 5127
rect 1353 5074 1367 5088
rect 1133 5013 1147 5027
rect 1113 4993 1127 5007
rect 1213 5013 1227 5027
rect 1193 4953 1207 4967
rect 1133 4913 1147 4927
rect 1113 4873 1127 4887
rect 953 4633 967 4647
rect 1013 4793 1027 4807
rect 1113 4773 1127 4787
rect 1073 4753 1087 4767
rect 1013 4653 1027 4667
rect 993 4593 1007 4607
rect 1093 4593 1107 4607
rect 1013 4554 1027 4568
rect 1053 4554 1067 4568
rect 953 4512 967 4526
rect 993 4512 1007 4526
rect 713 4333 727 4347
rect 953 4413 967 4427
rect 1153 4893 1167 4907
rect 1273 4993 1287 5007
rect 1233 4973 1247 4987
rect 1213 4854 1227 4868
rect 1253 4854 1267 4868
rect 1293 4893 1307 4907
rect 1333 4893 1347 4907
rect 1193 4812 1207 4826
rect 1253 4713 1267 4727
rect 1313 4812 1327 4826
rect 1233 4573 1247 4587
rect 1273 4573 1287 4587
rect 1133 4493 1147 4507
rect 1073 4453 1087 4467
rect 1153 4453 1167 4467
rect 1193 4453 1207 4467
rect 913 4353 927 4367
rect 973 4353 987 4367
rect 1093 4353 1107 4367
rect 653 4253 667 4267
rect 653 4193 667 4207
rect 573 3913 587 3927
rect 833 4253 847 4267
rect 1033 4334 1047 4348
rect 973 4292 987 4306
rect 1013 4292 1027 4306
rect 953 4253 967 4267
rect 993 4253 1007 4267
rect 1053 4253 1067 4267
rect 913 4113 927 4127
rect 673 4073 687 4087
rect 613 3873 627 3887
rect 653 3913 667 3927
rect 573 3813 587 3827
rect 713 4034 727 4048
rect 773 4034 787 4048
rect 813 4034 827 4048
rect 853 4034 867 4048
rect 893 4034 907 4048
rect 753 3973 767 3987
rect 813 3973 827 3987
rect 693 3913 707 3927
rect 733 3913 747 3927
rect 693 3873 707 3887
rect 673 3813 687 3827
rect 593 3772 607 3786
rect 713 3853 727 3867
rect 773 3853 787 3867
rect 933 3973 947 3987
rect 873 3873 887 3887
rect 1113 4113 1127 4127
rect 1053 4034 1067 4048
rect 1013 4013 1027 4027
rect 1033 3993 1047 4007
rect 1013 3953 1027 3967
rect 833 3853 847 3867
rect 993 3853 1007 3867
rect 1053 3853 1067 3867
rect 893 3814 907 3828
rect 953 3813 967 3827
rect 1273 4433 1287 4447
rect 1173 4373 1187 4387
rect 1533 5113 1547 5127
rect 1613 5113 1627 5127
rect 1513 5074 1527 5088
rect 1413 5032 1427 5046
rect 1473 5032 1487 5046
rect 1513 5033 1527 5047
rect 1573 5074 1587 5088
rect 1652 5074 1666 5088
rect 1673 5074 1687 5088
rect 1713 5074 1727 5088
rect 1413 4993 1427 5007
rect 1433 4953 1447 4967
rect 1413 4933 1427 4947
rect 1493 4893 1507 4907
rect 1433 4854 1447 4868
rect 1473 4813 1487 4827
rect 1453 4793 1467 4807
rect 1393 4753 1407 4767
rect 1353 4713 1367 4727
rect 1393 4713 1407 4727
rect 1333 4493 1347 4507
rect 1293 4353 1307 4367
rect 1313 4333 1327 4347
rect 1173 4293 1187 4307
rect 1213 4292 1227 4306
rect 1293 4293 1307 4307
rect 1293 4253 1307 4267
rect 1273 4113 1287 4127
rect 1233 4073 1247 4087
rect 1373 4433 1387 4447
rect 1473 4673 1487 4687
rect 1413 4573 1427 4587
rect 1453 4554 1467 4568
rect 1593 5032 1607 5046
rect 1633 5032 1647 5046
rect 1653 5013 1667 5027
rect 1693 5033 1707 5047
rect 1733 5032 1747 5046
rect 1673 4993 1687 5007
rect 1653 4953 1667 4967
rect 1673 4933 1687 4947
rect 1593 4893 1607 4907
rect 1673 4893 1687 4907
rect 1713 4854 1727 4868
rect 1773 4853 1787 4867
rect 1573 4793 1587 4807
rect 1733 4812 1747 4826
rect 1693 4793 1707 4807
rect 1633 4753 1647 4767
rect 1693 4753 1707 4767
rect 1513 4713 1527 4727
rect 1413 4512 1427 4526
rect 1473 4512 1487 4526
rect 1573 4554 1587 4568
rect 1613 4553 1627 4567
rect 1553 4512 1567 4526
rect 1613 4513 1627 4527
rect 1533 4473 1547 4487
rect 1473 4453 1487 4467
rect 1513 4453 1527 4467
rect 1393 4393 1407 4407
rect 1393 4372 1407 4386
rect 1433 4334 1447 4348
rect 1553 4433 1567 4447
rect 1493 4353 1507 4367
rect 1473 4253 1487 4267
rect 1373 4213 1387 4227
rect 1413 4213 1427 4227
rect 1593 4393 1607 4407
rect 1513 4292 1527 4306
rect 1513 4253 1527 4267
rect 1493 4153 1507 4167
rect 1453 4113 1467 4127
rect 1333 4033 1347 4047
rect 1213 3953 1227 3967
rect 1273 3953 1287 3967
rect 1213 3913 1227 3927
rect 1333 3913 1347 3927
rect 1153 3833 1167 3847
rect 1193 3813 1207 3827
rect 693 3753 707 3767
rect 633 3733 647 3747
rect 573 3593 587 3607
rect 693 3593 707 3607
rect 653 3533 667 3547
rect 833 3772 847 3786
rect 793 3753 807 3767
rect 873 3772 887 3786
rect 893 3753 907 3767
rect 853 3733 867 3747
rect 713 3573 727 3587
rect 773 3514 787 3528
rect 813 3514 827 3528
rect 853 3514 867 3528
rect 953 3772 967 3786
rect 993 3772 1007 3786
rect 913 3733 927 3747
rect 1033 3693 1047 3707
rect 1033 3653 1047 3667
rect 1013 3593 1027 3607
rect 993 3573 1007 3587
rect 933 3553 947 3567
rect 693 3472 707 3486
rect 793 3472 807 3486
rect 753 3433 767 3447
rect 793 3433 807 3447
rect 713 3373 727 3387
rect 593 3353 607 3367
rect 233 3252 247 3266
rect 353 3252 367 3266
rect 353 3193 367 3207
rect 393 3153 407 3167
rect 493 3252 507 3266
rect 533 3252 547 3266
rect 373 3113 387 3127
rect 433 3113 447 3127
rect 153 3013 167 3027
rect 273 3013 287 3027
rect 133 2993 147 3007
rect 213 2994 227 3008
rect 113 2952 127 2966
rect 213 2873 227 2887
rect 53 2853 67 2867
rect 133 2853 147 2867
rect 33 2793 47 2807
rect 13 2773 27 2787
rect 13 2733 27 2747
rect 93 2713 107 2727
rect 33 2673 47 2687
rect 153 2793 167 2807
rect 333 2952 347 2966
rect 593 3293 607 3307
rect 673 3294 687 3308
rect 753 3294 767 3308
rect 613 3252 627 3266
rect 493 3053 507 3067
rect 573 3053 587 3067
rect 393 2993 407 3007
rect 453 2994 467 3008
rect 433 2952 447 2966
rect 393 2913 407 2927
rect 353 2774 367 2788
rect 733 3233 747 3247
rect 953 3472 967 3486
rect 913 3433 927 3447
rect 873 3393 887 3407
rect 853 3373 867 3387
rect 953 3353 967 3367
rect 973 3333 987 3347
rect 1013 3513 1027 3527
rect 1073 3573 1087 3587
rect 1153 3772 1167 3786
rect 1193 3772 1207 3786
rect 1293 3873 1307 3887
rect 1273 3853 1287 3867
rect 1293 3813 1307 3827
rect 1333 3814 1347 3828
rect 1373 4053 1387 4067
rect 1393 4034 1407 4048
rect 1413 3873 1427 3887
rect 1213 3673 1227 3687
rect 1253 3673 1267 3687
rect 1213 3593 1227 3607
rect 1133 3573 1147 3587
rect 1093 3533 1107 3547
rect 1093 3472 1107 3486
rect 1173 3514 1187 3528
rect 1053 3433 1067 3447
rect 1053 3294 1067 3308
rect 1093 3294 1107 3308
rect 973 3253 987 3267
rect 1033 3252 1047 3266
rect 813 3233 827 3247
rect 793 3193 807 3207
rect 853 3193 867 3207
rect 793 3093 807 3107
rect 573 3032 587 3046
rect 673 3033 687 3047
rect 633 2994 647 3008
rect 693 2994 707 3008
rect 733 2994 747 3008
rect 773 2994 787 3008
rect 593 2952 607 2966
rect 633 2953 647 2967
rect 673 2952 687 2966
rect 913 3013 927 3027
rect 853 2994 867 3008
rect 713 2913 727 2927
rect 773 2913 787 2927
rect 493 2793 507 2807
rect 553 2793 567 2807
rect 433 2774 447 2788
rect 473 2773 487 2787
rect 333 2732 347 2746
rect 393 2733 407 2747
rect 453 2732 467 2746
rect 273 2673 287 2687
rect 153 2573 167 2587
rect 193 2573 207 2587
rect 73 2493 87 2507
rect 133 2493 147 2507
rect 73 2474 87 2488
rect 273 2553 287 2567
rect 313 2553 327 2567
rect 373 2553 387 2567
rect 213 2473 227 2487
rect 253 2474 267 2488
rect 873 2953 887 2967
rect 993 3193 1007 3207
rect 1093 3193 1107 3207
rect 1033 3173 1047 3187
rect 993 3013 1007 3027
rect 973 2952 987 2966
rect 1073 3073 1087 3087
rect 1193 3453 1207 3467
rect 1213 3433 1227 3447
rect 1213 3373 1227 3387
rect 1173 3294 1187 3308
rect 1233 3273 1247 3287
rect 1153 3233 1167 3247
rect 1113 3053 1127 3067
rect 1073 2994 1087 3008
rect 1113 2994 1127 3008
rect 913 2933 927 2947
rect 953 2933 967 2947
rect 893 2893 907 2907
rect 893 2793 907 2807
rect 993 2774 1007 2788
rect 573 2732 587 2746
rect 453 2493 467 2507
rect 493 2493 507 2507
rect 553 2493 567 2507
rect 433 2474 447 2488
rect 93 2432 107 2446
rect 133 2432 147 2446
rect 193 2432 207 2446
rect 73 2413 87 2427
rect 113 2293 127 2307
rect 213 2293 227 2307
rect 153 2254 167 2268
rect 192 2254 206 2268
rect 133 2212 147 2226
rect 93 2093 107 2107
rect 113 1973 127 1987
rect 153 1973 167 1987
rect 33 1954 47 1968
rect 73 1954 87 1968
rect 213 2253 227 2267
rect 273 2254 287 2268
rect 393 2254 407 2268
rect 453 2253 467 2267
rect 553 2432 567 2446
rect 673 2673 687 2687
rect 893 2732 907 2746
rect 853 2673 867 2687
rect 773 2533 787 2547
rect 673 2493 687 2507
rect 713 2493 727 2507
rect 613 2473 627 2487
rect 813 2474 827 2488
rect 1213 3213 1227 3227
rect 1373 3814 1387 3828
rect 1453 3833 1467 3847
rect 1593 4273 1607 4287
rect 1573 4233 1587 4247
rect 1713 4673 1727 4687
rect 1773 4793 1787 4807
rect 1853 5074 1867 5088
rect 1973 5332 1987 5346
rect 2093 5413 2107 5427
rect 2153 5373 2167 5387
rect 2053 5332 2067 5346
rect 2113 5293 2127 5307
rect 2033 5273 2047 5287
rect 2073 5273 2087 5287
rect 2053 5193 2067 5207
rect 1993 5133 2007 5147
rect 2013 5113 2027 5127
rect 1993 5093 2007 5107
rect 1973 5074 1987 5088
rect 1913 5052 1927 5066
rect 1833 5013 1847 5027
rect 1933 4913 1947 4927
rect 1833 4873 1847 4887
rect 1913 4873 1927 4887
rect 1793 4713 1807 4727
rect 1753 4553 1767 4567
rect 1793 4554 1807 4568
rect 1833 4573 1847 4587
rect 2113 5032 2127 5046
rect 2032 4913 2046 4927
rect 2053 4913 2067 4927
rect 2093 4913 2107 4927
rect 1933 4833 1947 4847
rect 1933 4793 1947 4807
rect 1913 4753 1927 4767
rect 2073 4753 2087 4767
rect 2053 4693 2067 4707
rect 2013 4593 2027 4607
rect 1993 4573 2007 4587
rect 1733 4533 1747 4547
rect 1773 4512 1787 4526
rect 1693 4473 1707 4487
rect 1633 4193 1647 4207
rect 1733 4213 1747 4227
rect 1933 4554 1947 4568
rect 1953 4512 1967 4526
rect 1993 4513 2007 4527
rect 1933 4473 1947 4487
rect 1913 4353 1927 4367
rect 2633 5433 2647 5447
rect 2573 5413 2587 5427
rect 2613 5413 2627 5427
rect 2593 5393 2607 5407
rect 2633 5393 2647 5407
rect 2193 5374 2207 5388
rect 2453 5374 2467 5388
rect 2553 5374 2567 5388
rect 2173 5333 2187 5347
rect 2233 5332 2247 5346
rect 2193 5213 2207 5227
rect 2333 5332 2347 5346
rect 2573 5332 2587 5346
rect 2493 5293 2507 5307
rect 2633 5293 2647 5307
rect 2273 5193 2287 5207
rect 2433 5133 2447 5147
rect 2353 5113 2367 5127
rect 2393 5113 2407 5127
rect 2373 5093 2387 5107
rect 2233 5074 2247 5088
rect 2293 5074 2307 5088
rect 2333 5074 2347 5088
rect 2213 5032 2227 5046
rect 2253 4993 2267 5007
rect 2193 4913 2207 4927
rect 2233 4913 2247 4927
rect 2353 5032 2367 5046
rect 2393 5032 2407 5046
rect 2333 4893 2347 4907
rect 2293 4854 2307 4868
rect 2233 4812 2247 4826
rect 2273 4812 2287 4826
rect 3253 5473 3267 5487
rect 3293 5473 3307 5487
rect 3033 5453 3047 5467
rect 3233 5453 3247 5467
rect 2733 5433 2747 5447
rect 2873 5433 2887 5447
rect 3013 5433 3027 5447
rect 2713 5413 2727 5427
rect 2693 5374 2707 5388
rect 2813 5413 2827 5427
rect 2793 5393 2807 5407
rect 2713 5332 2727 5346
rect 2753 5332 2767 5346
rect 2673 5293 2687 5307
rect 2653 5253 2667 5267
rect 2593 5173 2607 5187
rect 2493 5074 2507 5088
rect 2553 5073 2567 5087
rect 2693 5193 2707 5207
rect 2633 5074 2647 5088
rect 2673 5074 2687 5088
rect 2513 5032 2527 5046
rect 2433 4993 2447 5007
rect 2473 4993 2487 5007
rect 2513 4953 2527 4967
rect 2473 4913 2487 4927
rect 2413 4893 2427 4907
rect 2373 4854 2387 4868
rect 2753 5133 2767 5147
rect 2873 5332 2887 5346
rect 2853 5253 2867 5267
rect 2813 5193 2827 5207
rect 2813 5153 2827 5167
rect 2793 5073 2807 5087
rect 3013 5333 3027 5347
rect 3133 5413 3147 5427
rect 3213 5413 3227 5427
rect 3193 5393 3207 5407
rect 3093 5374 3107 5388
rect 3133 5374 3147 5388
rect 3193 5374 3207 5388
rect 3113 5313 3127 5327
rect 3153 5353 3167 5367
rect 3033 5293 3047 5307
rect 2953 5253 2967 5267
rect 2993 5253 3007 5267
rect 2913 5193 2927 5207
rect 2613 5032 2627 5046
rect 2693 5032 2707 5046
rect 2773 5032 2787 5046
rect 2813 5032 2827 5046
rect 2873 5013 2887 5027
rect 2653 4993 2667 5007
rect 2733 4993 2747 5007
rect 2793 4993 2807 5007
rect 2633 4953 2647 4967
rect 2753 4953 2767 4967
rect 2553 4873 2567 4887
rect 2593 4873 2607 4887
rect 2473 4854 2487 4868
rect 2533 4854 2547 4868
rect 2433 4812 2447 4826
rect 2173 4773 2187 4787
rect 2333 4773 2347 4787
rect 2133 4753 2147 4767
rect 2253 4753 2267 4767
rect 2093 4633 2107 4647
rect 2133 4633 2147 4647
rect 2093 4593 2107 4607
rect 2053 4554 2067 4568
rect 2193 4554 2207 4568
rect 2233 4554 2247 4568
rect 2073 4512 2087 4526
rect 2233 4473 2247 4487
rect 2373 4593 2387 4607
rect 2313 4512 2327 4526
rect 2353 4512 2367 4526
rect 2453 4733 2467 4747
rect 2553 4773 2567 4787
rect 2473 4713 2487 4727
rect 2513 4713 2527 4727
rect 2693 4893 2707 4907
rect 2633 4793 2647 4807
rect 2493 4653 2507 4667
rect 2593 4653 2607 4667
rect 2433 4512 2447 4526
rect 2373 4493 2387 4507
rect 2353 4473 2367 4487
rect 2413 4473 2427 4487
rect 2433 4433 2447 4447
rect 2333 4393 2347 4407
rect 2133 4373 2147 4387
rect 2253 4373 2267 4387
rect 2293 4373 2307 4387
rect 2013 4353 2027 4367
rect 2073 4353 2087 4367
rect 1893 4273 1907 4287
rect 1773 4213 1787 4227
rect 1873 4213 1887 4227
rect 1753 4173 1767 4187
rect 1693 4153 1707 4167
rect 1653 4113 1667 4127
rect 1573 4073 1587 4087
rect 1613 4034 1627 4048
rect 1753 4073 1767 4087
rect 1713 4034 1727 4048
rect 1753 4034 1767 4048
rect 1513 3993 1527 4007
rect 1553 3992 1567 4006
rect 1593 3992 1607 4006
rect 1753 3913 1767 3927
rect 1593 3893 1607 3907
rect 1973 4253 1987 4267
rect 1893 4034 1907 4048
rect 1933 4034 1947 4048
rect 2033 4213 2047 4227
rect 2013 4193 2027 4207
rect 2013 4034 2027 4048
rect 1813 3913 1827 3927
rect 1613 3873 1627 3887
rect 1773 3873 1787 3887
rect 1593 3853 1607 3867
rect 1333 3773 1347 3787
rect 1313 3573 1327 3587
rect 1273 3533 1287 3547
rect 1313 3533 1327 3547
rect 1533 3814 1547 3828
rect 1513 3772 1527 3786
rect 1553 3772 1567 3786
rect 1593 3773 1607 3787
rect 1573 3713 1587 3727
rect 1513 3693 1527 3707
rect 1533 3693 1547 3707
rect 1493 3633 1507 3647
rect 1433 3514 1447 3528
rect 1473 3514 1487 3528
rect 1393 3393 1407 3407
rect 1293 3333 1307 3347
rect 1333 3294 1347 3308
rect 1313 3252 1327 3266
rect 1393 3252 1407 3266
rect 1453 3252 1467 3266
rect 1253 3193 1267 3207
rect 1293 3193 1307 3207
rect 1353 3193 1367 3207
rect 1213 3173 1227 3187
rect 1273 3053 1287 3067
rect 1193 2994 1207 3008
rect 1233 2994 1247 3008
rect 1173 2953 1187 2967
rect 1093 2933 1107 2947
rect 1153 2933 1167 2947
rect 1133 2893 1147 2907
rect 1093 2793 1107 2807
rect 1033 2773 1047 2787
rect 1253 2952 1267 2966
rect 1213 2853 1227 2867
rect 1233 2833 1247 2847
rect 1273 2833 1287 2847
rect 1193 2793 1207 2807
rect 1133 2773 1147 2787
rect 1173 2773 1187 2787
rect 1033 2732 1047 2746
rect 1073 2732 1087 2746
rect 1113 2732 1127 2746
rect 1173 2733 1187 2747
rect 1013 2653 1027 2667
rect 913 2474 927 2488
rect 953 2474 967 2488
rect 653 2432 667 2446
rect 713 2432 727 2446
rect 753 2432 767 2446
rect 973 2433 987 2447
rect 1093 2533 1107 2547
rect 953 2393 967 2407
rect 1033 2432 1047 2446
rect 1073 2432 1087 2446
rect 613 2373 627 2387
rect 793 2373 807 2387
rect 973 2373 987 2387
rect 1073 2333 1087 2347
rect 613 2293 627 2307
rect 1013 2293 1027 2307
rect 533 2273 547 2287
rect 593 2273 607 2287
rect 573 2254 587 2268
rect 213 2212 227 2226
rect 253 2093 267 2107
rect 13 1893 27 1907
rect 13 1692 27 1706
rect 213 1954 227 1968
rect 253 1954 267 1968
rect 133 1893 147 1907
rect 193 1893 207 1907
rect 453 2173 467 2187
rect 413 2153 427 2167
rect 373 2093 387 2107
rect 373 1954 387 1968
rect 553 2173 567 2187
rect 953 2273 967 2287
rect 653 2254 667 2268
rect 693 2254 707 2268
rect 753 2253 767 2267
rect 793 2254 807 2268
rect 833 2254 847 2268
rect 893 2254 907 2268
rect 673 2193 687 2207
rect 693 2173 707 2187
rect 513 2133 527 2147
rect 613 2133 627 2147
rect 513 2093 527 2107
rect 533 2033 547 2047
rect 412 1953 426 1967
rect 433 1953 447 1967
rect 473 1954 487 1968
rect 393 1912 407 1926
rect 93 1853 107 1867
rect 53 1734 67 1748
rect 173 1734 187 1748
rect 33 1633 47 1647
rect 73 1692 87 1706
rect 73 1633 87 1647
rect 153 1633 167 1647
rect 13 1393 27 1407
rect 73 1493 87 1507
rect 113 1434 127 1448
rect 93 1392 107 1406
rect 33 1353 47 1367
rect 93 1353 107 1367
rect 13 1293 27 1307
rect 33 1233 47 1247
rect 273 1893 287 1907
rect 313 1893 327 1907
rect 213 1853 227 1867
rect 293 1853 307 1867
rect 253 1734 267 1748
rect 373 1833 387 1847
rect 353 1753 367 1767
rect 253 1673 267 1687
rect 213 1633 227 1647
rect 213 1434 227 1448
rect 293 1493 307 1507
rect 173 1393 187 1407
rect 333 1434 347 1448
rect 413 1813 427 1827
rect 573 1954 587 1968
rect 613 1954 627 1968
rect 673 1954 687 1968
rect 813 2212 827 2226
rect 853 2212 867 2226
rect 853 2193 867 2207
rect 813 2173 827 2187
rect 753 2153 767 2167
rect 1153 2474 1167 2488
rect 1213 2732 1227 2746
rect 1253 2713 1267 2727
rect 1333 3113 1347 3127
rect 1593 3573 1607 3587
rect 1593 3514 1607 3528
rect 1513 3393 1527 3407
rect 1553 3393 1567 3407
rect 1853 3993 1867 4007
rect 1833 3853 1847 3867
rect 1893 3913 1907 3927
rect 2033 3993 2047 4007
rect 1993 3953 2007 3967
rect 1953 3893 1967 3907
rect 1973 3853 1987 3867
rect 1873 3814 1887 3828
rect 1933 3814 1947 3828
rect 1973 3814 1987 3828
rect 1733 3693 1747 3707
rect 1713 3633 1727 3647
rect 1633 3593 1647 3607
rect 1613 3453 1627 3467
rect 1733 3613 1747 3627
rect 1773 3613 1787 3627
rect 1713 3573 1727 3587
rect 1653 3514 1667 3528
rect 1753 3472 1767 3486
rect 1773 3393 1787 3407
rect 1873 3713 1887 3727
rect 1833 3693 1847 3707
rect 1953 3772 1967 3786
rect 1913 3753 1927 3767
rect 2013 3773 2027 3787
rect 2053 3953 2067 3967
rect 2193 4292 2207 4306
rect 2233 4173 2247 4187
rect 2233 4113 2247 4127
rect 2173 4034 2187 4048
rect 2273 4093 2287 4107
rect 2313 4334 2327 4348
rect 2312 4293 2326 4307
rect 2393 4334 2407 4348
rect 2433 4334 2447 4348
rect 2533 4554 2547 4568
rect 2553 4473 2567 4487
rect 2593 4473 2607 4487
rect 2653 4753 2667 4767
rect 2653 4673 2667 4687
rect 2733 4812 2747 4826
rect 2733 4773 2747 4787
rect 2833 4854 2847 4868
rect 2893 4893 2907 4907
rect 2933 5133 2947 5147
rect 2973 5133 2987 5147
rect 3013 5133 3027 5147
rect 2993 5113 3007 5127
rect 3073 5113 3087 5127
rect 2953 5073 2967 5087
rect 3033 5074 3047 5088
rect 2933 5013 2947 5027
rect 3013 5032 3027 5046
rect 3313 5393 3327 5407
rect 3353 5374 3367 5388
rect 3413 5373 3427 5387
rect 3773 5413 3787 5427
rect 3833 5413 3847 5427
rect 3973 5413 3987 5427
rect 3733 5373 3747 5387
rect 3773 5374 3787 5388
rect 3893 5374 3907 5388
rect 3213 5313 3227 5327
rect 3153 5233 3167 5247
rect 3253 5173 3267 5187
rect 3173 5113 3187 5127
rect 3152 5074 3166 5088
rect 3173 5073 3187 5087
rect 3133 5032 3147 5046
rect 3172 5033 3186 5047
rect 3073 4953 3087 4967
rect 2973 4933 2987 4947
rect 3133 4913 3147 4927
rect 2953 4893 2967 4907
rect 3073 4893 3087 4907
rect 3113 4893 3127 4907
rect 2913 4853 2927 4867
rect 2893 4812 2907 4826
rect 3013 4854 3027 4868
rect 3053 4854 3067 4868
rect 3093 4853 3107 4867
rect 3133 4854 3147 4868
rect 3193 5032 3207 5046
rect 3193 4973 3207 4987
rect 3253 4973 3267 4987
rect 3173 4853 3187 4867
rect 2853 4793 2867 4807
rect 2793 4753 2807 4767
rect 2773 4713 2787 4727
rect 2693 4633 2707 4647
rect 2653 4593 2667 4607
rect 2713 4593 2727 4607
rect 2673 4553 2687 4567
rect 2733 4573 2747 4587
rect 2653 4513 2667 4527
rect 2593 4452 2607 4466
rect 2633 4453 2647 4467
rect 2533 4393 2547 4407
rect 2333 4292 2347 4306
rect 2373 4292 2387 4306
rect 2413 4233 2427 4247
rect 2393 4213 2407 4227
rect 2293 4073 2307 4087
rect 2273 3992 2287 4006
rect 2233 3973 2247 3987
rect 2053 3893 2067 3907
rect 2133 3893 2147 3907
rect 2093 3814 2107 3828
rect 2153 3814 2167 3828
rect 2193 3814 2207 3828
rect 2073 3772 2087 3786
rect 2053 3753 2067 3767
rect 1933 3733 1947 3747
rect 1993 3733 2007 3747
rect 1893 3673 1907 3687
rect 1833 3514 1847 3528
rect 1873 3514 1887 3528
rect 1853 3472 1867 3486
rect 1853 3453 1867 3467
rect 1813 3393 1827 3407
rect 1713 3373 1727 3387
rect 1793 3373 1807 3387
rect 1633 3333 1647 3347
rect 1733 3333 1747 3347
rect 1613 3252 1627 3266
rect 1673 3252 1687 3266
rect 1513 3193 1527 3207
rect 1573 3173 1587 3187
rect 1493 3093 1507 3107
rect 1333 2994 1347 3008
rect 1473 2993 1487 3007
rect 1513 2994 1527 3008
rect 1493 2933 1507 2947
rect 1473 2913 1487 2927
rect 1353 2893 1367 2907
rect 1393 2893 1407 2907
rect 1493 2893 1507 2907
rect 1793 3213 1807 3227
rect 1693 3113 1707 3127
rect 1633 3073 1647 3087
rect 1853 3373 1867 3387
rect 1833 3293 1847 3307
rect 1813 3053 1827 3067
rect 1833 3033 1847 3047
rect 1913 3472 1927 3486
rect 1893 3353 1907 3367
rect 1993 3633 2007 3647
rect 1993 3514 2007 3528
rect 2133 3773 2147 3787
rect 2113 3733 2127 3747
rect 2273 3813 2287 3827
rect 2153 3733 2167 3747
rect 2133 3693 2147 3707
rect 2073 3673 2087 3687
rect 1933 3413 1947 3427
rect 2013 3472 2027 3486
rect 2053 3413 2067 3427
rect 1973 3373 1987 3387
rect 2253 3772 2267 3786
rect 2353 4034 2367 4048
rect 2313 3953 2327 3967
rect 2333 3913 2347 3927
rect 2373 3873 2387 3887
rect 2313 3813 2327 3827
rect 2513 4292 2527 4306
rect 2473 4093 2487 4107
rect 2453 3992 2467 4006
rect 2453 3973 2467 3987
rect 2433 3913 2447 3927
rect 2413 3814 2427 3828
rect 2333 3772 2347 3786
rect 2393 3753 2407 3767
rect 2373 3733 2387 3747
rect 2293 3713 2307 3727
rect 2333 3713 2347 3727
rect 2413 3673 2427 3687
rect 2393 3613 2407 3627
rect 2213 3593 2227 3607
rect 2333 3593 2347 3607
rect 2133 3514 2147 3528
rect 2173 3514 2187 3528
rect 2233 3514 2247 3528
rect 2273 3514 2287 3528
rect 2313 3514 2327 3528
rect 2073 3393 2087 3407
rect 2013 3353 2027 3367
rect 1873 3294 1887 3308
rect 2013 3294 2027 3308
rect 1973 3252 1987 3266
rect 2033 3133 2047 3147
rect 2073 3133 2087 3147
rect 2013 3053 2027 3067
rect 1893 3033 1907 3047
rect 1633 2952 1647 2966
rect 1673 2952 1687 2966
rect 1693 2933 1707 2947
rect 1713 2913 1727 2927
rect 1853 2994 1867 3008
rect 1953 2994 1967 3008
rect 1693 2893 1707 2907
rect 1773 2893 1787 2907
rect 1613 2853 1627 2867
rect 1413 2793 1427 2807
rect 1493 2793 1507 2807
rect 1333 2774 1347 2788
rect 1393 2774 1407 2788
rect 1633 2793 1647 2807
rect 1533 2773 1547 2787
rect 1593 2774 1607 2788
rect 1653 2773 1667 2787
rect 1693 2774 1707 2788
rect 1733 2774 1747 2788
rect 1773 2774 1787 2788
rect 1413 2732 1427 2746
rect 1393 2713 1407 2727
rect 1293 2693 1307 2707
rect 1353 2693 1367 2707
rect 1253 2533 1267 2547
rect 1193 2474 1207 2488
rect 1293 2474 1307 2488
rect 1133 2432 1147 2446
rect 1193 2433 1207 2447
rect 1233 2432 1247 2446
rect 1313 2432 1327 2446
rect 1533 2713 1547 2727
rect 1613 2732 1627 2746
rect 1652 2732 1666 2746
rect 1713 2732 1727 2746
rect 1673 2713 1687 2727
rect 1653 2693 1667 2707
rect 1573 2673 1587 2687
rect 1473 2653 1487 2667
rect 1793 2593 1807 2607
rect 1733 2553 1747 2567
rect 1393 2533 1407 2547
rect 1733 2493 1747 2507
rect 1433 2474 1447 2488
rect 1492 2474 1506 2488
rect 1513 2474 1527 2488
rect 1473 2453 1487 2467
rect 1413 2432 1427 2446
rect 1433 2413 1447 2427
rect 1473 2413 1487 2427
rect 1273 2393 1287 2407
rect 1353 2393 1367 2407
rect 1253 2373 1267 2387
rect 1293 2373 1307 2387
rect 1093 2293 1107 2307
rect 1193 2274 1207 2288
rect 1113 2254 1127 2268
rect 1193 2253 1207 2267
rect 1233 2254 1247 2268
rect 1293 2254 1307 2268
rect 1373 2254 1387 2268
rect 933 2212 947 2226
rect 1013 2212 1027 2226
rect 1053 2212 1067 2226
rect 1253 2212 1267 2226
rect 1213 2193 1227 2207
rect 933 2173 947 2187
rect 1093 2173 1107 2187
rect 813 2133 827 2147
rect 893 2133 907 2147
rect 853 2093 867 2107
rect 893 2053 907 2067
rect 1073 2053 1087 2067
rect 1213 2053 1227 2067
rect 853 2033 867 2047
rect 713 2013 727 2027
rect 813 2013 827 2027
rect 493 1912 507 1926
rect 533 1912 547 1926
rect 493 1833 507 1847
rect 713 1954 727 1968
rect 753 1954 767 1968
rect 953 2013 967 2027
rect 693 1913 707 1927
rect 673 1853 687 1867
rect 473 1813 487 1827
rect 592 1813 606 1827
rect 613 1813 627 1827
rect 693 1813 707 1827
rect 433 1793 447 1807
rect 433 1753 447 1767
rect 593 1773 607 1787
rect 653 1773 667 1787
rect 513 1734 527 1748
rect 553 1734 567 1748
rect 613 1734 627 1748
rect 813 1913 827 1927
rect 773 1893 787 1907
rect 913 1912 927 1926
rect 1013 1973 1027 1987
rect 1053 1954 1067 1968
rect 1153 1973 1167 1987
rect 1093 1954 1107 1968
rect 1153 1954 1167 1968
rect 993 1912 1007 1926
rect 873 1893 887 1907
rect 953 1893 967 1907
rect 953 1853 967 1867
rect 853 1793 867 1807
rect 493 1693 507 1707
rect 433 1473 447 1487
rect 473 1473 487 1487
rect 573 1692 587 1706
rect 533 1653 547 1667
rect 732 1733 746 1747
rect 753 1733 767 1747
rect 813 1734 827 1748
rect 893 1773 907 1787
rect 853 1733 867 1747
rect 673 1692 687 1706
rect 533 1613 547 1627
rect 613 1613 627 1627
rect 593 1513 607 1527
rect 633 1434 647 1448
rect 153 1333 167 1347
rect 133 1233 147 1247
rect 233 1333 247 1347
rect 193 1293 207 1307
rect 173 1213 187 1227
rect 393 1392 407 1406
rect 273 1214 287 1228
rect 33 1172 47 1186
rect 73 1172 87 1186
rect 113 1172 127 1186
rect 173 1172 187 1186
rect 213 1172 227 1186
rect 13 873 27 887
rect 93 914 107 928
rect 153 933 167 947
rect 293 1172 307 1186
rect 493 1392 507 1406
rect 533 1393 547 1407
rect 573 1392 587 1406
rect 653 1393 667 1407
rect 653 1313 667 1327
rect 713 1673 727 1687
rect 1033 1893 1047 1907
rect 1353 2212 1367 2226
rect 1393 2212 1407 2226
rect 1393 2193 1407 2207
rect 1293 2173 1307 2187
rect 1333 2173 1347 2187
rect 1253 1993 1267 2007
rect 1273 1954 1287 1968
rect 1313 1954 1327 1968
rect 1553 2413 1567 2427
rect 1493 2353 1507 2367
rect 1473 2293 1487 2307
rect 1513 2254 1527 2268
rect 1573 2393 1587 2407
rect 1753 2474 1767 2488
rect 1893 2952 1907 2966
rect 1933 2952 1947 2966
rect 1973 2953 1987 2967
rect 1973 2893 1987 2907
rect 2013 2893 2027 2907
rect 2053 2893 2067 2907
rect 2033 2833 2047 2847
rect 1893 2793 1907 2807
rect 2013 2793 2027 2807
rect 1853 2774 1867 2788
rect 1893 2732 1907 2746
rect 1853 2673 1867 2687
rect 1953 2653 1967 2667
rect 1953 2593 1967 2607
rect 1893 2573 1907 2587
rect 1833 2553 1847 2567
rect 1853 2474 1867 2488
rect 1733 2432 1747 2446
rect 2173 3473 2187 3487
rect 2113 3353 2127 3367
rect 2133 3252 2147 3266
rect 2193 3233 2207 3247
rect 2193 3173 2207 3187
rect 2313 3413 2327 3427
rect 2253 3273 2267 3287
rect 2573 4153 2587 4167
rect 2733 4512 2747 4526
rect 2693 4473 2707 4487
rect 2653 4433 2667 4447
rect 2653 4393 2667 4407
rect 2693 4334 2707 4348
rect 2733 4334 2747 4348
rect 2713 4293 2727 4307
rect 2633 4253 2647 4267
rect 2733 4273 2747 4287
rect 2713 4213 2727 4227
rect 2693 4193 2707 4207
rect 2673 4173 2687 4187
rect 2593 4053 2607 4067
rect 2833 4693 2847 4707
rect 2813 4633 2827 4647
rect 2893 4673 2907 4687
rect 2833 4613 2847 4627
rect 2893 4593 2907 4607
rect 2833 4573 2847 4587
rect 2853 4512 2867 4526
rect 2833 4453 2847 4467
rect 2813 4393 2827 4407
rect 2793 4334 2807 4348
rect 2953 4812 2967 4826
rect 3033 4812 3047 4826
rect 2993 4793 3007 4807
rect 2973 4733 2987 4747
rect 2953 4653 2967 4667
rect 3033 4773 3047 4787
rect 3113 4793 3127 4807
rect 3173 4813 3187 4827
rect 3153 4793 3167 4807
rect 3173 4733 3187 4747
rect 3093 4693 3107 4707
rect 2993 4573 3007 4587
rect 3033 4573 3047 4587
rect 2953 4393 2967 4407
rect 2933 4353 2947 4367
rect 2973 4353 2987 4367
rect 2793 4273 2807 4287
rect 2753 4133 2767 4147
rect 2753 4073 2767 4087
rect 2673 4034 2687 4048
rect 2773 4033 2787 4047
rect 2593 3973 2607 3987
rect 2493 3833 2507 3847
rect 2533 3833 2547 3847
rect 2453 3814 2467 3828
rect 2873 4273 2887 4287
rect 2813 4213 2827 4227
rect 2913 4193 2927 4207
rect 2893 4073 2907 4087
rect 2793 3993 2807 4007
rect 2853 3992 2867 4006
rect 2773 3833 2787 3847
rect 2973 4273 2987 4287
rect 3333 5332 3347 5346
rect 3373 5332 3387 5346
rect 3413 5332 3427 5346
rect 3593 5332 3607 5346
rect 3653 5332 3667 5346
rect 3493 5213 3507 5227
rect 3553 5213 3567 5227
rect 3433 5193 3447 5207
rect 3293 5133 3307 5147
rect 3513 5173 3527 5187
rect 3373 5074 3387 5088
rect 3433 5074 3447 5088
rect 3393 5033 3407 5047
rect 3293 4993 3307 5007
rect 3233 4933 3247 4947
rect 3273 4933 3287 4947
rect 3213 4913 3227 4927
rect 3253 4893 3267 4907
rect 3293 4873 3307 4887
rect 3333 4873 3347 4887
rect 3253 4854 3267 4868
rect 3213 4813 3227 4827
rect 3273 4812 3287 4826
rect 3533 4893 3547 4907
rect 3433 4854 3447 4868
rect 3713 5313 3727 5327
rect 3953 5353 3967 5367
rect 3773 5333 3787 5347
rect 3813 5332 3827 5346
rect 3733 5293 3747 5307
rect 3813 5273 3827 5287
rect 3713 5193 3727 5207
rect 3773 5193 3787 5207
rect 3673 5074 3687 5088
rect 3713 5074 3727 5088
rect 3613 4993 3627 5007
rect 3653 4993 3667 5007
rect 3613 4953 3627 4967
rect 3553 4873 3567 4887
rect 3592 4873 3606 4887
rect 3613 4873 3627 4887
rect 3473 4833 3487 4847
rect 3413 4812 3427 4826
rect 3393 4733 3407 4747
rect 3213 4713 3227 4727
rect 3253 4713 3267 4727
rect 3193 4573 3207 4587
rect 3093 4554 3107 4568
rect 3133 4554 3147 4568
rect 3313 4673 3327 4687
rect 3273 4633 3287 4647
rect 3053 4512 3067 4526
rect 3033 4433 3047 4447
rect 3153 4512 3167 4526
rect 3213 4513 3227 4527
rect 3253 4512 3267 4526
rect 3113 4433 3127 4447
rect 3053 4413 3067 4427
rect 2993 4233 3007 4247
rect 2993 4193 3007 4207
rect 3513 4793 3527 4807
rect 3473 4693 3487 4707
rect 3753 4993 3767 5007
rect 3733 4953 3747 4967
rect 3753 4933 3767 4947
rect 3733 4893 3747 4907
rect 3653 4854 3667 4868
rect 3693 4854 3707 4868
rect 3633 4812 3647 4826
rect 3673 4773 3687 4787
rect 3693 4673 3707 4687
rect 3593 4653 3607 4667
rect 3673 4653 3687 4667
rect 3453 4633 3467 4647
rect 3533 4633 3547 4647
rect 3433 4593 3447 4607
rect 3353 4554 3367 4568
rect 3393 4554 3407 4568
rect 3333 4513 3347 4527
rect 3313 4473 3327 4487
rect 3373 4512 3387 4526
rect 3413 4493 3427 4507
rect 3333 4453 3347 4467
rect 3433 4413 3447 4427
rect 3233 4393 3247 4407
rect 3293 4393 3307 4407
rect 3093 4173 3107 4187
rect 3193 4173 3207 4187
rect 3173 4133 3187 4147
rect 2953 4093 2967 4107
rect 2953 4053 2967 4067
rect 3133 4053 3147 4067
rect 2953 4034 2967 4048
rect 2993 4034 3007 4048
rect 3053 4034 3067 4048
rect 2913 3993 2927 4007
rect 2973 3992 2987 4006
rect 3013 3992 3027 4006
rect 3193 4093 3207 4107
rect 3173 4033 3187 4047
rect 3333 4334 3347 4348
rect 3593 4613 3607 4627
rect 3653 4593 3667 4607
rect 3593 4573 3607 4587
rect 3553 4512 3567 4526
rect 3513 4473 3527 4487
rect 3653 4513 3667 4527
rect 3593 4453 3607 4467
rect 3653 4413 3667 4427
rect 3593 4353 3607 4367
rect 3433 4292 3447 4306
rect 3273 4233 3287 4247
rect 3373 4273 3387 4287
rect 3333 4233 3347 4247
rect 3313 4193 3327 4207
rect 3293 4133 3307 4147
rect 3253 4093 3267 4107
rect 3233 4053 3247 4067
rect 3313 4033 3327 4047
rect 3053 3893 3067 3907
rect 2893 3873 2907 3887
rect 3013 3873 3027 3887
rect 2613 3772 2627 3786
rect 2653 3772 2667 3786
rect 2713 3772 2727 3786
rect 2773 3772 2787 3786
rect 2833 3772 2847 3786
rect 2873 3772 2887 3786
rect 2493 3753 2507 3767
rect 2433 3633 2447 3647
rect 2953 3814 2967 3828
rect 3113 3992 3127 4006
rect 3193 3993 3207 4007
rect 3153 3953 3167 3967
rect 3273 3992 3287 4006
rect 3293 3973 3307 3987
rect 3233 3933 3247 3947
rect 3093 3873 3107 3887
rect 3073 3814 3087 3828
rect 3073 3772 3087 3786
rect 3373 4173 3387 4187
rect 3353 4033 3367 4047
rect 3413 4093 3427 4107
rect 3553 4334 3567 4348
rect 3953 5293 3967 5307
rect 3853 5193 3867 5207
rect 4313 5393 4327 5407
rect 4473 5393 4487 5407
rect 4193 5374 4207 5388
rect 4233 5374 4247 5388
rect 4453 5353 4467 5367
rect 4173 5332 4187 5346
rect 4313 5332 4327 5346
rect 4353 5332 4367 5346
rect 4073 5313 4087 5327
rect 4413 5313 4427 5327
rect 5453 5413 5467 5427
rect 5693 5413 5707 5427
rect 4673 5374 4687 5388
rect 4733 5374 4747 5388
rect 4773 5374 4787 5388
rect 4873 5374 4887 5388
rect 4913 5374 4927 5388
rect 4973 5374 4987 5388
rect 5053 5374 5067 5388
rect 5133 5374 5147 5388
rect 5173 5374 5187 5388
rect 5213 5374 5227 5388
rect 4473 5333 4487 5347
rect 4453 5293 4467 5307
rect 3993 5273 4007 5287
rect 4273 5233 4287 5247
rect 4013 5153 4027 5167
rect 3833 5113 3847 5127
rect 3973 5113 3987 5127
rect 3813 5073 3827 5087
rect 4113 5133 4127 5147
rect 3873 5074 3887 5088
rect 3933 5074 3947 5088
rect 3973 5074 3987 5088
rect 4013 5074 4027 5088
rect 3793 5033 3807 5047
rect 3773 4873 3787 4887
rect 3853 5032 3867 5046
rect 3913 5033 3927 5047
rect 3893 4873 3907 4887
rect 3793 4854 3807 4868
rect 3833 4854 3847 4868
rect 3893 4833 3907 4847
rect 3753 4813 3767 4827
rect 3813 4793 3827 4807
rect 3773 4693 3787 4707
rect 3793 4653 3807 4667
rect 3733 4633 3747 4647
rect 3773 4593 3787 4607
rect 3793 4553 3807 4567
rect 3733 4433 3747 4447
rect 3673 4353 3687 4367
rect 3693 4334 3707 4348
rect 3733 4334 3747 4348
rect 3773 4334 3787 4348
rect 3833 4693 3847 4707
rect 4053 5032 4067 5046
rect 3993 5013 4007 5027
rect 4033 5013 4047 5027
rect 4073 5013 4087 5027
rect 3933 4993 3947 5007
rect 4053 4993 4067 5007
rect 4013 4812 4027 4826
rect 3953 4793 3967 4807
rect 3913 4733 3927 4747
rect 3973 4733 3987 4747
rect 3953 4613 3967 4627
rect 3873 4573 3887 4587
rect 3933 4573 3947 4587
rect 3893 4554 3907 4568
rect 4013 4573 4027 4587
rect 3973 4553 3987 4567
rect 4073 4933 4087 4947
rect 4233 5093 4247 5107
rect 4133 5074 4147 5088
rect 4173 5074 4187 5088
rect 4133 4993 4147 5007
rect 4073 4733 4087 4747
rect 4053 4553 4067 4567
rect 3913 4512 3927 4526
rect 3953 4512 3967 4526
rect 3973 4492 3987 4506
rect 3873 4473 3887 4487
rect 3873 4393 3887 4407
rect 3833 4353 3847 4367
rect 3613 4313 3627 4327
rect 3593 4233 3607 4247
rect 3593 4193 3607 4207
rect 3573 4153 3587 4167
rect 3473 4073 3487 4087
rect 3553 4073 3567 4087
rect 3453 4053 3467 4067
rect 3533 4053 3547 4067
rect 3393 3992 3407 4006
rect 3453 3992 3467 4006
rect 3473 3953 3487 3967
rect 3333 3933 3347 3947
rect 3133 3772 3147 3786
rect 3093 3673 3107 3687
rect 3053 3653 3067 3667
rect 2413 3573 2427 3587
rect 2893 3573 2907 3587
rect 3033 3573 3047 3587
rect 2393 3514 2407 3528
rect 2473 3533 2487 3547
rect 2593 3533 2607 3547
rect 2433 3513 2447 3527
rect 2473 3514 2487 3528
rect 2513 3514 2527 3528
rect 2553 3514 2567 3528
rect 2713 3533 2727 3547
rect 2633 3514 2647 3528
rect 2673 3514 2687 3528
rect 2753 3514 2767 3528
rect 2793 3514 2807 3528
rect 2853 3514 2867 3528
rect 2893 3514 2907 3528
rect 3033 3514 3047 3528
rect 2353 3472 2367 3486
rect 2413 3472 2427 3486
rect 2493 3393 2507 3407
rect 2433 3233 2447 3247
rect 2313 3113 2327 3127
rect 2233 3073 2247 3087
rect 2193 3033 2207 3047
rect 2233 3033 2247 3047
rect 2153 3013 2167 3027
rect 2273 3013 2287 3027
rect 2413 3013 2427 3027
rect 2173 2952 2187 2966
rect 2233 2952 2247 2966
rect 2353 2952 2367 2966
rect 2293 2913 2307 2927
rect 2093 2893 2107 2907
rect 2073 2853 2087 2867
rect 2373 2853 2387 2867
rect 2413 2853 2427 2867
rect 2093 2833 2107 2847
rect 2053 2793 2067 2807
rect 2033 2773 2047 2787
rect 2373 2813 2387 2827
rect 2153 2793 2167 2807
rect 2033 2732 2047 2746
rect 2073 2732 2087 2746
rect 2173 2773 2187 2787
rect 2213 2774 2227 2788
rect 2273 2774 2287 2788
rect 2313 2774 2327 2788
rect 2373 2774 2387 2788
rect 2153 2732 2167 2746
rect 1973 2432 1987 2446
rect 2013 2432 2027 2446
rect 2233 2732 2247 2746
rect 2573 3453 2587 3467
rect 2493 3313 2507 3327
rect 2553 3313 2567 3327
rect 2613 3413 2627 3427
rect 2773 3473 2787 3487
rect 2733 3433 2747 3447
rect 2973 3472 2987 3486
rect 3033 3473 3047 3487
rect 2893 3453 2907 3467
rect 2773 3413 2787 3427
rect 2673 3373 2687 3387
rect 2713 3333 2727 3347
rect 2733 3313 2747 3327
rect 2713 3273 2727 3287
rect 2793 3294 2807 3308
rect 2833 3294 2847 3308
rect 2873 3294 2887 3308
rect 3333 3772 3347 3786
rect 3153 3633 3167 3647
rect 3193 3633 3207 3647
rect 3093 3514 3107 3528
rect 2973 3393 2987 3407
rect 3053 3393 3067 3407
rect 2933 3333 2947 3347
rect 3013 3294 3027 3308
rect 3073 3294 3087 3308
rect 2613 3252 2627 3266
rect 2733 3253 2747 3267
rect 2773 3252 2787 3266
rect 2453 3013 2467 3027
rect 2473 2994 2487 3008
rect 2573 3233 2587 3247
rect 2673 3233 2687 3247
rect 2673 3073 2687 3087
rect 2813 3073 2827 3087
rect 2633 3033 2647 3047
rect 2733 2994 2747 3008
rect 2773 2994 2787 3008
rect 2813 2994 2827 3008
rect 2653 2952 2667 2966
rect 2733 2953 2747 2967
rect 2793 2952 2807 2966
rect 2833 2952 2847 2966
rect 2913 3252 2927 3266
rect 2893 3033 2907 3047
rect 3073 3213 3087 3227
rect 3073 3153 3087 3167
rect 3073 3073 3087 3087
rect 3373 3913 3387 3927
rect 3493 3913 3507 3927
rect 3473 3893 3487 3907
rect 3373 3873 3387 3887
rect 3373 3813 3387 3827
rect 3433 3814 3447 3828
rect 3493 3814 3507 3828
rect 3413 3772 3427 3786
rect 3453 3772 3467 3786
rect 3413 3733 3427 3747
rect 3453 3713 3467 3727
rect 3373 3693 3387 3707
rect 3453 3633 3467 3647
rect 3353 3593 3367 3607
rect 3333 3573 3347 3587
rect 3213 3553 3227 3567
rect 3233 3472 3247 3486
rect 3273 3472 3287 3486
rect 3193 3453 3207 3467
rect 3333 3453 3347 3467
rect 3233 3413 3247 3427
rect 3153 3393 3167 3407
rect 3233 3392 3247 3406
rect 3133 3252 3147 3266
rect 3293 3353 3307 3367
rect 3393 3514 3407 3528
rect 3513 3613 3527 3627
rect 3493 3533 3507 3547
rect 3653 4193 3667 4207
rect 3613 4173 3627 4187
rect 3673 4133 3687 4147
rect 3713 4073 3727 4087
rect 3933 4433 3947 4447
rect 3913 4393 3927 4407
rect 3953 4393 3967 4407
rect 3893 4333 3907 4347
rect 4013 4473 4027 4487
rect 4013 4433 4027 4447
rect 3973 4373 3987 4387
rect 3793 4292 3807 4306
rect 3733 4053 3747 4067
rect 3773 4053 3787 4067
rect 3753 3992 3767 4006
rect 3793 3992 3807 4006
rect 3753 3973 3767 3987
rect 3733 3913 3747 3927
rect 3713 3813 3727 3827
rect 3613 3772 3627 3786
rect 3713 3772 3727 3786
rect 3673 3713 3687 3727
rect 3573 3653 3587 3667
rect 3873 4292 3887 4306
rect 3973 4292 3987 4306
rect 3953 4273 3967 4287
rect 3933 4253 3947 4267
rect 3913 4193 3927 4207
rect 3853 4133 3867 4147
rect 3893 4053 3907 4067
rect 3853 4033 3867 4047
rect 3913 3992 3927 4006
rect 3873 3973 3887 3987
rect 3893 3933 3907 3947
rect 3833 3873 3847 3887
rect 3793 3814 3807 3828
rect 3833 3814 3847 3828
rect 3873 3814 3887 3828
rect 3993 4253 4007 4267
rect 3993 4173 4007 4187
rect 3973 4133 3987 4147
rect 4053 4513 4067 4527
rect 4033 4413 4047 4427
rect 4073 4473 4087 4487
rect 4153 4853 4167 4867
rect 4253 4812 4267 4826
rect 4153 4773 4167 4787
rect 4133 4733 4147 4747
rect 4113 4554 4127 4568
rect 4613 5233 4627 5247
rect 4753 5332 4767 5346
rect 4713 5293 4727 5307
rect 4793 5273 4807 5287
rect 4853 5233 4867 5247
rect 4673 5193 4687 5207
rect 4513 5133 4527 5147
rect 4613 5133 4627 5147
rect 4553 5113 4567 5127
rect 4293 5093 4307 5107
rect 4333 5074 4347 5088
rect 4373 5074 4387 5088
rect 4433 5073 4447 5087
rect 4493 5074 4507 5088
rect 4653 5074 4667 5088
rect 4353 4993 4367 5007
rect 4573 5033 4587 5047
rect 4513 4953 4527 4967
rect 4473 4913 4487 4927
rect 4453 4873 4467 4887
rect 4353 4854 4367 4868
rect 4393 4854 4407 4868
rect 4293 4813 4307 4827
rect 4373 4793 4387 4807
rect 4413 4753 4427 4767
rect 4293 4733 4307 4747
rect 4293 4613 4307 4627
rect 4553 4913 4567 4927
rect 4493 4793 4507 4807
rect 4813 5153 4827 5167
rect 4753 5133 4767 5147
rect 4833 5133 4847 5147
rect 4813 5113 4827 5127
rect 4713 5074 4727 5088
rect 4933 5332 4947 5346
rect 4893 5193 4907 5207
rect 4913 5153 4927 5167
rect 4813 5073 4827 5087
rect 4853 5074 4867 5088
rect 4673 5033 4687 5047
rect 5033 5332 5047 5346
rect 5093 5273 5107 5287
rect 5513 5374 5527 5388
rect 5553 5374 5567 5388
rect 5593 5374 5607 5388
rect 5633 5374 5647 5388
rect 5133 5233 5147 5247
rect 5153 5173 5167 5187
rect 5013 5093 5027 5107
rect 5113 5093 5127 5107
rect 4953 5074 4967 5088
rect 4773 5032 4787 5046
rect 4813 5032 4827 5046
rect 4873 5032 4887 5046
rect 4912 5032 4926 5046
rect 4933 5033 4947 5047
rect 5073 5074 5087 5088
rect 5113 5074 5127 5088
rect 5233 5332 5247 5346
rect 5313 5332 5327 5346
rect 5373 5333 5387 5347
rect 5373 5173 5387 5187
rect 5473 5153 5487 5167
rect 5193 5133 5207 5147
rect 5573 5332 5587 5346
rect 5633 5332 5647 5346
rect 5673 5332 5687 5346
rect 5453 5113 5467 5127
rect 5513 5113 5527 5127
rect 5213 5074 5227 5088
rect 5273 5073 5287 5087
rect 5333 5074 5347 5088
rect 5393 5074 5407 5088
rect 5493 5074 5507 5088
rect 5533 5074 5547 5088
rect 5593 5074 5607 5088
rect 4733 4993 4747 5007
rect 4653 4933 4667 4947
rect 4593 4913 4607 4927
rect 4613 4893 4627 4907
rect 4573 4873 4587 4887
rect 4693 4893 4707 4907
rect 4773 4893 4787 4907
rect 4733 4873 4747 4887
rect 4913 4993 4927 5007
rect 4913 4933 4927 4947
rect 4813 4873 4827 4887
rect 4553 4753 4567 4767
rect 4453 4713 4467 4727
rect 4493 4713 4507 4727
rect 4473 4653 4487 4667
rect 4453 4613 4467 4627
rect 4413 4593 4427 4607
rect 4353 4554 4367 4568
rect 4393 4554 4407 4568
rect 4433 4554 4447 4568
rect 4213 4512 4227 4526
rect 4093 4433 4107 4447
rect 4113 4393 4127 4407
rect 4113 4353 4127 4367
rect 4133 4334 4147 4348
rect 4093 4292 4107 4306
rect 4053 4273 4067 4287
rect 4093 4253 4107 4267
rect 4033 4233 4047 4247
rect 4013 4153 4027 4167
rect 3993 4093 4007 4107
rect 3973 4073 3987 4087
rect 3973 4033 3987 4047
rect 4053 4113 4067 4127
rect 4153 4113 4167 4127
rect 4033 4034 4047 4048
rect 4073 4034 4087 4048
rect 4413 4512 4427 4526
rect 4313 4473 4327 4487
rect 4353 4473 4367 4487
rect 4373 4453 4387 4467
rect 4253 4292 4267 4306
rect 4313 4273 4327 4287
rect 4513 4633 4527 4647
rect 4672 4813 4686 4827
rect 4693 4813 4707 4827
rect 4633 4793 4647 4807
rect 4673 4773 4687 4787
rect 4753 4773 4767 4787
rect 4873 4812 4887 4826
rect 4633 4733 4647 4747
rect 4813 4733 4827 4747
rect 4573 4613 4587 4627
rect 4593 4593 4607 4607
rect 4472 4453 4486 4467
rect 4493 4453 4507 4467
rect 4533 4512 4547 4526
rect 4573 4512 4587 4526
rect 4613 4513 4627 4527
rect 4573 4473 4587 4487
rect 4593 4453 4607 4467
rect 4493 4393 4507 4407
rect 4413 4253 4427 4267
rect 4373 4233 4387 4247
rect 4493 4292 4507 4306
rect 4493 4273 4507 4287
rect 4453 4213 4467 4227
rect 4213 4133 4227 4147
rect 4313 4133 4327 4147
rect 4293 4073 4307 4087
rect 3953 3953 3967 3967
rect 3933 3933 3947 3947
rect 3973 3933 3987 3947
rect 3953 3913 3967 3927
rect 4053 3993 4067 4007
rect 3913 3873 3927 3887
rect 3953 3833 3967 3847
rect 3813 3713 3827 3727
rect 3773 3693 3787 3707
rect 3913 3814 3927 3828
rect 4193 4013 4207 4027
rect 4133 3933 4147 3947
rect 4173 3933 4187 3947
rect 4013 3893 4027 3907
rect 4053 3893 4067 3907
rect 3993 3813 4007 3827
rect 4073 3853 4087 3867
rect 3873 3733 3887 3747
rect 3833 3693 3847 3707
rect 3813 3673 3827 3687
rect 3733 3573 3747 3587
rect 3573 3553 3587 3567
rect 3653 3553 3667 3567
rect 3713 3553 3727 3567
rect 3773 3553 3787 3567
rect 3553 3533 3567 3547
rect 3613 3514 3627 3528
rect 3553 3472 3567 3486
rect 3513 3453 3527 3467
rect 3493 3333 3507 3347
rect 3553 3413 3567 3427
rect 3353 3313 3367 3327
rect 3393 3313 3407 3327
rect 3513 3313 3527 3327
rect 3333 3294 3347 3308
rect 3353 3252 3367 3266
rect 2933 2994 2947 3008
rect 2993 2993 3007 3007
rect 3033 2994 3047 3008
rect 3293 3193 3307 3207
rect 3233 3013 3247 3027
rect 3153 2994 3167 3008
rect 3193 2994 3207 3008
rect 2893 2952 2907 2966
rect 2693 2913 2707 2927
rect 2753 2913 2767 2927
rect 2873 2913 2887 2927
rect 2473 2853 2487 2867
rect 2473 2774 2487 2788
rect 2613 2773 2627 2787
rect 2653 2774 2667 2788
rect 2593 2753 2607 2767
rect 2493 2732 2507 2746
rect 2433 2713 2447 2727
rect 2453 2713 2467 2727
rect 2553 2713 2567 2727
rect 2613 2713 2627 2727
rect 2273 2693 2287 2707
rect 2333 2693 2347 2707
rect 2193 2673 2207 2687
rect 2453 2653 2467 2667
rect 2333 2613 2347 2627
rect 2093 2513 2107 2527
rect 2133 2474 2147 2488
rect 2173 2474 2187 2488
rect 2233 2474 2247 2488
rect 1913 2413 1927 2427
rect 1833 2353 1847 2367
rect 1893 2353 1907 2367
rect 1673 2333 1687 2347
rect 1573 2293 1587 2307
rect 1633 2293 1647 2307
rect 1753 2293 1767 2307
rect 1813 2293 1827 2307
rect 1553 2253 1567 2267
rect 1493 2212 1507 2226
rect 1533 2173 1547 2187
rect 1453 2013 1467 2027
rect 1413 1954 1427 1968
rect 1453 1954 1467 1968
rect 1493 1954 1507 1968
rect 1633 2254 1647 2268
rect 1613 2173 1627 2187
rect 1653 2113 1667 2127
rect 1573 2053 1587 2067
rect 1633 2013 1647 2027
rect 1353 1933 1367 1947
rect 1093 1833 1107 1847
rect 993 1773 1007 1787
rect 993 1734 1007 1748
rect 1033 1734 1047 1748
rect 1073 1734 1087 1748
rect 1133 1873 1147 1887
rect 1173 1873 1187 1887
rect 1213 1873 1227 1887
rect 753 1573 767 1587
rect 833 1692 847 1706
rect 893 1692 907 1706
rect 933 1692 947 1706
rect 833 1633 847 1647
rect 793 1553 807 1567
rect 753 1473 767 1487
rect 813 1473 827 1487
rect 713 1434 727 1448
rect 693 1393 707 1407
rect 693 1353 707 1367
rect 673 1293 687 1307
rect 613 1273 627 1287
rect 533 1253 547 1267
rect 593 1233 607 1247
rect 373 1214 387 1228
rect 413 1214 427 1228
rect 453 1214 467 1228
rect 493 1214 507 1228
rect 533 1214 547 1228
rect 333 1153 347 1167
rect 253 1113 267 1127
rect 253 933 267 947
rect 253 914 267 928
rect 313 914 327 928
rect 433 1153 447 1167
rect 413 1013 427 1027
rect 73 872 87 886
rect 133 853 147 867
rect 113 773 127 787
rect 73 733 87 747
rect 153 813 167 827
rect 173 793 187 807
rect 213 853 227 867
rect 193 773 207 787
rect 233 793 247 807
rect 273 793 287 807
rect 373 914 387 928
rect 412 914 426 928
rect 553 1172 567 1186
rect 453 1113 467 1127
rect 493 1113 507 1127
rect 433 913 447 927
rect 333 873 347 887
rect 333 813 347 827
rect 213 733 227 747
rect 153 693 167 707
rect 233 694 247 708
rect 93 652 107 666
rect 133 653 147 667
rect 173 652 187 666
rect 213 652 227 666
rect 253 653 267 667
rect 393 872 407 886
rect 653 1233 667 1247
rect 613 1213 627 1227
rect 733 1293 747 1307
rect 1033 1633 1047 1647
rect 1133 1692 1147 1706
rect 1213 1833 1227 1847
rect 1293 1912 1307 1926
rect 1313 1893 1327 1907
rect 1273 1833 1287 1847
rect 1253 1793 1267 1807
rect 1233 1734 1247 1748
rect 1293 1793 1307 1807
rect 1433 1873 1447 1887
rect 1413 1853 1427 1867
rect 1353 1833 1367 1847
rect 1313 1753 1327 1767
rect 1293 1733 1307 1747
rect 1133 1673 1147 1687
rect 973 1613 987 1627
rect 1093 1613 1107 1627
rect 953 1573 967 1587
rect 1113 1573 1127 1587
rect 913 1493 927 1507
rect 833 1433 847 1447
rect 873 1434 887 1448
rect 833 1393 847 1407
rect 853 1373 867 1387
rect 813 1273 827 1287
rect 773 1253 787 1267
rect 733 1213 747 1227
rect 773 1214 787 1228
rect 853 1313 867 1327
rect 933 1353 947 1367
rect 933 1313 947 1327
rect 893 1273 907 1287
rect 853 1213 867 1227
rect 673 1113 687 1127
rect 633 1093 647 1107
rect 833 1172 847 1186
rect 1073 1493 1087 1507
rect 1013 1473 1027 1487
rect 993 1373 1007 1387
rect 1153 1473 1167 1487
rect 1253 1692 1267 1706
rect 1393 1693 1407 1707
rect 1213 1653 1227 1667
rect 1313 1653 1327 1667
rect 1473 1853 1487 1867
rect 1533 1873 1547 1887
rect 1493 1813 1507 1827
rect 1473 1753 1487 1767
rect 1433 1733 1447 1747
rect 1333 1633 1347 1647
rect 1413 1633 1427 1647
rect 1273 1513 1287 1527
rect 1233 1434 1247 1448
rect 1313 1473 1327 1487
rect 1213 1393 1227 1407
rect 1093 1373 1107 1387
rect 1133 1373 1147 1387
rect 1193 1373 1207 1387
rect 1073 1353 1087 1367
rect 1033 1293 1047 1307
rect 1033 1233 1047 1247
rect 1073 1233 1087 1247
rect 913 1172 927 1186
rect 633 993 647 1007
rect 733 993 747 1007
rect 513 953 527 967
rect 693 953 707 967
rect 873 953 887 967
rect 593 932 607 946
rect 633 933 647 947
rect 553 914 567 928
rect 373 853 387 867
rect 413 853 427 867
rect 453 853 467 867
rect 353 753 367 767
rect 313 713 327 727
rect 353 713 367 727
rect 333 694 347 708
rect 393 753 407 767
rect 153 473 167 487
rect 113 394 127 408
rect 533 872 547 886
rect 653 914 667 928
rect 693 914 707 928
rect 733 914 747 928
rect 793 914 807 928
rect 833 914 847 928
rect 553 853 567 867
rect 593 853 607 867
rect 493 793 507 807
rect 453 713 467 727
rect 493 713 507 727
rect 533 653 547 667
rect 513 613 527 627
rect 413 553 427 567
rect 253 493 267 507
rect 413 493 427 507
rect 513 493 527 507
rect 193 473 207 487
rect 173 393 187 407
rect 33 353 47 367
rect 93 352 107 366
rect 113 333 127 347
rect 113 293 127 307
rect 93 253 107 267
rect 133 253 147 267
rect 213 433 227 447
rect 333 433 347 447
rect 293 394 307 408
rect 233 352 247 366
rect 253 333 267 347
rect 213 313 227 327
rect 333 353 347 367
rect 313 333 327 347
rect 273 313 287 327
rect 453 394 467 408
rect 493 394 507 408
rect 593 813 607 827
rect 673 872 687 886
rect 673 833 687 847
rect 693 813 707 827
rect 633 753 647 767
rect 753 873 767 887
rect 733 793 747 807
rect 753 733 767 747
rect 693 713 707 727
rect 633 694 647 708
rect 673 694 687 708
rect 653 652 667 666
rect 853 813 867 827
rect 813 793 827 807
rect 833 753 847 767
rect 813 733 827 747
rect 713 693 727 707
rect 753 694 767 708
rect 793 694 807 708
rect 553 633 567 647
rect 613 633 627 647
rect 693 652 707 666
rect 733 633 747 647
rect 673 613 687 627
rect 973 952 987 966
rect 933 914 947 928
rect 893 873 907 887
rect 1073 1133 1087 1147
rect 953 872 967 886
rect 1013 872 1027 886
rect 913 833 927 847
rect 893 793 907 807
rect 873 753 887 767
rect 853 733 867 747
rect 973 773 987 787
rect 1013 713 1027 727
rect 1193 1293 1207 1307
rect 1253 1353 1267 1367
rect 1213 1273 1227 1287
rect 1193 1233 1207 1247
rect 1153 1214 1167 1228
rect 1113 1172 1127 1186
rect 1193 1093 1207 1107
rect 1373 1533 1387 1547
rect 1493 1692 1507 1706
rect 1593 1913 1607 1927
rect 1773 2212 1787 2226
rect 1813 2212 1827 2226
rect 1733 2153 1747 2167
rect 1693 2013 1707 2027
rect 1673 1973 1687 1987
rect 1653 1954 1667 1968
rect 1873 2293 1887 2307
rect 1833 2193 1847 2207
rect 1773 2113 1787 2127
rect 1833 2093 1847 2107
rect 1753 2053 1767 2067
rect 1733 1973 1747 1987
rect 1833 2033 1847 2047
rect 1913 2193 1927 2207
rect 1893 2013 1907 2027
rect 1833 1954 1847 1968
rect 1873 1954 1887 1968
rect 1993 2254 2007 2268
rect 1993 2193 2007 2207
rect 1933 2153 1947 2167
rect 1973 2153 1987 2167
rect 1973 1993 1987 2007
rect 1913 1973 1927 1987
rect 1613 1873 1627 1887
rect 1553 1833 1567 1847
rect 1593 1833 1607 1847
rect 1673 1912 1687 1926
rect 1713 1912 1727 1926
rect 1753 1912 1767 1926
rect 1813 1912 1827 1926
rect 1833 1893 1847 1907
rect 1873 1893 1887 1907
rect 1673 1873 1687 1887
rect 1753 1873 1767 1887
rect 1653 1833 1667 1847
rect 1633 1793 1647 1807
rect 1593 1734 1607 1748
rect 1453 1493 1467 1507
rect 1413 1473 1427 1487
rect 1573 1692 1587 1706
rect 1693 1753 1707 1767
rect 1673 1734 1687 1748
rect 1533 1673 1547 1687
rect 1573 1613 1587 1627
rect 1533 1533 1547 1547
rect 1553 1473 1567 1487
rect 1473 1434 1487 1448
rect 1513 1434 1527 1448
rect 1593 1573 1607 1587
rect 1333 1373 1347 1387
rect 1273 1333 1287 1347
rect 1313 1333 1327 1347
rect 1253 1233 1267 1247
rect 1273 1214 1287 1228
rect 1393 1392 1407 1406
rect 1373 1373 1387 1387
rect 1353 1213 1367 1227
rect 1253 1172 1267 1186
rect 1333 1172 1347 1186
rect 1313 1133 1327 1147
rect 1293 1113 1307 1127
rect 1273 993 1287 1007
rect 1253 973 1267 987
rect 1093 913 1107 927
rect 1133 914 1147 928
rect 1113 853 1127 867
rect 1293 893 1307 907
rect 1233 853 1247 867
rect 1173 773 1187 787
rect 1293 773 1307 787
rect 1072 753 1086 767
rect 1093 753 1107 767
rect 1153 753 1167 767
rect 1053 733 1067 747
rect 1033 693 1047 707
rect 933 673 947 687
rect 833 633 847 647
rect 873 633 887 647
rect 953 653 967 667
rect 933 613 947 627
rect 773 593 787 607
rect 813 593 827 607
rect 773 473 787 487
rect 853 473 867 487
rect 773 433 787 447
rect 533 413 547 427
rect 633 413 647 427
rect 673 413 687 427
rect 573 394 587 408
rect 393 352 407 366
rect 353 313 367 327
rect 413 313 427 327
rect 313 293 327 307
rect 433 293 447 307
rect 473 293 487 307
rect 453 273 467 287
rect 433 253 447 267
rect 433 213 447 227
rect 353 174 367 188
rect 553 333 567 347
rect 593 333 607 347
rect 613 313 627 327
rect 593 293 607 307
rect 573 273 587 287
rect 493 193 507 207
rect 533 173 547 187
rect 713 394 727 408
rect 753 353 767 367
rect 693 313 707 327
rect 733 313 747 327
rect 753 233 767 247
rect 693 213 707 227
rect 733 213 747 227
rect 633 193 647 207
rect 213 132 227 146
rect 253 133 267 147
rect 293 132 307 146
rect 113 93 127 107
rect 333 93 347 107
rect 493 93 507 107
rect 573 132 587 146
rect 613 132 627 146
rect 693 173 707 187
rect 1133 733 1147 747
rect 1433 1333 1447 1347
rect 1393 1213 1407 1227
rect 1533 1392 1547 1406
rect 1533 1313 1547 1327
rect 1673 1613 1687 1627
rect 1653 1593 1667 1607
rect 1753 1734 1767 1748
rect 1793 1734 1807 1748
rect 1713 1673 1727 1687
rect 1693 1573 1707 1587
rect 1653 1553 1667 1567
rect 1773 1493 1787 1507
rect 1813 1673 1827 1687
rect 1913 1893 1927 1907
rect 1893 1853 1907 1867
rect 1853 1793 1867 1807
rect 1873 1653 1887 1667
rect 1853 1553 1867 1567
rect 1633 1473 1647 1487
rect 1793 1473 1807 1487
rect 1653 1434 1667 1448
rect 1693 1434 1707 1448
rect 1733 1434 1747 1448
rect 1773 1434 1787 1448
rect 1813 1434 1827 1448
rect 1853 1434 1867 1448
rect 1673 1313 1687 1327
rect 1553 1293 1567 1307
rect 1593 1293 1607 1307
rect 1473 1253 1487 1267
rect 1473 1214 1487 1228
rect 1373 1153 1387 1167
rect 1433 1153 1447 1167
rect 1413 1093 1427 1107
rect 1393 1053 1407 1067
rect 1393 914 1407 928
rect 1353 853 1367 867
rect 1333 813 1347 827
rect 1233 733 1247 747
rect 1313 733 1327 747
rect 1213 693 1227 707
rect 1113 652 1127 666
rect 1153 652 1167 666
rect 1053 633 1067 647
rect 1093 633 1107 647
rect 993 593 1007 607
rect 1053 553 1067 567
rect 1013 493 1027 507
rect 973 453 987 467
rect 953 433 967 447
rect 853 413 867 427
rect 872 394 886 408
rect 893 393 907 407
rect 1013 394 1027 408
rect 853 352 867 366
rect 993 352 1007 366
rect 953 313 967 327
rect 813 293 827 307
rect 993 293 1007 307
rect 1153 613 1167 627
rect 1193 593 1207 607
rect 1113 533 1127 547
rect 1193 453 1207 467
rect 1133 433 1147 447
rect 1093 413 1107 427
rect 1333 713 1347 727
rect 1413 873 1427 887
rect 1453 1133 1467 1147
rect 1493 1132 1507 1146
rect 1493 1093 1507 1107
rect 1793 1392 1807 1406
rect 1833 1392 1847 1406
rect 1813 1353 1827 1367
rect 1753 1293 1767 1307
rect 1733 1273 1747 1287
rect 1673 1253 1687 1267
rect 1553 1213 1567 1227
rect 1593 1214 1607 1228
rect 1653 1214 1667 1228
rect 1573 1172 1587 1186
rect 1573 1113 1587 1127
rect 1512 1053 1526 1067
rect 1533 1053 1547 1067
rect 1493 1033 1507 1047
rect 1473 973 1487 987
rect 1553 913 1567 927
rect 1513 872 1527 886
rect 1473 853 1487 867
rect 1633 1133 1647 1147
rect 1693 1172 1707 1186
rect 1653 1113 1667 1127
rect 1673 973 1687 987
rect 1593 913 1607 927
rect 1593 872 1607 886
rect 1653 872 1667 886
rect 1433 833 1447 847
rect 1533 833 1547 847
rect 1573 833 1587 847
rect 1413 813 1427 827
rect 1513 813 1527 827
rect 1373 773 1387 787
rect 1413 753 1427 767
rect 1473 753 1487 767
rect 1393 733 1407 747
rect 1273 694 1287 708
rect 1313 694 1327 708
rect 1352 694 1366 708
rect 1373 694 1387 708
rect 1233 652 1247 666
rect 1293 652 1307 666
rect 1433 694 1447 708
rect 1273 573 1287 587
rect 1333 513 1347 527
rect 1273 433 1287 447
rect 1173 393 1187 407
rect 1333 413 1347 427
rect 1053 273 1067 287
rect 893 253 907 267
rect 1033 253 1047 267
rect 853 233 867 247
rect 813 193 827 207
rect 713 132 727 146
rect 1033 213 1047 227
rect 993 193 1007 207
rect 1153 352 1167 366
rect 1173 313 1187 327
rect 1153 253 1167 267
rect 1093 173 1107 187
rect 1173 173 1187 187
rect 1293 352 1307 366
rect 1253 333 1267 347
rect 1313 273 1327 287
rect 1373 413 1387 427
rect 1353 393 1367 407
rect 1453 652 1467 666
rect 1493 652 1507 666
rect 1493 613 1507 627
rect 1492 553 1506 567
rect 1513 553 1527 567
rect 1713 1053 1727 1067
rect 1713 953 1727 967
rect 1573 793 1587 807
rect 1693 793 1707 807
rect 1733 913 1747 927
rect 1773 833 1787 847
rect 1793 773 1807 787
rect 1673 753 1687 767
rect 1713 753 1727 767
rect 1773 753 1787 767
rect 1573 733 1587 747
rect 1613 733 1627 747
rect 1593 652 1607 666
rect 1633 652 1647 666
rect 1753 733 1767 747
rect 1773 713 1787 727
rect 1793 693 1807 707
rect 1733 652 1747 666
rect 1773 652 1787 666
rect 1673 593 1687 607
rect 1653 573 1667 587
rect 1733 613 1747 627
rect 1713 573 1727 587
rect 1733 533 1747 547
rect 1593 493 1607 507
rect 1673 493 1687 507
rect 1613 473 1627 487
rect 1593 433 1607 447
rect 1553 413 1567 427
rect 1413 394 1427 408
rect 1473 393 1487 407
rect 1513 394 1527 408
rect 1393 352 1407 366
rect 1433 352 1447 366
rect 1413 313 1427 327
rect 1433 293 1447 307
rect 1413 273 1427 287
rect 1332 253 1346 267
rect 1353 253 1367 267
rect 1393 253 1407 267
rect 1233 213 1247 227
rect 1333 213 1347 227
rect 1273 193 1287 207
rect 1453 233 1467 247
rect 1433 213 1447 227
rect 1353 173 1367 187
rect 1413 174 1427 188
rect 1493 313 1507 327
rect 1493 273 1507 287
rect 1713 394 1727 408
rect 1953 1813 1967 1827
rect 1933 1734 1947 1748
rect 1993 1734 2007 1748
rect 2033 2053 2047 2067
rect 2033 2032 2047 2046
rect 2033 1913 2047 1927
rect 2033 1793 2047 1807
rect 1913 1653 1927 1667
rect 1893 1613 1907 1627
rect 1873 1353 1887 1367
rect 1913 1473 1927 1487
rect 1973 1673 1987 1687
rect 1993 1653 2007 1667
rect 1973 1573 1987 1587
rect 1973 1473 1987 1487
rect 1933 1453 1947 1467
rect 1913 1373 1927 1387
rect 1893 1333 1907 1347
rect 1953 1353 1967 1367
rect 1953 1293 1967 1307
rect 2013 1613 2027 1627
rect 2173 2433 2187 2447
rect 2113 2413 2127 2427
rect 2073 2373 2087 2387
rect 2173 2373 2187 2387
rect 2093 2353 2107 2367
rect 2073 2313 2087 2327
rect 2093 2273 2107 2287
rect 2113 2254 2127 2268
rect 2093 2212 2107 2226
rect 2213 2432 2227 2446
rect 2273 2432 2287 2446
rect 2233 2413 2247 2427
rect 2353 2474 2367 2488
rect 2393 2474 2407 2488
rect 2493 2573 2507 2587
rect 2353 2433 2367 2447
rect 2713 2732 2727 2746
rect 2673 2693 2687 2707
rect 2953 2873 2967 2887
rect 2973 2813 2987 2827
rect 2913 2793 2927 2807
rect 2953 2793 2967 2807
rect 2773 2773 2787 2787
rect 2833 2774 2847 2788
rect 2893 2773 2907 2787
rect 2773 2732 2787 2746
rect 2853 2732 2867 2746
rect 2893 2732 2907 2746
rect 2813 2713 2827 2727
rect 3053 2952 3067 2966
rect 3153 2953 3167 2967
rect 3093 2913 3107 2927
rect 2993 2773 3007 2787
rect 3253 2913 3267 2927
rect 3313 3113 3327 3127
rect 3453 3294 3467 3308
rect 3493 3294 3507 3308
rect 3433 3213 3447 3227
rect 3433 3173 3447 3187
rect 3393 3033 3407 3047
rect 3393 2952 3407 2966
rect 3313 2933 3327 2947
rect 3353 2933 3367 2947
rect 3333 2813 3347 2827
rect 3213 2773 3227 2787
rect 3133 2732 3147 2746
rect 3193 2732 3207 2746
rect 3273 2732 3287 2746
rect 3093 2693 3107 2707
rect 3033 2633 3047 2647
rect 3193 2633 3207 2647
rect 2933 2613 2947 2627
rect 2913 2533 2927 2547
rect 2973 2533 2987 2547
rect 2613 2513 2627 2527
rect 2653 2513 2667 2527
rect 2693 2513 2707 2527
rect 2753 2513 2767 2527
rect 2513 2474 2527 2488
rect 2553 2474 2567 2488
rect 2593 2474 2607 2488
rect 2733 2474 2747 2488
rect 2773 2473 2787 2487
rect 2813 2474 2827 2488
rect 2973 2493 2987 2507
rect 2933 2474 2947 2488
rect 3153 2593 3167 2607
rect 3133 2573 3147 2587
rect 3133 2513 3147 2527
rect 3093 2474 3107 2488
rect 3133 2473 3147 2487
rect 2573 2432 2587 2446
rect 2613 2432 2627 2446
rect 2653 2432 2667 2446
rect 2513 2393 2527 2407
rect 2713 2393 2727 2407
rect 2333 2373 2347 2387
rect 2373 2373 2387 2387
rect 2493 2373 2507 2387
rect 2573 2373 2587 2387
rect 2333 2333 2347 2347
rect 2273 2313 2287 2327
rect 2413 2293 2427 2307
rect 2473 2253 2487 2267
rect 2533 2254 2547 2268
rect 2593 2353 2607 2367
rect 2833 2432 2847 2446
rect 2893 2433 2907 2447
rect 2873 2333 2887 2347
rect 2673 2293 2687 2307
rect 2773 2293 2787 2307
rect 2833 2293 2847 2307
rect 2572 2253 2586 2267
rect 2593 2254 2607 2268
rect 2653 2253 2667 2267
rect 2193 2212 2207 2226
rect 2133 2193 2147 2207
rect 2173 2193 2187 2207
rect 2093 2173 2107 2187
rect 2173 2133 2187 2147
rect 2113 2113 2127 2127
rect 2073 1993 2087 2007
rect 2133 2073 2147 2087
rect 2253 2153 2267 2167
rect 2133 2033 2147 2047
rect 2193 2033 2207 2047
rect 2233 2033 2247 2047
rect 2153 2013 2167 2027
rect 2113 1793 2127 1807
rect 2133 1773 2147 1787
rect 2193 2012 2207 2026
rect 2213 1912 2227 1926
rect 2173 1773 2187 1787
rect 2113 1734 2127 1748
rect 2153 1734 2167 1748
rect 2053 1653 2067 1667
rect 2133 1692 2147 1706
rect 2233 1853 2247 1867
rect 2313 2213 2327 2227
rect 2293 1953 2307 1967
rect 2433 2212 2447 2226
rect 2473 2212 2487 2226
rect 2433 2173 2447 2187
rect 2413 2133 2427 2147
rect 2393 2073 2407 2087
rect 2313 1893 2327 1907
rect 2273 1773 2287 1787
rect 2253 1753 2267 1767
rect 2373 1912 2387 1926
rect 2553 2212 2567 2226
rect 2553 2173 2567 2187
rect 2593 2173 2607 2187
rect 2513 2133 2527 2147
rect 2553 2113 2567 2127
rect 2553 2073 2567 2087
rect 2453 2033 2467 2047
rect 2493 1954 2507 1968
rect 2533 1954 2547 1968
rect 2813 2273 2827 2287
rect 2673 2212 2687 2226
rect 2713 2212 2727 2226
rect 2673 2153 2687 2167
rect 2653 1973 2667 1987
rect 2633 1954 2647 1968
rect 2333 1853 2347 1867
rect 2353 1793 2367 1807
rect 2333 1753 2347 1767
rect 2173 1693 2187 1707
rect 2173 1613 2187 1627
rect 2073 1573 2087 1587
rect 2113 1553 2127 1567
rect 2033 1513 2047 1527
rect 2033 1492 2047 1506
rect 2073 1434 2087 1448
rect 2133 1453 2147 1467
rect 2013 1393 2027 1407
rect 1993 1373 2007 1387
rect 1853 1172 1867 1186
rect 1833 1153 1847 1167
rect 1893 1113 1907 1127
rect 1853 973 1867 987
rect 2053 1313 2067 1327
rect 2093 1313 2107 1327
rect 2253 1692 2267 1706
rect 2293 1692 2307 1706
rect 2193 1453 2207 1467
rect 2273 1453 2287 1467
rect 2213 1434 2227 1448
rect 2133 1333 2147 1347
rect 2113 1293 2127 1307
rect 2113 1253 2127 1267
rect 2053 1233 2067 1247
rect 2093 1233 2107 1247
rect 2013 1073 2027 1087
rect 1933 973 1947 987
rect 2073 1073 2087 1087
rect 2073 1033 2087 1047
rect 2033 953 2047 967
rect 1973 914 1987 928
rect 2013 914 2027 928
rect 1853 853 1867 867
rect 1833 793 1847 807
rect 1933 872 1947 886
rect 1993 872 2007 886
rect 2133 1214 2147 1228
rect 2233 1333 2247 1347
rect 2233 1312 2247 1326
rect 2193 1253 2207 1267
rect 2193 1214 2207 1228
rect 2413 1912 2427 1926
rect 2433 1853 2447 1867
rect 2373 1753 2387 1767
rect 2353 1733 2367 1747
rect 2393 1734 2407 1748
rect 2573 1912 2587 1926
rect 2573 1873 2587 1887
rect 2613 1873 2627 1887
rect 2533 1833 2547 1847
rect 2473 1813 2487 1827
rect 2513 1813 2527 1827
rect 2453 1733 2467 1747
rect 2513 1734 2527 1748
rect 2613 1773 2627 1787
rect 2553 1733 2567 1747
rect 2733 2133 2747 2147
rect 2693 2033 2707 2047
rect 2813 2173 2827 2187
rect 2773 2093 2787 2107
rect 2773 2013 2787 2027
rect 2733 1993 2747 2007
rect 2773 1954 2787 1968
rect 2693 1933 2707 1947
rect 2753 1912 2767 1926
rect 2793 1853 2807 1867
rect 2673 1753 2687 1767
rect 2653 1734 2667 1748
rect 2693 1733 2707 1747
rect 2753 1734 2767 1748
rect 2813 1793 2827 1807
rect 2413 1692 2427 1706
rect 2373 1673 2387 1687
rect 2353 1633 2367 1647
rect 2353 1593 2367 1607
rect 2333 1453 2347 1467
rect 2293 1433 2307 1447
rect 2413 1513 2427 1527
rect 2393 1473 2407 1487
rect 2333 1392 2347 1406
rect 2553 1553 2567 1567
rect 2433 1433 2447 1447
rect 2493 1453 2507 1467
rect 2513 1434 2527 1448
rect 2553 1434 2567 1448
rect 2593 1692 2607 1706
rect 2653 1673 2667 1687
rect 2633 1653 2647 1667
rect 2693 1653 2707 1667
rect 2733 1653 2747 1667
rect 2753 1633 2767 1647
rect 2693 1593 2707 1607
rect 2673 1493 2687 1507
rect 2633 1453 2647 1467
rect 2433 1393 2447 1407
rect 2413 1313 2427 1327
rect 2353 1293 2367 1307
rect 2393 1293 2407 1307
rect 2233 1213 2247 1227
rect 2133 1113 2147 1127
rect 2112 1013 2126 1027
rect 2133 1013 2147 1027
rect 2093 953 2107 967
rect 2213 1172 2227 1186
rect 2173 1132 2187 1146
rect 2213 1133 2227 1147
rect 2193 1113 2207 1127
rect 2233 1113 2247 1127
rect 2173 993 2187 1007
rect 2153 933 2167 947
rect 2133 914 2147 928
rect 1873 773 1887 787
rect 1873 752 1887 766
rect 2033 793 2047 807
rect 1953 773 1967 787
rect 1933 733 1947 747
rect 1913 694 1927 708
rect 1973 753 1987 767
rect 1953 693 1967 707
rect 1853 653 1867 667
rect 1813 593 1827 607
rect 1793 573 1807 587
rect 1813 453 1827 467
rect 1813 394 1827 408
rect 1933 652 1947 666
rect 2053 713 2067 727
rect 2113 853 2127 867
rect 2093 693 2107 707
rect 1893 613 1907 627
rect 1873 593 1887 607
rect 1853 573 1867 587
rect 1873 553 1887 567
rect 1973 652 1987 666
rect 2033 652 2047 666
rect 1953 513 1967 527
rect 1893 493 1907 507
rect 1853 433 1867 447
rect 1613 313 1627 327
rect 1653 313 1667 327
rect 1693 313 1707 327
rect 1533 253 1547 267
rect 1633 233 1647 247
rect 1533 213 1547 227
rect 1473 193 1487 207
rect 1613 193 1627 207
rect 873 132 887 146
rect 913 113 927 127
rect 1053 132 1067 146
rect 1093 132 1107 146
rect 1153 132 1167 146
rect 1193 133 1207 147
rect 1253 132 1267 146
rect 1293 132 1307 146
rect 1333 133 1347 147
rect 1393 132 1407 146
rect 1013 113 1027 127
rect 1433 113 1447 127
rect 573 93 587 107
rect 813 93 827 107
rect 1613 132 1627 146
rect 1653 174 1667 188
rect 1693 174 1707 188
rect 1793 352 1807 366
rect 2133 793 2147 807
rect 2173 873 2187 887
rect 2153 753 2167 767
rect 2233 1033 2247 1047
rect 2293 1253 2307 1267
rect 2333 1253 2347 1267
rect 2273 1214 2287 1228
rect 2413 1273 2427 1287
rect 2353 1233 2367 1247
rect 2333 1214 2347 1228
rect 2313 1172 2327 1186
rect 2493 1392 2507 1406
rect 2533 1393 2547 1407
rect 2473 1353 2487 1367
rect 2453 1273 2467 1287
rect 2593 1434 2607 1448
rect 2673 1433 2687 1447
rect 2553 1353 2567 1367
rect 2533 1333 2547 1347
rect 2513 1313 2527 1327
rect 2493 1293 2507 1307
rect 2473 1253 2487 1267
rect 2353 1133 2367 1147
rect 2353 1112 2367 1126
rect 2313 1093 2327 1107
rect 2253 933 2267 947
rect 2233 914 2247 928
rect 2333 1073 2347 1087
rect 2313 1053 2327 1067
rect 2193 813 2207 827
rect 2213 793 2227 807
rect 2173 713 2187 727
rect 2253 833 2267 847
rect 2233 713 2247 727
rect 2253 693 2267 707
rect 2153 633 2167 647
rect 2233 652 2247 666
rect 2293 813 2307 827
rect 2473 1053 2487 1067
rect 2513 1273 2527 1287
rect 2653 1392 2667 1406
rect 2713 1573 2727 1587
rect 2713 1513 2727 1527
rect 2813 1693 2827 1707
rect 2813 1613 2827 1627
rect 2813 1553 2827 1567
rect 2793 1493 2807 1507
rect 2773 1453 2787 1467
rect 2793 1433 2807 1447
rect 2613 1333 2627 1347
rect 2613 1253 2627 1267
rect 2513 1053 2527 1067
rect 2353 1033 2367 1047
rect 2332 1013 2346 1027
rect 2353 1012 2367 1026
rect 2333 992 2347 1006
rect 2333 913 2347 927
rect 2413 973 2427 987
rect 2393 953 2407 967
rect 2393 914 2407 928
rect 2493 1033 2507 1047
rect 2452 1013 2466 1027
rect 2473 1013 2487 1027
rect 2453 973 2467 987
rect 2493 953 2507 967
rect 2513 953 2527 967
rect 2473 914 2487 928
rect 2593 1113 2607 1127
rect 2573 933 2587 947
rect 2553 913 2567 927
rect 2433 893 2447 907
rect 2333 873 2347 887
rect 2753 1353 2767 1367
rect 2753 1332 2767 1346
rect 2793 1333 2807 1347
rect 2672 1273 2686 1287
rect 2693 1273 2707 1287
rect 2693 1233 2707 1247
rect 2633 1153 2647 1167
rect 2613 933 2627 947
rect 2693 1153 2707 1167
rect 2693 1013 2707 1027
rect 2733 1053 2747 1067
rect 2733 1013 2747 1027
rect 2713 973 2727 987
rect 2373 872 2387 886
rect 2353 853 2367 867
rect 2333 833 2347 847
rect 2313 693 2327 707
rect 2433 853 2447 867
rect 2533 872 2547 886
rect 2573 872 2587 886
rect 2713 933 2727 947
rect 2693 913 2707 927
rect 2793 1293 2807 1307
rect 2953 2413 2967 2427
rect 3133 2413 3147 2427
rect 2993 2333 3007 2347
rect 3133 2333 3147 2347
rect 2893 2273 2907 2287
rect 2933 2254 2947 2268
rect 3653 3413 3667 3427
rect 3593 3353 3607 3367
rect 3573 3333 3587 3347
rect 3553 3173 3567 3187
rect 3473 3113 3487 3127
rect 3473 3073 3487 3087
rect 3473 2994 3487 3008
rect 3493 2933 3507 2947
rect 3673 3313 3687 3327
rect 3633 3294 3647 3308
rect 3593 3193 3607 3207
rect 3593 3153 3607 3167
rect 3573 2933 3587 2947
rect 3453 2853 3467 2867
rect 3533 2853 3547 2867
rect 3453 2732 3467 2746
rect 3493 2732 3507 2746
rect 3553 2732 3567 2746
rect 3613 3033 3627 3047
rect 3293 2693 3307 2707
rect 3433 2693 3447 2707
rect 3473 2693 3487 2707
rect 3553 2693 3567 2707
rect 3533 2653 3547 2667
rect 3473 2593 3487 2607
rect 3313 2513 3327 2527
rect 3513 2513 3527 2527
rect 3353 2493 3367 2507
rect 3473 2493 3487 2507
rect 3393 2474 3407 2488
rect 3433 2474 3447 2488
rect 3233 2433 3247 2447
rect 3273 2433 3287 2447
rect 3213 2333 3227 2347
rect 3153 2293 3167 2307
rect 3013 2253 3027 2267
rect 3133 2253 3147 2267
rect 3173 2254 3187 2268
rect 2913 2213 2927 2227
rect 2993 2213 3007 2227
rect 2893 2153 2907 2167
rect 3133 2213 3147 2227
rect 3113 2193 3127 2207
rect 3012 2153 3026 2167
rect 3033 2153 3047 2167
rect 3113 2093 3127 2107
rect 3513 2473 3527 2487
rect 3333 2413 3347 2427
rect 3393 2413 3407 2427
rect 3493 2432 3507 2446
rect 3373 2393 3387 2407
rect 3453 2393 3467 2407
rect 3253 2333 3267 2347
rect 3233 2193 3247 2207
rect 3153 2093 3167 2107
rect 2913 2073 2927 2087
rect 3133 2073 3147 2087
rect 2893 2033 2907 2047
rect 3053 2053 3067 2067
rect 2933 1933 2947 1947
rect 2873 1912 2887 1926
rect 2853 1833 2867 1847
rect 2913 1813 2927 1827
rect 2973 2013 2987 2027
rect 2973 1973 2987 1987
rect 3032 1954 3046 1968
rect 3152 2033 3166 2047
rect 3173 2033 3187 2047
rect 3413 2373 3427 2387
rect 3393 2293 3407 2307
rect 3373 2253 3387 2267
rect 3272 2213 3286 2227
rect 3293 2212 3307 2226
rect 3453 2254 3467 2268
rect 3513 2393 3527 2407
rect 3513 2313 3527 2327
rect 3673 3252 3687 3266
rect 3733 3472 3747 3486
rect 3713 3413 3727 3427
rect 3713 3333 3727 3347
rect 3753 3393 3767 3407
rect 3733 3293 3747 3307
rect 3833 3533 3847 3547
rect 3853 3472 3867 3486
rect 3853 3433 3867 3447
rect 3813 3393 3827 3407
rect 3773 3353 3787 3367
rect 3973 3772 3987 3786
rect 4013 3653 4027 3667
rect 3933 3633 3947 3647
rect 4053 3633 4067 3647
rect 4013 3613 4027 3627
rect 4033 3593 4047 3607
rect 3953 3533 3967 3547
rect 3993 3514 4007 3528
rect 4013 3473 4027 3487
rect 3933 3433 3947 3447
rect 3893 3393 3907 3407
rect 4253 3992 4267 4006
rect 4293 3992 4307 4006
rect 4253 3933 4267 3947
rect 4233 3913 4247 3927
rect 4093 3833 4107 3847
rect 4133 3833 4147 3847
rect 4193 3833 4207 3847
rect 4093 3772 4107 3786
rect 4133 3772 4147 3786
rect 4193 3772 4207 3786
rect 4113 3733 4127 3747
rect 4093 3713 4107 3727
rect 4073 3553 4087 3567
rect 4053 3513 4067 3527
rect 4213 3733 4227 3747
rect 4233 3713 4247 3727
rect 4192 3673 4206 3687
rect 4213 3673 4227 3687
rect 4113 3653 4127 3667
rect 4173 3633 4187 3647
rect 4153 3593 4167 3607
rect 4133 3514 4147 3528
rect 4493 4113 4507 4127
rect 4473 4093 4487 4107
rect 4353 4073 4367 4087
rect 4433 4053 4447 4067
rect 4393 4034 4407 4048
rect 4973 5032 4987 5046
rect 5013 5032 5027 5046
rect 5093 5032 5107 5046
rect 5152 5032 5166 5046
rect 5173 5033 5187 5047
rect 5053 4953 5067 4967
rect 4993 4913 5007 4927
rect 4933 4893 4947 4907
rect 4933 4853 4947 4867
rect 5053 4893 5067 4907
rect 5133 4893 5147 4907
rect 4933 4793 4947 4807
rect 5093 4854 5107 4868
rect 5233 5032 5247 5046
rect 5273 5032 5287 5046
rect 5233 4973 5247 4987
rect 5273 4973 5287 4987
rect 5113 4812 5127 4826
rect 5173 4813 5187 4827
rect 5013 4773 5027 4787
rect 5053 4773 5067 4787
rect 5213 4773 5227 4787
rect 4873 4693 4887 4707
rect 4913 4693 4927 4707
rect 4853 4633 4867 4647
rect 4693 4554 4707 4568
rect 4753 4553 4767 4567
rect 4813 4554 4827 4568
rect 4853 4553 4867 4567
rect 4713 4512 4727 4526
rect 4753 4512 4767 4526
rect 4673 4493 4687 4507
rect 4673 4413 4687 4427
rect 4673 4373 4687 4387
rect 4893 4593 4907 4607
rect 4933 4593 4947 4607
rect 4973 4554 4987 4568
rect 4993 4513 5007 4527
rect 4953 4493 4967 4507
rect 4873 4453 4887 4467
rect 4833 4413 4847 4427
rect 4833 4373 4847 4387
rect 4973 4453 4987 4467
rect 4953 4353 4967 4367
rect 4793 4334 4807 4348
rect 4833 4333 4847 4347
rect 4873 4334 4887 4348
rect 4613 4292 4627 4306
rect 4773 4292 4787 4306
rect 4693 4273 4707 4287
rect 4593 4173 4607 4187
rect 4633 4153 4647 4167
rect 4573 4093 4587 4107
rect 4513 4073 4527 4087
rect 4493 4053 4507 4067
rect 4513 4034 4527 4048
rect 4553 4034 4567 4048
rect 4593 4034 4607 4048
rect 4773 4153 4787 4167
rect 4693 4133 4707 4147
rect 4893 4292 4907 4306
rect 4793 4093 4807 4107
rect 4753 4034 4767 4048
rect 4373 3992 4387 4006
rect 4433 3993 4447 4007
rect 4613 3992 4627 4006
rect 4593 3973 4607 3987
rect 4653 3973 4667 3987
rect 4493 3953 4507 3967
rect 4553 3953 4567 3967
rect 4273 3833 4287 3847
rect 4313 3833 4327 3847
rect 4333 3813 4347 3827
rect 4273 3773 4287 3787
rect 4293 3753 4307 3767
rect 4253 3693 4267 3707
rect 4193 3593 4207 3607
rect 4233 3593 4247 3607
rect 4173 3573 4187 3587
rect 4233 3533 4247 3547
rect 4273 3533 4287 3547
rect 4113 3472 4127 3486
rect 4273 3473 4287 3487
rect 4093 3453 4107 3467
rect 4073 3413 4087 3427
rect 4333 3753 4347 3767
rect 4313 3673 4327 3687
rect 4393 3514 4407 3528
rect 4353 3472 4367 3486
rect 4393 3473 4407 3487
rect 4293 3433 4307 3447
rect 4293 3393 4307 3407
rect 4193 3333 4207 3347
rect 4433 3772 4447 3786
rect 4493 3773 4507 3787
rect 4493 3713 4507 3727
rect 4573 3733 4587 3747
rect 4513 3633 4527 3647
rect 4813 3992 4827 4006
rect 4873 3992 4887 4006
rect 4793 3953 4807 3967
rect 4953 4293 4967 4307
rect 5153 4733 5167 4747
rect 5133 4673 5147 4687
rect 5033 4593 5047 4607
rect 5093 4554 5107 4568
rect 5133 4553 5147 4567
rect 5213 4554 5227 4568
rect 5253 4554 5267 4568
rect 5033 4512 5047 4526
rect 5113 4512 5127 4526
rect 5033 4413 5047 4427
rect 5013 4292 5027 4306
rect 4973 4213 4987 4227
rect 4993 4073 5007 4087
rect 5213 4473 5227 4487
rect 5193 4433 5207 4447
rect 5093 4413 5107 4427
rect 5173 4353 5187 4367
rect 5133 4334 5147 4348
rect 5153 4292 5167 4306
rect 5353 4973 5367 4987
rect 5713 5113 5727 5127
rect 5753 5113 5767 5127
rect 5653 5073 5667 5087
rect 5493 5013 5507 5027
rect 5433 4993 5447 5007
rect 5473 4993 5487 5007
rect 5393 4953 5407 4967
rect 5473 4953 5487 4967
rect 5313 4913 5327 4927
rect 5333 4812 5347 4826
rect 5373 4812 5387 4826
rect 5373 4733 5387 4747
rect 5393 4713 5407 4727
rect 5453 4713 5467 4727
rect 5373 4533 5387 4547
rect 5273 4512 5287 4526
rect 5333 4512 5347 4526
rect 5253 4433 5267 4447
rect 5373 4413 5387 4427
rect 5213 4333 5227 4347
rect 5253 4334 5267 4348
rect 5313 4333 5327 4347
rect 5353 4334 5367 4348
rect 5553 4893 5567 4907
rect 5653 4993 5667 5007
rect 5713 4913 5727 4927
rect 5693 4893 5707 4907
rect 5833 4913 5847 4927
rect 5713 4872 5727 4886
rect 5673 4854 5687 4868
rect 5493 4813 5507 4827
rect 5613 4813 5627 4827
rect 5473 4693 5487 4707
rect 5513 4693 5527 4707
rect 5453 4554 5467 4568
rect 5433 4512 5447 4526
rect 5433 4473 5447 4487
rect 5473 4453 5487 4467
rect 5573 4593 5587 4607
rect 5613 4593 5627 4607
rect 5553 4473 5567 4487
rect 5573 4453 5587 4467
rect 5513 4433 5527 4447
rect 5553 4433 5567 4447
rect 5433 4413 5447 4427
rect 5433 4373 5447 4387
rect 5553 4333 5567 4347
rect 5113 4173 5127 4187
rect 5033 4034 5047 4048
rect 5073 4032 5087 4046
rect 5173 4173 5187 4187
rect 5253 4113 5267 4127
rect 5173 4053 5187 4067
rect 4933 3992 4947 4006
rect 4973 3992 4987 4006
rect 5013 3953 5027 3967
rect 4853 3913 4867 3927
rect 4913 3913 4927 3927
rect 4653 3833 4667 3847
rect 4613 3813 4627 3827
rect 4693 3814 4707 3828
rect 4753 3813 4767 3827
rect 4813 3814 4827 3828
rect 5133 3992 5147 4006
rect 5113 3973 5127 3987
rect 4993 3893 5007 3907
rect 5073 3893 5087 3907
rect 4853 3813 4867 3827
rect 4973 3814 4987 3828
rect 4613 3772 4627 3786
rect 4673 3772 4687 3786
rect 4713 3772 4727 3786
rect 4753 3772 4767 3786
rect 4673 3753 4687 3767
rect 4793 3753 4807 3767
rect 4853 3773 4867 3787
rect 4833 3753 4847 3767
rect 4633 3693 4647 3707
rect 4873 3713 4887 3727
rect 4973 3753 4987 3767
rect 4953 3693 4967 3707
rect 5053 3814 5067 3828
rect 5093 3772 5107 3786
rect 5073 3753 5087 3767
rect 5073 3693 5087 3707
rect 4853 3653 4867 3667
rect 4993 3653 5007 3667
rect 4673 3633 4687 3647
rect 4613 3593 4627 3607
rect 4493 3553 4507 3567
rect 4593 3553 4607 3567
rect 4453 3514 4467 3528
rect 4573 3514 4587 3528
rect 4593 3472 4607 3486
rect 4733 3593 4747 3607
rect 4753 3573 4767 3587
rect 4733 3553 4747 3567
rect 4473 3433 4487 3447
rect 4713 3413 4727 3427
rect 4613 3393 4627 3407
rect 4413 3333 4427 3347
rect 4013 3293 4027 3307
rect 3713 3252 3727 3266
rect 3853 3252 3867 3266
rect 3893 3252 3907 3266
rect 3953 3252 3967 3266
rect 3873 3213 3887 3227
rect 3693 3113 3707 3127
rect 3773 3033 3787 3047
rect 3633 2994 3647 3008
rect 3813 2994 3827 3008
rect 4673 3333 4687 3347
rect 4333 3294 4347 3308
rect 4373 3294 4387 3308
rect 4433 3294 4447 3308
rect 4473 3294 4487 3308
rect 4193 3252 4207 3266
rect 4213 3153 4227 3167
rect 4113 3113 4127 3127
rect 4173 3113 4187 3127
rect 3933 3073 3947 3087
rect 4033 3073 4047 3087
rect 4013 3033 4027 3047
rect 3973 2994 3987 3008
rect 4013 2994 4027 3008
rect 4073 2994 4087 3008
rect 3673 2813 3687 2827
rect 3693 2813 3707 2827
rect 3733 2774 3747 2788
rect 3613 2693 3627 2707
rect 3673 2693 3687 2707
rect 3593 2533 3607 2547
rect 3653 2533 3667 2547
rect 3633 2474 3647 2488
rect 3833 2952 3847 2966
rect 3873 2953 3887 2967
rect 3913 2913 3927 2927
rect 4173 2994 4187 3008
rect 4333 3033 4347 3047
rect 4253 2994 4267 3008
rect 4293 2994 4307 3008
rect 4113 2953 4127 2967
rect 4153 2952 4167 2966
rect 3973 2913 3987 2927
rect 4013 2913 4027 2927
rect 4053 2913 4067 2927
rect 3953 2873 3967 2887
rect 3813 2813 3827 2827
rect 3953 2774 3967 2788
rect 3813 2733 3827 2747
rect 3853 2732 3867 2746
rect 3913 2732 3927 2746
rect 3793 2653 3807 2667
rect 3893 2613 3907 2627
rect 3753 2593 3767 2607
rect 3793 2593 3807 2607
rect 3713 2553 3727 2567
rect 3673 2513 3687 2527
rect 3773 2573 3787 2587
rect 3753 2493 3767 2507
rect 3573 2413 3587 2427
rect 3553 2373 3567 2387
rect 3553 2273 3567 2287
rect 3533 2253 3547 2267
rect 3413 2193 3427 2207
rect 3353 2173 3367 2187
rect 3093 2013 3107 2027
rect 3073 1993 3087 2007
rect 3053 1953 3067 1967
rect 2973 1913 2987 1927
rect 3133 1954 3147 1968
rect 3253 2033 3267 2047
rect 3272 1954 3286 1968
rect 3333 2113 3347 2127
rect 3413 2113 3427 2127
rect 3313 2093 3327 2107
rect 3293 1953 3307 1967
rect 2953 1833 2967 1847
rect 2953 1793 2967 1807
rect 2933 1753 2947 1767
rect 2853 1732 2867 1746
rect 2913 1734 2927 1748
rect 2853 1673 2867 1687
rect 2893 1673 2907 1687
rect 2873 1633 2887 1647
rect 2853 1513 2867 1527
rect 2873 1493 2887 1507
rect 2873 1453 2887 1467
rect 2933 1653 2947 1667
rect 2933 1632 2947 1646
rect 2933 1573 2947 1587
rect 3073 1912 3087 1926
rect 3113 1912 3127 1926
rect 3193 1913 3207 1927
rect 3293 1913 3307 1927
rect 3153 1893 3167 1907
rect 3153 1872 3167 1886
rect 3053 1853 3067 1867
rect 3053 1813 3067 1827
rect 3033 1734 3047 1748
rect 3073 1734 3087 1748
rect 3113 1734 3127 1748
rect 3273 1873 3287 1887
rect 3213 1833 3227 1847
rect 3193 1813 3207 1827
rect 3193 1734 3207 1748
rect 2993 1673 3007 1687
rect 2973 1593 2987 1607
rect 2953 1553 2967 1567
rect 2993 1493 3007 1507
rect 2933 1473 2947 1487
rect 2893 1434 2907 1448
rect 2833 1393 2847 1407
rect 2813 1253 2827 1267
rect 2873 1392 2887 1406
rect 2833 1233 2847 1247
rect 2753 933 2767 947
rect 2853 1214 2867 1228
rect 3053 1553 3067 1567
rect 3033 1533 3047 1547
rect 3053 1513 3067 1527
rect 3012 1473 3026 1487
rect 3033 1473 3047 1487
rect 2973 1434 2987 1448
rect 3033 1392 3047 1406
rect 3013 1333 3027 1347
rect 2993 1293 3007 1307
rect 2973 1273 2987 1287
rect 2933 1214 2947 1228
rect 2973 1213 2987 1227
rect 2873 1193 2887 1207
rect 2833 1073 2847 1087
rect 2893 1113 2907 1127
rect 2873 1073 2887 1087
rect 2853 1053 2867 1067
rect 2833 993 2847 1007
rect 2813 973 2827 987
rect 2493 853 2507 867
rect 2593 853 2607 867
rect 2673 873 2687 887
rect 2653 833 2667 847
rect 2513 793 2527 807
rect 2373 753 2387 767
rect 2413 753 2427 767
rect 2493 753 2507 767
rect 2173 613 2187 627
rect 2213 613 2227 627
rect 2273 612 2287 626
rect 2133 553 2147 567
rect 2153 493 2167 507
rect 2113 473 2127 487
rect 2013 453 2027 467
rect 1933 394 1947 408
rect 1853 352 1867 366
rect 1913 352 1927 366
rect 1793 293 1807 307
rect 1833 293 1847 307
rect 1973 333 1987 347
rect 1953 253 1967 267
rect 1853 193 1867 207
rect 2073 394 2087 408
rect 2193 473 2207 487
rect 2233 453 2247 467
rect 2193 394 2207 408
rect 2293 533 2307 547
rect 2313 473 2327 487
rect 2272 393 2286 407
rect 2293 394 2307 408
rect 2453 694 2467 708
rect 2373 613 2387 627
rect 2413 613 2427 627
rect 2373 592 2387 606
rect 2493 653 2507 667
rect 2453 613 2467 627
rect 2433 593 2447 607
rect 2393 573 2407 587
rect 2453 573 2467 587
rect 2373 553 2387 567
rect 2353 493 2367 507
rect 2433 553 2447 567
rect 2413 533 2427 547
rect 2393 513 2407 527
rect 2333 453 2347 467
rect 2373 473 2387 487
rect 2353 413 2367 427
rect 2093 352 2107 366
rect 2152 352 2166 366
rect 2173 353 2187 367
rect 2053 333 2067 347
rect 2013 293 2027 307
rect 2133 293 2147 307
rect 2053 233 2067 247
rect 2013 213 2027 227
rect 1913 173 1927 187
rect 1973 174 1987 188
rect 1793 153 1807 167
rect 2093 174 2107 188
rect 2213 333 2227 347
rect 2193 213 2207 227
rect 2333 394 2347 408
rect 2393 433 2407 447
rect 2413 393 2427 407
rect 2293 313 2307 327
rect 2353 352 2367 366
rect 2413 353 2427 367
rect 2573 753 2587 767
rect 2573 694 2587 708
rect 2773 873 2787 887
rect 2753 853 2767 867
rect 2693 753 2707 767
rect 2513 593 2527 607
rect 2493 533 2507 547
rect 2453 493 2467 507
rect 2593 652 2607 666
rect 2553 593 2567 607
rect 2553 533 2567 547
rect 2493 473 2507 487
rect 2533 473 2547 487
rect 2453 433 2467 447
rect 2533 433 2547 447
rect 2573 433 2587 447
rect 2633 433 2647 447
rect 2553 393 2567 407
rect 2393 313 2407 327
rect 2313 293 2327 307
rect 2473 333 2487 347
rect 2433 313 2447 327
rect 2473 293 2487 307
rect 2673 693 2687 707
rect 2733 753 2747 767
rect 2713 713 2727 727
rect 2793 833 2807 847
rect 2953 1172 2967 1186
rect 2993 1172 3007 1186
rect 3093 1693 3107 1707
rect 3133 1692 3147 1706
rect 3193 1692 3207 1706
rect 3193 1653 3207 1667
rect 3113 1633 3127 1647
rect 3093 1593 3107 1607
rect 3113 1573 3127 1587
rect 3113 1513 3127 1527
rect 3113 1473 3127 1487
rect 3153 1473 3167 1487
rect 3092 1433 3106 1447
rect 3113 1434 3127 1448
rect 3093 1393 3107 1407
rect 3073 1333 3087 1347
rect 3073 1293 3087 1307
rect 3033 1253 3047 1267
rect 3133 1353 3147 1367
rect 3093 1273 3107 1287
rect 3113 1253 3127 1267
rect 2953 1113 2967 1127
rect 2913 1093 2927 1107
rect 2933 1073 2947 1087
rect 2913 953 2927 967
rect 2913 914 2927 928
rect 2853 853 2867 867
rect 2812 813 2826 827
rect 2833 813 2847 827
rect 2793 753 2807 767
rect 3052 1153 3066 1167
rect 3073 1153 3087 1167
rect 3013 1093 3027 1107
rect 3053 1073 3067 1087
rect 3033 1053 3047 1067
rect 3033 1032 3047 1046
rect 2953 1013 2967 1027
rect 3013 1013 3027 1027
rect 2993 993 3007 1007
rect 2993 933 3007 947
rect 2973 914 2987 928
rect 3033 993 3047 1007
rect 3053 973 3067 987
rect 3033 872 3047 886
rect 2993 813 3007 827
rect 2933 793 2947 807
rect 2913 753 2927 767
rect 2993 753 3007 767
rect 2833 733 2847 747
rect 2973 733 2987 747
rect 3013 733 3027 747
rect 2813 693 2827 707
rect 2853 694 2867 708
rect 2933 694 2947 708
rect 2993 694 3007 708
rect 3033 694 3047 708
rect 2793 673 2807 687
rect 2673 653 2687 667
rect 2693 633 2707 647
rect 2673 433 2687 447
rect 2673 394 2687 408
rect 2773 653 2787 667
rect 2753 613 2767 627
rect 2713 493 2727 507
rect 2833 652 2847 666
rect 2873 652 2887 666
rect 2913 652 2927 666
rect 2953 633 2967 647
rect 2933 613 2947 627
rect 2913 513 2927 527
rect 3013 652 3027 666
rect 3053 633 3067 647
rect 2973 613 2987 627
rect 3013 593 3027 607
rect 3013 572 3027 586
rect 3033 553 3047 567
rect 2953 493 2967 507
rect 3013 493 3027 507
rect 2713 472 2727 486
rect 2773 473 2787 487
rect 2813 473 2827 487
rect 2993 473 3007 487
rect 2593 353 2607 367
rect 2533 293 2547 307
rect 2573 293 2587 307
rect 2293 273 2307 287
rect 2333 273 2347 287
rect 2413 273 2427 287
rect 2513 273 2527 287
rect 2173 173 2187 187
rect 2213 193 2227 207
rect 2252 193 2266 207
rect 2273 193 2287 207
rect 2293 174 2307 188
rect 1713 132 1727 146
rect 1753 132 1767 146
rect 1653 113 1667 127
rect 1633 73 1647 87
rect 1873 132 1887 146
rect 1913 132 1927 146
rect 1953 132 1967 146
rect 1833 93 1847 107
rect 1953 93 1967 107
rect 1653 53 1667 67
rect 2053 132 2067 146
rect 2153 132 2167 146
rect 2193 132 2207 146
rect 2133 93 2147 107
rect 2273 132 2287 146
rect 2233 93 2247 107
rect 2133 53 2147 67
rect 2193 53 2207 67
rect 533 33 547 47
rect 1433 33 1447 47
rect 1473 33 1487 47
rect 1993 33 2007 47
rect 2493 253 2507 267
rect 2373 233 2387 247
rect 2473 233 2487 247
rect 2553 233 2567 247
rect 2373 174 2387 188
rect 2413 174 2427 188
rect 2373 113 2387 127
rect 2433 132 2447 146
rect 2513 213 2527 227
rect 2553 174 2567 188
rect 2613 333 2627 347
rect 2613 273 2627 287
rect 2593 173 2607 187
rect 2533 132 2547 146
rect 2573 132 2587 146
rect 2473 113 2487 127
rect 2513 113 2527 127
rect 2673 333 2687 347
rect 2633 253 2647 267
rect 2673 273 2687 287
rect 2653 193 2667 207
rect 2973 453 2987 467
rect 2793 433 2807 447
rect 2773 413 2787 427
rect 2953 413 2967 427
rect 2813 394 2827 408
rect 2853 394 2867 408
rect 2913 394 2927 408
rect 2953 394 2967 408
rect 2733 353 2747 367
rect 2713 333 2727 347
rect 2733 293 2747 307
rect 2793 313 2807 327
rect 2753 233 2767 247
rect 2813 193 2827 207
rect 2753 173 2767 187
rect 2813 174 2827 188
rect 2853 313 2867 327
rect 2933 293 2947 307
rect 2933 233 2947 247
rect 2893 213 2907 227
rect 2653 132 2667 146
rect 2733 133 2747 147
rect 2693 113 2707 127
rect 2393 93 2407 107
rect 2573 93 2587 107
rect 2633 93 2647 107
rect 2373 33 2387 47
rect 2533 33 2547 47
rect 2333 13 2347 27
rect 2453 13 2467 27
rect 2673 93 2687 107
rect 2673 33 2687 47
rect 2793 113 2807 127
rect 2753 93 2767 107
rect 2573 13 2587 27
rect 2653 13 2667 27
rect 2693 13 2707 27
rect 2732 33 2746 47
rect 2753 33 2767 47
rect 2873 173 2887 187
rect 2973 213 2987 227
rect 2913 132 2927 146
rect 2953 132 2967 146
rect 3053 433 3067 447
rect 3033 413 3047 427
rect 3113 1173 3127 1187
rect 3233 1813 3247 1827
rect 3293 1773 3307 1787
rect 3393 1873 3407 1887
rect 3513 2212 3527 2226
rect 3513 2173 3527 2187
rect 3713 2474 3727 2488
rect 3773 2473 3787 2487
rect 3733 2432 3747 2446
rect 3753 2333 3767 2347
rect 3613 2293 3627 2307
rect 3673 2293 3687 2307
rect 3593 2273 3607 2287
rect 3933 2713 3947 2727
rect 3913 2533 3927 2547
rect 3893 2493 3907 2507
rect 3813 2474 3827 2488
rect 3853 2474 3867 2488
rect 4513 3293 4527 3307
rect 4573 3294 4587 3308
rect 4613 3294 4627 3308
rect 4673 3294 4687 3308
rect 4453 3252 4467 3266
rect 4433 3233 4447 3247
rect 4413 3153 4427 3167
rect 4553 3252 4567 3266
rect 4513 3193 4527 3207
rect 4913 3553 4927 3567
rect 4773 3514 4787 3528
rect 4833 3514 4847 3528
rect 4873 3514 4887 3528
rect 4953 3514 4967 3528
rect 4993 3513 5007 3527
rect 4773 3433 4787 3447
rect 4853 3472 4867 3486
rect 4913 3473 4927 3487
rect 4993 3473 5007 3487
rect 4853 3433 4867 3447
rect 4973 3433 4987 3447
rect 4813 3413 4827 3427
rect 4753 3373 4767 3387
rect 4813 3373 4827 3387
rect 4653 3233 4667 3247
rect 4713 3253 4727 3267
rect 4693 3233 4707 3247
rect 4793 3252 4807 3266
rect 4833 3252 4847 3266
rect 4893 3393 4907 3407
rect 4873 3313 4887 3327
rect 5073 3633 5087 3647
rect 5073 3553 5087 3567
rect 5353 4273 5367 4287
rect 5313 4253 5327 4267
rect 5353 4213 5367 4227
rect 5273 4093 5287 4107
rect 5313 4034 5327 4048
rect 5293 3992 5307 4006
rect 5453 4293 5467 4307
rect 5413 4273 5427 4287
rect 5393 4253 5407 4267
rect 5433 4253 5447 4267
rect 5393 4034 5407 4048
rect 5533 4273 5547 4287
rect 5473 4133 5487 4147
rect 5453 4033 5467 4047
rect 5533 4053 5547 4067
rect 5573 4273 5587 4287
rect 5553 4033 5567 4047
rect 5333 3973 5347 3987
rect 5373 3973 5387 3987
rect 5233 3913 5247 3927
rect 5353 3913 5367 3927
rect 5253 3873 5267 3887
rect 5173 3853 5187 3867
rect 5233 3853 5247 3867
rect 5133 3814 5147 3828
rect 5193 3814 5207 3828
rect 5113 3733 5127 3747
rect 5113 3653 5127 3667
rect 5113 3593 5127 3607
rect 5153 3772 5167 3786
rect 5313 3814 5327 3828
rect 5373 3813 5387 3827
rect 5153 3733 5167 3747
rect 5093 3472 5107 3486
rect 5013 3453 5027 3467
rect 5053 3453 5067 3467
rect 4933 3313 4947 3327
rect 4993 3294 5007 3308
rect 4913 3252 4927 3266
rect 4953 3233 4967 3247
rect 4753 3213 4767 3227
rect 4853 3213 4867 3227
rect 4533 3073 4547 3087
rect 4613 3033 4627 3047
rect 4613 2973 4627 2987
rect 4313 2952 4327 2966
rect 4373 2953 4387 2967
rect 4413 2952 4427 2966
rect 4453 2952 4467 2966
rect 4553 2952 4567 2966
rect 4193 2873 4207 2887
rect 4253 2873 4267 2887
rect 4373 2833 4387 2847
rect 3993 2813 4007 2827
rect 4013 2793 4027 2807
rect 4233 2793 4247 2807
rect 4333 2793 4347 2807
rect 4373 2793 4387 2807
rect 4113 2773 4127 2787
rect 4173 2774 4187 2788
rect 4033 2732 4047 2746
rect 3973 2713 3987 2727
rect 3953 2653 3967 2667
rect 4153 2732 4167 2746
rect 4053 2713 4067 2727
rect 4093 2693 4107 2707
rect 4052 2653 4066 2667
rect 4073 2653 4087 2667
rect 4033 2613 4047 2627
rect 3953 2533 3967 2547
rect 3933 2473 3947 2487
rect 4013 2474 4027 2488
rect 4053 2473 4067 2487
rect 3812 2433 3826 2447
rect 3833 2433 3847 2447
rect 3933 2433 3947 2447
rect 3793 2253 3807 2267
rect 3553 2153 3567 2167
rect 3493 2093 3507 2107
rect 3453 2073 3467 2087
rect 3473 1973 3487 1987
rect 3453 1913 3467 1927
rect 3433 1833 3447 1847
rect 3333 1813 3347 1827
rect 3353 1793 3367 1807
rect 3253 1734 3267 1748
rect 3313 1692 3327 1706
rect 3373 1773 3387 1787
rect 3413 1773 3427 1787
rect 3353 1653 3367 1667
rect 3333 1633 3347 1647
rect 3273 1593 3287 1607
rect 3553 1954 3567 1968
rect 3593 2212 3607 2226
rect 3693 2212 3707 2226
rect 3733 2212 3747 2226
rect 3773 2212 3787 2226
rect 3753 2173 3767 2187
rect 3693 2133 3707 2147
rect 3593 2113 3607 2127
rect 3613 2053 3627 2067
rect 3593 2013 3607 2027
rect 3713 2053 3727 2067
rect 3733 2033 3747 2047
rect 3653 1973 3667 1987
rect 3593 1953 3607 1967
rect 3733 1954 3747 1968
rect 3533 1893 3547 1907
rect 3573 1893 3587 1907
rect 3633 1912 3647 1926
rect 3673 1912 3687 1926
rect 3573 1872 3587 1886
rect 3552 1793 3566 1807
rect 3573 1793 3587 1807
rect 3533 1753 3547 1767
rect 3633 1873 3647 1887
rect 3613 1853 3627 1867
rect 3393 1692 3407 1706
rect 3373 1493 3387 1507
rect 3293 1473 3307 1487
rect 3353 1473 3367 1487
rect 3232 1433 3246 1447
rect 3253 1434 3267 1448
rect 3253 1373 3267 1387
rect 3213 1353 3227 1367
rect 3173 1293 3187 1307
rect 3153 1213 3167 1227
rect 3193 1214 3207 1228
rect 3133 1153 3147 1167
rect 3113 1133 3127 1147
rect 3173 1073 3187 1087
rect 3113 1033 3127 1047
rect 3153 1013 3167 1027
rect 3093 973 3107 987
rect 3313 1393 3327 1407
rect 3473 1693 3487 1707
rect 3453 1633 3467 1647
rect 3433 1434 3447 1448
rect 3493 1673 3507 1687
rect 3573 1673 3587 1687
rect 3593 1573 3607 1587
rect 3553 1553 3567 1567
rect 3573 1533 3587 1547
rect 3553 1493 3567 1507
rect 3573 1453 3587 1467
rect 3513 1434 3527 1448
rect 3613 1533 3627 1547
rect 3273 1313 3287 1327
rect 3353 1392 3367 1406
rect 3413 1392 3427 1406
rect 3473 1392 3487 1406
rect 3533 1392 3547 1406
rect 3593 1392 3607 1406
rect 3413 1353 3427 1367
rect 3333 1333 3347 1347
rect 3313 1293 3327 1307
rect 3333 1253 3347 1267
rect 3373 1253 3387 1267
rect 3273 1213 3287 1227
rect 3333 1214 3347 1228
rect 3273 1172 3287 1186
rect 3313 1172 3327 1186
rect 3333 1153 3347 1167
rect 3273 1133 3287 1147
rect 3393 1173 3407 1187
rect 3332 1073 3346 1087
rect 3353 1073 3367 1087
rect 3232 1033 3246 1047
rect 3253 1033 3267 1047
rect 3213 973 3227 987
rect 3193 953 3207 967
rect 3213 933 3227 947
rect 3293 1013 3307 1027
rect 3253 993 3267 1007
rect 3353 1033 3367 1047
rect 3333 973 3347 987
rect 3172 872 3186 886
rect 3193 873 3207 887
rect 3093 833 3107 847
rect 3133 833 3147 847
rect 3173 833 3187 847
rect 3133 793 3147 807
rect 3113 753 3127 767
rect 3193 773 3207 787
rect 3173 694 3187 708
rect 3333 914 3347 928
rect 3233 873 3247 887
rect 3193 652 3207 666
rect 3153 593 3167 607
rect 3113 493 3127 507
rect 3273 793 3287 807
rect 3353 873 3367 887
rect 3273 753 3287 767
rect 3313 753 3327 767
rect 3273 732 3287 746
rect 3393 1053 3407 1067
rect 3393 953 3407 967
rect 3433 1313 3447 1327
rect 3453 1293 3467 1307
rect 3613 1353 3627 1367
rect 3513 1333 3527 1347
rect 3473 1234 3487 1248
rect 3713 1853 3727 1867
rect 3713 1813 3727 1827
rect 3653 1793 3667 1807
rect 3713 1792 3727 1806
rect 3673 1773 3687 1787
rect 3673 1733 3687 1747
rect 3773 2093 3787 2107
rect 3873 2413 3887 2427
rect 3833 2393 3847 2407
rect 3913 2293 3927 2307
rect 4053 2413 4067 2427
rect 4093 2633 4107 2647
rect 4293 2774 4307 2788
rect 4273 2713 4287 2727
rect 4253 2673 4267 2687
rect 4193 2593 4207 2607
rect 4173 2513 4187 2527
rect 4153 2373 4167 2387
rect 4433 2774 4447 2788
rect 4493 2774 4507 2788
rect 4333 2673 4347 2687
rect 4393 2673 4407 2687
rect 4353 2653 4367 2667
rect 4273 2573 4287 2587
rect 4333 2573 4347 2587
rect 4293 2513 4307 2527
rect 4253 2474 4267 2488
rect 4053 2293 4067 2307
rect 3933 2273 3947 2287
rect 4013 2254 4027 2268
rect 3953 2212 3967 2226
rect 3993 2212 4007 2226
rect 4033 2212 4047 2226
rect 3813 2173 3827 2187
rect 3873 2173 3887 2187
rect 3993 2173 4007 2187
rect 3813 2133 3827 2147
rect 3853 2093 3867 2107
rect 3813 2073 3827 2087
rect 3773 1954 3787 1968
rect 3833 1954 3847 1968
rect 3753 1873 3767 1887
rect 3793 1833 3807 1847
rect 3773 1793 3787 1807
rect 3733 1753 3747 1767
rect 3693 1692 3707 1706
rect 3733 1692 3747 1706
rect 3993 2053 4007 2067
rect 3953 1954 3967 1968
rect 3993 1953 4007 1967
rect 3873 1893 3887 1907
rect 3913 1893 3927 1907
rect 3873 1853 3887 1867
rect 3813 1773 3827 1787
rect 3853 1773 3867 1787
rect 3833 1734 3847 1748
rect 3893 1813 3907 1827
rect 3673 1673 3687 1687
rect 3713 1653 3727 1667
rect 3693 1613 3707 1627
rect 3673 1473 3687 1487
rect 3653 1453 3667 1467
rect 3693 1434 3707 1448
rect 3653 1392 3667 1406
rect 3573 1313 3587 1327
rect 3633 1313 3647 1327
rect 3673 1313 3687 1327
rect 3452 1213 3466 1227
rect 3473 1213 3487 1227
rect 3513 1214 3527 1228
rect 3473 1153 3487 1167
rect 3433 993 3447 1007
rect 3413 933 3427 947
rect 3533 1172 3547 1186
rect 3613 1293 3627 1307
rect 3613 1233 3627 1247
rect 3633 1214 3647 1228
rect 3773 1692 3787 1706
rect 3813 1692 3827 1706
rect 3833 1613 3847 1627
rect 3853 1593 3867 1607
rect 3833 1573 3847 1587
rect 4053 2193 4067 2207
rect 4033 2133 4047 2147
rect 4213 2353 4227 2367
rect 4193 2293 4207 2307
rect 4193 2253 4207 2267
rect 4113 2213 4127 2227
rect 4093 2133 4107 2147
rect 4093 2112 4107 2126
rect 4053 2073 4067 2087
rect 4033 1993 4047 2007
rect 4173 2212 4187 2226
rect 4133 2193 4147 2207
rect 4153 2113 4167 2127
rect 4133 2033 4147 2047
rect 4113 1993 4127 2007
rect 4093 1973 4107 1987
rect 4033 1913 4047 1927
rect 3993 1773 4007 1787
rect 3933 1753 3947 1767
rect 3993 1734 4007 1748
rect 3973 1692 3987 1706
rect 3913 1653 3927 1667
rect 3933 1633 3947 1647
rect 3913 1573 3927 1587
rect 3773 1533 3787 1547
rect 3833 1533 3847 1547
rect 3733 1413 3747 1427
rect 3793 1392 3807 1406
rect 3793 1313 3807 1327
rect 3733 1253 3747 1267
rect 3793 1253 3807 1267
rect 3613 1172 3627 1186
rect 3493 1133 3507 1147
rect 3433 914 3447 928
rect 3473 914 3487 928
rect 3433 853 3447 867
rect 3413 833 3427 847
rect 3613 1133 3627 1147
rect 3613 1073 3627 1087
rect 3733 1172 3747 1186
rect 3773 1172 3787 1186
rect 3793 1093 3807 1107
rect 3753 1073 3767 1087
rect 3693 1053 3707 1067
rect 3733 1053 3747 1067
rect 3693 1013 3707 1027
rect 3773 993 3787 1007
rect 3653 953 3667 967
rect 3733 953 3747 967
rect 3533 914 3547 928
rect 3573 914 3587 928
rect 3613 914 3627 928
rect 3513 833 3527 847
rect 3372 753 3386 767
rect 3393 753 3407 767
rect 3353 713 3367 727
rect 3313 694 3327 708
rect 3253 653 3267 667
rect 3233 513 3247 527
rect 3213 493 3227 507
rect 3213 433 3227 447
rect 3153 413 3167 427
rect 3193 413 3207 427
rect 3293 652 3307 666
rect 3333 633 3347 647
rect 3433 813 3447 827
rect 3413 713 3427 727
rect 3473 773 3487 787
rect 3453 713 3467 727
rect 3413 652 3427 666
rect 3373 633 3387 647
rect 3353 613 3367 627
rect 3393 613 3407 627
rect 3453 613 3467 627
rect 3253 473 3267 487
rect 3093 394 3107 408
rect 3133 393 3147 407
rect 3012 353 3026 367
rect 3033 352 3047 366
rect 3073 352 3087 366
rect 3013 253 3027 267
rect 3053 174 3067 188
rect 3253 413 3267 427
rect 3293 413 3307 427
rect 3153 352 3167 366
rect 3173 313 3187 327
rect 3233 352 3247 366
rect 3233 313 3247 327
rect 3353 394 3367 408
rect 3593 872 3607 886
rect 3633 873 3647 887
rect 3593 833 3607 847
rect 3573 773 3587 787
rect 3553 753 3567 767
rect 3693 914 3707 928
rect 3773 913 3787 927
rect 3673 873 3687 887
rect 3653 833 3667 847
rect 3633 813 3647 827
rect 3613 793 3627 807
rect 3593 753 3607 767
rect 3533 694 3547 708
rect 3573 694 3587 708
rect 3633 753 3647 767
rect 3613 693 3627 707
rect 3513 633 3527 647
rect 3473 593 3487 607
rect 3533 573 3547 587
rect 3433 513 3447 527
rect 3473 394 3487 408
rect 3593 652 3607 666
rect 3593 593 3607 607
rect 3693 853 3707 867
rect 3693 773 3707 787
rect 3773 873 3787 887
rect 3753 813 3767 827
rect 3713 753 3727 767
rect 3693 733 3707 747
rect 3833 1133 3847 1147
rect 3873 1473 3887 1487
rect 3873 1392 3887 1406
rect 3933 1392 3947 1406
rect 3953 1373 3967 1387
rect 3893 1313 3907 1327
rect 3873 1293 3887 1307
rect 3873 1213 3887 1227
rect 4013 1673 4027 1687
rect 4113 1873 4127 1887
rect 4173 1954 4187 1968
rect 4253 2413 4267 2427
rect 4233 2293 4247 2307
rect 4413 2613 4427 2627
rect 4613 2933 4627 2947
rect 4673 3073 4687 3087
rect 4953 3073 4967 3087
rect 4913 3053 4927 3067
rect 4713 3033 4727 3047
rect 4673 2994 4687 3008
rect 4713 2994 4727 3008
rect 4753 2994 4767 3008
rect 4793 2994 4807 3008
rect 4693 2933 4707 2947
rect 4633 2913 4647 2927
rect 4873 2953 4887 2967
rect 4933 2952 4947 2966
rect 5073 3294 5087 3308
rect 5193 3553 5207 3567
rect 5193 3514 5207 3528
rect 5233 3514 5247 3528
rect 5173 3473 5187 3487
rect 5033 3252 5047 3266
rect 5113 3252 5127 3266
rect 5093 3153 5107 3167
rect 5073 3033 5087 3047
rect 5013 3013 5027 3027
rect 5033 2994 5047 3008
rect 5213 3472 5227 3486
rect 5253 3473 5267 3487
rect 5253 3433 5267 3447
rect 5433 3992 5447 4006
rect 5533 3973 5547 3987
rect 5573 3973 5587 3987
rect 5513 3893 5527 3907
rect 5433 3873 5447 3887
rect 5413 3814 5427 3828
rect 5473 3814 5487 3828
rect 5393 3753 5407 3767
rect 5333 3733 5347 3747
rect 5313 3593 5327 3607
rect 5353 3573 5367 3587
rect 5393 3513 5407 3527
rect 5453 3772 5467 3786
rect 5433 3733 5447 3747
rect 5513 3733 5527 3747
rect 5333 3472 5347 3486
rect 5413 3473 5427 3487
rect 5693 4673 5707 4687
rect 5693 4593 5707 4607
rect 5653 4554 5667 4568
rect 5713 4553 5727 4567
rect 5713 4513 5727 4527
rect 5673 4473 5687 4487
rect 5613 4453 5627 4467
rect 5673 4433 5687 4447
rect 5653 4413 5667 4427
rect 5693 4393 5707 4407
rect 5672 4373 5686 4387
rect 5673 4293 5687 4307
rect 5673 4033 5687 4047
rect 5633 3993 5647 4007
rect 5673 3993 5687 4007
rect 5653 3973 5667 3987
rect 5593 3913 5607 3927
rect 5573 3893 5587 3907
rect 5573 3693 5587 3707
rect 5613 3653 5627 3667
rect 5593 3573 5607 3587
rect 5553 3553 5567 3567
rect 5533 3533 5547 3547
rect 5493 3472 5507 3486
rect 5193 3413 5207 3427
rect 5273 3413 5287 3427
rect 5173 3313 5187 3327
rect 5353 3393 5367 3407
rect 5273 3353 5287 3367
rect 5233 3333 5247 3347
rect 5233 3294 5247 3308
rect 5213 3252 5227 3266
rect 5153 3233 5167 3247
rect 5133 3033 5147 3047
rect 5133 3012 5147 3026
rect 5113 2993 5127 3007
rect 5013 2953 5027 2967
rect 4813 2913 4827 2927
rect 4993 2913 5007 2927
rect 4753 2893 4767 2907
rect 4813 2892 4827 2906
rect 4593 2833 4607 2847
rect 4633 2833 4647 2847
rect 4753 2833 4767 2847
rect 4793 2833 4807 2847
rect 4593 2774 4607 2788
rect 4773 2813 4787 2827
rect 4733 2774 4747 2788
rect 4833 2873 4847 2887
rect 4813 2773 4827 2787
rect 4693 2753 4707 2767
rect 4453 2733 4467 2747
rect 4433 2573 4447 2587
rect 4413 2553 4427 2567
rect 4353 2473 4367 2487
rect 4393 2474 4407 2488
rect 4473 2713 4487 2727
rect 4553 2733 4567 2747
rect 4533 2693 4547 2707
rect 4513 2673 4527 2687
rect 4473 2573 4487 2587
rect 4333 2413 4347 2427
rect 4373 2393 4387 2407
rect 4353 2373 4367 2387
rect 4333 2353 4347 2367
rect 4273 2293 4287 2307
rect 4333 2273 4347 2287
rect 4293 2254 4307 2268
rect 4333 2213 4347 2227
rect 4333 2173 4347 2187
rect 4313 2153 4327 2167
rect 4273 2133 4287 2147
rect 4273 2073 4287 2087
rect 4313 2073 4327 2087
rect 4232 1953 4246 1967
rect 4253 1953 4267 1967
rect 4293 1954 4307 1968
rect 4333 1953 4347 1967
rect 4153 1913 4167 1927
rect 4133 1853 4147 1867
rect 4113 1833 4127 1847
rect 4133 1813 4147 1827
rect 4133 1773 4147 1787
rect 4113 1753 4127 1767
rect 4073 1734 4087 1748
rect 4113 1734 4127 1748
rect 4053 1653 4067 1667
rect 4033 1513 4047 1527
rect 4093 1692 4107 1706
rect 4093 1473 4107 1487
rect 4013 1373 4027 1387
rect 3952 1273 3966 1287
rect 3973 1273 3987 1287
rect 3993 1253 4007 1267
rect 3933 1214 3947 1228
rect 3873 1172 3887 1186
rect 3853 1093 3867 1107
rect 3813 1053 3827 1067
rect 3853 1053 3867 1067
rect 3813 913 3827 927
rect 3953 1172 3967 1186
rect 3953 1113 3967 1127
rect 3973 1073 3987 1087
rect 4133 1613 4147 1627
rect 4193 1912 4207 1926
rect 4233 1893 4247 1907
rect 4273 1913 4287 1927
rect 4253 1853 4267 1867
rect 4253 1832 4267 1846
rect 4173 1733 4187 1747
rect 4213 1734 4227 1748
rect 4313 1912 4327 1926
rect 4453 2413 4467 2427
rect 4413 2353 4427 2367
rect 4393 2254 4407 2268
rect 4513 2493 4527 2507
rect 4593 2633 4607 2647
rect 4573 2493 4587 2507
rect 4553 2432 4567 2446
rect 4673 2733 4687 2747
rect 4653 2693 4667 2707
rect 4693 2633 4707 2647
rect 4613 2573 4627 2587
rect 4673 2573 4687 2587
rect 4773 2713 4787 2727
rect 4753 2553 4767 2567
rect 4613 2533 4627 2547
rect 4733 2533 4747 2547
rect 4613 2473 4627 2487
rect 4653 2474 4667 2488
rect 4753 2493 4767 2507
rect 4813 2733 4827 2747
rect 4793 2553 4807 2567
rect 4713 2473 4727 2487
rect 4513 2413 4527 2427
rect 4373 2173 4387 2187
rect 4413 2133 4427 2147
rect 4393 2113 4407 2127
rect 4373 2053 4387 2067
rect 4393 2033 4407 2047
rect 4373 1993 4387 2007
rect 4473 2172 4487 2186
rect 4473 2093 4487 2107
rect 4473 2013 4487 2027
rect 4373 1953 4387 1967
rect 4433 1954 4447 1968
rect 4593 2413 4607 2427
rect 4573 2393 4587 2407
rect 4573 2333 4587 2347
rect 4633 2432 4647 2446
rect 4773 2432 4787 2446
rect 4893 2833 4907 2847
rect 5073 2933 5087 2947
rect 5053 2913 5067 2927
rect 5053 2833 5067 2847
rect 4913 2812 4927 2826
rect 4953 2813 4967 2827
rect 5013 2813 5027 2827
rect 4933 2793 4947 2807
rect 4873 2774 4887 2788
rect 4853 2733 4867 2747
rect 4913 2732 4927 2746
rect 5033 2713 5047 2727
rect 4853 2693 4867 2707
rect 4973 2633 4987 2647
rect 4953 2573 4967 2587
rect 4913 2553 4927 2567
rect 4873 2533 4887 2547
rect 4913 2474 4927 2488
rect 4733 2413 4747 2427
rect 4833 2413 4847 2427
rect 4692 2373 4706 2387
rect 4713 2373 4727 2387
rect 4613 2353 4627 2367
rect 4673 2353 4687 2367
rect 4553 2293 4567 2307
rect 4553 2254 4567 2268
rect 4533 2113 4547 2127
rect 4573 2173 4587 2187
rect 4553 2073 4567 2087
rect 4533 2033 4547 2047
rect 4593 2113 4607 2127
rect 4593 2053 4607 2067
rect 4573 2013 4587 2027
rect 4493 1953 4507 1967
rect 4553 1954 4567 1968
rect 4673 2332 4687 2346
rect 4633 2293 4647 2307
rect 4673 2254 4687 2268
rect 4713 2212 4727 2226
rect 4653 2153 4667 2167
rect 4753 2254 4767 2268
rect 4813 2254 4827 2268
rect 4853 2254 4867 2268
rect 4893 2393 4907 2407
rect 5253 3213 5267 3227
rect 5213 3193 5227 3207
rect 5213 3033 5227 3047
rect 5313 3294 5327 3308
rect 5273 3153 5287 3167
rect 5393 3252 5407 3266
rect 5313 3013 5327 3027
rect 5373 3013 5387 3027
rect 5353 2994 5367 3008
rect 5153 2933 5167 2947
rect 5133 2873 5147 2887
rect 5113 2793 5127 2807
rect 5153 2793 5167 2807
rect 5133 2774 5147 2788
rect 5213 2933 5227 2947
rect 5093 2733 5107 2747
rect 5113 2732 5127 2746
rect 5173 2732 5187 2746
rect 5193 2733 5207 2747
rect 5073 2713 5087 2727
rect 5133 2713 5147 2727
rect 5073 2653 5087 2667
rect 4993 2513 5007 2527
rect 5053 2513 5067 2527
rect 4973 2413 4987 2427
rect 4933 2333 4947 2347
rect 4893 2313 4907 2327
rect 4833 2212 4847 2226
rect 4873 2213 4887 2227
rect 4853 2173 4867 2187
rect 4793 2133 4807 2147
rect 4753 2113 4767 2127
rect 4693 2033 4707 2047
rect 4653 2013 4667 2027
rect 4673 1993 4687 2007
rect 4513 1932 4527 1946
rect 4373 1893 4387 1907
rect 4413 1893 4427 1907
rect 4493 1913 4507 1927
rect 4453 1893 4467 1907
rect 4293 1813 4307 1827
rect 4273 1773 4287 1787
rect 4273 1734 4287 1748
rect 4172 1693 4186 1707
rect 4153 1553 4167 1567
rect 4193 1692 4207 1706
rect 4213 1673 4227 1687
rect 4473 1873 4487 1887
rect 4433 1853 4447 1867
rect 4413 1833 4427 1847
rect 4313 1753 4327 1767
rect 4373 1753 4387 1767
rect 4353 1734 4367 1748
rect 4393 1734 4407 1748
rect 4233 1653 4247 1667
rect 4293 1653 4307 1667
rect 4413 1693 4427 1707
rect 4373 1633 4387 1647
rect 4333 1613 4347 1627
rect 4253 1573 4267 1587
rect 4173 1533 4187 1547
rect 4213 1473 4227 1487
rect 4173 1434 4187 1448
rect 4113 1373 4127 1387
rect 4113 1333 4127 1347
rect 4153 1392 4167 1406
rect 4232 1434 4246 1448
rect 4333 1572 4347 1586
rect 4293 1513 4307 1527
rect 4153 1371 4167 1385
rect 4213 1373 4227 1387
rect 4133 1313 4147 1327
rect 4133 1253 4147 1267
rect 4113 1233 4127 1247
rect 4053 1213 4067 1227
rect 4093 1214 4107 1228
rect 4053 1153 4067 1167
rect 3993 1053 4007 1067
rect 4013 1033 4027 1047
rect 3893 1013 3907 1027
rect 3973 1013 3987 1027
rect 3873 953 3887 967
rect 3933 973 3947 987
rect 3953 953 3967 967
rect 3953 913 3967 927
rect 4013 914 4027 928
rect 3873 872 3887 886
rect 3932 872 3946 886
rect 3953 873 3967 887
rect 3833 853 3847 867
rect 3993 872 4007 886
rect 3853 833 3867 847
rect 3953 833 3967 847
rect 3813 813 3827 827
rect 3793 733 3807 747
rect 3873 793 3887 807
rect 3673 652 3687 666
rect 3713 652 3727 666
rect 3633 573 3647 587
rect 3553 553 3567 567
rect 3573 413 3587 427
rect 3853 693 3867 707
rect 4013 753 4027 767
rect 3993 733 4007 747
rect 3933 694 3947 708
rect 3833 652 3847 666
rect 3873 652 3887 666
rect 3913 652 3927 666
rect 3793 493 3807 507
rect 3973 653 3987 667
rect 4073 1013 4087 1027
rect 4073 913 4087 927
rect 4113 914 4127 928
rect 4253 1433 4267 1447
rect 4473 1773 4487 1787
rect 4513 1873 4527 1887
rect 4553 1873 4567 1887
rect 4533 1793 4547 1807
rect 4513 1734 4527 1748
rect 4453 1693 4467 1707
rect 4453 1653 4467 1667
rect 4433 1633 4447 1647
rect 4413 1573 4427 1587
rect 4393 1553 4407 1567
rect 4352 1533 4366 1547
rect 4373 1533 4387 1547
rect 4333 1452 4347 1466
rect 4373 1493 4387 1507
rect 4413 1513 4427 1527
rect 4353 1433 4367 1447
rect 4273 1392 4287 1406
rect 4273 1353 4287 1367
rect 4253 1333 4267 1347
rect 4233 1313 4247 1327
rect 4253 1293 4267 1307
rect 4193 1273 4207 1287
rect 4173 1172 4187 1186
rect 4193 1153 4207 1167
rect 4253 1153 4267 1167
rect 4293 1313 4307 1327
rect 4533 1692 4547 1706
rect 4493 1613 4507 1627
rect 4493 1573 4507 1587
rect 4473 1473 4487 1487
rect 4413 1434 4427 1448
rect 4393 1393 4407 1407
rect 4373 1353 4387 1367
rect 4313 1273 4327 1287
rect 4333 1214 4347 1228
rect 4313 1172 4327 1186
rect 4373 1173 4387 1187
rect 4373 1133 4387 1147
rect 4353 1113 4367 1127
rect 4293 1093 4307 1107
rect 4273 1073 4287 1087
rect 4193 1033 4207 1047
rect 4213 993 4227 1007
rect 4213 953 4227 967
rect 4093 872 4107 886
rect 4213 914 4227 928
rect 4153 793 4167 807
rect 4053 733 4067 747
rect 4153 733 4167 747
rect 4073 694 4087 708
rect 4113 694 4127 708
rect 4013 652 4027 666
rect 4053 652 4067 666
rect 4133 653 4147 667
rect 3993 593 4007 607
rect 3973 573 3987 587
rect 4233 872 4247 886
rect 4433 1392 4447 1406
rect 4453 1333 4467 1347
rect 4673 1954 4687 1968
rect 4713 1954 4727 1968
rect 4773 2033 4787 2047
rect 4813 2033 4827 2047
rect 4693 1873 4707 1887
rect 4793 1993 4807 2007
rect 4793 1954 4807 1968
rect 5153 2693 5167 2707
rect 5213 2693 5227 2707
rect 5133 2633 5147 2647
rect 5093 2513 5107 2527
rect 5073 2493 5087 2507
rect 5053 2474 5067 2488
rect 4953 2293 4967 2307
rect 4993 2293 5007 2307
rect 4993 2254 5007 2268
rect 5073 2432 5087 2446
rect 5113 2432 5127 2446
rect 5053 2413 5067 2427
rect 5033 2333 5047 2347
rect 5033 2293 5047 2307
rect 4893 2133 4907 2147
rect 4973 2212 4987 2226
rect 4993 2173 5007 2187
rect 4933 2113 4947 2127
rect 4873 2073 4887 2087
rect 4873 2033 4887 2047
rect 4853 1993 4867 2007
rect 4913 1993 4927 2007
rect 4853 1954 4867 1968
rect 4773 1873 4787 1887
rect 4733 1853 4747 1867
rect 4713 1793 4727 1807
rect 4753 1773 4767 1787
rect 4633 1753 4647 1767
rect 4673 1753 4687 1767
rect 4713 1754 4727 1768
rect 4613 1734 4627 1748
rect 4573 1633 4587 1647
rect 4633 1692 4647 1706
rect 4593 1573 4607 1587
rect 4553 1533 4567 1547
rect 4653 1533 4667 1547
rect 4613 1513 4627 1527
rect 4713 1733 4727 1747
rect 4833 1912 4847 1926
rect 4873 1912 4887 1926
rect 4873 1833 4887 1847
rect 4833 1793 4847 1807
rect 4953 2033 4967 2047
rect 4993 1993 5007 2007
rect 4953 1953 4967 1967
rect 4993 1954 5007 1968
rect 4973 1912 4987 1926
rect 4953 1813 4967 1827
rect 4933 1753 4947 1767
rect 4693 1673 4707 1687
rect 4633 1473 4647 1487
rect 4673 1473 4687 1487
rect 4613 1453 4627 1467
rect 4513 1433 4527 1447
rect 4573 1434 4587 1448
rect 4593 1393 4607 1407
rect 4593 1353 4607 1367
rect 4553 1333 4567 1347
rect 4493 1313 4507 1327
rect 4533 1313 4547 1327
rect 4473 1293 4487 1307
rect 4493 1233 4507 1247
rect 4733 1573 4747 1587
rect 4733 1493 4747 1507
rect 4633 1433 4647 1447
rect 4713 1453 4727 1467
rect 4753 1473 4767 1487
rect 4733 1433 4747 1447
rect 4633 1393 4647 1407
rect 4613 1273 4627 1287
rect 4653 1333 4667 1347
rect 4593 1253 4607 1267
rect 4633 1253 4647 1267
rect 4673 1253 4687 1267
rect 4593 1214 4607 1228
rect 4633 1214 4647 1228
rect 4433 1172 4447 1186
rect 4393 1113 4407 1127
rect 4552 1172 4566 1186
rect 4573 1173 4587 1187
rect 4513 1113 4527 1127
rect 4553 1113 4567 1127
rect 4473 1093 4487 1107
rect 4653 1133 4667 1147
rect 4613 1093 4627 1107
rect 4473 1053 4487 1067
rect 4573 1053 4587 1067
rect 4473 1013 4487 1027
rect 4573 1013 4587 1027
rect 4613 1013 4627 1027
rect 4393 993 4407 1007
rect 4333 933 4347 947
rect 4333 914 4347 928
rect 4513 993 4527 1007
rect 4733 1393 4747 1407
rect 4733 1233 4747 1247
rect 4813 1693 4827 1707
rect 4853 1673 4867 1687
rect 4913 1693 4927 1707
rect 4893 1633 4907 1647
rect 4813 1493 4827 1507
rect 4893 1434 4907 1448
rect 4793 1392 4807 1406
rect 4812 1333 4826 1347
rect 4833 1333 4847 1347
rect 4752 1213 4766 1227
rect 4773 1213 4787 1227
rect 4713 1173 4727 1187
rect 4713 1133 4727 1147
rect 4853 1253 4867 1267
rect 4813 1213 4827 1227
rect 5133 2393 5147 2407
rect 5473 3433 5487 3447
rect 5493 3353 5507 3367
rect 5413 3213 5427 3227
rect 5453 3213 5467 3227
rect 5553 3513 5567 3527
rect 5613 3553 5627 3567
rect 5633 3532 5647 3546
rect 5673 3913 5687 3927
rect 5793 4812 5807 4826
rect 5793 4433 5807 4447
rect 5753 4373 5767 4387
rect 5793 4334 5807 4348
rect 5833 4333 5847 4347
rect 5733 4293 5747 4307
rect 5833 4293 5847 4307
rect 5733 4253 5747 4267
rect 5773 4253 5787 4267
rect 5753 4093 5767 4107
rect 5733 4033 5747 4047
rect 5813 4273 5827 4287
rect 5793 3993 5807 4007
rect 5753 3973 5767 3987
rect 5713 3873 5727 3887
rect 5693 3833 5707 3847
rect 5713 3814 5727 3828
rect 5773 3873 5787 3887
rect 5673 3773 5687 3787
rect 5733 3772 5747 3786
rect 5693 3653 5707 3667
rect 5673 3512 5687 3526
rect 5753 3514 5767 3528
rect 5793 3772 5807 3786
rect 5793 3733 5807 3747
rect 5613 3472 5627 3486
rect 5813 3633 5827 3647
rect 5573 3433 5587 3447
rect 5653 3393 5667 3407
rect 5733 3472 5747 3486
rect 5793 3473 5807 3487
rect 5693 3353 5707 3367
rect 5733 3353 5747 3367
rect 5553 3294 5567 3308
rect 5693 3294 5707 3308
rect 5493 3013 5507 3027
rect 5533 3013 5547 3027
rect 5413 2993 5427 3007
rect 5473 2994 5487 3008
rect 5493 2952 5507 2966
rect 5333 2873 5347 2887
rect 5413 2873 5427 2887
rect 5293 2833 5307 2847
rect 5293 2793 5307 2807
rect 5253 2732 5267 2746
rect 5313 2693 5327 2707
rect 5533 2933 5547 2947
rect 5593 3252 5607 3266
rect 5573 3213 5587 3227
rect 5693 3073 5707 3087
rect 5633 3033 5647 3047
rect 5653 2993 5667 3007
rect 5613 2952 5627 2966
rect 5653 2952 5667 2966
rect 5493 2893 5507 2907
rect 5553 2893 5567 2907
rect 5673 2893 5687 2907
rect 5473 2873 5487 2887
rect 5453 2833 5467 2847
rect 5413 2813 5427 2827
rect 5393 2732 5407 2746
rect 5433 2693 5447 2707
rect 5393 2653 5407 2667
rect 5333 2633 5347 2647
rect 5453 2633 5467 2647
rect 5213 2474 5227 2488
rect 5193 2432 5207 2446
rect 5193 2373 5207 2387
rect 5153 2333 5167 2347
rect 5193 2333 5207 2347
rect 5113 2293 5127 2307
rect 5153 2254 5167 2268
rect 5053 2212 5067 2226
rect 5073 2153 5087 2167
rect 5133 2212 5147 2226
rect 5272 2513 5286 2527
rect 5293 2513 5307 2527
rect 5273 2474 5287 2488
rect 5313 2474 5327 2488
rect 5433 2473 5447 2487
rect 5413 2432 5427 2446
rect 5253 2413 5267 2427
rect 5293 2412 5307 2426
rect 5253 2373 5267 2387
rect 5253 2293 5267 2307
rect 5253 2254 5267 2268
rect 5553 2833 5567 2847
rect 5813 3073 5827 3087
rect 5773 3033 5787 3047
rect 5733 2994 5747 3008
rect 5773 2994 5787 3008
rect 5813 2994 5827 3008
rect 5753 2933 5767 2947
rect 5693 2833 5707 2847
rect 5793 2833 5807 2847
rect 5653 2774 5667 2788
rect 5733 2774 5747 2788
rect 5493 2733 5507 2747
rect 5513 2713 5527 2727
rect 5633 2693 5647 2707
rect 5553 2673 5567 2687
rect 5653 2673 5667 2687
rect 5553 2533 5567 2547
rect 5513 2493 5527 2507
rect 5473 2473 5487 2487
rect 5533 2474 5547 2488
rect 5593 2474 5607 2488
rect 5633 2474 5647 2488
rect 5753 2713 5767 2727
rect 5753 2653 5767 2667
rect 5753 2593 5767 2607
rect 5753 2533 5767 2547
rect 5733 2474 5747 2488
rect 5773 2473 5787 2487
rect 5333 2373 5347 2387
rect 5333 2333 5347 2347
rect 5433 2393 5447 2407
rect 5433 2333 5447 2347
rect 5413 2313 5427 2327
rect 5333 2293 5347 2307
rect 5373 2293 5387 2307
rect 5373 2272 5387 2286
rect 5293 2253 5307 2267
rect 5333 2253 5347 2267
rect 5493 2432 5507 2446
rect 5513 2353 5527 2367
rect 5493 2333 5507 2347
rect 5553 2432 5567 2446
rect 5533 2313 5547 2327
rect 5473 2293 5487 2307
rect 5513 2293 5527 2307
rect 5453 2273 5467 2287
rect 5153 2133 5167 2147
rect 5133 2113 5147 2127
rect 5093 2073 5107 2087
rect 5093 2033 5107 2047
rect 5133 2033 5147 2047
rect 5073 2013 5087 2027
rect 5053 1993 5067 2007
rect 5113 1973 5127 1987
rect 5053 1953 5067 1967
rect 5093 1954 5107 1968
rect 5153 2013 5167 2027
rect 5153 1953 5167 1967
rect 5073 1873 5087 1887
rect 5093 1853 5107 1867
rect 5053 1793 5067 1807
rect 5033 1754 5047 1768
rect 5033 1733 5047 1747
rect 4953 1533 4967 1547
rect 5013 1692 5027 1706
rect 5033 1673 5047 1687
rect 4973 1513 4987 1527
rect 5013 1513 5027 1527
rect 4993 1493 5007 1507
rect 5013 1473 5027 1487
rect 4993 1453 5007 1467
rect 4953 1434 4967 1448
rect 4993 1392 5007 1406
rect 5033 1353 5047 1367
rect 4953 1253 4967 1267
rect 5013 1253 5027 1267
rect 4813 1173 4827 1187
rect 4733 1093 4747 1107
rect 4793 1093 4807 1107
rect 4753 993 4767 1007
rect 4693 953 4707 967
rect 4613 933 4627 947
rect 4633 914 4647 928
rect 4673 912 4687 926
rect 4713 914 4727 928
rect 4353 872 4367 886
rect 4293 813 4307 827
rect 4273 753 4287 767
rect 4193 694 4207 708
rect 4233 694 4247 708
rect 4533 872 4547 886
rect 4573 872 4587 886
rect 4613 872 4627 886
rect 4433 853 4447 867
rect 4493 853 4507 867
rect 4273 693 4287 707
rect 4253 553 4267 567
rect 4373 694 4387 708
rect 4313 653 4327 667
rect 4293 513 4307 527
rect 4093 473 4107 487
rect 4133 473 4147 487
rect 3833 453 3847 467
rect 3893 453 3907 467
rect 3613 394 3627 408
rect 3653 394 3667 408
rect 3713 394 3727 408
rect 3753 394 3767 408
rect 3453 352 3467 366
rect 3333 333 3347 347
rect 3193 273 3207 287
rect 3293 273 3307 287
rect 3173 253 3187 267
rect 3313 253 3327 267
rect 3393 253 3407 267
rect 3253 233 3267 247
rect 3253 174 3267 188
rect 3053 113 3067 127
rect 3033 93 3047 107
rect 3013 33 3027 47
rect 3213 132 3227 146
rect 3253 133 3267 147
rect 3173 113 3187 127
rect 3533 353 3547 367
rect 3593 352 3607 366
rect 3633 353 3647 367
rect 3553 253 3567 267
rect 3493 233 3507 247
rect 3513 173 3527 187
rect 3593 213 3607 227
rect 3633 173 3647 187
rect 3293 132 3307 146
rect 3273 93 3287 107
rect 3393 132 3407 146
rect 3433 132 3447 146
rect 3793 393 3807 407
rect 3853 394 3867 408
rect 3793 352 3807 366
rect 3833 352 3847 366
rect 3813 293 3827 307
rect 3733 253 3747 267
rect 3693 213 3707 227
rect 3733 174 3747 188
rect 3773 174 3787 188
rect 3613 93 3627 107
rect 3653 93 3667 107
rect 3073 73 3087 87
rect 3353 73 3367 87
rect 3473 73 3487 87
rect 3573 73 3587 87
rect 3053 53 3067 67
rect 3753 132 3767 146
rect 3073 33 3087 47
rect 3713 33 3727 47
rect 2993 13 3007 27
rect 3973 433 3987 447
rect 4053 433 4067 447
rect 3913 393 3927 407
rect 4013 394 4027 408
rect 3913 352 3927 366
rect 3953 352 3967 366
rect 4113 433 4127 447
rect 4293 433 4307 447
rect 4153 394 4167 408
rect 4253 394 4267 408
rect 4353 652 4367 666
rect 4393 652 4407 666
rect 4573 793 4587 807
rect 4633 793 4647 807
rect 4533 753 4547 767
rect 4453 713 4467 727
rect 4493 694 4507 708
rect 4373 553 4387 567
rect 4353 433 4367 447
rect 3893 293 3907 307
rect 3893 253 3907 267
rect 3853 174 3867 188
rect 3953 193 3967 207
rect 4233 352 4247 366
rect 4133 313 4147 327
rect 4313 353 4327 367
rect 4273 313 4287 327
rect 4313 273 4327 287
rect 4233 253 4247 267
rect 4293 233 4307 247
rect 4293 193 4307 207
rect 3833 132 3847 146
rect 3873 132 3887 146
rect 3913 132 3927 146
rect 3913 93 3927 107
rect 3993 174 4007 188
rect 4033 174 4047 188
rect 4093 174 4107 188
rect 3973 132 3987 146
rect 4013 132 4027 146
rect 4053 132 4067 146
rect 3953 33 3967 47
rect 4173 174 4187 188
rect 4233 173 4247 187
rect 4273 174 4287 188
rect 4433 652 4447 666
rect 4373 393 4387 407
rect 4513 652 4527 666
rect 4733 872 4747 886
rect 4773 872 4787 886
rect 4873 1172 4887 1186
rect 4833 1113 4847 1127
rect 4893 1073 4907 1087
rect 4933 1213 4947 1227
rect 4973 1214 4987 1228
rect 5153 1913 5167 1927
rect 5153 1853 5167 1867
rect 5113 1813 5127 1827
rect 5233 2173 5247 2187
rect 5193 2153 5207 2167
rect 5193 2093 5207 2107
rect 5193 2053 5207 2067
rect 5233 1993 5247 2007
rect 5193 1953 5207 1967
rect 5273 1954 5287 1968
rect 5313 2213 5327 2227
rect 5393 2212 5407 2226
rect 5433 2213 5447 2227
rect 5393 2193 5407 2207
rect 5333 2173 5347 2187
rect 5313 2113 5327 2127
rect 5313 2033 5327 2047
rect 5353 2133 5367 2147
rect 5333 2013 5347 2027
rect 5333 1973 5347 1987
rect 5253 1912 5267 1926
rect 5213 1893 5227 1907
rect 5233 1873 5247 1887
rect 5113 1773 5127 1787
rect 5173 1773 5187 1787
rect 5153 1734 5167 1748
rect 5533 2273 5547 2287
rect 5593 2393 5607 2407
rect 5573 2353 5587 2367
rect 5573 2313 5587 2327
rect 5573 2292 5587 2306
rect 5573 2253 5587 2267
rect 5533 2212 5547 2226
rect 5493 2173 5507 2187
rect 5453 2133 5467 2147
rect 5452 2112 5466 2126
rect 5473 2113 5487 2127
rect 5433 2093 5447 2107
rect 5353 1954 5367 1968
rect 5353 1893 5367 1907
rect 5313 1873 5327 1887
rect 5253 1793 5267 1807
rect 5293 1793 5307 1807
rect 5213 1733 5227 1747
rect 5333 1853 5347 1867
rect 5333 1813 5347 1827
rect 5313 1753 5327 1767
rect 5293 1734 5307 1748
rect 5093 1673 5107 1687
rect 5173 1692 5187 1706
rect 5213 1692 5227 1706
rect 5193 1673 5207 1687
rect 5133 1633 5147 1647
rect 5093 1613 5107 1627
rect 5193 1573 5207 1587
rect 5233 1573 5247 1587
rect 5113 1553 5127 1567
rect 5153 1473 5167 1487
rect 5193 1434 5207 1448
rect 5073 1353 5087 1367
rect 5173 1392 5187 1406
rect 5133 1373 5147 1387
rect 5113 1333 5127 1347
rect 5093 1313 5107 1327
rect 5133 1253 5147 1267
rect 5113 1233 5127 1247
rect 4913 1033 4927 1047
rect 4933 1013 4947 1027
rect 4833 914 4847 928
rect 4873 914 4887 928
rect 4833 873 4847 887
rect 4893 853 4907 867
rect 4833 833 4847 847
rect 4813 793 4827 807
rect 4853 753 4867 767
rect 4913 753 4927 767
rect 4673 714 4687 728
rect 4713 713 4727 727
rect 4673 693 4687 707
rect 4493 553 4507 567
rect 4573 553 4587 567
rect 4413 352 4427 366
rect 4353 313 4367 327
rect 4333 213 4347 227
rect 4653 613 4667 627
rect 4613 533 4627 547
rect 4553 473 4567 487
rect 4753 694 4767 708
rect 4793 694 4807 708
rect 4753 593 4767 607
rect 4633 433 4647 447
rect 4713 433 4727 447
rect 4593 394 4607 408
rect 4513 352 4527 366
rect 4493 333 4507 347
rect 4573 352 4587 366
rect 4533 313 4547 327
rect 4453 293 4467 307
rect 4513 293 4527 307
rect 4373 253 4387 267
rect 4353 173 4367 187
rect 4153 132 4167 146
rect 4193 132 4207 146
rect 4293 132 4307 146
rect 4333 132 4347 146
rect 4433 253 4447 267
rect 4393 173 4407 187
rect 4513 233 4527 247
rect 4473 193 4487 207
rect 4413 132 4427 146
rect 4492 133 4506 147
rect 4613 193 4627 207
rect 4573 174 4587 188
rect 4613 174 4627 188
rect 4813 652 4827 666
rect 4993 1172 5007 1186
rect 5093 1214 5107 1228
rect 4993 993 5007 1007
rect 5053 993 5067 1007
rect 5053 953 5067 967
rect 4973 913 4987 927
rect 5013 914 5027 928
rect 5093 914 5107 928
rect 5153 1172 5167 1186
rect 5153 1073 5167 1087
rect 5173 1053 5187 1067
rect 5133 914 5147 928
rect 5253 1353 5267 1367
rect 5312 1653 5326 1667
rect 5333 1653 5347 1667
rect 5373 1853 5387 1867
rect 5433 1913 5447 1927
rect 5413 1833 5427 1847
rect 5373 1813 5387 1827
rect 5413 1812 5427 1826
rect 5513 2053 5527 2067
rect 5473 1953 5487 1967
rect 5573 2113 5587 2127
rect 5533 1973 5547 1987
rect 5553 1954 5567 1968
rect 5653 2432 5667 2446
rect 5692 2433 5706 2447
rect 5713 2433 5727 2447
rect 5613 2353 5627 2367
rect 5673 2353 5687 2367
rect 5613 2313 5627 2327
rect 5633 2293 5647 2307
rect 5693 2293 5707 2307
rect 5613 2212 5627 2226
rect 5593 1933 5607 1947
rect 5493 1912 5507 1926
rect 5453 1833 5467 1847
rect 5433 1753 5447 1767
rect 5453 1734 5467 1748
rect 5393 1692 5407 1706
rect 5393 1633 5407 1647
rect 5573 1913 5587 1927
rect 5533 1833 5547 1847
rect 5573 1813 5587 1827
rect 5533 1793 5547 1807
rect 5633 2193 5647 2207
rect 5733 2293 5747 2307
rect 5713 2193 5727 2207
rect 5673 2133 5687 2147
rect 5713 1973 5727 1987
rect 5693 1893 5707 1907
rect 5653 1853 5667 1867
rect 5653 1813 5667 1827
rect 5613 1773 5627 1787
rect 5573 1734 5587 1748
rect 5633 1734 5647 1748
rect 5693 1753 5707 1767
rect 5513 1693 5527 1707
rect 5673 1734 5687 1748
rect 5713 1733 5727 1747
rect 5493 1653 5507 1667
rect 5513 1633 5527 1647
rect 5433 1593 5447 1607
rect 5353 1573 5367 1587
rect 5413 1573 5427 1587
rect 5393 1453 5407 1467
rect 5293 1434 5307 1448
rect 5373 1392 5387 1406
rect 5553 1553 5567 1567
rect 5533 1533 5547 1547
rect 5493 1513 5507 1527
rect 5533 1493 5547 1507
rect 5472 1473 5486 1487
rect 5493 1473 5507 1487
rect 5433 1434 5447 1448
rect 5453 1392 5467 1406
rect 5313 1373 5327 1387
rect 5373 1353 5387 1367
rect 5433 1353 5447 1367
rect 5273 1333 5287 1347
rect 5313 1333 5327 1347
rect 5213 1233 5227 1247
rect 5273 1214 5287 1228
rect 5213 1173 5227 1187
rect 5213 1133 5227 1147
rect 5253 1133 5267 1147
rect 5333 1253 5347 1267
rect 5333 1213 5347 1227
rect 5413 1214 5427 1228
rect 5353 1172 5367 1186
rect 5313 1093 5327 1107
rect 5253 1073 5267 1087
rect 5353 1073 5367 1087
rect 5193 1033 5207 1047
rect 5233 993 5247 1007
rect 4993 872 5007 886
rect 5033 872 5047 886
rect 4973 853 4987 867
rect 5013 853 5027 867
rect 5153 853 5167 867
rect 5153 813 5167 827
rect 5112 753 5126 767
rect 5133 753 5147 767
rect 5073 733 5087 747
rect 5093 713 5107 727
rect 4913 694 4927 708
rect 4953 694 4967 708
rect 4993 693 5007 707
rect 5053 694 5067 708
rect 4853 593 4867 607
rect 4933 652 4947 666
rect 4913 613 4927 627
rect 4773 573 4787 587
rect 4893 573 4907 587
rect 4913 553 4927 567
rect 4953 533 4967 547
rect 4813 433 4827 447
rect 4713 394 4727 408
rect 4753 394 4767 408
rect 4693 352 4707 366
rect 4693 293 4707 307
rect 4673 253 4687 267
rect 4853 394 4867 408
rect 4893 394 4907 408
rect 4833 352 4847 366
rect 4893 353 4907 367
rect 5433 1173 5447 1187
rect 5433 1133 5447 1147
rect 5393 1053 5407 1067
rect 5513 1353 5527 1367
rect 5493 1313 5507 1327
rect 5473 1233 5487 1247
rect 5453 1113 5467 1127
rect 5353 1033 5367 1047
rect 5433 1033 5447 1047
rect 5313 953 5327 967
rect 5273 914 5287 928
rect 5313 914 5327 928
rect 5233 813 5247 827
rect 5193 753 5207 767
rect 5173 713 5187 727
rect 5213 694 5227 708
rect 5293 793 5307 807
rect 5293 733 5307 747
rect 5273 713 5287 727
rect 4933 352 4947 366
rect 4993 352 5007 366
rect 4793 293 4807 307
rect 4733 253 4747 267
rect 4773 253 4787 267
rect 4873 253 4887 267
rect 4793 233 4807 247
rect 4693 213 4707 227
rect 4733 213 4747 227
rect 4093 93 4107 107
rect 4373 93 4387 107
rect 4453 93 4467 107
rect 4073 73 4087 87
rect 4513 132 4527 146
rect 4553 132 4567 146
rect 4593 93 4607 107
rect 4693 174 4707 188
rect 5073 652 5087 666
rect 5133 652 5147 666
rect 5053 394 5067 408
rect 5093 394 5107 408
rect 5133 394 5147 408
rect 5073 352 5087 366
rect 5113 333 5127 347
rect 5013 313 5027 327
rect 4973 273 4987 287
rect 4753 132 4767 146
rect 4793 132 4807 146
rect 4713 113 4727 127
rect 4893 113 4907 127
rect 4653 73 4667 87
rect 4833 73 4847 87
rect 5053 233 5067 247
rect 5133 233 5147 247
rect 5073 213 5087 227
rect 5013 174 5027 188
rect 5053 173 5067 187
rect 4933 153 4947 167
rect 4993 132 5007 146
rect 4933 113 4947 127
rect 4973 111 4987 125
rect 5193 652 5207 666
rect 5213 513 5227 527
rect 5293 693 5307 707
rect 5373 973 5387 987
rect 5573 1434 5587 1448
rect 5653 1673 5667 1687
rect 5713 1693 5727 1707
rect 5693 1673 5707 1687
rect 5653 1434 5667 1448
rect 5813 2693 5827 2707
rect 5813 2653 5827 2667
rect 5793 2273 5807 2287
rect 5753 2254 5767 2268
rect 5793 2212 5807 2226
rect 5753 2193 5767 2207
rect 5773 2173 5787 2187
rect 5753 2153 5767 2167
rect 5773 2133 5787 2147
rect 5833 2613 5847 2627
rect 5833 2473 5847 2487
rect 5833 2433 5847 2447
rect 5833 2313 5847 2327
rect 5833 2273 5847 2287
rect 5733 1493 5747 1507
rect 5813 1952 5827 1966
rect 5793 1933 5807 1947
rect 5773 1773 5787 1787
rect 5813 1893 5827 1907
rect 5813 1853 5827 1867
rect 5793 1553 5807 1567
rect 5773 1434 5787 1448
rect 5813 1433 5827 1447
rect 5593 1392 5607 1406
rect 5693 1392 5707 1406
rect 5653 1373 5667 1387
rect 5633 1313 5647 1327
rect 5533 1293 5547 1307
rect 5613 1293 5627 1307
rect 5513 1273 5527 1287
rect 5553 1253 5567 1267
rect 5633 1273 5647 1287
rect 5673 1313 5687 1327
rect 5613 1233 5627 1247
rect 5653 1233 5667 1247
rect 5593 1093 5607 1107
rect 5493 973 5507 987
rect 5473 933 5487 947
rect 5393 872 5407 886
rect 5433 872 5447 886
rect 5393 833 5407 847
rect 5373 793 5387 807
rect 5353 753 5367 767
rect 5333 713 5347 727
rect 5393 773 5407 787
rect 5412 713 5426 727
rect 5433 713 5447 727
rect 5393 693 5407 707
rect 5273 633 5287 647
rect 5373 633 5387 647
rect 5253 593 5267 607
rect 5373 593 5387 607
rect 5233 453 5247 467
rect 5233 413 5247 427
rect 5293 553 5307 567
rect 5253 394 5267 408
rect 5193 352 5207 366
rect 5233 352 5247 366
rect 5273 353 5287 367
rect 5173 313 5187 327
rect 5153 193 5167 207
rect 5313 433 5327 447
rect 5313 393 5327 407
rect 5353 394 5367 408
rect 5393 394 5407 408
rect 5493 914 5507 928
rect 5533 914 5547 928
rect 5573 933 5587 947
rect 5633 1033 5647 1047
rect 5613 1013 5627 1027
rect 5593 913 5607 927
rect 5493 773 5507 787
rect 5593 873 5607 887
rect 5593 833 5607 847
rect 5513 753 5527 767
rect 5493 713 5507 727
rect 5473 694 5487 708
rect 5513 694 5527 708
rect 5553 793 5567 807
rect 5753 1392 5767 1406
rect 5793 1392 5807 1406
rect 5713 1293 5727 1307
rect 5753 1293 5767 1307
rect 5733 1253 5747 1267
rect 5813 1273 5827 1287
rect 5753 1233 5767 1247
rect 5673 1193 5687 1207
rect 5793 1113 5807 1127
rect 5673 1053 5687 1067
rect 5653 973 5667 987
rect 5753 973 5767 987
rect 5673 953 5687 967
rect 5713 953 5727 967
rect 5633 913 5647 927
rect 5653 872 5667 886
rect 5673 833 5687 847
rect 5633 793 5647 807
rect 5573 773 5587 787
rect 5613 773 5627 787
rect 5593 713 5607 727
rect 5693 793 5707 807
rect 5433 653 5447 667
rect 5473 633 5487 647
rect 5453 613 5467 627
rect 5533 613 5547 627
rect 5493 593 5507 607
rect 5633 694 5647 708
rect 5573 613 5587 627
rect 5553 433 5567 447
rect 5313 353 5327 367
rect 5293 333 5307 347
rect 5333 333 5347 347
rect 5413 353 5427 367
rect 5373 253 5387 267
rect 5413 233 5427 247
rect 5313 192 5327 206
rect 5213 173 5227 187
rect 5273 174 5287 188
rect 5153 132 5167 146
rect 5513 394 5527 408
rect 5453 353 5467 367
rect 5493 313 5507 327
rect 5453 273 5467 287
rect 5513 253 5527 267
rect 5473 213 5487 227
rect 5393 174 5407 188
rect 5433 174 5447 188
rect 5673 653 5687 667
rect 5653 633 5667 647
rect 5613 453 5627 467
rect 5633 453 5647 467
rect 5653 413 5667 427
rect 5733 652 5747 666
rect 5793 653 5807 667
rect 5693 613 5707 627
rect 5713 573 5727 587
rect 5673 394 5687 408
rect 5613 352 5627 366
rect 5653 352 5667 366
rect 5573 313 5587 327
rect 5593 293 5607 307
rect 5573 273 5587 287
rect 5533 233 5547 247
rect 5553 173 5567 187
rect 5593 193 5607 207
rect 5673 333 5687 347
rect 5693 233 5707 247
rect 5673 193 5687 207
rect 5833 1133 5847 1147
rect 5753 413 5767 427
rect 5813 413 5827 427
rect 5773 313 5787 327
rect 5833 313 5847 327
rect 5713 193 5727 207
rect 5773 193 5787 207
rect 5253 132 5267 146
rect 5313 133 5327 147
rect 5373 132 5387 146
rect 5533 132 5547 146
rect 5633 132 5647 146
rect 5673 132 5687 146
rect 5713 133 5727 147
rect 5753 132 5767 146
rect 5033 93 5047 107
rect 5073 93 5087 107
rect 5213 93 5227 107
rect 4913 33 4927 47
rect 3973 13 3987 27
rect 4493 13 4507 27
<< metal3 >>
rect 2047 5476 2093 5484
rect 2187 5476 2213 5484
rect 2667 5476 2833 5484
rect 3267 5476 3293 5484
rect 3047 5456 3233 5464
rect 2647 5436 2733 5444
rect 2887 5436 3013 5444
rect 1387 5416 1453 5424
rect 1867 5416 2093 5424
rect 2107 5416 2573 5424
rect 2627 5416 2713 5424
rect 2827 5416 3133 5424
rect 3227 5416 3773 5424
rect 3847 5416 3973 5424
rect 5467 5416 5693 5424
rect 667 5396 753 5404
rect 2607 5396 2633 5404
rect 2807 5396 3193 5404
rect 4327 5396 4473 5404
rect 347 5376 373 5384
rect 627 5377 693 5385
rect 716 5376 813 5384
rect 216 5364 224 5374
rect 216 5356 273 5364
rect 376 5347 384 5374
rect 367 5336 384 5347
rect 367 5333 380 5336
rect 507 5336 613 5344
rect 716 5346 724 5376
rect 1327 5376 1413 5384
rect 1427 5376 1444 5384
rect 1436 5364 1444 5376
rect 1487 5377 1513 5385
rect 1627 5376 1673 5384
rect 1807 5376 1933 5384
rect 1947 5376 2013 5384
rect 2167 5376 2193 5384
rect 2216 5376 2453 5384
rect 1436 5356 1733 5364
rect 2216 5364 2224 5376
rect 2467 5376 2553 5384
rect 2576 5376 2693 5384
rect 2576 5364 2584 5376
rect 3107 5377 3133 5385
rect 3313 5384 3327 5393
rect 3207 5376 3304 5384
rect 3313 5380 3353 5384
rect 3316 5376 3353 5380
rect 2076 5356 2224 5364
rect 2336 5356 2584 5364
rect 2756 5356 3153 5364
rect 1047 5336 1073 5344
rect 1207 5336 1373 5344
rect 1447 5336 1533 5344
rect 1587 5335 1613 5343
rect 1827 5335 1853 5343
rect 1987 5336 2053 5344
rect 327 5316 673 5324
rect 967 5316 1133 5324
rect 2076 5324 2084 5356
rect 2336 5346 2344 5356
rect 2756 5346 2764 5356
rect 3296 5364 3304 5376
rect 3427 5376 3733 5384
rect 3787 5377 3893 5385
rect 4207 5376 4233 5384
rect 4687 5377 4733 5385
rect 4787 5376 4873 5384
rect 4927 5377 4973 5385
rect 4987 5376 5053 5384
rect 5147 5377 5173 5385
rect 5196 5376 5213 5384
rect 3296 5356 3344 5364
rect 2187 5336 2233 5344
rect 2587 5336 2713 5344
rect 2887 5336 3013 5344
rect 3336 5346 3344 5356
rect 3967 5356 4453 5364
rect 3387 5335 3413 5343
rect 3607 5335 3653 5343
rect 4176 5346 4184 5356
rect 5196 5364 5204 5376
rect 5527 5377 5553 5385
rect 5607 5377 5633 5385
rect 5036 5356 5204 5364
rect 3787 5336 3813 5344
rect 4327 5335 4353 5343
rect 5036 5346 5044 5356
rect 4487 5336 4753 5344
rect 4947 5336 5033 5344
rect 5247 5336 5313 5344
rect 5387 5336 5573 5344
rect 5647 5335 5673 5343
rect 1847 5316 2084 5324
rect 3127 5316 3213 5324
rect 3727 5316 4073 5324
rect 4087 5316 4413 5324
rect 1747 5296 1773 5304
rect 1787 5296 2113 5304
rect 2507 5296 2633 5304
rect 2687 5296 3033 5304
rect 3747 5296 3953 5304
rect 4467 5296 4713 5304
rect 687 5276 713 5284
rect 767 5276 793 5284
rect 807 5276 1473 5284
rect 1807 5276 1833 5284
rect 2047 5276 2073 5284
rect 3827 5276 3993 5284
rect 4807 5276 5093 5284
rect 1147 5260 1304 5264
rect 1147 5256 1307 5260
rect 1293 5247 1307 5256
rect 2667 5256 2853 5264
rect 2967 5256 2993 5264
rect 47 5236 553 5244
rect 567 5236 593 5244
rect 607 5236 693 5244
rect 707 5236 953 5244
rect 1487 5236 1653 5244
rect 1667 5236 1793 5244
rect 3167 5236 4273 5244
rect 4287 5236 4613 5244
rect 4867 5236 5133 5244
rect 1047 5216 2193 5224
rect 3507 5216 3553 5224
rect 1307 5196 2053 5204
rect 2067 5196 2273 5204
rect 2707 5196 2813 5204
rect 2927 5196 3433 5204
rect 3447 5196 3713 5204
rect 3727 5196 3773 5204
rect 3867 5196 4673 5204
rect 4687 5196 4893 5204
rect 87 5176 113 5184
rect 1087 5176 1113 5184
rect 1227 5176 2593 5184
rect 3267 5176 3513 5184
rect 5167 5176 5373 5184
rect 2827 5156 4013 5164
rect 4827 5156 4913 5164
rect 4927 5156 5473 5164
rect 287 5136 973 5144
rect 1147 5136 1253 5144
rect 1427 5136 1753 5144
rect 1767 5136 1993 5144
rect 2447 5136 2753 5144
rect 2947 5136 2973 5144
rect 3027 5136 3293 5144
rect 4127 5136 4513 5144
rect 4627 5136 4753 5144
rect 4847 5136 5193 5144
rect 1007 5116 1173 5124
rect 1187 5116 1393 5124
rect 1547 5116 1613 5124
rect 2027 5116 2353 5124
rect 2407 5116 2993 5124
rect 3087 5116 3173 5124
rect 3847 5116 3973 5124
rect 4567 5116 4813 5124
rect 5467 5116 5513 5124
rect 5527 5116 5713 5124
rect 5727 5116 5753 5124
rect 567 5096 813 5104
rect 2007 5096 2373 5104
rect 4247 5096 4293 5104
rect 5027 5096 5113 5104
rect 67 5077 113 5085
rect 167 5077 193 5085
rect 236 5047 244 5074
rect 327 5076 393 5084
rect 467 5077 513 5085
rect 776 5076 873 5084
rect 76 5040 133 5044
rect 73 5036 133 5040
rect 73 5027 87 5036
rect 227 5036 244 5047
rect 227 5033 240 5036
rect 347 5036 373 5044
rect 656 5044 664 5074
rect 776 5046 784 5076
rect 1087 5077 1133 5085
rect 1367 5077 1513 5085
rect 1587 5077 1652 5085
rect 1687 5077 1713 5085
rect 1736 5076 1853 5084
rect 973 5064 987 5073
rect 1736 5064 1744 5076
rect 1936 5076 1973 5084
rect 1936 5067 1944 5076
rect 2307 5077 2333 5085
rect 2507 5076 2553 5084
rect 1920 5066 1944 5067
rect 973 5060 1024 5064
rect 976 5056 1024 5060
rect 547 5036 664 5044
rect 787 5036 933 5044
rect 1016 5046 1024 5056
rect 1636 5056 1744 5064
rect 1427 5035 1473 5043
rect 1636 5046 1644 5056
rect 1927 5056 1944 5066
rect 1927 5053 1940 5056
rect 1527 5036 1593 5044
rect 1707 5036 1733 5044
rect 2127 5036 2213 5044
rect 2236 5044 2244 5074
rect 2647 5077 2673 5085
rect 2793 5064 2807 5073
rect 2596 5060 2807 5064
rect 2596 5056 2804 5060
rect 2236 5036 2353 5044
rect 2407 5036 2513 5044
rect 2596 5044 2604 5056
rect 2527 5036 2604 5044
rect 2627 5035 2693 5043
rect 2787 5035 2813 5043
rect 2956 5044 2964 5073
rect 2956 5036 3013 5044
rect 3036 5044 3044 5074
rect 3156 5047 3164 5074
rect 3187 5084 3200 5087
rect 3187 5073 3204 5084
rect 3387 5076 3433 5084
rect 3687 5077 3713 5085
rect 3887 5077 3933 5085
rect 4027 5076 4064 5084
rect 3036 5036 3133 5044
rect 3156 5036 3172 5047
rect 3160 5033 3172 5036
rect 3196 5046 3204 5073
rect 3407 5036 3793 5044
rect 3816 5044 3824 5073
rect 3816 5036 3853 5044
rect 3976 5044 3984 5074
rect 4056 5046 4064 5076
rect 4147 5077 4173 5085
rect 3927 5036 3984 5044
rect 827 5016 893 5024
rect 1007 5016 1053 5024
rect 1147 5016 1213 5024
rect 1667 5016 1833 5024
rect 2887 5016 2933 5024
rect 4007 5016 4033 5024
rect 4336 5024 4344 5074
rect 4087 5016 4344 5024
rect 207 4996 253 5004
rect 707 4996 793 5004
rect 1127 4996 1273 5004
rect 1427 4996 1673 5004
rect 2267 4996 2433 5004
rect 2487 4996 2653 5004
rect 2747 4996 2793 5004
rect 3307 4996 3613 5004
rect 3667 4996 3753 5004
rect 3947 4996 4053 5004
rect 4147 4996 4353 5004
rect 4376 5004 4384 5074
rect 4447 5076 4493 5084
rect 4667 5077 4713 5085
rect 4827 5076 4853 5084
rect 4936 5076 4953 5084
rect 4936 5047 4944 5076
rect 5127 5076 5213 5084
rect 5076 5064 5084 5074
rect 5287 5076 5333 5084
rect 5407 5077 5493 5085
rect 5607 5076 5653 5084
rect 5076 5060 5184 5064
rect 5076 5056 5187 5060
rect 5173 5047 5187 5056
rect 4587 5036 4673 5044
rect 4787 5035 4813 5043
rect 4887 5035 4912 5043
rect 4987 5035 5013 5043
rect 5107 5035 5152 5043
rect 5247 5035 5273 5043
rect 5536 5024 5544 5074
rect 5507 5016 5544 5024
rect 4376 4996 4733 5004
rect 4927 4996 5433 5004
rect 5487 4996 5653 5004
rect 427 4976 653 4984
rect 667 4976 853 4984
rect 947 4976 1233 4984
rect 3207 4976 3253 4984
rect 5247 4976 5273 4984
rect 5287 4976 5353 4984
rect 727 4956 753 4964
rect 987 4956 1193 4964
rect 1447 4956 1653 4964
rect 2527 4956 2633 4964
rect 2767 4956 3073 4964
rect 3627 4956 3733 4964
rect 4527 4956 5053 4964
rect 5407 4956 5473 4964
rect 107 4936 213 4944
rect 227 4936 493 4944
rect 507 4936 953 4944
rect 967 4936 1413 4944
rect 1687 4936 2973 4944
rect 3247 4936 3273 4944
rect 3767 4936 4073 4944
rect 4667 4936 4913 4944
rect 727 4916 1133 4924
rect 1947 4916 2032 4924
rect 2067 4916 2093 4924
rect 2207 4916 2233 4924
rect 2247 4916 2473 4924
rect 3147 4916 3213 4924
rect 4487 4916 4553 4924
rect 4567 4916 4593 4924
rect 5007 4916 5313 4924
rect 5727 4916 5833 4924
rect 247 4896 273 4904
rect 287 4896 313 4904
rect 1167 4896 1293 4904
rect 1347 4896 1493 4904
rect 1607 4896 1673 4904
rect 1687 4896 1844 4904
rect 1836 4887 1844 4896
rect 2347 4896 2413 4904
rect 2707 4896 2893 4904
rect 2967 4896 3073 4904
rect 3127 4896 3253 4904
rect 3547 4896 3733 4904
rect 4627 4896 4693 4904
rect 4787 4896 4933 4904
rect 5067 4896 5133 4904
rect 5567 4896 5693 4904
rect 587 4876 753 4884
rect 847 4876 893 4884
rect 907 4876 1113 4884
rect 1847 4876 1913 4884
rect 2567 4876 2593 4884
rect 3307 4876 3333 4884
rect 3567 4876 3592 4884
rect 3787 4876 3893 4884
rect 4467 4876 4573 4884
rect 4747 4876 4813 4884
rect 107 4856 153 4864
rect 207 4856 313 4864
rect 367 4856 413 4864
rect 56 4827 64 4853
rect 316 4844 324 4854
rect 1227 4857 1253 4865
rect 1727 4856 1773 4864
rect 316 4836 484 4844
rect 287 4815 333 4823
rect 427 4815 453 4823
rect 476 4824 484 4836
rect 476 4816 593 4824
rect 616 4824 624 4854
rect 616 4816 733 4824
rect 747 4816 833 4824
rect 1207 4816 1313 4824
rect 1436 4824 1444 4854
rect 2387 4857 2473 4865
rect 2496 4856 2533 4864
rect 1920 4844 1933 4847
rect 1916 4833 1933 4844
rect 1436 4816 1473 4824
rect 1916 4824 1924 4833
rect 1747 4816 1924 4824
rect 2247 4815 2273 4823
rect 2296 4824 2304 4854
rect 2496 4844 2504 4856
rect 2736 4856 2833 4864
rect 2436 4836 2504 4844
rect 2436 4826 2444 4836
rect 2736 4826 2744 4856
rect 2927 4856 3013 4864
rect 3067 4856 3093 4864
rect 3116 4856 3133 4864
rect 2296 4816 2364 4824
rect 1467 4796 1573 4804
rect 1587 4796 1693 4804
rect 1787 4796 1933 4804
rect 2356 4804 2364 4816
rect 2907 4815 2953 4823
rect 3116 4824 3124 4856
rect 3267 4856 3404 4864
rect 3176 4827 3184 4853
rect 3396 4844 3404 4856
rect 3613 4864 3627 4873
rect 3447 4856 3464 4864
rect 3613 4860 3653 4864
rect 3616 4856 3653 4860
rect 3396 4836 3424 4844
rect 3047 4816 3124 4824
rect 3416 4826 3424 4836
rect 3227 4816 3273 4824
rect 2356 4796 2633 4804
rect 2867 4796 2993 4804
rect 3127 4796 3153 4804
rect 3456 4804 3464 4856
rect 3807 4856 3833 4864
rect 3696 4844 3704 4854
rect 4167 4856 4353 4864
rect 3487 4836 3704 4844
rect 4396 4844 4404 4854
rect 4947 4856 5093 4864
rect 5107 4856 5344 4864
rect 3907 4836 4024 4844
rect 4396 4836 4664 4844
rect 3647 4816 3753 4824
rect 4016 4826 4024 4836
rect 4656 4827 4664 4836
rect 4267 4816 4293 4824
rect 4656 4816 4672 4827
rect 4660 4813 4672 4816
rect 4707 4816 4873 4824
rect 5127 4816 5173 4824
rect 5336 4826 5344 4856
rect 5713 4864 5727 4872
rect 5687 4860 5727 4864
rect 5687 4856 5724 4860
rect 5387 4816 5493 4824
rect 5627 4816 5793 4824
rect 3456 4796 3513 4804
rect 3827 4796 3953 4804
rect 4387 4796 4493 4804
rect 4647 4796 4933 4804
rect 167 4776 493 4784
rect 507 4776 693 4784
rect 1013 4784 1027 4793
rect 1013 4780 1113 4784
rect 1016 4776 1113 4780
rect 2187 4776 2333 4784
rect 2567 4776 2733 4784
rect 3047 4776 3673 4784
rect 3687 4776 4153 4784
rect 4687 4776 4753 4784
rect 5027 4776 5053 4784
rect 5067 4776 5213 4784
rect 807 4756 1073 4764
rect 1407 4756 1633 4764
rect 1707 4756 1913 4764
rect 1927 4756 2073 4764
rect 2147 4756 2253 4764
rect 2667 4756 2793 4764
rect 4427 4756 4553 4764
rect 2467 4736 2973 4744
rect 2987 4736 3173 4744
rect 3187 4736 3393 4744
rect 3407 4736 3913 4744
rect 3987 4736 4073 4744
rect 4087 4736 4133 4744
rect 4307 4736 4633 4744
rect 4647 4736 4813 4744
rect 4827 4736 5153 4744
rect 5167 4736 5373 4744
rect 667 4716 893 4724
rect 1267 4716 1353 4724
rect 1367 4716 1393 4724
rect 1527 4716 1793 4724
rect 2487 4716 2513 4724
rect 2527 4716 2773 4724
rect 3227 4716 3253 4724
rect 4467 4716 4493 4724
rect 5407 4716 5453 4724
rect 2067 4696 2833 4704
rect 3107 4696 3473 4704
rect 3787 4696 3833 4704
rect 4887 4696 4913 4704
rect 5487 4696 5513 4704
rect 1487 4676 1713 4684
rect 2667 4676 2893 4684
rect 3327 4676 3693 4684
rect 5147 4676 5693 4684
rect 707 4656 1013 4664
rect 2507 4656 2593 4664
rect 2607 4656 2953 4664
rect 3607 4656 3673 4664
rect 3807 4656 4473 4664
rect 747 4636 953 4644
rect 2107 4636 2133 4644
rect 2707 4636 2813 4644
rect 3287 4636 3453 4644
rect 3547 4636 3733 4644
rect 4527 4636 4853 4644
rect 2847 4616 3593 4624
rect 3967 4616 4293 4624
rect 4467 4616 4573 4624
rect 127 4596 373 4604
rect 387 4596 433 4604
rect 1007 4596 1093 4604
rect 2027 4596 2093 4604
rect 2387 4596 2653 4604
rect 2667 4596 2713 4604
rect 2907 4596 3424 4604
rect 1247 4576 1273 4584
rect 1427 4576 1833 4584
rect 1847 4576 1993 4584
rect 2747 4576 2833 4584
rect 3007 4576 3033 4584
rect 3156 4576 3193 4584
rect 87 4556 153 4564
rect 167 4556 213 4564
rect 287 4557 313 4565
rect 367 4557 393 4565
rect 527 4557 573 4565
rect 627 4557 653 4565
rect 747 4556 764 4564
rect 476 4544 484 4554
rect 436 4536 484 4544
rect 107 4515 153 4523
rect 247 4516 273 4524
rect 436 4524 444 4536
rect 756 4527 764 4556
rect 1027 4557 1053 4565
rect 1467 4556 1564 4564
rect 347 4516 444 4524
rect 467 4516 513 4524
rect 836 4524 844 4554
rect 1556 4526 1564 4556
rect 1587 4556 1613 4564
rect 1767 4564 1780 4567
rect 1767 4553 1784 4564
rect 1807 4556 1933 4564
rect 1956 4556 2053 4564
rect 1616 4540 1733 4544
rect 1613 4536 1733 4540
rect 1613 4527 1627 4536
rect 816 4516 844 4524
rect 816 4504 824 4516
rect 967 4515 993 4523
rect 1427 4515 1473 4523
rect 1776 4526 1784 4553
rect 1956 4526 1964 4556
rect 2207 4557 2233 4565
rect 2007 4516 2073 4524
rect 2327 4515 2353 4523
rect 2536 4524 2544 4554
rect 3107 4557 3133 4565
rect 2676 4527 2684 4553
rect 2447 4516 2544 4524
rect 2667 4516 2684 4527
rect 3156 4526 3164 4576
rect 3416 4584 3424 4596
rect 3447 4596 3653 4604
rect 3787 4596 3824 4604
rect 3416 4576 3584 4584
rect 3336 4556 3353 4564
rect 3336 4527 3344 4556
rect 3576 4564 3584 4576
rect 3607 4584 3620 4587
rect 3816 4584 3824 4596
rect 4427 4596 4464 4604
rect 3607 4573 3624 4584
rect 3816 4576 3873 4584
rect 4027 4576 4104 4584
rect 3616 4564 3624 4573
rect 3407 4556 3564 4564
rect 3576 4556 3604 4564
rect 3616 4556 3793 4564
rect 2667 4513 2680 4516
rect 2747 4516 2853 4524
rect 2867 4515 3053 4523
rect 3227 4516 3253 4524
rect 3556 4526 3564 4556
rect 3596 4544 3604 4556
rect 3933 4564 3947 4573
rect 3907 4560 3947 4564
rect 3907 4556 3944 4560
rect 4096 4564 4104 4576
rect 4096 4556 4113 4564
rect 4367 4557 4393 4565
rect 4416 4556 4433 4564
rect 3596 4536 3644 4544
rect 3387 4520 3424 4524
rect 3387 4516 3427 4520
rect 3413 4507 3427 4516
rect 607 4496 824 4504
rect 1147 4496 1333 4504
rect 2216 4496 2373 4504
rect 207 4476 393 4484
rect 1547 4476 1693 4484
rect 2216 4484 2224 4496
rect 3636 4504 3644 4536
rect 3667 4516 3913 4524
rect 3927 4515 3953 4523
rect 3976 4506 3984 4553
rect 4056 4527 4064 4553
rect 4416 4544 4424 4556
rect 4216 4536 4424 4544
rect 4456 4544 4464 4596
rect 4607 4596 4893 4604
rect 4947 4596 5033 4604
rect 5047 4596 5573 4604
rect 5627 4596 5693 4604
rect 4616 4556 4693 4564
rect 4456 4536 4564 4544
rect 4216 4526 4224 4536
rect 4427 4516 4533 4524
rect 4556 4524 4564 4536
rect 4616 4527 4624 4556
rect 4767 4556 4813 4564
rect 4867 4556 4973 4564
rect 4987 4556 5093 4564
rect 5227 4557 5253 4565
rect 5396 4556 5453 4564
rect 5133 4544 5147 4553
rect 5396 4547 5404 4556
rect 4996 4540 5147 4544
rect 4993 4536 5144 4540
rect 4993 4527 5007 4536
rect 5387 4536 5404 4547
rect 5656 4544 5664 4554
rect 5556 4536 5664 4544
rect 5387 4533 5400 4536
rect 4556 4516 4573 4524
rect 4727 4515 4753 4523
rect 5047 4515 5113 4523
rect 5287 4515 5333 4523
rect 5556 4524 5564 4536
rect 5716 4527 5724 4553
rect 5447 4516 5564 4524
rect 3636 4496 3864 4504
rect 3856 4487 3864 4496
rect 4687 4496 4953 4504
rect 1947 4476 2224 4484
rect 2247 4476 2353 4484
rect 2427 4476 2553 4484
rect 2607 4476 2693 4484
rect 3327 4476 3513 4484
rect 3856 4476 3873 4487
rect 3860 4473 3873 4476
rect 4027 4476 4073 4484
rect 4327 4476 4353 4484
rect 4367 4476 4573 4484
rect 5227 4476 5433 4484
rect 5567 4476 5673 4484
rect 667 4456 1073 4464
rect 1167 4456 1193 4464
rect 1207 4456 1473 4464
rect 1487 4456 1513 4464
rect 2607 4456 2633 4464
rect 2847 4456 3333 4464
rect 3347 4456 3593 4464
rect 4387 4456 4472 4464
rect 4507 4456 4593 4464
rect 4887 4456 4973 4464
rect 5487 4456 5573 4464
rect 5587 4456 5613 4464
rect 287 4436 373 4444
rect 1287 4436 1373 4444
rect 1387 4436 1553 4444
rect 2447 4436 2653 4444
rect 2667 4436 3033 4444
rect 3047 4436 3113 4444
rect 3127 4436 3733 4444
rect 3947 4436 4013 4444
rect 4027 4436 4093 4444
rect 5207 4436 5253 4444
rect 5527 4436 5553 4444
rect 5687 4436 5793 4444
rect 567 4416 953 4424
rect 3067 4416 3433 4424
rect 3556 4416 3653 4424
rect 407 4396 493 4404
rect 1407 4396 1593 4404
rect 2347 4396 2533 4404
rect 2667 4396 2813 4404
rect 2967 4396 3233 4404
rect 3247 4396 3293 4404
rect 3556 4404 3564 4416
rect 4047 4416 4673 4424
rect 4847 4416 5033 4424
rect 5107 4416 5373 4424
rect 5447 4416 5653 4424
rect 3307 4396 3564 4404
rect 3887 4396 3913 4404
rect 3967 4396 4104 4404
rect 67 4376 313 4384
rect 567 4376 613 4384
rect 1187 4376 1393 4384
rect 2147 4376 2253 4384
rect 2307 4376 3973 4384
rect 4096 4384 4104 4396
rect 4127 4396 4493 4404
rect 4096 4376 4204 4384
rect 487 4356 633 4364
rect 647 4356 693 4364
rect 927 4356 973 4364
rect 987 4356 1093 4364
rect 1307 4356 1493 4364
rect 1927 4356 2013 4364
rect 2027 4356 2073 4364
rect 2947 4356 2973 4364
rect 3607 4356 3673 4364
rect 3796 4356 3833 4364
rect 107 4336 253 4344
rect 456 4336 593 4344
rect 87 4296 193 4304
rect 267 4295 293 4303
rect 416 4304 424 4334
rect 367 4296 424 4304
rect 456 4304 464 4336
rect 656 4336 713 4344
rect 656 4324 664 4336
rect 1047 4336 1313 4344
rect 2327 4337 2393 4345
rect 2447 4336 2524 4344
rect 536 4316 664 4324
rect 536 4306 544 4316
rect 447 4296 464 4304
rect 987 4295 1013 4303
rect 1187 4296 1213 4304
rect 1436 4304 1444 4334
rect 1307 4296 1513 4304
rect 2207 4296 2312 4304
rect 2516 4306 2524 4336
rect 2747 4337 2793 4345
rect 3347 4336 3424 4344
rect 2696 4307 2704 4334
rect 2347 4295 2373 4303
rect 2696 4296 2713 4307
rect 2700 4293 2713 4296
rect 3416 4304 3424 4336
rect 3616 4336 3693 4344
rect 3556 4324 3564 4334
rect 3616 4327 3624 4336
rect 3747 4337 3773 4345
rect 3556 4316 3613 4324
rect 3796 4306 3804 4356
rect 4100 4364 4113 4367
rect 4096 4353 4113 4364
rect 4196 4364 4204 4376
rect 4687 4376 4833 4384
rect 5447 4376 5672 4384
rect 5693 4384 5707 4393
rect 5693 4380 5753 4384
rect 5696 4376 5753 4380
rect 4196 4356 4224 4364
rect 4096 4344 4104 4353
rect 3907 4336 4104 4344
rect 3416 4296 3433 4304
rect 3887 4295 3973 4303
rect 4136 4304 4144 4334
rect 4107 4296 4144 4304
rect 4216 4304 4224 4356
rect 4807 4336 4833 4344
rect 4856 4336 4873 4344
rect 4856 4324 4864 4336
rect 4953 4344 4967 4353
rect 4936 4340 4967 4344
rect 4936 4336 4964 4340
rect 4936 4324 4944 4336
rect 5173 4344 5187 4353
rect 5147 4340 5187 4344
rect 5147 4336 5184 4340
rect 5267 4336 5313 4344
rect 4796 4316 4864 4324
rect 4896 4316 4944 4324
rect 4216 4296 4253 4304
rect 4507 4295 4613 4303
rect 4796 4304 4804 4316
rect 4896 4306 4904 4316
rect 4787 4296 4804 4304
rect 4967 4296 5013 4304
rect 5216 4304 5224 4333
rect 5167 4296 5224 4304
rect 5356 4304 5364 4334
rect 5356 4296 5453 4304
rect 5556 4304 5564 4333
rect 5556 4296 5673 4304
rect 5796 4304 5804 4334
rect 5836 4307 5844 4333
rect 5747 4296 5804 4304
rect 1607 4276 1893 4284
rect 2747 4276 2793 4284
rect 2887 4276 2973 4284
rect 2987 4276 3373 4284
rect 3967 4276 4053 4284
rect 4327 4276 4493 4284
rect 4507 4276 4693 4284
rect 5367 4276 5413 4284
rect 5587 4276 5813 4284
rect 667 4256 833 4264
rect 967 4256 993 4264
rect 1007 4256 1053 4264
rect 1067 4256 1293 4264
rect 1487 4256 1513 4264
rect 1987 4256 2633 4264
rect 3947 4256 3993 4264
rect 4107 4256 4413 4264
rect 5327 4256 5393 4264
rect 5533 4264 5547 4273
rect 5447 4260 5547 4264
rect 5447 4256 5544 4260
rect 5747 4256 5773 4264
rect 1587 4236 2413 4244
rect 2427 4236 2993 4244
rect 3287 4236 3333 4244
rect 3347 4236 3593 4244
rect 4047 4236 4373 4244
rect 1387 4216 1413 4224
rect 1747 4216 1773 4224
rect 1787 4216 1873 4224
rect 2047 4216 2393 4224
rect 2727 4216 2813 4224
rect 4467 4216 4973 4224
rect 4987 4216 5353 4224
rect 587 4196 653 4204
rect 1647 4196 2013 4204
rect 2707 4196 2913 4204
rect 3007 4196 3313 4204
rect 3327 4196 3593 4204
rect 3667 4196 3913 4204
rect 3927 4196 4124 4204
rect 1656 4176 1753 4184
rect 387 4156 413 4164
rect 1656 4164 1664 4176
rect 2247 4176 2673 4184
rect 3107 4176 3193 4184
rect 3207 4176 3373 4184
rect 3627 4176 3993 4184
rect 4116 4184 4124 4196
rect 4116 4176 4593 4184
rect 4607 4176 5113 4184
rect 5127 4176 5173 4184
rect 1507 4156 1664 4164
rect 1707 4156 2573 4164
rect 2587 4156 3573 4164
rect 3587 4156 4013 4164
rect 4647 4156 4773 4164
rect 2767 4136 3173 4144
rect 3307 4136 3673 4144
rect 3867 4136 3973 4144
rect 4227 4136 4313 4144
rect 4707 4136 5473 4144
rect 127 4116 373 4124
rect 927 4116 1113 4124
rect 1127 4116 1273 4124
rect 1287 4116 1453 4124
rect 1467 4116 1653 4124
rect 1667 4116 2233 4124
rect 4067 4116 4153 4124
rect 4507 4116 5253 4124
rect 2287 4096 2473 4104
rect 2967 4096 3193 4104
rect 3267 4096 3413 4104
rect 4007 4096 4473 4104
rect 4587 4096 4793 4104
rect 5287 4096 5753 4104
rect 487 4076 673 4084
rect 1247 4076 1573 4084
rect 1767 4076 2293 4084
rect 2767 4076 2893 4084
rect 3487 4076 3553 4084
rect 3567 4076 3713 4084
rect 3987 4076 4293 4084
rect 4307 4076 4353 4084
rect 4527 4076 4993 4084
rect 1360 4064 1373 4067
rect 1356 4053 1373 4064
rect 2967 4056 3133 4064
rect 3247 4056 3453 4064
rect 3547 4056 3733 4064
rect 3787 4056 3893 4064
rect 4447 4056 4493 4064
rect 5136 4056 5173 4064
rect 167 4036 193 4044
rect 207 4036 233 4044
rect 587 4036 713 4044
rect 787 4036 804 4044
rect 276 4024 284 4034
rect 796 4024 804 4036
rect 827 4037 853 4045
rect 1036 4036 1053 4044
rect 896 4024 904 4034
rect 276 4016 384 4024
rect 796 4016 1013 4024
rect 207 3995 353 4003
rect 376 4004 384 4016
rect 1036 4007 1044 4036
rect 1356 4047 1364 4053
rect 1347 4036 1364 4047
rect 1347 4033 1360 4036
rect 1407 4036 1604 4044
rect 376 3996 433 4004
rect 1596 4006 1604 4036
rect 1727 4037 1753 4045
rect 1907 4037 1933 4045
rect 2593 4044 2607 4053
rect 2367 4040 2607 4044
rect 2367 4036 2604 4040
rect 1527 3996 1553 4004
rect 1616 4004 1624 4034
rect 2016 4007 2024 4034
rect 1616 3996 1853 4004
rect 2016 3996 2033 4007
rect 2020 3993 2033 3996
rect 267 3976 313 3984
rect 767 3976 813 3984
rect 827 3976 933 3984
rect 2176 3984 2184 4034
rect 2476 4024 2484 4036
rect 2687 4036 2773 4044
rect 2796 4036 2953 4044
rect 2796 4024 2804 4036
rect 3007 4037 3053 4045
rect 3300 4044 3313 4047
rect 3296 4033 3313 4044
rect 4407 4036 4513 4044
rect 4567 4037 4593 4045
rect 4616 4036 4753 4044
rect 2476 4016 2804 4024
rect 2287 3995 2453 4003
rect 2807 3996 2853 4004
rect 2927 3996 2973 4004
rect 3027 3996 3113 4004
rect 3176 4004 3184 4033
rect 3127 3996 3184 4004
rect 3207 3996 3273 4004
rect 3296 3987 3304 4033
rect 3356 4004 3364 4033
rect 3356 3996 3393 4004
rect 3467 3995 3753 4003
rect 3856 4004 3864 4033
rect 3807 3996 3864 4004
rect 3976 4004 3984 4033
rect 4036 4024 4044 4034
rect 4076 4024 4084 4034
rect 4036 4020 4064 4024
rect 4036 4016 4067 4020
rect 4076 4016 4193 4024
rect 3927 3996 3984 4004
rect 4053 4007 4067 4016
rect 4267 3995 4293 4003
rect 4387 3996 4433 4004
rect 2176 3976 2233 3984
rect 2467 3976 2593 3984
rect 3767 3976 3873 3984
rect 4516 3984 4524 4034
rect 4616 4006 4624 4036
rect 5047 4037 5073 4045
rect 5136 4006 5144 4056
rect 5296 4056 5533 4064
rect 5296 4006 5304 4056
rect 5327 4037 5393 4045
rect 5416 4036 5453 4044
rect 4827 3995 4873 4003
rect 4947 3995 4973 4003
rect 4516 3976 4593 3984
rect 4607 3976 4653 3984
rect 5127 3976 5333 3984
rect 5416 3984 5424 4036
rect 5747 4036 5804 4044
rect 5553 4024 5567 4033
rect 5436 4020 5644 4024
rect 5436 4016 5647 4020
rect 5436 4006 5444 4016
rect 5633 4007 5647 4016
rect 5676 4007 5684 4033
rect 5796 4007 5804 4036
rect 5387 3976 5424 3984
rect 5547 3976 5573 3984
rect 5667 3976 5753 3984
rect 147 3956 313 3964
rect 1027 3956 1213 3964
rect 1227 3956 1273 3964
rect 2007 3956 2053 3964
rect 2067 3956 2313 3964
rect 3167 3956 3473 3964
rect 3487 3956 3953 3964
rect 4507 3956 4553 3964
rect 4807 3956 5013 3964
rect 3247 3936 3333 3944
rect 3907 3936 3933 3944
rect 3987 3936 4133 3944
rect 4187 3936 4253 3944
rect 507 3916 573 3924
rect 587 3916 653 3924
rect 667 3916 693 3924
rect 707 3916 733 3924
rect 1227 3916 1333 3924
rect 1767 3916 1813 3924
rect 1907 3916 2333 3924
rect 2347 3916 2433 3924
rect 3387 3916 3493 3924
rect 3507 3916 3733 3924
rect 3967 3916 4233 3924
rect 4867 3916 4913 3924
rect 5247 3916 5353 3924
rect 5607 3916 5673 3924
rect 247 3896 293 3904
rect 307 3896 353 3904
rect 1607 3896 1953 3904
rect 2067 3896 2133 3904
rect 3067 3896 3473 3904
rect 4027 3896 4053 3904
rect 5007 3896 5073 3904
rect 5527 3896 5573 3904
rect 407 3876 493 3884
rect 547 3876 613 3884
rect 627 3876 693 3884
rect 707 3876 873 3884
rect 1307 3876 1413 3884
rect 1627 3876 1773 3884
rect 2387 3876 2893 3884
rect 3027 3876 3093 3884
rect 3107 3876 3373 3884
rect 3847 3876 3913 3884
rect 5267 3876 5433 3884
rect 5727 3876 5773 3884
rect 267 3856 293 3864
rect 727 3856 773 3864
rect 847 3856 993 3864
rect 1007 3856 1053 3864
rect 1287 3856 1593 3864
rect 1847 3856 1973 3864
rect 4087 3856 4324 3864
rect 4316 3847 4324 3856
rect 5187 3856 5233 3864
rect 327 3836 453 3844
rect 616 3836 1153 3844
rect 167 3817 193 3825
rect 476 3816 573 3824
rect 396 3787 404 3813
rect 436 3787 444 3813
rect 127 3776 153 3784
rect 267 3775 293 3783
rect 476 3786 484 3816
rect 616 3824 624 3836
rect 2507 3836 2533 3844
rect 3967 3836 4093 3844
rect 4207 3836 4273 3844
rect 4327 3836 4653 3844
rect 5680 3844 5693 3847
rect 5676 3833 5693 3844
rect 596 3816 624 3824
rect 596 3786 604 3816
rect 687 3816 884 3824
rect 876 3804 884 3816
rect 907 3816 953 3824
rect 1207 3816 1293 3824
rect 1347 3817 1373 3825
rect 1453 3824 1467 3833
rect 1453 3820 1533 3824
rect 1456 3816 1533 3820
rect 1887 3817 1933 3825
rect 2107 3816 2144 3824
rect 1976 3804 1984 3814
rect 876 3796 904 3804
rect 1976 3796 2064 3804
rect 847 3775 873 3783
rect 896 3767 904 3796
rect 967 3775 993 3783
rect 1167 3775 1193 3783
rect 1347 3776 1513 3784
rect 1567 3776 1593 3784
rect 1967 3776 2013 3784
rect 2056 3784 2064 3796
rect 2136 3787 2144 3816
rect 2167 3817 2193 3825
rect 2260 3824 2273 3827
rect 2256 3813 2273 3824
rect 2427 3817 2453 3825
rect 2056 3776 2073 3784
rect 2256 3786 2264 3813
rect 2316 3784 2324 3813
rect 2776 3786 2784 3833
rect 2967 3817 3073 3825
rect 3387 3816 3433 3824
rect 2316 3776 2333 3784
rect 2627 3775 2653 3783
rect 2727 3776 2773 3784
rect 2847 3775 2873 3783
rect 3087 3775 3133 3783
rect 3347 3776 3413 3784
rect 3496 3784 3504 3814
rect 3727 3816 3793 3824
rect 3847 3816 3873 3824
rect 3887 3817 3913 3825
rect 3980 3824 3993 3827
rect 3976 3813 3993 3824
rect 4133 3824 4147 3833
rect 4133 3820 4333 3824
rect 4136 3816 4333 3820
rect 4627 3816 4693 3824
rect 4767 3816 4813 3824
rect 4987 3817 5053 3825
rect 5147 3817 5193 3825
rect 3976 3786 3984 3813
rect 4856 3787 4864 3813
rect 3467 3776 3504 3784
rect 3627 3775 3713 3783
rect 4107 3775 4133 3783
rect 4207 3776 4273 3784
rect 4287 3776 4433 3784
rect 4447 3776 4493 3784
rect 4627 3775 4673 3783
rect 4727 3775 4753 3783
rect 5107 3775 5153 3783
rect 707 3756 793 3764
rect 1927 3756 2053 3764
rect 2407 3756 2493 3764
rect 4307 3756 4333 3764
rect 4687 3756 4793 3764
rect 4847 3756 4973 3764
rect 4987 3756 5073 3764
rect 5316 3764 5324 3814
rect 5427 3817 5473 3825
rect 5376 3784 5384 3813
rect 5676 3787 5684 3833
rect 5376 3776 5453 3784
rect 5316 3756 5393 3764
rect 207 3736 313 3744
rect 387 3736 633 3744
rect 867 3736 913 3744
rect 1947 3736 1993 3744
rect 2127 3736 2153 3744
rect 2167 3736 2373 3744
rect 2387 3736 3413 3744
rect 3427 3736 3873 3744
rect 4127 3736 4213 3744
rect 4587 3736 5113 3744
rect 5167 3736 5333 3744
rect 5447 3736 5513 3744
rect 5716 3744 5724 3814
rect 5747 3775 5793 3783
rect 5716 3736 5793 3744
rect 1587 3716 1873 3724
rect 2307 3716 2333 3724
rect 3467 3716 3673 3724
rect 3687 3716 3813 3724
rect 4107 3716 4233 3724
rect 4507 3716 4873 3724
rect 87 3696 213 3704
rect 547 3696 1033 3704
rect 1527 3696 1533 3704
rect 1547 3696 1733 3704
rect 1847 3696 2133 3704
rect 3387 3696 3773 3704
rect 3847 3696 4253 3704
rect 4647 3696 4953 3704
rect 5087 3696 5573 3704
rect 1227 3676 1253 3684
rect 1907 3676 2073 3684
rect 2427 3676 3093 3684
rect 3827 3676 4192 3684
rect 4227 3676 4313 3684
rect 407 3656 1033 3664
rect 3067 3656 3573 3664
rect 4027 3656 4113 3664
rect 4867 3656 4993 3664
rect 5127 3656 5613 3664
rect 5627 3656 5693 3664
rect 1507 3636 1713 3644
rect 2007 3636 2433 3644
rect 3167 3636 3193 3644
rect 3207 3636 3453 3644
rect 3947 3636 4053 3644
rect 4187 3636 4513 3644
rect 4527 3636 4673 3644
rect 5087 3636 5813 3644
rect 27 3616 533 3624
rect 1747 3616 1773 3624
rect 1787 3616 2393 3624
rect 3527 3616 4013 3624
rect 587 3596 693 3604
rect 1027 3596 1213 3604
rect 1647 3596 2213 3604
rect 2347 3596 3324 3604
rect 3316 3587 3324 3596
rect 3367 3596 4033 3604
rect 4167 3596 4193 3604
rect 4247 3596 4613 3604
rect 4747 3596 5113 3604
rect 5127 3596 5313 3604
rect 727 3576 993 3584
rect 1087 3576 1133 3584
rect 1327 3576 1593 3584
rect 1727 3576 2413 3584
rect 2907 3576 3033 3584
rect 3316 3576 3333 3587
rect 3320 3573 3333 3576
rect 3747 3576 4173 3584
rect 4767 3576 5353 3584
rect 5536 3576 5593 3584
rect 447 3556 533 3564
rect 547 3556 933 3564
rect 3227 3556 3573 3564
rect 3667 3556 3713 3564
rect 3787 3556 4073 3564
rect 4507 3556 4593 3564
rect 4607 3556 4733 3564
rect 4927 3556 5073 3564
rect 5536 3564 5544 3576
rect 5207 3556 5544 3564
rect 5567 3556 5613 3564
rect 327 3536 353 3544
rect 367 3536 653 3544
rect 667 3536 1093 3544
rect 1107 3536 1273 3544
rect 1287 3536 1313 3544
rect 2487 3536 2593 3544
rect 2607 3536 2713 3544
rect 3507 3536 3553 3544
rect 3847 3536 3953 3544
rect 4247 3536 4273 3544
rect 5096 3536 5224 3544
rect 127 3516 213 3524
rect 447 3516 773 3524
rect 827 3517 853 3525
rect 56 3487 64 3513
rect 256 3467 264 3514
rect 1136 3516 1173 3524
rect 427 3475 453 3483
rect 707 3475 793 3483
rect 1016 3484 1024 3513
rect 967 3476 1024 3484
rect 1136 3484 1144 3516
rect 1447 3517 1473 3525
rect 1607 3517 1653 3525
rect 1667 3516 1833 3524
rect 1887 3516 1993 3524
rect 2147 3517 2173 3525
rect 2187 3516 2233 3524
rect 2287 3517 2313 3525
rect 2407 3516 2433 3524
rect 2447 3516 2473 3524
rect 2527 3517 2553 3525
rect 2647 3517 2673 3525
rect 2867 3517 2893 3525
rect 3047 3517 3093 3525
rect 2756 3487 2764 3514
rect 1107 3476 1144 3484
rect 1767 3476 1784 3484
rect 87 3456 133 3464
rect 1207 3456 1613 3464
rect 1776 3464 1784 3476
rect 1867 3475 1913 3483
rect 2027 3476 2173 3484
rect 2367 3475 2413 3483
rect 2756 3476 2773 3487
rect 2760 3473 2773 3476
rect 1776 3456 1853 3464
rect 2796 3464 2804 3514
rect 2987 3476 3033 3484
rect 3247 3476 3273 3484
rect 3396 3484 3404 3514
rect 3616 3504 3624 3514
rect 3616 3496 3724 3504
rect 3396 3476 3553 3484
rect 3716 3484 3724 3496
rect 3996 3487 4004 3514
rect 4147 3517 4393 3525
rect 4416 3516 4453 3524
rect 3716 3476 3733 3484
rect 3747 3476 3853 3484
rect 3996 3476 4013 3487
rect 4000 3473 4013 3476
rect 2587 3456 2804 3464
rect 2907 3456 3193 3464
rect 3347 3456 3513 3464
rect 4056 3464 4064 3513
rect 4416 3504 4424 3516
rect 4467 3516 4573 3524
rect 4787 3517 4833 3525
rect 4887 3516 4953 3524
rect 4356 3496 4424 3504
rect 4127 3476 4273 3484
rect 4356 3486 4364 3496
rect 4996 3487 5004 3513
rect 4407 3476 4593 3484
rect 4867 3476 4913 3484
rect 5096 3486 5104 3536
rect 5176 3516 5193 3524
rect 5176 3487 5184 3516
rect 5216 3486 5224 3536
rect 5547 3536 5633 3544
rect 5236 3487 5244 3514
rect 5393 3504 5407 3513
rect 5393 3500 5444 3504
rect 5396 3496 5444 3500
rect 5236 3476 5253 3487
rect 5240 3473 5253 3476
rect 5347 3476 5413 3484
rect 5436 3484 5444 3496
rect 5436 3476 5493 3484
rect 5556 3484 5564 3513
rect 5687 3517 5753 3525
rect 5556 3476 5613 3484
rect 5747 3476 5793 3484
rect 4056 3456 4093 3464
rect 5027 3456 5053 3464
rect 767 3436 793 3444
rect 927 3436 1053 3444
rect 1227 3436 2733 3444
rect 3867 3436 3933 3444
rect 4307 3436 4473 3444
rect 4787 3436 4853 3444
rect 4987 3436 5253 3444
rect 5267 3436 5473 3444
rect 5487 3436 5573 3444
rect 1947 3416 2053 3424
rect 2327 3416 2613 3424
rect 2787 3416 3233 3424
rect 3567 3416 3653 3424
rect 3727 3416 4073 3424
rect 4727 3416 4813 3424
rect 5207 3416 5273 3424
rect 187 3396 353 3404
rect 887 3396 1393 3404
rect 1527 3396 1553 3404
rect 1787 3396 1813 3404
rect 2087 3396 2493 3404
rect 2987 3396 3053 3404
rect 3167 3396 3233 3404
rect 3576 3396 3753 3404
rect 487 3376 713 3384
rect 867 3376 1213 3384
rect 1727 3376 1793 3384
rect 1867 3376 1973 3384
rect 3576 3384 3584 3396
rect 3767 3396 3813 3404
rect 3907 3396 4293 3404
rect 4627 3396 4893 3404
rect 5367 3396 5653 3404
rect 2687 3376 3584 3384
rect 4767 3376 4813 3384
rect 107 3356 193 3364
rect 607 3356 953 3364
rect 967 3356 1893 3364
rect 2027 3356 2113 3364
rect 3307 3356 3593 3364
rect 3607 3356 3773 3364
rect 5287 3356 5493 3364
rect 5707 3356 5733 3364
rect 987 3336 1293 3344
rect 1647 3336 1733 3344
rect 2727 3336 2933 3344
rect 3507 3336 3573 3344
rect 3587 3336 3713 3344
rect 4207 3336 4413 3344
rect 4687 3336 5233 3344
rect 87 3324 100 3327
rect 87 3313 104 3324
rect 2507 3316 2553 3324
rect 2567 3316 2733 3324
rect 3367 3316 3393 3324
rect 3527 3316 3673 3324
rect 4887 3316 4933 3324
rect 56 3267 64 3293
rect 96 3247 104 3313
rect 216 3284 224 3294
rect 327 3296 373 3304
rect 447 3297 473 3305
rect 496 3296 593 3304
rect 216 3276 264 3284
rect 167 3255 233 3263
rect 256 3264 264 3276
rect 496 3266 504 3296
rect 687 3297 753 3305
rect 1067 3297 1093 3305
rect 1107 3296 1173 3304
rect 1347 3296 1464 3304
rect 1247 3276 1404 3284
rect 256 3256 353 3264
rect 547 3256 613 3264
rect 1396 3266 1404 3276
rect 1456 3266 1464 3296
rect 1847 3296 1873 3304
rect 2807 3296 2824 3304
rect 987 3256 1033 3264
rect 1296 3256 1313 3264
rect 87 3236 104 3247
rect 87 3233 100 3236
rect 747 3236 813 3244
rect 1296 3244 1304 3256
rect 1627 3255 1673 3263
rect 2016 3264 2024 3294
rect 2176 3276 2253 3284
rect 1987 3256 2024 3264
rect 2176 3264 2184 3276
rect 2616 3276 2713 3284
rect 2616 3266 2624 3276
rect 2816 3284 2824 3296
rect 2847 3297 2873 3305
rect 3027 3297 3073 3305
rect 3256 3296 3333 3304
rect 3256 3284 3264 3296
rect 3376 3296 3453 3304
rect 3376 3284 3384 3296
rect 3507 3297 3633 3305
rect 3647 3296 3733 3304
rect 3747 3296 4013 3304
rect 4347 3297 4373 3305
rect 4487 3296 4513 3304
rect 2816 3276 2904 3284
rect 2147 3256 2184 3264
rect 2747 3256 2773 3264
rect 2896 3264 2904 3276
rect 3136 3276 3264 3284
rect 3356 3276 3384 3284
rect 3136 3266 3144 3276
rect 3356 3266 3364 3276
rect 2896 3256 2913 3264
rect 3687 3255 3713 3263
rect 3867 3255 3893 3263
rect 3967 3255 4193 3263
rect 4436 3247 4444 3294
rect 4587 3297 4613 3305
rect 4687 3296 4924 3304
rect 4467 3256 4553 3264
rect 4567 3256 4713 3264
rect 4916 3266 4924 3296
rect 5007 3297 5073 3305
rect 4807 3255 4833 3263
rect 5047 3255 5113 3263
rect 5176 3264 5184 3313
rect 5247 3296 5313 3304
rect 5567 3297 5693 3305
rect 5176 3256 5213 3264
rect 5407 3255 5593 3263
rect 1167 3236 1304 3244
rect 2207 3236 2433 3244
rect 2447 3236 2573 3244
rect 2587 3236 2673 3244
rect 4667 3236 4693 3244
rect 4967 3236 5153 3244
rect 1227 3216 1793 3224
rect 3087 3216 3433 3224
rect 3887 3216 4753 3224
rect 4767 3216 4853 3224
rect 5267 3216 5413 3224
rect 5467 3216 5573 3224
rect 147 3196 353 3204
rect 367 3196 793 3204
rect 807 3196 853 3204
rect 1007 3196 1093 3204
rect 1267 3196 1293 3204
rect 1367 3196 1513 3204
rect 3307 3196 3593 3204
rect 4527 3196 5213 3204
rect 1047 3176 1213 3184
rect 1587 3176 2193 3184
rect 3447 3176 3553 3184
rect 407 3156 3073 3164
rect 3607 3156 4213 3164
rect 4227 3156 4413 3164
rect 5107 3156 5273 3164
rect 2047 3136 2073 3144
rect 387 3116 433 3124
rect 1347 3116 1693 3124
rect 2327 3116 3313 3124
rect 3487 3116 3693 3124
rect 4127 3116 4173 3124
rect 807 3096 1493 3104
rect 1087 3076 1633 3084
rect 1647 3076 2233 3084
rect 2687 3076 2813 3084
rect 2827 3076 3073 3084
rect 3087 3076 3473 3084
rect 3947 3076 4033 3084
rect 4047 3076 4533 3084
rect 4687 3076 4953 3084
rect 5707 3076 5813 3084
rect 507 3056 573 3064
rect 1127 3056 1273 3064
rect 1827 3056 2013 3064
rect 4596 3056 4913 3064
rect 587 3036 673 3044
rect 1847 3036 1893 3044
rect 2207 3036 2233 3044
rect 2247 3036 2633 3044
rect 2907 3036 3393 3044
rect 3627 3036 3773 3044
rect 4027 3036 4333 3044
rect 4596 3044 4604 3056
rect 4347 3036 4604 3044
rect 4627 3036 4713 3044
rect 5087 3036 5133 3044
rect 5147 3036 5213 3044
rect 5647 3036 5773 3044
rect 47 3016 113 3024
rect 167 3016 273 3024
rect 927 3016 993 3024
rect 2167 3016 2273 3024
rect 2287 3016 2413 3024
rect 2427 3016 2453 3024
rect 2936 3016 3233 3024
rect 2936 3008 2944 3016
rect 5027 3016 5133 3024
rect 5327 3016 5373 3024
rect 5387 3016 5493 3024
rect 5507 3016 5533 3024
rect -24 2996 73 3004
rect 120 3004 133 3007
rect 116 2993 133 3004
rect 227 2996 393 3004
rect 467 2996 633 3004
rect 647 2997 693 3005
rect 747 2997 773 3005
rect 867 2996 1073 3004
rect 1096 2996 1113 3004
rect 116 2966 124 2993
rect 1096 2984 1104 2996
rect 1127 2996 1193 3004
rect 676 2976 724 2984
rect 347 2956 433 2964
rect 607 2956 633 2964
rect 676 2966 684 2976
rect 716 2964 724 2976
rect 1076 2976 1104 2984
rect 716 2956 873 2964
rect 1076 2964 1084 2976
rect 987 2956 1084 2964
rect 1236 2964 1244 2994
rect 1187 2956 1244 2964
rect 1336 2964 1344 2994
rect 1487 2996 1513 3004
rect 1867 2996 1953 3004
rect 2487 2997 2733 3005
rect 2827 2996 2933 3004
rect 2776 2984 2784 2994
rect 3007 2996 3033 3004
rect 3167 2997 3193 3005
rect 3396 2996 3473 3004
rect 2716 2976 2784 2984
rect 1267 2956 1344 2964
rect 1647 2955 1673 2963
rect 1907 2955 1933 2963
rect 1987 2956 2173 2964
rect 2247 2955 2353 2963
rect 2716 2964 2724 2976
rect 2667 2956 2724 2964
rect 2747 2956 2793 2964
rect 2847 2955 2893 2963
rect 3067 2956 3153 2964
rect 3396 2966 3404 2996
rect 3487 2996 3633 3004
rect 3987 2997 4013 3005
rect 4087 2996 4173 3004
rect 4267 2997 4293 3005
rect 4727 2996 4753 3004
rect 4767 2997 4793 3005
rect 5076 2996 5113 3004
rect 927 2936 953 2944
rect 1107 2936 1153 2944
rect 1276 2936 1493 2944
rect 407 2916 713 2924
rect 1276 2924 1284 2936
rect 1707 2936 1764 2944
rect 787 2916 1284 2924
rect 1487 2916 1713 2924
rect 1756 2924 1764 2936
rect 3327 2936 3353 2944
rect 3507 2936 3573 2944
rect 1756 2916 2293 2924
rect 2707 2916 2753 2924
rect 2767 2916 2873 2924
rect 2887 2916 3093 2924
rect 3496 2924 3504 2933
rect 3267 2916 3504 2924
rect 3816 2924 3824 2994
rect 4516 2976 4613 2984
rect 3847 2956 3873 2964
rect 4127 2956 4153 2964
rect 4327 2956 4373 2964
rect 4387 2956 4413 2964
rect 4516 2964 4524 2976
rect 4467 2956 4524 2964
rect 4676 2964 4684 2994
rect 5036 2967 5044 2994
rect 4567 2956 4684 2964
rect 4887 2956 4933 2964
rect 5027 2956 5044 2967
rect 5027 2953 5040 2956
rect 5076 2947 5084 2996
rect 5356 2964 5364 2994
rect 5427 2996 5473 3004
rect 5667 2996 5733 3004
rect 5787 2997 5813 3005
rect 5356 2956 5493 2964
rect 5627 2955 5653 2963
rect 4627 2936 4693 2944
rect 5167 2936 5213 2944
rect 5547 2936 5753 2944
rect 3816 2916 3913 2924
rect 3987 2916 4013 2924
rect 4027 2916 4053 2924
rect 4647 2916 4813 2924
rect 5007 2916 5053 2924
rect 907 2896 1133 2904
rect 1147 2896 1353 2904
rect 1367 2896 1393 2904
rect 1507 2896 1693 2904
rect 1787 2896 1973 2904
rect 2027 2896 2053 2904
rect 2107 2896 2804 2904
rect 2796 2884 2804 2896
rect 4767 2896 4813 2904
rect 5507 2896 5553 2904
rect 5567 2896 5673 2904
rect 227 2876 2084 2884
rect 2796 2876 2953 2884
rect 2076 2867 2084 2876
rect 3967 2876 4193 2884
rect 4207 2876 4253 2884
rect 4267 2876 4833 2884
rect 5147 2876 5333 2884
rect 5427 2876 5473 2884
rect 67 2856 133 2864
rect 1227 2856 1613 2864
rect 2087 2856 2373 2864
rect 2427 2856 2473 2864
rect 3467 2856 3533 2864
rect 1247 2836 1273 2844
rect 2047 2836 2093 2844
rect 4387 2836 4593 2844
rect 4647 2836 4753 2844
rect 4807 2836 4893 2844
rect 5067 2836 5293 2844
rect 5467 2836 5553 2844
rect 5707 2836 5793 2844
rect 2387 2816 2973 2824
rect 2987 2816 3333 2824
rect 3347 2816 3673 2824
rect 3687 2816 3693 2824
rect 3827 2816 3993 2824
rect 4787 2816 4913 2824
rect 4967 2816 5013 2824
rect 5027 2816 5413 2824
rect 47 2796 153 2804
rect 507 2796 553 2804
rect 1107 2796 1193 2804
rect 1427 2796 1493 2804
rect 1507 2796 1633 2804
rect 1907 2796 2013 2804
rect 2067 2796 2153 2804
rect 2927 2796 2953 2804
rect 4027 2796 4233 2804
rect 4347 2796 4373 2804
rect 4947 2796 5113 2804
rect 5167 2796 5293 2804
rect 367 2776 433 2784
rect 447 2776 473 2784
rect 16 2747 24 2773
rect -24 2724 -16 2744
rect 347 2736 393 2744
rect 896 2746 904 2793
rect 1007 2776 1033 2784
rect 1120 2784 1133 2787
rect 1116 2773 1133 2784
rect 1347 2777 1393 2785
rect 1547 2776 1593 2784
rect 1667 2776 1693 2784
rect 1747 2776 1773 2784
rect 1787 2777 1853 2785
rect 1896 2776 2033 2784
rect 1116 2746 1124 2773
rect 1176 2747 1184 2773
rect 467 2735 573 2743
rect 1047 2735 1073 2743
rect 1896 2746 1904 2776
rect 2187 2776 2213 2784
rect 2287 2777 2313 2785
rect 2327 2776 2373 2784
rect 2487 2777 2613 2785
rect 2627 2777 2653 2785
rect 2787 2776 2833 2784
rect 2907 2776 2993 2784
rect 3136 2776 3213 2784
rect 2536 2756 2593 2764
rect 1227 2735 1413 2743
rect 1627 2735 1652 2743
rect 1676 2740 1713 2744
rect 1673 2736 1713 2740
rect 1673 2727 1687 2736
rect 2047 2735 2073 2743
rect 2167 2735 2233 2743
rect 2536 2744 2544 2756
rect 3136 2746 3144 2776
rect 3747 2777 3953 2785
rect 4127 2776 4173 2784
rect 4307 2777 4433 2785
rect 4456 2776 4493 2784
rect 4456 2764 4464 2776
rect 4607 2776 4733 2784
rect 5667 2777 5733 2785
rect 3276 2756 3924 2764
rect 3276 2746 3284 2756
rect 3556 2746 3564 2756
rect 2507 2736 2544 2744
rect 2727 2735 2773 2743
rect 2867 2735 2893 2743
rect 3207 2735 3273 2743
rect 3467 2735 3493 2743
rect 3916 2746 3924 2756
rect 4456 2756 4693 2764
rect 4456 2747 4464 2756
rect 4816 2747 4824 2773
rect 4876 2747 4884 2774
rect 3827 2736 3853 2744
rect 4047 2736 4153 2744
rect 4567 2736 4673 2744
rect 4867 2736 4884 2747
rect 4867 2733 4880 2736
rect 4927 2735 5093 2743
rect 5107 2735 5113 2743
rect 5136 2727 5144 2774
rect 5187 2736 5193 2744
rect 5207 2736 5253 2744
rect 5407 2736 5493 2744
rect -24 2716 93 2724
rect 1267 2716 1393 2724
rect 1407 2716 1533 2724
rect 2447 2716 2453 2724
rect 2467 2716 2553 2724
rect 2627 2716 2813 2724
rect 3947 2716 3973 2724
rect 4067 2716 4144 2724
rect 1307 2696 1353 2704
rect 1667 2696 2273 2704
rect 2347 2696 2673 2704
rect 3107 2696 3293 2704
rect 3447 2696 3473 2704
rect 3567 2696 3613 2704
rect 3687 2696 4093 2704
rect 4136 2704 4144 2716
rect 4287 2716 4473 2724
rect 4487 2716 4773 2724
rect 5047 2716 5073 2724
rect 5527 2716 5753 2724
rect 4136 2696 4404 2704
rect 4396 2687 4404 2696
rect 4547 2696 4653 2704
rect 4667 2696 4853 2704
rect 5167 2696 5213 2704
rect 5327 2696 5433 2704
rect 5447 2696 5633 2704
rect 5876 2704 5884 2744
rect 5827 2696 5884 2704
rect 47 2676 273 2684
rect 287 2676 673 2684
rect 687 2676 853 2684
rect 1587 2676 1853 2684
rect 1867 2676 2193 2684
rect 4267 2676 4333 2684
rect 4407 2676 4513 2684
rect 5567 2676 5653 2684
rect 1027 2656 1473 2664
rect 1967 2656 2453 2664
rect 3547 2656 3793 2664
rect 3967 2656 4052 2664
rect 4087 2656 4353 2664
rect 5087 2656 5393 2664
rect 5767 2656 5813 2664
rect 3047 2636 3193 2644
rect 4107 2636 4593 2644
rect 4707 2636 4973 2644
rect 4987 2636 5133 2644
rect 5347 2636 5453 2644
rect 2347 2616 2933 2624
rect 3907 2616 4033 2624
rect 4427 2616 5833 2624
rect 1807 2596 1953 2604
rect 2476 2596 3153 2604
rect 167 2576 193 2584
rect 2476 2584 2484 2596
rect 3487 2596 3753 2604
rect 3807 2596 4193 2604
rect 4207 2596 5753 2604
rect 1907 2576 2484 2584
rect 2507 2576 3133 2584
rect 3787 2576 4273 2584
rect 4287 2576 4333 2584
rect 4447 2576 4473 2584
rect 4487 2576 4613 2584
rect 4687 2576 4953 2584
rect 287 2556 313 2564
rect 327 2556 373 2564
rect 1747 2556 1833 2564
rect 3727 2556 4413 2564
rect 4716 2556 4753 2564
rect 787 2536 1093 2544
rect 1107 2536 1253 2544
rect 1267 2536 1393 2544
rect 2927 2536 2973 2544
rect 3607 2536 3653 2544
rect 3927 2536 3953 2544
rect 4716 2544 4724 2556
rect 4807 2556 4913 2564
rect 4627 2536 4724 2544
rect 4747 2536 4873 2544
rect 5567 2536 5753 2544
rect 2107 2516 2613 2524
rect 2667 2516 2693 2524
rect 2707 2516 2753 2524
rect 3147 2516 3313 2524
rect 3527 2516 3673 2524
rect 4187 2516 4293 2524
rect 5007 2516 5053 2524
rect 5107 2516 5272 2524
rect 5307 2516 5664 2524
rect 87 2496 133 2504
rect 467 2496 493 2504
rect 567 2496 673 2504
rect 687 2496 713 2504
rect 2987 2496 3353 2504
rect 3367 2496 3473 2504
rect 3767 2496 3893 2504
rect 4527 2504 4540 2507
rect 4527 2493 4544 2504
rect 4587 2496 4753 2504
rect 5656 2504 5664 2516
rect 5656 2496 5804 2504
rect 76 2427 84 2474
rect 227 2476 253 2484
rect 447 2476 613 2484
rect 927 2477 953 2485
rect 1167 2477 1193 2485
rect 1447 2477 1492 2485
rect 107 2436 133 2444
rect 147 2435 193 2443
rect 567 2436 653 2444
rect 727 2435 753 2443
rect 816 2444 824 2474
rect 1296 2464 1304 2474
rect 1296 2456 1473 2464
rect 816 2436 973 2444
rect 1047 2435 1073 2443
rect 1087 2436 1133 2444
rect 1207 2436 1233 2444
rect 1327 2436 1413 2444
rect 1447 2416 1473 2424
rect 1516 2424 1524 2474
rect 1736 2446 1744 2493
rect 1767 2476 1853 2484
rect 2147 2477 2173 2485
rect 2367 2477 2393 2485
rect 2527 2477 2553 2485
rect 2576 2476 2593 2484
rect 2236 2464 2244 2474
rect 2576 2464 2584 2476
rect 2747 2476 2773 2484
rect 2787 2476 2813 2484
rect 3107 2476 3133 2484
rect 2936 2464 2944 2474
rect 3407 2477 3433 2485
rect 3647 2476 3713 2484
rect 3827 2477 3853 2485
rect 3920 2484 3933 2487
rect 2236 2456 2584 2464
rect 2876 2456 2944 2464
rect 3016 2456 3304 2464
rect 1987 2435 2013 2443
rect 2187 2436 2213 2444
rect 2227 2436 2273 2444
rect 1516 2416 1553 2424
rect 1927 2416 2113 2424
rect 2296 2424 2304 2456
rect 2367 2436 2573 2444
rect 2627 2435 2653 2443
rect 2876 2444 2884 2456
rect 2847 2436 2884 2444
rect 3016 2444 3024 2456
rect 2907 2436 3024 2444
rect 3247 2436 3273 2444
rect 3296 2444 3304 2456
rect 3296 2436 3493 2444
rect 3516 2444 3524 2473
rect 3773 2464 3787 2473
rect 3916 2473 3933 2484
rect 4027 2476 4053 2484
rect 3916 2464 3924 2473
rect 3716 2460 3787 2464
rect 3716 2456 3784 2460
rect 3896 2456 3924 2464
rect 3716 2444 3724 2456
rect 3507 2436 3524 2444
rect 3656 2436 3724 2444
rect 2247 2416 2304 2424
rect 2967 2416 3133 2424
rect 3347 2416 3393 2424
rect 3656 2424 3664 2436
rect 3747 2436 3812 2444
rect 3896 2444 3904 2456
rect 3847 2436 3904 2444
rect 3947 2436 4204 2444
rect 3587 2416 3664 2424
rect 3887 2416 4053 2424
rect 4196 2424 4204 2436
rect 4256 2427 4264 2474
rect 4353 2464 4367 2473
rect 4396 2464 4404 2474
rect 4353 2460 4404 2464
rect 4356 2456 4404 2460
rect 4196 2416 4244 2424
rect 967 2396 1273 2404
rect 1367 2396 1573 2404
rect 2527 2396 2713 2404
rect 3387 2396 3453 2404
rect 3527 2396 3833 2404
rect 4236 2404 4244 2416
rect 4347 2416 4453 2424
rect 4476 2416 4513 2424
rect 4236 2396 4373 2404
rect 4476 2404 4484 2416
rect 4536 2424 4544 2493
rect 4667 2476 4713 2484
rect 4856 2476 4913 2484
rect 4616 2444 4624 2473
rect 4567 2436 4633 2444
rect 4856 2444 4864 2476
rect 4927 2476 5053 2484
rect 5076 2446 5084 2493
rect 5116 2476 5213 2484
rect 5116 2446 5124 2476
rect 5287 2477 5313 2485
rect 5447 2476 5473 2484
rect 5516 2464 5524 2493
rect 5547 2477 5593 2485
rect 5647 2476 5733 2484
rect 5496 2456 5524 2464
rect 5496 2446 5504 2456
rect 4787 2436 4864 2444
rect 5207 2436 5413 2444
rect 5567 2435 5653 2443
rect 5667 2436 5692 2444
rect 5776 2444 5784 2473
rect 5796 2464 5804 2496
rect 5847 2476 5884 2484
rect 5796 2456 5824 2464
rect 5727 2436 5784 2444
rect 5816 2447 5824 2456
rect 5816 2436 5833 2447
rect 5820 2433 5833 2436
rect 4536 2416 4593 2424
rect 4747 2416 4833 2424
rect 4987 2416 5053 2424
rect 5267 2416 5293 2424
rect 4387 2396 4484 2404
rect 4496 2396 4573 2404
rect 627 2376 793 2384
rect 987 2376 1253 2384
rect 1307 2376 2073 2384
rect 2187 2376 2333 2384
rect 2347 2376 2373 2384
rect 2507 2376 2573 2384
rect 3427 2376 3553 2384
rect 4167 2376 4353 2384
rect 4496 2384 4504 2396
rect 4907 2396 5133 2404
rect 5447 2396 5593 2404
rect 4367 2376 4504 2384
rect 4556 2376 4692 2384
rect 1507 2356 1833 2364
rect 1847 2356 1893 2364
rect 2107 2356 2593 2364
rect 4227 2356 4333 2364
rect 4556 2364 4564 2376
rect 4727 2376 5193 2384
rect 5267 2376 5333 2384
rect 4427 2356 4564 2364
rect 4627 2356 4673 2364
rect 5527 2356 5573 2364
rect 5627 2356 5673 2364
rect 1087 2336 1673 2344
rect 2347 2336 2873 2344
rect 2887 2336 2993 2344
rect 3147 2336 3213 2344
rect 3267 2336 3753 2344
rect 4587 2344 4600 2347
rect 4587 2333 4604 2344
rect 2087 2316 2273 2324
rect 3213 2324 3227 2333
rect 3213 2320 3513 2324
rect 3216 2316 3513 2320
rect 4596 2324 4604 2333
rect 4687 2336 4933 2344
rect 4947 2336 5033 2344
rect 5167 2336 5193 2344
rect 5347 2336 5433 2344
rect 5447 2336 5493 2344
rect 4596 2316 4893 2324
rect 5427 2316 5533 2324
rect 5587 2316 5613 2324
rect 5847 2316 5884 2324
rect 127 2296 213 2304
rect 627 2296 1013 2304
rect 1027 2296 1093 2304
rect 1487 2296 1573 2304
rect 1587 2296 1633 2304
rect 1647 2296 1753 2304
rect 1827 2296 1873 2304
rect 1887 2296 2024 2304
rect 547 2276 593 2284
rect 967 2276 1193 2284
rect 1207 2284 1220 2287
rect 2016 2284 2024 2296
rect 2427 2296 2673 2304
rect 2787 2296 2833 2304
rect 3167 2296 3393 2304
rect 3687 2296 3913 2304
rect 3927 2296 4053 2304
rect 4067 2296 4193 2304
rect 4207 2296 4233 2304
rect 4287 2296 4553 2304
rect 4647 2296 4953 2304
rect 5007 2296 5033 2304
rect 5127 2296 5253 2304
rect 5347 2296 5373 2304
rect 5487 2296 5513 2304
rect 1207 2276 1224 2284
rect 2016 2276 2093 2284
rect 1207 2274 1220 2276
rect 1200 2273 1220 2274
rect 2827 2276 2893 2284
rect 3567 2276 3593 2284
rect 167 2257 192 2265
rect 227 2256 273 2264
rect 407 2256 453 2264
rect 587 2256 653 2264
rect 147 2215 213 2223
rect 696 2224 704 2254
rect 767 2256 793 2264
rect 847 2257 893 2265
rect 1127 2256 1193 2264
rect 1247 2257 1293 2265
rect 1307 2256 1373 2264
rect 1527 2256 1553 2264
rect 1567 2256 1633 2264
rect 2127 2256 2324 2264
rect 696 2216 813 2224
rect 867 2216 933 2224
rect 1027 2215 1053 2223
rect 1267 2216 1353 2224
rect 1407 2216 1493 2224
rect 1787 2215 1813 2223
rect 1996 2207 2004 2254
rect 2316 2227 2324 2256
rect 2487 2256 2533 2264
rect 2560 2264 2572 2267
rect 2556 2253 2572 2264
rect 2607 2256 2653 2264
rect 2107 2215 2193 2223
rect 2556 2226 2564 2253
rect 2936 2227 2944 2254
rect 3027 2256 3133 2264
rect 3360 2264 3373 2267
rect 2447 2215 2473 2223
rect 2687 2215 2713 2223
rect 2927 2216 2944 2227
rect 2927 2213 2940 2216
rect 3007 2216 3133 2224
rect 3176 2224 3184 2254
rect 3356 2253 3373 2264
rect 3176 2216 3272 2224
rect 3356 2224 3364 2253
rect 3456 2224 3464 2254
rect 3616 2264 3624 2293
rect 5587 2296 5633 2304
rect 5707 2296 5733 2304
rect 5876 2296 5884 2316
rect 3596 2256 3624 2264
rect 3307 2216 3364 2224
rect 3416 2220 3464 2224
rect 3413 2216 3464 2220
rect 3413 2207 3427 2216
rect 3536 2224 3544 2253
rect 3596 2226 3604 2256
rect 3527 2216 3544 2224
rect 3707 2215 3733 2223
rect 3796 2224 3804 2253
rect 3936 2244 3944 2273
rect 4180 2264 4193 2267
rect 4027 2256 4044 2264
rect 4036 2244 4044 2256
rect 4176 2253 4193 2264
rect 4333 2264 4347 2273
rect 5387 2276 5453 2284
rect 5547 2276 5624 2284
rect 4307 2260 4347 2264
rect 4307 2256 4344 2260
rect 4567 2256 4673 2264
rect 4767 2257 4813 2265
rect 4867 2256 4884 2264
rect 3936 2236 4024 2244
rect 4036 2236 4064 2244
rect 3787 2216 3804 2224
rect 3967 2215 3993 2223
rect 4016 2224 4024 2236
rect 4016 2216 4033 2224
rect 4056 2224 4064 2236
rect 4056 2216 4113 2224
rect 4176 2226 4184 2253
rect 4396 2244 4404 2254
rect 4376 2236 4404 2244
rect 4376 2224 4384 2236
rect 4876 2227 4884 2256
rect 5007 2256 5153 2264
rect 5167 2256 5253 2264
rect 5347 2264 5360 2267
rect 5347 2253 5364 2264
rect 5296 2227 5304 2253
rect 5356 2244 5364 2253
rect 5436 2256 5573 2264
rect 5356 2236 5404 2244
rect 4347 2216 4384 2224
rect 4727 2216 4833 2224
rect 4987 2216 5053 2224
rect 5067 2215 5133 2223
rect 5296 2216 5313 2227
rect 5300 2213 5313 2216
rect 5396 2226 5404 2236
rect 5436 2227 5444 2256
rect 5616 2226 5624 2276
rect 5807 2276 5833 2284
rect 687 2196 853 2204
rect 1227 2196 1393 2204
rect 1847 2196 1913 2204
rect 2147 2196 2173 2204
rect 3127 2196 3233 2204
rect 4067 2196 4133 2204
rect 5536 2204 5544 2212
rect 5756 2207 5764 2254
rect 5876 2244 5884 2264
rect 5876 2236 5904 2244
rect 5807 2216 5884 2224
rect 5407 2196 5544 2204
rect 5647 2196 5713 2204
rect 467 2176 553 2184
rect 707 2176 813 2184
rect 947 2176 1093 2184
rect 1307 2176 1333 2184
rect 1547 2176 1613 2184
rect 1627 2176 2093 2184
rect 2447 2176 2553 2184
rect 2607 2176 2813 2184
rect 3236 2184 3244 2193
rect 3236 2176 3353 2184
rect 3527 2176 3753 2184
rect 3827 2176 3873 2184
rect 4007 2176 4333 2184
rect 4387 2176 4473 2184
rect 4587 2176 4853 2184
rect 5007 2176 5233 2184
rect 5347 2176 5493 2184
rect 5896 2184 5904 2236
rect 5787 2176 5904 2184
rect 427 2156 753 2164
rect 1747 2156 1933 2164
rect 1947 2156 1973 2164
rect 2267 2156 2673 2164
rect 2907 2156 3012 2164
rect 3047 2156 3553 2164
rect 4327 2156 4653 2164
rect 5087 2156 5193 2164
rect 5236 2156 5753 2164
rect 527 2136 613 2144
rect 827 2136 893 2144
rect 2187 2136 2413 2144
rect 2427 2136 2513 2144
rect 2527 2136 2733 2144
rect 3707 2136 3813 2144
rect 4047 2136 4093 2144
rect 4107 2136 4273 2144
rect 4427 2136 4793 2144
rect 4907 2136 4964 2144
rect 1667 2116 1773 2124
rect 2127 2116 2553 2124
rect 3347 2116 3413 2124
rect 3607 2116 4093 2124
rect 4167 2116 4393 2124
rect 4547 2116 4593 2124
rect 4767 2116 4933 2124
rect 4956 2124 4964 2136
rect 5236 2144 5244 2156
rect 5167 2136 5244 2144
rect 5367 2136 5453 2144
rect 5687 2136 5773 2144
rect 4956 2116 5133 2124
rect 5327 2116 5452 2124
rect 107 2096 253 2104
rect 267 2096 373 2104
rect 387 2096 513 2104
rect 867 2096 1833 2104
rect 2787 2096 3113 2104
rect 3167 2096 3313 2104
rect 3327 2096 3493 2104
rect 3507 2096 3773 2104
rect 3867 2096 4464 2104
rect 2147 2076 2393 2084
rect 2567 2076 2913 2084
rect 3147 2076 3453 2084
rect 3467 2076 3804 2084
rect 907 2056 1073 2064
rect 1227 2056 1573 2064
rect 1767 2056 2033 2064
rect 3067 2056 3613 2064
rect 3627 2056 3713 2064
rect 3796 2064 3804 2076
rect 3827 2076 4053 2084
rect 4287 2076 4313 2084
rect 4456 2084 4464 2096
rect 4933 2104 4947 2113
rect 5487 2116 5573 2124
rect 4487 2100 4947 2104
rect 4487 2096 4944 2100
rect 5207 2096 5433 2104
rect 4456 2076 4553 2084
rect 4887 2076 5093 2084
rect 3796 2056 3993 2064
rect 4387 2056 4593 2064
rect 5207 2056 5513 2064
rect 547 2036 853 2044
rect 1847 2036 2033 2044
rect 2056 2036 2133 2044
rect 727 2016 813 2024
rect 967 2016 1453 2024
rect 1647 2016 1693 2024
rect 2056 2024 2064 2036
rect 2207 2036 2233 2044
rect 2247 2036 2453 2044
rect 2476 2036 2693 2044
rect 1907 2016 2064 2024
rect 2167 2016 2193 2024
rect 2476 2024 2484 2036
rect 2907 2036 3152 2044
rect 3187 2036 3253 2044
rect 3747 2036 4133 2044
rect 4407 2036 4533 2044
rect 4707 2036 4773 2044
rect 4787 2036 4813 2044
rect 4827 2036 4873 2044
rect 4967 2036 5093 2044
rect 5147 2036 5313 2044
rect 2207 2016 2484 2024
rect 2787 2016 2973 2024
rect 3107 2016 3593 2024
rect 4487 2016 4573 2024
rect 4667 2016 5073 2024
rect 5167 2016 5333 2024
rect 1267 1996 1304 2004
rect 127 1976 153 1984
rect 1027 1976 1153 1984
rect 47 1957 73 1965
rect 87 1956 213 1964
rect 267 1956 373 1964
rect 400 1964 412 1967
rect 396 1953 412 1964
rect 447 1956 473 1964
rect 487 1956 573 1964
rect 627 1957 673 1965
rect 1067 1957 1093 1965
rect 1167 1956 1273 1964
rect 396 1926 404 1953
rect 716 1927 724 1954
rect 756 1944 764 1954
rect 756 1936 944 1944
rect 507 1915 533 1923
rect 707 1916 724 1927
rect 707 1913 720 1916
rect 827 1916 913 1924
rect 936 1924 944 1936
rect 1296 1926 1304 1996
rect 1987 1996 2073 2004
rect 2747 1996 3073 2004
rect 3756 1996 4033 2004
rect 1687 1984 1700 1987
rect 1720 1984 1733 1987
rect 1687 1973 1704 1984
rect 1467 1957 1493 1965
rect 1596 1956 1653 1964
rect 1316 1944 1324 1954
rect 1316 1936 1353 1944
rect 936 1916 993 1924
rect 27 1896 133 1904
rect 207 1896 273 1904
rect 287 1896 313 1904
rect 787 1896 873 1904
rect 967 1896 1033 1904
rect 1416 1904 1424 1954
rect 1596 1927 1604 1956
rect 1696 1924 1704 1973
rect 1716 1973 1733 1984
rect 2667 1976 2764 1984
rect 1716 1926 1724 1973
rect 1847 1957 1873 1965
rect 1687 1916 1704 1924
rect 1767 1915 1813 1923
rect 1916 1907 1924 1973
rect 2507 1957 2533 1965
rect 2756 1964 2764 1976
rect 3487 1976 3653 1984
rect 3756 1984 3764 1996
rect 4127 1996 4373 2004
rect 4687 1996 4793 2004
rect 4867 1996 4913 2004
rect 4927 1996 4993 2004
rect 5067 1996 5233 2004
rect 3667 1976 3764 1984
rect 4107 1976 4284 1984
rect 2756 1956 2773 1964
rect 2973 1964 2987 1973
rect 2973 1960 3032 1964
rect 2976 1956 3032 1960
rect 2047 1916 2213 1924
rect 2296 1907 2304 1953
rect 2387 1915 2413 1923
rect 2427 1916 2573 1924
rect 2636 1924 2644 1954
rect 3147 1956 3204 1964
rect 2707 1936 2933 1944
rect 3053 1944 3067 1953
rect 2956 1940 3067 1944
rect 2956 1936 3064 1940
rect 2956 1927 2964 1936
rect 3196 1927 3204 1956
rect 2636 1916 2753 1924
rect 2956 1924 2973 1927
rect 2887 1916 2973 1924
rect 2960 1913 2973 1916
rect 3087 1915 3113 1923
rect 1327 1896 1424 1904
rect 1847 1896 1873 1904
rect 2296 1896 2313 1907
rect 2300 1893 2313 1896
rect 3276 1904 3284 1954
rect 3567 1956 3593 1964
rect 3747 1957 3773 1965
rect 3847 1956 3953 1964
rect 3967 1956 3993 1964
rect 4276 1967 4284 1976
rect 5127 1976 5333 1984
rect 5547 1976 5713 1984
rect 3296 1927 3304 1953
rect 4176 1944 4184 1954
rect 4246 1953 4247 1960
rect 4267 1964 4284 1967
rect 4267 1956 4293 1964
rect 4267 1953 4280 1956
rect 4347 1956 4373 1964
rect 4156 1940 4184 1944
rect 4233 1944 4247 1953
rect 4233 1940 4264 1944
rect 4153 1936 4184 1940
rect 4235 1936 4264 1940
rect 4153 1927 4167 1936
rect 3467 1916 3633 1924
rect 3687 1916 4033 1924
rect 4256 1927 4264 1936
rect 4207 1920 4244 1924
rect 4207 1916 4247 1920
rect 4256 1916 4273 1927
rect 4233 1907 4247 1916
rect 4260 1913 4273 1916
rect 4436 1924 4444 1954
rect 4567 1956 4673 1964
rect 4807 1957 4853 1965
rect 4493 1947 4507 1953
rect 4493 1946 4520 1947
rect 4493 1940 4513 1946
rect 4496 1936 4513 1940
rect 4500 1933 4513 1936
rect 4327 1916 4493 1924
rect 3167 1896 3284 1904
rect 3547 1896 3573 1904
rect 3887 1896 3913 1904
rect 4387 1896 4413 1904
rect 4556 1904 4564 1954
rect 4716 1924 4724 1954
rect 5007 1956 5053 1964
rect 5067 1956 5093 1964
rect 5367 1956 5444 1964
rect 4716 1916 4833 1924
rect 4956 1924 4964 1953
rect 5156 1927 5164 1953
rect 5193 1944 5207 1953
rect 5193 1940 5244 1944
rect 5196 1936 5244 1940
rect 4887 1916 4973 1924
rect 5236 1924 5244 1936
rect 5236 1916 5253 1924
rect 5276 1924 5284 1954
rect 5436 1927 5444 1956
rect 5276 1916 5344 1924
rect 5336 1907 5344 1916
rect 5476 1924 5484 1953
rect 5556 1927 5564 1954
rect 5827 1956 5884 1964
rect 5607 1936 5793 1944
rect 5476 1916 5493 1924
rect 5556 1916 5573 1927
rect 5560 1913 5573 1916
rect 4467 1896 4564 1904
rect 5076 1896 5213 1904
rect 5076 1887 5084 1896
rect 5336 1896 5353 1907
rect 5340 1893 5353 1896
rect 5707 1896 5813 1904
rect 1147 1876 1173 1884
rect 1227 1876 1433 1884
rect 1547 1876 1613 1884
rect 1687 1876 1753 1884
rect 2587 1876 2613 1884
rect 3167 1876 3273 1884
rect 3407 1876 3573 1884
rect 3647 1876 3753 1884
rect 4127 1876 4473 1884
rect 4527 1876 4553 1884
rect 4707 1876 4773 1884
rect 4816 1876 5073 1884
rect 107 1856 213 1864
rect 307 1856 673 1864
rect 687 1856 953 1864
rect 1427 1856 1473 1864
rect 1907 1856 2233 1864
rect 2347 1856 2433 1864
rect 2807 1856 3053 1864
rect 3627 1856 3713 1864
rect 3887 1856 4133 1864
rect 4267 1856 4433 1864
rect 4816 1864 4824 1876
rect 5247 1876 5313 1884
rect 4747 1856 4824 1864
rect 5107 1856 5153 1864
rect 5347 1856 5373 1864
rect 5667 1856 5813 1864
rect 387 1836 493 1844
rect 1107 1836 1213 1844
rect 1287 1836 1353 1844
rect 1367 1836 1553 1844
rect 1607 1836 1653 1844
rect 2547 1836 2684 1844
rect 427 1816 473 1824
rect 487 1816 592 1824
rect 627 1816 693 1824
rect 1507 1816 1953 1824
rect 2487 1816 2513 1824
rect 2676 1824 2684 1836
rect 2867 1836 2953 1844
rect 3227 1836 3433 1844
rect 3807 1836 4113 1844
rect 4267 1836 4413 1844
rect 4887 1836 5204 1844
rect 2676 1816 2913 1824
rect 3067 1816 3193 1824
rect 3247 1816 3333 1824
rect 3727 1816 3893 1824
rect 4147 1816 4293 1824
rect 4967 1816 5113 1824
rect 5196 1824 5204 1836
rect 5427 1836 5453 1844
rect 5467 1836 5533 1844
rect 5196 1816 5333 1824
rect 5387 1816 5413 1824
rect 5587 1816 5653 1824
rect 447 1796 853 1804
rect 1267 1796 1293 1804
rect 1307 1796 1633 1804
rect 1867 1796 2033 1804
rect 2047 1796 2113 1804
rect 2256 1796 2353 1804
rect 607 1776 653 1784
rect 907 1776 993 1784
rect 1776 1776 2133 1784
rect 367 1756 433 1764
rect 1327 1756 1473 1764
rect 1776 1764 1784 1776
rect 2256 1784 2264 1796
rect 2827 1796 2953 1804
rect 3367 1796 3552 1804
rect 3587 1796 3653 1804
rect 3727 1796 3773 1804
rect 4547 1796 4713 1804
rect 4756 1796 4833 1804
rect 4756 1787 4764 1796
rect 5067 1796 5253 1804
rect 5307 1796 5533 1804
rect 2187 1776 2264 1784
rect 2287 1776 2613 1784
rect 2956 1776 3284 1784
rect 2956 1767 2964 1776
rect 1707 1756 1784 1764
rect 2347 1756 2373 1764
rect 2687 1756 2784 1764
rect 67 1737 173 1745
rect 496 1736 513 1744
rect 27 1695 73 1703
rect 256 1687 264 1734
rect 496 1707 504 1736
rect 567 1737 613 1745
rect 767 1736 813 1744
rect 840 1744 853 1747
rect 836 1733 853 1744
rect 1007 1736 1033 1744
rect 1047 1737 1073 1745
rect 1136 1736 1233 1744
rect 587 1696 673 1704
rect 735 1704 743 1733
rect 836 1706 844 1733
rect 1136 1706 1144 1736
rect 1256 1736 1293 1744
rect 1256 1706 1264 1736
rect 1607 1737 1673 1745
rect 1767 1737 1793 1745
rect 1947 1737 1993 1745
rect 2127 1737 2153 1745
rect 687 1696 743 1704
rect 907 1695 933 1703
rect 1436 1704 1444 1733
rect 1407 1696 1444 1704
rect 1507 1696 1573 1704
rect 2147 1696 2173 1704
rect 2256 1706 2264 1753
rect 2367 1744 2380 1747
rect 2367 1733 2384 1744
rect 2407 1736 2453 1744
rect 2527 1736 2544 1744
rect 2376 1724 2384 1733
rect 2536 1724 2544 1736
rect 2567 1736 2653 1744
rect 2707 1736 2753 1744
rect 2376 1716 2424 1724
rect 2536 1716 2604 1724
rect 2416 1706 2424 1716
rect 2596 1706 2604 1716
rect 2307 1696 2413 1704
rect 2776 1704 2784 1756
rect 2947 1756 2964 1767
rect 3276 1764 3284 1776
rect 3307 1776 3373 1784
rect 3427 1776 3673 1784
rect 3687 1776 3813 1784
rect 3827 1776 3853 1784
rect 4007 1776 4133 1784
rect 4487 1776 4753 1784
rect 5127 1776 5173 1784
rect 5627 1776 5773 1784
rect 3416 1764 3424 1773
rect 3276 1756 3424 1764
rect 3496 1756 3533 1764
rect 2947 1753 2960 1756
rect 2867 1737 2913 1745
rect 3087 1737 3113 1745
rect 3207 1737 3253 1745
rect 3496 1744 3504 1756
rect 3947 1756 3984 1764
rect 3476 1736 3504 1744
rect 3036 1724 3044 1734
rect 3036 1716 3064 1724
rect 2776 1696 2813 1704
rect 3056 1704 3064 1716
rect 3476 1707 3484 1736
rect 3687 1744 3700 1747
rect 3687 1733 3704 1744
rect 3056 1696 3093 1704
rect 3147 1695 3193 1703
rect 3327 1696 3393 1704
rect 3696 1706 3704 1733
rect 3736 1706 3744 1753
rect 3847 1736 3904 1744
rect 3787 1695 3813 1703
rect 3896 1704 3904 1736
rect 3976 1706 3984 1756
rect 4273 1764 4287 1773
rect 4127 1756 4204 1764
rect 4273 1760 4304 1764
rect 4276 1756 4304 1760
rect 4087 1737 4113 1745
rect 3896 1696 3964 1704
rect 727 1676 1133 1684
rect 1547 1676 1713 1684
rect 1727 1676 1813 1684
rect 1827 1676 1973 1684
rect 2387 1676 2653 1684
rect 2867 1676 2893 1684
rect 3007 1676 3493 1684
rect 3507 1676 3573 1684
rect 3587 1676 3673 1684
rect 3956 1684 3964 1696
rect 3996 1704 4004 1734
rect 4176 1707 4184 1733
rect 3996 1696 4093 1704
rect 4196 1706 4204 1756
rect 4227 1737 4273 1745
rect 3956 1676 4013 1684
rect 4296 1684 4304 1756
rect 4647 1756 4673 1764
rect 4727 1756 4804 1764
rect 4313 1744 4327 1753
rect 4313 1740 4353 1744
rect 4316 1736 4353 1740
rect 4376 1704 4384 1753
rect 4407 1736 4513 1744
rect 4456 1707 4464 1736
rect 4627 1736 4713 1744
rect 4796 1744 4804 1756
rect 4947 1756 5033 1764
rect 5396 1756 5433 1764
rect 4727 1736 4784 1744
rect 4796 1736 4824 1744
rect 4776 1724 4784 1736
rect 4776 1716 4804 1724
rect 4376 1696 4413 1704
rect 4547 1695 4633 1703
rect 4227 1676 4304 1684
rect 4796 1684 4804 1716
rect 4816 1707 4824 1736
rect 5056 1736 5153 1744
rect 5036 1724 5044 1733
rect 4916 1720 5044 1724
rect 4913 1716 5044 1720
rect 4913 1707 4927 1716
rect 5056 1704 5064 1736
rect 5227 1736 5293 1744
rect 5027 1696 5064 1704
rect 5187 1695 5213 1703
rect 5316 1704 5324 1753
rect 5396 1706 5404 1756
rect 5467 1736 5573 1744
rect 5647 1737 5673 1745
rect 5296 1696 5324 1704
rect 4707 1676 4853 1684
rect 5047 1676 5093 1684
rect 5296 1684 5304 1696
rect 5696 1704 5704 1753
rect 5716 1707 5724 1733
rect 5527 1696 5704 1704
rect 5207 1676 5304 1684
rect 5667 1676 5693 1684
rect 716 1664 724 1673
rect 547 1656 724 1664
rect 1227 1656 1313 1664
rect 1887 1656 1913 1664
rect 2007 1656 2053 1664
rect 2647 1656 2693 1664
rect 2747 1656 2933 1664
rect 3207 1656 3353 1664
rect 3727 1656 3913 1664
rect 4067 1656 4233 1664
rect 4307 1656 4453 1664
rect 4556 1656 5312 1664
rect 47 1636 73 1644
rect 167 1636 213 1644
rect 847 1636 1033 1644
rect 1347 1636 1413 1644
rect 2736 1644 2744 1653
rect 2367 1636 2744 1644
rect 2767 1636 2873 1644
rect 2947 1636 3113 1644
rect 3347 1636 3453 1644
rect 3947 1636 4373 1644
rect 4556 1644 4564 1656
rect 5347 1656 5493 1664
rect 4447 1636 4564 1644
rect 4587 1636 4893 1644
rect 5336 1644 5344 1653
rect 5147 1636 5344 1644
rect 5407 1636 5513 1644
rect 547 1616 613 1624
rect 987 1616 1093 1624
rect 1107 1616 1573 1624
rect 1687 1616 1893 1624
rect 2027 1616 2173 1624
rect 2827 1616 3284 1624
rect 3276 1607 3284 1616
rect 3707 1616 3833 1624
rect 4147 1616 4333 1624
rect 4507 1616 5093 1624
rect 1667 1596 2353 1604
rect 2707 1596 2804 1604
rect 767 1576 953 1584
rect 1127 1576 1593 1584
rect 1607 1576 1693 1584
rect 1987 1576 2073 1584
rect 2087 1576 2713 1584
rect 2796 1584 2804 1596
rect 2987 1596 3093 1604
rect 3287 1596 3853 1604
rect 4336 1604 4344 1613
rect 4336 1596 5433 1604
rect 2796 1576 2933 1584
rect 3127 1576 3593 1584
rect 3847 1576 3913 1584
rect 4267 1576 4333 1584
rect 4427 1576 4493 1584
rect 4507 1576 4593 1584
rect 4747 1576 5193 1584
rect 5247 1576 5353 1584
rect 5367 1576 5413 1584
rect 807 1556 1653 1564
rect 1867 1556 2104 1564
rect 1387 1536 1533 1544
rect 2096 1544 2104 1556
rect 2127 1556 2553 1564
rect 2827 1556 2953 1564
rect 3067 1564 3080 1567
rect 3067 1553 3084 1564
rect 3567 1556 4153 1564
rect 4167 1556 4393 1564
rect 4916 1556 5113 1564
rect 2096 1536 3033 1544
rect 3076 1544 3084 1553
rect 3076 1536 3573 1544
rect 3627 1536 3773 1544
rect 3847 1536 4173 1544
rect 4187 1536 4352 1544
rect 4387 1536 4553 1544
rect 4916 1544 4924 1556
rect 5567 1556 5793 1564
rect 4667 1536 4924 1544
rect 4967 1536 5533 1544
rect 607 1516 924 1524
rect 916 1507 924 1516
rect 1287 1516 1464 1524
rect 1456 1507 1464 1516
rect 2047 1516 2413 1524
rect 2727 1516 2853 1524
rect 2867 1516 3053 1524
rect 3127 1516 4033 1524
rect 4047 1516 4293 1524
rect 4427 1516 4613 1524
rect 4987 1516 5013 1524
rect 5136 1516 5493 1524
rect 87 1496 293 1504
rect 927 1496 1073 1504
rect 1467 1496 1773 1504
rect 1787 1496 2033 1504
rect 2687 1496 2793 1504
rect 2887 1496 2993 1504
rect 3387 1496 3553 1504
rect 4387 1496 4733 1504
rect 4827 1496 4993 1504
rect 5136 1504 5144 1516
rect 5007 1496 5144 1504
rect 5547 1496 5733 1504
rect 447 1476 473 1484
rect 767 1476 813 1484
rect 827 1476 1013 1484
rect 1167 1476 1313 1484
rect 1427 1476 1544 1484
rect 1536 1464 1544 1476
rect 1567 1476 1633 1484
rect 1696 1476 1793 1484
rect 1696 1464 1704 1476
rect 1807 1476 1913 1484
rect 1987 1476 2393 1484
rect 2947 1476 3012 1484
rect 3047 1476 3113 1484
rect 3167 1476 3293 1484
rect 3307 1476 3353 1484
rect 3687 1476 3873 1484
rect 4107 1476 4213 1484
rect 4487 1476 4633 1484
rect 4687 1476 4753 1484
rect 5027 1476 5124 1484
rect 1536 1456 1704 1464
rect 2147 1456 2193 1464
rect 2287 1456 2333 1464
rect 2647 1456 2773 1464
rect 2787 1456 2873 1464
rect 3587 1456 3653 1464
rect 127 1436 184 1444
rect 176 1407 184 1436
rect 227 1436 333 1444
rect 636 1407 644 1434
rect 716 1407 724 1434
rect 1487 1437 1513 1445
rect 1747 1437 1773 1445
rect 1827 1437 1853 1445
rect 836 1407 844 1433
rect 27 1396 93 1404
rect 407 1395 493 1403
rect 547 1396 573 1404
rect 636 1396 653 1407
rect 640 1393 653 1396
rect 707 1396 724 1407
rect 707 1393 720 1396
rect 876 1387 884 1434
rect 1236 1407 1244 1434
rect 1227 1396 1244 1407
rect 1256 1396 1393 1404
rect 1227 1393 1240 1396
rect 867 1376 884 1387
rect 867 1373 880 1376
rect 1007 1376 1093 1384
rect 1107 1376 1133 1384
rect 1256 1384 1264 1396
rect 1656 1404 1664 1434
rect 1547 1396 1664 1404
rect 1696 1404 1704 1434
rect 1936 1424 1944 1453
rect 2227 1436 2244 1444
rect 1896 1416 1944 1424
rect 1696 1396 1793 1404
rect 1896 1404 1904 1416
rect 1847 1396 1904 1404
rect 2076 1404 2084 1434
rect 2027 1396 2084 1404
rect 2236 1404 2244 1436
rect 2296 1404 2304 1433
rect 2436 1407 2444 1433
rect 2236 1396 2264 1404
rect 2296 1396 2333 1404
rect 1207 1376 1264 1384
rect 1347 1376 1373 1384
rect 1927 1376 1993 1384
rect 2256 1384 2264 1396
rect 2496 1406 2504 1453
rect 4347 1456 4544 1464
rect 2567 1437 2593 1445
rect 2516 1407 2524 1434
rect 3036 1436 3092 1444
rect 2516 1396 2533 1407
rect 2520 1393 2533 1396
rect 2676 1404 2684 1433
rect 2793 1424 2807 1433
rect 2896 1424 2904 1434
rect 2793 1420 2904 1424
rect 2796 1416 2904 1420
rect 2667 1396 2684 1404
rect 2833 1407 2847 1416
rect 2976 1404 2984 1434
rect 3036 1406 3044 1436
rect 3116 1407 3124 1434
rect 3447 1436 3513 1444
rect 4187 1437 4232 1445
rect 2887 1396 2984 1404
rect 3107 1396 3124 1407
rect 3107 1393 3120 1396
rect 3235 1387 3243 1433
rect 3256 1424 3264 1434
rect 3696 1424 3704 1434
rect 4367 1436 4413 1444
rect 4427 1436 4513 1444
rect 3256 1416 3284 1424
rect 3696 1416 3724 1424
rect 3276 1404 3284 1416
rect 3276 1396 3313 1404
rect 3367 1395 3413 1403
rect 3487 1395 3533 1403
rect 3607 1395 3653 1403
rect 3716 1404 3724 1416
rect 4253 1424 4267 1433
rect 4416 1424 4424 1434
rect 3747 1420 4267 1424
rect 4396 1420 4424 1424
rect 3747 1416 4264 1420
rect 4393 1416 4424 1420
rect 4393 1407 4407 1416
rect 3716 1396 3793 1404
rect 3887 1395 3933 1403
rect 4167 1396 4273 1404
rect 4536 1404 4544 1456
rect 4627 1456 4713 1464
rect 5116 1464 5124 1476
rect 5167 1476 5472 1484
rect 5507 1476 5884 1484
rect 5007 1456 5084 1464
rect 5116 1456 5184 1464
rect 4576 1407 4584 1434
rect 4907 1437 4953 1445
rect 5076 1444 5084 1456
rect 5076 1436 5164 1444
rect 4636 1407 4644 1433
rect 4736 1407 4744 1433
rect 4447 1396 4564 1404
rect 4576 1396 4593 1407
rect 2256 1376 2564 1384
rect 3235 1376 3253 1387
rect 2556 1367 2564 1376
rect 3240 1373 3253 1376
rect 3967 1376 4013 1384
rect 4027 1376 4113 1384
rect 4167 1376 4213 1384
rect 4556 1384 4564 1396
rect 4580 1393 4593 1396
rect 4807 1396 4993 1404
rect 4796 1384 4804 1392
rect 5156 1387 5164 1436
rect 5176 1406 5184 1456
rect 5407 1456 5764 1464
rect 5207 1436 5293 1444
rect 5447 1436 5573 1444
rect 5756 1444 5764 1456
rect 5756 1436 5773 1444
rect 5387 1395 5453 1403
rect 5467 1396 5593 1404
rect 5656 1387 5664 1434
rect 5876 1436 5884 1476
rect 5707 1395 5753 1403
rect 5816 1404 5824 1433
rect 5807 1396 5824 1404
rect 4556 1376 4804 1384
rect 5147 1384 5164 1387
rect 5147 1376 5313 1384
rect 5147 1373 5160 1376
rect 47 1356 93 1364
rect 707 1356 933 1364
rect 1087 1356 1253 1364
rect 1827 1356 1873 1364
rect 1967 1356 2473 1364
rect 2567 1356 2753 1364
rect 3147 1356 3213 1364
rect 3427 1356 3613 1364
rect 4287 1356 4373 1364
rect 4607 1356 4784 1364
rect 167 1336 233 1344
rect 1287 1336 1313 1344
rect 1327 1336 1433 1344
rect 1447 1336 1893 1344
rect 2147 1336 2233 1344
rect 2547 1336 2613 1344
rect 2767 1336 2793 1344
rect 3027 1336 3073 1344
rect 3347 1336 3513 1344
rect 3796 1336 4113 1344
rect 3796 1327 3804 1336
rect 4267 1336 4453 1344
rect 4567 1336 4653 1344
rect 4776 1344 4784 1356
rect 5047 1356 5073 1364
rect 5267 1356 5373 1364
rect 5447 1356 5513 1364
rect 4776 1336 4812 1344
rect 4847 1336 5113 1344
rect 5287 1336 5313 1344
rect 667 1316 853 1324
rect 947 1316 1533 1324
rect 1687 1316 2053 1324
rect 2107 1316 2233 1324
rect 2427 1316 2513 1324
rect 3287 1316 3433 1324
rect 3587 1316 3633 1324
rect 3687 1316 3793 1324
rect 3907 1316 4133 1324
rect 4247 1316 4293 1324
rect 4307 1316 4493 1324
rect 4507 1316 4533 1324
rect 5107 1316 5493 1324
rect 5507 1316 5633 1324
rect 5647 1316 5673 1324
rect 27 1296 193 1304
rect 687 1296 733 1304
rect 1047 1296 1193 1304
rect 1567 1296 1593 1304
rect 1767 1296 1953 1304
rect 2127 1296 2353 1304
rect 2407 1296 2493 1304
rect 2576 1296 2793 1304
rect 627 1276 813 1284
rect 827 1276 893 1284
rect 1227 1276 1733 1284
rect 2427 1276 2453 1284
rect 2576 1284 2584 1296
rect 3007 1296 3073 1304
rect 3087 1296 3173 1304
rect 3187 1296 3313 1304
rect 3467 1296 3613 1304
rect 3716 1296 3824 1304
rect 2527 1276 2584 1284
rect 2596 1276 2672 1284
rect 547 1256 773 1264
rect 1487 1256 1673 1264
rect 2127 1256 2193 1264
rect 2307 1256 2333 1264
rect 2596 1264 2604 1276
rect 2707 1276 2864 1284
rect 2487 1256 2604 1264
rect 2627 1256 2813 1264
rect 2856 1264 2864 1276
rect 2987 1276 3093 1284
rect 3716 1284 3724 1296
rect 3676 1276 3724 1284
rect 3816 1284 3824 1296
rect 3887 1296 4104 1304
rect 3816 1276 3952 1284
rect 2856 1256 3033 1264
rect 3127 1256 3333 1264
rect 3676 1264 3684 1276
rect 4096 1284 4104 1296
rect 4267 1296 4473 1304
rect 5547 1296 5613 1304
rect 5727 1296 5753 1304
rect 3987 1276 4084 1284
rect 4096 1276 4193 1284
rect 3387 1256 3684 1264
rect 3807 1256 3993 1264
rect 4076 1264 4084 1276
rect 4327 1276 4613 1284
rect 5527 1276 5633 1284
rect 5647 1276 5813 1284
rect 4076 1256 4133 1264
rect 4580 1264 4593 1267
rect 4576 1253 4593 1264
rect 4647 1256 4673 1264
rect 4867 1256 4953 1264
rect 4967 1256 5013 1264
rect 5147 1256 5333 1264
rect 5496 1256 5553 1264
rect 47 1236 133 1244
rect 607 1236 653 1244
rect 1047 1236 1073 1244
rect 1207 1236 1253 1244
rect 2067 1236 2093 1244
rect 2367 1236 2693 1244
rect 2847 1236 3473 1244
rect 3733 1244 3747 1253
rect 3627 1240 3747 1244
rect 3627 1236 3744 1240
rect 4127 1236 4493 1244
rect 4576 1244 4584 1253
rect 5496 1247 5504 1256
rect 5676 1256 5733 1264
rect 4507 1236 4584 1244
rect 5127 1236 5213 1244
rect 5487 1236 5504 1247
rect 5487 1233 5500 1236
rect 5627 1236 5653 1244
rect 187 1216 264 1224
rect 256 1204 264 1216
rect 287 1216 373 1224
rect 427 1217 453 1225
rect 507 1217 533 1225
rect 747 1216 773 1224
rect 1167 1216 1273 1224
rect 1316 1216 1353 1224
rect 256 1196 304 1204
rect 296 1186 304 1196
rect 47 1175 73 1183
rect 127 1176 173 1184
rect 187 1175 213 1183
rect 616 1184 624 1213
rect 567 1176 624 1184
rect 856 1184 864 1213
rect 847 1176 913 1184
rect 1127 1176 1253 1184
rect 1316 1184 1324 1216
rect 1407 1216 1473 1224
rect 1607 1217 1653 1225
rect 2147 1217 2193 1225
rect 2287 1217 2333 1225
rect 2867 1217 2933 1225
rect 2987 1216 3153 1224
rect 3207 1216 3273 1224
rect 1553 1204 1567 1213
rect 1553 1200 1584 1204
rect 1556 1196 1584 1200
rect 1576 1186 1584 1196
rect 1316 1176 1333 1184
rect 1707 1175 1853 1183
rect 2236 1184 2244 1213
rect 2316 1196 2873 1204
rect 2316 1186 2324 1196
rect 2227 1176 2244 1184
rect 2967 1175 2993 1183
rect 3056 1180 3113 1184
rect 3053 1176 3113 1180
rect 3053 1167 3067 1176
rect 3287 1175 3313 1183
rect 3336 1184 3344 1214
rect 3527 1216 3633 1224
rect 3647 1216 3873 1224
rect 3336 1176 3393 1184
rect 347 1156 433 1164
rect 1387 1156 1433 1164
rect 1847 1156 2633 1164
rect 2707 1156 3044 1164
rect 1087 1136 1313 1144
rect 1327 1136 1453 1144
rect 1507 1136 1633 1144
rect 1647 1136 2173 1144
rect 2227 1136 2353 1144
rect 3036 1144 3044 1156
rect 3066 1160 3067 1167
rect 3087 1156 3133 1164
rect 3455 1164 3463 1213
rect 3476 1167 3484 1213
rect 3776 1186 3784 1216
rect 3947 1216 4053 1224
rect 4076 1216 4093 1224
rect 4076 1204 4084 1216
rect 4347 1216 4364 1224
rect 4056 1196 4084 1204
rect 3547 1176 3613 1184
rect 3627 1175 3733 1183
rect 3887 1175 3953 1183
rect 4056 1167 4064 1196
rect 4356 1187 4364 1216
rect 4733 1224 4747 1233
rect 4647 1216 4724 1224
rect 4733 1220 4752 1224
rect 4736 1216 4752 1220
rect 4596 1187 4604 1214
rect 4716 1187 4724 1216
rect 4947 1216 4973 1224
rect 5216 1224 5224 1233
rect 5156 1216 5224 1224
rect 4187 1176 4313 1184
rect 4356 1176 4373 1187
rect 4360 1173 4373 1176
rect 4447 1175 4552 1183
rect 4587 1176 4604 1187
rect 4587 1173 4600 1176
rect 4776 1184 4784 1213
rect 4813 1204 4827 1213
rect 4813 1200 4884 1204
rect 4816 1196 4884 1200
rect 4776 1176 4813 1184
rect 4876 1186 4884 1196
rect 5096 1184 5104 1214
rect 5156 1186 5164 1216
rect 5007 1176 5104 1184
rect 5276 1184 5284 1214
rect 5347 1224 5360 1227
rect 5347 1213 5364 1224
rect 5356 1186 5364 1213
rect 5416 1187 5424 1214
rect 5676 1207 5684 1256
rect 5767 1236 5844 1244
rect 5227 1176 5284 1184
rect 5416 1176 5433 1187
rect 5420 1173 5433 1176
rect 3347 1156 3463 1164
rect 4207 1156 4253 1164
rect 5836 1147 5844 1236
rect 3036 1136 3113 1144
rect 3287 1136 3493 1144
rect 3627 1136 3833 1144
rect 4387 1136 4653 1144
rect 4727 1136 5213 1144
rect 5267 1136 5433 1144
rect 267 1116 453 1124
rect 507 1116 673 1124
rect 687 1116 1293 1124
rect 1587 1116 1653 1124
rect 1907 1116 2133 1124
rect 2207 1116 2233 1124
rect 2367 1116 2593 1124
rect 2776 1116 2893 1124
rect 647 1096 1193 1104
rect 1427 1096 1493 1104
rect 2776 1104 2784 1116
rect 2967 1116 3264 1124
rect 2327 1096 2784 1104
rect 2927 1096 3013 1104
rect 3256 1104 3264 1116
rect 3967 1116 4353 1124
rect 4407 1116 4513 1124
rect 4567 1116 4833 1124
rect 5467 1116 5793 1124
rect 3256 1096 3364 1104
rect 3356 1087 3364 1096
rect 3807 1096 3853 1104
rect 3876 1096 4293 1104
rect 2027 1076 2073 1084
rect 2347 1076 2833 1084
rect 2887 1076 2933 1084
rect 3067 1076 3173 1084
rect 3187 1076 3332 1084
rect 3367 1076 3613 1084
rect 3876 1084 3884 1096
rect 4487 1096 4613 1104
rect 4747 1096 4793 1104
rect 5327 1096 5593 1104
rect 3767 1076 3884 1084
rect 3987 1076 4273 1084
rect 4907 1076 5153 1084
rect 5267 1076 5353 1084
rect 1407 1056 1512 1064
rect 1547 1056 1713 1064
rect 2327 1056 2473 1064
rect 2527 1056 2733 1064
rect 2867 1056 3033 1064
rect 3407 1056 3693 1064
rect 3747 1056 3813 1064
rect 3867 1056 3993 1064
rect 4007 1056 4224 1064
rect 1507 1036 2073 1044
rect 2247 1036 2353 1044
rect 2507 1036 3033 1044
rect 3127 1036 3232 1044
rect 3267 1036 3353 1044
rect 4027 1036 4193 1044
rect 4216 1044 4224 1056
rect 4487 1056 4573 1064
rect 5187 1056 5393 1064
rect 5407 1056 5673 1064
rect 4216 1036 4784 1044
rect 427 1016 2112 1024
rect 2147 1016 2332 1024
rect 2367 1016 2452 1024
rect 2487 1016 2693 1024
rect 2747 1016 2953 1024
rect 3027 1016 3153 1024
rect 3167 1016 3293 1024
rect 3707 1016 3893 1024
rect 3907 1016 3973 1024
rect 4087 1016 4473 1024
rect 4587 1016 4613 1024
rect 4776 1024 4784 1036
rect 4927 1036 5184 1044
rect 4776 1016 4933 1024
rect 5176 1024 5184 1036
rect 5207 1036 5353 1044
rect 5447 1036 5633 1044
rect 5176 1016 5613 1024
rect 647 996 733 1004
rect 1287 996 1684 1004
rect 1676 987 1684 996
rect 2187 996 2333 1004
rect 2847 996 2993 1004
rect 3047 996 3253 1004
rect 3447 996 3773 1004
rect 4227 996 4393 1004
rect 4527 996 4753 1004
rect 4767 996 4993 1004
rect 5067 996 5233 1004
rect 1267 976 1473 984
rect 1687 976 1853 984
rect 1947 976 2413 984
rect 2467 976 2713 984
rect 2727 976 2813 984
rect 2827 976 3053 984
rect 3107 976 3213 984
rect 3347 976 3933 984
rect 5387 976 5493 984
rect 5667 976 5753 984
rect 527 956 693 964
rect 887 956 973 964
rect 1727 956 2033 964
rect 2107 956 2393 964
rect 2507 953 2513 967
rect 2927 956 3193 964
rect 3207 956 3393 964
rect 3667 956 3733 964
rect 3776 956 3873 964
rect 167 936 253 944
rect 607 936 633 944
rect 2587 936 2613 944
rect 2727 936 2753 944
rect 3007 936 3184 944
rect 327 917 373 925
rect 396 916 412 924
rect 27 876 73 884
rect 96 864 104 914
rect 256 884 264 914
rect 396 904 404 916
rect 567 916 653 924
rect 707 917 733 925
rect 947 916 1093 924
rect 376 896 404 904
rect 256 876 333 884
rect 376 867 384 896
rect 436 884 444 913
rect 407 876 444 884
rect 547 876 673 884
rect 796 884 804 914
rect 767 876 804 884
rect 836 884 844 914
rect 836 876 893 884
rect 967 875 1013 883
rect 1096 884 1104 913
rect 1136 904 1144 914
rect 1136 896 1293 904
rect 1396 887 1404 914
rect 1567 916 1593 924
rect 2027 916 2133 924
rect 1733 904 1747 913
rect 1976 904 1984 914
rect 1733 900 1984 904
rect 1736 896 1984 900
rect 1096 876 1144 884
rect 1396 876 1413 887
rect 96 856 133 864
rect 227 856 373 864
rect 427 856 453 864
rect 567 856 593 864
rect 1016 864 1024 872
rect 1016 856 1113 864
rect 1136 864 1144 876
rect 1400 873 1413 876
rect 1527 876 1593 884
rect 1607 875 1653 883
rect 1856 867 1864 896
rect 1947 875 1993 883
rect 1136 856 1233 864
rect 1367 856 1473 864
rect 2156 864 2164 933
rect 2176 916 2233 924
rect 2176 887 2184 916
rect 2253 924 2267 933
rect 2253 920 2324 924
rect 2256 916 2324 920
rect 2127 856 2164 864
rect 2316 864 2324 916
rect 2347 916 2393 924
rect 2396 904 2404 914
rect 2336 900 2433 904
rect 2333 896 2433 900
rect 2333 887 2347 896
rect 2476 884 2484 914
rect 2567 916 2693 924
rect 2927 917 2973 925
rect 3176 904 3184 936
rect 3227 944 3240 947
rect 3227 933 3244 944
rect 3776 944 3784 956
rect 3967 956 4213 964
rect 4707 956 5053 964
rect 5067 956 5313 964
rect 5687 956 5713 964
rect 3427 936 3784 944
rect 3176 900 3204 904
rect 3176 896 3207 900
rect 3193 887 3207 896
rect 3236 887 3244 933
rect 3487 916 3504 924
rect 3336 887 3344 914
rect 2387 876 2484 884
rect 2547 875 2573 883
rect 2687 876 2773 884
rect 3047 876 3172 884
rect 3336 876 3353 887
rect 3340 873 3353 876
rect 3436 867 3444 914
rect 3496 884 3504 916
rect 3547 917 3573 925
rect 3616 887 3624 914
rect 3696 887 3704 914
rect 3496 876 3593 884
rect 3616 876 3633 887
rect 3620 873 3633 876
rect 3687 876 3704 887
rect 3687 873 3700 876
rect 2316 856 2353 864
rect 2447 856 2493 864
rect 2607 856 2753 864
rect 2767 856 2853 864
rect 3756 864 3764 936
rect 4347 936 4613 944
rect 5487 936 5573 944
rect 3827 916 3953 924
rect 3776 887 3784 913
rect 4016 904 4024 914
rect 4127 916 4213 924
rect 4227 916 4333 924
rect 4456 916 4633 924
rect 3976 896 4024 904
rect 3976 887 3984 896
rect 3887 875 3932 883
rect 3967 876 3984 887
rect 3967 873 3980 876
rect 4076 884 4084 913
rect 4456 904 4464 916
rect 4647 916 4664 924
rect 4376 896 4464 904
rect 4007 876 4093 884
rect 4247 876 4353 884
rect 4376 884 4384 896
rect 4367 876 4384 884
rect 4547 876 4573 884
rect 4587 875 4613 883
rect 4656 884 4664 916
rect 4687 917 4713 925
rect 4847 917 4873 925
rect 4987 924 5000 927
rect 4987 913 5004 924
rect 5027 917 5093 925
rect 5327 916 5444 924
rect 4656 876 4733 884
rect 4787 876 4833 884
rect 4996 886 5004 913
rect 5136 884 5144 914
rect 5047 876 5144 884
rect 5276 884 5284 914
rect 5436 886 5444 916
rect 5507 917 5533 925
rect 5647 924 5660 927
rect 5647 913 5664 924
rect 5596 887 5604 913
rect 5276 876 5393 884
rect 5656 886 5664 913
rect 3707 856 3764 864
rect 3796 856 3833 864
rect 687 836 913 844
rect 1447 836 1533 844
rect 1587 836 1773 844
rect 2267 836 2333 844
rect 2667 836 2793 844
rect 3107 836 3133 844
rect 3187 836 3413 844
rect 3527 836 3593 844
rect 3796 844 3804 856
rect 4447 856 4493 864
rect 4907 856 4973 864
rect 5027 856 5153 864
rect 3667 836 3804 844
rect 3867 836 3953 844
rect 4847 836 5393 844
rect 5607 836 5673 844
rect 167 816 333 824
rect 347 816 593 824
rect 707 816 853 824
rect 1347 816 1404 824
rect 187 796 233 804
rect 247 796 273 804
rect 287 796 493 804
rect 747 796 813 804
rect 1396 804 1404 816
rect 1427 816 1513 824
rect 2207 816 2293 824
rect 2416 816 2812 824
rect 907 796 1184 804
rect 1396 796 1573 804
rect 1176 787 1184 796
rect 1707 796 1833 804
rect 2047 796 2133 804
rect 2416 804 2424 816
rect 2847 816 2993 824
rect 3447 816 3633 824
rect 3647 816 3753 824
rect 3767 816 3813 824
rect 4307 816 4404 824
rect 2227 796 2424 804
rect 2527 796 2933 804
rect 2947 796 3133 804
rect 3287 796 3613 804
rect 3887 796 4153 804
rect 4396 804 4404 816
rect 5167 816 5233 824
rect 4396 796 4573 804
rect 4647 796 4813 804
rect 5307 796 5373 804
rect 5387 796 5553 804
rect 5647 796 5693 804
rect 127 776 193 784
rect 987 776 1104 784
rect 1096 767 1104 776
rect 1187 776 1293 784
rect 1307 776 1373 784
rect 1807 776 1873 784
rect 1887 776 1953 784
rect 3207 776 3473 784
rect 3587 776 3693 784
rect 5407 776 5493 784
rect 5587 776 5613 784
rect 367 756 393 764
rect 407 756 633 764
rect 847 756 873 764
rect 896 756 1072 764
rect 87 736 213 744
rect 767 736 813 744
rect 896 744 904 756
rect 1107 756 1153 764
rect 1427 756 1473 764
rect 1687 756 1713 764
rect 1787 756 1873 764
rect 1987 756 2153 764
rect 2167 756 2373 764
rect 2427 756 2493 764
rect 2587 756 2693 764
rect 2747 756 2793 764
rect 2807 756 2864 764
rect 867 736 904 744
rect 1067 736 1133 744
rect 1247 736 1313 744
rect 1407 736 1573 744
rect 1627 736 1753 744
rect 1767 736 1933 744
rect 2616 736 2833 744
rect 216 716 313 724
rect 167 704 180 707
rect 167 693 184 704
rect 107 656 133 664
rect 176 666 184 693
rect 216 666 224 716
rect 367 716 453 724
rect 507 716 693 724
rect 1027 716 1064 724
rect 247 696 264 704
rect 256 667 264 696
rect 347 696 404 704
rect 396 664 404 696
rect 647 697 673 705
rect 727 696 753 704
rect 956 696 1033 704
rect 796 684 804 694
rect 796 676 933 684
rect 956 667 964 696
rect 396 656 533 664
rect 667 655 693 663
rect 1056 664 1064 716
rect 1296 716 1333 724
rect 1227 696 1273 704
rect 1296 666 1304 716
rect 1496 716 1773 724
rect 1327 697 1352 705
rect 1387 697 1433 705
rect 1356 684 1364 694
rect 1356 676 1444 684
rect 1056 656 1113 664
rect 1167 655 1233 663
rect 1436 664 1444 676
rect 1496 666 1504 716
rect 2067 716 2173 724
rect 2196 716 2233 724
rect 1780 704 1793 707
rect 1596 696 1793 704
rect 1596 666 1604 696
rect 1776 693 1793 696
rect 1856 696 1913 704
rect 1776 666 1784 693
rect 1856 667 1864 696
rect 2196 704 2204 716
rect 2107 696 2204 704
rect 2467 696 2573 704
rect 1436 656 1453 664
rect 1647 656 1733 664
rect 1956 664 1964 693
rect 1947 656 1964 664
rect 1987 655 2033 663
rect 2256 664 2264 693
rect 2247 656 2264 664
rect 2316 664 2324 693
rect 2316 656 2493 664
rect 2616 664 2624 736
rect 2856 744 2864 756
rect 2927 756 2993 764
rect 3127 756 3273 764
rect 3327 756 3372 764
rect 3407 756 3553 764
rect 3607 756 3633 764
rect 3727 756 4013 764
rect 4027 756 4273 764
rect 4547 756 4853 764
rect 5100 764 5112 767
rect 4927 756 5112 764
rect 5096 753 5112 756
rect 5147 756 5193 764
rect 5367 756 5513 764
rect 2856 736 2973 744
rect 3027 736 3273 744
rect 2660 704 2673 707
rect 2607 656 2624 664
rect 2656 693 2673 704
rect 2656 667 2664 693
rect 2656 656 2673 667
rect 2660 653 2673 656
rect 567 636 613 644
rect 747 636 833 644
rect 847 636 873 644
rect 1067 636 1093 644
rect 1976 644 1984 652
rect 2716 647 2724 713
rect 2776 696 2813 704
rect 2776 667 2784 696
rect 2867 697 2933 705
rect 2807 684 2820 687
rect 2807 673 2824 684
rect 2816 664 2824 673
rect 2816 656 2833 664
rect 2887 655 2913 663
rect 2996 664 3004 694
rect 3016 666 3024 733
rect 3396 736 3693 744
rect 3296 716 3353 724
rect 3047 696 3164 704
rect 3156 684 3164 696
rect 3187 696 3264 704
rect 3156 676 3204 684
rect 3196 666 3204 676
rect 3256 667 3264 696
rect 2927 656 3004 664
rect 3296 666 3304 716
rect 3396 724 3404 736
rect 3807 736 3993 744
rect 4067 736 4153 744
rect 4167 736 5073 744
rect 5096 744 5104 753
rect 5096 736 5293 744
rect 3367 716 3404 724
rect 3427 716 3453 724
rect 4687 716 4713 724
rect 5107 716 5173 724
rect 5187 716 5273 724
rect 5347 716 5412 724
rect 5507 716 5593 724
rect 3327 696 3533 704
rect 3416 666 3424 696
rect 3576 684 3584 694
rect 3840 704 3853 707
rect 3627 696 3853 704
rect 3836 693 3853 696
rect 4127 696 4193 704
rect 3576 676 3724 684
rect 3716 666 3724 676
rect 3836 666 3844 693
rect 3936 684 3944 694
rect 4076 684 4084 694
rect 4236 684 4244 694
rect 4287 696 4364 704
rect 3936 680 3984 684
rect 3936 676 3987 680
rect 4076 676 4124 684
rect 4236 680 4324 684
rect 4236 676 4327 680
rect 3973 667 3987 676
rect 3607 656 3673 664
rect 3887 655 3913 663
rect 4116 667 4124 676
rect 4313 667 4327 676
rect 4027 655 4053 663
rect 4116 656 4133 667
rect 4120 653 4133 656
rect 4356 666 4364 696
rect 4453 704 4467 713
rect 4387 696 4493 704
rect 4687 696 4753 704
rect 4807 696 4913 704
rect 4967 696 4993 704
rect 5016 696 5053 704
rect 5016 684 5024 696
rect 5227 696 5284 704
rect 4936 676 5024 684
rect 5276 684 5284 696
rect 5307 696 5393 704
rect 5433 704 5447 713
rect 5433 700 5473 704
rect 5436 696 5473 700
rect 5527 696 5544 704
rect 5393 684 5407 693
rect 5276 676 5384 684
rect 5393 680 5484 684
rect 5396 676 5484 680
rect 4936 666 4944 676
rect 4407 655 4433 663
rect 4447 656 4513 664
rect 4827 656 4933 664
rect 5087 656 5133 664
rect 5147 655 5193 663
rect 5376 664 5384 676
rect 5376 656 5433 664
rect 5476 647 5484 676
rect 5536 664 5544 696
rect 5647 696 5684 704
rect 5676 667 5684 696
rect 5536 656 5644 664
rect 5636 647 5644 656
rect 5747 656 5793 664
rect 1756 636 1984 644
rect 1756 627 1764 636
rect 2167 640 2224 644
rect 2167 636 2227 640
rect 2213 627 2227 636
rect 2707 636 2724 647
rect 2707 633 2720 636
rect 2967 636 3053 644
rect 3347 636 3373 644
rect 3387 636 3513 644
rect 5287 636 5373 644
rect 5636 636 5653 647
rect 5640 633 5653 636
rect 527 616 673 624
rect 947 616 1153 624
rect 1507 616 1724 624
rect 787 596 813 604
rect 827 596 993 604
rect 1207 596 1673 604
rect 1716 604 1724 616
rect 1747 616 1764 627
rect 1747 613 1760 616
rect 1907 616 2173 624
rect 2287 616 2373 624
rect 2427 616 2453 624
rect 2767 616 2933 624
rect 2947 616 2973 624
rect 2987 616 3353 624
rect 3407 616 3453 624
rect 4667 616 4913 624
rect 5467 616 5533 624
rect 5587 616 5693 624
rect 1716 596 1813 604
rect 1887 596 2373 604
rect 2447 596 2513 604
rect 2527 596 2553 604
rect 3027 596 3153 604
rect 3487 596 3593 604
rect 4007 596 4753 604
rect 4867 596 5253 604
rect 5387 596 5493 604
rect 1287 576 1653 584
rect 1727 576 1793 584
rect 1867 576 2393 584
rect 2467 576 3013 584
rect 3547 576 3633 584
rect 3987 576 4773 584
rect 4787 576 4893 584
rect 4907 576 5713 584
rect 427 556 1053 564
rect 1067 556 1492 564
rect 1527 556 1873 564
rect 2147 556 2373 564
rect 2447 556 3033 564
rect 3567 556 4253 564
rect 4267 556 4373 564
rect 4507 556 4573 564
rect 4927 556 5293 564
rect 1127 536 1733 544
rect 2307 536 2413 544
rect 2507 536 2553 544
rect 4627 536 4953 544
rect 1347 516 1953 524
rect 2407 516 2913 524
rect 3247 516 3433 524
rect 4307 516 5213 524
rect 267 496 413 504
rect 427 496 513 504
rect 1027 496 1593 504
rect 1687 496 1893 504
rect 2167 496 2353 504
rect 2467 496 2713 504
rect 2727 496 2953 504
rect 3027 496 3113 504
rect 3227 496 3793 504
rect 167 476 193 484
rect 207 476 773 484
rect 867 476 984 484
rect 976 467 984 476
rect 1627 476 2113 484
rect 2207 476 2313 484
rect 2387 476 2493 484
rect 2507 476 2533 484
rect 2727 476 2773 484
rect 2827 476 2993 484
rect 3267 476 4093 484
rect 4147 476 4553 484
rect 987 456 1193 464
rect 1827 456 2013 464
rect 2247 456 2333 464
rect 2347 456 2973 464
rect 3847 456 3893 464
rect 5247 456 5613 464
rect 5627 456 5633 464
rect 227 436 333 444
rect 787 436 953 444
rect 1147 436 1273 444
rect 1607 436 1853 444
rect 2407 436 2453 444
rect 2547 436 2573 444
rect 2587 436 2633 444
rect 2687 436 2793 444
rect 3067 436 3213 444
rect 3987 436 4053 444
rect 4127 436 4293 444
rect 4307 436 4353 444
rect 4647 436 4713 444
rect 4727 436 4813 444
rect 5327 436 5553 444
rect 547 416 633 424
rect 647 416 673 424
rect 1107 416 1333 424
rect 1347 416 1373 424
rect 1387 416 1553 424
rect 2787 416 2953 424
rect 3167 416 3193 424
rect 3207 416 3253 424
rect 3307 416 3573 424
rect 5767 416 5813 424
rect 47 356 93 364
rect 116 347 124 394
rect 467 397 493 405
rect 176 364 184 393
rect 176 356 233 364
rect 296 364 304 394
rect 576 384 584 394
rect 716 384 724 394
rect 576 376 724 384
rect 256 360 304 364
rect 253 356 304 360
rect 253 347 267 356
rect 347 356 393 364
rect 716 364 724 376
rect 716 356 753 364
rect 856 366 864 413
rect 876 364 884 394
rect 907 396 1013 404
rect 1160 404 1173 407
rect 876 356 993 364
rect 327 336 553 344
rect 1016 344 1024 394
rect 1156 393 1173 404
rect 1427 396 1473 404
rect 1487 396 1513 404
rect 1727 396 1804 404
rect 1156 366 1164 393
rect 1167 356 1293 364
rect 1356 364 1364 393
rect 1796 384 1804 396
rect 1827 396 1933 404
rect 2087 396 2193 404
rect 2216 396 2272 404
rect 2216 384 2224 396
rect 2307 397 2333 405
rect 1436 376 1804 384
rect 2176 380 2224 384
rect 1436 366 1444 376
rect 1796 366 1804 376
rect 2173 376 2224 380
rect 2173 367 2187 376
rect 1356 356 1393 364
rect 1867 355 1913 363
rect 2107 355 2152 363
rect 2356 366 2364 413
rect 2687 396 2813 404
rect 2416 367 2424 393
rect 2556 364 2564 393
rect 2736 367 2744 396
rect 2867 397 2913 405
rect 2556 356 2593 364
rect 2956 364 2964 394
rect 2956 356 3012 364
rect 3036 366 3044 413
rect 3107 396 3133 404
rect 3367 396 3473 404
rect 3667 397 3713 405
rect 3767 396 3793 404
rect 3616 367 3624 394
rect 3867 396 3913 404
rect 3087 355 3153 363
rect 3247 356 3453 364
rect 3547 356 3593 364
rect 3616 356 3633 367
rect 3620 353 3633 356
rect 3807 355 3833 363
rect 3927 355 3953 363
rect 4016 364 4024 394
rect 4156 384 4164 394
rect 4256 384 4264 394
rect 4387 396 4424 404
rect 4156 376 4264 384
rect 4016 356 4233 364
rect 4256 364 4264 376
rect 4256 356 4313 364
rect 4416 366 4424 396
rect 4607 396 4713 404
rect 4767 397 4853 405
rect 4907 397 5053 405
rect 5107 397 5133 405
rect 4716 384 4724 394
rect 4716 376 5204 384
rect 4527 355 4573 363
rect 4587 356 4693 364
rect 4716 364 4724 376
rect 4716 356 4833 364
rect 5196 366 5204 376
rect 5236 366 5244 413
rect 5267 396 5284 404
rect 5276 367 5284 396
rect 5316 367 5324 393
rect 4907 356 4933 364
rect 5007 355 5073 363
rect 5356 364 5364 394
rect 5396 384 5404 394
rect 5396 376 5444 384
rect 5436 367 5444 376
rect 5356 356 5413 364
rect 5436 356 5453 367
rect 5440 353 5453 356
rect 5516 364 5524 394
rect 5656 366 5664 413
rect 5516 356 5613 364
rect 607 336 744 344
rect 1016 336 1253 344
rect 736 327 744 336
rect 1987 336 2053 344
rect 2156 344 2164 352
rect 2156 336 2213 344
rect 2296 336 2464 344
rect 2296 327 2304 336
rect 227 316 273 324
rect 367 316 413 324
rect 627 316 693 324
rect 747 316 953 324
rect 1187 316 1413 324
rect 1507 316 1613 324
rect 1627 316 1653 324
rect 1707 316 2293 324
rect 2407 316 2433 324
rect 2456 324 2464 336
rect 2487 336 2613 344
rect 2687 336 2713 344
rect 3156 344 3164 352
rect 5676 347 5684 394
rect 3156 336 3333 344
rect 4507 336 5113 344
rect 5307 336 5333 344
rect 2456 316 2793 324
rect 2807 316 2853 324
rect 3187 316 3233 324
rect 4147 316 4273 324
rect 4287 316 4353 324
rect 4367 316 4533 324
rect 5027 316 5173 324
rect 5507 316 5573 324
rect 5787 316 5833 324
rect 127 296 313 304
rect 447 296 473 304
rect 487 296 593 304
rect 607 296 813 304
rect 1007 296 1433 304
rect 1807 296 1833 304
rect 2027 296 2133 304
rect 2327 296 2473 304
rect 2547 296 2573 304
rect 2747 296 2933 304
rect 3827 296 3893 304
rect 4467 296 4513 304
rect 4707 296 4793 304
rect 5176 304 5184 313
rect 5176 296 5593 304
rect 467 276 573 284
rect 1067 276 1313 284
rect 1427 276 1493 284
rect 2136 284 2144 293
rect 2136 276 2293 284
rect 2347 276 2413 284
rect 2527 276 2613 284
rect 2627 276 2673 284
rect 3207 276 3293 284
rect 4327 276 4973 284
rect 5467 276 5573 284
rect 107 256 133 264
rect 147 256 433 264
rect 907 256 1033 264
rect 1167 256 1332 264
rect 1367 256 1393 264
rect 1407 256 1533 264
rect 1967 256 2493 264
rect 2647 256 3013 264
rect 3027 256 3173 264
rect 3327 256 3393 264
rect 3407 256 3553 264
rect 3747 256 3893 264
rect 3907 256 4233 264
rect 4387 256 4433 264
rect 4687 256 4733 264
rect 4787 256 4873 264
rect 5387 256 5513 264
rect 767 236 853 244
rect 876 236 1453 244
rect 447 216 693 224
rect 876 224 884 236
rect 1596 236 1633 244
rect 747 216 884 224
rect 1047 216 1233 224
rect 1347 216 1433 224
rect 1520 224 1533 227
rect 1516 213 1533 224
rect 1596 224 1604 236
rect 2067 236 2244 244
rect 1547 216 1604 224
rect 2027 216 2193 224
rect 2236 224 2244 236
rect 2387 236 2473 244
rect 2567 236 2753 244
rect 2947 236 3253 244
rect 3507 236 4293 244
rect 4307 236 4513 244
rect 4807 236 5053 244
rect 5147 236 5344 244
rect 2236 216 2513 224
rect 2907 216 2973 224
rect 3607 216 3693 224
rect 4347 216 4693 224
rect 4747 216 5073 224
rect 5336 224 5344 236
rect 5427 236 5533 244
rect 5547 236 5693 244
rect 5336 216 5473 224
rect 620 204 633 207
rect 507 196 564 204
rect 367 176 533 184
rect 227 136 253 144
rect 267 136 293 144
rect 556 144 564 196
rect 616 193 633 204
rect 827 196 993 204
rect 1287 196 1473 204
rect 616 146 624 193
rect 707 184 720 187
rect 707 173 724 184
rect 1107 176 1173 184
rect 1296 176 1353 184
rect 716 146 724 173
rect 556 136 573 144
rect 887 136 1053 144
rect 1067 135 1093 143
rect 1167 136 1193 144
rect 1296 146 1304 176
rect 1516 184 1524 213
rect 1627 196 1853 204
rect 2227 196 2252 204
rect 2667 204 2680 207
rect 2667 193 2684 204
rect 2827 196 2964 204
rect 1427 176 1524 184
rect 1667 177 1693 185
rect 1927 176 1973 184
rect 2076 176 2093 184
rect 1756 156 1793 164
rect 1207 136 1253 144
rect 1756 146 1764 156
rect 2076 164 2084 176
rect 2187 176 2244 184
rect 1807 156 2084 164
rect 1347 136 1393 144
rect 1627 135 1713 143
rect 1887 135 1913 143
rect 1967 135 2053 143
rect 2167 135 2193 143
rect 927 116 1013 124
rect 1447 116 1653 124
rect 2236 124 2244 176
rect 2276 146 2284 193
rect 2307 176 2373 184
rect 2427 176 2553 184
rect 2676 184 2684 193
rect 2676 176 2744 184
rect 2447 136 2533 144
rect 2596 144 2604 173
rect 2736 147 2744 176
rect 2767 177 2813 185
rect 2887 176 2924 184
rect 2587 136 2653 144
rect 2916 146 2924 176
rect 2956 146 2964 196
rect 3967 196 4204 204
rect 3067 177 3253 185
rect 3527 176 3633 184
rect 3647 176 3733 184
rect 3787 176 3853 184
rect 3876 176 3993 184
rect 3876 164 3884 176
rect 3216 156 3404 164
rect 3216 146 3224 156
rect 3396 146 3404 156
rect 3756 156 3884 164
rect 3756 146 3764 156
rect 4016 146 4024 196
rect 4047 177 4093 185
rect 4107 176 4173 184
rect 4196 146 4204 196
rect 4487 196 4613 204
rect 5167 196 5313 204
rect 4247 176 4273 184
rect 4296 146 4304 193
rect 5727 196 5773 204
rect 4340 184 4353 187
rect 4336 173 4353 184
rect 4336 146 4344 173
rect 4393 164 4407 173
rect 4495 176 4573 184
rect 4393 160 4424 164
rect 4396 156 4424 160
rect 4416 146 4424 156
rect 4495 147 4503 176
rect 4627 176 4693 184
rect 5040 184 5053 187
rect 5016 164 5024 174
rect 4947 156 5024 164
rect 5036 173 5053 184
rect 5227 176 5273 184
rect 5407 177 5433 185
rect 5540 184 5553 187
rect 5536 173 5553 184
rect 3267 136 3293 144
rect 3407 135 3433 143
rect 3847 135 3873 143
rect 3927 135 3973 143
rect 4067 136 4153 144
rect 4527 135 4553 143
rect 4767 135 4793 143
rect 5036 144 5044 173
rect 5007 136 5044 144
rect 5167 136 5253 144
rect 5536 146 5544 173
rect 5596 164 5604 193
rect 5596 156 5644 164
rect 5636 146 5644 156
rect 5676 146 5684 193
rect 5327 136 5373 144
rect 5727 136 5753 144
rect 2236 116 2373 124
rect 2487 116 2513 124
rect 2707 116 2793 124
rect 3067 116 3173 124
rect 4727 116 4893 124
rect 4907 116 4933 124
rect 4947 116 4973 124
rect 127 96 333 104
rect 507 96 573 104
rect 587 96 813 104
rect 1847 96 1953 104
rect 2147 96 2233 104
rect 2407 96 2573 104
rect 2647 96 2673 104
rect 2767 96 3033 104
rect 3287 96 3613 104
rect 3667 96 3913 104
rect 4107 96 4373 104
rect 4467 96 4593 104
rect 5047 96 5073 104
rect 5087 96 5213 104
rect 1647 76 3073 84
rect 3367 76 3473 84
rect 3587 76 4073 84
rect 4667 76 4833 84
rect 1667 56 2133 64
rect 2207 56 3053 64
rect 547 36 1433 44
rect 1487 36 1993 44
rect 2387 36 2533 44
rect 2687 36 2732 44
rect 2767 36 3013 44
rect 3087 36 3713 44
rect 3967 36 4913 44
rect 2347 16 2453 24
rect 2587 16 2653 24
rect 2707 16 2993 24
rect 3987 16 4493 24
use NOR2X1  _723_
timestamp 0
transform 1 0 2730 0 1 4950
box -6 -8 66 268
use INVX2  _724_
timestamp 0
transform -1 0 2670 0 -1 4950
box -6 -8 46 268
use NOR2X1  _725_
timestamp 0
transform -1 0 2390 0 1 3910
box -6 -8 66 268
use OAI21X1  _726_
timestamp 0
transform -1 0 2410 0 1 4950
box -6 -8 86 268
use INVX2  _727_
timestamp 0
transform 1 0 3090 0 1 3390
box -6 -8 46 268
use NOR2X1  _728_
timestamp 0
transform -1 0 3750 0 1 3390
box -6 -8 66 268
use AOI22X1  _729_
timestamp 0
transform -1 0 1090 0 1 4950
box -6 -8 106 268
use OAI21X1  _730_
timestamp 0
transform -1 0 2270 0 1 4950
box -6 -8 86 268
use INVX1  _731_
timestamp 0
transform -1 0 2310 0 -1 4950
box -6 -8 46 268
use INVX1  _732_
timestamp 0
transform -1 0 4210 0 -1 5470
box -6 -8 46 268
use NAND2X1  _733_
timestamp 0
transform 1 0 3330 0 -1 5470
box -6 -8 66 268
use OAI21X1  _734_
timestamp 0
transform 1 0 3190 0 -1 5470
box -6 -8 86 268
use AOI22X1  _735_
timestamp 0
transform -1 0 1270 0 1 4950
box -6 -8 106 268
use OAI21X1  _736_
timestamp 0
transform -1 0 2670 0 1 4950
box -6 -8 86 268
use INVX1  _737_
timestamp 0
transform -1 0 2770 0 -1 4950
box -6 -8 46 268
use NAND2X1  _738_
timestamp 0
transform 1 0 2510 0 -1 4950
box -6 -8 66 268
use OAI21X1  _739_
timestamp 0
transform 1 0 2370 0 -1 4950
box -6 -8 86 268
use AOI22X1  _740_
timestamp 0
transform -1 0 2010 0 -1 3910
box -6 -8 106 268
use OAI21X1  _741_
timestamp 0
transform -1 0 2210 0 -1 4950
box -6 -8 86 268
use NOR2X1  _742_
timestamp 0
transform 1 0 2790 0 -1 4430
box -6 -8 66 268
use OAI21X1  _743_
timestamp 0
transform -1 0 3030 0 1 3910
box -6 -8 86 268
use AOI22X1  _744_
timestamp 0
transform 1 0 1930 0 1 3910
box -6 -8 106 268
use OAI21X1  _745_
timestamp 0
transform -1 0 2710 0 -1 4430
box -6 -8 86 268
use INVX2  _746_
timestamp 0
transform -1 0 2910 0 -1 2350
box -6 -8 46 268
use NAND2X1  _747_
timestamp 0
transform -1 0 2150 0 -1 2350
box -6 -8 66 268
use OAI21X1  _748_
timestamp 0
transform -1 0 2390 0 1 1830
box -6 -8 86 268
use INVX1  _749_
timestamp 0
transform -1 0 4770 0 -1 1310
box -6 -8 46 268
use NAND2X1  _750_
timestamp 0
transform 1 0 2730 0 1 1830
box -6 -8 66 268
use OAI21X1  _751_
timestamp 0
transform 1 0 2570 0 1 1830
box -6 -8 86 268
use INVX2  _752_
timestamp 0
transform -1 0 4410 0 -1 2870
box -6 -8 46 268
use NAND2X1  _753_
timestamp 0
transform -1 0 4190 0 -1 2350
box -6 -8 66 268
use OAI21X1  _754_
timestamp 0
transform 1 0 4230 0 1 2350
box -6 -8 86 268
use INVX2  _755_
timestamp 0
transform -1 0 4190 0 1 1310
box -6 -8 46 268
use NAND2X1  _756_
timestamp 0
transform -1 0 3910 0 -1 2350
box -6 -8 66 268
use OAI21X1  _757_
timestamp 0
transform -1 0 4070 0 -1 2350
box -6 -8 86 268
use NAND2X1  _758_
timestamp 0
transform 1 0 2810 0 1 2350
box -6 -8 66 268
use OAI21X1  _759_
timestamp 0
transform -1 0 3010 0 1 2350
box -6 -8 86 268
use NAND2X1  _760_
timestamp 0
transform 1 0 3310 0 1 2350
box -6 -8 66 268
use OAI21X1  _761_
timestamp 0
transform -1 0 3510 0 1 2350
box -6 -8 86 268
use NAND2X1  _762_
timestamp 0
transform -1 0 4210 0 -1 2870
box -6 -8 66 268
use OAI21X1  _763_
timestamp 0
transform 1 0 4010 0 -1 2870
box -6 -8 86 268
use NAND2X1  _764_
timestamp 0
transform 1 0 3710 0 1 2350
box -6 -8 66 268
use OAI21X1  _765_
timestamp 0
transform -1 0 3930 0 1 2350
box -6 -8 86 268
use INVX1  _766_
timestamp 0
transform 1 0 410 0 1 3390
box -6 -8 46 268
use NAND2X1  _767_
timestamp 0
transform -1 0 2770 0 1 3390
box -6 -8 66 268
use OAI21X1  _768_
timestamp 0
transform 1 0 750 0 1 3390
box -6 -8 86 268
use INVX1  _769_
timestamp 0
transform -1 0 350 0 -1 5470
box -6 -8 46 268
use NAND2X1  _770_
timestamp 0
transform 1 0 790 0 -1 5470
box -6 -8 66 268
use OAI21X1  _771_
timestamp 0
transform 1 0 650 0 -1 5470
box -6 -8 86 268
use INVX1  _772_
timestamp 0
transform 1 0 2110 0 1 3390
box -6 -8 46 268
use NAND2X1  _773_
timestamp 0
transform 1 0 2590 0 1 3390
box -6 -8 66 268
use OAI21X1  _774_
timestamp 0
transform 1 0 2210 0 1 3390
box -6 -8 86 268
use INVX1  _775_
timestamp 0
transform 1 0 430 0 1 2870
box -6 -8 46 268
use NAND2X1  _776_
timestamp 0
transform 1 0 2270 0 1 2870
box -6 -8 66 268
use OAI21X1  _777_
timestamp 0
transform 1 0 670 0 1 2870
box -6 -8 86 268
use INVX1  _778_
timestamp 0
transform 1 0 70 0 1 3390
box -6 -8 46 268
use NAND2X1  _779_
timestamp 0
transform 1 0 350 0 -1 3390
box -6 -8 66 268
use OAI21X1  _780_
timestamp 0
transform 1 0 210 0 -1 3390
box -6 -8 86 268
use INVX1  _781_
timestamp 0
transform 1 0 1210 0 1 3910
box -6 -8 46 268
use NAND2X1  _782_
timestamp 0
transform 1 0 2470 0 1 3390
box -6 -8 66 268
use OAI21X1  _783_
timestamp 0
transform 1 0 1550 0 1 3910
box -6 -8 86 268
use INVX1  _784_
timestamp 0
transform -1 0 1370 0 1 2870
box -6 -8 46 268
use NAND2X1  _785_
timestamp 0
transform 1 0 2150 0 1 2870
box -6 -8 66 268
use OAI21X1  _786_
timestamp 0
transform 1 0 1670 0 1 2870
box -6 -8 86 268
use INVX1  _787_
timestamp 0
transform 1 0 2310 0 -1 2870
box -6 -8 46 268
use NAND2X1  _788_
timestamp 0
transform 1 0 2810 0 -1 2870
box -6 -8 66 268
use OAI21X1  _789_
timestamp 0
transform 1 0 2650 0 -1 2870
box -6 -8 86 268
use INVX1  _790_
timestamp 0
transform 1 0 1410 0 -1 5470
box -6 -8 46 268
use NAND2X1  _791_
timestamp 0
transform 1 0 1650 0 -1 5470
box -6 -8 66 268
use OAI21X1  _792_
timestamp 0
transform 1 0 1510 0 -1 5470
box -6 -8 86 268
use INVX1  _793_
timestamp 0
transform 1 0 2010 0 -1 4430
box -6 -8 46 268
use NAND2X1  _794_
timestamp 0
transform 1 0 2510 0 -1 4430
box -6 -8 66 268
use OAI21X1  _795_
timestamp 0
transform -1 0 2450 0 -1 4430
box -6 -8 86 268
use INVX1  _796_
timestamp 0
transform -1 0 4810 0 -1 4430
box -6 -8 46 268
use NAND2X1  _797_
timestamp 0
transform -1 0 4530 0 1 3910
box -6 -8 66 268
use OAI21X1  _798_
timestamp 0
transform -1 0 4670 0 1 3910
box -6 -8 86 268
use INVX1  _799_
timestamp 0
transform -1 0 5450 0 1 3910
box -6 -8 46 268
use NAND2X1  _800_
timestamp 0
transform -1 0 4410 0 1 3910
box -6 -8 66 268
use OAI21X1  _801_
timestamp 0
transform -1 0 5350 0 1 3910
box -6 -8 86 268
use INVX1  _802_
timestamp 0
transform -1 0 5790 0 1 270
box -6 -8 46 268
use NAND2X1  _803_
timestamp 0
transform -1 0 5630 0 -1 3910
box -6 -8 66 268
use OAI21X1  _804_
timestamp 0
transform 1 0 5430 0 1 4950
box -6 -8 86 268
use INVX1  _805_
timestamp 0
transform 1 0 5310 0 -1 4950
box -6 -8 46 268
use NAND2X1  _806_
timestamp 0
transform -1 0 4470 0 -1 4430
box -6 -8 66 268
use OAI21X1  _807_
timestamp 0
transform -1 0 4670 0 -1 4950
box -6 -8 86 268
use INVX1  _808_
timestamp 0
transform -1 0 3750 0 1 4950
box -6 -8 46 268
use NAND2X1  _809_
timestamp 0
transform 1 0 3150 0 -1 4430
box -6 -8 66 268
use OAI21X1  _810_
timestamp 0
transform 1 0 3110 0 1 4430
box -6 -8 86 268
use INVX1  _811_
timestamp 0
transform -1 0 3810 0 -1 4950
box -6 -8 46 268
use NAND2X1  _812_
timestamp 0
transform -1 0 4510 0 1 3390
box -6 -8 66 268
use OAI21X1  _813_
timestamp 0
transform 1 0 3770 0 -1 4430
box -6 -8 86 268
use INVX1  _814_
timestamp 0
transform 1 0 650 0 1 2350
box -6 -8 46 268
use NAND3X1  _815_
timestamp 0
transform -1 0 2150 0 1 2350
box -6 -8 86 268
use OAI21X1  _816_
timestamp 0
transform 1 0 750 0 1 2350
box -6 -8 86 268
use INVX8  _817_
timestamp 0
transform 1 0 1170 0 1 4430
box -6 -8 106 268
use NAND2X1  _818_
timestamp 0
transform 1 0 1610 0 -1 2350
box -6 -8 66 268
use NAND2X1  _819_
timestamp 0
transform -1 0 1790 0 -1 2350
box -6 -8 66 268
use XNOR2X1  _820_
timestamp 0
transform 1 0 1510 0 1 2350
box -6 -8 126 268
use NAND2X1  _821_
timestamp 0
transform 1 0 1010 0 -1 4430
box -6 -8 66 268
use OAI21X1  _822_
timestamp 0
transform -1 0 1450 0 -1 4430
box -6 -8 86 268
use NOR2X1  _823_
timestamp 0
transform -1 0 1530 0 -1 2350
box -6 -8 66 268
use NAND2X1  _824_
timestamp 0
transform 1 0 1530 0 1 1830
box -6 -8 66 268
use NAND2X1  _825_
timestamp 0
transform 1 0 1370 0 1 1310
box -6 -8 66 268
use NOR2X1  _826_
timestamp 0
transform -1 0 1190 0 1 1830
box -6 -8 66 268
use AOI22X1  _827_
timestamp 0
transform 1 0 1650 0 1 1830
box -6 -8 106 268
use OAI21X1  _828_
timestamp 0
transform 1 0 1250 0 1 1830
box -6 -8 86 268
use INVX1  _829_
timestamp 0
transform 1 0 1350 0 -1 1830
box -6 -8 46 268
use AND2X2  _830_
timestamp 0
transform -1 0 1650 0 -1 1830
box -6 -8 86 268
use AND2X2  _831_
timestamp 0
transform 1 0 1710 0 -1 1830
box -6 -8 86 268
use NAND2X1  _832_
timestamp 0
transform -1 0 1510 0 -1 1830
box -6 -8 66 268
use INVX1  _833_
timestamp 0
transform 1 0 1870 0 -1 2350
box -6 -8 46 268
use INVX1  _834_
timestamp 0
transform 1 0 1810 0 1 1830
box -6 -8 46 268
use NAND2X1  _835_
timestamp 0
transform -1 0 2030 0 -1 2350
box -6 -8 66 268
use OAI21X1  _836_
timestamp 0
transform 1 0 1910 0 1 1830
box -6 -8 86 268
use NAND3X1  _837_
timestamp 0
transform -1 0 1470 0 1 1830
box -6 -8 86 268
use NAND3X1  _838_
timestamp 0
transform -1 0 1410 0 -1 2350
box -6 -8 86 268
use INVX1  _839_
timestamp 0
transform -1 0 970 0 -1 2350
box -6 -8 46 268
use AOI21X1  _840_
timestamp 0
transform -1 0 1270 0 -1 2350
box -6 -8 86 268
use OAI21X1  _841_
timestamp 0
transform -1 0 1130 0 -1 2350
box -6 -8 86 268
use INVX1  _842_
timestamp 0
transform 1 0 1930 0 1 2870
box -6 -8 46 268
use NAND2X1  _843_
timestamp 0
transform -1 0 1870 0 1 2870
box -6 -8 66 268
use AND2X2  _844_
timestamp 0
transform 1 0 1690 0 1 2350
box -6 -8 86 268
use INVX1  _845_
timestamp 0
transform 1 0 430 0 -1 2870
box -6 -8 46 268
use NAND2X1  _846_
timestamp 0
transform -1 0 2250 0 1 1830
box -6 -8 66 268
use AOI21X1  _847_
timestamp 0
transform -1 0 1070 0 1 1830
box -6 -8 86 268
use NAND2X1  _848_
timestamp 0
transform -1 0 1570 0 1 1310
box -6 -8 66 268
use NAND2X1  _849_
timestamp 0
transform 1 0 1110 0 1 1310
box -6 -8 66 268
use NOR2X1  _850_
timestamp 0
transform -1 0 1050 0 1 1310
box -6 -8 66 268
use AOI22X1  _851_
timestamp 0
transform -1 0 1350 0 -1 1310
box -6 -8 106 268
use OAI21X1  _852_
timestamp 0
transform -1 0 790 0 1 1310
box -6 -8 86 268
use INVX1  _853_
timestamp 0
transform -1 0 950 0 -1 1310
box -6 -8 46 268
use AND2X2  _854_
timestamp 0
transform 1 0 1110 0 -1 1310
box -6 -8 86 268
use NAND2X1  _855_
timestamp 0
transform -1 0 1290 0 1 1310
box -6 -8 66 268
use INVX1  _856_
timestamp 0
transform 1 0 530 0 -1 1310
box -6 -8 46 268
use NAND3X1  _857_
timestamp 0
transform -1 0 650 0 1 1310
box -6 -8 86 268
use NAND3X1  _858_
timestamp 0
transform 1 0 710 0 1 1830
box -6 -8 86 268
use OAI21X1  _859_
timestamp 0
transform -1 0 1290 0 -1 1830
box -6 -8 86 268
use AOI21X1  _860_
timestamp 0
transform -1 0 930 0 1 1310
box -6 -8 86 268
use INVX2  _861_
timestamp 0
transform 1 0 1970 0 -1 1830
box -6 -8 46 268
use OAI21X1  _862_
timestamp 0
transform -1 0 1850 0 1 1310
box -6 -8 86 268
use INVX2  _863_
timestamp 0
transform -1 0 2910 0 1 1830
box -6 -8 46 268
use INVX1  _864_
timestamp 0
transform -1 0 2770 0 1 790
box -6 -8 46 268
use OAI21X1  _865_
timestamp 0
transform -1 0 2110 0 1 1310
box -6 -8 86 268
use AOI21X1  _866_
timestamp 0
transform -1 0 1710 0 1 1310
box -6 -8 86 268
use OAI21X1  _867_
timestamp 0
transform 1 0 1070 0 -1 1830
box -6 -8 86 268
use NAND3X1  _868_
timestamp 0
transform 1 0 850 0 1 1830
box -6 -8 86 268
use INVX1  _869_
timestamp 0
transform -1 0 510 0 1 1830
box -6 -8 46 268
use NAND3X1  _870_
timestamp 0
transform -1 0 730 0 -1 1830
box -6 -8 86 268
use OAI21X1  _871_
timestamp 0
transform -1 0 1010 0 -1 1830
box -6 -8 86 268
use NAND3X1  _872_
timestamp 0
transform 1 0 570 0 1 1830
box -6 -8 86 268
use AOI21X1  _873_
timestamp 0
transform -1 0 730 0 -1 2350
box -6 -8 86 268
use NAND3X1  _874_
timestamp 0
transform -1 0 870 0 -1 2350
box -6 -8 86 268
use NAND2X1  _875_
timestamp 0
transform 1 0 370 0 -1 2350
box -6 -8 66 268
use OAI22X1  _876_
timestamp 0
transform 1 0 490 0 -1 2350
box -6 -8 106 268
use INVX1  _877_
timestamp 0
transform -1 0 110 0 1 2350
box -6 -8 46 268
use INVX1  _878_
timestamp 0
transform -1 0 410 0 1 1830
box -6 -8 46 268
use AOI21X1  _879_
timestamp 0
transform -1 0 590 0 -1 1830
box -6 -8 86 268
use OAI21X1  _880_
timestamp 0
transform -1 0 510 0 1 1310
box -6 -8 86 268
use OAI21X1  _881_
timestamp 0
transform -1 0 710 0 -1 1310
box -6 -8 86 268
use AND2X2  _882_
timestamp 0
transform 1 0 1610 0 1 790
box -6 -8 86 268
use NAND2X1  _883_
timestamp 0
transform 1 0 1210 0 1 790
box -6 -8 66 268
use AOI22X1  _884_
timestamp 0
transform 1 0 1410 0 -1 1310
box -6 -8 106 268
use INVX1  _885_
timestamp 0
transform -1 0 1050 0 -1 1310
box -6 -8 46 268
use NAND2X1  _886_
timestamp 0
transform 1 0 1350 0 1 790
box -6 -8 66 268
use INVX1  _887_
timestamp 0
transform -1 0 910 0 -1 790
box -6 -8 46 268
use NAND3X1  _888_
timestamp 0
transform -1 0 990 0 1 790
box -6 -8 86 268
use NAND2X1  _889_
timestamp 0
transform -1 0 2410 0 1 790
box -6 -8 66 268
use NOR2X1  _890_
timestamp 0
transform 1 0 970 0 -1 790
box -6 -8 66 268
use OAI21X1  _891_
timestamp 0
transform 1 0 770 0 1 790
box -6 -8 86 268
use AOI21X1  _892_
timestamp 0
transform -1 0 710 0 1 790
box -6 -8 86 268
use AOI21X1  _893_
timestamp 0
transform -1 0 850 0 -1 1310
box -6 -8 86 268
use NAND3X1  _894_
timestamp 0
transform -1 0 1150 0 1 790
box -6 -8 86 268
use OAI21X1  _895_
timestamp 0
transform -1 0 810 0 -1 790
box -6 -8 86 268
use AOI21X1  _896_
timestamp 0
transform -1 0 530 0 -1 790
box -6 -8 86 268
use NAND2X1  _897_
timestamp 0
transform 1 0 2730 0 1 1310
box -6 -8 66 268
use INVX1  _898_
timestamp 0
transform 1 0 2210 0 1 2350
box -6 -8 46 268
use INVX2  _899_
timestamp 0
transform 1 0 4270 0 -1 2870
box -6 -8 46 268
use NAND2X1  _900_
timestamp 0
transform -1 0 2370 0 1 1310
box -6 -8 66 268
use OAI21X1  _901_
timestamp 0
transform 1 0 2230 0 -1 2350
box -6 -8 86 268
use OAI21X1  _902_
timestamp 0
transform -1 0 2250 0 1 1310
box -6 -8 86 268
use OAI21X1  _903_
timestamp 0
transform 1 0 350 0 1 790
box -6 -8 86 268
use NAND3X1  _904_
timestamp 0
transform -1 0 670 0 -1 790
box -6 -8 86 268
use NAND3X1  _905_
timestamp 0
transform -1 0 570 0 1 790
box -6 -8 86 268
use INVX1  _906_
timestamp 0
transform 1 0 70 0 -1 790
box -6 -8 46 268
use NAND3X1  _907_
timestamp 0
transform 1 0 210 0 1 790
box -6 -8 86 268
use NAND3X1  _908_
timestamp 0
transform -1 0 450 0 -1 1310
box -6 -8 86 268
use INVX1  _909_
timestamp 0
transform 1 0 410 0 -1 1830
box -6 -8 46 268
use AOI21X1  _910_
timestamp 0
transform -1 0 330 0 -1 1830
box -6 -8 86 268
use AOI21X1  _911_
timestamp 0
transform -1 0 150 0 1 790
box -6 -8 86 268
use INVX1  _912_
timestamp 0
transform -1 0 370 0 1 1310
box -6 -8 46 268
use OAI21X1  _913_
timestamp 0
transform 1 0 190 0 1 1310
box -6 -8 86 268
use AOI21X1  _914_
timestamp 0
transform 1 0 70 0 1 1830
box -6 -8 86 268
use NAND3X1  _915_
timestamp 0
transform 1 0 210 0 1 1830
box -6 -8 86 268
use NAND2X1  _916_
timestamp 0
transform 1 0 250 0 -1 2350
box -6 -8 66 268
use OAI22X1  _917_
timestamp 0
transform 1 0 70 0 -1 2350
box -6 -8 106 268
use AND2X2  _918_
timestamp 0
transform 1 0 2870 0 -1 1830
box -6 -8 86 268
use NAND2X1  _919_
timestamp 0
transform 1 0 790 0 -1 1830
box -6 -8 66 268
use INVX1  _920_
timestamp 0
transform 1 0 190 0 -1 270
box -6 -8 46 268
use AOI21X1  _921_
timestamp 0
transform 1 0 170 0 -1 790
box -6 -8 86 268
use NAND2X1  _922_
timestamp 0
transform 1 0 2450 0 1 1830
box -6 -8 66 268
use AND2X2  _923_
timestamp 0
transform 1 0 2070 0 -1 1830
box -6 -8 86 268
use OAI21X1  _924_
timestamp 0
transform 1 0 2230 0 -1 1830
box -6 -8 86 268
use INVX2  _925_
timestamp 0
transform 1 0 3910 0 1 1310
box -6 -8 46 268
use OAI21X1  _926_
timestamp 0
transform -1 0 2810 0 -1 1830
box -6 -8 86 268
use NAND3X1  _927_
timestamp 0
transform 1 0 2590 0 -1 1830
box -6 -8 86 268
use INVX1  _928_
timestamp 0
transform -1 0 2530 0 -1 1830
box -6 -8 46 268
use NAND2X1  _929_
timestamp 0
transform 1 0 2370 0 -1 1830
box -6 -8 66 268
use OAI21X1  _930_
timestamp 0
transform -1 0 2670 0 1 1310
box -6 -8 86 268
use NAND3X1  _931_
timestamp 0
transform -1 0 2530 0 1 1310
box -6 -8 86 268
use NAND2X1  _932_
timestamp 0
transform -1 0 2230 0 -1 1310
box -6 -8 66 268
use OAI22X1  _933_
timestamp 0
transform 1 0 1090 0 -1 790
box -6 -8 106 268
use INVX1  _934_
timestamp 0
transform 1 0 1130 0 -1 270
box -6 -8 46 268
use NAND2X1  _935_
timestamp 0
transform 1 0 1570 0 -1 1310
box -6 -8 66 268
use NAND3X1  _936_
timestamp 0
transform -1 0 2090 0 -1 790
box -6 -8 86 268
use NAND2X1  _937_
timestamp 0
transform -1 0 2290 0 1 790
box -6 -8 66 268
use NAND3X1  _938_
timestamp 0
transform -1 0 1550 0 1 790
box -6 -8 86 268
use NAND3X1  _939_
timestamp 0
transform -1 0 1510 0 -1 790
box -6 -8 86 268
use INVX1  _940_
timestamp 0
transform -1 0 1790 0 1 790
box -6 -8 46 268
use AND2X2  _941_
timestamp 0
transform -1 0 2910 0 1 790
box -6 -8 86 268
use NAND2X1  _942_
timestamp 0
transform 1 0 1850 0 1 790
box -6 -8 66 268
use OAI21X1  _943_
timestamp 0
transform -1 0 2550 0 1 790
box -6 -8 86 268
use NAND3X1  _944_
timestamp 0
transform -1 0 1650 0 -1 790
box -6 -8 86 268
use NAND3X1  _945_
timestamp 0
transform -1 0 1310 0 -1 270
box -6 -8 86 268
use AOI21X1  _946_
timestamp 0
transform -1 0 1790 0 -1 790
box -6 -8 86 268
use AOI21X1  _947_
timestamp 0
transform -1 0 1350 0 -1 790
box -6 -8 86 268
use OAI21X1  _948_
timestamp 0
transform -1 0 1170 0 1 270
box -6 -8 86 268
use NAND3X1  _949_
timestamp 0
transform -1 0 1070 0 -1 270
box -6 -8 86 268
use AND2X2  _950_
timestamp 0
transform -1 0 2110 0 -1 1310
box -6 -8 86 268
use NAND3X1  _951_
timestamp 0
transform 1 0 1370 0 1 270
box -6 -8 86 268
use OAI21X1  _952_
timestamp 0
transform -1 0 1310 0 1 270
box -6 -8 86 268
use NAND3X1  _953_
timestamp 0
transform -1 0 890 0 1 270
box -6 -8 86 268
use NAND3X1  _954_
timestamp 0
transform -1 0 470 0 1 270
box -6 -8 86 268
use OAI21X1  _955_
timestamp 0
transform -1 0 390 0 -1 790
box -6 -8 86 268
use AOI21X1  _956_
timestamp 0
transform -1 0 1030 0 1 270
box -6 -8 86 268
use AOI21X1  _957_
timestamp 0
transform -1 0 930 0 -1 270
box -6 -8 86 268
use OAI21X1  _958_
timestamp 0
transform -1 0 750 0 1 270
box -6 -8 86 268
use NAND3X1  _959_
timestamp 0
transform -1 0 310 0 1 270
box -6 -8 86 268
use NAND3X1  _960_
timestamp 0
transform -1 0 510 0 -1 270
box -6 -8 86 268
use OAI21X1  _961_
timestamp 0
transform -1 0 610 0 1 270
box -6 -8 86 268
use NAND3X1  _962_
timestamp 0
transform -1 0 170 0 1 270
box -6 -8 86 268
use NAND2X1  _963_
timestamp 0
transform -1 0 130 0 -1 1310
box -6 -8 66 268
use NAND2X1  _964_
timestamp 0
transform 1 0 70 0 1 1310
box -6 -8 66 268
use XNOR2X1  _965_
timestamp 0
transform 1 0 70 0 -1 1830
box -6 -8 126 268
use NAND2X1  _966_
timestamp 0
transform -1 0 930 0 -1 3910
box -6 -8 66 268
use OAI21X1  _967_
timestamp 0
transform -1 0 1070 0 -1 3910
box -6 -8 86 268
use INVX1  _968_
timestamp 0
transform 1 0 1130 0 1 2350
box -6 -8 46 268
use AOI22X1  _969_
timestamp 0
transform 1 0 210 0 -1 1310
box -6 -8 106 268
use AOI21X1  _970_
timestamp 0
transform 1 0 570 0 -1 270
box -6 -8 86 268
use OAI21X1  _971_
timestamp 0
transform -1 0 790 0 -1 270
box -6 -8 86 268
use NAND2X1  _972_
timestamp 0
transform 1 0 2850 0 1 1310
box -6 -8 66 268
use OAI21X1  _973_
timestamp 0
transform 1 0 2290 0 -1 1310
box -6 -8 86 268
use INVX1  _974_
timestamp 0
transform 1 0 2310 0 -1 790
box -6 -8 46 268
use INVX1  _975_
timestamp 0
transform 1 0 1790 0 1 270
box -6 -8 46 268
use AOI21X1  _976_
timestamp 0
transform 1 0 1890 0 1 270
box -6 -8 86 268
use NAND2X1  _977_
timestamp 0
transform 1 0 2990 0 1 1830
box -6 -8 66 268
use AND2X2  _978_
timestamp 0
transform -1 0 3470 0 -1 1830
box -6 -8 86 268
use OAI21X1  _979_
timestamp 0
transform 1 0 3250 0 -1 1830
box -6 -8 86 268
use AND2X2  _980_
timestamp 0
transform -1 0 3590 0 1 1310
box -6 -8 86 268
use OAI21X1  _981_
timestamp 0
transform -1 0 3610 0 -1 1830
box -6 -8 86 268
use NAND3X1  _982_
timestamp 0
transform -1 0 3190 0 -1 1830
box -6 -8 86 268
use INVX1  _983_
timestamp 0
transform -1 0 3050 0 -1 1830
box -6 -8 46 268
use NAND2X1  _984_
timestamp 0
transform -1 0 3450 0 1 1310
box -6 -8 66 268
use OAI21X1  _985_
timestamp 0
transform -1 0 3050 0 1 1310
box -6 -8 86 268
use NAND3X1  _986_
timestamp 0
transform 1 0 3110 0 1 1310
box -6 -8 86 268
use NAND2X1  _987_
timestamp 0
transform -1 0 2970 0 -1 1310
box -6 -8 66 268
use NOR2X1  _988_
timestamp 0
transform -1 0 2170 0 1 790
box -6 -8 66 268
use AOI21X1  _989_
timestamp 0
transform 1 0 1970 0 1 790
box -6 -8 86 268
use NAND2X1  _990_
timestamp 0
transform 1 0 3790 0 -1 790
box -6 -8 66 268
use NAND2X1  _991_
timestamp 0
transform -1 0 3230 0 -1 1310
box -6 -8 66 268
use NAND3X1  _992_
timestamp 0
transform -1 0 3550 0 -1 1310
box -6 -8 86 268
use NAND2X1  _993_
timestamp 0
transform -1 0 3830 0 -1 1310
box -6 -8 66 268
use NAND3X1  _994_
timestamp 0
transform -1 0 3910 0 1 790
box -6 -8 86 268
use NAND3X1  _995_
timestamp 0
transform -1 0 3630 0 1 790
box -6 -8 86 268
use INVX1  _996_
timestamp 0
transform -1 0 3450 0 -1 790
box -6 -8 46 268
use AND2X2  _997_
timestamp 0
transform -1 0 3850 0 1 1310
box -6 -8 86 268
use NAND2X1  _998_
timestamp 0
transform 1 0 3670 0 -1 790
box -6 -8 66 268
use OAI21X1  _999_
timestamp 0
transform -1 0 3390 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1000_
timestamp 0
transform -1 0 3350 0 -1 790
box -6 -8 86 268
use NAND3X1  _1001_
timestamp 0
transform -1 0 2770 0 -1 790
box -6 -8 86 268
use AOI22X1  _1002_
timestamp 0
transform -1 0 2250 0 -1 790
box -6 -8 106 268
use OAI21X1  _1003_
timestamp 0
transform 1 0 1870 0 -1 790
box -6 -8 86 268
use AOI22X1  _1004_
timestamp 0
transform 1 0 3250 0 1 790
box -6 -8 106 268
use AOI21X1  _1005_
timestamp 0
transform -1 0 3490 0 1 790
box -6 -8 86 268
use OAI21X1  _1006_
timestamp 0
transform -1 0 3050 0 1 790
box -6 -8 86 268
use NAND3X1  _1007_
timestamp 0
transform 1 0 2550 0 -1 790
box -6 -8 86 268
use AND2X2  _1008_
timestamp 0
transform 1 0 3030 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1009_
timestamp 0
transform 1 0 2970 0 -1 790
box -6 -8 86 268
use OAI21X1  _1010_
timestamp 0
transform -1 0 3190 0 1 790
box -6 -8 86 268
use NAND3X1  _1011_
timestamp 0
transform -1 0 3270 0 1 270
box -6 -8 86 268
use NAND3X1  _1012_
timestamp 0
transform -1 0 2690 0 1 270
box -6 -8 86 268
use AOI21X1  _1013_
timestamp 0
transform 1 0 1510 0 1 270
box -6 -8 86 268
use OAI21X1  _1014_
timestamp 0
transform 1 0 1650 0 1 270
box -6 -8 86 268
use AOI21X1  _1015_
timestamp 0
transform -1 0 3110 0 1 270
box -6 -8 86 268
use AOI21X1  _1016_
timestamp 0
transform -1 0 2490 0 -1 790
box -6 -8 86 268
use OAI21X1  _1017_
timestamp 0
transform -1 0 2410 0 1 270
box -6 -8 86 268
use NAND3X1  _1018_
timestamp 0
transform -1 0 2130 0 1 270
box -6 -8 86 268
use NAND3X1  _1019_
timestamp 0
transform -1 0 2830 0 1 270
box -6 -8 86 268
use OAI21X1  _1020_
timestamp 0
transform 1 0 2470 0 1 270
box -6 -8 86 268
use NAND3X1  _1021_
timestamp 0
transform -1 0 2590 0 -1 270
box -6 -8 86 268
use NAND2X1  _1022_
timestamp 0
transform 1 0 1830 0 -1 270
box -6 -8 66 268
use XNOR2X1  _1023_
timestamp 0
transform -1 0 1610 0 -1 270
box -6 -8 126 268
use NOR2X1  _1024_
timestamp 0
transform 1 0 1370 0 -1 270
box -6 -8 66 268
use NAND3X1  _1025_
timestamp 0
transform 1 0 1950 0 -1 270
box -6 -8 86 268
use INVX1  _1026_
timestamp 0
transform 1 0 90 0 -1 270
box -6 -8 46 268
use AOI21X1  _1027_
timestamp 0
transform 1 0 290 0 -1 270
box -6 -8 86 268
use AOI21X1  _1028_
timestamp 0
transform -1 0 2450 0 -1 270
box -6 -8 86 268
use AOI21X1  _1029_
timestamp 0
transform 1 0 2190 0 1 270
box -6 -8 86 268
use OAI21X1  _1030_
timestamp 0
transform -1 0 2310 0 -1 270
box -6 -8 86 268
use NAND3X1  _1031_
timestamp 0
transform -1 0 2170 0 -1 270
box -6 -8 86 268
use NAND2X1  _1032_
timestamp 0
transform 1 0 1390 0 1 2350
box -6 -8 66 268
use OAI22X1  _1033_
timestamp 0
transform 1 0 1230 0 1 2350
box -6 -8 106 268
use OAI21X1  _1034_
timestamp 0
transform 1 0 1690 0 -1 270
box -6 -8 86 268
use INVX1  _1035_
timestamp 0
transform -1 0 2830 0 -1 270
box -6 -8 46 268
use AOI21X1  _1036_
timestamp 0
transform 1 0 2650 0 -1 270
box -6 -8 86 268
use NAND2X1  _1037_
timestamp 0
transform -1 0 3310 0 1 1310
box -6 -8 66 268
use INVX1  _1038_
timestamp 0
transform 1 0 3830 0 1 270
box -6 -8 46 268
use INVX1  _1039_
timestamp 0
transform 1 0 3330 0 1 270
box -6 -8 46 268
use AOI21X1  _1040_
timestamp 0
transform 1 0 3430 0 1 270
box -6 -8 86 268
use NAND2X1  _1041_
timestamp 0
transform 1 0 4050 0 1 1830
box -6 -8 66 268
use AND2X2  _1042_
timestamp 0
transform 1 0 3770 0 1 1830
box -6 -8 86 268
use OAI21X1  _1043_
timestamp 0
transform -1 0 4410 0 -1 1830
box -6 -8 86 268
use AND2X2  _1044_
timestamp 0
transform 1 0 3490 0 1 1830
box -6 -8 86 268
use OAI21X1  _1045_
timestamp 0
transform 1 0 3630 0 1 1830
box -6 -8 86 268
use NAND3X1  _1046_
timestamp 0
transform 1 0 4190 0 -1 1830
box -6 -8 86 268
use INVX1  _1047_
timestamp 0
transform -1 0 4130 0 -1 1830
box -6 -8 46 268
use NAND2X1  _1048_
timestamp 0
transform 1 0 3910 0 1 1830
box -6 -8 66 268
use NAND2X1  _1049_
timestamp 0
transform -1 0 3750 0 -1 1830
box -6 -8 66 268
use OAI21X1  _1050_
timestamp 0
transform -1 0 3890 0 -1 1830
box -6 -8 86 268
use NAND3X1  _1051_
timestamp 0
transform -1 0 4030 0 -1 1830
box -6 -8 86 268
use NAND2X1  _1052_
timestamp 0
transform -1 0 4870 0 1 270
box -6 -8 66 268
use AOI22X1  _1053_
timestamp 0
transform -1 0 3610 0 -1 790
box -6 -8 106 268
use NAND2X1  _1054_
timestamp 0
transform 1 0 3970 0 1 790
box -6 -8 66 268
use NAND2X1  _1055_
timestamp 0
transform 1 0 4830 0 -1 1310
box -6 -8 66 268
use NOR2X1  _1056_
timestamp 0
transform 1 0 4970 0 -1 1310
box -6 -8 66 268
use AOI22X1  _1057_
timestamp 0
transform -1 0 4530 0 -1 1310
box -6 -8 106 268
use OAI21X1  _1058_
timestamp 0
transform -1 0 4550 0 1 790
box -6 -8 86 268
use INVX1  _1059_
timestamp 0
transform 1 0 4090 0 1 790
box -6 -8 46 268
use AND2X2  _1060_
timestamp 0
transform -1 0 4250 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1061_
timestamp 0
transform -1 0 4370 0 -1 1310
box -6 -8 66 268
use INVX1  _1062_
timestamp 0
transform 1 0 4610 0 1 790
box -6 -8 46 268
use NAND3X1  _1063_
timestamp 0
transform 1 0 4330 0 1 790
box -6 -8 86 268
use NAND3X1  _1064_
timestamp 0
transform 1 0 4390 0 1 270
box -6 -8 86 268
use AOI22X1  _1065_
timestamp 0
transform -1 0 3710 0 -1 1310
box -6 -8 106 268
use OAI21X1  _1066_
timestamp 0
transform -1 0 3770 0 1 790
box -6 -8 86 268
use AOI21X1  _1067_
timestamp 0
transform -1 0 4270 0 1 790
box -6 -8 86 268
use OAI21X1  _1068_
timestamp 0
transform 1 0 4010 0 1 1310
box -6 -8 86 268
use OAI21X1  _1069_
timestamp 0
transform 1 0 3890 0 -1 1310
box -6 -8 86 268
use AOI21X1  _1070_
timestamp 0
transform 1 0 4030 0 -1 1310
box -6 -8 86 268
use OAI21X1  _1071_
timestamp 0
transform -1 0 4130 0 -1 790
box -6 -8 86 268
use NAND3X1  _1072_
timestamp 0
transform -1 0 4610 0 1 270
box -6 -8 86 268
use AND2X2  _1073_
timestamp 0
transform 1 0 4830 0 -1 270
box -6 -8 86 268
use NAND3X1  _1074_
timestamp 0
transform 1 0 4470 0 -1 790
box -6 -8 86 268
use OAI21X1  _1075_
timestamp 0
transform 1 0 4190 0 -1 790
box -6 -8 86 268
use NAND3X1  _1076_
timestamp 0
transform -1 0 5050 0 -1 270
box -6 -8 86 268
use NAND3X1  _1077_
timestamp 0
transform -1 0 4350 0 -1 270
box -6 -8 86 268
use AOI21X1  _1078_
timestamp 0
transform 1 0 2830 0 -1 790
box -6 -8 86 268
use OAI21X1  _1079_
timestamp 0
transform 1 0 3130 0 -1 790
box -6 -8 86 268
use AOI21X1  _1080_
timestamp 0
transform -1 0 4770 0 -1 270
box -6 -8 86 268
use AOI21X1  _1081_
timestamp 0
transform 1 0 4670 0 1 270
box -6 -8 86 268
use OAI21X1  _1082_
timestamp 0
transform -1 0 4490 0 -1 270
box -6 -8 86 268
use AOI21X1  _1083_
timestamp 0
transform -1 0 4070 0 -1 270
box -6 -8 86 268
use NAND3X1  _1084_
timestamp 0
transform -1 0 4310 0 1 270
box -6 -8 86 268
use OAI21X1  _1085_
timestamp 0
transform -1 0 4630 0 -1 270
box -6 -8 86 268
use AOI21X1  _1086_
timestamp 0
transform -1 0 3930 0 -1 270
box -6 -8 86 268
use OAI21X1  _1087_
timestamp 0
transform -1 0 3790 0 -1 270
box -6 -8 86 268
use AOI21X1  _1088_
timestamp 0
transform -1 0 2970 0 1 270
box -6 -8 86 268
use OAI21X1  _1089_
timestamp 0
transform 1 0 2890 0 -1 270
box -6 -8 86 268
use NAND3X1  _1090_
timestamp 0
transform -1 0 3770 0 1 270
box -6 -8 86 268
use NAND3X1  _1091_
timestamp 0
transform -1 0 4210 0 -1 270
box -6 -8 86 268
use NAND3X1  _1092_
timestamp 0
transform -1 0 3630 0 -1 270
box -6 -8 86 268
use NAND2X1  _1093_
timestamp 0
transform 1 0 3430 0 -1 270
box -6 -8 66 268
use XOR2X1  _1094_
timestamp 0
transform 1 0 1850 0 -1 1310
box -6 -8 126 268
use NAND2X1  _1095_
timestamp 0
transform 1 0 2190 0 -1 2870
box -6 -8 66 268
use OAI21X1  _1096_
timestamp 0
transform 1 0 2050 0 -1 2870
box -6 -8 86 268
use NAND2X1  _1097_
timestamp 0
transform 1 0 3810 0 -1 5470
box -6 -8 66 268
use NAND2X1  _1098_
timestamp 0
transform -1 0 3230 0 -1 270
box -6 -8 66 268
use NAND2X1  _1099_
timestamp 0
transform -1 0 3630 0 1 270
box -6 -8 66 268
use OAI21X1  _1100_
timestamp 0
transform 1 0 3450 0 -1 2350
box -6 -8 86 268
use AOI21X1  _1101_
timestamp 0
transform -1 0 4170 0 1 270
box -6 -8 86 268
use OAI21X1  _1102_
timestamp 0
transform 1 0 3950 0 1 270
box -6 -8 86 268
use NAND2X1  _1103_
timestamp 0
transform 1 0 3910 0 -1 790
box -6 -8 66 268
use INVX1  _1104_
timestamp 0
transform -1 0 5790 0 -1 270
box -6 -8 46 268
use INVX1  _1105_
timestamp 0
transform -1 0 5290 0 -1 270
box -6 -8 46 268
use AOI21X1  _1106_
timestamp 0
transform 1 0 5110 0 -1 270
box -6 -8 86 268
use INVX2  _1107_
timestamp 0
transform 1 0 4290 0 1 1830
box -6 -8 46 268
use NOR2X1  _1108_
timestamp 0
transform -1 0 4530 0 -1 1830
box -6 -8 66 268
use AND2X2  _1109_
timestamp 0
transform 1 0 5290 0 1 1310
box -6 -8 86 268
use AOI22X1  _1110_
timestamp 0
transform 1 0 5110 0 1 1310
box -6 -8 106 268
use AOI21X1  _1111_
timestamp 0
transform 1 0 5430 0 1 1310
box -6 -8 86 268
use XNOR2X1  _1112_
timestamp 0
transform -1 0 5810 0 -1 1310
box -6 -8 126 268
use AOI21X1  _1113_
timestamp 0
transform 1 0 4710 0 1 790
box -6 -8 86 268
use NAND2X1  _1114_
timestamp 0
transform 1 0 4530 0 1 1310
box -6 -8 66 268
use NAND2X1  _1115_
timestamp 0
transform 1 0 4590 0 -1 1830
box -6 -8 66 268
use NAND2X1  _1116_
timestamp 0
transform 1 0 4410 0 1 1310
box -6 -8 66 268
use OAI21X1  _1117_
timestamp 0
transform 1 0 4270 0 1 1310
box -6 -8 86 268
use OAI21X1  _1118_
timestamp 0
transform 1 0 4650 0 1 1310
box -6 -8 86 268
use NOR2X1  _1119_
timestamp 0
transform -1 0 5450 0 1 790
box -6 -8 66 268
use OAI21X1  _1120_
timestamp 0
transform 1 0 4590 0 -1 1310
box -6 -8 86 268
use XOR2X1  _1121_
timestamp 0
transform -1 0 4910 0 1 1310
box -6 -8 126 268
use NOR2X1  _1122_
timestamp 0
transform -1 0 5290 0 -1 1310
box -6 -8 66 268
use OAI21X1  _1123_
timestamp 0
transform 1 0 5650 0 1 790
box -6 -8 86 268
use XOR2X1  _1124_
timestamp 0
transform -1 0 5630 0 -1 1310
box -6 -8 126 268
use OAI21X1  _1125_
timestamp 0
transform 1 0 5090 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1126_
timestamp 0
transform -1 0 5330 0 1 790
box -6 -8 66 268
use NAND3X1  _1127_
timestamp 0
transform 1 0 5450 0 -1 790
box -6 -8 86 268
use NAND3X1  _1128_
timestamp 0
transform -1 0 5690 0 -1 270
box -6 -8 86 268
use AOI21X1  _1129_
timestamp 0
transform -1 0 4410 0 -1 790
box -6 -8 86 268
use OAI21X1  _1130_
timestamp 0
transform 1 0 5190 0 1 270
box -6 -8 86 268
use AOI21X1  _1131_
timestamp 0
transform -1 0 5390 0 -1 790
box -6 -8 86 268
use NAND2X1  _1132_
timestamp 0
transform -1 0 4930 0 1 790
box -6 -8 66 268
use OAI21X1  _1133_
timestamp 0
transform 1 0 4990 0 1 790
box -6 -8 86 268
use AOI21X1  _1134_
timestamp 0
transform 1 0 5130 0 1 790
box -6 -8 86 268
use OAI21X1  _1135_
timestamp 0
transform 1 0 5170 0 -1 790
box -6 -8 86 268
use NAND3X1  _1136_
timestamp 0
transform -1 0 5550 0 -1 270
box -6 -8 86 268
use NAND3X1  _1137_
timestamp 0
transform -1 0 5670 0 -1 790
box -6 -8 86 268
use OAI21X1  _1138_
timestamp 0
transform -1 0 5110 0 -1 790
box -6 -8 86 268
use NAND3X1  _1139_
timestamp 0
transform 1 0 4890 0 -1 790
box -6 -8 86 268
use NAND3X1  _1140_
timestamp 0
transform 1 0 5050 0 1 270
box -6 -8 86 268
use INVX1  _1141_
timestamp 0
transform 1 0 4930 0 1 270
box -6 -8 46 268
use AOI21X1  _1142_
timestamp 0
transform -1 0 4830 0 -1 790
box -6 -8 86 268
use AOI21X1  _1143_
timestamp 0
transform -1 0 5410 0 1 270
box -6 -8 86 268
use OAI21X1  _1144_
timestamp 0
transform -1 0 4690 0 -1 790
box -6 -8 86 268
use NAND2X1  _1145_
timestamp 0
transform -1 0 4350 0 1 2870
box -6 -8 66 268
use XOR2X1  _1146_
timestamp 0
transform 1 0 4230 0 -1 3390
box -6 -8 126 268
use OAI21X1  _1147_
timestamp 0
transform -1 0 3910 0 1 4950
box -6 -8 86 268
use INVX1  _1148_
timestamp 0
transform 1 0 4050 0 1 2870
box -6 -8 46 268
use AOI21X1  _1149_
timestamp 0
transform -1 0 4230 0 1 2870
box -6 -8 86 268
use AOI22X1  _1150_
timestamp 0
transform 1 0 5570 0 1 1310
box -6 -8 106 268
use INVX1  _1151_
timestamp 0
transform 1 0 5670 0 -1 1830
box -6 -8 46 268
use OAI21X1  _1152_
timestamp 0
transform -1 0 5430 0 -1 1310
box -6 -8 86 268
use NOR2X1  _1153_
timestamp 0
transform 1 0 4390 0 -1 2350
box -6 -8 66 268
use NAND2X1  _1154_
timestamp 0
transform 1 0 4170 0 1 1830
box -6 -8 66 268
use NAND2X1  _1155_
timestamp 0
transform 1 0 4530 0 -1 2350
box -6 -8 66 268
use OR2X2  _1156_
timestamp 0
transform 1 0 4650 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1157_
timestamp 0
transform 1 0 4250 0 -1 2350
box -6 -8 86 268
use NAND3X1  _1158_
timestamp 0
transform 1 0 4790 0 -1 2350
box -6 -8 86 268
use NAND2X1  _1159_
timestamp 0
transform -1 0 5290 0 -1 2350
box -6 -8 66 268
use NAND2X1  _1160_
timestamp 0
transform -1 0 4530 0 -1 2870
box -6 -8 66 268
use OAI21X1  _1161_
timestamp 0
transform -1 0 5010 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1162_
timestamp 0
transform 1 0 4410 0 1 1830
box -6 -8 86 268
use NAND2X1  _1163_
timestamp 0
transform -1 0 4610 0 1 1830
box -6 -8 66 268
use OAI21X1  _1164_
timestamp 0
transform 1 0 4830 0 -1 1830
box -6 -8 86 268
use NOR2X1  _1165_
timestamp 0
transform 1 0 4710 0 -1 1830
box -6 -8 66 268
use NAND3X1  _1166_
timestamp 0
transform 1 0 4810 0 1 1830
box -6 -8 86 268
use NAND3X1  _1167_
timestamp 0
transform 1 0 5350 0 1 1830
box -6 -8 86 268
use AOI21X1  _1168_
timestamp 0
transform -1 0 5590 0 1 790
box -6 -8 86 268
use AOI21X1  _1169_
timestamp 0
transform 1 0 4670 0 1 1830
box -6 -8 86 268
use INVX1  _1170_
timestamp 0
transform 1 0 4970 0 1 1830
box -6 -8 46 268
use OAI21X1  _1171_
timestamp 0
transform 1 0 5210 0 1 1830
box -6 -8 86 268
use NAND3X1  _1172_
timestamp 0
transform -1 0 5570 0 1 1830
box -6 -8 86 268
use NAND3X1  _1173_
timestamp 0
transform 1 0 5390 0 -1 1830
box -6 -8 86 268
use OAI21X1  _1174_
timestamp 0
transform 1 0 5070 0 1 1830
box -6 -8 86 268
use NAND3X1  _1175_
timestamp 0
transform -1 0 5610 0 -1 1830
box -6 -8 86 268
use NAND2X1  _1176_
timestamp 0
transform 1 0 5130 0 -1 1830
box -6 -8 66 268
use NAND3X1  _1177_
timestamp 0
transform -1 0 5070 0 -1 1830
box -6 -8 86 268
use AOI21X1  _1178_
timestamp 0
transform -1 0 5690 0 1 270
box -6 -8 86 268
use OAI21X1  _1179_
timestamp 0
transform -1 0 5550 0 1 270
box -6 -8 86 268
use NAND3X1  _1180_
timestamp 0
transform -1 0 5330 0 -1 1830
box -6 -8 86 268
use AND2X2  _1181_
timestamp 0
transform -1 0 4610 0 1 2870
box -6 -8 86 268
use XOR2X1  _1182_
timestamp 0
transform -1 0 4170 0 -1 3390
box -6 -8 126 268
use NAND2X1  _1183_
timestamp 0
transform -1 0 4050 0 1 3910
box -6 -8 66 268
use OAI21X1  _1184_
timestamp 0
transform 1 0 3910 0 -1 3910
box -6 -8 86 268
use INVX1  _1185_
timestamp 0
transform -1 0 5050 0 -1 4430
box -6 -8 46 268
use NAND2X1  _1186_
timestamp 0
transform 1 0 4670 0 1 2870
box -6 -8 66 268
use NOR2X1  _1187_
timestamp 0
transform -1 0 4470 0 1 2870
box -6 -8 66 268
use NAND2X1  _1188_
timestamp 0
transform -1 0 4970 0 1 2870
box -6 -8 66 268
use NAND2X1  _1189_
timestamp 0
transform 1 0 4790 0 1 2870
box -6 -8 66 268
use INVX1  _1190_
timestamp 0
transform -1 0 4590 0 -1 3390
box -6 -8 46 268
use AOI21X1  _1191_
timestamp 0
transform 1 0 4410 0 -1 3390
box -6 -8 86 268
use NAND2X1  _1192_
timestamp 0
transform 1 0 5650 0 -1 4950
box -6 -8 66 268
use OAI21X1  _1193_
timestamp 0
transform -1 0 5170 0 -1 2350
box -6 -8 86 268
use INVX1  _1194_
timestamp 0
transform 1 0 5490 0 1 2350
box -6 -8 46 268
use OR2X2  _1195_
timestamp 0
transform 1 0 4970 0 1 1310
box -6 -8 86 268
use NOR2X1  _1196_
timestamp 0
transform -1 0 4690 0 1 2350
box -6 -8 66 268
use OAI21X1  _1197_
timestamp 0
transform 1 0 4370 0 1 2350
box -6 -8 86 268
use NAND2X1  _1198_
timestamp 0
transform 1 0 4750 0 1 2350
box -6 -8 66 268
use OAI21X1  _1199_
timestamp 0
transform -1 0 4950 0 1 2350
box -6 -8 86 268
use XOR2X1  _1200_
timestamp 0
transform 1 0 5310 0 1 2350
box -6 -8 126 268
use AOI21X1  _1201_
timestamp 0
transform 1 0 5490 0 -1 2350
box -6 -8 86 268
use NAND3X1  _1202_
timestamp 0
transform 1 0 5350 0 -1 2350
box -6 -8 86 268
use INVX1  _1203_
timestamp 0
transform -1 0 5770 0 1 2350
box -6 -8 46 268
use OAI21X1  _1204_
timestamp 0
transform -1 0 5670 0 1 2350
box -6 -8 86 268
use INVX1  _1205_
timestamp 0
transform -1 0 5770 0 -1 790
box -6 -8 46 268
use NAND3X1  _1206_
timestamp 0
transform 1 0 5730 0 1 1310
box -6 -8 86 268
use AND2X2  _1207_
timestamp 0
transform -1 0 5710 0 1 1830
box -6 -8 86 268
use NAND2X1  _1208_
timestamp 0
transform 1 0 5730 0 1 2870
box -6 -8 66 268
use OR2X2  _1209_
timestamp 0
transform -1 0 5650 0 1 2870
box -6 -8 86 268
use NAND2X1  _1210_
timestamp 0
transform -1 0 5510 0 -1 3390
box -6 -8 66 268
use NAND2X1  _1211_
timestamp 0
transform -1 0 5250 0 1 3390
box -6 -8 66 268
use AND2X2  _1212_
timestamp 0
transform -1 0 3370 0 -1 270
box -6 -8 86 268
use NAND3X1  _1213_
timestamp 0
transform 1 0 3030 0 -1 270
box -6 -8 86 268
use NAND3X1  _1214_
timestamp 0
transform -1 0 3990 0 1 2870
box -6 -8 86 268
use AOI21X1  _1215_
timestamp 0
transform 1 0 3770 0 1 2870
box -6 -8 86 268
use INVX1  _1216_
timestamp 0
transform -1 0 4990 0 1 3390
box -6 -8 46 268
use OAI21X1  _1217_
timestamp 0
transform 1 0 4810 0 1 3390
box -6 -8 86 268
use NAND3X1  _1218_
timestamp 0
transform -1 0 5130 0 1 3390
box -6 -8 86 268
use OAI21X1  _1219_
timestamp 0
transform 1 0 4970 0 1 3910
box -6 -8 86 268
use NAND2X1  _1220_
timestamp 0
transform -1 0 5170 0 -1 4430
box -6 -8 66 268
use AOI21X1  _1221_
timestamp 0
transform -1 0 5770 0 -1 2870
box -6 -8 86 268
use INVX1  _1222_
timestamp 0
transform 1 0 5190 0 1 2350
box -6 -8 46 268
use OAI22X1  _1223_
timestamp 0
transform 1 0 5030 0 1 2350
box -6 -8 106 268
use OAI21X1  _1224_
timestamp 0
transform 1 0 4730 0 -1 2870
box -6 -8 86 268
use NOR2X1  _1225_
timestamp 0
transform 1 0 4510 0 1 2350
box -6 -8 66 268
use INVX1  _1226_
timestamp 0
transform 1 0 4870 0 -1 2870
box -6 -8 46 268
use OR2X2  _1227_
timestamp 0
transform 1 0 5110 0 -1 2870
box -6 -8 86 268
use AND2X2  _1228_
timestamp 0
transform 1 0 5250 0 -1 2870
box -6 -8 86 268
use XNOR2X1  _1229_
timestamp 0
transform -1 0 5630 0 -1 2870
box -6 -8 126 268
use XOR2X1  _1230_
timestamp 0
transform 1 0 5590 0 -1 3390
box -6 -8 126 268
use INVX1  _1231_
timestamp 0
transform 1 0 5750 0 1 3910
box -6 -8 46 268
use NAND3X1  _1232_
timestamp 0
transform -1 0 5830 0 -1 4430
box -6 -8 86 268
use OAI21X1  _1233_
timestamp 0
transform 1 0 5570 0 1 3390
box -6 -8 86 268
use NAND2X1  _1234_
timestamp 0
transform -1 0 5770 0 1 3390
box -6 -8 66 268
use NAND3X1  _1235_
timestamp 0
transform 1 0 5690 0 -1 3910
box -6 -8 86 268
use NAND2X1  _1236_
timestamp 0
transform 1 0 5230 0 -1 4430
box -6 -8 66 268
use INVX1  _1237_
timestamp 0
transform 1 0 5770 0 -1 4950
box -6 -8 46 268
use NOR2X1  _1238_
timestamp 0
transform -1 0 5510 0 1 2870
box -6 -8 66 268
use AOI21X1  _1239_
timestamp 0
transform -1 0 5370 0 1 2870
box -6 -8 86 268
use NOR2X1  _1240_
timestamp 0
transform -1 0 5410 0 -1 270
box -6 -8 66 268
use NAND3X1  _1241_
timestamp 0
transform -1 0 5390 0 -1 3390
box -6 -8 86 268
use OAI21X1  _1242_
timestamp 0
transform -1 0 5250 0 -1 3390
box -6 -8 86 268
use NAND2X1  _1243_
timestamp 0
transform 1 0 5390 0 -1 2870
box -6 -8 66 268
use OAI21X1  _1244_
timestamp 0
transform 1 0 4590 0 -1 2870
box -6 -8 86 268
use OR2X2  _1245_
timestamp 0
transform 1 0 4970 0 -1 2870
box -6 -8 86 268
use INVX1  _1246_
timestamp 0
transform 1 0 5190 0 1 2870
box -6 -8 46 268
use OAI21X1  _1247_
timestamp 0
transform -1 0 5110 0 1 2870
box -6 -8 86 268
use AND2X2  _1248_
timestamp 0
transform 1 0 5030 0 -1 3390
box -6 -8 86 268
use NOR2X1  _1249_
timestamp 0
transform -1 0 5490 0 -1 3910
box -6 -8 66 268
use INVX1  _1250_
timestamp 0
transform -1 0 4690 0 -1 3390
box -6 -8 46 268
use OAI21X1  _1251_
timestamp 0
transform 1 0 4890 0 -1 3390
box -6 -8 86 268
use AOI21X1  _1252_
timestamp 0
transform 1 0 4750 0 -1 3390
box -6 -8 86 268
use INVX1  _1253_
timestamp 0
transform -1 0 5510 0 1 3390
box -6 -8 46 268
use OAI21X1  _1254_
timestamp 0
transform -1 0 5390 0 1 3390
box -6 -8 86 268
use OAI22X1  _1255_
timestamp 0
transform -1 0 5450 0 -1 4430
box -6 -8 106 268
use INVX1  _1256_
timestamp 0
transform -1 0 5250 0 -1 4950
box -6 -8 46 268
use AOI21X1  _1257_
timestamp 0
transform 1 0 5290 0 -1 3910
box -6 -8 86 268
use AND2X2  _1258_
timestamp 0
transform 1 0 5150 0 -1 3910
box -6 -8 86 268
use AOI22X1  _1259_
timestamp 0
transform 1 0 5110 0 1 3910
box -6 -8 106 268
use NOR2X1  _1260_
timestamp 0
transform -1 0 250 0 1 4430
box -6 -8 66 268
use INVX1  _1261_
timestamp 0
transform 1 0 90 0 1 4430
box -6 -8 46 268
use NAND2X1  _1262_
timestamp 0
transform 1 0 310 0 1 4430
box -6 -8 66 268
use NAND2X1  _1263_
timestamp 0
transform -1 0 490 0 1 4430
box -6 -8 66 268
use NAND2X1  _1264_
timestamp 0
transform -1 0 1110 0 1 4430
box -6 -8 66 268
use OAI21X1  _1265_
timestamp 0
transform 1 0 550 0 1 4430
box -6 -8 86 268
use INVX1  _1266_
timestamp 0
transform -1 0 870 0 -1 4950
box -6 -8 46 268
use NOR2X1  _1267_
timestamp 0
transform 1 0 570 0 -1 4950
box -6 -8 66 268
use NOR2X1  _1268_
timestamp 0
transform 1 0 370 0 1 4950
box -6 -8 66 268
use NOR2X1  _1269_
timestamp 0
transform -1 0 250 0 -1 4950
box -6 -8 66 268
use NAND2X1  _1270_
timestamp 0
transform 1 0 70 0 -1 4950
box -6 -8 66 268
use OAI21X1  _1271_
timestamp 0
transform 1 0 310 0 -1 4950
box -6 -8 86 268
use NAND2X1  _1272_
timestamp 0
transform 1 0 450 0 -1 4950
box -6 -8 66 268
use NAND2X1  _1273_
timestamp 0
transform 1 0 870 0 1 4950
box -6 -8 66 268
use OAI21X1  _1274_
timestamp 0
transform 1 0 490 0 1 4950
box -6 -8 86 268
use OAI21X1  _1275_
timestamp 0
transform -1 0 770 0 -1 4950
box -6 -8 86 268
use XOR2X1  _1276_
timestamp 0
transform -1 0 1990 0 -1 3390
box -6 -8 126 268
use XNOR2X1  _1277_
timestamp 0
transform 1 0 1650 0 1 3390
box -6 -8 126 268
use NAND2X1  _1278_
timestamp 0
transform 1 0 2070 0 -1 3910
box -6 -8 66 268
use OAI21X1  _1279_
timestamp 0
transform 1 0 1770 0 -1 3910
box -6 -8 86 268
use NOR2X1  _1280_
timestamp 0
transform -1 0 2030 0 1 3390
box -6 -8 66 268
use AOI21X1  _1281_
timestamp 0
transform 1 0 1830 0 1 3390
box -6 -8 86 268
use NOR2X1  _1282_
timestamp 0
transform 1 0 310 0 -1 2870
box -6 -8 66 268
use NOR2X1  _1283_
timestamp 0
transform -1 0 610 0 1 2870
box -6 -8 66 268
use NOR2X1  _1284_
timestamp 0
transform 1 0 710 0 -1 3390
box -6 -8 66 268
use XOR2X1  _1285_
timestamp 0
transform -1 0 950 0 -1 3390
box -6 -8 126 268
use NAND2X1  _1286_
timestamp 0
transform -1 0 1570 0 -1 3910
box -6 -8 66 268
use OAI21X1  _1287_
timestamp 0
transform 1 0 1370 0 -1 3910
box -6 -8 86 268
use NAND2X1  _1288_
timestamp 0
transform -1 0 290 0 1 4950
box -6 -8 66 268
use NAND2X1  _1289_
timestamp 0
transform -1 0 130 0 -1 3910
box -6 -8 66 268
use NAND2X1  _1290_
timestamp 0
transform 1 0 70 0 -1 3390
box -6 -8 66 268
use AND2X2  _1291_
timestamp 0
transform 1 0 90 0 1 3910
box -6 -8 86 268
use INVX1  _1292_
timestamp 0
transform 1 0 350 0 1 3910
box -6 -8 46 268
use INVX1  _1293_
timestamp 0
transform -1 0 650 0 -1 3390
box -6 -8 46 268
use OAI21X1  _1294_
timestamp 0
transform 1 0 470 0 -1 3390
box -6 -8 86 268
use INVX1  _1295_
timestamp 0
transform -1 0 230 0 -1 4430
box -6 -8 46 268
use NAND2X1  _1296_
timestamp 0
transform -1 0 130 0 -1 4430
box -6 -8 66 268
use NAND2X1  _1297_
timestamp 0
transform 1 0 230 0 1 3910
box -6 -8 66 268
use NAND2X1  _1298_
timestamp 0
transform -1 0 350 0 -1 4430
box -6 -8 66 268
use OAI21X1  _1299_
timestamp 0
transform 1 0 90 0 1 4950
box -6 -8 86 268
use NAND2X1  _1300_
timestamp 0
transform -1 0 750 0 1 4430
box -6 -8 66 268
use OAI21X1  _1301_
timestamp 0
transform 1 0 190 0 -1 3910
box -6 -8 86 268
use OR2X2  _1302_
timestamp 0
transform -1 0 790 0 1 3910
box -6 -8 86 268
use NAND2X1  _1303_
timestamp 0
transform -1 0 910 0 1 3910
box -6 -8 66 268
use AND2X2  _1304_
timestamp 0
transform 1 0 570 0 1 3910
box -6 -8 86 268
use NOR2X1  _1305_
timestamp 0
transform -1 0 470 0 -1 4430
box -6 -8 66 268
use INVX1  _1306_
timestamp 0
transform 1 0 350 0 -1 3910
box -6 -8 46 268
use INVX1  _1307_
timestamp 0
transform -1 0 710 0 -1 4430
box -6 -8 46 268
use OAI21X1  _1308_
timestamp 0
transform -1 0 670 0 -1 3910
box -6 -8 86 268
use OAI21X1  _1309_
timestamp 0
transform -1 0 610 0 -1 4430
box -6 -8 86 268
use NAND2X1  _1310_
timestamp 0
transform -1 0 1590 0 1 3390
box -6 -8 66 268
use OAI21X1  _1311_
timestamp 0
transform 1 0 730 0 -1 3910
box -6 -8 86 268
use XOR2X1  _1312_
timestamp 0
transform 1 0 890 0 -1 2870
box -6 -8 126 268
use NOR2X1  _1313_
timestamp 0
transform -1 0 1070 0 -1 3390
box -6 -8 66 268
use NAND2X1  _1314_
timestamp 0
transform -1 0 1010 0 1 2870
box -6 -8 66 268
use NAND2X1  _1315_
timestamp 0
transform 1 0 1070 0 1 2870
box -6 -8 66 268
use OAI21X1  _1316_
timestamp 0
transform 1 0 1290 0 -1 3390
box -6 -8 86 268
use OAI21X1  _1317_
timestamp 0
transform -1 0 1270 0 1 2870
box -6 -8 86 268
use NOR2X1  _1318_
timestamp 0
transform 1 0 1690 0 -1 2870
box -6 -8 66 268
use NAND2X1  _1319_
timestamp 0
transform -1 0 1630 0 -1 2870
box -6 -8 66 268
use INVX1  _1320_
timestamp 0
transform 1 0 1330 0 -1 2870
box -6 -8 46 268
use NOR2X1  _1321_
timestamp 0
transform -1 0 1510 0 -1 2870
box -6 -8 66 268
use XNOR2X1  _1322_
timestamp 0
transform 1 0 1670 0 -1 3390
box -6 -8 126 268
use NAND2X1  _1323_
timestamp 0
transform 1 0 2330 0 -1 3910
box -6 -8 66 268
use OAI21X1  _1324_
timestamp 0
transform 1 0 2190 0 -1 3910
box -6 -8 86 268
use NAND2X1  _1325_
timestamp 0
transform -1 0 1770 0 1 4950
box -6 -8 66 268
use OAI21X1  _1326_
timestamp 0
transform 1 0 450 0 -1 3910
box -6 -8 86 268
use NAND2X1  _1327_
timestamp 0
transform -1 0 1130 0 -1 2870
box -6 -8 66 268
use OAI21X1  _1328_
timestamp 0
transform 1 0 1190 0 -1 2870
box -6 -8 86 268
use AND2X2  _1329_
timestamp 0
transform -1 0 1230 0 -1 3390
box -6 -8 86 268
use AOI21X1  _1330_
timestamp 0
transform 1 0 1030 0 1 3390
box -6 -8 86 268
use NOR2X1  _1331_
timestamp 0
transform -1 0 510 0 1 3910
box -6 -8 66 268
use NAND3X1  _1332_
timestamp 0
transform 1 0 890 0 1 3390
box -6 -8 86 268
use NAND2X1  _1333_
timestamp 0
transform 1 0 1170 0 1 3390
box -6 -8 66 268
use OR2X2  _1334_
timestamp 0
transform -1 0 2130 0 -1 5470
box -6 -8 86 268
use NAND2X1  _1335_
timestamp 0
transform 1 0 1770 0 -1 5470
box -6 -8 66 268
use AND2X2  _1336_
timestamp 0
transform -1 0 1990 0 -1 5470
box -6 -8 86 268
use NOR2X1  _1337_
timestamp 0
transform -1 0 1890 0 1 4950
box -6 -8 66 268
use INVX1  _1338_
timestamp 0
transform 1 0 1430 0 -1 4950
box -6 -8 46 268
use INVX1  _1339_
timestamp 0
transform 1 0 1950 0 1 4950
box -6 -8 46 268
use OAI21X1  _1340_
timestamp 0
transform -1 0 1610 0 -1 4950
box -6 -8 86 268
use OAI21X1  _1341_
timestamp 0
transform -1 0 1650 0 1 4950
box -6 -8 86 268
use OAI21X1  _1342_
timestamp 0
transform 1 0 1670 0 -1 4950
box -6 -8 86 268
use NOR2X1  _1343_
timestamp 0
transform 1 0 1910 0 1 4430
box -6 -8 66 268
use NAND2X1  _1344_
timestamp 0
transform -1 0 2110 0 1 4430
box -6 -8 66 268
use INVX1  _1345_
timestamp 0
transform -1 0 1490 0 1 4430
box -6 -8 46 268
use NOR2X1  _1346_
timestamp 0
transform -1 0 1610 0 1 4430
box -6 -8 66 268
use INVX1  _1347_
timestamp 0
transform 1 0 1670 0 1 4430
box -6 -8 46 268
use XOR2X1  _1348_
timestamp 0
transform 1 0 1950 0 -1 4950
box -6 -8 126 268
use NAND2X1  _1349_
timestamp 0
transform 1 0 3110 0 1 4950
box -6 -8 66 268
use OAI21X1  _1350_
timestamp 0
transform 1 0 2970 0 1 4950
box -6 -8 86 268
use NAND2X1  _1351_
timestamp 0
transform 1 0 2410 0 1 4430
box -6 -8 66 268
use NOR2X1  _1352_
timestamp 0
transform -1 0 1890 0 -1 4950
box -6 -8 66 268
use OAI21X1  _1353_
timestamp 0
transform 1 0 1770 0 1 4430
box -6 -8 86 268
use AOI21X1  _1354_
timestamp 0
transform 1 0 1870 0 -1 4430
box -6 -8 86 268
use NOR2X1  _1355_
timestamp 0
transform 1 0 4790 0 1 4430
box -6 -8 66 268
use NOR2X1  _1356_
timestamp 0
transform 1 0 4870 0 -1 4430
box -6 -8 66 268
use NOR2X1  _1357_
timestamp 0
transform -1 0 4730 0 1 4430
box -6 -8 66 268
use INVX1  _1358_
timestamp 0
transform -1 0 4330 0 1 4430
box -6 -8 46 268
use AND2X2  _1359_
timestamp 0
transform -1 0 2910 0 1 4430
box -6 -8 86 268
use OAI21X1  _1360_
timestamp 0
transform -1 0 2750 0 1 4430
box -6 -8 86 268
use OAI21X1  _1361_
timestamp 0
transform -1 0 2610 0 1 4430
box -6 -8 86 268
use NOR2X1  _1362_
timestamp 0
transform -1 0 3930 0 1 4430
box -6 -8 66 268
use NOR2X1  _1363_
timestamp 0
transform -1 0 4050 0 1 4430
box -6 -8 66 268
use NOR2X1  _1364_
timestamp 0
transform -1 0 5490 0 1 4430
box -6 -8 66 268
use NAND2X1  _1365_
timestamp 0
transform -1 0 5710 0 1 4430
box -6 -8 66 268
use INVX1  _1366_
timestamp 0
transform 1 0 5550 0 1 4430
box -6 -8 46 268
use NOR2X1  _1367_
timestamp 0
transform 1 0 5070 0 1 4430
box -6 -8 66 268
use XOR2X1  _1368_
timestamp 0
transform 1 0 4110 0 1 4430
box -6 -8 126 268
use NAND2X1  _1369_
timestamp 0
transform -1 0 3470 0 -1 3910
box -6 -8 66 268
use OAI21X1  _1370_
timestamp 0
transform -1 0 3850 0 -1 3910
box -6 -8 86 268
use NAND2X1  _1371_
timestamp 0
transform -1 0 4030 0 1 4950
box -6 -8 66 268
use AOI21X1  _1372_
timestamp 0
transform -1 0 4990 0 1 4430
box -6 -8 86 268
use NAND2X1  _1373_
timestamp 0
transform -1 0 4450 0 1 4430
box -6 -8 66 268
use OAI21X1  _1374_
timestamp 0
transform 1 0 4530 0 1 4430
box -6 -8 86 268
use NAND2X1  _1375_
timestamp 0
transform -1 0 5730 0 -1 5470
box -6 -8 66 268
use NOR2X1  _1376_
timestamp 0
transform 1 0 5550 0 -1 5470
box -6 -8 66 268
use INVX1  _1377_
timestamp 0
transform -1 0 5350 0 -1 5470
box -6 -8 46 268
use AND2X2  _1378_
timestamp 0
transform 1 0 5410 0 -1 5470
box -6 -8 86 268
use NOR2X1  _1379_
timestamp 0
transform -1 0 4530 0 1 4950
box -6 -8 66 268
use INVX1  _1380_
timestamp 0
transform 1 0 4590 0 1 4950
box -6 -8 46 268
use INVX1  _1381_
timestamp 0
transform -1 0 4890 0 1 4950
box -6 -8 46 268
use OAI21X1  _1382_
timestamp 0
transform -1 0 4790 0 1 4950
box -6 -8 86 268
use OAI21X1  _1383_
timestamp 0
transform -1 0 4410 0 1 4950
box -6 -8 86 268
use OAI21X1  _1384_
timestamp 0
transform 1 0 5170 0 -1 5470
box -6 -8 86 268
use NOR2X1  _1385_
timestamp 0
transform 1 0 5310 0 1 4950
box -6 -8 66 268
use NOR2X1  _1386_
timestamp 0
transform 1 0 5090 0 -1 4950
box -6 -8 66 268
use NOR2X1  _1387_
timestamp 0
transform -1 0 5250 0 1 4950
box -6 -8 66 268
use INVX1  _1388_
timestamp 0
transform -1 0 4990 0 1 4950
box -6 -8 46 268
use OR2X2  _1389_
timestamp 0
transform 1 0 5030 0 -1 5470
box -6 -8 86 268
use AOI21X1  _1390_
timestamp 0
transform -1 0 4950 0 -1 5470
box -6 -8 86 268
use AOI22X1  _1391_
timestamp 0
transform 1 0 4710 0 -1 5470
box -6 -8 106 268
use AOI21X1  _1392_
timestamp 0
transform -1 0 5130 0 1 4950
box -6 -8 86 268
use INVX1  _1393_
timestamp 0
transform -1 0 4530 0 -1 4950
box -6 -8 46 268
use NOR2X1  _1394_
timestamp 0
transform -1 0 4790 0 -1 4950
box -6 -8 66 268
use AOI21X1  _1395_
timestamp 0
transform -1 0 4430 0 -1 4950
box -6 -8 86 268
use INVX1  _1396_
timestamp 0
transform 1 0 3130 0 -1 4950
box -6 -8 46 268
use NOR2X1  _1397_
timestamp 0
transform -1 0 3310 0 -1 4950
box -6 -8 66 268
use OAI21X1  _1398_
timestamp 0
transform -1 0 3070 0 -1 4950
box -6 -8 86 268
use OAI22X1  _1399_
timestamp 0
transform 1 0 2830 0 -1 4950
box -6 -8 106 268
use NAND2X1  _1400_
timestamp 0
transform 1 0 3350 0 1 4430
box -6 -8 66 268
use NAND3X1  _1401_
timestamp 0
transform 1 0 3370 0 -1 4950
box -6 -8 86 268
use OAI21X1  _1402_
timestamp 0
transform -1 0 3710 0 -1 4950
box -6 -8 86 268
use NAND2X1  _1403_
timestamp 0
transform -1 0 3570 0 -1 4950
box -6 -8 66 268
use OAI21X1  _1404_
timestamp 0
transform -1 0 3570 0 1 4430
box -6 -8 86 268
use INVX1  _1405_
timestamp 0
transform -1 0 4650 0 -1 5470
box -6 -8 46 268
use NAND3X1  _1406_
timestamp 0
transform 1 0 3090 0 1 3910
box -6 -8 86 268
use NAND2X1  _1407_
timestamp 0
transform -1 0 4850 0 -1 3910
box -6 -8 66 268
use OAI21X1  _1408_
timestamp 0
transform 1 0 4650 0 -1 3910
box -6 -8 86 268
use INVX1  _1409_
timestamp 0
transform -1 0 4550 0 -1 5470
box -6 -8 46 268
use NAND2X1  _1410_
timestamp 0
transform -1 0 4110 0 -1 4430
box -6 -8 66 268
use OAI21X1  _1411_
timestamp 0
transform 1 0 3910 0 -1 4430
box -6 -8 86 268
use INVX1  _1412_
timestamp 0
transform 1 0 3470 0 -1 5470
box -6 -8 46 268
use NAND2X1  _1413_
timestamp 0
transform 1 0 3370 0 1 3910
box -6 -8 66 268
use OAI21X1  _1414_
timestamp 0
transform 1 0 3230 0 1 3910
box -6 -8 86 268
use INVX1  _1415_
timestamp 0
transform 1 0 3250 0 1 4430
box -6 -8 46 268
use NAND2X1  _1416_
timestamp 0
transform 1 0 4570 0 1 3390
box -6 -8 66 268
use OAI21X1  _1417_
timestamp 0
transform 1 0 4070 0 1 3390
box -6 -8 86 268
use NOR2X1  _1418_
timestamp 0
transform -1 0 2530 0 1 4950
box -6 -8 66 268
use NOR2X1  _1419_
timestamp 0
transform 1 0 2550 0 -1 5470
box -6 -8 66 268
use AOI21X1  _1420_
timestamp 0
transform -1 0 2770 0 -1 5470
box -6 -8 86 268
use NOR2X1  _1421_
timestamp 0
transform -1 0 2510 0 1 3910
box -6 -8 66 268
use AOI21X1  _1422_
timestamp 0
transform 1 0 2570 0 1 3910
box -6 -8 86 268
use NOR2X1  _1423_
timestamp 0
transform -1 0 3710 0 -1 4430
box -6 -8 66 268
use AOI21X1  _1424_
timestamp 0
transform 1 0 3270 0 -1 4430
box -6 -8 86 268
use NOR2X1  _1425_
timestamp 0
transform -1 0 3930 0 1 3910
box -6 -8 66 268
use AOI21X1  _1426_
timestamp 0
transform 1 0 3730 0 1 3910
box -6 -8 86 268
use INVX1  _1427_
timestamp 0
transform -1 0 2970 0 1 2870
box -6 -8 46 268
use OAI21X1  _1428_
timestamp 0
transform -1 0 3510 0 -1 3390
box -6 -8 86 268
use OAI21X1  _1429_
timestamp 0
transform 1 0 3290 0 -1 3390
box -6 -8 86 268
use OAI21X1  _1430_
timestamp 0
transform -1 0 2850 0 -1 3390
box -6 -8 86 268
use OAI21X1  _1431_
timestamp 0
transform -1 0 2990 0 -1 3390
box -6 -8 86 268
use OAI21X1  _1432_
timestamp 0
transform -1 0 2710 0 1 2870
box -6 -8 86 268
use OAI21X1  _1433_
timestamp 0
transform -1 0 2850 0 1 2870
box -6 -8 86 268
use OAI21X1  _1434_
timestamp 0
transform -1 0 3110 0 1 2870
box -6 -8 86 268
use OAI21X1  _1435_
timestamp 0
transform -1 0 3270 0 1 2870
box -6 -8 86 268
use NOR2X1  _1436_
timestamp 0
transform 1 0 3190 0 1 3390
box -6 -8 66 268
use AOI21X1  _1437_
timestamp 0
transform -1 0 3630 0 1 3390
box -6 -8 86 268
use NOR2X1  _1438_
timestamp 0
transform -1 0 1230 0 -1 4950
box -6 -8 66 268
use AOI21X1  _1439_
timestamp 0
transform -1 0 1370 0 -1 4950
box -6 -8 86 268
use NOR2X1  _1440_
timestamp 0
transform -1 0 3870 0 1 3390
box -6 -8 66 268
use AOI21X1  _1441_
timestamp 0
transform -1 0 4010 0 1 3390
box -6 -8 86 268
use NOR2X1  _1442_
timestamp 0
transform -1 0 3410 0 1 2870
box -6 -8 66 268
use AOI21X1  _1443_
timestamp 0
transform 1 0 3470 0 1 2870
box -6 -8 86 268
use NAND2X1  _1444_
timestamp 0
transform 1 0 2690 0 1 2350
box -6 -8 66 268
use OAI21X1  _1445_
timestamp 0
transform -1 0 2630 0 1 2350
box -6 -8 86 268
use NAND2X1  _1446_
timestamp 0
transform 1 0 2510 0 -1 2350
box -6 -8 66 268
use OAI21X1  _1447_
timestamp 0
transform 1 0 2370 0 -1 2350
box -6 -8 86 268
use NAND2X1  _1448_
timestamp 0
transform 1 0 3730 0 -1 2350
box -6 -8 66 268
use OAI21X1  _1449_
timestamp 0
transform 1 0 3110 0 1 1830
box -6 -8 86 268
use NAND2X1  _1450_
timestamp 0
transform 1 0 3590 0 1 2350
box -6 -8 66 268
use OAI21X1  _1451_
timestamp 0
transform -1 0 3670 0 -1 2350
box -6 -8 86 268
use DFFPOSX1  _1452_
timestamp 0
transform 1 0 3010 0 1 2350
box -6 -8 246 268
use DFFPOSX1  _1453_
timestamp 0
transform -1 0 3390 0 -1 2350
box -6 -8 246 268
use DFFPOSX1  _1454_
timestamp 0
transform -1 0 3950 0 -1 2870
box -6 -8 246 268
use DFFPOSX1  _1455_
timestamp 0
transform 1 0 3930 0 1 2350
box -6 -8 246 268
use DFFPOSX1  _1456_
timestamp 0
transform -1 0 690 0 1 3390
box -6 -8 246 268
use DFFPOSX1  _1457_
timestamp 0
transform -1 0 590 0 -1 5470
box -6 -8 246 268
use DFFPOSX1  _1458_
timestamp 0
transform -1 0 2230 0 -1 3390
box -6 -8 246 268
use DFFPOSX1  _1459_
timestamp 0
transform 1 0 130 0 1 2870
box -6 -8 246 268
use DFFPOSX1  _1460_
timestamp 0
transform -1 0 350 0 1 3390
box -6 -8 246 268
use DFFPOSX1  _1461_
timestamp 0
transform -1 0 1490 0 1 3910
box -6 -8 246 268
use DFFPOSX1  _1462_
timestamp 0
transform -1 0 1610 0 1 2870
box -6 -8 246 268
use DFFPOSX1  _1463_
timestamp 0
transform -1 0 2590 0 -1 2870
box -6 -8 246 268
use DFFPOSX1  _1464_
timestamp 0
transform 1 0 1110 0 -1 5470
box -6 -8 246 268
use DFFPOSX1  _1465_
timestamp 0
transform -1 0 2290 0 -1 4430
box -6 -8 246 268
use DFFPOSX1  _1466_
timestamp 0
transform 1 0 4670 0 1 3910
box -6 -8 246 268
use DFFPOSX1  _1467_
timestamp 0
transform 1 0 5450 0 1 3910
box -6 -8 246 268
use DFFPOSX1  _1468_
timestamp 0
transform 1 0 5510 0 1 4950
box -6 -8 246 268
use DFFPOSX1  _1469_
timestamp 0
transform 1 0 4790 0 -1 4950
box -6 -8 246 268
use DFFPOSX1  _1470_
timestamp 0
transform 1 0 3410 0 1 4950
box -6 -8 246 268
use DFFPOSX1  _1471_
timestamp 0
transform -1 0 4050 0 -1 4950
box -6 -8 246 268
use DFFPOSX1  _1472_
timestamp 0
transform 1 0 350 0 1 2350
box -6 -8 246 268
use DFFPOSX1  _1473_
timestamp 0
transform -1 0 1310 0 -1 4430
box -6 -8 246 268
use DFFPOSX1  _1474_
timestamp 0
transform 1 0 1770 0 1 2350
box -6 -8 246 268
use DFFPOSX1  _1475_
timestamp 0
transform -1 0 710 0 -1 2870
box -6 -8 246 268
use DFFPOSX1  _1476_
timestamp 0
transform -1 0 350 0 1 2350
box -6 -8 246 268
use DFFPOSX1  _1477_
timestamp 0
transform -1 0 1150 0 1 3910
box -6 -8 246 268
use DFFPOSX1  _1478_
timestamp 0
transform 1 0 830 0 1 2350
box -6 -8 246 268
use DFFPOSX1  _1479_
timestamp 0
transform -1 0 1990 0 -1 2870
box -6 -8 246 268
use DFFPOSX1  _1480_
timestamp 0
transform -1 0 4110 0 -1 5470
box -6 -8 246 268
use DFFPOSX1  _1481_
timestamp 0
transform -1 0 4230 0 -1 3910
box -6 -8 246 268
use DFFPOSX1  _1482_
timestamp 0
transform 1 0 4470 0 -1 4430
box -6 -8 246 268
use DFFPOSX1  _1483_
timestamp 0
transform 1 0 5450 0 -1 4430
box -6 -8 246 268
use DFFPOSX1  _1484_
timestamp 0
transform 1 0 5350 0 -1 4950
box -6 -8 246 268
use DFFPOSX1  _1485_
timestamp 0
transform 1 0 5130 0 1 4430
box -6 -8 246 268
use DFFPOSX1  _1486_
timestamp 0
transform 1 0 750 0 1 4430
box -6 -8 246 268
use DFFPOSX1  _1487_
timestamp 0
transform 1 0 570 0 1 4950
box -6 -8 246 268
use DFFPOSX1  _1488_
timestamp 0
transform 1 0 1630 0 1 3910
box -6 -8 246 268
use DFFPOSX1  _1489_
timestamp 0
transform 1 0 1070 0 -1 3910
box -6 -8 246 268
use DFFPOSX1  _1490_
timestamp 0
transform 1 0 10 0 -1 5470
box -6 -8 246 268
use DFFPOSX1  _1491_
timestamp 0
transform -1 0 950 0 -1 4430
box -6 -8 246 268
use DFFPOSX1  _1492_
timestamp 0
transform 1 0 1370 0 -1 3390
box -6 -8 246 268
use DFFPOSX1  _1493_
timestamp 0
transform -1 0 2270 0 1 3910
box -6 -8 246 268
use DFFPOSX1  _1494_
timestamp 0
transform 1 0 1270 0 1 4950
box -6 -8 246 268
use DFFPOSX1  _1495_
timestamp 0
transform 1 0 2890 0 -1 5470
box -6 -8 246 268
use DFFPOSX1  _1496_
timestamp 0
transform 1 0 2110 0 1 4430
box -6 -8 246 268
use DFFPOSX1  _1497_
timestamp 0
transform -1 0 3710 0 -1 3910
box -6 -8 246 268
use DFFPOSX1  _1498_
timestamp 0
transform -1 0 4270 0 1 4950
box -6 -8 246 268
use DFFPOSX1  _1499_
timestamp 0
transform -1 0 4450 0 -1 5470
box -6 -8 246 268
use DFFPOSX1  _1500_
timestamp 0
transform -1 0 3410 0 1 4950
box -6 -8 246 268
use DFFPOSX1  _1501_
timestamp 0
transform -1 0 3810 0 1 4430
box -6 -8 246 268
use DFFPOSX1  _1502_
timestamp 0
transform 1 0 4850 0 -1 3910
box -6 -8 246 268
use DFFPOSX1  _1503_
timestamp 0
transform -1 0 4350 0 -1 4430
box -6 -8 246 268
use DFFPOSX1  _1504_
timestamp 0
transform 1 0 2850 0 -1 4430
box -6 -8 246 268
use DFFPOSX1  _1505_
timestamp 0
transform 1 0 4150 0 1 3390
box -6 -8 246 268
use DFFPOSX1  _1506_
timestamp 0
transform 1 0 2250 0 -1 5470
box -6 -8 246 268
use DFFPOSX1  _1507_
timestamp 0
transform -1 0 2750 0 -1 3910
box -6 -8 246 268
use DFFPOSX1  _1508_
timestamp 0
transform 1 0 3350 0 -1 4430
box -6 -8 246 268
use DFFPOSX1  _1509_
timestamp 0
transform 1 0 4050 0 1 3910
box -6 -8 246 268
use DFFPOSX1  _1510_
timestamp 0
transform -1 0 3230 0 -1 3390
box -6 -8 246 268
use DFFPOSX1  _1511_
timestamp 0
transform -1 0 2710 0 -1 3390
box -6 -8 246 268
use DFFPOSX1  _1512_
timestamp 0
transform -1 0 2570 0 1 2870
box -6 -8 246 268
use DFFPOSX1  _1513_
timestamp 0
transform -1 0 3230 0 -1 2870
box -6 -8 246 268
use DFFPOSX1  _1514_
timestamp 0
transform -1 0 3490 0 1 3390
box -6 -8 246 268
use DFFPOSX1  _1515_
timestamp 0
transform -1 0 1110 0 -1 4950
box -6 -8 246 268
use DFFPOSX1  _1516_
timestamp 0
transform -1 0 3990 0 -1 3390
box -6 -8 246 268
use DFFPOSX1  _1517_
timestamp 0
transform -1 0 3590 0 -1 2870
box -6 -8 246 268
use DFFPOSX1  _1518_
timestamp 0
transform -1 0 2490 0 1 2350
box -6 -8 246 268
use DFFPOSX1  _1519_
timestamp 0
transform -1 0 2810 0 -1 2350
box -6 -8 246 268
use DFFPOSX1  _1520_
timestamp 0
transform 1 0 3190 0 1 1830
box -6 -8 246 268
use DFFPOSX1  _1521_
timestamp 0
transform -1 0 3150 0 -1 2350
box -6 -8 246 268
use DFFPOSX1  _1522_
timestamp 0
transform 1 0 10 0 -1 2870
box -6 -8 246 268
use DFFPOSX1  _1523_
timestamp 0
transform 1 0 2770 0 1 3390
box -6 -8 246 268
use DFFPOSX1  _1524_
timestamp 0
transform 1 0 2650 0 1 3910
box -6 -8 246 268
use DFFPOSX1  _1525_
timestamp 0
transform 1 0 2750 0 -1 3910
box -6 -8 246 268
use DFFPOSX1  _1526_
timestamp 0
transform -1 0 3230 0 -1 3910
box -6 -8 246 268
use BUFX2  _1527_
timestamp 0
transform -1 0 130 0 1 2870
box -6 -8 66 268
use BUFX2  _1528_
timestamp 0
transform 1 0 2430 0 -1 1310
box -6 -8 66 268
use BUFX2  _1529_
timestamp 0
transform -1 0 2610 0 -1 1310
box -6 -8 66 268
use BUFX2  _1530_
timestamp 0
transform 1 0 5750 0 -1 2350
box -6 -8 66 268
use BUFX2  _1531_
timestamp 0
transform 1 0 5630 0 -1 2350
box -6 -8 66 268
use BUFX2  _1532_
timestamp 0
transform -1 0 2130 0 1 4950
box -6 -8 66 268
use BUFX2  _1533_
timestamp 0
transform 1 0 2830 0 -1 5470
box -6 -8 66 268
use BUFX2  _1534_
timestamp 0
transform 1 0 2190 0 -1 5470
box -6 -8 66 268
use BUFX2  _1535_
timestamp 0
transform -1 0 2910 0 1 4950
box -6 -8 66 268
use BUFX2  BUFX2_insert0
timestamp 0
transform 1 0 810 0 1 2870
box -6 -8 66 268
use BUFX2  BUFX2_insert1
timestamp 0
transform 1 0 4530 0 -1 3910
box -6 -8 66 268
use BUFX2  BUFX2_insert2
timestamp 0
transform 1 0 2350 0 1 3390
box -6 -8 66 268
use BUFX2  BUFX2_insert3
timestamp 0
transform -1 0 1710 0 -1 3910
box -6 -8 66 268
use BUFX2  BUFX2_insert4
timestamp 0
transform -1 0 830 0 -1 2870
box -6 -8 66 268
use BUFX2  BUFX2_insert5
timestamp 0
transform 1 0 4690 0 1 3390
box -6 -8 66 268
use BUFX2  BUFX2_insert6
timestamp 0
transform 1 0 3490 0 1 3910
box -6 -8 66 268
use BUFX2  BUFX2_insert15
timestamp 0
transform 1 0 2790 0 -1 1310
box -6 -8 66 268
use BUFX2  BUFX2_insert16
timestamp 0
transform 1 0 1850 0 -1 1830
box -6 -8 66 268
use BUFX2  BUFX2_insert17
timestamp 0
transform -1 0 2670 0 1 790
box -6 -8 66 268
use BUFX2  BUFX2_insert18
timestamp 0
transform -1 0 2130 0 1 1830
box -6 -8 66 268
use BUFX2  BUFX2_insert19
timestamp 0
transform 1 0 2450 0 -1 3910
box -6 -8 66 268
use BUFX2  BUFX2_insert20
timestamp 0
transform -1 0 1570 0 -1 4430
box -6 -8 66 268
use BUFX2  BUFX2_insert21
timestamp 0
transform 1 0 3290 0 -1 3910
box -6 -8 66 268
use BUFX2  BUFX2_insert22
timestamp 0
transform -1 0 1390 0 1 4430
box -6 -8 66 268
use BUFX2  BUFX2_insert23
timestamp 0
transform -1 0 3030 0 1 4430
box -6 -8 66 268
use BUFX2  BUFX2_insert24
timestamp 0
transform 1 0 3610 0 1 3910
box -6 -8 66 268
use BUFX2  BUFX2_insert25
timestamp 0
transform -1 0 3710 0 -1 2870
box -6 -8 66 268
use BUFX2  BUFX2_insert26
timestamp 0
transform -1 0 3690 0 1 2870
box -6 -8 66 268
use BUFX2  BUFX2_insert27
timestamp 0
transform -1 0 3350 0 -1 2870
box -6 -8 66 268
use BUFX2  BUFX2_insert28
timestamp 0
transform -1 0 2990 0 -1 2870
box -6 -8 66 268
use BUFX2  BUFX2_insert29
timestamp 0
transform -1 0 2090 0 1 2870
box -6 -8 66 268
use BUFX2  BUFX2_insert30
timestamp 0
transform -1 0 1970 0 1 1310
box -6 -8 66 268
use BUFX2  BUFX2_insert31
timestamp 0
transform 1 0 3650 0 1 1310
box -6 -8 66 268
use BUFX2  BUFX2_insert32
timestamp 0
transform 1 0 2670 0 -1 1310
box -6 -8 66 268
use BUFX2  BUFX2_insert33
timestamp 0
transform -1 0 1770 0 -1 1310
box -6 -8 66 268
use CLKBUF1  CLKBUF1_insert7
timestamp 0
transform -1 0 1470 0 1 3390
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert8
timestamp 0
transform -1 0 1810 0 -1 4430
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert9
timestamp 0
transform 1 0 4110 0 -1 4950
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert10
timestamp 0
transform -1 0 3750 0 -1 3390
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert11
timestamp 0
transform -1 0 1110 0 -1 5470
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert12
timestamp 0
transform 1 0 3570 0 -1 5470
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert13
timestamp 0
transform 1 0 4290 0 -1 3910
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert14
timestamp 0
transform 1 0 2290 0 -1 3390
box -6 -8 186 268
use FILL  FILL85650x23550
timestamp 0
transform -1 0 5730 0 -1 1830
box -6 -8 26 268
use FILL  FILL85650x27450
timestamp 0
transform 1 0 5710 0 1 1830
box -6 -8 26 268
use FILL  FILL85650x46950
timestamp 0
transform -1 0 5730 0 -1 3390
box -6 -8 26 268
use FILL  FILL85650x66450
timestamp 0
transform 1 0 5710 0 1 4430
box -6 -8 26 268
use FILL  FILL85950x11850
timestamp 0
transform 1 0 5730 0 1 790
box -6 -8 26 268
use FILL  FILL85950x23550
timestamp 0
transform -1 0 5750 0 -1 1830
box -6 -8 26 268
use FILL  FILL85950x27450
timestamp 0
transform 1 0 5730 0 1 1830
box -6 -8 26 268
use FILL  FILL85950x46950
timestamp 0
transform -1 0 5750 0 -1 3390
box -6 -8 26 268
use FILL  FILL85950x66450
timestamp 0
transform 1 0 5730 0 1 4430
box -6 -8 26 268
use FILL  FILL85950x78150
timestamp 0
transform -1 0 5750 0 -1 5470
box -6 -8 26 268
use FILL  FILL86250x11850
timestamp 0
transform 1 0 5750 0 1 790
box -6 -8 26 268
use FILL  FILL86250x23550
timestamp 0
transform -1 0 5770 0 -1 1830
box -6 -8 26 268
use FILL  FILL86250x27450
timestamp 0
transform 1 0 5750 0 1 1830
box -6 -8 26 268
use FILL  FILL86250x46950
timestamp 0
transform -1 0 5770 0 -1 3390
box -6 -8 26 268
use FILL  FILL86250x66450
timestamp 0
transform 1 0 5750 0 1 4430
box -6 -8 26 268
use FILL  FILL86250x74250
timestamp 0
transform 1 0 5750 0 1 4950
box -6 -8 26 268
use FILL  FILL86250x78150
timestamp 0
transform -1 0 5770 0 -1 5470
box -6 -8 26 268
use FILL  FILL86550x7950
timestamp 0
transform -1 0 5790 0 -1 790
box -6 -8 26 268
use FILL  FILL86550x11850
timestamp 0
transform 1 0 5770 0 1 790
box -6 -8 26 268
use FILL  FILL86550x23550
timestamp 0
transform -1 0 5790 0 -1 1830
box -6 -8 26 268
use FILL  FILL86550x27450
timestamp 0
transform 1 0 5770 0 1 1830
box -6 -8 26 268
use FILL  FILL86550x35250
timestamp 0
transform 1 0 5770 0 1 2350
box -6 -8 26 268
use FILL  FILL86550x39150
timestamp 0
transform -1 0 5790 0 -1 2870
box -6 -8 26 268
use FILL  FILL86550x46950
timestamp 0
transform -1 0 5790 0 -1 3390
box -6 -8 26 268
use FILL  FILL86550x50850
timestamp 0
transform 1 0 5770 0 1 3390
box -6 -8 26 268
use FILL  FILL86550x54750
timestamp 0
transform -1 0 5790 0 -1 3910
box -6 -8 26 268
use FILL  FILL86550x66450
timestamp 0
transform 1 0 5770 0 1 4430
box -6 -8 26 268
use FILL  FILL86550x74250
timestamp 0
transform 1 0 5770 0 1 4950
box -6 -8 26 268
use FILL  FILL86550x78150
timestamp 0
transform -1 0 5790 0 -1 5470
box -6 -8 26 268
use FILL  FILL86850x150
timestamp 0
transform -1 0 5810 0 -1 270
box -6 -8 26 268
use FILL  FILL86850x4050
timestamp 0
transform 1 0 5790 0 1 270
box -6 -8 26 268
use FILL  FILL86850x7950
timestamp 0
transform -1 0 5810 0 -1 790
box -6 -8 26 268
use FILL  FILL86850x11850
timestamp 0
transform 1 0 5790 0 1 790
box -6 -8 26 268
use FILL  FILL86850x23550
timestamp 0
transform -1 0 5810 0 -1 1830
box -6 -8 26 268
use FILL  FILL86850x27450
timestamp 0
transform 1 0 5790 0 1 1830
box -6 -8 26 268
use FILL  FILL86850x35250
timestamp 0
transform 1 0 5790 0 1 2350
box -6 -8 26 268
use FILL  FILL86850x39150
timestamp 0
transform -1 0 5810 0 -1 2870
box -6 -8 26 268
use FILL  FILL86850x43050
timestamp 0
transform 1 0 5790 0 1 2870
box -6 -8 26 268
use FILL  FILL86850x46950
timestamp 0
transform -1 0 5810 0 -1 3390
box -6 -8 26 268
use FILL  FILL86850x50850
timestamp 0
transform 1 0 5790 0 1 3390
box -6 -8 26 268
use FILL  FILL86850x54750
timestamp 0
transform -1 0 5810 0 -1 3910
box -6 -8 26 268
use FILL  FILL86850x58650
timestamp 0
transform 1 0 5790 0 1 3910
box -6 -8 26 268
use FILL  FILL86850x66450
timestamp 0
transform 1 0 5790 0 1 4430
box -6 -8 26 268
use FILL  FILL86850x74250
timestamp 0
transform 1 0 5790 0 1 4950
box -6 -8 26 268
use FILL  FILL86850x78150
timestamp 0
transform -1 0 5810 0 -1 5470
box -6 -8 26 268
use FILL  FILL87150x150
timestamp 0
transform -1 0 5830 0 -1 270
box -6 -8 26 268
use FILL  FILL87150x4050
timestamp 0
transform 1 0 5810 0 1 270
box -6 -8 26 268
use FILL  FILL87150x7950
timestamp 0
transform -1 0 5830 0 -1 790
box -6 -8 26 268
use FILL  FILL87150x11850
timestamp 0
transform 1 0 5810 0 1 790
box -6 -8 26 268
use FILL  FILL87150x15750
timestamp 0
transform -1 0 5830 0 -1 1310
box -6 -8 26 268
use FILL  FILL87150x19650
timestamp 0
transform 1 0 5810 0 1 1310
box -6 -8 26 268
use FILL  FILL87150x23550
timestamp 0
transform -1 0 5830 0 -1 1830
box -6 -8 26 268
use FILL  FILL87150x27450
timestamp 0
transform 1 0 5810 0 1 1830
box -6 -8 26 268
use FILL  FILL87150x31350
timestamp 0
transform -1 0 5830 0 -1 2350
box -6 -8 26 268
use FILL  FILL87150x35250
timestamp 0
transform 1 0 5810 0 1 2350
box -6 -8 26 268
use FILL  FILL87150x39150
timestamp 0
transform -1 0 5830 0 -1 2870
box -6 -8 26 268
use FILL  FILL87150x43050
timestamp 0
transform 1 0 5810 0 1 2870
box -6 -8 26 268
use FILL  FILL87150x46950
timestamp 0
transform -1 0 5830 0 -1 3390
box -6 -8 26 268
use FILL  FILL87150x50850
timestamp 0
transform 1 0 5810 0 1 3390
box -6 -8 26 268
use FILL  FILL87150x54750
timestamp 0
transform -1 0 5830 0 -1 3910
box -6 -8 26 268
use FILL  FILL87150x58650
timestamp 0
transform 1 0 5810 0 1 3910
box -6 -8 26 268
use FILL  FILL87150x66450
timestamp 0
transform 1 0 5810 0 1 4430
box -6 -8 26 268
use FILL  FILL87150x70350
timestamp 0
transform -1 0 5830 0 -1 4950
box -6 -8 26 268
use FILL  FILL87150x74250
timestamp 0
transform 1 0 5810 0 1 4950
box -6 -8 26 268
use FILL  FILL87150x78150
timestamp 0
transform -1 0 5830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__723_
timestamp 0
transform 1 0 2670 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__724_
timestamp 0
transform -1 0 2590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__725_
timestamp 0
transform -1 0 2290 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__726_
timestamp 0
transform -1 0 2290 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__727_
timestamp 0
transform 1 0 3010 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__728_
timestamp 0
transform -1 0 3650 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__729_
timestamp 0
transform -1 0 950 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__730_
timestamp 0
transform -1 0 2150 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__731_
timestamp 0
transform -1 0 2230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__732_
timestamp 0
transform -1 0 4130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__733_
timestamp 0
transform 1 0 3270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__734_
timestamp 0
transform 1 0 3130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__735_
timestamp 0
transform -1 0 1110 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__736_
timestamp 0
transform -1 0 2550 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__737_
timestamp 0
transform -1 0 2690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__738_
timestamp 0
transform 1 0 2450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__739_
timestamp 0
transform 1 0 2310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__740_
timestamp 0
transform -1 0 1870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__741_
timestamp 0
transform -1 0 2090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__742_
timestamp 0
transform 1 0 2710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__743_
timestamp 0
transform -1 0 2910 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__744_
timestamp 0
transform 1 0 1870 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__745_
timestamp 0
transform -1 0 2590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__746_
timestamp 0
transform -1 0 2830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__747_
timestamp 0
transform -1 0 2050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__748_
timestamp 0
transform -1 0 2270 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__749_
timestamp 0
transform -1 0 4690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__750_
timestamp 0
transform 1 0 2650 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__751_
timestamp 0
transform 1 0 2510 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__752_
timestamp 0
transform -1 0 4330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__753_
timestamp 0
transform -1 0 4090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__754_
timestamp 0
transform 1 0 4170 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__755_
timestamp 0
transform -1 0 4110 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__756_
timestamp 0
transform -1 0 3810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__757_
timestamp 0
transform -1 0 3930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__758_
timestamp 0
transform 1 0 2750 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__759_
timestamp 0
transform -1 0 2890 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__760_
timestamp 0
transform 1 0 3250 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__761_
timestamp 0
transform -1 0 3390 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__762_
timestamp 0
transform -1 0 4110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__763_
timestamp 0
transform 1 0 3950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__764_
timestamp 0
transform 1 0 3650 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__765_
timestamp 0
transform -1 0 3790 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__766_
timestamp 0
transform 1 0 350 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__767_
timestamp 0
transform -1 0 2670 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__768_
timestamp 0
transform 1 0 690 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__769_
timestamp 0
transform -1 0 270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__770_
timestamp 0
transform 1 0 730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__771_
timestamp 0
transform 1 0 590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__772_
timestamp 0
transform 1 0 2030 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__773_
timestamp 0
transform 1 0 2530 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__774_
timestamp 0
transform 1 0 2150 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__775_
timestamp 0
transform 1 0 370 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__776_
timestamp 0
transform 1 0 2210 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__777_
timestamp 0
transform 1 0 610 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__778_
timestamp 0
transform 1 0 10 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__779_
timestamp 0
transform 1 0 290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__780_
timestamp 0
transform 1 0 130 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__781_
timestamp 0
transform 1 0 1150 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__782_
timestamp 0
transform 1 0 2410 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__783_
timestamp 0
transform 1 0 1490 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__784_
timestamp 0
transform -1 0 1290 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__785_
timestamp 0
transform 1 0 2090 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__786_
timestamp 0
transform 1 0 1610 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__787_
timestamp 0
transform 1 0 2250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__788_
timestamp 0
transform 1 0 2730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__789_
timestamp 0
transform 1 0 2590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__790_
timestamp 0
transform 1 0 1350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__791_
timestamp 0
transform 1 0 1590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__792_
timestamp 0
transform 1 0 1450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__793_
timestamp 0
transform 1 0 1950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__794_
timestamp 0
transform 1 0 2450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__795_
timestamp 0
transform -1 0 2310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__796_
timestamp 0
transform -1 0 4730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__797_
timestamp 0
transform -1 0 4430 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__798_
timestamp 0
transform -1 0 4550 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__799_
timestamp 0
transform -1 0 5370 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__800_
timestamp 0
transform -1 0 4310 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__801_
timestamp 0
transform -1 0 5230 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__802_
timestamp 0
transform -1 0 5710 0 1 270
box -6 -8 26 268
use FILL  FILL_0__803_
timestamp 0
transform -1 0 5510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__804_
timestamp 0
transform 1 0 5370 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__805_
timestamp 0
transform 1 0 5250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__806_
timestamp 0
transform -1 0 4370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__807_
timestamp 0
transform -1 0 4550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__808_
timestamp 0
transform -1 0 3670 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__809_
timestamp 0
transform 1 0 3090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__810_
timestamp 0
transform 1 0 3030 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__811_
timestamp 0
transform -1 0 3730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__812_
timestamp 0
transform -1 0 4410 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__813_
timestamp 0
transform 1 0 3710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__814_
timestamp 0
transform 1 0 590 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__815_
timestamp 0
transform -1 0 2030 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__816_
timestamp 0
transform 1 0 690 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__817_
timestamp 0
transform 1 0 1110 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__818_
timestamp 0
transform 1 0 1530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__819_
timestamp 0
transform -1 0 1690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__820_
timestamp 0
transform 1 0 1450 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__821_
timestamp 0
transform 1 0 950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__822_
timestamp 0
transform -1 0 1330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__823_
timestamp 0
transform -1 0 1430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__824_
timestamp 0
transform 1 0 1470 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__825_
timestamp 0
transform 1 0 1290 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__826_
timestamp 0
transform -1 0 1090 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__827_
timestamp 0
transform 1 0 1590 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__828_
timestamp 0
transform 1 0 1190 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__829_
timestamp 0
transform 1 0 1290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__830_
timestamp 0
transform -1 0 1530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__831_
timestamp 0
transform 1 0 1650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__832_
timestamp 0
transform -1 0 1410 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__833_
timestamp 0
transform 1 0 1790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__834_
timestamp 0
transform 1 0 1750 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__835_
timestamp 0
transform -1 0 1930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__836_
timestamp 0
transform 1 0 1850 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__837_
timestamp 0
transform -1 0 1350 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__838_
timestamp 0
transform -1 0 1290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__839_
timestamp 0
transform -1 0 890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__840_
timestamp 0
transform -1 0 1150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__841_
timestamp 0
transform -1 0 990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__842_
timestamp 0
transform 1 0 1870 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__843_
timestamp 0
transform -1 0 1770 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__844_
timestamp 0
transform 1 0 1630 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__845_
timestamp 0
transform 1 0 370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__846_
timestamp 0
transform -1 0 2150 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__847_
timestamp 0
transform -1 0 950 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__848_
timestamp 0
transform -1 0 1450 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__849_
timestamp 0
transform 1 0 1050 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__850_
timestamp 0
transform -1 0 950 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__851_
timestamp 0
transform -1 0 1210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__852_
timestamp 0
transform -1 0 670 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__853_
timestamp 0
transform -1 0 870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__854_
timestamp 0
transform 1 0 1050 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__855_
timestamp 0
transform -1 0 1190 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__856_
timestamp 0
transform 1 0 450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__857_
timestamp 0
transform -1 0 530 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__858_
timestamp 0
transform 1 0 650 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__859_
timestamp 0
transform -1 0 1170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__860_
timestamp 0
transform -1 0 810 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__861_
timestamp 0
transform 1 0 1910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__862_
timestamp 0
transform -1 0 1730 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__863_
timestamp 0
transform -1 0 2810 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__864_
timestamp 0
transform -1 0 2690 0 1 790
box -6 -8 26 268
use FILL  FILL_0__865_
timestamp 0
transform -1 0 1990 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__866_
timestamp 0
transform -1 0 1590 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__867_
timestamp 0
transform 1 0 1010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__868_
timestamp 0
transform 1 0 790 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__869_
timestamp 0
transform -1 0 430 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__870_
timestamp 0
transform -1 0 610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__871_
timestamp 0
transform -1 0 870 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__872_
timestamp 0
transform 1 0 510 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__873_
timestamp 0
transform -1 0 610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__874_
timestamp 0
transform -1 0 750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__875_
timestamp 0
transform 1 0 310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__876_
timestamp 0
transform 1 0 430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__877_
timestamp 0
transform -1 0 30 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__878_
timestamp 0
transform -1 0 310 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__879_
timestamp 0
transform -1 0 470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__880_
timestamp 0
transform -1 0 390 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__881_
timestamp 0
transform -1 0 590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__882_
timestamp 0
transform 1 0 1550 0 1 790
box -6 -8 26 268
use FILL  FILL_0__883_
timestamp 0
transform 1 0 1150 0 1 790
box -6 -8 26 268
use FILL  FILL_0__884_
timestamp 0
transform 1 0 1350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__885_
timestamp 0
transform -1 0 970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__886_
timestamp 0
transform 1 0 1270 0 1 790
box -6 -8 26 268
use FILL  FILL_0__887_
timestamp 0
transform -1 0 830 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__888_
timestamp 0
transform -1 0 870 0 1 790
box -6 -8 26 268
use FILL  FILL_0__889_
timestamp 0
transform -1 0 2310 0 1 790
box -6 -8 26 268
use FILL  FILL_0__890_
timestamp 0
transform 1 0 910 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__891_
timestamp 0
transform 1 0 710 0 1 790
box -6 -8 26 268
use FILL  FILL_0__892_
timestamp 0
transform -1 0 590 0 1 790
box -6 -8 26 268
use FILL  FILL_0__893_
timestamp 0
transform -1 0 730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__894_
timestamp 0
transform -1 0 1010 0 1 790
box -6 -8 26 268
use FILL  FILL_0__895_
timestamp 0
transform -1 0 690 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__896_
timestamp 0
transform -1 0 410 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__897_
timestamp 0
transform 1 0 2670 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__898_
timestamp 0
transform 1 0 2150 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__899_
timestamp 0
transform 1 0 4210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__900_
timestamp 0
transform -1 0 2270 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__901_
timestamp 0
transform 1 0 2150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__902_
timestamp 0
transform -1 0 2130 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__903_
timestamp 0
transform 1 0 290 0 1 790
box -6 -8 26 268
use FILL  FILL_0__904_
timestamp 0
transform -1 0 550 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__905_
timestamp 0
transform -1 0 450 0 1 790
box -6 -8 26 268
use FILL  FILL_0__906_
timestamp 0
transform 1 0 10 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__907_
timestamp 0
transform 1 0 150 0 1 790
box -6 -8 26 268
use FILL  FILL_0__908_
timestamp 0
transform -1 0 330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__909_
timestamp 0
transform 1 0 330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__910_
timestamp 0
transform -1 0 210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__911_
timestamp 0
transform -1 0 30 0 1 790
box -6 -8 26 268
use FILL  FILL_0__912_
timestamp 0
transform -1 0 290 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__913_
timestamp 0
transform 1 0 130 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__914_
timestamp 0
transform 1 0 10 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__915_
timestamp 0
transform 1 0 150 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__916_
timestamp 0
transform 1 0 170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__917_
timestamp 0
transform 1 0 10 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__918_
timestamp 0
transform 1 0 2810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__919_
timestamp 0
transform 1 0 730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__920_
timestamp 0
transform 1 0 130 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__921_
timestamp 0
transform 1 0 110 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__922_
timestamp 0
transform 1 0 2390 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__923_
timestamp 0
transform 1 0 2010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__924_
timestamp 0
transform 1 0 2150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__925_
timestamp 0
transform 1 0 3850 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__926_
timestamp 0
transform -1 0 2690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__927_
timestamp 0
transform 1 0 2530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__928_
timestamp 0
transform -1 0 2450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__929_
timestamp 0
transform 1 0 2310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__930_
timestamp 0
transform -1 0 2550 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__931_
timestamp 0
transform -1 0 2390 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__932_
timestamp 0
transform -1 0 2130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__933_
timestamp 0
transform 1 0 1030 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__934_
timestamp 0
transform 1 0 1070 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__935_
timestamp 0
transform 1 0 1510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__936_
timestamp 0
transform -1 0 1970 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__937_
timestamp 0
transform -1 0 2190 0 1 790
box -6 -8 26 268
use FILL  FILL_0__938_
timestamp 0
transform -1 0 1430 0 1 790
box -6 -8 26 268
use FILL  FILL_0__939_
timestamp 0
transform -1 0 1370 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__940_
timestamp 0
transform -1 0 1710 0 1 790
box -6 -8 26 268
use FILL  FILL_0__941_
timestamp 0
transform -1 0 2790 0 1 790
box -6 -8 26 268
use FILL  FILL_0__942_
timestamp 0
transform 1 0 1790 0 1 790
box -6 -8 26 268
use FILL  FILL_0__943_
timestamp 0
transform -1 0 2430 0 1 790
box -6 -8 26 268
use FILL  FILL_0__944_
timestamp 0
transform -1 0 1530 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__945_
timestamp 0
transform -1 0 1190 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__946_
timestamp 0
transform -1 0 1670 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__947_
timestamp 0
transform -1 0 1210 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__948_
timestamp 0
transform -1 0 1050 0 1 270
box -6 -8 26 268
use FILL  FILL_0__949_
timestamp 0
transform -1 0 950 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__950_
timestamp 0
transform -1 0 1990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__951_
timestamp 0
transform 1 0 1310 0 1 270
box -6 -8 26 268
use FILL  FILL_0__952_
timestamp 0
transform -1 0 1190 0 1 270
box -6 -8 26 268
use FILL  FILL_0__953_
timestamp 0
transform -1 0 770 0 1 270
box -6 -8 26 268
use FILL  FILL_0__954_
timestamp 0
transform -1 0 330 0 1 270
box -6 -8 26 268
use FILL  FILL_0__955_
timestamp 0
transform -1 0 270 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__956_
timestamp 0
transform -1 0 910 0 1 270
box -6 -8 26 268
use FILL  FILL_0__957_
timestamp 0
transform -1 0 810 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__958_
timestamp 0
transform -1 0 630 0 1 270
box -6 -8 26 268
use FILL  FILL_0__959_
timestamp 0
transform -1 0 190 0 1 270
box -6 -8 26 268
use FILL  FILL_0__960_
timestamp 0
transform -1 0 390 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__961_
timestamp 0
transform -1 0 490 0 1 270
box -6 -8 26 268
use FILL  FILL_0__962_
timestamp 0
transform -1 0 30 0 1 270
box -6 -8 26 268
use FILL  FILL_0__963_
timestamp 0
transform -1 0 30 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__964_
timestamp 0
transform 1 0 10 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__965_
timestamp 0
transform 1 0 10 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__966_
timestamp 0
transform -1 0 830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__967_
timestamp 0
transform -1 0 950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__968_
timestamp 0
transform 1 0 1070 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__969_
timestamp 0
transform 1 0 130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__970_
timestamp 0
transform 1 0 510 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__971_
timestamp 0
transform -1 0 670 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__972_
timestamp 0
transform 1 0 2790 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__973_
timestamp 0
transform 1 0 2230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__974_
timestamp 0
transform 1 0 2250 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__975_
timestamp 0
transform 1 0 1730 0 1 270
box -6 -8 26 268
use FILL  FILL_0__976_
timestamp 0
transform 1 0 1830 0 1 270
box -6 -8 26 268
use FILL  FILL_0__977_
timestamp 0
transform 1 0 2910 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__978_
timestamp 0
transform -1 0 3350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__979_
timestamp 0
transform 1 0 3190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__980_
timestamp 0
transform -1 0 3470 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__981_
timestamp 0
transform -1 0 3490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__982_
timestamp 0
transform -1 0 3070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__983_
timestamp 0
transform -1 0 2970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__984_
timestamp 0
transform -1 0 3330 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__985_
timestamp 0
transform -1 0 2930 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__986_
timestamp 0
transform 1 0 3050 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__987_
timestamp 0
transform -1 0 2870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__988_
timestamp 0
transform -1 0 2070 0 1 790
box -6 -8 26 268
use FILL  FILL_0__989_
timestamp 0
transform 1 0 1910 0 1 790
box -6 -8 26 268
use FILL  FILL_0__990_
timestamp 0
transform 1 0 3730 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__991_
timestamp 0
transform -1 0 3130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__992_
timestamp 0
transform -1 0 3410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__993_
timestamp 0
transform -1 0 3730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__994_
timestamp 0
transform -1 0 3790 0 1 790
box -6 -8 26 268
use FILL  FILL_0__995_
timestamp 0
transform -1 0 3510 0 1 790
box -6 -8 26 268
use FILL  FILL_0__996_
timestamp 0
transform -1 0 3370 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__997_
timestamp 0
transform -1 0 3730 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__998_
timestamp 0
transform 1 0 3610 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__999_
timestamp 0
transform -1 0 3250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1000_
timestamp 0
transform -1 0 3230 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1001_
timestamp 0
transform -1 0 2650 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1002_
timestamp 0
transform -1 0 2110 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1003_
timestamp 0
transform 1 0 1790 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1004_
timestamp 0
transform 1 0 3190 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1005_
timestamp 0
transform -1 0 3370 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1006_
timestamp 0
transform -1 0 2930 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1007_
timestamp 0
transform 1 0 2490 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1008_
timestamp 0
transform 1 0 2970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1009_
timestamp 0
transform 1 0 2910 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1010_
timestamp 0
transform -1 0 3070 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1011_
timestamp 0
transform -1 0 3130 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1012_
timestamp 0
transform -1 0 2570 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1013_
timestamp 0
transform 1 0 1450 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1014_
timestamp 0
transform 1 0 1590 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1015_
timestamp 0
transform -1 0 2990 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1016_
timestamp 0
transform -1 0 2370 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1017_
timestamp 0
transform -1 0 2290 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1018_
timestamp 0
transform -1 0 1990 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1019_
timestamp 0
transform -1 0 2710 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1020_
timestamp 0
transform 1 0 2410 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1021_
timestamp 0
transform -1 0 2470 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1022_
timestamp 0
transform 1 0 1770 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1023_
timestamp 0
transform -1 0 1450 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1024_
timestamp 0
transform 1 0 1310 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1025_
timestamp 0
transform 1 0 1890 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1026_
timestamp 0
transform 1 0 10 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1027_
timestamp 0
transform 1 0 230 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1028_
timestamp 0
transform -1 0 2330 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1029_
timestamp 0
transform 1 0 2130 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1030_
timestamp 0
transform -1 0 2190 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1031_
timestamp 0
transform -1 0 2050 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1032_
timestamp 0
transform 1 0 1330 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1033_
timestamp 0
transform 1 0 1170 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1034_
timestamp 0
transform 1 0 1610 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1035_
timestamp 0
transform -1 0 2750 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1036_
timestamp 0
transform 1 0 2590 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1037_
timestamp 0
transform -1 0 3210 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1038_
timestamp 0
transform 1 0 3770 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1039_
timestamp 0
transform 1 0 3270 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1040_
timestamp 0
transform 1 0 3370 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1041_
timestamp 0
transform 1 0 3970 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1042_
timestamp 0
transform 1 0 3710 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1043_
timestamp 0
transform -1 0 4290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1044_
timestamp 0
transform 1 0 3430 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1045_
timestamp 0
transform 1 0 3570 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1046_
timestamp 0
transform 1 0 4130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1047_
timestamp 0
transform -1 0 4050 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1048_
timestamp 0
transform 1 0 3850 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1049_
timestamp 0
transform -1 0 3630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1050_
timestamp 0
transform -1 0 3770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1051_
timestamp 0
transform -1 0 3910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1052_
timestamp 0
transform -1 0 4770 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1053_
timestamp 0
transform -1 0 3470 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1054_
timestamp 0
transform 1 0 3910 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1055_
timestamp 0
transform 1 0 4770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1056_
timestamp 0
transform 1 0 4890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1057_
timestamp 0
transform -1 0 4390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1058_
timestamp 0
transform -1 0 4430 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1059_
timestamp 0
transform 1 0 4030 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1060_
timestamp 0
transform -1 0 4130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1061_
timestamp 0
transform -1 0 4270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1062_
timestamp 0
transform 1 0 4550 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1063_
timestamp 0
transform 1 0 4270 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1064_
timestamp 0
transform 1 0 4310 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1065_
timestamp 0
transform -1 0 3570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1066_
timestamp 0
transform -1 0 3650 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1067_
timestamp 0
transform -1 0 4150 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1068_
timestamp 0
transform 1 0 3950 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1069_
timestamp 0
transform 1 0 3830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1070_
timestamp 0
transform 1 0 3970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1071_
timestamp 0
transform -1 0 3990 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1072_
timestamp 0
transform -1 0 4490 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1073_
timestamp 0
transform 1 0 4770 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1074_
timestamp 0
transform 1 0 4410 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1075_
timestamp 0
transform 1 0 4130 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1076_
timestamp 0
transform -1 0 4930 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1077_
timestamp 0
transform -1 0 4230 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1078_
timestamp 0
transform 1 0 2770 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1079_
timestamp 0
transform 1 0 3050 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1080_
timestamp 0
transform -1 0 4650 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1081_
timestamp 0
transform 1 0 4610 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1082_
timestamp 0
transform -1 0 4370 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1083_
timestamp 0
transform -1 0 3950 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1084_
timestamp 0
transform -1 0 4190 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1085_
timestamp 0
transform -1 0 4510 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1086_
timestamp 0
transform -1 0 3810 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1087_
timestamp 0
transform -1 0 3650 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1088_
timestamp 0
transform -1 0 2850 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1089_
timestamp 0
transform 1 0 2830 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1090_
timestamp 0
transform -1 0 3650 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1091_
timestamp 0
transform -1 0 4090 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1092_
timestamp 0
transform -1 0 3510 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1093_
timestamp 0
transform 1 0 3370 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1094_
timestamp 0
transform 1 0 1770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1095_
timestamp 0
transform 1 0 2130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1096_
timestamp 0
transform 1 0 1990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1097_
timestamp 0
transform 1 0 3750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1098_
timestamp 0
transform -1 0 3130 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1099_
timestamp 0
transform -1 0 3530 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1100_
timestamp 0
transform 1 0 3390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1101_
timestamp 0
transform -1 0 4050 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1102_
timestamp 0
transform 1 0 3870 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1103_
timestamp 0
transform 1 0 3850 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1104_
timestamp 0
transform -1 0 5710 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1105_
timestamp 0
transform -1 0 5210 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1106_
timestamp 0
transform 1 0 5050 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1107_
timestamp 0
transform 1 0 4230 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1108_
timestamp 0
transform -1 0 4430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1109_
timestamp 0
transform 1 0 5210 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1110_
timestamp 0
transform 1 0 5050 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1111_
timestamp 0
transform 1 0 5370 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1112_
timestamp 0
transform -1 0 5650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1113_
timestamp 0
transform 1 0 4650 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1114_
timestamp 0
transform 1 0 4470 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1115_
timestamp 0
transform 1 0 4530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1116_
timestamp 0
transform 1 0 4350 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1117_
timestamp 0
transform 1 0 4190 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1118_
timestamp 0
transform 1 0 4590 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1119_
timestamp 0
transform -1 0 5350 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1120_
timestamp 0
transform 1 0 4530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1121_
timestamp 0
transform -1 0 4750 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1122_
timestamp 0
transform -1 0 5190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1123_
timestamp 0
transform 1 0 5590 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1124_
timestamp 0
transform -1 0 5450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1125_
timestamp 0
transform 1 0 5030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1126_
timestamp 0
transform -1 0 5230 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1127_
timestamp 0
transform 1 0 5390 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1128_
timestamp 0
transform -1 0 5570 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1129_
timestamp 0
transform -1 0 4290 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1130_
timestamp 0
transform 1 0 5130 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1131_
timestamp 0
transform -1 0 5270 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1132_
timestamp 0
transform -1 0 4810 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1133_
timestamp 0
transform 1 0 4930 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1134_
timestamp 0
transform 1 0 5070 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1135_
timestamp 0
transform 1 0 5110 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1136_
timestamp 0
transform -1 0 5430 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1137_
timestamp 0
transform -1 0 5550 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1138_
timestamp 0
transform -1 0 4990 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1139_
timestamp 0
transform 1 0 4830 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1140_
timestamp 0
transform 1 0 4970 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1141_
timestamp 0
transform 1 0 4870 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1142_
timestamp 0
transform -1 0 4710 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1143_
timestamp 0
transform -1 0 5290 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1144_
timestamp 0
transform -1 0 4570 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1145_
timestamp 0
transform -1 0 4250 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1146_
timestamp 0
transform 1 0 4170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1147_
timestamp 0
transform -1 0 3770 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1148_
timestamp 0
transform 1 0 3990 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1149_
timestamp 0
transform -1 0 4110 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1150_
timestamp 0
transform 1 0 5510 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1151_
timestamp 0
transform 1 0 5610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1152_
timestamp 0
transform -1 0 5310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1153_
timestamp 0
transform 1 0 4330 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1154_
timestamp 0
transform 1 0 4110 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1155_
timestamp 0
transform 1 0 4450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1156_
timestamp 0
transform 1 0 4590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1157_
timestamp 0
transform 1 0 4190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1158_
timestamp 0
transform 1 0 4730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1159_
timestamp 0
transform -1 0 5190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1160_
timestamp 0
transform -1 0 4430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1161_
timestamp 0
transform -1 0 4890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1162_
timestamp 0
transform 1 0 4330 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1163_
timestamp 0
transform -1 0 4510 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1164_
timestamp 0
transform 1 0 4770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1165_
timestamp 0
transform 1 0 4650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1166_
timestamp 0
transform 1 0 4750 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1167_
timestamp 0
transform 1 0 5290 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1168_
timestamp 0
transform -1 0 5470 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1169_
timestamp 0
transform 1 0 4610 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1170_
timestamp 0
transform 1 0 4890 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1171_
timestamp 0
transform 1 0 5150 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1172_
timestamp 0
transform -1 0 5450 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1173_
timestamp 0
transform 1 0 5330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1174_
timestamp 0
transform 1 0 5010 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1175_
timestamp 0
transform -1 0 5490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1176_
timestamp 0
transform 1 0 5070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1177_
timestamp 0
transform -1 0 4930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1178_
timestamp 0
transform -1 0 5570 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1179_
timestamp 0
transform -1 0 5430 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1180_
timestamp 0
transform -1 0 5210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1181_
timestamp 0
transform -1 0 4490 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1182_
timestamp 0
transform -1 0 4010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1183_
timestamp 0
transform -1 0 3950 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1184_
timestamp 0
transform 1 0 3850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1185_
timestamp 0
transform -1 0 4950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1186_
timestamp 0
transform 1 0 4610 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1187_
timestamp 0
transform -1 0 4370 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1188_
timestamp 0
transform -1 0 4870 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1189_
timestamp 0
transform 1 0 4730 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1190_
timestamp 0
transform -1 0 4510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1191_
timestamp 0
transform 1 0 4350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1192_
timestamp 0
transform 1 0 5590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1193_
timestamp 0
transform -1 0 5030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1194_
timestamp 0
transform 1 0 5430 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1195_
timestamp 0
transform 1 0 4910 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1196_
timestamp 0
transform -1 0 4590 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1197_
timestamp 0
transform 1 0 4310 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1198_
timestamp 0
transform 1 0 4690 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1199_
timestamp 0
transform -1 0 4830 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1200_
timestamp 0
transform 1 0 5230 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1201_
timestamp 0
transform 1 0 5430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1202_
timestamp 0
transform 1 0 5290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1203_
timestamp 0
transform -1 0 5690 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1204_
timestamp 0
transform -1 0 5550 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1205_
timestamp 0
transform -1 0 5690 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1206_
timestamp 0
transform 1 0 5670 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1207_
timestamp 0
transform -1 0 5590 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1208_
timestamp 0
transform 1 0 5650 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1209_
timestamp 0
transform -1 0 5530 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1210_
timestamp 0
transform -1 0 5410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1211_
timestamp 0
transform -1 0 5150 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1212_
timestamp 0
transform -1 0 3250 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1213_
timestamp 0
transform 1 0 2970 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1214_
timestamp 0
transform -1 0 3870 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1215_
timestamp 0
transform 1 0 3690 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1216_
timestamp 0
transform -1 0 4910 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1217_
timestamp 0
transform 1 0 4750 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1218_
timestamp 0
transform -1 0 5010 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1219_
timestamp 0
transform 1 0 4910 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1220_
timestamp 0
transform -1 0 5070 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1221_
timestamp 0
transform -1 0 5650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1222_
timestamp 0
transform 1 0 5130 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1223_
timestamp 0
transform 1 0 4950 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1224_
timestamp 0
transform 1 0 4670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1225_
timestamp 0
transform 1 0 4450 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1226_
timestamp 0
transform 1 0 4810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1227_
timestamp 0
transform 1 0 5050 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1228_
timestamp 0
transform 1 0 5190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1229_
timestamp 0
transform -1 0 5470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1230_
timestamp 0
transform 1 0 5510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1231_
timestamp 0
transform 1 0 5690 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1232_
timestamp 0
transform -1 0 5710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1233_
timestamp 0
transform 1 0 5510 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1234_
timestamp 0
transform -1 0 5670 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1235_
timestamp 0
transform 1 0 5630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1236_
timestamp 0
transform 1 0 5170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1237_
timestamp 0
transform 1 0 5710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1238_
timestamp 0
transform -1 0 5390 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1239_
timestamp 0
transform -1 0 5250 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1240_
timestamp 0
transform -1 0 5310 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1241_
timestamp 0
transform -1 0 5270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1242_
timestamp 0
transform -1 0 5130 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1243_
timestamp 0
transform 1 0 5330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1244_
timestamp 0
transform 1 0 4530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1245_
timestamp 0
transform 1 0 4910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1246_
timestamp 0
transform 1 0 5110 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1247_
timestamp 0
transform -1 0 4990 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1248_
timestamp 0
transform 1 0 4970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1249_
timestamp 0
transform -1 0 5390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1250_
timestamp 0
transform -1 0 4610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1251_
timestamp 0
transform 1 0 4830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1252_
timestamp 0
transform 1 0 4690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1253_
timestamp 0
transform -1 0 5410 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1254_
timestamp 0
transform -1 0 5270 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1255_
timestamp 0
transform -1 0 5310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1256_
timestamp 0
transform -1 0 5170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1257_
timestamp 0
transform 1 0 5230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1258_
timestamp 0
transform 1 0 5090 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1259_
timestamp 0
transform 1 0 5050 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1260_
timestamp 0
transform -1 0 150 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1261_
timestamp 0
transform 1 0 10 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1262_
timestamp 0
transform 1 0 250 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1263_
timestamp 0
transform -1 0 390 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1264_
timestamp 0
transform -1 0 1010 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1265_
timestamp 0
transform 1 0 490 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1266_
timestamp 0
transform -1 0 790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1267_
timestamp 0
transform 1 0 510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1268_
timestamp 0
transform 1 0 290 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1269_
timestamp 0
transform -1 0 150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1270_
timestamp 0
transform 1 0 10 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1271_
timestamp 0
transform 1 0 250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1272_
timestamp 0
transform 1 0 390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1273_
timestamp 0
transform 1 0 810 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1274_
timestamp 0
transform 1 0 430 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1275_
timestamp 0
transform -1 0 650 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1276_
timestamp 0
transform -1 0 1810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1277_
timestamp 0
transform 1 0 1590 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1278_
timestamp 0
transform 1 0 2010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1279_
timestamp 0
transform 1 0 1710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1280_
timestamp 0
transform -1 0 1930 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1281_
timestamp 0
transform 1 0 1770 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1282_
timestamp 0
transform 1 0 250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1283_
timestamp 0
transform -1 0 490 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1284_
timestamp 0
transform 1 0 650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1285_
timestamp 0
transform -1 0 790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1286_
timestamp 0
transform -1 0 1470 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1287_
timestamp 0
transform 1 0 1310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1288_
timestamp 0
transform -1 0 190 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1289_
timestamp 0
transform -1 0 30 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1290_
timestamp 0
transform 1 0 10 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1291_
timestamp 0
transform 1 0 10 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1292_
timestamp 0
transform 1 0 290 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1293_
timestamp 0
transform -1 0 570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1294_
timestamp 0
transform 1 0 410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1295_
timestamp 0
transform -1 0 150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1296_
timestamp 0
transform -1 0 30 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1297_
timestamp 0
transform 1 0 170 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1298_
timestamp 0
transform -1 0 250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1299_
timestamp 0
transform 1 0 10 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1300_
timestamp 0
transform -1 0 650 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1301_
timestamp 0
transform 1 0 130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1302_
timestamp 0
transform -1 0 670 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1303_
timestamp 0
transform -1 0 810 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1304_
timestamp 0
transform 1 0 510 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1305_
timestamp 0
transform -1 0 370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1306_
timestamp 0
transform 1 0 270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1307_
timestamp 0
transform -1 0 630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1308_
timestamp 0
transform -1 0 550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1309_
timestamp 0
transform -1 0 490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1310_
timestamp 0
transform -1 0 1490 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1311_
timestamp 0
transform 1 0 670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1312_
timestamp 0
transform 1 0 830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1313_
timestamp 0
transform -1 0 970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1314_
timestamp 0
transform -1 0 890 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1315_
timestamp 0
transform 1 0 1010 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1316_
timestamp 0
transform 1 0 1230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1317_
timestamp 0
transform -1 0 1150 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1318_
timestamp 0
transform 1 0 1630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1319_
timestamp 0
transform -1 0 1530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1320_
timestamp 0
transform 1 0 1270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1321_
timestamp 0
transform -1 0 1390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1322_
timestamp 0
transform 1 0 1610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1323_
timestamp 0
transform 1 0 2270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1324_
timestamp 0
transform 1 0 2130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1325_
timestamp 0
transform -1 0 1670 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1326_
timestamp 0
transform 1 0 390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1327_
timestamp 0
transform -1 0 1030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1328_
timestamp 0
transform 1 0 1130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1329_
timestamp 0
transform -1 0 1090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1330_
timestamp 0
transform 1 0 970 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1331_
timestamp 0
transform -1 0 410 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1332_
timestamp 0
transform 1 0 830 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1333_
timestamp 0
transform 1 0 1110 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1334_
timestamp 0
transform -1 0 2010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1335_
timestamp 0
transform 1 0 1710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1336_
timestamp 0
transform -1 0 1850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1337_
timestamp 0
transform -1 0 1790 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1338_
timestamp 0
transform 1 0 1370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1339_
timestamp 0
transform 1 0 1890 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1340_
timestamp 0
transform -1 0 1490 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1341_
timestamp 0
transform -1 0 1530 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1342_
timestamp 0
transform 1 0 1610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1343_
timestamp 0
transform 1 0 1850 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1344_
timestamp 0
transform -1 0 1990 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1345_
timestamp 0
transform -1 0 1410 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1346_
timestamp 0
transform -1 0 1510 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1347_
timestamp 0
transform 1 0 1610 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1348_
timestamp 0
transform 1 0 1890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1349_
timestamp 0
transform 1 0 3050 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1350_
timestamp 0
transform 1 0 2910 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1351_
timestamp 0
transform 1 0 2350 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1352_
timestamp 0
transform -1 0 1770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1353_
timestamp 0
transform 1 0 1710 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1354_
timestamp 0
transform 1 0 1810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1355_
timestamp 0
transform 1 0 4730 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1356_
timestamp 0
transform 1 0 4810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1357_
timestamp 0
transform -1 0 4630 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1358_
timestamp 0
transform -1 0 4250 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1359_
timestamp 0
transform -1 0 2770 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1360_
timestamp 0
transform -1 0 2630 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1361_
timestamp 0
transform -1 0 2490 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1362_
timestamp 0
transform -1 0 3830 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1363_
timestamp 0
transform -1 0 3950 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1364_
timestamp 0
transform -1 0 5390 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1365_
timestamp 0
transform -1 0 5610 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1366_
timestamp 0
transform 1 0 5490 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1367_
timestamp 0
transform 1 0 4990 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1368_
timestamp 0
transform 1 0 4050 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1369_
timestamp 0
transform -1 0 3370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1370_
timestamp 0
transform -1 0 3730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1371_
timestamp 0
transform -1 0 3930 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1372_
timestamp 0
transform -1 0 4870 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1373_
timestamp 0
transform -1 0 4350 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1374_
timestamp 0
transform 1 0 4450 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1375_
timestamp 0
transform -1 0 5630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1376_
timestamp 0
transform 1 0 5490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1377_
timestamp 0
transform -1 0 5270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1378_
timestamp 0
transform 1 0 5350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1379_
timestamp 0
transform -1 0 4430 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1380_
timestamp 0
transform 1 0 4530 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1381_
timestamp 0
transform -1 0 4810 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1382_
timestamp 0
transform -1 0 4650 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1383_
timestamp 0
transform -1 0 4290 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1384_
timestamp 0
transform 1 0 5110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1385_
timestamp 0
transform 1 0 5250 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1386_
timestamp 0
transform 1 0 5030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1387_
timestamp 0
transform -1 0 5150 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1388_
timestamp 0
transform -1 0 4910 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1389_
timestamp 0
transform 1 0 4950 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1390_
timestamp 0
transform -1 0 4830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1391_
timestamp 0
transform 1 0 4650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1392_
timestamp 0
transform -1 0 5010 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1393_
timestamp 0
transform -1 0 4450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1394_
timestamp 0
transform -1 0 4690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1395_
timestamp 0
transform -1 0 4310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1396_
timestamp 0
transform 1 0 3070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1397_
timestamp 0
transform -1 0 3190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1398_
timestamp 0
transform -1 0 2950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1399_
timestamp 0
transform 1 0 2770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1400_
timestamp 0
transform 1 0 3290 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1401_
timestamp 0
transform 1 0 3310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1402_
timestamp 0
transform -1 0 3590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1403_
timestamp 0
transform -1 0 3470 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1404_
timestamp 0
transform -1 0 3430 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1405_
timestamp 0
transform -1 0 4570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1406_
timestamp 0
transform 1 0 3030 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1407_
timestamp 0
transform -1 0 4750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1408_
timestamp 0
transform 1 0 4590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1409_
timestamp 0
transform -1 0 4470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1410_
timestamp 0
transform -1 0 4010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1411_
timestamp 0
transform 1 0 3850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1412_
timestamp 0
transform 1 0 3390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1413_
timestamp 0
transform 1 0 3310 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1414_
timestamp 0
transform 1 0 3170 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1415_
timestamp 0
transform 1 0 3190 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1416_
timestamp 0
transform 1 0 4510 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1417_
timestamp 0
transform 1 0 4010 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1418_
timestamp 0
transform -1 0 2430 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1419_
timestamp 0
transform 1 0 2490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1420_
timestamp 0
transform -1 0 2630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1421_
timestamp 0
transform -1 0 2410 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1422_
timestamp 0
transform 1 0 2510 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1423_
timestamp 0
transform -1 0 3610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1424_
timestamp 0
transform 1 0 3210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1425_
timestamp 0
transform -1 0 3830 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1426_
timestamp 0
transform 1 0 3670 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1427_
timestamp 0
transform -1 0 2870 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1428_
timestamp 0
transform -1 0 3390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1429_
timestamp 0
transform 1 0 3230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1430_
timestamp 0
transform -1 0 2730 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1431_
timestamp 0
transform -1 0 2870 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1432_
timestamp 0
transform -1 0 2590 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1433_
timestamp 0
transform -1 0 2730 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1434_
timestamp 0
transform -1 0 2990 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1435_
timestamp 0
transform -1 0 3130 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1436_
timestamp 0
transform 1 0 3130 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1437_
timestamp 0
transform -1 0 3510 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1438_
timestamp 0
transform -1 0 1130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1439_
timestamp 0
transform -1 0 1250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1440_
timestamp 0
transform -1 0 3770 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1441_
timestamp 0
transform -1 0 3890 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1442_
timestamp 0
transform -1 0 3290 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1443_
timestamp 0
transform 1 0 3410 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1444_
timestamp 0
transform 1 0 2630 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1445_
timestamp 0
transform -1 0 2510 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1446_
timestamp 0
transform 1 0 2450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1447_
timestamp 0
transform 1 0 2310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1448_
timestamp 0
transform 1 0 3670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1449_
timestamp 0
transform 1 0 3050 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1450_
timestamp 0
transform 1 0 3510 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1451_
timestamp 0
transform -1 0 3550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1527_
timestamp 0
transform -1 0 30 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1528_
timestamp 0
transform 1 0 2370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1529_
timestamp 0
transform -1 0 2510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1530_
timestamp 0
transform 1 0 5690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1531_
timestamp 0
transform 1 0 5570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1532_
timestamp 0
transform -1 0 2010 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1533_
timestamp 0
transform 1 0 2770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1534_
timestamp 0
transform 1 0 2130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1535_
timestamp 0
transform -1 0 2810 0 1 4950
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert0
timestamp 0
transform 1 0 750 0 1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert1
timestamp 0
transform 1 0 4470 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert2
timestamp 0
transform 1 0 2290 0 1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert3
timestamp 0
transform -1 0 1590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert4
timestamp 0
transform -1 0 730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert5
timestamp 0
transform 1 0 4630 0 1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert6
timestamp 0
transform 1 0 3430 0 1 3910
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert15
timestamp 0
transform 1 0 2730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert16
timestamp 0
transform 1 0 1790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert17
timestamp 0
transform -1 0 2570 0 1 790
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert18
timestamp 0
transform -1 0 2010 0 1 1830
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert19
timestamp 0
transform 1 0 2390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert20
timestamp 0
transform -1 0 1470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert21
timestamp 0
transform 1 0 3230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert22
timestamp 0
transform -1 0 1290 0 1 4430
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert23
timestamp 0
transform -1 0 2930 0 1 4430
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert24
timestamp 0
transform 1 0 3550 0 1 3910
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert25
timestamp 0
transform -1 0 3610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert26
timestamp 0
transform -1 0 3570 0 1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert27
timestamp 0
transform -1 0 3250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert28
timestamp 0
transform -1 0 2890 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert29
timestamp 0
transform -1 0 1990 0 1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert30
timestamp 0
transform -1 0 1870 0 1 1310
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert31
timestamp 0
transform 1 0 3590 0 1 1310
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert32
timestamp 0
transform 1 0 2610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert33
timestamp 0
transform -1 0 1650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert7
timestamp 0
transform -1 0 1250 0 1 3390
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert8
timestamp 0
transform -1 0 1590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert9
timestamp 0
transform 1 0 4050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert10
timestamp 0
transform -1 0 3530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert11
timestamp 0
transform -1 0 870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert12
timestamp 0
transform 1 0 3510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert13
timestamp 0
transform 1 0 4230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert14
timestamp 0
transform 1 0 2230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__723_
timestamp 0
transform 1 0 2690 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__724_
timestamp 0
transform -1 0 2610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__725_
timestamp 0
transform -1 0 2310 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__726_
timestamp 0
transform -1 0 2310 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__727_
timestamp 0
transform 1 0 3030 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__728_
timestamp 0
transform -1 0 3670 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__729_
timestamp 0
transform -1 0 970 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__730_
timestamp 0
transform -1 0 2170 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__731_
timestamp 0
transform -1 0 2250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__732_
timestamp 0
transform -1 0 4150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__733_
timestamp 0
transform 1 0 3290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__734_
timestamp 0
transform 1 0 3150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__735_
timestamp 0
transform -1 0 1130 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__736_
timestamp 0
transform -1 0 2570 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__737_
timestamp 0
transform -1 0 2710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__738_
timestamp 0
transform 1 0 2470 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__739_
timestamp 0
transform 1 0 2330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__740_
timestamp 0
transform -1 0 1890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__741_
timestamp 0
transform -1 0 2110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__742_
timestamp 0
transform 1 0 2730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__743_
timestamp 0
transform -1 0 2930 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__744_
timestamp 0
transform 1 0 1890 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__745_
timestamp 0
transform -1 0 2610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__746_
timestamp 0
transform -1 0 2850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__747_
timestamp 0
transform -1 0 2070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__748_
timestamp 0
transform -1 0 2290 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__749_
timestamp 0
transform -1 0 4710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__750_
timestamp 0
transform 1 0 2670 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__751_
timestamp 0
transform 1 0 2530 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__752_
timestamp 0
transform -1 0 4350 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__753_
timestamp 0
transform -1 0 4110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__754_
timestamp 0
transform 1 0 4190 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__755_
timestamp 0
transform -1 0 4130 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__756_
timestamp 0
transform -1 0 3830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__757_
timestamp 0
transform -1 0 3950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__758_
timestamp 0
transform 1 0 2770 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__759_
timestamp 0
transform -1 0 2910 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__760_
timestamp 0
transform 1 0 3270 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__761_
timestamp 0
transform -1 0 3410 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__762_
timestamp 0
transform -1 0 4130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__763_
timestamp 0
transform 1 0 3970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__764_
timestamp 0
transform 1 0 3670 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__765_
timestamp 0
transform -1 0 3810 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__766_
timestamp 0
transform 1 0 370 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__767_
timestamp 0
transform -1 0 2690 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__768_
timestamp 0
transform 1 0 710 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__769_
timestamp 0
transform -1 0 290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__770_
timestamp 0
transform 1 0 750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__771_
timestamp 0
transform 1 0 610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__772_
timestamp 0
transform 1 0 2050 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__773_
timestamp 0
transform 1 0 2550 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__774_
timestamp 0
transform 1 0 2170 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__775_
timestamp 0
transform 1 0 390 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__776_
timestamp 0
transform 1 0 2230 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__777_
timestamp 0
transform 1 0 630 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__778_
timestamp 0
transform 1 0 30 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__779_
timestamp 0
transform 1 0 310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__780_
timestamp 0
transform 1 0 150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__781_
timestamp 0
transform 1 0 1170 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__782_
timestamp 0
transform 1 0 2430 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__783_
timestamp 0
transform 1 0 1510 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__784_
timestamp 0
transform -1 0 1310 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__785_
timestamp 0
transform 1 0 2110 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__786_
timestamp 0
transform 1 0 1630 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__787_
timestamp 0
transform 1 0 2270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__788_
timestamp 0
transform 1 0 2750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__789_
timestamp 0
transform 1 0 2610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__790_
timestamp 0
transform 1 0 1370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__791_
timestamp 0
transform 1 0 1610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__792_
timestamp 0
transform 1 0 1470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__793_
timestamp 0
transform 1 0 1970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__794_
timestamp 0
transform 1 0 2470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__795_
timestamp 0
transform -1 0 2330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__796_
timestamp 0
transform -1 0 4750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__797_
timestamp 0
transform -1 0 4450 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__798_
timestamp 0
transform -1 0 4570 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__799_
timestamp 0
transform -1 0 5390 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__800_
timestamp 0
transform -1 0 4330 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__801_
timestamp 0
transform -1 0 5250 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__802_
timestamp 0
transform -1 0 5730 0 1 270
box -6 -8 26 268
use FILL  FILL_1__803_
timestamp 0
transform -1 0 5530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__804_
timestamp 0
transform 1 0 5390 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__805_
timestamp 0
transform 1 0 5270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__806_
timestamp 0
transform -1 0 4390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__807_
timestamp 0
transform -1 0 4570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__808_
timestamp 0
transform -1 0 3690 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__809_
timestamp 0
transform 1 0 3110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__810_
timestamp 0
transform 1 0 3050 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__811_
timestamp 0
transform -1 0 3750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__812_
timestamp 0
transform -1 0 4430 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__813_
timestamp 0
transform 1 0 3730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__814_
timestamp 0
transform 1 0 610 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__815_
timestamp 0
transform -1 0 2050 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__816_
timestamp 0
transform 1 0 710 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__817_
timestamp 0
transform 1 0 1130 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__818_
timestamp 0
transform 1 0 1550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__819_
timestamp 0
transform -1 0 1710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__820_
timestamp 0
transform 1 0 1470 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__821_
timestamp 0
transform 1 0 970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__822_
timestamp 0
transform -1 0 1350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__823_
timestamp 0
transform -1 0 1450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__824_
timestamp 0
transform 1 0 1490 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__825_
timestamp 0
transform 1 0 1310 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__826_
timestamp 0
transform -1 0 1110 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__827_
timestamp 0
transform 1 0 1610 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__828_
timestamp 0
transform 1 0 1210 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__829_
timestamp 0
transform 1 0 1310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__830_
timestamp 0
transform -1 0 1550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__831_
timestamp 0
transform 1 0 1670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__832_
timestamp 0
transform -1 0 1430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__833_
timestamp 0
transform 1 0 1810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__834_
timestamp 0
transform 1 0 1770 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__835_
timestamp 0
transform -1 0 1950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__836_
timestamp 0
transform 1 0 1870 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__837_
timestamp 0
transform -1 0 1370 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__838_
timestamp 0
transform -1 0 1310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__839_
timestamp 0
transform -1 0 910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__840_
timestamp 0
transform -1 0 1170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__841_
timestamp 0
transform -1 0 1010 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__842_
timestamp 0
transform 1 0 1890 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__843_
timestamp 0
transform -1 0 1790 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__844_
timestamp 0
transform 1 0 1650 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__845_
timestamp 0
transform 1 0 390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__846_
timestamp 0
transform -1 0 2170 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__847_
timestamp 0
transform -1 0 970 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__848_
timestamp 0
transform -1 0 1470 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__849_
timestamp 0
transform 1 0 1070 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__850_
timestamp 0
transform -1 0 970 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__851_
timestamp 0
transform -1 0 1230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__852_
timestamp 0
transform -1 0 690 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__853_
timestamp 0
transform -1 0 890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__854_
timestamp 0
transform 1 0 1070 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__855_
timestamp 0
transform -1 0 1210 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__856_
timestamp 0
transform 1 0 470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__857_
timestamp 0
transform -1 0 550 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__858_
timestamp 0
transform 1 0 670 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__859_
timestamp 0
transform -1 0 1190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__860_
timestamp 0
transform -1 0 830 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__861_
timestamp 0
transform 1 0 1930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__862_
timestamp 0
transform -1 0 1750 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__863_
timestamp 0
transform -1 0 2830 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__864_
timestamp 0
transform -1 0 2710 0 1 790
box -6 -8 26 268
use FILL  FILL_1__865_
timestamp 0
transform -1 0 2010 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__866_
timestamp 0
transform -1 0 1610 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__867_
timestamp 0
transform 1 0 1030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__868_
timestamp 0
transform 1 0 810 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__869_
timestamp 0
transform -1 0 450 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__870_
timestamp 0
transform -1 0 630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__871_
timestamp 0
transform -1 0 890 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__872_
timestamp 0
transform 1 0 530 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__873_
timestamp 0
transform -1 0 630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__874_
timestamp 0
transform -1 0 770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__875_
timestamp 0
transform 1 0 330 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__876_
timestamp 0
transform 1 0 450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__877_
timestamp 0
transform -1 0 50 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__878_
timestamp 0
transform -1 0 330 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__879_
timestamp 0
transform -1 0 490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__880_
timestamp 0
transform -1 0 410 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__881_
timestamp 0
transform -1 0 610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__882_
timestamp 0
transform 1 0 1570 0 1 790
box -6 -8 26 268
use FILL  FILL_1__883_
timestamp 0
transform 1 0 1170 0 1 790
box -6 -8 26 268
use FILL  FILL_1__884_
timestamp 0
transform 1 0 1370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__885_
timestamp 0
transform -1 0 990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__886_
timestamp 0
transform 1 0 1290 0 1 790
box -6 -8 26 268
use FILL  FILL_1__887_
timestamp 0
transform -1 0 850 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__888_
timestamp 0
transform -1 0 890 0 1 790
box -6 -8 26 268
use FILL  FILL_1__889_
timestamp 0
transform -1 0 2330 0 1 790
box -6 -8 26 268
use FILL  FILL_1__890_
timestamp 0
transform 1 0 930 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__891_
timestamp 0
transform 1 0 730 0 1 790
box -6 -8 26 268
use FILL  FILL_1__892_
timestamp 0
transform -1 0 610 0 1 790
box -6 -8 26 268
use FILL  FILL_1__893_
timestamp 0
transform -1 0 750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__894_
timestamp 0
transform -1 0 1030 0 1 790
box -6 -8 26 268
use FILL  FILL_1__895_
timestamp 0
transform -1 0 710 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__896_
timestamp 0
transform -1 0 430 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__897_
timestamp 0
transform 1 0 2690 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__898_
timestamp 0
transform 1 0 2170 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__899_
timestamp 0
transform 1 0 4230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__900_
timestamp 0
transform -1 0 2290 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__901_
timestamp 0
transform 1 0 2170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__902_
timestamp 0
transform -1 0 2150 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__903_
timestamp 0
transform 1 0 310 0 1 790
box -6 -8 26 268
use FILL  FILL_1__904_
timestamp 0
transform -1 0 570 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__905_
timestamp 0
transform -1 0 470 0 1 790
box -6 -8 26 268
use FILL  FILL_1__906_
timestamp 0
transform 1 0 30 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__907_
timestamp 0
transform 1 0 170 0 1 790
box -6 -8 26 268
use FILL  FILL_1__908_
timestamp 0
transform -1 0 350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__909_
timestamp 0
transform 1 0 350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__910_
timestamp 0
transform -1 0 230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__911_
timestamp 0
transform -1 0 50 0 1 790
box -6 -8 26 268
use FILL  FILL_1__912_
timestamp 0
transform -1 0 310 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__913_
timestamp 0
transform 1 0 150 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__914_
timestamp 0
transform 1 0 30 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__915_
timestamp 0
transform 1 0 170 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__916_
timestamp 0
transform 1 0 190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__917_
timestamp 0
transform 1 0 30 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__918_
timestamp 0
transform 1 0 2830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__919_
timestamp 0
transform 1 0 750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__920_
timestamp 0
transform 1 0 150 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__921_
timestamp 0
transform 1 0 130 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__922_
timestamp 0
transform 1 0 2410 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__923_
timestamp 0
transform 1 0 2030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__924_
timestamp 0
transform 1 0 2170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__925_
timestamp 0
transform 1 0 3870 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__926_
timestamp 0
transform -1 0 2710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__927_
timestamp 0
transform 1 0 2550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__928_
timestamp 0
transform -1 0 2470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__929_
timestamp 0
transform 1 0 2330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__930_
timestamp 0
transform -1 0 2570 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__931_
timestamp 0
transform -1 0 2410 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__932_
timestamp 0
transform -1 0 2150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__933_
timestamp 0
transform 1 0 1050 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__934_
timestamp 0
transform 1 0 1090 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__935_
timestamp 0
transform 1 0 1530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__936_
timestamp 0
transform -1 0 1990 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__937_
timestamp 0
transform -1 0 2210 0 1 790
box -6 -8 26 268
use FILL  FILL_1__938_
timestamp 0
transform -1 0 1450 0 1 790
box -6 -8 26 268
use FILL  FILL_1__939_
timestamp 0
transform -1 0 1390 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__940_
timestamp 0
transform -1 0 1730 0 1 790
box -6 -8 26 268
use FILL  FILL_1__941_
timestamp 0
transform -1 0 2810 0 1 790
box -6 -8 26 268
use FILL  FILL_1__942_
timestamp 0
transform 1 0 1810 0 1 790
box -6 -8 26 268
use FILL  FILL_1__943_
timestamp 0
transform -1 0 2450 0 1 790
box -6 -8 26 268
use FILL  FILL_1__944_
timestamp 0
transform -1 0 1550 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__945_
timestamp 0
transform -1 0 1210 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__946_
timestamp 0
transform -1 0 1690 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__947_
timestamp 0
transform -1 0 1230 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__948_
timestamp 0
transform -1 0 1070 0 1 270
box -6 -8 26 268
use FILL  FILL_1__949_
timestamp 0
transform -1 0 970 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__950_
timestamp 0
transform -1 0 2010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__951_
timestamp 0
transform 1 0 1330 0 1 270
box -6 -8 26 268
use FILL  FILL_1__952_
timestamp 0
transform -1 0 1210 0 1 270
box -6 -8 26 268
use FILL  FILL_1__953_
timestamp 0
transform -1 0 790 0 1 270
box -6 -8 26 268
use FILL  FILL_1__954_
timestamp 0
transform -1 0 350 0 1 270
box -6 -8 26 268
use FILL  FILL_1__955_
timestamp 0
transform -1 0 290 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__956_
timestamp 0
transform -1 0 930 0 1 270
box -6 -8 26 268
use FILL  FILL_1__957_
timestamp 0
transform -1 0 830 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__958_
timestamp 0
transform -1 0 650 0 1 270
box -6 -8 26 268
use FILL  FILL_1__959_
timestamp 0
transform -1 0 210 0 1 270
box -6 -8 26 268
use FILL  FILL_1__960_
timestamp 0
transform -1 0 410 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__961_
timestamp 0
transform -1 0 510 0 1 270
box -6 -8 26 268
use FILL  FILL_1__962_
timestamp 0
transform -1 0 50 0 1 270
box -6 -8 26 268
use FILL  FILL_1__963_
timestamp 0
transform -1 0 50 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__964_
timestamp 0
transform 1 0 30 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__965_
timestamp 0
transform 1 0 30 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__966_
timestamp 0
transform -1 0 850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__967_
timestamp 0
transform -1 0 970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__968_
timestamp 0
transform 1 0 1090 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__969_
timestamp 0
transform 1 0 150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__970_
timestamp 0
transform 1 0 530 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__971_
timestamp 0
transform -1 0 690 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__972_
timestamp 0
transform 1 0 2810 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__973_
timestamp 0
transform 1 0 2250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__974_
timestamp 0
transform 1 0 2270 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__975_
timestamp 0
transform 1 0 1750 0 1 270
box -6 -8 26 268
use FILL  FILL_1__976_
timestamp 0
transform 1 0 1850 0 1 270
box -6 -8 26 268
use FILL  FILL_1__977_
timestamp 0
transform 1 0 2930 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__978_
timestamp 0
transform -1 0 3370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__979_
timestamp 0
transform 1 0 3210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__980_
timestamp 0
transform -1 0 3490 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__981_
timestamp 0
transform -1 0 3510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__982_
timestamp 0
transform -1 0 3090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__983_
timestamp 0
transform -1 0 2990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__984_
timestamp 0
transform -1 0 3350 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__985_
timestamp 0
transform -1 0 2950 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__986_
timestamp 0
transform 1 0 3070 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__987_
timestamp 0
transform -1 0 2890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__988_
timestamp 0
transform -1 0 2090 0 1 790
box -6 -8 26 268
use FILL  FILL_1__989_
timestamp 0
transform 1 0 1930 0 1 790
box -6 -8 26 268
use FILL  FILL_1__990_
timestamp 0
transform 1 0 3750 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__991_
timestamp 0
transform -1 0 3150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__992_
timestamp 0
transform -1 0 3430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__993_
timestamp 0
transform -1 0 3750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__994_
timestamp 0
transform -1 0 3810 0 1 790
box -6 -8 26 268
use FILL  FILL_1__995_
timestamp 0
transform -1 0 3530 0 1 790
box -6 -8 26 268
use FILL  FILL_1__996_
timestamp 0
transform -1 0 3390 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__997_
timestamp 0
transform -1 0 3750 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__998_
timestamp 0
transform 1 0 3630 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__999_
timestamp 0
transform -1 0 3270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1000_
timestamp 0
transform -1 0 3250 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1001_
timestamp 0
transform -1 0 2670 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1002_
timestamp 0
transform -1 0 2130 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1003_
timestamp 0
transform 1 0 1810 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1004_
timestamp 0
transform 1 0 3210 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1005_
timestamp 0
transform -1 0 3390 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1006_
timestamp 0
transform -1 0 2950 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1007_
timestamp 0
transform 1 0 2510 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1008_
timestamp 0
transform 1 0 2990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1009_
timestamp 0
transform 1 0 2930 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1010_
timestamp 0
transform -1 0 3090 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1011_
timestamp 0
transform -1 0 3150 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1012_
timestamp 0
transform -1 0 2590 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1013_
timestamp 0
transform 1 0 1470 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1014_
timestamp 0
transform 1 0 1610 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1015_
timestamp 0
transform -1 0 3010 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1016_
timestamp 0
transform -1 0 2390 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1017_
timestamp 0
transform -1 0 2310 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1018_
timestamp 0
transform -1 0 2010 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1019_
timestamp 0
transform -1 0 2730 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1020_
timestamp 0
transform 1 0 2430 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1021_
timestamp 0
transform -1 0 2490 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1022_
timestamp 0
transform 1 0 1790 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1023_
timestamp 0
transform -1 0 1470 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1024_
timestamp 0
transform 1 0 1330 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1025_
timestamp 0
transform 1 0 1910 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1026_
timestamp 0
transform 1 0 30 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1027_
timestamp 0
transform 1 0 250 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1028_
timestamp 0
transform -1 0 2350 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1029_
timestamp 0
transform 1 0 2150 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1030_
timestamp 0
transform -1 0 2210 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1031_
timestamp 0
transform -1 0 2070 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1032_
timestamp 0
transform 1 0 1350 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1033_
timestamp 0
transform 1 0 1190 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1034_
timestamp 0
transform 1 0 1630 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1035_
timestamp 0
transform -1 0 2770 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1036_
timestamp 0
transform 1 0 2610 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1037_
timestamp 0
transform -1 0 3230 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1038_
timestamp 0
transform 1 0 3790 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1039_
timestamp 0
transform 1 0 3290 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1040_
timestamp 0
transform 1 0 3390 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1041_
timestamp 0
transform 1 0 3990 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1042_
timestamp 0
transform 1 0 3730 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1043_
timestamp 0
transform -1 0 4310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1044_
timestamp 0
transform 1 0 3450 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1045_
timestamp 0
transform 1 0 3590 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1046_
timestamp 0
transform 1 0 4150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1047_
timestamp 0
transform -1 0 4070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1048_
timestamp 0
transform 1 0 3870 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1049_
timestamp 0
transform -1 0 3650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1050_
timestamp 0
transform -1 0 3790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1051_
timestamp 0
transform -1 0 3930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1052_
timestamp 0
transform -1 0 4790 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1053_
timestamp 0
transform -1 0 3490 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1054_
timestamp 0
transform 1 0 3930 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1055_
timestamp 0
transform 1 0 4790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1056_
timestamp 0
transform 1 0 4910 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1057_
timestamp 0
transform -1 0 4410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1058_
timestamp 0
transform -1 0 4450 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1059_
timestamp 0
transform 1 0 4050 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1060_
timestamp 0
transform -1 0 4150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1061_
timestamp 0
transform -1 0 4290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1062_
timestamp 0
transform 1 0 4570 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1063_
timestamp 0
transform 1 0 4290 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1064_
timestamp 0
transform 1 0 4330 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1065_
timestamp 0
transform -1 0 3590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1066_
timestamp 0
transform -1 0 3670 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1067_
timestamp 0
transform -1 0 4170 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1068_
timestamp 0
transform 1 0 3970 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1069_
timestamp 0
transform 1 0 3850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1070_
timestamp 0
transform 1 0 3990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1071_
timestamp 0
transform -1 0 4010 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1072_
timestamp 0
transform -1 0 4510 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1073_
timestamp 0
transform 1 0 4790 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1074_
timestamp 0
transform 1 0 4430 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1075_
timestamp 0
transform 1 0 4150 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1076_
timestamp 0
transform -1 0 4950 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1077_
timestamp 0
transform -1 0 4250 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1078_
timestamp 0
transform 1 0 2790 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1079_
timestamp 0
transform 1 0 3070 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1080_
timestamp 0
transform -1 0 4670 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1081_
timestamp 0
transform 1 0 4630 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1082_
timestamp 0
transform -1 0 4390 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1083_
timestamp 0
transform -1 0 3970 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1084_
timestamp 0
transform -1 0 4210 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1085_
timestamp 0
transform -1 0 4530 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1086_
timestamp 0
transform -1 0 3830 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1087_
timestamp 0
transform -1 0 3670 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1088_
timestamp 0
transform -1 0 2870 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1089_
timestamp 0
transform 1 0 2850 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1090_
timestamp 0
transform -1 0 3670 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1091_
timestamp 0
transform -1 0 4110 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1092_
timestamp 0
transform -1 0 3530 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1093_
timestamp 0
transform 1 0 3390 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1094_
timestamp 0
transform 1 0 1790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1095_
timestamp 0
transform 1 0 2150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1096_
timestamp 0
transform 1 0 2010 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1097_
timestamp 0
transform 1 0 3770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1098_
timestamp 0
transform -1 0 3150 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1099_
timestamp 0
transform -1 0 3550 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1100_
timestamp 0
transform 1 0 3410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1101_
timestamp 0
transform -1 0 4070 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1102_
timestamp 0
transform 1 0 3890 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1103_
timestamp 0
transform 1 0 3870 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1104_
timestamp 0
transform -1 0 5730 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1105_
timestamp 0
transform -1 0 5230 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1106_
timestamp 0
transform 1 0 5070 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1107_
timestamp 0
transform 1 0 4250 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1108_
timestamp 0
transform -1 0 4450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1109_
timestamp 0
transform 1 0 5230 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1110_
timestamp 0
transform 1 0 5070 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1111_
timestamp 0
transform 1 0 5390 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1112_
timestamp 0
transform -1 0 5670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1113_
timestamp 0
transform 1 0 4670 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1114_
timestamp 0
transform 1 0 4490 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1115_
timestamp 0
transform 1 0 4550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1116_
timestamp 0
transform 1 0 4370 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1117_
timestamp 0
transform 1 0 4210 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1118_
timestamp 0
transform 1 0 4610 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1119_
timestamp 0
transform -1 0 5370 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1120_
timestamp 0
transform 1 0 4550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1121_
timestamp 0
transform -1 0 4770 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1122_
timestamp 0
transform -1 0 5210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1123_
timestamp 0
transform 1 0 5610 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1124_
timestamp 0
transform -1 0 5470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1125_
timestamp 0
transform 1 0 5050 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1126_
timestamp 0
transform -1 0 5250 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1127_
timestamp 0
transform 1 0 5410 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1128_
timestamp 0
transform -1 0 5590 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1129_
timestamp 0
transform -1 0 4310 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1130_
timestamp 0
transform 1 0 5150 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1131_
timestamp 0
transform -1 0 5290 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1132_
timestamp 0
transform -1 0 4830 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1133_
timestamp 0
transform 1 0 4950 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1134_
timestamp 0
transform 1 0 5090 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1135_
timestamp 0
transform 1 0 5130 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1136_
timestamp 0
transform -1 0 5450 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1137_
timestamp 0
transform -1 0 5570 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1138_
timestamp 0
transform -1 0 5010 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1139_
timestamp 0
transform 1 0 4850 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1140_
timestamp 0
transform 1 0 4990 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1141_
timestamp 0
transform 1 0 4890 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1142_
timestamp 0
transform -1 0 4730 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1143_
timestamp 0
transform -1 0 5310 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1144_
timestamp 0
transform -1 0 4590 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1145_
timestamp 0
transform -1 0 4270 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1146_
timestamp 0
transform 1 0 4190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1147_
timestamp 0
transform -1 0 3790 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1148_
timestamp 0
transform 1 0 4010 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1149_
timestamp 0
transform -1 0 4130 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1150_
timestamp 0
transform 1 0 5530 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1151_
timestamp 0
transform 1 0 5630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1152_
timestamp 0
transform -1 0 5330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1153_
timestamp 0
transform 1 0 4350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1154_
timestamp 0
transform 1 0 4130 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1155_
timestamp 0
transform 1 0 4470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1156_
timestamp 0
transform 1 0 4610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1157_
timestamp 0
transform 1 0 4210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1158_
timestamp 0
transform 1 0 4750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1159_
timestamp 0
transform -1 0 5210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1160_
timestamp 0
transform -1 0 4450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1161_
timestamp 0
transform -1 0 4910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1162_
timestamp 0
transform 1 0 4350 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1163_
timestamp 0
transform -1 0 4530 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1164_
timestamp 0
transform 1 0 4790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1165_
timestamp 0
transform 1 0 4670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1166_
timestamp 0
transform 1 0 4770 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1167_
timestamp 0
transform 1 0 5310 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1168_
timestamp 0
transform -1 0 5490 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1169_
timestamp 0
transform 1 0 4630 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1170_
timestamp 0
transform 1 0 4910 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1171_
timestamp 0
transform 1 0 5170 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1172_
timestamp 0
transform -1 0 5470 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1173_
timestamp 0
transform 1 0 5350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1174_
timestamp 0
transform 1 0 5030 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1175_
timestamp 0
transform -1 0 5510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1176_
timestamp 0
transform 1 0 5090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1177_
timestamp 0
transform -1 0 4950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1178_
timestamp 0
transform -1 0 5590 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1179_
timestamp 0
transform -1 0 5450 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1180_
timestamp 0
transform -1 0 5230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1181_
timestamp 0
transform -1 0 4510 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1182_
timestamp 0
transform -1 0 4030 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1183_
timestamp 0
transform -1 0 3970 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1184_
timestamp 0
transform 1 0 3870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1185_
timestamp 0
transform -1 0 4970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1186_
timestamp 0
transform 1 0 4630 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1187_
timestamp 0
transform -1 0 4390 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1188_
timestamp 0
transform -1 0 4890 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1189_
timestamp 0
transform 1 0 4750 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1190_
timestamp 0
transform -1 0 4530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1191_
timestamp 0
transform 1 0 4370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1192_
timestamp 0
transform 1 0 5610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1193_
timestamp 0
transform -1 0 5050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1194_
timestamp 0
transform 1 0 5450 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1195_
timestamp 0
transform 1 0 4930 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1196_
timestamp 0
transform -1 0 4610 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1197_
timestamp 0
transform 1 0 4330 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1198_
timestamp 0
transform 1 0 4710 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1199_
timestamp 0
transform -1 0 4850 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1200_
timestamp 0
transform 1 0 5250 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1201_
timestamp 0
transform 1 0 5450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1202_
timestamp 0
transform 1 0 5310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1203_
timestamp 0
transform -1 0 5710 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1204_
timestamp 0
transform -1 0 5570 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1205_
timestamp 0
transform -1 0 5710 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1206_
timestamp 0
transform 1 0 5690 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1207_
timestamp 0
transform -1 0 5610 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1208_
timestamp 0
transform 1 0 5670 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1209_
timestamp 0
transform -1 0 5550 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1210_
timestamp 0
transform -1 0 5430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1211_
timestamp 0
transform -1 0 5170 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1212_
timestamp 0
transform -1 0 3270 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1213_
timestamp 0
transform 1 0 2990 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1214_
timestamp 0
transform -1 0 3890 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1215_
timestamp 0
transform 1 0 3710 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1216_
timestamp 0
transform -1 0 4930 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1217_
timestamp 0
transform 1 0 4770 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1218_
timestamp 0
transform -1 0 5030 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1219_
timestamp 0
transform 1 0 4930 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1220_
timestamp 0
transform -1 0 5090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1221_
timestamp 0
transform -1 0 5670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1222_
timestamp 0
transform 1 0 5150 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1223_
timestamp 0
transform 1 0 4970 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1224_
timestamp 0
transform 1 0 4690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1225_
timestamp 0
transform 1 0 4470 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1226_
timestamp 0
transform 1 0 4830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1227_
timestamp 0
transform 1 0 5070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1228_
timestamp 0
transform 1 0 5210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1229_
timestamp 0
transform -1 0 5490 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1230_
timestamp 0
transform 1 0 5530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1231_
timestamp 0
transform 1 0 5710 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1232_
timestamp 0
transform -1 0 5730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1233_
timestamp 0
transform 1 0 5530 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1234_
timestamp 0
transform -1 0 5690 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1235_
timestamp 0
transform 1 0 5650 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1236_
timestamp 0
transform 1 0 5190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1237_
timestamp 0
transform 1 0 5730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1238_
timestamp 0
transform -1 0 5410 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1239_
timestamp 0
transform -1 0 5270 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1240_
timestamp 0
transform -1 0 5330 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1241_
timestamp 0
transform -1 0 5290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1242_
timestamp 0
transform -1 0 5150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1243_
timestamp 0
transform 1 0 5350 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1244_
timestamp 0
transform 1 0 4550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1245_
timestamp 0
transform 1 0 4930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1246_
timestamp 0
transform 1 0 5130 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1247_
timestamp 0
transform -1 0 5010 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1248_
timestamp 0
transform 1 0 4990 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1249_
timestamp 0
transform -1 0 5410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1250_
timestamp 0
transform -1 0 4630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1251_
timestamp 0
transform 1 0 4850 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1252_
timestamp 0
transform 1 0 4710 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1253_
timestamp 0
transform -1 0 5430 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1254_
timestamp 0
transform -1 0 5290 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1255_
timestamp 0
transform -1 0 5330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1256_
timestamp 0
transform -1 0 5190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1257_
timestamp 0
transform 1 0 5250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1258_
timestamp 0
transform 1 0 5110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1259_
timestamp 0
transform 1 0 5070 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1260_
timestamp 0
transform -1 0 170 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1261_
timestamp 0
transform 1 0 30 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1262_
timestamp 0
transform 1 0 270 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1263_
timestamp 0
transform -1 0 410 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1264_
timestamp 0
transform -1 0 1030 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1265_
timestamp 0
transform 1 0 510 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1266_
timestamp 0
transform -1 0 810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1267_
timestamp 0
transform 1 0 530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1268_
timestamp 0
transform 1 0 310 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1269_
timestamp 0
transform -1 0 170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1270_
timestamp 0
transform 1 0 30 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1271_
timestamp 0
transform 1 0 270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1272_
timestamp 0
transform 1 0 410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1273_
timestamp 0
transform 1 0 830 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1274_
timestamp 0
transform 1 0 450 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1275_
timestamp 0
transform -1 0 670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1276_
timestamp 0
transform -1 0 1830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1277_
timestamp 0
transform 1 0 1610 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1278_
timestamp 0
transform 1 0 2030 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1279_
timestamp 0
transform 1 0 1730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1280_
timestamp 0
transform -1 0 1950 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1281_
timestamp 0
transform 1 0 1790 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1282_
timestamp 0
transform 1 0 270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1283_
timestamp 0
transform -1 0 510 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1284_
timestamp 0
transform 1 0 670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1285_
timestamp 0
transform -1 0 810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1286_
timestamp 0
transform -1 0 1490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1287_
timestamp 0
transform 1 0 1330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1288_
timestamp 0
transform -1 0 210 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1289_
timestamp 0
transform -1 0 50 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1290_
timestamp 0
transform 1 0 30 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1291_
timestamp 0
transform 1 0 30 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1292_
timestamp 0
transform 1 0 310 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1293_
timestamp 0
transform -1 0 590 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1294_
timestamp 0
transform 1 0 430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1295_
timestamp 0
transform -1 0 170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1296_
timestamp 0
transform -1 0 50 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1297_
timestamp 0
transform 1 0 190 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1298_
timestamp 0
transform -1 0 270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1299_
timestamp 0
transform 1 0 30 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1300_
timestamp 0
transform -1 0 670 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1301_
timestamp 0
transform 1 0 150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1302_
timestamp 0
transform -1 0 690 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1303_
timestamp 0
transform -1 0 830 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1304_
timestamp 0
transform 1 0 530 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1305_
timestamp 0
transform -1 0 390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1306_
timestamp 0
transform 1 0 290 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1307_
timestamp 0
transform -1 0 650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1308_
timestamp 0
transform -1 0 570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1309_
timestamp 0
transform -1 0 510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1310_
timestamp 0
transform -1 0 1510 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1311_
timestamp 0
transform 1 0 690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1312_
timestamp 0
transform 1 0 850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1313_
timestamp 0
transform -1 0 990 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1314_
timestamp 0
transform -1 0 910 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1315_
timestamp 0
transform 1 0 1030 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1316_
timestamp 0
transform 1 0 1250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1317_
timestamp 0
transform -1 0 1170 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1318_
timestamp 0
transform 1 0 1650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1319_
timestamp 0
transform -1 0 1550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1320_
timestamp 0
transform 1 0 1290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1321_
timestamp 0
transform -1 0 1410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1322_
timestamp 0
transform 1 0 1630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1323_
timestamp 0
transform 1 0 2290 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1324_
timestamp 0
transform 1 0 2150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1325_
timestamp 0
transform -1 0 1690 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1326_
timestamp 0
transform 1 0 410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1327_
timestamp 0
transform -1 0 1050 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1328_
timestamp 0
transform 1 0 1150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1329_
timestamp 0
transform -1 0 1110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1330_
timestamp 0
transform 1 0 990 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1331_
timestamp 0
transform -1 0 430 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1332_
timestamp 0
transform 1 0 850 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1333_
timestamp 0
transform 1 0 1130 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1334_
timestamp 0
transform -1 0 2030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1335_
timestamp 0
transform 1 0 1730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1336_
timestamp 0
transform -1 0 1870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1337_
timestamp 0
transform -1 0 1810 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1338_
timestamp 0
transform 1 0 1390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1339_
timestamp 0
transform 1 0 1910 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1340_
timestamp 0
transform -1 0 1510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1341_
timestamp 0
transform -1 0 1550 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1342_
timestamp 0
transform 1 0 1630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1343_
timestamp 0
transform 1 0 1870 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1344_
timestamp 0
transform -1 0 2010 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1345_
timestamp 0
transform -1 0 1430 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1346_
timestamp 0
transform -1 0 1530 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1347_
timestamp 0
transform 1 0 1630 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1348_
timestamp 0
transform 1 0 1910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1349_
timestamp 0
transform 1 0 3070 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1350_
timestamp 0
transform 1 0 2930 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1351_
timestamp 0
transform 1 0 2370 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1352_
timestamp 0
transform -1 0 1790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1353_
timestamp 0
transform 1 0 1730 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1354_
timestamp 0
transform 1 0 1830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1355_
timestamp 0
transform 1 0 4750 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1356_
timestamp 0
transform 1 0 4830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1357_
timestamp 0
transform -1 0 4650 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1358_
timestamp 0
transform -1 0 4270 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1359_
timestamp 0
transform -1 0 2790 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1360_
timestamp 0
transform -1 0 2650 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1361_
timestamp 0
transform -1 0 2510 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1362_
timestamp 0
transform -1 0 3850 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1363_
timestamp 0
transform -1 0 3970 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1364_
timestamp 0
transform -1 0 5410 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1365_
timestamp 0
transform -1 0 5630 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1366_
timestamp 0
transform 1 0 5510 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1367_
timestamp 0
transform 1 0 5010 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1368_
timestamp 0
transform 1 0 4070 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1369_
timestamp 0
transform -1 0 3390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1370_
timestamp 0
transform -1 0 3750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1371_
timestamp 0
transform -1 0 3950 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1372_
timestamp 0
transform -1 0 4890 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1373_
timestamp 0
transform -1 0 4370 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1374_
timestamp 0
transform 1 0 4470 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1375_
timestamp 0
transform -1 0 5650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1376_
timestamp 0
transform 1 0 5510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1377_
timestamp 0
transform -1 0 5290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1378_
timestamp 0
transform 1 0 5370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1379_
timestamp 0
transform -1 0 4450 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1380_
timestamp 0
transform 1 0 4550 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1381_
timestamp 0
transform -1 0 4830 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1382_
timestamp 0
transform -1 0 4670 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1383_
timestamp 0
transform -1 0 4310 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1384_
timestamp 0
transform 1 0 5130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1385_
timestamp 0
transform 1 0 5270 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1386_
timestamp 0
transform 1 0 5050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1387_
timestamp 0
transform -1 0 5170 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1388_
timestamp 0
transform -1 0 4930 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1389_
timestamp 0
transform 1 0 4970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1390_
timestamp 0
transform -1 0 4850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1391_
timestamp 0
transform 1 0 4670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1392_
timestamp 0
transform -1 0 5030 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1393_
timestamp 0
transform -1 0 4470 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1394_
timestamp 0
transform -1 0 4710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1395_
timestamp 0
transform -1 0 4330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1396_
timestamp 0
transform 1 0 3090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1397_
timestamp 0
transform -1 0 3210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1398_
timestamp 0
transform -1 0 2970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1399_
timestamp 0
transform 1 0 2790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1400_
timestamp 0
transform 1 0 3310 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1401_
timestamp 0
transform 1 0 3330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1402_
timestamp 0
transform -1 0 3610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1403_
timestamp 0
transform -1 0 3490 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1404_
timestamp 0
transform -1 0 3450 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1405_
timestamp 0
transform -1 0 4590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1406_
timestamp 0
transform 1 0 3050 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1407_
timestamp 0
transform -1 0 4770 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1408_
timestamp 0
transform 1 0 4610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1409_
timestamp 0
transform -1 0 4490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1410_
timestamp 0
transform -1 0 4030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1411_
timestamp 0
transform 1 0 3870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1412_
timestamp 0
transform 1 0 3410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1413_
timestamp 0
transform 1 0 3330 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1414_
timestamp 0
transform 1 0 3190 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1415_
timestamp 0
transform 1 0 3210 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1416_
timestamp 0
transform 1 0 4530 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1417_
timestamp 0
transform 1 0 4030 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1418_
timestamp 0
transform -1 0 2450 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1419_
timestamp 0
transform 1 0 2510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1420_
timestamp 0
transform -1 0 2650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1421_
timestamp 0
transform -1 0 2430 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1422_
timestamp 0
transform 1 0 2530 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1423_
timestamp 0
transform -1 0 3630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1424_
timestamp 0
transform 1 0 3230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1425_
timestamp 0
transform -1 0 3850 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1426_
timestamp 0
transform 1 0 3690 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1427_
timestamp 0
transform -1 0 2890 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1428_
timestamp 0
transform -1 0 3410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1429_
timestamp 0
transform 1 0 3250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1430_
timestamp 0
transform -1 0 2750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1431_
timestamp 0
transform -1 0 2890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1432_
timestamp 0
transform -1 0 2610 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1433_
timestamp 0
transform -1 0 2750 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1434_
timestamp 0
transform -1 0 3010 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1435_
timestamp 0
transform -1 0 3150 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1436_
timestamp 0
transform 1 0 3150 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1437_
timestamp 0
transform -1 0 3530 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1438_
timestamp 0
transform -1 0 1150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1439_
timestamp 0
transform -1 0 1270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1440_
timestamp 0
transform -1 0 3790 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1441_
timestamp 0
transform -1 0 3910 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1442_
timestamp 0
transform -1 0 3310 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1443_
timestamp 0
transform 1 0 3430 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1444_
timestamp 0
transform 1 0 2650 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1445_
timestamp 0
transform -1 0 2530 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1446_
timestamp 0
transform 1 0 2470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1447_
timestamp 0
transform 1 0 2330 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1448_
timestamp 0
transform 1 0 3690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1449_
timestamp 0
transform 1 0 3070 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1450_
timestamp 0
transform 1 0 3530 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1451_
timestamp 0
transform -1 0 3570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1527_
timestamp 0
transform -1 0 50 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1528_
timestamp 0
transform 1 0 2390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1529_
timestamp 0
transform -1 0 2530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1530_
timestamp 0
transform 1 0 5710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1531_
timestamp 0
transform 1 0 5590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1532_
timestamp 0
transform -1 0 2030 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1533_
timestamp 0
transform 1 0 2790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1534_
timestamp 0
transform 1 0 2150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1535_
timestamp 0
transform -1 0 2830 0 1 4950
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert0
timestamp 0
transform 1 0 770 0 1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert1
timestamp 0
transform 1 0 4490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert2
timestamp 0
transform 1 0 2310 0 1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert3
timestamp 0
transform -1 0 1610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert4
timestamp 0
transform -1 0 750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert5
timestamp 0
transform 1 0 4650 0 1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert6
timestamp 0
transform 1 0 3450 0 1 3910
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert15
timestamp 0
transform 1 0 2750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert16
timestamp 0
transform 1 0 1810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert17
timestamp 0
transform -1 0 2590 0 1 790
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert18
timestamp 0
transform -1 0 2030 0 1 1830
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert19
timestamp 0
transform 1 0 2410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert20
timestamp 0
transform -1 0 1490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert21
timestamp 0
transform 1 0 3250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert22
timestamp 0
transform -1 0 1310 0 1 4430
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert23
timestamp 0
transform -1 0 2950 0 1 4430
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert24
timestamp 0
transform 1 0 3570 0 1 3910
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert25
timestamp 0
transform -1 0 3630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert26
timestamp 0
transform -1 0 3590 0 1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert27
timestamp 0
transform -1 0 3270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert28
timestamp 0
transform -1 0 2910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert29
timestamp 0
transform -1 0 2010 0 1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert30
timestamp 0
transform -1 0 1890 0 1 1310
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert31
timestamp 0
transform 1 0 3610 0 1 1310
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert32
timestamp 0
transform 1 0 2630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert33
timestamp 0
transform -1 0 1670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert7
timestamp 0
transform -1 0 1270 0 1 3390
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert8
timestamp 0
transform -1 0 1610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert9
timestamp 0
transform 1 0 4070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert10
timestamp 0
transform -1 0 3550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert11
timestamp 0
transform -1 0 890 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert12
timestamp 0
transform 1 0 3530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert13
timestamp 0
transform 1 0 4250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert14
timestamp 0
transform 1 0 2250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__723_
timestamp 0
transform 1 0 2710 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__724_
timestamp 0
transform -1 0 2630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__725_
timestamp 0
transform -1 0 2330 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__726_
timestamp 0
transform -1 0 2330 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__727_
timestamp 0
transform 1 0 3050 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__728_
timestamp 0
transform -1 0 3690 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__729_
timestamp 0
transform -1 0 990 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__730_
timestamp 0
transform -1 0 2190 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__731_
timestamp 0
transform -1 0 2270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__732_
timestamp 0
transform -1 0 4170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__733_
timestamp 0
transform 1 0 3310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__734_
timestamp 0
transform 1 0 3170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__735_
timestamp 0
transform -1 0 1150 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__736_
timestamp 0
transform -1 0 2590 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__737_
timestamp 0
transform -1 0 2730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__738_
timestamp 0
transform 1 0 2490 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__739_
timestamp 0
transform 1 0 2350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__740_
timestamp 0
transform -1 0 1910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__741_
timestamp 0
transform -1 0 2130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__742_
timestamp 0
transform 1 0 2750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__743_
timestamp 0
transform -1 0 2950 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__744_
timestamp 0
transform 1 0 1910 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__745_
timestamp 0
transform -1 0 2630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__746_
timestamp 0
transform -1 0 2870 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__747_
timestamp 0
transform -1 0 2090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__748_
timestamp 0
transform -1 0 2310 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__749_
timestamp 0
transform -1 0 4730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__750_
timestamp 0
transform 1 0 2690 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__751_
timestamp 0
transform 1 0 2550 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__752_
timestamp 0
transform -1 0 4370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__753_
timestamp 0
transform -1 0 4130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__754_
timestamp 0
transform 1 0 4210 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__755_
timestamp 0
transform -1 0 4150 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__756_
timestamp 0
transform -1 0 3850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__757_
timestamp 0
transform -1 0 3970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__758_
timestamp 0
transform 1 0 2790 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__759_
timestamp 0
transform -1 0 2930 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__760_
timestamp 0
transform 1 0 3290 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__761_
timestamp 0
transform -1 0 3430 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__762_
timestamp 0
transform -1 0 4150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__763_
timestamp 0
transform 1 0 3990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__764_
timestamp 0
transform 1 0 3690 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__765_
timestamp 0
transform -1 0 3830 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__766_
timestamp 0
transform 1 0 390 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__767_
timestamp 0
transform -1 0 2710 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__768_
timestamp 0
transform 1 0 730 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__769_
timestamp 0
transform -1 0 310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__770_
timestamp 0
transform 1 0 770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__771_
timestamp 0
transform 1 0 630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__772_
timestamp 0
transform 1 0 2070 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__773_
timestamp 0
transform 1 0 2570 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__774_
timestamp 0
transform 1 0 2190 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__775_
timestamp 0
transform 1 0 410 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__776_
timestamp 0
transform 1 0 2250 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__777_
timestamp 0
transform 1 0 650 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__778_
timestamp 0
transform 1 0 50 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__779_
timestamp 0
transform 1 0 330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__780_
timestamp 0
transform 1 0 170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__781_
timestamp 0
transform 1 0 1190 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__782_
timestamp 0
transform 1 0 2450 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__783_
timestamp 0
transform 1 0 1530 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__784_
timestamp 0
transform -1 0 1330 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__785_
timestamp 0
transform 1 0 2130 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__786_
timestamp 0
transform 1 0 1650 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__787_
timestamp 0
transform 1 0 2290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__788_
timestamp 0
transform 1 0 2770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__789_
timestamp 0
transform 1 0 2630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__790_
timestamp 0
transform 1 0 1390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__791_
timestamp 0
transform 1 0 1630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__792_
timestamp 0
transform 1 0 1490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__793_
timestamp 0
transform 1 0 1990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__794_
timestamp 0
transform 1 0 2490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__795_
timestamp 0
transform -1 0 2350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__796_
timestamp 0
transform -1 0 4770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__797_
timestamp 0
transform -1 0 4470 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__798_
timestamp 0
transform -1 0 4590 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__799_
timestamp 0
transform -1 0 5410 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__800_
timestamp 0
transform -1 0 4350 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__801_
timestamp 0
transform -1 0 5270 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__802_
timestamp 0
transform -1 0 5750 0 1 270
box -6 -8 26 268
use FILL  FILL_2__803_
timestamp 0
transform -1 0 5550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__804_
timestamp 0
transform 1 0 5410 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__805_
timestamp 0
transform 1 0 5290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__806_
timestamp 0
transform -1 0 4410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__807_
timestamp 0
transform -1 0 4590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__808_
timestamp 0
transform -1 0 3710 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__809_
timestamp 0
transform 1 0 3130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__810_
timestamp 0
transform 1 0 3070 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__811_
timestamp 0
transform -1 0 3770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__812_
timestamp 0
transform -1 0 4450 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__813_
timestamp 0
transform 1 0 3750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__814_
timestamp 0
transform 1 0 630 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__815_
timestamp 0
transform -1 0 2070 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__816_
timestamp 0
transform 1 0 730 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__817_
timestamp 0
transform 1 0 1150 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__818_
timestamp 0
transform 1 0 1570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__819_
timestamp 0
transform -1 0 1730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__820_
timestamp 0
transform 1 0 1490 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__821_
timestamp 0
transform 1 0 990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__822_
timestamp 0
transform -1 0 1370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__823_
timestamp 0
transform -1 0 1470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__824_
timestamp 0
transform 1 0 1510 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__825_
timestamp 0
transform 1 0 1330 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__826_
timestamp 0
transform -1 0 1130 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__827_
timestamp 0
transform 1 0 1630 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__828_
timestamp 0
transform 1 0 1230 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__829_
timestamp 0
transform 1 0 1330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__830_
timestamp 0
transform -1 0 1570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__831_
timestamp 0
transform 1 0 1690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__832_
timestamp 0
transform -1 0 1450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__833_
timestamp 0
transform 1 0 1830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__834_
timestamp 0
transform 1 0 1790 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__835_
timestamp 0
transform -1 0 1970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__836_
timestamp 0
transform 1 0 1890 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__837_
timestamp 0
transform -1 0 1390 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__838_
timestamp 0
transform -1 0 1330 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__839_
timestamp 0
transform -1 0 930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__840_
timestamp 0
transform -1 0 1190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__841_
timestamp 0
transform -1 0 1030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__842_
timestamp 0
transform 1 0 1910 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__843_
timestamp 0
transform -1 0 1810 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__844_
timestamp 0
transform 1 0 1670 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__845_
timestamp 0
transform 1 0 410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__846_
timestamp 0
transform -1 0 2190 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__847_
timestamp 0
transform -1 0 990 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__848_
timestamp 0
transform -1 0 1490 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__849_
timestamp 0
transform 1 0 1090 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__850_
timestamp 0
transform -1 0 990 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__851_
timestamp 0
transform -1 0 1250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__852_
timestamp 0
transform -1 0 710 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__853_
timestamp 0
transform -1 0 910 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__854_
timestamp 0
transform 1 0 1090 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__855_
timestamp 0
transform -1 0 1230 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__856_
timestamp 0
transform 1 0 490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__857_
timestamp 0
transform -1 0 570 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__858_
timestamp 0
transform 1 0 690 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__859_
timestamp 0
transform -1 0 1210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__860_
timestamp 0
transform -1 0 850 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__861_
timestamp 0
transform 1 0 1950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__862_
timestamp 0
transform -1 0 1770 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__863_
timestamp 0
transform -1 0 2850 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__864_
timestamp 0
transform -1 0 2730 0 1 790
box -6 -8 26 268
use FILL  FILL_2__865_
timestamp 0
transform -1 0 2030 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__866_
timestamp 0
transform -1 0 1630 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__867_
timestamp 0
transform 1 0 1050 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__868_
timestamp 0
transform 1 0 830 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__869_
timestamp 0
transform -1 0 470 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__870_
timestamp 0
transform -1 0 650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__871_
timestamp 0
transform -1 0 910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__872_
timestamp 0
transform 1 0 550 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__873_
timestamp 0
transform -1 0 650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__874_
timestamp 0
transform -1 0 790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__875_
timestamp 0
transform 1 0 350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__876_
timestamp 0
transform 1 0 470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__877_
timestamp 0
transform -1 0 70 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__878_
timestamp 0
transform -1 0 350 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__879_
timestamp 0
transform -1 0 510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__880_
timestamp 0
transform -1 0 430 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__881_
timestamp 0
transform -1 0 630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__882_
timestamp 0
transform 1 0 1590 0 1 790
box -6 -8 26 268
use FILL  FILL_2__883_
timestamp 0
transform 1 0 1190 0 1 790
box -6 -8 26 268
use FILL  FILL_2__884_
timestamp 0
transform 1 0 1390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__885_
timestamp 0
transform -1 0 1010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__886_
timestamp 0
transform 1 0 1310 0 1 790
box -6 -8 26 268
use FILL  FILL_2__887_
timestamp 0
transform -1 0 870 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__888_
timestamp 0
transform -1 0 910 0 1 790
box -6 -8 26 268
use FILL  FILL_2__889_
timestamp 0
transform -1 0 2350 0 1 790
box -6 -8 26 268
use FILL  FILL_2__890_
timestamp 0
transform 1 0 950 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__891_
timestamp 0
transform 1 0 750 0 1 790
box -6 -8 26 268
use FILL  FILL_2__892_
timestamp 0
transform -1 0 630 0 1 790
box -6 -8 26 268
use FILL  FILL_2__893_
timestamp 0
transform -1 0 770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__894_
timestamp 0
transform -1 0 1050 0 1 790
box -6 -8 26 268
use FILL  FILL_2__895_
timestamp 0
transform -1 0 730 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__896_
timestamp 0
transform -1 0 450 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__897_
timestamp 0
transform 1 0 2710 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__898_
timestamp 0
transform 1 0 2190 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__899_
timestamp 0
transform 1 0 4250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__900_
timestamp 0
transform -1 0 2310 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__901_
timestamp 0
transform 1 0 2190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__902_
timestamp 0
transform -1 0 2170 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__903_
timestamp 0
transform 1 0 330 0 1 790
box -6 -8 26 268
use FILL  FILL_2__904_
timestamp 0
transform -1 0 590 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__905_
timestamp 0
transform -1 0 490 0 1 790
box -6 -8 26 268
use FILL  FILL_2__906_
timestamp 0
transform 1 0 50 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__907_
timestamp 0
transform 1 0 190 0 1 790
box -6 -8 26 268
use FILL  FILL_2__908_
timestamp 0
transform -1 0 370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__909_
timestamp 0
transform 1 0 370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__910_
timestamp 0
transform -1 0 250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__911_
timestamp 0
transform -1 0 70 0 1 790
box -6 -8 26 268
use FILL  FILL_2__912_
timestamp 0
transform -1 0 330 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__913_
timestamp 0
transform 1 0 170 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__914_
timestamp 0
transform 1 0 50 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__915_
timestamp 0
transform 1 0 190 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__916_
timestamp 0
transform 1 0 210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__917_
timestamp 0
transform 1 0 50 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__918_
timestamp 0
transform 1 0 2850 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__919_
timestamp 0
transform 1 0 770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__920_
timestamp 0
transform 1 0 170 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__921_
timestamp 0
transform 1 0 150 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__922_
timestamp 0
transform 1 0 2430 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__923_
timestamp 0
transform 1 0 2050 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__924_
timestamp 0
transform 1 0 2190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__925_
timestamp 0
transform 1 0 3890 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__926_
timestamp 0
transform -1 0 2730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__927_
timestamp 0
transform 1 0 2570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__928_
timestamp 0
transform -1 0 2490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__929_
timestamp 0
transform 1 0 2350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__930_
timestamp 0
transform -1 0 2590 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__931_
timestamp 0
transform -1 0 2430 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__932_
timestamp 0
transform -1 0 2170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__933_
timestamp 0
transform 1 0 1070 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__934_
timestamp 0
transform 1 0 1110 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__935_
timestamp 0
transform 1 0 1550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__936_
timestamp 0
transform -1 0 2010 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__937_
timestamp 0
transform -1 0 2230 0 1 790
box -6 -8 26 268
use FILL  FILL_2__938_
timestamp 0
transform -1 0 1470 0 1 790
box -6 -8 26 268
use FILL  FILL_2__939_
timestamp 0
transform -1 0 1410 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__940_
timestamp 0
transform -1 0 1750 0 1 790
box -6 -8 26 268
use FILL  FILL_2__941_
timestamp 0
transform -1 0 2830 0 1 790
box -6 -8 26 268
use FILL  FILL_2__942_
timestamp 0
transform 1 0 1830 0 1 790
box -6 -8 26 268
use FILL  FILL_2__943_
timestamp 0
transform -1 0 2470 0 1 790
box -6 -8 26 268
use FILL  FILL_2__944_
timestamp 0
transform -1 0 1570 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__945_
timestamp 0
transform -1 0 1230 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__946_
timestamp 0
transform -1 0 1710 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__947_
timestamp 0
transform -1 0 1250 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__948_
timestamp 0
transform -1 0 1090 0 1 270
box -6 -8 26 268
use FILL  FILL_2__949_
timestamp 0
transform -1 0 990 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__950_
timestamp 0
transform -1 0 2030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__951_
timestamp 0
transform 1 0 1350 0 1 270
box -6 -8 26 268
use FILL  FILL_2__952_
timestamp 0
transform -1 0 1230 0 1 270
box -6 -8 26 268
use FILL  FILL_2__953_
timestamp 0
transform -1 0 810 0 1 270
box -6 -8 26 268
use FILL  FILL_2__954_
timestamp 0
transform -1 0 370 0 1 270
box -6 -8 26 268
use FILL  FILL_2__955_
timestamp 0
transform -1 0 310 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__956_
timestamp 0
transform -1 0 950 0 1 270
box -6 -8 26 268
use FILL  FILL_2__957_
timestamp 0
transform -1 0 850 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__958_
timestamp 0
transform -1 0 670 0 1 270
box -6 -8 26 268
use FILL  FILL_2__959_
timestamp 0
transform -1 0 230 0 1 270
box -6 -8 26 268
use FILL  FILL_2__960_
timestamp 0
transform -1 0 430 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__961_
timestamp 0
transform -1 0 530 0 1 270
box -6 -8 26 268
use FILL  FILL_2__962_
timestamp 0
transform -1 0 70 0 1 270
box -6 -8 26 268
use FILL  FILL_2__963_
timestamp 0
transform -1 0 70 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__964_
timestamp 0
transform 1 0 50 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__965_
timestamp 0
transform 1 0 50 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__966_
timestamp 0
transform -1 0 870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__967_
timestamp 0
transform -1 0 990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__968_
timestamp 0
transform 1 0 1110 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__969_
timestamp 0
transform 1 0 170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__970_
timestamp 0
transform 1 0 550 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__971_
timestamp 0
transform -1 0 710 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__972_
timestamp 0
transform 1 0 2830 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__973_
timestamp 0
transform 1 0 2270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__974_
timestamp 0
transform 1 0 2290 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__975_
timestamp 0
transform 1 0 1770 0 1 270
box -6 -8 26 268
use FILL  FILL_2__976_
timestamp 0
transform 1 0 1870 0 1 270
box -6 -8 26 268
use FILL  FILL_2__977_
timestamp 0
transform 1 0 2950 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__978_
timestamp 0
transform -1 0 3390 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__979_
timestamp 0
transform 1 0 3230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__980_
timestamp 0
transform -1 0 3510 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__981_
timestamp 0
transform -1 0 3530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__982_
timestamp 0
transform -1 0 3110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__983_
timestamp 0
transform -1 0 3010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__984_
timestamp 0
transform -1 0 3370 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__985_
timestamp 0
transform -1 0 2970 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__986_
timestamp 0
transform 1 0 3090 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__987_
timestamp 0
transform -1 0 2910 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__988_
timestamp 0
transform -1 0 2110 0 1 790
box -6 -8 26 268
use FILL  FILL_2__989_
timestamp 0
transform 1 0 1950 0 1 790
box -6 -8 26 268
use FILL  FILL_2__990_
timestamp 0
transform 1 0 3770 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__991_
timestamp 0
transform -1 0 3170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__992_
timestamp 0
transform -1 0 3450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__993_
timestamp 0
transform -1 0 3770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__994_
timestamp 0
transform -1 0 3830 0 1 790
box -6 -8 26 268
use FILL  FILL_2__995_
timestamp 0
transform -1 0 3550 0 1 790
box -6 -8 26 268
use FILL  FILL_2__996_
timestamp 0
transform -1 0 3410 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__997_
timestamp 0
transform -1 0 3770 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__998_
timestamp 0
transform 1 0 3650 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__999_
timestamp 0
transform -1 0 3290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1000_
timestamp 0
transform -1 0 3270 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1001_
timestamp 0
transform -1 0 2690 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1002_
timestamp 0
transform -1 0 2150 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1003_
timestamp 0
transform 1 0 1830 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1004_
timestamp 0
transform 1 0 3230 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1005_
timestamp 0
transform -1 0 3410 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1006_
timestamp 0
transform -1 0 2970 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1007_
timestamp 0
transform 1 0 2530 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1008_
timestamp 0
transform 1 0 3010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1009_
timestamp 0
transform 1 0 2950 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1010_
timestamp 0
transform -1 0 3110 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1011_
timestamp 0
transform -1 0 3170 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1012_
timestamp 0
transform -1 0 2610 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1013_
timestamp 0
transform 1 0 1490 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1014_
timestamp 0
transform 1 0 1630 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1015_
timestamp 0
transform -1 0 3030 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1016_
timestamp 0
transform -1 0 2410 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1017_
timestamp 0
transform -1 0 2330 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1018_
timestamp 0
transform -1 0 2030 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1019_
timestamp 0
transform -1 0 2750 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1020_
timestamp 0
transform 1 0 2450 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1021_
timestamp 0
transform -1 0 2510 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1022_
timestamp 0
transform 1 0 1810 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1023_
timestamp 0
transform -1 0 1490 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1024_
timestamp 0
transform 1 0 1350 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1025_
timestamp 0
transform 1 0 1930 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1026_
timestamp 0
transform 1 0 50 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1027_
timestamp 0
transform 1 0 270 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1028_
timestamp 0
transform -1 0 2370 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1029_
timestamp 0
transform 1 0 2170 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1030_
timestamp 0
transform -1 0 2230 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1031_
timestamp 0
transform -1 0 2090 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1032_
timestamp 0
transform 1 0 1370 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1033_
timestamp 0
transform 1 0 1210 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1034_
timestamp 0
transform 1 0 1650 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1035_
timestamp 0
transform -1 0 2790 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1036_
timestamp 0
transform 1 0 2630 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1037_
timestamp 0
transform -1 0 3250 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1038_
timestamp 0
transform 1 0 3810 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1039_
timestamp 0
transform 1 0 3310 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1040_
timestamp 0
transform 1 0 3410 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1041_
timestamp 0
transform 1 0 4010 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1042_
timestamp 0
transform 1 0 3750 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1043_
timestamp 0
transform -1 0 4330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1044_
timestamp 0
transform 1 0 3470 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1045_
timestamp 0
transform 1 0 3610 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1046_
timestamp 0
transform 1 0 4170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1047_
timestamp 0
transform -1 0 4090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1048_
timestamp 0
transform 1 0 3890 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1049_
timestamp 0
transform -1 0 3670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1050_
timestamp 0
transform -1 0 3810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1051_
timestamp 0
transform -1 0 3950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1052_
timestamp 0
transform -1 0 4810 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1053_
timestamp 0
transform -1 0 3510 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1054_
timestamp 0
transform 1 0 3950 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1055_
timestamp 0
transform 1 0 4810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1056_
timestamp 0
transform 1 0 4930 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1057_
timestamp 0
transform -1 0 4430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1058_
timestamp 0
transform -1 0 4470 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1059_
timestamp 0
transform 1 0 4070 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1060_
timestamp 0
transform -1 0 4170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1061_
timestamp 0
transform -1 0 4310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1062_
timestamp 0
transform 1 0 4590 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1063_
timestamp 0
transform 1 0 4310 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1064_
timestamp 0
transform 1 0 4350 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1065_
timestamp 0
transform -1 0 3610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1066_
timestamp 0
transform -1 0 3690 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1067_
timestamp 0
transform -1 0 4190 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1068_
timestamp 0
transform 1 0 3990 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1069_
timestamp 0
transform 1 0 3870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1070_
timestamp 0
transform 1 0 4010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1071_
timestamp 0
transform -1 0 4030 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1072_
timestamp 0
transform -1 0 4530 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1073_
timestamp 0
transform 1 0 4810 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1074_
timestamp 0
transform 1 0 4450 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1075_
timestamp 0
transform 1 0 4170 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1076_
timestamp 0
transform -1 0 4970 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1077_
timestamp 0
transform -1 0 4270 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1078_
timestamp 0
transform 1 0 2810 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1079_
timestamp 0
transform 1 0 3090 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1080_
timestamp 0
transform -1 0 4690 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1081_
timestamp 0
transform 1 0 4650 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1082_
timestamp 0
transform -1 0 4410 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1083_
timestamp 0
transform -1 0 3990 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1084_
timestamp 0
transform -1 0 4230 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1085_
timestamp 0
transform -1 0 4550 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1086_
timestamp 0
transform -1 0 3850 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1087_
timestamp 0
transform -1 0 3690 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1088_
timestamp 0
transform -1 0 2890 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1089_
timestamp 0
transform 1 0 2870 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1090_
timestamp 0
transform -1 0 3690 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1091_
timestamp 0
transform -1 0 4130 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1092_
timestamp 0
transform -1 0 3550 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1093_
timestamp 0
transform 1 0 3410 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1094_
timestamp 0
transform 1 0 1810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1095_
timestamp 0
transform 1 0 2170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1096_
timestamp 0
transform 1 0 2030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1097_
timestamp 0
transform 1 0 3790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1098_
timestamp 0
transform -1 0 3170 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1099_
timestamp 0
transform -1 0 3570 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1100_
timestamp 0
transform 1 0 3430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1101_
timestamp 0
transform -1 0 4090 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1102_
timestamp 0
transform 1 0 3910 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1103_
timestamp 0
transform 1 0 3890 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1104_
timestamp 0
transform -1 0 5750 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1105_
timestamp 0
transform -1 0 5250 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1106_
timestamp 0
transform 1 0 5090 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1107_
timestamp 0
transform 1 0 4270 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1108_
timestamp 0
transform -1 0 4470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1109_
timestamp 0
transform 1 0 5250 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1110_
timestamp 0
transform 1 0 5090 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1111_
timestamp 0
transform 1 0 5410 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1112_
timestamp 0
transform -1 0 5690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1113_
timestamp 0
transform 1 0 4690 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1114_
timestamp 0
transform 1 0 4510 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1115_
timestamp 0
transform 1 0 4570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1116_
timestamp 0
transform 1 0 4390 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1117_
timestamp 0
transform 1 0 4230 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1118_
timestamp 0
transform 1 0 4630 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1119_
timestamp 0
transform -1 0 5390 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1120_
timestamp 0
transform 1 0 4570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1121_
timestamp 0
transform -1 0 4790 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1122_
timestamp 0
transform -1 0 5230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1123_
timestamp 0
transform 1 0 5630 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1124_
timestamp 0
transform -1 0 5490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1125_
timestamp 0
transform 1 0 5070 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1126_
timestamp 0
transform -1 0 5270 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1127_
timestamp 0
transform 1 0 5430 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1128_
timestamp 0
transform -1 0 5610 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1129_
timestamp 0
transform -1 0 4330 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1130_
timestamp 0
transform 1 0 5170 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1131_
timestamp 0
transform -1 0 5310 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1132_
timestamp 0
transform -1 0 4850 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1133_
timestamp 0
transform 1 0 4970 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1134_
timestamp 0
transform 1 0 5110 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1135_
timestamp 0
transform 1 0 5150 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1136_
timestamp 0
transform -1 0 5470 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1137_
timestamp 0
transform -1 0 5590 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1138_
timestamp 0
transform -1 0 5030 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1139_
timestamp 0
transform 1 0 4870 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1140_
timestamp 0
transform 1 0 5010 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1141_
timestamp 0
transform 1 0 4910 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1142_
timestamp 0
transform -1 0 4750 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1143_
timestamp 0
transform -1 0 5330 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1144_
timestamp 0
transform -1 0 4610 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1145_
timestamp 0
transform -1 0 4290 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1146_
timestamp 0
transform 1 0 4210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1147_
timestamp 0
transform -1 0 3810 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1148_
timestamp 0
transform 1 0 4030 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1149_
timestamp 0
transform -1 0 4150 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1150_
timestamp 0
transform 1 0 5550 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1151_
timestamp 0
transform 1 0 5650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1152_
timestamp 0
transform -1 0 5350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1153_
timestamp 0
transform 1 0 4370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1154_
timestamp 0
transform 1 0 4150 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1155_
timestamp 0
transform 1 0 4490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1156_
timestamp 0
transform 1 0 4630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1157_
timestamp 0
transform 1 0 4230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1158_
timestamp 0
transform 1 0 4770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1159_
timestamp 0
transform -1 0 5230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1160_
timestamp 0
transform -1 0 4470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1161_
timestamp 0
transform -1 0 4930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1162_
timestamp 0
transform 1 0 4370 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1163_
timestamp 0
transform -1 0 4550 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1164_
timestamp 0
transform 1 0 4810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1165_
timestamp 0
transform 1 0 4690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1166_
timestamp 0
transform 1 0 4790 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1167_
timestamp 0
transform 1 0 5330 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1168_
timestamp 0
transform -1 0 5510 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1169_
timestamp 0
transform 1 0 4650 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1170_
timestamp 0
transform 1 0 4930 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1171_
timestamp 0
transform 1 0 5190 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1172_
timestamp 0
transform -1 0 5490 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1173_
timestamp 0
transform 1 0 5370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1174_
timestamp 0
transform 1 0 5050 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1175_
timestamp 0
transform -1 0 5530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1176_
timestamp 0
transform 1 0 5110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1177_
timestamp 0
transform -1 0 4970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1178_
timestamp 0
transform -1 0 5610 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1179_
timestamp 0
transform -1 0 5470 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1180_
timestamp 0
transform -1 0 5250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1181_
timestamp 0
transform -1 0 4530 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1182_
timestamp 0
transform -1 0 4050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1183_
timestamp 0
transform -1 0 3990 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1184_
timestamp 0
transform 1 0 3890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1185_
timestamp 0
transform -1 0 4990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1186_
timestamp 0
transform 1 0 4650 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1187_
timestamp 0
transform -1 0 4410 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1188_
timestamp 0
transform -1 0 4910 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1189_
timestamp 0
transform 1 0 4770 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1190_
timestamp 0
transform -1 0 4550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1191_
timestamp 0
transform 1 0 4390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1192_
timestamp 0
transform 1 0 5630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1193_
timestamp 0
transform -1 0 5070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1194_
timestamp 0
transform 1 0 5470 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1195_
timestamp 0
transform 1 0 4950 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1196_
timestamp 0
transform -1 0 4630 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1197_
timestamp 0
transform 1 0 4350 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1198_
timestamp 0
transform 1 0 4730 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1199_
timestamp 0
transform -1 0 4870 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1200_
timestamp 0
transform 1 0 5270 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1201_
timestamp 0
transform 1 0 5470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1202_
timestamp 0
transform 1 0 5330 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1203_
timestamp 0
transform -1 0 5730 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1204_
timestamp 0
transform -1 0 5590 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1205_
timestamp 0
transform -1 0 5730 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1206_
timestamp 0
transform 1 0 5710 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1207_
timestamp 0
transform -1 0 5630 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1208_
timestamp 0
transform 1 0 5690 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1209_
timestamp 0
transform -1 0 5570 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1210_
timestamp 0
transform -1 0 5450 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1211_
timestamp 0
transform -1 0 5190 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1212_
timestamp 0
transform -1 0 3290 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1213_
timestamp 0
transform 1 0 3010 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1214_
timestamp 0
transform -1 0 3910 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1215_
timestamp 0
transform 1 0 3730 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1216_
timestamp 0
transform -1 0 4950 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1217_
timestamp 0
transform 1 0 4790 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1218_
timestamp 0
transform -1 0 5050 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1219_
timestamp 0
transform 1 0 4950 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1220_
timestamp 0
transform -1 0 5110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1221_
timestamp 0
transform -1 0 5690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1222_
timestamp 0
transform 1 0 5170 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1223_
timestamp 0
transform 1 0 4990 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1224_
timestamp 0
transform 1 0 4710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1225_
timestamp 0
transform 1 0 4490 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1226_
timestamp 0
transform 1 0 4850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1227_
timestamp 0
transform 1 0 5090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1228_
timestamp 0
transform 1 0 5230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1229_
timestamp 0
transform -1 0 5510 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1230_
timestamp 0
transform 1 0 5550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1231_
timestamp 0
transform 1 0 5730 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1232_
timestamp 0
transform -1 0 5750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1233_
timestamp 0
transform 1 0 5550 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1234_
timestamp 0
transform -1 0 5710 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1235_
timestamp 0
transform 1 0 5670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1236_
timestamp 0
transform 1 0 5210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1237_
timestamp 0
transform 1 0 5750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1238_
timestamp 0
transform -1 0 5430 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1239_
timestamp 0
transform -1 0 5290 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1240_
timestamp 0
transform -1 0 5350 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1241_
timestamp 0
transform -1 0 5310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1242_
timestamp 0
transform -1 0 5170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1243_
timestamp 0
transform 1 0 5370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1244_
timestamp 0
transform 1 0 4570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1245_
timestamp 0
transform 1 0 4950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1246_
timestamp 0
transform 1 0 5150 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1247_
timestamp 0
transform -1 0 5030 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1248_
timestamp 0
transform 1 0 5010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1249_
timestamp 0
transform -1 0 5430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1250_
timestamp 0
transform -1 0 4650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1251_
timestamp 0
transform 1 0 4870 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1252_
timestamp 0
transform 1 0 4730 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1253_
timestamp 0
transform -1 0 5450 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1254_
timestamp 0
transform -1 0 5310 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1255_
timestamp 0
transform -1 0 5350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1256_
timestamp 0
transform -1 0 5210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1257_
timestamp 0
transform 1 0 5270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1258_
timestamp 0
transform 1 0 5130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1259_
timestamp 0
transform 1 0 5090 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1260_
timestamp 0
transform -1 0 190 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1261_
timestamp 0
transform 1 0 50 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1262_
timestamp 0
transform 1 0 290 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1263_
timestamp 0
transform -1 0 430 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1264_
timestamp 0
transform -1 0 1050 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1265_
timestamp 0
transform 1 0 530 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1266_
timestamp 0
transform -1 0 830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1267_
timestamp 0
transform 1 0 550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1268_
timestamp 0
transform 1 0 330 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1269_
timestamp 0
transform -1 0 190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1270_
timestamp 0
transform 1 0 50 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1271_
timestamp 0
transform 1 0 290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1272_
timestamp 0
transform 1 0 430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1273_
timestamp 0
transform 1 0 850 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1274_
timestamp 0
transform 1 0 470 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1275_
timestamp 0
transform -1 0 690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1276_
timestamp 0
transform -1 0 1850 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1277_
timestamp 0
transform 1 0 1630 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1278_
timestamp 0
transform 1 0 2050 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1279_
timestamp 0
transform 1 0 1750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1280_
timestamp 0
transform -1 0 1970 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1281_
timestamp 0
transform 1 0 1810 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1282_
timestamp 0
transform 1 0 290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1283_
timestamp 0
transform -1 0 530 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1284_
timestamp 0
transform 1 0 690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1285_
timestamp 0
transform -1 0 830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1286_
timestamp 0
transform -1 0 1510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1287_
timestamp 0
transform 1 0 1350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1288_
timestamp 0
transform -1 0 230 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1289_
timestamp 0
transform -1 0 70 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1290_
timestamp 0
transform 1 0 50 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1291_
timestamp 0
transform 1 0 50 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1292_
timestamp 0
transform 1 0 330 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1293_
timestamp 0
transform -1 0 610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1294_
timestamp 0
transform 1 0 450 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1295_
timestamp 0
transform -1 0 190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1296_
timestamp 0
transform -1 0 70 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1297_
timestamp 0
transform 1 0 210 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1298_
timestamp 0
transform -1 0 290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1299_
timestamp 0
transform 1 0 50 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1300_
timestamp 0
transform -1 0 690 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1301_
timestamp 0
transform 1 0 170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1302_
timestamp 0
transform -1 0 710 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1303_
timestamp 0
transform -1 0 850 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1304_
timestamp 0
transform 1 0 550 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1305_
timestamp 0
transform -1 0 410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1306_
timestamp 0
transform 1 0 310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1307_
timestamp 0
transform -1 0 670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1308_
timestamp 0
transform -1 0 590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1309_
timestamp 0
transform -1 0 530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1310_
timestamp 0
transform -1 0 1530 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1311_
timestamp 0
transform 1 0 710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1312_
timestamp 0
transform 1 0 870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1313_
timestamp 0
transform -1 0 1010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1314_
timestamp 0
transform -1 0 930 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1315_
timestamp 0
transform 1 0 1050 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1316_
timestamp 0
transform 1 0 1270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1317_
timestamp 0
transform -1 0 1190 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1318_
timestamp 0
transform 1 0 1670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1319_
timestamp 0
transform -1 0 1570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1320_
timestamp 0
transform 1 0 1310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1321_
timestamp 0
transform -1 0 1430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1322_
timestamp 0
transform 1 0 1650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1323_
timestamp 0
transform 1 0 2310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1324_
timestamp 0
transform 1 0 2170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1325_
timestamp 0
transform -1 0 1710 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1326_
timestamp 0
transform 1 0 430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1327_
timestamp 0
transform -1 0 1070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1328_
timestamp 0
transform 1 0 1170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1329_
timestamp 0
transform -1 0 1130 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1330_
timestamp 0
transform 1 0 1010 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1331_
timestamp 0
transform -1 0 450 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1332_
timestamp 0
transform 1 0 870 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1333_
timestamp 0
transform 1 0 1150 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1334_
timestamp 0
transform -1 0 2050 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1335_
timestamp 0
transform 1 0 1750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1336_
timestamp 0
transform -1 0 1890 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1337_
timestamp 0
transform -1 0 1830 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1338_
timestamp 0
transform 1 0 1410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1339_
timestamp 0
transform 1 0 1930 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1340_
timestamp 0
transform -1 0 1530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1341_
timestamp 0
transform -1 0 1570 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1342_
timestamp 0
transform 1 0 1650 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1343_
timestamp 0
transform 1 0 1890 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1344_
timestamp 0
transform -1 0 2030 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1345_
timestamp 0
transform -1 0 1450 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1346_
timestamp 0
transform -1 0 1550 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1347_
timestamp 0
transform 1 0 1650 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1348_
timestamp 0
transform 1 0 1930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1349_
timestamp 0
transform 1 0 3090 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1350_
timestamp 0
transform 1 0 2950 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1351_
timestamp 0
transform 1 0 2390 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1352_
timestamp 0
transform -1 0 1810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1353_
timestamp 0
transform 1 0 1750 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1354_
timestamp 0
transform 1 0 1850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1355_
timestamp 0
transform 1 0 4770 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1356_
timestamp 0
transform 1 0 4850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1357_
timestamp 0
transform -1 0 4670 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1358_
timestamp 0
transform -1 0 4290 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1359_
timestamp 0
transform -1 0 2810 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1360_
timestamp 0
transform -1 0 2670 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1361_
timestamp 0
transform -1 0 2530 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1362_
timestamp 0
transform -1 0 3870 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1363_
timestamp 0
transform -1 0 3990 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1364_
timestamp 0
transform -1 0 5430 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1365_
timestamp 0
transform -1 0 5650 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1366_
timestamp 0
transform 1 0 5530 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1367_
timestamp 0
transform 1 0 5030 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1368_
timestamp 0
transform 1 0 4090 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1369_
timestamp 0
transform -1 0 3410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1370_
timestamp 0
transform -1 0 3770 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1371_
timestamp 0
transform -1 0 3970 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1372_
timestamp 0
transform -1 0 4910 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1373_
timestamp 0
transform -1 0 4390 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1374_
timestamp 0
transform 1 0 4490 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1375_
timestamp 0
transform -1 0 5670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1376_
timestamp 0
transform 1 0 5530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1377_
timestamp 0
transform -1 0 5310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1378_
timestamp 0
transform 1 0 5390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1379_
timestamp 0
transform -1 0 4470 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1380_
timestamp 0
transform 1 0 4570 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1381_
timestamp 0
transform -1 0 4850 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1382_
timestamp 0
transform -1 0 4690 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1383_
timestamp 0
transform -1 0 4330 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1384_
timestamp 0
transform 1 0 5150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1385_
timestamp 0
transform 1 0 5290 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1386_
timestamp 0
transform 1 0 5070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1387_
timestamp 0
transform -1 0 5190 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1388_
timestamp 0
transform -1 0 4950 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1389_
timestamp 0
transform 1 0 4990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1390_
timestamp 0
transform -1 0 4870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1391_
timestamp 0
transform 1 0 4690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1392_
timestamp 0
transform -1 0 5050 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1393_
timestamp 0
transform -1 0 4490 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1394_
timestamp 0
transform -1 0 4730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1395_
timestamp 0
transform -1 0 4350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1396_
timestamp 0
transform 1 0 3110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1397_
timestamp 0
transform -1 0 3230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1398_
timestamp 0
transform -1 0 2990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1399_
timestamp 0
transform 1 0 2810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1400_
timestamp 0
transform 1 0 3330 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1401_
timestamp 0
transform 1 0 3350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1402_
timestamp 0
transform -1 0 3630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1403_
timestamp 0
transform -1 0 3510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1404_
timestamp 0
transform -1 0 3470 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1405_
timestamp 0
transform -1 0 4610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1406_
timestamp 0
transform 1 0 3070 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1407_
timestamp 0
transform -1 0 4790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1408_
timestamp 0
transform 1 0 4630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1409_
timestamp 0
transform -1 0 4510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1410_
timestamp 0
transform -1 0 4050 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1411_
timestamp 0
transform 1 0 3890 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1412_
timestamp 0
transform 1 0 3430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1413_
timestamp 0
transform 1 0 3350 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1414_
timestamp 0
transform 1 0 3210 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1415_
timestamp 0
transform 1 0 3230 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1416_
timestamp 0
transform 1 0 4550 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1417_
timestamp 0
transform 1 0 4050 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1418_
timestamp 0
transform -1 0 2470 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1419_
timestamp 0
transform 1 0 2530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1420_
timestamp 0
transform -1 0 2670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1421_
timestamp 0
transform -1 0 2450 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1422_
timestamp 0
transform 1 0 2550 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1423_
timestamp 0
transform -1 0 3650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1424_
timestamp 0
transform 1 0 3250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1425_
timestamp 0
transform -1 0 3870 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1426_
timestamp 0
transform 1 0 3710 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1427_
timestamp 0
transform -1 0 2910 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1428_
timestamp 0
transform -1 0 3430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1429_
timestamp 0
transform 1 0 3270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1430_
timestamp 0
transform -1 0 2770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1431_
timestamp 0
transform -1 0 2910 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1432_
timestamp 0
transform -1 0 2630 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1433_
timestamp 0
transform -1 0 2770 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1434_
timestamp 0
transform -1 0 3030 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1435_
timestamp 0
transform -1 0 3170 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1436_
timestamp 0
transform 1 0 3170 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1437_
timestamp 0
transform -1 0 3550 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1438_
timestamp 0
transform -1 0 1170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1439_
timestamp 0
transform -1 0 1290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1440_
timestamp 0
transform -1 0 3810 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1441_
timestamp 0
transform -1 0 3930 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1442_
timestamp 0
transform -1 0 3330 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1443_
timestamp 0
transform 1 0 3450 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1444_
timestamp 0
transform 1 0 2670 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1445_
timestamp 0
transform -1 0 2550 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1446_
timestamp 0
transform 1 0 2490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1447_
timestamp 0
transform 1 0 2350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1448_
timestamp 0
transform 1 0 3710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1449_
timestamp 0
transform 1 0 3090 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1450_
timestamp 0
transform 1 0 3550 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1451_
timestamp 0
transform -1 0 3590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1527_
timestamp 0
transform -1 0 70 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1528_
timestamp 0
transform 1 0 2410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1529_
timestamp 0
transform -1 0 2550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1530_
timestamp 0
transform 1 0 5730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1531_
timestamp 0
transform 1 0 5610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1532_
timestamp 0
transform -1 0 2050 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1533_
timestamp 0
transform 1 0 2810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1534_
timestamp 0
transform 1 0 2170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1535_
timestamp 0
transform -1 0 2850 0 1 4950
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert0
timestamp 0
transform 1 0 790 0 1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert1
timestamp 0
transform 1 0 4510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert2
timestamp 0
transform 1 0 2330 0 1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert3
timestamp 0
transform -1 0 1630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert4
timestamp 0
transform -1 0 770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert5
timestamp 0
transform 1 0 4670 0 1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert6
timestamp 0
transform 1 0 3470 0 1 3910
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert15
timestamp 0
transform 1 0 2770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert16
timestamp 0
transform 1 0 1830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert17
timestamp 0
transform -1 0 2610 0 1 790
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert18
timestamp 0
transform -1 0 2050 0 1 1830
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert19
timestamp 0
transform 1 0 2430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert20
timestamp 0
transform -1 0 1510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert21
timestamp 0
transform 1 0 3270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert22
timestamp 0
transform -1 0 1330 0 1 4430
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert23
timestamp 0
transform -1 0 2970 0 1 4430
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert24
timestamp 0
transform 1 0 3590 0 1 3910
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert25
timestamp 0
transform -1 0 3650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert26
timestamp 0
transform -1 0 3610 0 1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert27
timestamp 0
transform -1 0 3290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert28
timestamp 0
transform -1 0 2930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert29
timestamp 0
transform -1 0 2030 0 1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert30
timestamp 0
transform -1 0 1910 0 1 1310
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert31
timestamp 0
transform 1 0 3630 0 1 1310
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert32
timestamp 0
transform 1 0 2650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert33
timestamp 0
transform -1 0 1690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert7
timestamp 0
transform -1 0 1290 0 1 3390
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert8
timestamp 0
transform -1 0 1630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert9
timestamp 0
transform 1 0 4090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert10
timestamp 0
transform -1 0 3570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert11
timestamp 0
transform -1 0 910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert12
timestamp 0
transform 1 0 3550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert13
timestamp 0
transform 1 0 4270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert14
timestamp 0
transform 1 0 2270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__727_
timestamp 0
transform 1 0 3070 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__735_
timestamp 0
transform -1 0 1170 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__742_
timestamp 0
transform 1 0 2770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__750_
timestamp 0
transform 1 0 2710 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__757_
timestamp 0
transform -1 0 3990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__765_
timestamp 0
transform -1 0 3850 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__772_
timestamp 0
transform 1 0 2090 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__780_
timestamp 0
transform 1 0 190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__788_
timestamp 0
transform 1 0 2790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__795_
timestamp 0
transform -1 0 2370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__803_
timestamp 0
transform -1 0 5570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__810_
timestamp 0
transform 1 0 3090 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__818_
timestamp 0
transform 1 0 1590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__825_
timestamp 0
transform 1 0 1350 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__833_
timestamp 0
transform 1 0 1850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__841_
timestamp 0
transform -1 0 1050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__848_
timestamp 0
transform -1 0 1510 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__856_
timestamp 0
transform 1 0 510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__863_
timestamp 0
transform -1 0 2870 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__871_
timestamp 0
transform -1 0 930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__878_
timestamp 0
transform -1 0 370 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__886_
timestamp 0
transform 1 0 1330 0 1 790
box -6 -8 26 268
use FILL  FILL_3__894_
timestamp 0
transform -1 0 1070 0 1 790
box -6 -8 26 268
use FILL  FILL_3__901_
timestamp 0
transform 1 0 2210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__909_
timestamp 0
transform 1 0 390 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__916_
timestamp 0
transform 1 0 230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__924_
timestamp 0
transform 1 0 2210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__931_
timestamp 0
transform -1 0 2450 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__939_
timestamp 0
transform -1 0 1430 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__947_
timestamp 0
transform -1 0 1270 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__954_
timestamp 0
transform -1 0 390 0 1 270
box -6 -8 26 268
use FILL  FILL_3__962_
timestamp 0
transform -1 0 90 0 1 270
box -6 -8 26 268
use FILL  FILL_3__969_
timestamp 0
transform 1 0 190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__977_
timestamp 0
transform 1 0 2970 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__984_
timestamp 0
transform -1 0 3390 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__992_
timestamp 0
transform -1 0 3470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__999_
timestamp 0
transform -1 0 3310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1003_
timestamp 0
transform 1 0 1850 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1011_
timestamp 0
transform -1 0 3190 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1018_
timestamp 0
transform -1 0 2050 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1026_
timestamp 0
transform 1 0 70 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1034_
timestamp 0
transform 1 0 1670 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1041_
timestamp 0
transform 1 0 4030 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1049_
timestamp 0
transform -1 0 3690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1056_
timestamp 0
transform 1 0 4950 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1064_
timestamp 0
transform 1 0 4370 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1071_
timestamp 0
transform -1 0 4050 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1079_
timestamp 0
transform 1 0 3110 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1087_
timestamp 0
transform -1 0 3710 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1094_
timestamp 0
transform 1 0 1830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1102_
timestamp 0
transform 1 0 3930 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1109_
timestamp 0
transform 1 0 5270 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1117_
timestamp 0
transform 1 0 4250 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1124_
timestamp 0
transform -1 0 5510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1132_
timestamp 0
transform -1 0 4870 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1140_
timestamp 0
transform 1 0 5030 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1147_
timestamp 0
transform -1 0 3830 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1155_
timestamp 0
transform 1 0 4510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1162_
timestamp 0
transform 1 0 4390 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1170_
timestamp 0
transform 1 0 4950 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1177_
timestamp 0
transform -1 0 4990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1185_
timestamp 0
transform -1 0 5010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1193_
timestamp 0
transform -1 0 5090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1200_
timestamp 0
transform 1 0 5290 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1208_
timestamp 0
transform 1 0 5710 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1215_
timestamp 0
transform 1 0 3750 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1223_
timestamp 0
transform 1 0 5010 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1230_
timestamp 0
transform 1 0 5570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1238_
timestamp 0
transform -1 0 5450 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1246_
timestamp 0
transform 1 0 5170 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1253_
timestamp 0
transform -1 0 5470 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1261_
timestamp 0
transform 1 0 70 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1268_
timestamp 0
transform 1 0 350 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1276_
timestamp 0
transform -1 0 1870 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1283_
timestamp 0
transform -1 0 550 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1291_
timestamp 0
transform 1 0 70 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1299_
timestamp 0
transform 1 0 70 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1306_
timestamp 0
transform 1 0 330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1314_
timestamp 0
transform -1 0 950 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1321_
timestamp 0
transform -1 0 1450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1329_
timestamp 0
transform -1 0 1150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1336_
timestamp 0
transform -1 0 1910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1344_
timestamp 0
transform -1 0 2050 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1352_
timestamp 0
transform -1 0 1830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1359_
timestamp 0
transform -1 0 2830 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1367_
timestamp 0
transform 1 0 5050 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1374_
timestamp 0
transform 1 0 4510 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1382_
timestamp 0
transform -1 0 4710 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1389_
timestamp 0
transform 1 0 5010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1397_
timestamp 0
transform -1 0 3250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1404_
timestamp 0
transform -1 0 3490 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1412_
timestamp 0
transform 1 0 3450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1420_
timestamp 0
transform -1 0 2690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1427_
timestamp 0
transform -1 0 2930 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1435_
timestamp 0
transform -1 0 3190 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1442_
timestamp 0
transform -1 0 3350 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1450_
timestamp 0
transform 1 0 3570 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1532_
timestamp 0
transform -1 0 2070 0 1 4950
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert3
timestamp 0
transform -1 0 1650 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert18
timestamp 0
transform -1 0 2070 0 1 1830
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert26
timestamp 0
transform -1 0 3630 0 1 2870
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert33
timestamp 0
transform -1 0 1710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert11
timestamp 0
transform -1 0 930 0 -1 5470
box -6 -8 26 268
<< labels >>
flabel metal1 s 5843 2 5903 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -63 2 -3 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal3 s 5876 1956 5884 1964 3 FreeSans 16 0 0 0 Cin[5]
port 2 nsew
flabel metal3 s 5876 1436 5884 1444 3 FreeSans 16 0 0 0 Cin[4]
port 3 nsew
flabel metal3 s 5876 2296 5884 2304 3 FreeSans 16 0 0 0 Cin[3]
port 4 nsew
flabel metal2 s 3837 -23 3843 -17 7 FreeSans 16 270 0 0 Cin[2]
port 5 nsew
flabel metal2 s 2697 -23 2703 -17 7 FreeSans 16 270 0 0 Cin[1]
port 6 nsew
flabel metal2 s 2657 -23 2663 -17 7 FreeSans 16 270 0 0 Cin[0]
port 7 nsew
flabel metal3 s -24 2736 -16 2744 7 FreeSans 16 0 0 0 Rdy
port 8 nsew
flabel metal3 s -24 2996 -16 3004 7 FreeSans 16 0 0 0 Vld
port 9 nsew
flabel metal3 s 5876 2476 5884 2484 3 FreeSans 16 0 0 0 Xin[3]
port 10 nsew
flabel metal3 s 5876 2736 5884 2744 3 FreeSans 16 0 0 0 Xin[2]
port 11 nsew
flabel metal2 s 2537 -23 2543 -17 7 FreeSans 16 270 0 0 Xin[1]
port 12 nsew
flabel metal2 s 2837 -23 2843 -17 7 FreeSans 16 270 0 0 Xin[0]
port 13 nsew
flabel metal3 s 5876 2256 5884 2264 3 FreeSans 16 0 0 0 Xout[3]
port 14 nsew
flabel metal3 s 5876 2216 5884 2224 3 FreeSans 16 0 0 0 Xout[2]
port 15 nsew
flabel metal2 s 2577 -23 2583 -17 7 FreeSans 16 270 0 0 Xout[1]
port 16 nsew
flabel metal2 s 2457 -23 2463 -17 7 FreeSans 16 270 0 0 Xout[0]
port 17 nsew
flabel metal2 s 3257 5517 3263 5523 3 FreeSans 16 90 0 0 Yin[3]
port 18 nsew
flabel metal2 s 3477 5517 3483 5523 3 FreeSans 16 90 0 0 Yin[2]
port 19 nsew
flabel metal2 s 4517 5517 4523 5523 3 FreeSans 16 90 0 0 Yin[1]
port 20 nsew
flabel metal2 s 4617 5517 4623 5523 3 FreeSans 16 90 0 0 Yin[0]
port 21 nsew
flabel metal2 s 2837 5517 2843 5523 3 FreeSans 16 90 0 0 Yout[3]
port 22 nsew
flabel metal2 s 2217 5517 2223 5523 3 FreeSans 16 90 0 0 Yout[2]
port 23 nsew
flabel metal2 s 2877 5517 2883 5523 3 FreeSans 16 90 0 0 Yout[1]
port 24 nsew
flabel metal2 s 2097 5517 2103 5523 3 FreeSans 16 90 0 0 Yout[0]
port 25 nsew
flabel metal2 s 1037 5517 1043 5523 3 FreeSans 16 90 0 0 clk
port 26 nsew
<< properties >>
string FIXED_BBOX -40 -40 5880 5520
<< end >>
