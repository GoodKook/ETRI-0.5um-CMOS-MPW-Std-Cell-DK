magic
tech scmos
magscale 1 2
timestamp 1702311544
<< nwell >>
rect -13 154 94 272
<< ntransistor >>
rect 18 14 22 54
rect 28 14 32 54
rect 48 14 52 34
<< ptransistor >>
rect 18 206 22 246
rect 38 206 42 246
rect 58 206 62 246
<< ndiffusion >>
rect 16 14 18 54
rect 22 14 28 54
rect 32 14 34 54
rect 46 14 48 34
rect 52 14 54 34
<< pdiffusion >>
rect 16 206 18 246
rect 22 206 24 246
rect 36 206 38 246
rect 42 206 44 246
rect 56 206 58 246
rect 62 206 64 246
<< ndcontact >>
rect 4 14 16 54
rect 34 14 46 54
rect 54 14 66 34
<< pdcontact >>
rect 4 206 16 246
rect 24 206 36 246
rect 44 206 56 246
rect 64 206 76 246
<< psubstratepcontact >>
rect -6 -6 86 6
<< nsubstratencontact >>
rect -6 254 86 266
<< polysilicon >>
rect 18 246 22 250
rect 38 246 42 250
rect 58 246 62 250
rect 18 54 22 206
rect 38 97 42 206
rect 28 85 38 97
rect 28 54 32 85
rect 58 72 62 206
rect 60 60 62 72
rect 48 34 52 60
rect 18 10 22 14
rect 28 10 32 14
rect 48 10 52 14
<< polycontact >>
rect 6 105 18 117
rect 38 85 50 97
rect 48 60 60 72
<< metal1 >>
rect -6 266 86 268
rect -6 252 86 254
rect 4 246 16 252
rect 44 246 56 252
rect 3 123 17 137
rect 6 117 17 123
rect 24 72 30 206
rect 66 137 74 206
rect 63 123 77 137
rect 43 103 57 117
rect 43 97 52 103
rect 50 85 52 97
rect 4 64 48 72
rect 4 54 16 64
rect 66 40 74 123
rect 54 34 74 40
rect 34 8 46 14
rect -6 6 86 8
rect -6 -8 86 -6
<< m1p >>
rect -6 252 86 268
rect 3 123 17 137
rect 63 123 77 137
rect 43 103 57 117
rect -6 -8 86 8
<< labels >>
rlabel nsubstratencontact 40 260 40 260 0 vdd
port 4 nsew power bidirectional abutment
rlabel psubstratepcontact 40 0 40 0 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal1 10 127 10 127 1 A
port 1 n signal input
rlabel metal1 50 107 50 107 5 B
port 2 n signal input
rlabel metal1 70 127 70 127 1 Y
port 3 n signal output
<< properties >>
string FIXED_BBOX 0 0 80 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
