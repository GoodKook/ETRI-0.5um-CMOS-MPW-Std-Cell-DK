magic
tech scmos
magscale 1 3
timestamp 1725338299
<< checkpaint >>
rect -25 299 275 300
rect -29 279 279 299
rect -49 275 299 279
rect -49 -25 300 275
rect -49 -29 299 -25
rect -29 -49 279 -29
rect -25 -50 275 -49
<< ndiffusion >>
rect 75 75 175 175
<< psubstratepdiff >>
rect 10 220 240 240
rect 10 30 30 220
rect 220 30 240 220
rect 10 10 240 30
<< genericcontact >>
rect 35 220 215 240
rect 10 35 30 215
rect 75 75 175 175
rect 220 35 240 215
rect 35 10 215 30
<< metal1 >>
rect 10 220 240 240
rect 10 30 30 220
rect 75 75 175 175
rect 220 30 240 220
rect 10 10 240 30
<< end >>
