magic
tech scmos
magscale 1 2
timestamp 1727495774
<< nwell >>
rect -6 154 126 272
<< ntransistor >>
rect 20 14 24 54
rect 40 14 44 54
rect 60 14 64 54
rect 80 14 84 54
<< ptransistor >>
rect 20 166 24 246
rect 30 166 34 246
rect 60 166 64 246
rect 70 166 74 246
<< ndiffusion >>
rect 18 14 20 54
rect 24 44 40 54
rect 24 14 26 44
rect 38 14 40 44
rect 44 14 46 54
rect 58 14 60 54
rect 64 26 66 54
rect 78 26 80 54
rect 64 14 80 26
rect 84 14 86 54
<< pdiffusion >>
rect 18 166 20 246
rect 24 166 30 246
rect 34 166 36 246
rect 58 166 60 246
rect 64 166 70 246
rect 74 166 76 246
<< ndcontact >>
rect 6 14 18 54
rect 26 14 38 44
rect 46 14 58 54
rect 66 26 78 54
rect 86 14 98 54
<< pdcontact >>
rect 6 166 18 246
rect 36 166 58 246
rect 76 166 88 246
<< psubstratepcontact >>
rect 0 -6 120 6
<< nsubstratencontact >>
rect 0 254 120 266
<< polysilicon >>
rect 20 246 24 250
rect 30 246 34 250
rect 60 246 64 250
rect 70 246 74 250
rect 20 162 24 166
rect 10 158 24 162
rect 30 162 34 166
rect 30 158 44 162
rect 10 129 16 158
rect 40 123 44 158
rect 10 82 16 117
rect 36 111 44 123
rect 10 76 24 82
rect 20 54 24 76
rect 40 54 44 111
rect 60 54 64 166
rect 70 162 74 166
rect 70 158 88 162
rect 84 129 88 158
rect 84 82 88 117
rect 80 76 88 82
rect 80 54 84 76
rect 20 10 24 14
rect 40 10 44 14
rect 60 10 64 14
rect 80 10 84 14
<< polycontact >>
rect 4 117 16 129
rect 24 111 36 123
rect 64 111 76 123
rect 84 117 96 129
<< metal1 >>
rect 0 266 120 268
rect 0 252 120 254
rect 6 246 18 252
rect 76 246 88 252
rect 44 117 52 166
rect 43 72 52 103
rect 43 64 74 72
rect 6 54 58 56
rect 68 54 74 64
rect 18 50 46 54
rect 58 14 86 20
rect 26 8 38 14
rect 0 6 120 8
rect 0 -8 120 -6
<< m2contact >>
rect 23 123 37 137
rect 3 103 17 117
rect 63 123 77 137
rect 43 103 57 117
rect 83 103 97 117
<< metal2 >>
rect 23 137 37 157
rect 63 137 77 157
rect 3 83 17 103
rect 43 83 57 103
rect 83 83 97 103
<< m2p >>
rect 23 143 37 157
rect 63 143 77 157
rect 3 83 17 97
rect 43 83 57 97
rect 83 83 97 97
<< labels >>
rlabel metal2 3 83 17 97 0 A
port 0 nsew signal input
rlabel metal2 23 143 37 157 0 B
port 1 nsew signal input
rlabel metal2 63 143 77 157 0 D
port 3 nsew signal input
rlabel metal2 83 83 97 97 0 C
port 2 nsew signal input
rlabel metal2 43 83 57 97 0 Y
port 4 nsew signal output
rlabel metal1 0 266 120 268 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal1 0 254 120 266 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal1 0 252 120 254 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal1 0 6 120 8 0 gnd
port 6 nsew ground bidirectional abutment
rlabel metal1 0 -6 120 6 0 gnd
port 6 nsew ground bidirectional abutment
rlabel metal1 0 -8 120 -6 0 gnd
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 120 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
