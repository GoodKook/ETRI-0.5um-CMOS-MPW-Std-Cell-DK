magic
tech scmos
magscale 1 60
timestamp 1709422372
<< checkpaint >>
rect 147100 672200 952620 677000
rect 140100 605700 952620 672200
rect 140100 600900 663108 605700
rect 147040 596560 663108 600900
rect 141400 596320 663108 596560
rect 135220 585368 663108 596320
rect 128800 584900 663108 585368
rect 128800 573954 663400 584900
rect 674260 577720 726780 590260
rect 128800 561414 666414 573954
rect 128800 555112 663400 561414
rect 110500 462584 663400 555112
rect 110500 444584 767640 462584
rect 110500 404530 663400 444584
rect 110500 316292 672200 404530
rect 82768 315260 672200 316292
rect 59274 288860 672200 315260
rect 62160 288654 672200 288860
rect 75556 278350 672200 288654
rect 110500 238750 672200 278350
rect 124042 235112 672200 238750
rect 110500 206750 672200 235112
rect 124042 173948 672200 206750
rect 101586 147100 672200 173948
rect 101586 128800 553500 147100
rect 558558 146716 645594 147100
rect 558558 130540 611800 146716
rect 558558 130300 611500 130540
rect 558558 130000 610540 130300
rect 558558 128800 587340 130000
rect 101586 127840 552958 128800
rect 101586 126030 182410 127840
rect 110910 113416 182410 126030
rect 109300 109300 111702 111702
rect 204796 110500 232958 127840
rect 236796 110500 265158 127840
rect 268796 110500 297158 127840
rect 300796 110500 552958 127840
use IOFILLER10  IOFILLER10_0 ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/chip_top/pads_ETRI050
timestamp 1537935238
transform 1 0 444678 0 1 148301
box -70 0 2070 50120
use IOFILLER10  IOFILLER10_1
timestamp 1537935238
transform 1 0 473438 0 1 148301
box -70 0 2070 50120
use IOFILLER10  IOFILLER10_2
timestamp 1537935238
transform 1 0 443038 0 1 148301
box -70 0 2070 50120
use IOFILLER10  IOFILLER10_3
timestamp 1537935238
transform 1 0 441438 0 1 148301
box -70 0 2070 50120
use IOFILLER10  IOFILLER10_4
timestamp 1537935238
transform 1 0 476678 0 1 148301
box -70 0 2070 50120
use IOFILLER10  IOFILLER10_5
timestamp 1537935238
transform 1 0 475038 0 1 148301
box -70 0 2070 50120
use IOFILLER40  IOFILLER40_0 ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/chip_top/pads_ETRI050
timestamp 1709340318
transform 1 0 263648 0 1 148300
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_1
timestamp 1709340318
transform 1 0 231648 0 1 148300
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_2
timestamp 1709340318
transform 1 0 327648 0 1 148300
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_3
timestamp 1709340318
transform 1 0 295648 0 1 148300
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_4
timestamp 1709340318
transform 1 0 391648 0 1 148300
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_5
timestamp 1709340318
transform 1 0 359648 0 1 148300
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_6
timestamp 1709340318
transform 1 0 455648 0 1 148300
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_7
timestamp 1709340318
transform 1 0 423648 0 1 148300
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_8
timestamp 1709340318
transform 1 0 519648 0 1 148300
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_9
timestamp 1709340318
transform 1 0 487648 0 1 148300
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_11
timestamp 1709340318
transform 1 0 263648 0 -1 611560
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_12
timestamp 1709340318
transform 1 0 231648 0 -1 611560
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_13
timestamp 1709340318
transform 1 0 327648 0 -1 611560
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_14
timestamp 1709340318
transform 1 0 295648 0 -1 611560
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_15
timestamp 1709340318
transform 1 0 391648 0 -1 611560
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_16
timestamp 1709340318
transform 1 0 359648 0 -1 611560
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_17
timestamp 1709340318
transform 1 0 455648 0 -1 611560
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_18
timestamp 1709340318
transform 1 0 423648 0 -1 611560
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_19
timestamp 1709340318
transform 1 0 519648 0 -1 611560
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_20
timestamp 1709340318
transform 1 0 487648 0 -1 611560
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_22
timestamp 1709340318
transform 0 1 148300 -1 0 304380
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_23
timestamp 1709340318
transform 0 1 148300 -1 0 240380
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_24
timestamp 1709340318
transform 0 1 148300 -1 0 272380
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_25
timestamp 1709340318
transform 0 1 148300 -1 0 400380
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_26
timestamp 1709340318
transform 0 1 148300 -1 0 336380
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_27
timestamp 1709340318
transform 0 1 148300 -1 0 368380
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_28
timestamp 1709340318
transform 0 1 148300 -1 0 464380
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_29
timestamp 1709340318
transform 0 1 148300 -1 0 432380
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_31
timestamp 1709340318
transform 0 1 148300 -1 0 496380
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_32
timestamp 1709340318
transform 0 1 148300 -1 0 528380
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_33
timestamp 1709340318
transform 0 -1 611610 1 0 295640
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_34
timestamp 1709340318
transform 0 -1 611610 1 0 231640
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_35
timestamp 1709340318
transform 0 -1 611610 1 0 263640
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_36
timestamp 1709340318
transform 0 -1 611610 1 0 391640
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_37
timestamp 1709340318
transform 0 -1 611610 1 0 327640
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_38
timestamp 1709340318
transform 0 -1 611610 1 0 359640
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_39
timestamp 1709340318
transform 0 -1 611610 1 0 455640
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_40
timestamp 1709340318
transform 0 -1 611610 1 0 423640
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_42
timestamp 1709340318
transform 0 -1 611610 1 0 487640
box 0 0 8720 50120
use IOFILLER40  IOFILLER40_43
timestamp 1709340318
transform 0 -1 611610 1 0 519640
box 0 0 8720 50120
use IOFILLER50  IOFILLER50_0 ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/chip_top/pads_ETRI050
timestamp 1537935238
transform 1 0 198120 0 1 148300
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_1
timestamp 1537935238
transform 1 0 551650 0 1 148300
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_2
timestamp 1537935238
transform 1 0 551650 0 -1 611560
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_3
timestamp 1537935238
transform 1 0 198128 0 -1 611560
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_4
timestamp 1537935238
transform 0 1 148300 -1 0 208260
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_5
timestamp 1537935238
transform 0 1 148300 -1 0 561780
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_6
timestamp 1537935238
transform 0 -1 611610 -1 0 208260
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_7
timestamp 1537935238
transform 0 -1 611608 -1 0 561832
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_8
timestamp 1537935238
transform 1 0 463818 0 1 148301
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_9
timestamp 1537935238
transform 1 0 446198 0 1 148300
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_10
timestamp 1537935238
transform 1 0 431818 0 1 148301
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_11
timestamp 1537935238
transform 1 0 478198 0 1 148300
box -70 0 10070 50120
use PCORNER  PCORNER_0 ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/chip_top/pads_ETRI050
timestamp 1537935238
transform 1 0 148300 0 1 148300
box 0 0 50600 50600
use PCORNER  PCORNER_1
timestamp 1537935238
transform 1 0 148302 0 -1 611560
box 0 0 50600 50600
use PCORNER  PCORNER_2
timestamp 1537935238
transform 0 -1 611610 1 0 148300
box 0 0 50600 50600
use PCORNER  PCORNER_3
timestamp 1537935238
transform -1 0 611608 0 -1 611560
box 0 0 50600 50600
use PAD80  PAD80_0 ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/chip_top/pads_ETRI050
timestamp 1709379016
transform 1 0 467458 0 1 130000
box 0 0 17000 17000
use PAD80  PAD80_1
timestamp 1709379016
transform 1 0 435458 0 1 130000
box 0 0 17000 17000
use PIC  CLK ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/chip_top/pads_ETRI050
timestamp 1537935238
transform 0 -1 611610 1 0 303950
box -200 -18300 24200 50600
use PIC  DI[0]
timestamp 1537935238
transform 1 0 399958 0 1 148300
box -200 -18300 24200 50600
use PIC  DI[1]
timestamp 1537935238
transform 0 -1 611610 1 0 431950
box -200 -18300 24200 50600
use PIC  DI[2]
timestamp 1537935238
transform 1 0 335958 0 1 148300
box -200 -18300 24200 50600
use PIC  DI[3]
timestamp 1537935238
transform 0 1 148300 -1 0 423950
box -200 -18300 24200 50600
use PIC  DI[4]
timestamp 1537935238
transform 1 0 239958 0 1 148300
box -200 -18300 24200 50600
use PIC  DI[5]
timestamp 1537935238
transform 0 1 148300 -1 0 455950
box -200 -18300 24200 50600
use PIC  DI[6]
timestamp 1537935238
transform 0 1 148300 -1 0 487950
box -200 -18300 24200 50600
use PIC  DI[7]
timestamp 1537935238
transform 0 1 148300 -1 0 551950
box -200 -18300 24200 50600
use PIC  IRQ
timestamp 1537935238
transform 0 -1 611610 1 0 207950
box -200 -18300 24200 50600
use PIC  NMI
timestamp 1537935238
transform 1 0 495958 0 1 148300
box -200 -18300 24200 50600
use PIC  RDY
timestamp 1537935238
transform 0 1 148300 -1 0 391950
box -200 -18300 24200 50600
use PIC  RESET
timestamp 1537935238
transform 0 -1 611610 1 0 239950
box -200 -18300 24200 50600
use POB8  AB[0] ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/chip_top/pads_ETRI050
timestamp 1537935238
transform 0 -1 611610 1 0 271950
box -200 -18300 24200 50600
use POB8  AB[1]
timestamp 1537935238
transform 1 0 271958 0 -1 611560
box -200 -18300 24200 50600
use POB8  AB[2]
timestamp 1537935238
transform 1 0 303958 0 -1 611560
box -200 -18300 24200 50600
use POB8  AB[3]
timestamp 1537935238
transform 1 0 463958 0 -1 611560
box -200 -18300 24200 50600
use POB8  AB[4]
timestamp 1537935238
transform 1 0 239958 0 -1 611560
box -200 -18300 24200 50600
use POB8  AB[5]
timestamp 1537935238
transform 1 0 399958 0 -1 611560
box -200 -18300 24200 50600
use POB8  AB[6]
timestamp 1537935238
transform 1 0 495958 0 -1 611560
box -200 -18300 24200 50600
use POB8  AB[7]
timestamp 1537935238
transform 1 0 431958 0 -1 611560
box -200 -18300 24200 50600
use POB8  AB[8]
timestamp 1537935238
transform 1 0 303958 0 1 148300
box -200 -18300 24200 50600
use POB8  AB[9]
timestamp 1537935238
transform 0 1 148300 -1 0 231950
box -200 -18300 24200 50600
use POB8  AB[10]
timestamp 1537935238
transform 1 0 271958 0 1 148300
box -200 -18300 24200 50600
use POB8  AB[11]
timestamp 1537935238
transform 0 1 148300 -1 0 263950
box -200 -18300 24200 50600
use POB8  AB[12]
timestamp 1537935238
transform 0 1 148300 -1 0 295950
box -200 -18300 24200 50600
use POB8  AB[13]
timestamp 1537935238
transform 0 1 148300 -1 0 327950
box -200 -18300 24200 50600
use POB8  AB[14]
timestamp 1537935238
transform 0 1 148300 -1 0 519950
box -200 -18300 24200 50600
use POB8  AB[15]
timestamp 1537935238
transform 0 1 148300 -1 0 359950
box -200 -18300 24200 50600
use POB8  DO[0]
timestamp 1537935238
transform 1 0 367958 0 -1 611560
box -200 -18300 24200 50600
use POB8  DO[1]
timestamp 1537935238
transform 0 -1 611610 1 0 335950
box -200 -18300 24200 50600
use POB8  DO[2]
timestamp 1537935238
transform 0 -1 611610 1 0 495950
box -200 -18300 24200 50600
use POB8  DO[3]
timestamp 1537935238
transform 0 -1 611610 1 0 367950
box -200 -18300 24200 50600
use POB8  DO[4]
timestamp 1537935238
transform 1 0 335958 0 -1 611560
box -200 -18300 24200 50600
use POB8  DO[5]
timestamp 1537935238
transform 0 -1 611610 1 0 527950
box -200 -18300 24200 50600
use POB8  DO[6]
timestamp 1537935238
transform 0 -1 611610 1 0 399950
box -200 -18300 24200 50600
use POB8  DO[7]
timestamp 1537935238
transform 0 -1 611610 1 0 463950
box -200 -18300 24200 50600
use POB8  WE
timestamp 1537935238
transform 1 0 367958 0 1 148300
box -200 -18300 24200 50600
use PVSS  PVSS_0 ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/chip_top/pads_ETRI050
timestamp 1537935238
transform 1 0 527958 0 -1 611560
box 0 -18300 24000 50600
use PVSS  PVSS_1
timestamp 1537935238
transform 1 0 527958 0 1 148300
box 0 -18300 24000 50600
use PVDD  PVDD_0 ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/chip_top/pads_ETRI050
timestamp 1537935238
transform 1 0 207958 0 -1 611560
box 0 -18300 24000 50600
use PVDD  PVDD_1
timestamp 1537935238
transform 1 0 207758 0 1 148300
box 0 -18300 24000 50600
use MY_LOGO  MY_LOGO_0
timestamp 1706263538
transform 1 0 555820 0 1 131500
box 14100 240 54780 15240
<< end >>