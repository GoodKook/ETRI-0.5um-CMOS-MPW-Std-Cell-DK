magic
tech scmos
magscale 1 3
timestamp 1537935238
<< checkpaint >>
rect -60 -60 78 100
<< genericcontact >>
rect 6 23 12 29
rect 6 11 12 17
<< metal1 >>
rect 0 0 18 40
<< pseudo_rpoly2 >>
rect 1 1 17 39
<< end >>
