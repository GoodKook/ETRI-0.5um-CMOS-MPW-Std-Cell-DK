VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO NOR3X1
  CLASS BLOCK ;
  FOREIGN NOR3X1 ;
  ORIGIN 2.100 0.900 ;
  SIZE 22.500 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 12.600000 ;
    PORT
      LAYER metal1 ;
        RECT 3.000 6.900 5.700 8.100 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 12.600000 ;
    PORT
      LAYER metal1 ;
        RECT 5.400 9.900 7.800 11.100 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 12.600000 ;
    PORT
      LAYER metal1 ;
        RECT 7.800 12.900 10.200 14.100 ;
    END
  END C
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 15.000 18.000 16.200 26.400 ;
        RECT 15.000 17.100 15.900 18.000 ;
        RECT 15.000 16.800 16.200 17.100 ;
        RECT 11.100 15.900 16.200 16.800 ;
        RECT 11.100 6.000 12.000 15.900 ;
        RECT 6.000 5.100 12.000 6.000 ;
        RECT 6.000 4.800 6.900 5.100 ;
        RECT 5.400 3.900 6.900 4.800 ;
        RECT 10.200 4.800 12.000 5.100 ;
        RECT 5.400 1.800 6.600 3.900 ;
        RECT 10.200 1.800 11.400 4.800 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 19.800 30.900 ;
        RECT 3.000 19.200 4.200 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 3.000 0.900 4.200 4.800 ;
        RECT 7.800 0.900 9.000 4.200 ;
        RECT -0.600 -0.900 19.800 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 19.200 1.800 28.200 ;
        RECT 0.900 18.300 1.800 19.200 ;
        RECT 5.400 27.300 11.400 28.200 ;
        RECT 5.400 19.200 6.600 27.300 ;
        RECT 7.800 19.200 9.000 26.400 ;
        RECT 10.200 19.500 11.400 27.300 ;
        RECT 12.900 27.300 18.300 28.200 ;
        RECT 12.900 27.000 13.800 27.300 ;
        RECT 5.400 18.300 6.300 19.200 ;
        RECT 0.900 17.400 6.300 18.300 ;
        RECT 8.100 18.600 9.000 19.200 ;
        RECT 12.600 18.600 13.800 27.000 ;
        RECT 8.100 18.000 13.800 18.600 ;
        RECT 17.400 27.000 18.300 27.300 ;
        RECT 17.400 18.000 18.600 27.000 ;
        RECT 8.100 17.700 13.500 18.000 ;
  END
END NOR3X1
MACRO DFFNEGX1
  CLASS BLOCK ;
  FOREIGN DFFNEGX1 ;
  ORIGIN 2.400 0.900 ;
  SIZE 33.600 BY 32.400 ;
  PIN D
    ANTENNAGATEAREA 5.400000 ;
    PORT
      LAYER metal1 ;
        RECT 10.200 13.800 11.400 14.100 ;
        RECT 4.200 12.900 11.400 13.800 ;
        RECT 4.200 12.600 5.400 12.900 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 21.600000 ;
    PORT
      LAYER metal1 ;
        RECT 8.100 20.100 9.300 21.300 ;
        RECT 7.800 18.900 9.000 20.100 ;
        RECT 7.800 11.100 9.000 11.400 ;
        RECT 1.800 10.200 19.200 11.100 ;
        RECT 1.800 9.900 4.200 10.200 ;
        RECT 6.000 8.100 7.200 10.200 ;
        RECT 18.000 9.900 19.200 10.200 ;
        RECT 6.300 6.900 7.500 8.100 ;
      LAYER via1 ;
        RECT 7.800 10.200 9.000 11.400 ;
      LAYER metal2 ;
        RECT 7.800 10.200 9.000 20.100 ;
    END
  END CLK
  PIN Q
    ANTENNAGATEAREA 3.600000 ;
    PORT
      LAYER metal1 ;
        RECT 27.000 15.300 28.200 28.200 ;
        RECT 21.900 14.400 28.200 15.300 ;
        RECT 21.900 14.100 23.100 14.400 ;
        RECT 27.000 9.300 28.200 14.400 ;
        RECT 22.500 8.400 28.200 9.300 ;
        RECT 22.500 8.100 23.700 8.400 ;
        RECT 27.000 1.800 28.200 8.400 ;
    END
  END Q
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 29.400 30.900 ;
        RECT 3.000 16.500 4.200 29.100 ;
        RECT 11.400 22.200 12.600 29.100 ;
        RECT 16.200 22.200 17.400 29.100 ;
        RECT 24.600 16.200 25.800 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 3.000 0.900 4.200 7.800 ;
        RECT 11.100 0.900 12.600 4.800 ;
        RECT 16.200 0.900 17.400 4.800 ;
        RECT 24.600 0.900 25.800 7.500 ;
        RECT -0.600 -0.900 29.400 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 15.600 1.800 28.200 ;
        RECT 7.200 23.100 8.400 28.200 ;
        RECT 5.400 22.200 8.400 23.100 ;
        RECT 13.800 22.200 15.000 28.200 ;
        RECT 20.100 22.200 21.900 28.200 ;
        RECT 5.400 21.000 6.600 22.200 ;
        RECT 13.800 21.300 14.700 22.200 ;
        RECT 10.500 20.400 15.900 21.300 ;
        RECT 19.800 21.000 21.000 22.200 ;
        RECT 10.500 20.100 11.700 20.400 ;
        RECT 14.700 20.100 15.900 20.400 ;
        RECT 5.400 18.000 6.600 18.300 ;
        RECT 12.300 18.000 13.500 18.300 ;
        RECT 5.400 17.100 13.500 18.000 ;
        RECT 16.200 18.000 17.700 18.300 ;
        RECT 20.700 18.000 21.900 18.300 ;
        RECT 16.200 17.100 21.900 18.000 ;
        RECT 16.200 16.200 17.100 17.100 ;
        RECT 6.300 15.600 17.100 16.200 ;
        RECT 0.600 15.300 17.100 15.600 ;
        RECT 0.600 14.700 7.500 15.300 ;
        RECT 24.300 13.200 25.500 13.500 ;
        RECT 19.800 12.300 25.500 13.200 ;
        RECT 19.800 12.000 21.000 12.300 ;
        RECT 0.600 1.800 1.800 9.000 ;
        RECT 10.500 6.600 11.700 6.900 ;
        RECT 5.400 4.800 6.600 6.000 ;
        RECT 10.500 5.700 14.700 6.600 ;
        RECT 13.800 4.800 14.700 5.700 ;
        RECT 19.800 4.800 21.000 6.000 ;
        RECT 5.400 3.900 8.400 4.800 ;
        RECT 7.200 1.800 8.400 3.900 ;
        RECT 13.800 1.800 15.000 4.800 ;
        RECT 19.800 3.900 21.900 4.800 ;
        RECT 20.100 1.800 21.900 3.900 ;
      LAYER via1 ;
        RECT 0.600 15.000 1.800 16.200 ;
        RECT 0.600 7.800 1.800 9.000 ;
      LAYER metal2 ;
        RECT 5.400 16.200 6.600 22.200 ;
        RECT 19.800 18.300 21.000 22.200 ;
        RECT 19.800 17.100 20.700 18.300 ;
        RECT 0.600 7.800 1.800 16.200 ;
        RECT 5.400 15.000 6.300 16.200 ;
        RECT 5.400 4.800 6.600 15.000 ;
        RECT 19.800 4.800 21.000 17.100 ;
  END
END DFFNEGX1
MACRO FILL
  CLASS BLOCK ;
  FOREIGN FILL ;
  ORIGIN 2.400 0.900 ;
  SIZE 7.200 BY 32.400 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 3.000 30.900 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT -0.600 -0.900 3.000 0.900 ;
    END
  END gnd
END FILL
MACRO BUFX4
  CLASS BLOCK ;
  FOREIGN BUFX4 ;
  ORIGIN 2.700 0.900 ;
  SIZE 13.800 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 8.100000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 12.900 2.100 14.100 ;
        RECT 0.900 11.700 2.100 12.900 ;
    END
  END A
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 5.400 17.700 6.600 28.200 ;
        RECT 5.400 16.200 6.900 17.700 ;
        RECT 6.000 11.100 6.900 16.200 ;
        RECT 5.400 9.900 6.900 11.100 ;
        RECT 6.000 7.800 6.900 9.900 ;
        RECT 5.400 6.900 6.900 7.800 ;
        RECT 5.400 1.800 6.600 6.900 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 10.200 30.900 ;
        RECT 3.000 18.000 4.200 29.100 ;
        RECT 7.800 16.200 9.000 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 3.000 0.900 4.200 7.800 ;
        RECT 7.800 0.900 9.000 7.800 ;
        RECT -0.600 -0.900 10.200 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 17.100 1.800 28.200 ;
        RECT 0.600 16.200 4.500 17.100 ;
        RECT 3.600 13.200 4.500 16.200 ;
        RECT 3.600 12.000 5.100 13.200 ;
        RECT 3.600 9.600 4.500 12.000 ;
        RECT 0.600 8.700 4.500 9.600 ;
        RECT 0.600 1.800 1.800 8.700 ;
  END
END BUFX4
MACRO BUFX2
  CLASS BLOCK ;
  FOREIGN BUFX2 ;
  ORIGIN 1.500 0.900 ;
  SIZE 9.900 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 5.400000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 11.700 1.800 14.100 ;
    END
  END A
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 5.400 16.200 6.600 28.200 ;
        RECT 5.700 12.900 6.600 16.200 ;
        RECT 5.400 1.800 6.600 12.900 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 7.800 30.900 ;
        RECT 3.000 18.000 4.200 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 3.000 0.900 4.200 7.800 ;
        RECT -0.600 -0.900 7.800 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 17.100 1.800 28.200 ;
        RECT 0.600 16.200 3.900 17.100 ;
        RECT 3.000 15.300 3.900 16.200 ;
        RECT 3.000 14.100 4.800 15.300 ;
        RECT 3.000 9.600 3.900 14.100 ;
        RECT 0.600 8.700 3.900 9.600 ;
        RECT 0.600 1.800 1.800 8.700 ;
  END
END BUFX2
MACRO AOI22X1
  CLASS BLOCK ;
  FOREIGN AOI22X1 ;
  ORIGIN 2.400 0.900 ;
  SIZE 16.200 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 10.800000 ;
    PORT
      LAYER metal1 ;
        RECT 1.800 14.100 3.000 14.700 ;
        RECT 0.600 13.200 3.000 14.100 ;
        RECT 0.600 12.900 1.800 13.200 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 10.800000 ;
    PORT
      LAYER metal1 ;
        RECT 3.000 9.900 4.200 12.300 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 10.800000 ;
    PORT
      LAYER metal1 ;
        RECT 10.200 12.900 11.400 15.300 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA 10.800000 ;
    PORT
      LAYER metal1 ;
        RECT 7.500 11.700 8.700 12.900 ;
        RECT 7.800 11.100 8.700 11.700 ;
        RECT 7.800 9.900 9.000 11.100 ;
    END
  END D
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 7.800 16.200 9.000 26.400 ;
        RECT 7.800 15.300 8.700 16.200 ;
        RECT 5.700 14.400 8.700 15.300 ;
        RECT 5.700 14.100 6.600 14.400 ;
        RECT 5.400 12.900 6.600 14.100 ;
        RECT 5.700 7.800 6.600 12.900 ;
        RECT 5.100 1.800 7.500 7.800 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 12.600 30.900 ;
        RECT 3.000 18.000 4.200 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 1.200 0.900 2.400 7.800 ;
        RECT 10.200 0.900 11.400 7.800 ;
        RECT -0.600 -0.900 12.600 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 17.100 1.800 28.200 ;
        RECT 5.400 27.300 11.400 28.200 ;
        RECT 5.400 17.100 6.600 27.300 ;
        RECT 0.600 16.200 6.600 17.100 ;
        RECT 10.200 16.200 11.400 27.300 ;
  END
END AOI22X1
MACRO AOI21X1
  CLASS BLOCK ;
  FOREIGN AOI21X1 ;
  ORIGIN 2.100 0.900 ;
  SIZE 13.800 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 10.800000 ;
    PORT
      LAYER metal1 ;
        RECT 1.800 14.100 3.000 14.700 ;
        RECT 0.600 13.200 3.000 14.100 ;
        RECT 0.600 12.900 1.800 13.200 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 10.800000 ;
    PORT
      LAYER metal1 ;
        RECT 3.000 9.900 4.200 12.300 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 9.000000 ;
    PORT
      LAYER metal1 ;
        RECT 7.800 6.900 9.000 8.100 ;
        RECT 7.500 5.700 8.700 6.900 ;
    END
  END C
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 7.800 16.200 9.000 28.200 ;
        RECT 7.800 14.100 8.700 16.200 ;
        RECT 5.400 13.200 9.000 14.100 ;
        RECT 5.400 7.800 6.300 13.200 ;
        RECT 7.800 12.900 9.000 13.200 ;
        RECT 5.400 1.800 6.600 7.800 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 10.200 30.900 ;
        RECT 3.000 18.000 4.200 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 1.500 0.900 2.700 7.800 ;
        RECT 7.800 0.900 9.000 4.800 ;
        RECT -0.600 -0.900 10.200 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 17.100 1.800 28.200 ;
        RECT 5.400 17.100 6.600 28.200 ;
        RECT 0.600 16.200 6.600 17.100 ;
  END
END AOI21X1
MACRO AND2X2
  CLASS BLOCK ;
  FOREIGN AND2X2 ;
  ORIGIN 2.400 0.900 ;
  SIZE 14.400 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 7.200000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 9.900 1.800 12.300 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 7.200000 ;
    PORT
      LAYER metal1 ;
        RECT 3.000 12.900 4.200 14.100 ;
        RECT 3.300 11.700 4.200 12.900 ;
        RECT 3.300 10.800 4.800 11.700 ;
        RECT 3.600 10.500 4.800 10.800 ;
    END
  END B
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 7.800 16.200 9.000 28.200 ;
        RECT 8.100 14.100 9.000 16.200 ;
        RECT 7.800 12.900 9.000 14.100 ;
        RECT 8.100 7.800 9.000 12.900 ;
        RECT 6.900 6.300 9.000 7.800 ;
        RECT 6.900 1.800 8.100 6.300 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 10.200 30.900 ;
        RECT 0.600 22.200 1.800 29.100 ;
        RECT 5.400 16.800 6.600 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 4.500 0.900 5.700 7.500 ;
        RECT -0.600 -0.900 10.200 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 3.000 22.200 4.200 28.200 ;
        RECT 3.300 15.900 4.200 22.200 ;
        RECT 3.300 15.000 6.900 15.900 ;
        RECT 6.000 9.900 6.900 15.000 ;
        RECT 6.000 9.600 7.200 9.900 ;
        RECT 2.700 9.000 7.200 9.600 ;
        RECT 0.900 8.700 7.200 9.000 ;
        RECT 0.900 8.100 3.600 8.700 ;
        RECT 0.900 7.800 1.800 8.100 ;
        RECT 0.600 1.800 1.800 7.800 ;
  END
END AND2X2
MACRO AND2X1
  CLASS BLOCK ;
  FOREIGN AND2X1 ;
  ORIGIN 2.400 0.900 ;
  SIZE 14.400 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 7.200000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 9.900 1.800 12.300 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 7.200000 ;
    PORT
      LAYER metal1 ;
        RECT 3.000 15.900 5.100 17.100 ;
        RECT 3.900 14.700 5.100 15.900 ;
    END
  END B
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 7.800 22.200 9.000 28.200 ;
        RECT 8.100 20.100 9.000 22.200 ;
        RECT 7.800 18.900 9.000 20.100 ;
        RECT 8.100 5.700 9.000 18.900 ;
        RECT 6.900 4.800 9.000 5.700 ;
        RECT 6.900 1.800 8.100 4.800 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 10.200 30.900 ;
        RECT 0.600 22.200 1.800 29.100 ;
        RECT 5.400 22.200 6.600 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 4.500 0.900 5.700 7.800 ;
        RECT -0.600 -0.900 10.200 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 3.000 22.200 4.200 28.200 ;
        RECT 3.300 21.300 4.200 22.200 ;
        RECT 3.300 20.400 6.900 21.300 ;
        RECT 6.000 9.900 6.900 20.400 ;
        RECT 2.700 9.000 7.200 9.900 ;
        RECT 2.700 8.700 3.600 9.000 ;
        RECT 6.000 8.700 7.200 9.000 ;
        RECT 0.900 7.800 3.600 8.700 ;
        RECT 0.600 1.800 1.800 7.800 ;
  END
END AND2X1
MACRO INVX8
  CLASS BLOCK ;
  FOREIGN INVX8 ;
  ORIGIN 2.700 0.900 ;
  SIZE 16.200 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 43.200001 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 8.700 1.800 11.100 ;
    END
  END A
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 3.000 15.300 4.200 28.200 ;
        RECT 7.800 15.300 9.000 28.200 ;
        RECT 3.000 14.100 9.000 15.300 ;
        RECT 7.800 9.900 9.000 14.100 ;
        RECT 3.000 8.700 9.000 9.900 ;
        RECT 3.000 1.800 4.200 8.700 ;
        RECT 7.800 1.800 9.000 8.700 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 12.600 30.900 ;
        RECT 0.600 16.200 1.800 29.100 ;
        RECT 5.400 16.200 6.600 29.100 ;
        RECT 10.200 16.200 11.400 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 0.900 1.800 7.800 ;
        RECT 5.400 0.900 6.600 7.800 ;
        RECT 10.200 0.900 11.400 7.800 ;
        RECT -0.600 -0.900 12.600 0.900 ;
    END
  END gnd
END INVX8
MACRO INVX4
  CLASS BLOCK ;
  FOREIGN INVX4 ;
  ORIGIN 2.700 0.900 ;
  SIZE 11.100 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 21.600000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 8.700 1.800 11.100 ;
    END
  END A
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 3.000 1.800 4.200 28.200 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 7.800 30.900 ;
        RECT 0.600 16.200 1.800 29.100 ;
        RECT 5.400 16.200 6.600 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 0.900 1.800 7.800 ;
        RECT 5.400 0.900 6.600 7.800 ;
        RECT -0.600 -0.900 7.800 0.900 ;
    END
  END gnd
END INVX4
MACRO INVX2
  CLASS BLOCK ;
  FOREIGN INVX2 ;
  ORIGIN 2.700 0.900 ;
  SIZE 10.500 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 10.800000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 8.700 1.800 11.100 ;
    END
  END A
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 3.000 1.800 4.200 28.200 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 5.400 30.900 ;
        RECT 0.600 16.200 1.800 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 0.900 1.800 7.800 ;
        RECT -0.600 -0.900 5.400 0.900 ;
    END
  END gnd
END INVX2
MACRO INVX1
  CLASS BLOCK ;
  FOREIGN INVX1 ;
  ORIGIN 2.700 0.900 ;
  SIZE 10.500 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 5.400000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 5.700 1.800 8.100 ;
    END
  END A
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 3.000 1.800 4.200 28.200 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 5.400 30.900 ;
        RECT 0.600 22.200 1.800 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 0.900 1.800 4.800 ;
        RECT -0.600 -0.900 5.400 0.900 ;
    END
  END gnd
END INVX1
MACRO HAX1
  CLASS BLOCK ;
  FOREIGN HAX1 ;
  ORIGIN 1.500 0.900 ;
  SIZE 26.700 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 18.000000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 9.900 1.800 11.100 ;
        RECT 15.000 10.800 16.200 11.100 ;
        RECT 12.600 9.900 16.200 10.800 ;
        RECT 0.600 9.000 13.500 9.900 ;
        RECT 1.200 8.700 2.400 9.000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 18.000000 ;
    PORT
      LAYER metal1 ;
        RECT 3.000 12.900 4.200 14.100 ;
        RECT 3.300 12.000 4.500 12.900 ;
        RECT 12.600 12.600 13.800 12.900 ;
        RECT 3.600 11.700 4.800 12.000 ;
        RECT 10.800 11.700 13.800 12.600 ;
        RECT 3.600 10.800 11.700 11.700 ;
    END
  END B
  PIN YC
    PORT
      LAYER metal1 ;
        RECT 7.800 12.600 9.000 28.200 ;
        RECT 6.900 1.800 8.100 6.000 ;
      LAYER via1 ;
        RECT 6.900 4.800 8.100 6.000 ;
      LAYER metal2 ;
        RECT 7.800 12.600 9.000 13.800 ;
        RECT 8.100 6.000 9.000 12.600 ;
        RECT 6.900 4.800 9.000 6.000 ;
    END
  END YC
  PIN YS
    PORT
      LAYER metal1 ;
        RECT 21.300 22.200 22.500 28.200 ;
        RECT 21.600 21.300 22.500 22.200 ;
        RECT 20.100 20.400 22.500 21.300 ;
        RECT 20.100 17.100 21.000 20.400 ;
        RECT 19.800 15.900 21.000 17.100 ;
        RECT 20.100 6.900 21.000 15.900 ;
        RECT 20.100 6.000 22.500 6.900 ;
        RECT 21.600 4.800 22.500 6.000 ;
        RECT 21.300 1.800 22.500 4.800 ;
    END
  END YS
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 24.600 30.900 ;
        RECT 3.000 22.800 4.200 29.100 ;
        RECT 10.200 22.200 11.400 29.100 ;
        RECT 16.500 16.200 17.700 29.100 ;
        RECT 18.900 22.200 20.100 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 0.900 1.800 7.800 ;
        RECT 9.300 0.900 10.500 7.500 ;
        RECT 18.900 0.900 20.100 4.800 ;
        RECT -0.600 -0.900 24.600 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 22.200 1.800 28.200 ;
        RECT 0.900 21.900 1.800 22.200 ;
        RECT 5.400 21.900 6.600 28.200 ;
        RECT 0.900 21.000 6.600 21.900 ;
        RECT 5.700 13.800 6.600 21.000 ;
        RECT 12.600 16.200 13.800 28.200 ;
        RECT 12.900 15.300 13.800 16.200 ;
        RECT 12.900 14.400 18.000 15.300 ;
        RECT 5.700 12.600 6.900 13.800 ;
        RECT 17.100 9.300 18.000 14.400 ;
        RECT 17.100 9.000 18.900 9.300 ;
        RECT 14.400 8.100 18.900 9.000 ;
        RECT 5.700 7.800 8.400 8.100 ;
        RECT 14.400 7.800 15.300 8.100 ;
        RECT 4.500 6.900 8.400 7.800 ;
        RECT 4.500 1.800 5.700 6.900 ;
        RECT 11.700 2.700 12.900 7.800 ;
        RECT 14.100 3.600 15.300 7.800 ;
        RECT 16.500 2.700 17.700 7.200 ;
        RECT 11.700 1.800 17.700 2.700 ;
      LAYER via1 ;
        RECT 5.700 6.900 6.900 8.100 ;
      LAYER metal2 ;
        RECT 5.700 12.600 6.900 13.800 ;
        RECT 5.700 8.100 6.600 12.600 ;
        RECT 5.700 6.900 6.900 8.100 ;
  END
END HAX1
MACRO FAX1
  CLASS BLOCK ;
  FOREIGN FAX1 ;
  ORIGIN 1.500 0.900 ;
  SIZE 39.300 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 44.640003 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 9.900 1.800 11.100 ;
        RECT 26.700 10.200 27.900 11.400 ;
        RECT 0.900 9.600 3.000 9.900 ;
        RECT 0.900 9.300 12.300 9.600 ;
        RECT 26.700 9.300 27.600 10.200 ;
        RECT 0.900 9.000 27.600 9.300 ;
        RECT 1.800 8.700 27.600 9.000 ;
        RECT 11.100 8.400 27.600 8.700 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 43.920002 ;
    PORT
      LAYER metal1 ;
        RECT 3.000 12.900 4.200 14.100 ;
        RECT 3.300 11.700 4.200 12.900 ;
        RECT 3.300 11.400 5.400 11.700 ;
        RECT 8.700 11.400 9.900 11.700 ;
        RECT 3.300 11.100 15.300 11.400 ;
        RECT 24.000 11.100 25.200 11.400 ;
        RECT 3.300 10.800 25.200 11.100 ;
        RECT 4.200 10.500 25.200 10.800 ;
        RECT 14.100 10.200 25.200 10.500 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 33.120003 ;
    PORT
      LAYER metal1 ;
        RECT 5.400 13.800 7.800 14.100 ;
        RECT 5.400 13.500 16.500 13.800 ;
        RECT 5.400 13.200 17.700 13.500 ;
        RECT 5.400 12.900 22.800 13.200 ;
        RECT 15.600 12.300 22.800 12.900 ;
        RECT 21.600 12.000 22.800 12.300 ;
    END
  END C
  PIN YS
    PORT
      LAYER metal1 ;
        RECT 29.400 23.100 30.600 28.200 ;
        RECT 29.100 22.200 30.600 23.100 ;
        RECT 29.100 14.700 30.000 22.200 ;
        RECT 29.100 13.800 32.100 14.700 ;
        RECT 31.200 8.100 32.100 13.800 ;
        RECT 31.200 6.900 33.000 8.100 ;
        RECT 31.200 6.600 32.100 6.900 ;
        RECT 29.700 5.700 32.100 6.600 ;
        RECT 29.700 4.800 30.600 5.700 ;
        RECT 29.400 1.800 30.600 4.800 ;
    END
  END YS
  PIN YC
    PORT
      LAYER metal1 ;
        RECT 34.200 22.200 35.400 28.200 ;
        RECT 34.500 11.100 35.400 22.200 ;
        RECT 34.200 9.900 35.400 11.100 ;
        RECT 34.500 4.800 35.400 9.900 ;
        RECT 34.200 1.800 35.400 4.800 ;
    END
  END YC
  OBS
      LAYER metal1 ;
        RECT -0.600 29.100 36.600 30.900 ;
        RECT 0.600 17.100 1.800 28.200 ;
        RECT 3.000 18.000 4.200 29.100 ;
        RECT 5.400 17.100 6.600 28.200 ;
        RECT 0.600 16.200 6.600 17.100 ;
        RECT 7.800 16.200 9.000 28.200 ;
        RECT 11.700 16.200 12.900 29.100 ;
        RECT 14.100 18.300 15.300 28.200 ;
        RECT 16.500 19.200 17.700 29.100 ;
        RECT 18.900 18.300 20.100 28.200 ;
        RECT 14.100 17.400 20.100 18.300 ;
        RECT 14.100 16.200 15.300 17.400 ;
        RECT 18.000 15.300 19.200 15.600 ;
        RECT 21.300 15.300 22.800 28.200 ;
        RECT 18.000 14.400 20.400 15.300 ;
        RECT 19.200 14.100 20.400 14.400 ;
        RECT 21.600 14.100 22.800 15.300 ;
        RECT 27.000 13.800 28.200 29.100 ;
        RECT 31.800 22.200 33.000 29.100 ;
        RECT 31.200 15.900 33.600 17.100 ;
        RECT 29.100 10.500 30.300 12.900 ;
        RECT 0.600 6.900 6.600 7.800 ;
        RECT 0.600 1.800 1.800 6.900 ;
        RECT 3.000 0.900 4.200 6.000 ;
        RECT 5.400 1.800 6.600 6.900 ;
        RECT 7.800 1.800 9.000 7.800 ;
        RECT 11.700 0.900 12.900 7.200 ;
        RECT 14.100 6.600 20.100 7.500 ;
        RECT 14.100 1.800 15.300 6.600 ;
        RECT 16.500 0.900 17.700 5.700 ;
        RECT 18.900 1.800 20.100 6.600 ;
        RECT 21.600 6.300 22.800 7.500 ;
        RECT 21.300 1.800 22.800 6.300 ;
        RECT 27.000 0.900 28.200 7.500 ;
        RECT 31.800 0.900 33.000 4.800 ;
        RECT -0.600 -0.900 36.600 0.900 ;
      LAYER via1 ;
        RECT 29.100 11.700 30.300 12.900 ;
        RECT 7.800 6.600 9.000 7.800 ;
      LAYER metal2 ;
        RECT 7.800 17.100 9.000 17.400 ;
        RECT 7.800 16.200 32.400 17.100 ;
        RECT 8.100 7.800 9.000 16.200 ;
        RECT 18.000 14.400 19.200 16.200 ;
        RECT 31.200 15.900 32.400 16.200 ;
        RECT 21.600 14.100 22.800 15.300 ;
        RECT 7.800 6.600 9.000 7.800 ;
        RECT 21.900 12.600 22.800 14.100 ;
        RECT 29.100 12.600 30.300 12.900 ;
        RECT 21.900 11.700 30.300 12.600 ;
        RECT 21.900 7.500 22.800 11.700 ;
        RECT 21.600 6.300 22.800 7.500 ;
  END
END FAX1
MACRO DFFPOSX1
  CLASS BLOCK ;
  FOREIGN DFFPOSX1 ;
  ORIGIN 2.400 0.900 ;
  SIZE 33.600 BY 32.400 ;
  PIN D
    ANTENNAGATEAREA 5.400000 ;
    PORT
      LAYER metal1 ;
        RECT 10.200 13.800 11.400 14.100 ;
        RECT 3.900 12.900 11.400 13.800 ;
        RECT 3.900 12.600 5.100 12.900 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 19.800001 ;
    PORT
      LAYER metal1 ;
        RECT 20.100 18.300 22.200 19.500 ;
        RECT 20.100 16.800 21.000 18.300 ;
        RECT 17.400 15.900 21.000 16.800 ;
        RECT 6.300 11.100 7.500 11.400 ;
        RECT 17.400 11.100 18.300 15.900 ;
        RECT 1.800 10.200 18.300 11.100 ;
        RECT 1.800 9.900 4.200 10.200 ;
        RECT 8.100 6.900 9.000 10.200 ;
        RECT 16.500 9.900 17.700 10.200 ;
        RECT 7.800 5.700 9.000 6.900 ;
    END
  END CLK
  PIN Q
    ANTENNAGATEAREA 3.600000 ;
    PORT
      LAYER metal1 ;
        RECT 27.000 15.300 28.200 28.200 ;
        RECT 21.900 14.400 28.200 15.300 ;
        RECT 21.900 14.100 23.100 14.400 ;
        RECT 27.000 9.300 28.200 14.400 ;
        RECT 22.500 8.400 28.200 9.300 ;
        RECT 22.500 8.100 23.700 8.400 ;
        RECT 27.000 1.800 28.200 8.400 ;
    END
  END Q
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 29.400 30.900 ;
        RECT 3.000 16.500 4.200 29.100 ;
        RECT 11.400 22.200 12.600 29.100 ;
        RECT 16.200 22.200 17.400 29.100 ;
        RECT 24.600 16.200 25.800 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 3.000 0.900 4.200 7.800 ;
        RECT 11.100 0.900 12.600 4.800 ;
        RECT 16.200 0.900 17.400 4.800 ;
        RECT 24.600 0.900 25.800 7.500 ;
        RECT -0.600 -0.900 29.400 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 15.600 1.800 28.200 ;
        RECT 7.200 23.100 8.400 28.200 ;
        RECT 5.400 22.200 8.400 23.100 ;
        RECT 13.800 22.200 15.000 28.200 ;
        RECT 20.100 22.200 21.900 28.200 ;
        RECT 5.400 21.000 6.600 22.200 ;
        RECT 13.800 21.300 14.700 22.200 ;
        RECT 10.500 20.400 15.900 21.300 ;
        RECT 19.800 21.000 21.000 22.200 ;
        RECT 10.500 20.100 11.700 20.400 ;
        RECT 14.700 20.100 15.900 20.400 ;
        RECT 5.400 18.000 6.600 18.300 ;
        RECT 12.300 18.000 13.500 18.300 ;
        RECT 5.400 17.100 13.500 18.000 ;
        RECT 14.400 18.000 17.700 18.900 ;
        RECT 14.400 16.200 15.300 18.000 ;
        RECT 16.500 17.700 17.700 18.000 ;
        RECT 8.100 15.600 15.300 16.200 ;
        RECT 0.600 15.300 15.300 15.600 ;
        RECT 0.600 15.000 9.300 15.300 ;
        RECT 0.600 14.700 9.000 15.000 ;
        RECT 24.300 13.200 25.500 13.500 ;
        RECT 19.800 12.300 25.500 13.200 ;
        RECT 19.800 12.000 21.000 12.300 ;
        RECT 0.600 1.800 1.800 9.000 ;
        RECT 10.500 6.600 11.700 6.900 ;
        RECT 5.400 4.800 6.600 6.000 ;
        RECT 10.500 5.700 14.700 6.600 ;
        RECT 13.800 4.800 14.700 5.700 ;
        RECT 19.800 4.800 21.000 6.000 ;
        RECT 5.400 3.900 8.400 4.800 ;
        RECT 7.200 1.800 8.400 3.900 ;
        RECT 13.800 1.800 15.000 4.800 ;
        RECT 19.800 3.900 21.900 4.800 ;
        RECT 20.100 1.800 21.900 3.900 ;
      LAYER via1 ;
        RECT 0.600 7.800 1.800 9.000 ;
      LAYER metal2 ;
        RECT 0.600 7.800 1.800 16.200 ;
        RECT 5.400 4.800 6.600 22.200 ;
        RECT 19.800 4.800 21.000 22.200 ;
  END
END DFFPOSX1
MACRO MUX2X1
  CLASS BLOCK ;
  FOREIGN MUX2X1 ;
  ORIGIN 1.500 0.900 ;
  SIZE 17.400 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 10.800000 ;
    PORT
      LAYER metal1 ;
        RECT 10.200 12.900 11.400 15.300 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 10.800000 ;
    PORT
      LAYER metal1 ;
        RECT 3.000 11.700 4.200 14.100 ;
    END
  END B
  PIN S
    ANTENNAGATEAREA 16.200001 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 11.700 1.800 14.100 ;
    END
  END S
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 6.900 17.700 8.100 28.200 ;
        RECT 6.900 16.800 9.300 17.700 ;
        RECT 8.400 11.100 9.300 16.800 ;
        RECT 8.400 9.900 11.400 11.100 ;
        RECT 8.400 9.000 9.300 9.900 ;
        RECT 8.100 8.400 9.300 9.000 ;
        RECT 6.900 7.500 9.300 8.400 ;
        RECT 6.900 3.000 8.100 7.500 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 15.000 30.900 ;
        RECT 3.000 16.800 4.200 29.100 ;
        RECT 10.800 16.200 12.000 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 3.000 0.900 4.200 8.400 ;
        RECT 10.800 0.900 12.000 9.000 ;
        RECT -0.600 -0.900 15.000 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 21.000 1.800 27.000 ;
        RECT 0.600 15.900 1.500 21.000 ;
        RECT 0.600 15.000 6.300 15.900 ;
        RECT 5.400 12.000 6.300 15.000 ;
        RECT 5.400 10.800 7.500 12.000 ;
        RECT 5.400 10.200 6.900 10.800 ;
        RECT 0.600 9.300 6.900 10.200 ;
        RECT 0.600 6.000 1.500 9.300 ;
        RECT 0.600 3.000 1.800 6.000 ;
  END
END MUX2X1
MACRO XOR2X1
  CLASS BLOCK ;
  FOREIGN XOR2X1 ;
  ORIGIN 2.400 0.900 ;
  SIZE 21.600 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 21.600000 ;
    PORT
      LAYER metal1 ;
        RECT 6.000 11.400 7.200 11.700 ;
        RECT 3.000 11.100 7.200 11.400 ;
        RECT 0.600 10.500 7.200 11.100 ;
        RECT 0.600 10.200 3.900 10.500 ;
        RECT 0.600 9.900 3.000 10.200 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 21.600000 ;
    PORT
      LAYER metal1 ;
        RECT 13.800 9.900 16.200 11.100 ;
    END
  END B
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 7.200 16.200 9.600 28.200 ;
        RECT 8.100 14.100 9.000 16.200 ;
        RECT 7.800 12.900 9.000 14.100 ;
        RECT 8.100 11.100 9.000 12.900 ;
        RECT 8.100 10.200 9.600 11.100 ;
        RECT 8.700 7.200 9.600 10.200 ;
        RECT 7.200 1.800 9.600 7.200 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 17.400 30.900 ;
        RECT 3.300 28.200 4.500 29.100 ;
        RECT 3.000 18.300 4.500 28.200 ;
        RECT 12.300 18.300 13.800 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 3.000 1.800 4.500 6.900 ;
        RECT 3.300 0.900 4.500 1.800 ;
        RECT 12.300 0.900 13.800 6.900 ;
        RECT -0.600 -0.900 17.400 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 17.100 1.800 28.200 ;
        RECT 3.300 17.100 4.500 17.400 ;
        RECT 0.600 16.200 4.500 17.100 ;
        RECT 12.600 17.100 13.800 17.400 ;
        RECT 15.000 17.100 16.200 28.200 ;
        RECT 12.600 16.200 16.200 17.100 ;
        RECT 5.100 14.100 6.300 14.400 ;
        RECT 3.900 13.200 6.300 14.100 ;
        RECT 3.900 12.900 5.100 13.200 ;
        RECT 10.800 9.900 12.000 11.100 ;
        RECT 10.800 9.300 11.700 9.900 ;
        RECT 3.300 8.700 4.500 9.000 ;
        RECT 0.600 7.800 4.500 8.700 ;
        RECT 5.400 8.100 7.800 9.300 ;
        RECT 10.500 8.100 11.700 9.300 ;
        RECT 12.600 8.700 13.800 9.000 ;
        RECT 12.600 7.800 16.200 8.700 ;
        RECT 0.600 1.800 1.800 7.800 ;
        RECT 15.000 1.800 16.200 7.800 ;
      LAYER via1 ;
        RECT 3.300 16.200 4.500 17.400 ;
        RECT 5.100 13.200 6.300 14.400 ;
        RECT 3.300 7.800 4.500 9.000 ;
      LAYER metal2 ;
        RECT 3.300 16.200 4.500 17.400 ;
        RECT 12.600 16.200 13.800 17.400 ;
        RECT 3.300 9.000 4.200 16.200 ;
        RECT 5.100 13.200 6.300 14.400 ;
        RECT 5.400 11.100 6.300 13.200 ;
        RECT 12.900 11.100 13.800 16.200 ;
        RECT 5.400 10.200 13.800 11.100 ;
        RECT 5.400 9.000 6.600 9.300 ;
        RECT 10.500 9.000 11.700 9.300 ;
        RECT 12.900 9.000 13.800 10.200 ;
        RECT 3.300 8.100 11.700 9.000 ;
        RECT 3.300 7.800 4.500 8.100 ;
        RECT 12.600 7.800 13.800 9.000 ;
  END
END XOR2X1
MACRO TBUFX2
  CLASS BLOCK ;
  FOREIGN TBUFX2 ;
  ORIGIN 1.500 0.900 ;
  SIZE 19.500 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 21.600000 ;
    PORT
      LAYER metal1 ;
        RECT 13.500 9.900 16.200 11.100 ;
    END
  END A
  PIN EN
    ANTENNAGATEAREA 18.000000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 12.900 1.800 15.300 ;
        RECT 0.600 9.900 1.500 12.900 ;
        RECT 0.600 8.700 2.100 9.900 ;
    END
  END EN
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 7.800 16.200 9.000 26.400 ;
        RECT 7.800 14.100 8.700 16.200 ;
        RECT 7.800 12.900 9.000 14.100 ;
        RECT 7.800 7.800 8.700 12.900 ;
        RECT 7.800 3.600 9.000 7.800 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 17.400 30.900 ;
        RECT 0.600 16.200 1.800 29.100 ;
        RECT 12.600 18.300 13.800 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 0.900 1.800 7.800 ;
        RECT 12.600 0.900 13.800 6.900 ;
        RECT -0.600 -0.900 17.400 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 3.000 16.200 4.200 28.200 ;
        RECT 5.400 27.300 11.400 28.200 ;
        RECT 5.400 16.200 6.600 27.300 ;
        RECT 10.200 17.400 11.400 27.300 ;
        RECT 15.000 17.400 16.200 28.200 ;
        RECT 10.200 16.200 16.200 17.400 ;
        RECT 3.000 13.500 3.900 16.200 ;
        RECT 3.000 12.300 4.200 13.500 ;
        RECT 3.000 7.800 3.900 12.300 ;
        RECT 10.200 7.800 16.200 8.700 ;
        RECT 3.000 1.800 4.200 7.800 ;
        RECT 5.400 2.700 6.600 7.800 ;
        RECT 10.200 2.700 11.400 7.800 ;
        RECT 15.300 6.900 16.200 7.800 ;
        RECT 5.400 1.800 11.400 2.700 ;
        RECT 15.000 1.800 16.200 6.900 ;
  END
END TBUFX2
MACRO TBUFX1
  CLASS BLOCK ;
  FOREIGN TBUFX1 ;
  ORIGIN 1.500 0.900 ;
  SIZE 14.100 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 10.800000 ;
    PORT
      LAYER metal1 ;
        RECT 9.000 9.900 11.400 11.100 ;
    END
  END A
  PIN EN
    ANTENNAGATEAREA 9.000000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 18.900 3.000 20.100 ;
    END
  END EN
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 5.700 16.200 6.900 28.200 ;
        RECT 6.000 14.100 6.900 16.200 ;
        RECT 5.400 12.900 6.900 14.100 ;
        RECT 6.000 7.800 6.900 12.900 ;
        RECT 5.700 1.800 6.900 7.800 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 12.600 30.900 ;
        RECT 0.600 22.200 1.800 29.100 ;
        RECT 9.600 16.200 10.800 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 0.900 1.800 4.800 ;
        RECT 9.600 0.900 10.800 7.800 ;
        RECT -0.600 -0.900 12.600 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 3.000 23.100 4.200 28.200 ;
        RECT 3.000 22.200 4.800 23.100 ;
        RECT 3.900 15.900 4.800 22.200 ;
        RECT 3.600 15.000 4.800 15.900 ;
        RECT 3.600 12.000 4.500 15.000 ;
        RECT 3.600 11.100 4.800 12.000 ;
        RECT 3.900 9.900 5.100 11.100 ;
        RECT 3.900 4.800 4.800 9.900 ;
        RECT 3.000 3.600 4.800 4.800 ;
        RECT 3.000 1.800 4.200 3.600 ;
  END
END TBUFX1
MACRO OR2X2
  CLASS BLOCK ;
  FOREIGN OR2X2 ;
  ORIGIN 2.100 0.900 ;
  SIZE 12.600 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 9.000000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 5.700 1.800 8.100 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 9.000000 ;
    PORT
      LAYER metal1 ;
        RECT 3.600 11.100 4.800 12.300 ;
        RECT 3.000 9.900 4.500 11.100 ;
    END
  END B
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 6.900 17.100 8.100 28.200 ;
        RECT 6.900 16.200 9.000 17.100 ;
        RECT 8.100 14.100 9.000 16.200 ;
        RECT 7.800 12.900 9.000 14.100 ;
        RECT 8.100 7.800 9.000 12.900 ;
        RECT 7.800 1.800 9.000 7.800 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 10.200 30.900 ;
        RECT 4.500 16.200 5.700 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 0.900 1.800 4.800 ;
        RECT 5.400 0.900 6.600 7.200 ;
        RECT -0.600 -0.900 10.200 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 15.300 1.800 28.200 ;
        RECT 0.600 14.700 6.600 15.300 ;
        RECT 0.600 14.400 6.900 14.700 ;
        RECT 5.700 13.500 6.900 14.400 ;
        RECT 6.000 9.000 6.900 13.500 ;
        RECT 3.300 8.100 6.900 9.000 ;
        RECT 3.300 4.800 4.200 8.100 ;
        RECT 3.000 1.800 4.200 4.800 ;
  END
END OR2X2
MACRO OR2X1
  CLASS BLOCK ;
  FOREIGN OR2X1 ;
  ORIGIN 2.400 0.900 ;
  SIZE 14.400 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 9.000000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 5.700 1.800 8.100 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 9.000000 ;
    PORT
      LAYER metal1 ;
        RECT 3.000 9.900 4.200 11.100 ;
        RECT 3.300 8.700 5.400 9.900 ;
    END
  END B
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 6.900 22.200 8.100 28.200 ;
        RECT 7.200 21.300 9.000 22.200 ;
        RECT 8.100 14.100 9.000 21.300 ;
        RECT 7.800 12.900 9.000 14.100 ;
        RECT 8.100 4.800 9.000 12.900 ;
        RECT 7.800 1.800 9.000 4.800 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 10.200 30.900 ;
        RECT 4.500 16.200 5.700 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 0.900 1.800 4.800 ;
        RECT 5.400 0.900 6.600 4.800 ;
        RECT -0.600 -0.900 10.200 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 15.300 1.800 28.200 ;
        RECT 0.600 14.400 6.900 15.300 ;
        RECT 5.700 14.100 6.900 14.400 ;
        RECT 5.700 11.700 6.600 14.100 ;
        RECT 5.700 10.800 7.200 11.700 ;
        RECT 6.300 7.200 7.200 10.800 ;
        RECT 3.300 6.300 7.200 7.200 ;
        RECT 3.300 4.800 4.200 6.300 ;
        RECT 3.000 1.800 4.200 4.800 ;
  END
END OR2X1
MACRO OAI22X1
  CLASS BLOCK ;
  FOREIGN OAI22X1 ;
  ORIGIN 2.400 0.900 ;
  SIZE 16.200 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 10.800000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 10.800 1.800 11.100 ;
        RECT 0.600 9.900 3.000 10.800 ;
        RECT 1.800 9.300 3.000 9.900 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 10.800000 ;
    PORT
      LAYER metal1 ;
        RECT 3.000 11.700 4.200 14.100 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 10.800000 ;
    PORT
      LAYER metal1 ;
        RECT 10.200 9.900 11.400 12.300 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA 10.800000 ;
    PORT
      LAYER metal1 ;
        RECT 7.800 11.700 9.000 14.100 ;
    END
  END D
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 4.500 16.200 7.500 28.200 ;
        RECT 5.400 11.100 6.300 16.200 ;
        RECT 5.400 10.800 6.600 11.100 ;
        RECT 5.400 9.900 9.000 10.800 ;
        RECT 8.100 7.800 9.000 9.900 ;
        RECT 7.800 3.600 9.000 7.800 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 12.600 30.900 ;
        RECT 0.600 16.200 1.800 29.100 ;
        RECT 10.200 16.200 11.400 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 3.000 0.900 4.200 6.600 ;
        RECT -0.600 -0.900 12.600 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.900 7.800 6.300 8.400 ;
        RECT 0.600 7.500 6.600 7.800 ;
        RECT 0.600 1.800 1.800 7.500 ;
        RECT 5.400 2.700 6.600 7.500 ;
        RECT 10.200 2.700 11.400 7.800 ;
        RECT 5.400 1.800 11.400 2.700 ;
  END
END OAI22X1
MACRO OAI21X1
  CLASS BLOCK ;
  FOREIGN OAI21X1 ;
  ORIGIN 2.400 0.900 ;
  SIZE 12.600 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 10.800000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 10.800 1.800 11.100 ;
        RECT 0.600 9.900 3.000 10.800 ;
        RECT 1.800 9.300 3.000 9.900 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 10.800000 ;
    PORT
      LAYER metal1 ;
        RECT 3.000 11.700 4.200 14.100 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 7.200000 ;
    PORT
      LAYER metal1 ;
        RECT 6.600 18.900 7.800 20.100 ;
        RECT 6.900 17.100 7.800 18.900 ;
        RECT 6.900 16.200 9.000 17.100 ;
        RECT 7.800 15.900 9.000 16.200 ;
    END
  END C
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 4.500 17.100 5.700 28.200 ;
        RECT 4.500 16.200 6.000 17.100 ;
        RECT 5.100 11.100 6.000 16.200 ;
        RECT 5.100 9.900 9.000 11.100 ;
        RECT 7.800 7.800 8.700 9.900 ;
        RECT 7.800 1.800 9.000 7.800 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 10.200 30.900 ;
        RECT 0.600 16.200 1.800 29.100 ;
        RECT 6.900 22.200 8.100 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 3.000 0.900 4.200 6.600 ;
        RECT -0.600 -0.900 10.200 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.900 7.800 6.300 8.400 ;
        RECT 0.600 7.500 6.600 7.800 ;
        RECT 0.600 1.800 1.800 7.500 ;
        RECT 5.400 1.800 6.600 7.500 ;
  END
END OAI21X1
MACRO NOR2X1
  CLASS BLOCK ;
  FOREIGN NOR2X1 ;
  ORIGIN 2.400 0.900 ;
  SIZE 12.000 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 9.000000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 5.700 1.800 8.100 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 9.000000 ;
    PORT
      LAYER metal1 ;
        RECT 5.400 12.900 6.600 15.300 ;
    END
  END B
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 4.500 17.400 5.700 28.200 ;
        RECT 3.000 16.200 5.700 17.400 ;
        RECT 3.300 11.100 4.200 16.200 ;
        RECT 3.000 9.900 4.200 11.100 ;
        RECT 3.300 4.800 4.200 9.900 ;
        RECT 3.000 1.800 4.200 4.800 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 7.800 30.900 ;
        RECT 0.600 16.200 1.800 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 0.900 1.800 4.800 ;
        RECT 5.400 0.900 6.600 4.800 ;
        RECT -0.600 -0.900 7.800 0.900 ;
    END
  END gnd
END NOR2X1
MACRO NAND3X1
  CLASS BLOCK ;
  FOREIGN NAND3X1 ;
  ORIGIN 2.400 0.900 ;
  SIZE 14.400 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 9.000000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 14.700 1.800 17.100 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 9.000000 ;
    PORT
      LAYER metal1 ;
        RECT 3.000 12.900 5.400 14.100 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 9.000000 ;
    PORT
      LAYER metal1 ;
        RECT 5.400 17.700 6.600 20.100 ;
    END
  END C
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 3.000 22.200 4.200 28.200 ;
        RECT 3.300 21.900 4.200 22.200 ;
        RECT 7.800 22.200 9.000 28.200 ;
        RECT 7.800 21.900 8.700 22.200 ;
        RECT 3.300 21.000 8.700 21.900 ;
        RECT 7.800 17.100 8.700 21.000 ;
        RECT 7.800 15.900 9.000 17.100 ;
        RECT 7.800 11.100 8.700 15.900 ;
        RECT 6.300 10.800 8.700 11.100 ;
        RECT 6.000 10.200 8.700 10.800 ;
        RECT 6.000 1.800 7.200 10.200 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 10.200 30.900 ;
        RECT 0.600 22.200 1.800 29.100 ;
        RECT 5.400 22.800 6.600 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 0.900 1.800 10.800 ;
        RECT -0.600 -0.900 10.200 0.900 ;
    END
  END gnd
END NAND3X1
MACRO NAND2X1
  CLASS BLOCK ;
  FOREIGN NAND2X1 ;
  ORIGIN 2.400 0.900 ;
  SIZE 12.000 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 7.200000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 8.700 1.800 11.100 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 7.200000 ;
    PORT
      LAYER metal1 ;
        RECT 5.400 15.900 6.600 18.300 ;
    END
  END B
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 3.000 7.800 4.200 28.200 ;
        RECT 3.000 6.900 5.700 7.800 ;
        RECT 4.500 1.800 5.700 6.900 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 7.800 30.900 ;
        RECT 0.600 22.200 1.800 29.100 ;
        RECT 5.400 22.200 6.600 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 0.900 1.800 7.800 ;
        RECT -0.600 -0.900 7.800 0.900 ;
    END
  END gnd
END NAND2X1
MACRO XNOR2X1
  CLASS BLOCK ;
  FOREIGN XNOR2X1 ;
  ORIGIN 2.400 0.900 ;
  SIZE 21.600 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 21.600000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 10.800 3.000 11.100 ;
        RECT 0.600 9.900 5.700 10.800 ;
        RECT 4.800 9.300 5.700 9.900 ;
        RECT 10.800 9.900 12.000 11.100 ;
        RECT 10.800 9.300 11.700 9.900 ;
        RECT 4.800 8.400 7.800 9.300 ;
        RECT 5.400 8.100 7.800 8.400 ;
        RECT 10.500 8.100 11.700 9.300 ;
      LAYER metal2 ;
        RECT 5.400 9.000 6.600 9.300 ;
        RECT 10.500 9.000 11.700 9.300 ;
        RECT 5.400 8.100 11.700 9.000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 21.600000 ;
    PORT
      LAYER metal1 ;
        RECT 13.800 9.900 16.200 11.100 ;
    END
  END B
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 7.200 17.100 9.600 28.200 ;
        RECT 7.200 16.200 10.200 17.100 ;
        RECT 9.300 14.100 10.200 16.200 ;
        RECT 9.300 13.200 11.400 14.100 ;
        RECT 8.700 12.900 11.400 13.200 ;
        RECT 8.700 12.300 10.200 12.900 ;
        RECT 8.700 7.200 9.600 12.300 ;
        RECT 7.200 1.800 9.600 7.200 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 17.400 30.900 ;
        RECT 3.300 28.200 4.500 29.100 ;
        RECT 3.000 18.300 4.500 28.200 ;
        RECT 12.300 18.300 13.800 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 3.000 1.800 4.500 6.900 ;
        RECT 3.300 0.900 4.500 1.800 ;
        RECT 12.300 0.900 13.800 6.900 ;
        RECT -0.600 -0.900 17.400 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 17.100 1.800 28.200 ;
        RECT 2.700 17.100 3.900 17.400 ;
        RECT 0.600 16.200 3.900 17.100 ;
        RECT 12.600 17.100 13.800 17.400 ;
        RECT 15.000 17.100 16.200 28.200 ;
        RECT 12.600 16.200 16.200 17.100 ;
        RECT 3.000 15.300 3.900 16.200 ;
        RECT 3.000 14.400 8.100 15.300 ;
        RECT 6.900 14.100 8.100 14.400 ;
        RECT 3.600 13.200 4.800 13.500 ;
        RECT 3.600 12.300 7.500 13.200 ;
        RECT 6.600 11.400 7.500 12.300 ;
        RECT 6.600 10.200 7.800 11.400 ;
        RECT 2.700 8.700 3.900 9.000 ;
        RECT 0.600 7.800 3.900 8.700 ;
        RECT 12.600 8.700 13.800 9.000 ;
        RECT 12.600 7.800 16.200 8.700 ;
        RECT 0.600 1.800 1.800 7.800 ;
        RECT 15.000 1.800 16.200 7.800 ;
      LAYER via1 ;
        RECT 2.700 16.200 3.900 17.400 ;
        RECT 2.700 7.800 3.900 9.000 ;
      LAYER metal2 ;
        RECT 2.700 16.200 3.900 17.400 ;
        RECT 12.600 16.200 13.800 17.400 ;
        RECT 2.700 9.000 3.600 16.200 ;
        RECT 6.600 11.100 7.800 11.400 ;
        RECT 12.900 11.100 13.800 16.200 ;
        RECT 6.600 10.200 13.800 11.100 ;
        RECT 12.900 9.000 13.800 10.200 ;
        RECT 2.700 7.800 3.900 9.000 ;
        RECT 12.600 7.800 13.800 9.000 ;
  END
END XNOR2X1
MACRO LATCH
  CLASS BLOCK ;
  FOREIGN LATCH ;
  ORIGIN 2.400 0.900 ;
  SIZE 21.600 BY 32.400 ;
  PIN D
    ANTENNAGATEAREA 5.400000 ;
    PORT
      LAYER metal1 ;
        RECT 5.400 15.300 6.600 17.100 ;
        RECT 3.900 14.100 6.600 15.300 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 14.400001 ;
    PORT
      LAYER metal1 ;
        RECT 1.800 10.800 4.200 11.100 ;
        RECT 8.700 10.800 9.900 12.300 ;
        RECT 1.800 9.900 9.900 10.800 ;
        RECT 6.600 6.900 7.800 9.900 ;
    END
  END CLK
  PIN Q
    ANTENNAGATEAREA 3.600000 ;
    PORT
      LAYER metal1 ;
        RECT 15.000 12.600 16.200 28.200 ;
        RECT 11.100 11.400 16.200 12.600 ;
        RECT 15.000 1.800 16.200 11.400 ;
    END
  END Q
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 17.400 30.900 ;
        RECT 3.000 16.200 4.200 29.100 ;
        RECT 12.600 16.200 13.800 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 3.000 0.900 4.200 7.800 ;
        RECT 12.600 0.900 13.800 7.800 ;
        RECT -0.600 -0.900 17.400 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 14.700 1.800 28.200 ;
        RECT 7.500 22.200 9.300 28.200 ;
        RECT 7.800 21.000 9.000 22.200 ;
        RECT 7.800 14.100 14.100 15.300 ;
        RECT 0.600 12.900 1.800 13.200 ;
        RECT 6.300 12.900 7.500 13.200 ;
        RECT 0.600 12.000 7.500 12.900 ;
        RECT 0.600 1.800 1.800 9.000 ;
        RECT 7.800 4.800 9.000 6.000 ;
        RECT 7.500 1.800 9.300 4.800 ;
      LAYER via1 ;
        RECT 0.600 15.000 1.800 16.200 ;
        RECT 0.600 7.800 1.800 9.000 ;
      LAYER metal2 ;
        RECT 0.600 7.800 1.800 16.200 ;
        RECT 7.800 4.800 9.000 22.200 ;
  END
END LATCH
MACRO DFFSR
  CLASS BLOCK ;
  FOREIGN DFFSR ;
  ORIGIN 2.400 0.900 ;
  SIZE 57.600 BY 32.400 ;
  PIN D
    ANTENNAGATEAREA 5.400000 ;
    PORT
      LAYER metal1 ;
        RECT 19.800 8.700 21.000 11.100 ;
    END
  END D
  PIN S
    ANTENNAGATEAREA 14.400001 ;
    PORT
      LAYER metal1 ;
        RECT 5.400 16.200 6.600 17.100 ;
        RECT 10.500 16.200 11.700 16.500 ;
        RECT 5.400 15.300 45.900 16.200 ;
        RECT 44.700 15.000 45.900 15.300 ;
    END
  END S
  PIN R
    ANTENNAGATEAREA 14.400001 ;
    PORT
      LAYER metal1 ;
        RECT 2.700 13.500 37.800 14.400 ;
        RECT 2.700 13.200 3.900 13.500 ;
        RECT 10.200 12.900 11.400 13.500 ;
        RECT 36.600 12.600 37.800 13.500 ;
    END
  END R
  PIN CLK
    ANTENNAGATEAREA 5.400000 ;
    PORT
      LAYER metal1 ;
        RECT 24.600 6.900 27.000 8.100 ;
    END
  END CLK
  PIN Q
    PORT
      LAYER metal1 ;
        RECT 48.600 16.500 49.800 28.200 ;
        RECT 48.600 15.300 50.100 16.500 ;
        RECT 48.900 8.700 50.100 15.300 ;
        RECT 48.600 7.500 50.100 8.700 ;
        RECT 48.600 1.800 49.800 7.500 ;
    END
  END Q
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 53.400 30.900 ;
        RECT 0.600 22.200 1.800 29.100 ;
        RECT 5.400 22.200 6.600 29.100 ;
        RECT 10.200 22.200 11.400 29.100 ;
        RECT 19.800 22.200 21.000 29.100 ;
        RECT 24.600 22.200 25.800 29.100 ;
        RECT 36.600 22.200 37.800 29.100 ;
        RECT 41.400 22.200 42.600 29.100 ;
        RECT 46.200 22.200 47.400 29.100 ;
        RECT 51.000 22.200 52.200 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 5.400 0.900 6.600 7.800 ;
        RECT 19.800 0.900 21.000 4.800 ;
        RECT 24.600 0.900 25.800 4.800 ;
        RECT 41.400 0.900 42.600 7.800 ;
        RECT 51.000 0.900 52.200 4.800 ;
        RECT -0.600 -0.900 53.400 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 3.000 23.100 4.200 28.200 ;
        RECT 2.700 22.200 4.200 23.100 ;
        RECT 2.700 21.300 3.600 22.200 ;
        RECT 7.800 21.300 9.000 28.200 ;
        RECT 12.600 24.000 13.800 28.200 ;
        RECT 15.000 24.000 16.200 28.200 ;
        RECT 0.600 20.400 3.600 21.300 ;
        RECT 0.600 12.000 1.800 20.400 ;
        RECT 4.500 20.100 10.800 21.300 ;
        RECT 17.400 21.000 18.600 28.200 ;
        RECT 22.200 21.000 23.400 28.200 ;
        RECT 4.500 19.500 5.400 20.100 ;
        RECT 3.000 18.300 5.400 19.500 ;
        RECT 9.900 19.200 18.600 20.100 ;
        RECT 6.900 18.300 9.000 19.200 ;
        RECT 6.900 18.000 16.200 18.300 ;
        RECT 8.100 17.400 16.200 18.000 ;
        RECT 15.000 17.100 16.200 17.400 ;
        RECT 17.700 18.000 18.600 19.200 ;
        RECT 19.500 18.900 23.400 20.100 ;
        RECT 27.000 18.900 28.200 28.200 ;
        RECT 29.400 24.000 30.600 28.200 ;
        RECT 31.800 24.000 33.000 28.200 ;
        RECT 34.200 24.000 35.400 28.200 ;
        RECT 31.800 20.100 38.100 21.300 ;
        RECT 39.000 20.100 40.200 28.200 ;
        RECT 43.800 21.300 45.000 28.200 ;
        RECT 43.800 20.400 47.700 21.300 ;
        RECT 39.000 18.900 42.900 20.100 ;
        RECT 29.400 18.000 30.600 18.300 ;
        RECT 17.700 17.100 30.600 18.000 ;
        RECT 34.200 18.000 35.400 18.300 ;
        RECT 46.800 18.000 47.700 20.400 ;
        RECT 34.200 17.100 47.700 18.000 ;
        RECT 46.800 14.400 47.700 17.100 ;
        RECT 46.800 13.500 48.000 14.400 ;
        RECT 0.600 10.800 13.800 12.000 ;
        RECT 14.700 11.400 17.700 12.600 ;
        RECT 23.400 11.400 28.200 12.600 ;
        RECT 0.600 1.800 1.800 10.800 ;
        RECT 4.200 8.700 8.700 9.900 ;
        RECT 7.500 7.800 8.700 8.700 ;
        RECT 16.500 7.800 17.700 11.400 ;
        RECT 27.600 10.200 28.800 10.500 ;
        RECT 22.200 9.300 28.800 10.200 ;
        RECT 22.200 9.000 23.400 9.300 ;
        RECT 31.800 8.100 33.000 12.300 ;
        RECT 40.500 11.400 46.200 12.600 ;
        RECT 40.500 9.600 41.700 11.400 ;
        RECT 47.100 10.500 48.000 13.500 ;
        RECT 22.200 7.800 23.400 8.100 ;
        RECT 7.500 6.600 11.400 7.800 ;
        RECT 16.500 6.900 23.400 7.800 ;
        RECT 31.500 6.900 33.000 8.100 ;
        RECT 39.000 8.700 41.700 9.600 ;
        RECT 46.200 9.600 48.000 10.500 ;
        RECT 39.000 7.800 40.200 8.700 ;
        RECT 10.200 1.800 11.400 6.600 ;
        RECT 36.600 6.600 40.200 7.800 ;
        RECT 12.600 1.800 13.800 6.000 ;
        RECT 15.000 1.800 16.200 6.000 ;
        RECT 17.400 1.800 18.600 6.000 ;
        RECT 22.200 1.800 23.400 6.000 ;
        RECT 27.000 1.800 28.200 6.000 ;
        RECT 29.400 1.800 30.600 6.000 ;
        RECT 31.800 1.800 33.000 6.000 ;
        RECT 34.200 1.800 35.400 6.000 ;
        RECT 36.600 1.800 37.800 6.600 ;
        RECT 46.200 1.800 47.400 9.600 ;
      LAYER via1 ;
        RECT 27.000 21.000 28.200 22.200 ;
        RECT 22.200 18.900 23.400 20.100 ;
        RECT 29.400 17.100 30.600 18.300 ;
        RECT 12.600 10.800 13.800 12.000 ;
        RECT 27.000 11.400 28.200 12.600 ;
        RECT 12.600 4.800 13.800 6.000 ;
        RECT 15.000 4.800 16.200 6.000 ;
        RECT 17.400 4.800 18.600 6.000 ;
        RECT 22.200 4.800 23.400 6.000 ;
        RECT 27.000 4.800 28.200 6.000 ;
        RECT 29.400 4.800 30.600 6.000 ;
        RECT 31.800 4.800 33.000 6.000 ;
        RECT 34.200 4.800 35.400 6.000 ;
      LAYER metal2 ;
        RECT 12.600 4.800 13.800 25.200 ;
        RECT 15.000 4.800 16.200 25.200 ;
        RECT 17.400 4.800 18.600 22.200 ;
        RECT 22.200 4.800 23.400 22.200 ;
        RECT 27.000 4.800 28.200 22.200 ;
        RECT 29.400 4.800 30.600 25.200 ;
        RECT 31.800 4.800 33.000 25.200 ;
        RECT 34.200 4.800 35.400 25.200 ;
  END
END DFFSR
MACRO CLKBUF3
  CLASS BLOCK ;
  FOREIGN CLKBUF3 ;
  ORIGIN 2.400 0.900 ;
  SIZE 45.600 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 21.600000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 10.800 3.300 12.000 ;
        RECT 0.600 9.900 1.800 10.800 ;
    END
  END A
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 36.600 15.300 37.800 28.200 ;
        RECT 36.600 14.100 40.200 15.300 ;
        RECT 39.000 9.900 40.200 14.100 ;
        RECT 36.600 8.700 40.200 9.900 ;
        RECT 36.600 1.800 37.800 8.700 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 41.400 30.900 ;
        RECT 0.600 16.200 1.800 29.100 ;
        RECT 5.400 16.200 6.600 29.100 ;
        RECT 10.200 16.200 11.400 29.100 ;
        RECT 15.000 16.200 16.200 29.100 ;
        RECT 19.800 16.200 21.000 29.100 ;
        RECT 24.600 16.200 25.800 29.100 ;
        RECT 29.400 16.200 30.600 29.100 ;
        RECT 34.200 16.200 35.400 29.100 ;
        RECT 39.000 16.200 40.200 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 0.900 1.800 7.800 ;
        RECT 5.400 0.900 6.600 7.800 ;
        RECT 10.200 0.900 11.400 7.800 ;
        RECT 15.000 0.900 16.200 7.800 ;
        RECT 19.800 0.900 21.000 7.800 ;
        RECT 24.600 0.900 25.800 7.800 ;
        RECT 29.400 0.900 30.600 7.800 ;
        RECT 34.200 0.900 35.400 7.800 ;
        RECT 39.000 0.900 40.200 7.800 ;
        RECT -0.600 -0.900 41.400 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 3.000 15.300 4.200 28.200 ;
        RECT 7.800 15.300 9.000 28.200 ;
        RECT 12.600 15.300 13.800 28.200 ;
        RECT 17.400 15.300 18.600 28.200 ;
        RECT 22.200 15.300 23.400 28.200 ;
        RECT 27.000 15.300 28.200 28.200 ;
        RECT 31.800 15.300 33.000 28.200 ;
        RECT 3.000 14.100 5.700 15.300 ;
        RECT 7.800 14.100 11.100 15.300 ;
        RECT 12.600 14.100 15.900 15.300 ;
        RECT 17.400 14.100 21.000 15.300 ;
        RECT 22.200 14.100 24.900 15.300 ;
        RECT 27.000 14.100 30.300 15.300 ;
        RECT 31.800 14.100 35.100 15.300 ;
        RECT 4.500 12.000 5.700 14.100 ;
        RECT 9.900 12.000 11.100 14.100 ;
        RECT 14.700 12.000 15.900 14.100 ;
        RECT 19.800 12.000 21.000 14.100 ;
        RECT 23.700 12.000 24.900 14.100 ;
        RECT 29.100 12.000 30.300 14.100 ;
        RECT 33.900 12.000 35.100 14.100 ;
        RECT 4.500 10.800 8.400 12.000 ;
        RECT 9.900 10.800 13.500 12.000 ;
        RECT 14.700 10.800 18.600 12.000 ;
        RECT 19.800 10.800 22.500 12.000 ;
        RECT 23.700 10.800 27.600 12.000 ;
        RECT 29.100 10.800 32.700 12.000 ;
        RECT 33.900 10.800 37.800 12.000 ;
        RECT 4.500 9.900 5.700 10.800 ;
        RECT 9.900 9.900 11.100 10.800 ;
        RECT 14.700 9.900 15.900 10.800 ;
        RECT 19.800 9.900 21.000 10.800 ;
        RECT 23.700 9.900 24.900 10.800 ;
        RECT 29.100 9.900 30.300 10.800 ;
        RECT 33.900 9.900 35.100 10.800 ;
        RECT 3.000 8.700 5.700 9.900 ;
        RECT 7.800 8.700 11.100 9.900 ;
        RECT 12.600 8.700 15.900 9.900 ;
        RECT 17.400 8.700 21.000 9.900 ;
        RECT 22.200 8.700 24.900 9.900 ;
        RECT 27.000 8.700 30.300 9.900 ;
        RECT 31.800 8.700 35.100 9.900 ;
        RECT 3.000 1.800 4.200 8.700 ;
        RECT 7.800 1.800 9.000 8.700 ;
        RECT 12.600 1.800 13.800 8.700 ;
        RECT 17.400 1.800 18.600 8.700 ;
        RECT 22.200 1.800 23.400 8.700 ;
        RECT 27.000 1.800 28.200 8.700 ;
        RECT 31.800 1.800 33.000 8.700 ;
  END
END CLKBUF3
MACRO CLKBUF2
  CLASS BLOCK ;
  FOREIGN CLKBUF2 ;
  ORIGIN 2.400 0.900 ;
  SIZE 36.000 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 21.600000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 10.800 3.300 12.000 ;
        RECT 0.600 9.900 1.800 10.800 ;
    END
  END A
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 27.000 15.300 28.200 28.200 ;
        RECT 27.000 14.100 30.600 15.300 ;
        RECT 29.400 9.900 30.600 14.100 ;
        RECT 27.000 8.700 30.600 9.900 ;
        RECT 27.000 1.800 28.200 8.700 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 31.800 30.900 ;
        RECT 0.600 16.200 1.800 29.100 ;
        RECT 5.400 16.200 6.600 29.100 ;
        RECT 10.200 16.200 11.400 29.100 ;
        RECT 15.000 16.200 16.200 29.100 ;
        RECT 19.800 16.200 21.000 29.100 ;
        RECT 24.600 16.200 25.800 29.100 ;
        RECT 29.400 16.200 30.600 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 0.900 1.800 7.800 ;
        RECT 5.400 0.900 6.600 7.800 ;
        RECT 10.200 0.900 11.400 7.800 ;
        RECT 15.000 0.900 16.200 7.800 ;
        RECT 19.800 0.900 21.000 7.800 ;
        RECT 24.600 0.900 25.800 7.800 ;
        RECT 29.400 0.900 30.600 7.800 ;
        RECT -0.600 -0.900 31.800 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 3.000 15.300 4.200 28.200 ;
        RECT 7.800 15.300 9.000 28.200 ;
        RECT 12.600 15.300 13.800 28.200 ;
        RECT 17.400 15.300 18.600 28.200 ;
        RECT 22.200 15.300 23.400 28.200 ;
        RECT 3.000 14.100 5.700 15.300 ;
        RECT 7.800 14.100 11.100 15.300 ;
        RECT 12.600 14.100 15.900 15.300 ;
        RECT 17.400 14.100 21.000 15.300 ;
        RECT 22.200 14.100 24.900 15.300 ;
        RECT 4.500 12.000 5.700 14.100 ;
        RECT 9.900 12.000 11.100 14.100 ;
        RECT 14.700 12.000 15.900 14.100 ;
        RECT 19.800 12.000 21.000 14.100 ;
        RECT 23.700 12.000 24.900 14.100 ;
        RECT 4.500 10.800 8.400 12.000 ;
        RECT 9.900 10.800 13.500 12.000 ;
        RECT 14.700 10.800 18.600 12.000 ;
        RECT 19.800 10.800 22.500 12.000 ;
        RECT 23.700 10.800 27.600 12.000 ;
        RECT 4.500 9.900 5.700 10.800 ;
        RECT 9.900 9.900 11.100 10.800 ;
        RECT 14.700 9.900 15.900 10.800 ;
        RECT 19.800 9.900 21.000 10.800 ;
        RECT 23.700 9.900 24.900 10.800 ;
        RECT 3.000 8.700 5.700 9.900 ;
        RECT 7.800 8.700 11.100 9.900 ;
        RECT 12.600 8.700 15.900 9.900 ;
        RECT 17.400 8.700 21.000 9.900 ;
        RECT 22.200 8.700 24.900 9.900 ;
        RECT 3.000 1.800 4.200 8.700 ;
        RECT 7.800 1.800 9.000 8.700 ;
        RECT 12.600 1.800 13.800 8.700 ;
        RECT 17.400 1.800 18.600 8.700 ;
        RECT 22.200 1.800 23.400 8.700 ;
  END
END CLKBUF2
MACRO CLKBUF1
  CLASS BLOCK ;
  FOREIGN CLKBUF1 ;
  ORIGIN 2.400 0.900 ;
  SIZE 26.400 BY 32.400 ;
  PIN A
    ANTENNAGATEAREA 21.600000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 10.800 3.300 12.000 ;
        RECT 0.600 9.900 1.800 10.800 ;
    END
  END A
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 17.400 15.300 18.600 28.200 ;
        RECT 17.400 14.100 21.000 15.300 ;
        RECT 19.800 9.900 21.000 14.100 ;
        RECT 17.400 8.700 21.000 9.900 ;
        RECT 17.400 1.800 18.600 8.700 ;
    END
  END Y
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.600 29.100 22.200 30.900 ;
        RECT 0.600 16.200 1.800 29.100 ;
        RECT 5.400 16.200 6.600 29.100 ;
        RECT 10.200 16.200 11.400 29.100 ;
        RECT 15.000 16.200 16.200 29.100 ;
        RECT 19.800 16.200 21.000 29.100 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 0.900 1.800 7.800 ;
        RECT 5.400 0.900 6.600 7.800 ;
        RECT 10.200 0.900 11.400 7.800 ;
        RECT 15.000 0.900 16.200 7.800 ;
        RECT 19.800 0.900 21.000 7.800 ;
        RECT -0.600 -0.900 22.200 0.900 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 3.000 15.300 4.200 28.200 ;
        RECT 7.800 15.300 9.000 28.200 ;
        RECT 12.600 15.300 13.800 28.200 ;
        RECT 3.000 14.100 5.700 15.300 ;
        RECT 7.800 14.100 11.100 15.300 ;
        RECT 12.600 14.100 15.900 15.300 ;
        RECT 4.500 12.000 5.700 14.100 ;
        RECT 9.900 12.000 11.100 14.100 ;
        RECT 14.700 12.000 15.900 14.100 ;
        RECT 4.500 10.800 8.400 12.000 ;
        RECT 9.900 10.800 13.500 12.000 ;
        RECT 14.700 10.800 18.600 12.000 ;
        RECT 4.500 9.900 5.700 10.800 ;
        RECT 9.900 9.900 11.100 10.800 ;
        RECT 14.700 9.900 15.900 10.800 ;
        RECT 3.000 8.700 5.700 9.900 ;
        RECT 7.800 8.700 11.100 9.900 ;
        RECT 12.600 8.700 15.900 9.900 ;
        RECT 3.000 1.800 4.200 8.700 ;
        RECT 7.800 1.800 9.000 8.700 ;
        RECT 12.600 1.800 13.800 8.700 ;
  END
END CLKBUF1
END LIBRARY

