** sch_path: /home/goodkook/ETRI050_DesignKit/Tutorials/1-4_StdCell_DFFSR/Sch/NAND2X1.sch
**.subckt NAND2X1 B A Y vdd gnd
*.ipin A
*.ipin B
*.opin Y
*.iopin vdd
*.iopin gnd
M1 Y A net1 GND nfet w=6u l=0.6u m=1
M2 Y A vdd VDD pfet w=6u l=0.6u m=1
M3 net1 B gnd GND nfet w=6u l=0.6u m=1
M4 Y B vdd VDD pfet w=6u l=0.6u m=1
**.ends
.end
