magic
tech scmos
magscale 1 2
timestamp 1702310384
<< nwell >>
rect -12 154 273 272
<< ntransistor >>
rect 18 14 22 54
rect 38 14 42 54
rect 58 14 62 54
rect 78 14 82 54
rect 98 14 102 54
rect 118 14 122 54
rect 138 14 142 54
rect 158 14 162 54
rect 178 14 182 54
rect 198 14 202 54
rect 218 14 222 54
rect 238 14 242 54
<< ptransistor >>
rect 18 166 22 246
rect 38 166 42 246
rect 58 166 62 246
rect 78 166 82 246
rect 98 166 102 246
rect 118 166 122 246
rect 138 166 142 246
rect 158 166 162 246
rect 178 166 182 246
rect 198 166 202 246
rect 218 166 222 246
rect 238 166 242 246
<< ndiffusion >>
rect 16 14 18 54
rect 22 14 24 54
rect 36 14 38 54
rect 42 14 44 54
rect 56 14 58 54
rect 62 14 64 54
rect 76 14 78 54
rect 82 14 84 54
rect 96 14 98 54
rect 102 14 104 54
rect 116 14 118 54
rect 122 14 124 54
rect 136 14 138 54
rect 142 14 144 54
rect 156 14 158 54
rect 162 14 164 54
rect 176 14 178 54
rect 182 14 184 54
rect 196 14 198 54
rect 202 14 204 54
rect 216 14 218 54
rect 222 14 224 54
rect 236 14 238 54
rect 242 14 244 54
<< pdiffusion >>
rect 16 166 18 246
rect 22 166 24 246
rect 36 166 38 246
rect 42 166 44 246
rect 56 166 58 246
rect 62 166 64 246
rect 76 166 78 246
rect 82 166 84 246
rect 96 166 98 246
rect 102 166 104 246
rect 116 166 118 246
rect 122 166 124 246
rect 136 166 138 246
rect 142 166 144 246
rect 156 166 158 246
rect 162 166 164 246
rect 176 166 178 246
rect 182 166 184 246
rect 196 166 198 246
rect 202 166 204 246
rect 216 166 218 246
rect 222 166 224 246
rect 236 166 238 246
rect 242 166 244 246
<< ndcontact >>
rect 4 14 16 54
rect 24 14 36 54
rect 44 14 56 54
rect 64 14 76 54
rect 84 14 96 54
rect 104 14 116 54
rect 124 14 136 54
rect 144 14 156 54
rect 164 14 176 54
rect 184 14 196 54
rect 204 14 216 54
rect 224 14 236 54
rect 244 14 256 54
<< pdcontact >>
rect 4 166 16 246
rect 24 166 36 246
rect 44 166 56 246
rect 64 166 76 246
rect 84 166 96 246
rect 104 166 116 246
rect 124 166 136 246
rect 144 166 156 246
rect 164 166 176 246
rect 184 166 196 246
rect 204 166 216 246
rect 224 166 236 246
rect 244 166 256 246
<< psubstratepcontact >>
rect -6 -6 266 6
<< nsubstratencontact >>
rect -6 254 266 266
<< polysilicon >>
rect 18 246 22 250
rect 38 246 42 250
rect 58 246 62 250
rect 78 246 82 250
rect 98 246 102 250
rect 118 246 122 250
rect 138 246 142 250
rect 158 246 162 250
rect 178 246 182 250
rect 198 246 202 250
rect 218 246 222 250
rect 238 246 242 250
rect 18 117 22 166
rect 38 117 42 166
rect 18 108 42 117
rect 18 54 22 108
rect 38 54 42 108
rect 58 122 62 166
rect 78 118 82 166
rect 70 110 82 118
rect 58 54 62 110
rect 78 54 82 110
rect 98 122 102 166
rect 118 118 122 166
rect 110 110 122 118
rect 98 54 102 110
rect 118 54 122 110
rect 138 122 142 166
rect 158 118 162 166
rect 150 110 162 118
rect 138 54 142 110
rect 158 54 162 110
rect 178 122 182 166
rect 198 118 202 166
rect 190 110 202 118
rect 178 54 182 110
rect 198 54 202 110
rect 218 122 222 166
rect 238 118 242 166
rect 230 110 242 118
rect 218 54 222 110
rect 238 54 242 110
rect 18 10 22 14
rect 38 10 42 14
rect 58 10 62 14
rect 78 10 82 14
rect 98 10 102 14
rect 118 10 122 14
rect 138 10 142 14
rect 158 10 162 14
rect 178 10 182 14
rect 198 10 202 14
rect 218 10 222 14
rect 238 10 242 14
<< polycontact >>
rect 6 105 18 117
rect 58 110 70 122
rect 98 110 110 122
rect 138 110 150 122
rect 178 110 190 122
rect 218 110 230 122
<< metal1 >>
rect -6 266 266 268
rect -6 252 266 254
rect 4 246 16 252
rect 44 246 56 252
rect 84 246 96 252
rect 124 246 136 252
rect 164 246 176 252
rect 204 246 216 252
rect 244 246 256 252
rect 24 160 36 166
rect 64 160 76 166
rect 104 160 116 166
rect 144 160 156 166
rect 184 160 196 166
rect 224 160 236 166
rect 24 152 46 160
rect 64 152 90 160
rect 104 152 130 160
rect 144 152 172 160
rect 184 152 206 160
rect 224 152 254 160
rect 3 123 17 137
rect 6 117 17 123
rect 38 118 46 152
rect 38 110 58 118
rect 82 118 90 152
rect 82 110 98 118
rect 122 118 130 152
rect 122 110 138 118
rect 164 118 172 152
rect 164 110 178 118
rect 198 118 206 152
rect 246 137 254 152
rect 243 123 257 137
rect 198 110 218 118
rect 38 68 46 110
rect 82 68 90 110
rect 122 68 130 110
rect 164 68 172 110
rect 198 68 206 110
rect 246 68 254 123
rect 24 60 46 68
rect 64 60 90 68
rect 104 60 130 68
rect 144 60 172 68
rect 184 60 206 68
rect 224 60 254 68
rect 24 54 36 60
rect 64 54 76 60
rect 104 54 116 60
rect 144 54 156 60
rect 184 54 196 60
rect 224 54 236 60
rect 4 8 16 14
rect 44 8 56 14
rect 84 8 96 14
rect 124 8 136 14
rect 164 8 176 14
rect 204 8 216 14
rect 244 8 256 14
rect -6 6 266 8
rect -6 -8 266 -6
<< m1p >>
rect -6 252 266 268
rect 3 123 17 137
rect 243 123 257 137
rect -6 -8 266 8
<< labels >>
rlabel nsubstratencontact 130 260 130 260 0 vdd
port 3 nsew power bidirectional abutment
rlabel psubstratepcontact 130 0 130 0 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 10 131 10 131 0 A
port 1 nsew signal input
rlabel metal1 250 131 250 131 0 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 260 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
