magic
tech scmos
magscale 1 30
timestamp 1756369954
<< checkpaint >>
rect 9150 9150 180850 180850
use IOFILLER18  IOFILLER18_6 ~/ETRI050_DesignKit/pads_ETRI
timestamp 1741148472
transform 1 0 73845 0 1 18900
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_7
timestamp 1741148472
transform 1 0 60345 0 1 18900
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_8
timestamp 1741148472
transform 1 0 100845 0 1 18900
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_9
timestamp 1741148472
transform 1 0 87345 0 1 18900
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_10
timestamp 1741148472
transform 1 0 127845 0 1 18900
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_11
timestamp 1741148472
transform 1 0 114345 0 1 18900
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_12
timestamp 1741148472
transform 0 1 18899 -1 0 75655
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_13
timestamp 1741148472
transform 0 1 18899 -1 0 62155
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_14
timestamp 1741148472
transform 0 1 18900 -1 0 102655
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_15
timestamp 1741148472
transform 0 1 18900 -1 0 89155
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_16
timestamp 1741148472
transform 1 0 73845 0 -1 171100
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_17
timestamp 1741148472
transform 0 1 18897 -1 0 116155
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_18
timestamp 1741148472
transform 0 1 18900 -1 0 129655
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_19
timestamp 1741148472
transform 1 0 60345 0 -1 171101
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_20
timestamp 1741148472
transform 1 0 100845 0 -1 171100
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_21
timestamp 1741148472
transform 1 0 87344 0 -1 171100
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_22
timestamp 1741148472
transform 1 0 127845 0 -1 171100
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_23
timestamp 1741148472
transform 1 0 114345 0 -1 171100
box 30 0 1770 25060
use IOFILLER50  IOFILLER50_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 43621 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_3
timestamp 1569139307
transform 1 0 43638 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_4
timestamp 1569139307
transform 0 1 18900 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_5
timestamp 1569139307
transform 0 1 18900 -1 0 146379
box -35 0 5035 25060
use PCORNER  PCORNER_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 18900 0 1 18900
box 0 0 25300 25300
use PCORNER  PCORNER_1
timestamp 1569139307
transform 1 0 18900 0 -1 171100
box 0 0 25300 25300
use PAD_80__0  PAD_80_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1740657577
transform 0 -1 176000 1 0 135500
box -4250 -4250 4250 4900
use PAD_80__0  PAD_80_1
timestamp 1740657577
transform 0 -1 176000 1 0 122000
box -4250 -4250 4250 4900
use PAD_80__0  PAD_80_2
timestamp 1740657577
transform 0 -1 176000 1 0 108500
box -4250 -4250 4250 4900
use PAD_80__0  PAD_80_3
timestamp 1740657577
transform 0 -1 176000 1 0 95000
box -4250 -4250 4250 4900
use PAD_80__0  PAD_80_4
timestamp 1740657577
transform 0 -1 176000 1 0 81500
box -4250 -4250 4250 4900
use PAD_80__0  PAD_80_5
timestamp 1740657577
transform 0 -1 176000 1 0 68000
box -4250 -4250 4250 4900
use PAD_80__0  PAD_80_6
timestamp 1740657577
transform 0 -1 176000 1 0 54500
box -4250 -4250 4250 4900
use PIC  CLK ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1756352440
transform 0 1 18900 -1 0 114500
box -100 -9150 12100 25300
use PIC  RST
timestamp 1756352440
transform 0 1 18900 -1 0 128000
box -100 -9150 12100 25300
use PIC  X_0
timestamp 1756352440
transform 1 0 75500 0 -1 171100
box -100 -9150 12100 25300
use PIC  X_1
timestamp 1756352440
transform 1 0 48500 0 -1 171100
box -100 -9150 12100 25300
use PIC  X_2
timestamp 1756352440
transform 1 0 116000 0 -1 171100
box -100 -9150 12100 25300
use PIC  X_3
timestamp 1756352440
transform 0 1 18900 -1 0 87500
box -100 -9150 12100 25300
use PIC  X_4
timestamp 1756352440
transform 1 0 89000 0 -1 171100
box -100 -9150 12100 25300
use PIC  X_5
timestamp 1756352440
transform 0 1 18900 -1 0 101000
box -100 -9150 12100 25300
use PIC  X_6
timestamp 1756352440
transform 1 0 62000 0 -1 171100
box -100 -9150 12100 25300
use PIC  X_7
timestamp 1756352440
transform 1 0 102500 0 -1 171100
box -100 -9150 12100 25300
use POB8  READY ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 0 1 18900 -1 0 141500
box -100 -9150 12100 25300
use POB8  Y_0
timestamp 1569139307
transform 1 0 89000 0 1 18900
box -100 -9150 12100 25300
use POB8  Y_1
timestamp 1569139307
transform 0 1 18900 -1 0 74000
box -100 -9150 12100 25300
use POB8  Y_2
timestamp 1569139307
transform 0 1 18900 -1 0 60500
box -100 -9150 12100 25300
use POB8  Y_3
timestamp 1569139307
transform 1 0 75500 0 1 18900
box -100 -9150 12100 25300
use POB8  Y_4
timestamp 1569139307
transform 1 0 102500 0 1 18900
box -100 -9150 12100 25300
use POB8  Y_5
timestamp 1569139307
transform 1 0 62000 0 1 18900
box -100 -9150 12100 25300
use POB8  Y_6
timestamp 1569139307
transform 1 0 116000 0 1 18900
box -100 -9150 12100 25300
use POB8  Y_7
timestamp 1569139307
transform 1 0 129500 0 1 18900
box -100 -9150 12100 25300
use PVSS  GND ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 129500 0 -1 171100
box 0 -9150 12000 25300
use PVDD  VDD ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 48500 0 1 18900
box 0 -9150 12000 25300
use MY_LOGO  MY_LOGO_0
timestamp 1756367991
transform 1 0 -610 0 1 -230
box 152200 14900 178300 173120
<< end >>