magic
tech scmos
magscale 1 30
timestamp 1727178187
<< checkpaint >>
rect 18300 186927 44800 197000
rect 13915 181835 44800 186927
rect 46919 186419 142100 190000
rect 46919 181835 143266 186419
rect 6771 176042 185015 181835
rect 6771 175958 328570 176042
rect 205 167042 328570 175958
rect 205 160774 185015 167042
rect 6771 143081 185015 160774
rect 0 142100 185015 143081
rect 0 102896 190000 142100
rect -13866 102380 190000 102896
rect -25613 89180 190000 102380
rect -24170 89077 190000 89180
rect -17472 83925 190000 89077
rect 0 47900 190000 83925
rect 6771 46919 190000 47900
rect 6771 32547 185015 46919
rect 6771 31724 186496 32547
rect -4457 10781 186496 31724
rect -4457 8670 185015 10781
rect -4457 7765 35955 8670
rect 205 1458 35955 7765
rect -600 -600 630 630
rect 46919 0 142100 8670
<< metal1 >>
rect 45400 132100 49000 138900
rect 140400 130800 144600 140200
rect 45400 51100 49000 57800
<< m2contact >>
rect 44200 132100 45400 138900
rect 144600 130800 145800 140200
rect 44200 51100 45400 57800
<< metal2 >>
rect 59800 145100 60200 145900
rect 62000 141100 62400 143900
rect 73300 141900 73700 145900
rect 86800 142500 87200 145900
rect 100300 143100 100700 145900
rect 113800 143700 114200 145900
rect 127300 143700 127700 145900
rect 100300 142800 109100 143100
rect 98000 142200 103100 142500
rect 86800 141600 94100 141900
rect 93800 141100 94100 141600
rect 102800 141100 103100 142200
rect 120100 141100 120400 142800
rect 120800 141100 121100 143400
rect 122300 141100 122600 143400
rect 140800 143100 141200 145900
rect 122900 142800 127800 143100
rect 122900 141100 123300 142800
rect 44100 132100 44200 138900
rect 145800 130800 145900 140200
rect 144300 116900 144600 118300
rect 44100 116300 46300 116700
rect 144300 116500 145900 116900
rect 46000 112100 46300 116300
rect 44100 102800 46000 103200
rect 46600 98100 46900 105700
rect 143300 103400 143600 108700
rect 143300 103000 145900 103400
rect 44100 89300 46600 89700
rect 47200 88500 47500 94800
rect 142700 89900 143000 100400
rect 142700 89500 145900 89900
rect 44100 75800 47200 76200
rect 47800 75200 48100 82500
rect 142100 76400 142400 87400
rect 142100 76000 145900 76400
rect 44100 62300 47800 62700
rect 142400 62500 145900 62900
rect 143100 59800 145900 60200
rect 51200 45400 51600 50300
rect 55100 46000 55500 50300
rect 57200 46600 57600 50400
rect 64100 47200 64500 50300
rect 78200 47800 78600 50300
rect 93800 48400 94200 50300
rect 100700 49000 101100 50300
rect 102200 49600 102600 50300
rect 102200 49300 115800 49600
rect 129300 49300 142200 49600
rect 115900 48700 127400 49000
rect 102800 48100 114100 48400
rect 78200 47500 94900 47800
rect 64100 46900 73100 47200
rect 57200 46300 64600 46600
rect 49000 45100 51600 45400
rect 49000 44100 49400 45100
rect 62500 44100 62900 45700
rect 76000 44100 76400 46300
rect 89500 44100 89900 46900
rect 113800 44100 114200 47500
rect 127300 44100 127700 48100
rect 140800 44100 141200 48700
<< m3contact >>
rect 59800 144300 60200 145100
rect 62000 143900 62400 144700
rect 113800 143400 114700 143700
rect 120200 143400 121100 143700
rect 109100 142800 110000 143100
rect 119500 142800 120400 143100
rect 86800 142200 87700 142500
rect 97100 142200 98000 142500
rect 73300 141600 74200 141900
rect 85900 141600 86800 141900
rect 122300 143400 123200 143700
rect 126800 143400 127700 143700
rect 127800 142800 128700 143100
rect 140300 142800 141200 143100
rect 144300 118300 144600 119200
rect 46000 111200 46300 112100
rect 143300 108700 143600 109600
rect 46600 105700 46900 106600
rect 46000 102800 46300 103700
rect 46600 97200 46900 98100
rect 142700 100400 143000 101300
rect 47200 94800 47500 95700
rect 46600 89300 46900 90200
rect 47200 87600 47500 88500
rect 142100 87400 142400 88300
rect 47800 82500 48100 83400
rect 47200 75800 47500 76700
rect 47800 74300 48100 75200
rect 47800 62300 48100 63200
rect 142100 61900 142400 62900
rect 142800 59300 143100 60200
rect 115800 49300 116700 49600
rect 128400 49300 129300 49600
rect 142200 49300 143100 49600
rect 100700 48700 101600 49000
rect 115000 48700 115900 49000
rect 127400 48700 128300 49000
rect 140300 48700 141200 49000
rect 93800 48100 94700 48400
rect 101900 48100 102800 48400
rect 114100 48100 115000 48400
rect 126800 48100 127700 48400
rect 94900 47500 95800 47800
rect 113300 47500 114200 47800
rect 73100 46900 74000 47200
rect 89000 46900 89900 47200
rect 64600 46300 65500 46600
rect 75500 46300 76400 46600
rect 55100 45700 56000 46000
rect 62000 45700 62900 46000
<< metal3 >>
rect 60200 144300 62000 144700
rect 114700 143400 120200 143700
rect 123200 143400 126800 143700
rect 110000 142800 119500 143100
rect 128700 142800 140300 143100
rect 87700 142200 97100 142500
rect 74200 141600 85900 141900
rect 140100 118800 144300 119200
rect 140100 115200 143600 115600
rect 46000 108700 46300 111200
rect 140100 111000 143000 111300
rect 46000 108300 49600 108700
rect 46000 107600 49600 108000
rect 46000 103700 46300 107600
rect 46900 106200 49600 106600
rect 142700 101300 143000 111000
rect 143300 109600 143600 115200
rect 140100 99300 142400 99600
rect 46600 90200 46900 97200
rect 47500 95300 49600 95700
rect 47200 76700 47500 87600
rect 142100 88300 142400 99300
rect 48100 83000 49600 83400
rect 47800 63200 48100 74300
rect 142100 56700 142400 61900
rect 140100 56400 142400 56700
rect 142800 49600 143100 59300
rect 116700 49300 128400 49600
rect 101600 48700 115000 49000
rect 128300 48700 140300 49000
rect 94700 48100 101900 48400
rect 115000 48100 126800 48400
rect 95800 47500 113300 47800
rect 74000 46900 89000 47200
rect 65500 46300 75500 46600
rect 56000 45700 62000 46000
use PIC  CIN_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1555589239
transform 1 0 62000 0 -1 171100
box -100 -9150 12100 25300
use PIC  CIN_1
timestamp 1555589239
transform 1 0 75500 0 -1 171100
box -100 -9150 12100 25300
use PIC  CIN_2
timestamp 1555589239
transform 1 0 89000 0 -1 171100
box -100 -9150 12100 25300
use PIC  CIN_3
timestamp 1555589239
transform 1 0 102500 0 -1 171100
box -100 -9150 12100 25300
use PIC  CIN_4
timestamp 1555589239
transform 1 0 116000 0 -1 171100
box -100 -9150 12100 25300
use PIC  CIN_5
timestamp 1555589239
transform 1 0 129500 0 -1 171100
box -100 -9150 12100 25300
use PIC  CLK
timestamp 1555589239
transform 1 0 48500 0 -1 171100
box -100 -9150 12100 25300
use fir_pe_Core  fir_pe_Core_0
timestamp 1727167961
transform 1 0 49845 0 1 50560
box -945 -360 90645 90660
use IOFILLER18  IOFILLER18_0 ~/ETRI050_DesignKit/pads_ETRI050
timestamp 1725930584
transform 0 -1 171100 -1 0 75646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_1
timestamp 1725930584
transform 0 -1 171098 -1 0 62146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_2
timestamp 1725930584
transform 0 -1 171100 -1 0 102646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_3
timestamp 1725930584
transform 0 -1 171100 -1 0 89146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_4
timestamp 1725930584
transform 0 -1 171102 -1 0 129646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_5
timestamp 1725930584
transform 0 -1 171100 -1 0 116146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_6
timestamp 1725930584
transform 1 0 73845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_7
timestamp 1725930584
transform 1 0 60345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_8
timestamp 1725930584
transform 1 0 100845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_9
timestamp 1725930584
transform 1 0 87345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_10
timestamp 1725930584
transform 1 0 127845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_11
timestamp 1725930584
transform 1 0 114345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_12
timestamp 1725930584
transform 0 1 18899 -1 0 75655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_13
timestamp 1725930584
transform 0 1 18899 -1 0 62155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_14
timestamp 1725930584
transform 0 1 18900 -1 0 102655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_15
timestamp 1725930584
transform 0 1 18900 -1 0 89155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_16
timestamp 1725930584
transform 1 0 73845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_17
timestamp 1725930584
transform 0 1 18897 -1 0 116155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_18
timestamp 1725930584
transform 0 1 18900 -1 0 129655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_19
timestamp 1725930584
transform 1 0 60345 0 -1 171101
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_20
timestamp 1725930584
transform 1 0 100845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_21
timestamp 1725930584
transform 1 0 87344 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_22
timestamp 1725930584
transform 1 0 127845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_23
timestamp 1725930584
transform 1 0 114345 0 -1 171100
box -60 0 1860 25060
use IOFILLER50  IOFILLER50_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1555589239
transform 1 0 43621 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_1
timestamp 1555589239
transform 1 0 141360 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_2
timestamp 1555589239
transform 1 0 141345 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_3
timestamp 1555589239
transform 1 0 43638 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_4
timestamp 1555589239
transform 0 1 18900 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_5
timestamp 1555589239
transform 0 1 18900 -1 0 146379
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_6
timestamp 1555589239
transform 0 -1 171100 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_7
timestamp 1555589239
transform 0 -1 171100 -1 0 146346
box -35 0 5035 25060
use MY_LOGO  MY_LOGO_0
timestamp 1724157349
transform 1 0 149420 0 1 9675
box 180 225 21510 9045
use PCORNER  PCORNER_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1555589239
transform 1 0 18900 0 1 18900
box 0 0 25300 25300
use PCORNER  PCORNER_1
timestamp 1555589239
transform 1 0 18900 0 -1 171100
box 0 0 25300 25300
use PCORNER  PCORNER_2
timestamp 1555589239
transform 0 -1 171100 1 0 18900
box 0 0 25300 25300
use PCORNER  PCORNER_3
timestamp 1555589239
transform -1 0 171100 0 -1 171100
box 0 0 25300 25300
use PIC  RDY_I
timestamp 1555589239
transform 0 1 18900 -1 0 74000
box -100 -9150 12100 25300
use PVDD  VDD_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1555589239
transform 0 1 18900 -1 0 141500
box -100 -9150 12100 25300
use PVDD  VDD_1
timestamp 1555589239
transform 0 1 18900 -1 0 60500
box -100 -9150 12100 25300
use POB8  VLD_O ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1555589239
transform 0 -1 171100 1 0 62000
box -100 -9150 12100 25300
use PVSS  VSS_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1555589239
transform 0 -1 171100 1 0 129500
box -100 -9150 12100 25300
use PIC  XIN_0
timestamp 1555589239
transform 0 1 18900 -1 0 87500
box -100 -9150 12100 25300
use PIC  XIN_1
timestamp 1555589239
transform 0 1 18900 -1 0 101000
box -100 -9150 12100 25300
use PIC  XIN_2
timestamp 1555589239
transform 0 1 18900 -1 0 114500
box -100 -9150 12100 25300
use PIC  XIN_3
timestamp 1555589239
transform 0 1 18900 -1 0 128000
box -100 -9150 12100 25300
use POB8  XOUT_0
timestamp 1555589239
transform 0 -1 171100 1 0 75500
box -100 -9150 12100 25300
use POB8  XOUT_1
timestamp 1555589239
transform 0 -1 171100 1 0 89000
box -100 -9150 12100 25300
use POB8  XOUT_2
timestamp 1555589239
transform 0 -1 171100 1 0 102500
box -100 -9150 12100 25300
use POB8  XOUT_3
timestamp 1555589239
transform 0 -1 171100 1 0 116000
box -100 -9150 12100 25300
use PIC  YIN_0
timestamp 1555589239
transform 0 -1 171100 1 0 48500
box -100 -9150 12100 25300
use PIC  YIN_1
timestamp 1555589239
transform 1 0 129500 0 1 18900
box -100 -9150 12100 25300
use PIC  YIN_2
timestamp 1555589239
transform 1 0 116000 0 1 18900
box -100 -9150 12100 25300
use PIC  YIN_3
timestamp 1555589239
transform 1 0 102500 0 1 18900
box -100 -9150 12100 25300
use POB8  YOUT_0
timestamp 1555589239
transform 1 0 89000 0 1 18900
box -100 -9150 12100 25300
use POB8  YOUT_1
timestamp 1555589239
transform 1 0 75500 0 1 18900
box -100 -9150 12100 25300
use POB8  YOUT_2
timestamp 1555589239
transform 1 0 62000 0 1 18900
box -100 -9150 12100 25300
use POB8  YOUT_3
timestamp 1555589239
transform 1 0 48500 0 1 18900
box -100 -9150 12100 25300
<< end >>
