magic
tech scmos
timestamp 1701862152
<< checkpaint >>
rect -7 81 37 89
rect -7 49 57 81
rect 13 40 57 49
rect 73 29 117 69
rect 163 40 237 81
<< nwell >>
rect -6 97 237 136
<< ntransistor >>
rect 12 7 14 27
rect 18 7 20 27
rect 30 7 32 27
rect 36 7 38 27
rect 61 7 63 17
rect 71 7 73 17
rect 81 7 83 17
rect 106 7 108 17
rect 116 7 118 17
rect 136 7 138 17
rect 146 7 148 17
rect 171 7 173 27
rect 177 7 179 27
rect 188 7 190 27
rect 194 7 196 27
rect 217 7 219 17
<< ptransistor >>
rect 11 103 13 123
rect 21 103 23 123
rect 31 103 33 123
rect 41 103 43 123
rect 63 113 65 123
rect 73 113 75 123
rect 83 103 85 123
rect 106 103 108 123
rect 116 103 118 123
rect 136 113 138 123
rect 146 113 148 123
rect 166 103 168 123
rect 176 103 178 123
rect 186 103 188 123
rect 196 103 198 123
rect 217 103 219 123
<< ndiffusion >>
rect 10 7 12 27
rect 14 7 18 27
rect 20 7 22 27
rect 28 7 30 27
rect 32 7 36 27
rect 38 7 40 27
rect 60 7 61 17
rect 63 7 64 17
rect 70 7 71 17
rect 73 7 74 17
rect 80 7 81 17
rect 83 7 84 17
rect 105 7 106 17
rect 108 7 109 17
rect 115 7 116 17
rect 118 7 119 17
rect 135 7 136 17
rect 138 7 139 17
rect 145 7 146 17
rect 148 7 149 17
rect 169 7 171 27
rect 173 7 177 27
rect 179 7 180 27
rect 186 7 188 27
rect 190 7 194 27
rect 196 7 198 27
rect 216 7 217 17
rect 219 7 220 17
<< pdiffusion >>
rect 10 103 11 123
rect 13 103 14 123
rect 20 103 21 123
rect 23 103 24 123
rect 30 103 31 123
rect 33 103 34 123
rect 40 103 41 123
rect 43 103 44 123
rect 62 113 63 123
rect 65 113 66 123
rect 72 113 73 123
rect 75 113 76 123
rect 82 103 83 123
rect 85 103 86 123
rect 105 103 106 123
rect 108 103 109 123
rect 115 103 116 123
rect 118 103 119 123
rect 135 113 136 123
rect 138 113 139 123
rect 145 113 146 123
rect 148 113 149 123
rect 165 103 166 123
rect 168 103 169 123
rect 175 103 176 123
rect 178 103 179 123
rect 185 103 186 123
rect 188 103 189 123
rect 195 103 196 123
rect 198 103 199 123
rect 216 103 217 123
rect 219 103 220 123
<< ndcontact >>
rect 4 7 10 27
rect 22 7 28 27
rect 40 7 46 27
rect 54 7 60 17
rect 64 7 70 17
rect 74 7 80 17
rect 84 7 90 17
rect 99 7 105 17
rect 109 7 115 17
rect 119 7 125 17
rect 129 7 135 17
rect 139 7 145 17
rect 149 7 155 17
rect 163 7 169 27
rect 180 7 186 27
rect 198 7 204 27
rect 210 7 216 17
rect 220 7 226 17
<< pdcontact >>
rect 4 103 10 123
rect 14 103 20 123
rect 24 103 30 123
rect 34 103 40 123
rect 44 103 50 123
rect 56 113 62 123
rect 66 113 72 123
rect 76 103 82 123
rect 86 103 92 123
rect 99 103 105 123
rect 109 103 115 123
rect 119 103 125 123
rect 129 113 135 123
rect 139 113 145 123
rect 149 113 155 123
rect 159 103 165 123
rect 169 103 175 123
rect 179 103 185 123
rect 189 103 195 123
rect 199 103 205 123
rect 210 103 216 123
rect 220 103 226 123
<< psubstratepcontact >>
rect -3 -3 233 3
<< nsubstratencontact >>
rect -3 127 233 133
<< polysilicon >>
rect 11 123 13 125
rect 21 123 23 125
rect 31 123 33 125
rect 41 123 43 125
rect 63 123 65 125
rect 73 123 75 125
rect 83 123 85 125
rect 106 123 108 125
rect 116 123 118 125
rect 136 123 138 125
rect 146 123 148 125
rect 166 123 168 125
rect 176 123 178 125
rect 186 123 188 125
rect 196 123 198 125
rect 217 123 219 125
rect 11 58 13 103
rect 21 94 23 103
rect 11 52 12 58
rect 12 27 14 52
rect 22 36 24 88
rect 31 86 33 103
rect 18 27 20 30
rect 30 27 32 80
rect 41 68 43 103
rect 41 42 43 62
rect 63 49 65 113
rect 73 66 75 113
rect 36 40 43 42
rect 36 27 38 40
rect 73 39 75 60
rect 83 45 85 103
rect 106 71 108 103
rect 116 83 118 103
rect 136 96 138 113
rect 128 90 138 96
rect 116 80 130 83
rect 106 66 115 71
rect 61 37 75 39
rect 61 17 63 37
rect 71 17 73 27
rect 81 17 83 39
rect 106 27 108 66
rect 128 58 130 80
rect 116 56 130 58
rect 116 40 118 56
rect 136 55 138 90
rect 146 72 148 113
rect 166 97 168 103
rect 148 66 155 69
rect 136 52 148 55
rect 93 23 108 27
rect 106 17 108 23
rect 116 17 118 34
rect 136 17 138 27
rect 146 17 148 52
rect 152 33 155 66
rect 160 42 163 94
rect 176 83 178 103
rect 186 95 188 103
rect 168 80 178 83
rect 168 67 171 80
rect 186 75 188 89
rect 196 80 198 103
rect 181 72 188 75
rect 160 39 165 42
rect 162 30 165 39
rect 168 34 171 61
rect 181 44 183 72
rect 196 51 198 74
rect 182 38 183 44
rect 168 32 179 34
rect 162 28 173 30
rect 171 27 173 28
rect 177 27 179 32
rect 181 30 183 38
rect 186 48 198 51
rect 186 34 188 48
rect 217 44 219 103
rect 198 38 219 44
rect 186 32 196 34
rect 181 28 190 30
rect 188 27 190 28
rect 194 27 196 32
rect 217 17 219 38
rect 12 5 14 7
rect 18 5 20 7
rect 30 5 32 7
rect 36 5 38 7
rect 61 5 63 7
rect 71 5 73 7
rect 81 5 83 7
rect 106 5 108 7
rect 116 5 118 7
rect 136 5 138 7
rect 146 5 148 7
rect 171 5 173 7
rect 177 5 179 7
rect 188 5 190 7
rect 194 5 196 7
rect 217 5 219 7
<< polycontact >>
rect 19 88 25 94
rect 12 52 18 58
rect 18 30 24 36
rect 30 80 36 86
rect 38 62 44 68
rect 73 60 79 66
rect 63 43 69 49
rect 122 90 128 96
rect 81 39 87 45
rect 71 27 77 33
rect 115 65 121 71
rect 142 66 148 72
rect 160 94 166 100
rect 112 34 118 40
rect 87 20 93 27
rect 136 27 142 33
rect 182 89 188 95
rect 192 74 198 80
rect 168 61 174 67
rect 152 27 158 33
rect 176 38 182 44
rect 192 38 198 44
<< metal1 >>
rect -3 133 233 134
rect -3 126 233 127
rect 4 123 10 126
rect 24 123 30 126
rect 44 123 50 126
rect 86 123 92 126
rect 109 123 115 126
rect 159 123 165 126
rect 179 123 185 126
rect 199 123 205 126
rect 220 123 226 126
rect 13 103 14 106
rect 13 100 16 103
rect 4 97 16 100
rect 4 43 8 97
rect 34 93 40 103
rect 99 98 105 103
rect 25 89 83 93
rect 99 91 103 98
rect 119 96 121 103
rect 146 96 160 100
rect 119 90 122 96
rect 169 93 173 103
rect 191 100 195 103
rect 191 97 204 100
rect 79 87 83 89
rect 36 80 63 84
rect 79 83 131 87
rect 169 89 182 93
rect 201 86 204 97
rect 156 83 204 86
rect 79 76 192 80
rect 79 74 83 76
rect 38 71 83 74
rect 38 68 44 71
rect 12 58 18 61
rect 79 62 103 66
rect 145 62 148 66
rect 103 59 148 62
rect 157 61 168 67
rect 157 56 160 61
rect 18 52 160 56
rect 181 52 186 61
rect 4 39 53 43
rect 4 27 8 39
rect 24 30 46 34
rect 41 27 46 30
rect 63 33 66 43
rect 87 42 91 45
rect 164 47 186 52
rect 119 42 169 47
rect 172 38 176 44
rect 182 38 192 44
rect 63 29 71 33
rect 77 29 87 33
rect 84 23 87 29
rect 142 27 152 33
rect 172 27 177 38
rect 201 27 204 83
rect 99 20 101 27
rect 99 17 105 20
rect 169 23 177 27
rect 210 68 215 103
rect 210 61 211 68
rect 210 17 215 61
rect 22 4 28 7
rect 84 4 90 7
rect 109 4 115 7
rect 180 4 186 7
rect 220 4 226 7
rect -3 3 233 4
rect -3 -4 233 -3
<< m2contact >>
rect 56 106 63 113
rect 66 106 73 113
rect 129 106 136 113
rect 139 106 146 113
rect 149 106 156 113
rect 74 96 81 103
rect 103 91 110 98
rect 121 96 128 103
rect 139 96 146 103
rect 63 79 70 86
rect 131 83 138 90
rect 149 83 156 90
rect 11 61 18 68
rect 31 61 38 68
rect 103 62 110 69
rect 121 65 128 72
rect 181 61 188 68
rect 53 36 60 43
rect 91 41 98 48
rect 112 40 119 47
rect 54 17 61 24
rect 64 17 71 24
rect 74 17 81 24
rect 101 20 108 27
rect 119 17 126 24
rect 129 17 136 24
rect 139 17 146 24
rect 149 17 156 24
rect 211 61 218 68
<< metal2 >>
rect 53 106 56 113
rect 13 68 17 77
rect 33 53 37 61
rect 53 43 58 106
rect 66 86 70 106
rect 56 24 60 36
rect 66 24 70 79
rect 74 24 78 96
rect 103 69 106 91
rect 122 72 126 96
rect 131 90 136 106
rect 139 103 146 106
rect 93 48 97 57
rect 103 27 106 62
rect 122 24 126 65
rect 131 24 136 83
rect 142 24 146 96
rect 149 90 154 106
rect 149 24 154 83
rect 183 53 187 61
rect 213 53 217 61
<< m1p >>
rect -3 126 233 134
rect -3 -4 233 4
<< m2p >>
rect 13 69 17 77
rect 33 53 37 60
rect 93 49 97 57
rect 183 53 187 60
rect 213 53 217 60
<< labels >>
rlabel metal2 94 56 94 56 1 D
port 1 n signal input
rlabel metal2 35 54 35 54 7 S
port 2 n signal input
rlabel metal2 15 76 15 76 1 R
port 3 n signal input
rlabel metal2 185 54 185 54 3 CLK
port 4 n signal input
rlabel metal2 215 54 215 54 1 Q
port 5 n signal output
rlabel metal1 -3 126 233 134 0 vdd
port 6 nsew power bidirectional abutment
rlabel metal1 -3 -4 233 4 0 gnd
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 230 130
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
