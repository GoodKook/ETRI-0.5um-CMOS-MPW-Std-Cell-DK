magic
tech scmos
magscale 1 2
timestamp 1702307569
<< nwell >>
rect -13 154 93 272
<< ntransistor >>
rect 18 14 22 54
rect 38 14 42 54
rect 58 14 62 54
<< ptransistor >>
rect 21 166 25 246
rect 35 166 39 246
rect 55 206 59 246
<< ndiffusion >>
rect 16 14 18 54
rect 22 45 38 54
rect 22 14 24 45
rect 36 14 38 45
rect 42 14 44 54
rect 56 14 58 54
rect 62 14 64 54
<< pdiffusion >>
rect 19 166 21 246
rect 25 166 35 246
rect 39 166 41 246
rect 53 206 55 246
rect 59 206 61 246
<< ndcontact >>
rect 4 14 16 54
rect 24 14 36 45
rect 44 14 56 54
rect 64 14 76 54
<< pdcontact >>
rect 7 166 19 246
rect 41 166 53 246
rect 61 206 73 246
<< psubstratepcontact >>
rect -7 -6 87 6
<< nsubstratencontact >>
rect -7 254 87 266
<< polysilicon >>
rect 21 246 25 250
rect 35 246 39 250
rect 55 246 59 250
rect 55 190 59 206
rect 55 184 62 190
rect 21 164 25 166
rect 15 160 25 164
rect 35 164 39 166
rect 35 160 42 164
rect 15 117 19 160
rect 17 105 19 117
rect 15 68 19 105
rect 38 97 42 160
rect 39 85 42 97
rect 15 64 22 68
rect 18 54 22 64
rect 38 54 42 85
rect 58 97 62 184
rect 58 85 63 97
rect 58 54 62 85
rect 18 10 22 14
rect 38 10 42 14
rect 58 10 62 14
<< polycontact >>
rect 5 105 17 117
rect 27 85 39 97
rect 63 85 75 97
<< metal1 >>
rect -7 266 87 268
rect -7 252 87 254
rect 7 246 19 252
rect 61 246 73 252
rect 53 166 54 174
rect 46 137 54 166
rect 3 123 17 137
rect 43 123 57 137
rect 5 117 17 123
rect 23 103 37 117
rect 27 97 37 103
rect 46 69 54 123
rect 63 103 77 117
rect 63 97 75 103
rect 46 63 72 69
rect 4 54 56 57
rect 16 51 44 54
rect 64 54 72 63
rect 24 8 36 14
rect -7 6 87 8
rect -7 -8 87 -6
<< m1p >>
rect -7 252 87 268
rect 3 123 17 137
rect 43 123 57 137
rect 23 103 37 117
rect 63 103 77 117
rect -7 -8 87 8
<< labels >>
rlabel nsubstratencontact 40 260 40 260 0 vdd
port 5 nsew power bidirectional abutment
rlabel psubstratepcontact 40 0 40 0 0 gnd
port 6 nsew ground bidirectional abutment
rlabel metal1 10 127 10 127 0 A
port 1 nsew signal input
rlabel metal1 50 131 50 131 0 Y
port 4 nsew signal output
rlabel metal1 30 107 30 107 0 B
port 2 nsew signal input
rlabel metal1 70 111 70 111 0 C
port 3 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 80 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
