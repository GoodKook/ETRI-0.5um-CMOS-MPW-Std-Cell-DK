magic
tech scmos
magscale 1 2
timestamp 1728305240
<< nwell >>
rect -13 134 112 252
<< ntransistor >>
rect 21 14 25 34
rect 41 14 45 34
rect 61 14 65 34
<< ptransistor >>
rect 21 146 25 226
rect 31 146 35 226
rect 53 186 57 226
<< ndiffusion >>
rect 19 14 21 34
rect 25 14 27 34
rect 39 14 41 34
rect 45 14 47 34
rect 59 14 61 34
rect 65 14 67 34
<< pdiffusion >>
rect 19 146 21 226
rect 25 146 31 226
rect 35 146 37 226
rect 49 186 53 226
rect 57 186 59 226
<< ndcontact >>
rect 7 14 19 34
rect 27 14 39 34
rect 47 14 59 34
rect 67 14 79 34
<< pdcontact >>
rect 7 146 19 226
rect 37 146 49 226
rect 59 186 71 226
<< psubstratepcontact >>
rect -7 -6 106 6
<< nsubstratencontact >>
rect -7 234 106 246
<< polysilicon >>
rect 21 226 25 230
rect 31 226 35 230
rect 53 226 57 230
rect 21 124 25 146
rect 12 118 25 124
rect 12 103 16 118
rect 12 45 16 91
rect 31 69 35 146
rect 53 140 57 186
rect 36 57 45 69
rect 12 40 25 45
rect 21 34 25 40
rect 41 34 45 57
rect 61 34 65 44
rect 21 10 25 14
rect 41 10 45 14
rect 61 10 65 14
<< polycontact >>
rect 4 91 16 103
rect 51 128 63 140
rect 24 57 36 69
rect 53 44 65 56
<< metal1 >>
rect -7 246 106 248
rect -7 232 106 234
rect 37 226 49 232
rect 59 180 77 186
rect 7 140 19 146
rect 7 134 51 140
rect 49 128 51 134
rect 49 56 57 128
rect 69 83 77 180
rect 77 69 79 83
rect 49 50 53 56
rect 29 44 53 50
rect 29 34 35 44
rect 71 34 79 69
rect 7 8 19 14
rect 47 8 59 14
rect -7 6 106 8
rect -7 -8 106 -6
<< m2contact >>
rect 3 77 17 91
rect 23 69 37 83
rect 63 69 77 83
<< metal2 >>
rect 3 63 17 77
rect 23 83 37 97
rect 63 83 77 97
<< m1p >>
rect -7 232 106 248
rect -7 -8 106 8
<< m2p >>
rect 23 83 37 97
rect 63 83 77 97
rect 3 63 17 77
<< labels >>
rlabel metal1 -7 -8 106 8 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 -7 232 106 248 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal2 3 63 17 77 0 A
port 0 nsew signal input
rlabel metal2 63 83 77 97 0 Y
port 2 nsew signal output
rlabel metal2 23 83 37 97 0 B
port 1 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
