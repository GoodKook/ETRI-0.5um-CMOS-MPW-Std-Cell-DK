magic
tech scmos
magscale 1 2
timestamp 1702508443
<< nwell >>
rect -13 154 94 272
<< ntransistor >>
rect 18 14 22 54
rect 28 14 32 54
rect 48 14 52 34
<< ptransistor >>
rect 18 206 22 246
rect 38 206 42 246
rect 58 206 62 246
<< ndiffusion >>
rect 16 14 18 54
rect 22 14 28 54
rect 32 14 34 54
rect 46 14 48 34
rect 52 14 54 34
<< pdiffusion >>
rect 16 206 18 246
rect 22 206 24 246
rect 36 206 38 246
rect 42 206 44 246
rect 56 206 58 246
rect 62 206 64 246
<< ndcontact >>
rect 4 14 16 54
rect 34 14 46 54
rect 54 14 66 34
<< pdcontact >>
rect 4 206 16 246
rect 24 206 36 246
rect 44 206 56 246
rect 64 206 76 246
<< psubstratepcontact >>
rect -6 -6 86 6
<< nsubstratencontact >>
rect -6 254 86 266
<< polysilicon >>
rect 18 246 22 250
rect 38 246 42 250
rect 58 246 62 250
rect 18 54 22 206
rect 38 129 42 206
rect 38 85 42 117
rect 28 80 42 85
rect 28 54 32 80
rect 58 72 62 206
rect 60 60 62 72
rect 48 34 52 60
rect 18 10 22 14
rect 28 10 32 14
rect 48 10 52 14
<< polycontact >>
rect 6 91 18 103
rect 38 117 50 129
rect 48 60 60 72
<< metal1 >>
rect -6 266 86 268
rect -6 252 86 254
rect 4 246 16 252
rect 44 246 56 252
rect 25 72 32 206
rect 64 117 72 206
rect 4 64 48 72
rect 4 54 16 64
rect 66 40 72 103
rect 54 34 72 40
rect 34 8 42 14
rect -6 6 86 8
rect -6 -8 86 -6
<< m2contact >>
rect 5 103 19 117
rect 40 103 54 117
rect 60 103 74 117
<< metal2 >>
rect 6 117 14 134
rect 66 117 74 134
rect 46 86 54 103
<< m1p >>
rect -6 252 86 268
rect -6 -8 86 8
<< m2p >>
rect 6 119 14 134
rect 66 119 74 134
rect 46 86 54 101
<< labels >>
rlabel metal2 10 131 10 131 1 A
port 1 n signal input
rlabel metal2 50 89 50 89 1 B
port 2 n signal input
rlabel metal2 70 131 70 131 5 Y
port 3 n signal output
rlabel metal1 -6 252 86 268 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 -6 -8 86 8 0 gnd
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 80 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
